module basic_750_5000_1000_5_levels_1xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_543,In_596);
or U1 (N_1,In_511,In_466);
and U2 (N_2,In_316,In_108);
nand U3 (N_3,In_566,In_548);
and U4 (N_4,In_186,In_154);
or U5 (N_5,In_461,In_724);
and U6 (N_6,In_609,In_103);
nand U7 (N_7,In_169,In_87);
nor U8 (N_8,In_68,In_326);
or U9 (N_9,In_202,In_734);
and U10 (N_10,In_669,In_293);
and U11 (N_11,In_612,In_7);
nor U12 (N_12,In_567,In_505);
nor U13 (N_13,In_400,In_586);
nand U14 (N_14,In_340,In_502);
nand U15 (N_15,In_294,In_83);
nand U16 (N_16,In_331,In_574);
nor U17 (N_17,In_525,In_419);
or U18 (N_18,In_638,In_9);
nand U19 (N_19,In_41,In_238);
or U20 (N_20,In_193,In_743);
and U21 (N_21,In_675,In_179);
or U22 (N_22,In_300,In_627);
and U23 (N_23,In_350,In_591);
or U24 (N_24,In_11,In_506);
and U25 (N_25,In_335,In_580);
and U26 (N_26,In_613,In_545);
and U27 (N_27,In_50,In_381);
nor U28 (N_28,In_38,In_366);
and U29 (N_29,In_386,In_618);
and U30 (N_30,In_392,In_454);
or U31 (N_31,In_464,In_82);
nand U32 (N_32,In_710,In_291);
nor U33 (N_33,In_504,In_65);
xnor U34 (N_34,In_721,In_700);
nor U35 (N_35,In_157,In_571);
and U36 (N_36,In_218,In_537);
or U37 (N_37,In_195,In_289);
nand U38 (N_38,In_29,In_64);
nor U39 (N_39,In_369,In_501);
nor U40 (N_40,In_346,In_190);
and U41 (N_41,In_465,In_557);
or U42 (N_42,In_544,In_277);
nor U43 (N_43,In_474,In_483);
and U44 (N_44,In_705,In_363);
and U45 (N_45,In_124,In_281);
nor U46 (N_46,In_744,In_244);
nor U47 (N_47,In_717,In_579);
and U48 (N_48,In_560,In_237);
nand U49 (N_49,In_211,In_128);
and U50 (N_50,In_347,In_563);
nor U51 (N_51,In_739,In_98);
and U52 (N_52,In_372,In_262);
or U53 (N_53,In_147,In_726);
nor U54 (N_54,In_480,In_46);
or U55 (N_55,In_167,In_456);
and U56 (N_56,In_549,In_684);
and U57 (N_57,In_603,In_79);
nor U58 (N_58,In_200,In_418);
nor U59 (N_59,In_655,In_679);
nor U60 (N_60,In_641,In_119);
nand U61 (N_61,In_703,In_180);
nor U62 (N_62,In_257,In_5);
or U63 (N_63,In_359,In_223);
and U64 (N_64,In_408,In_106);
and U65 (N_65,In_182,In_16);
and U66 (N_66,In_714,In_733);
nand U67 (N_67,In_707,In_630);
nor U68 (N_68,In_2,In_94);
nand U69 (N_69,In_607,In_336);
nor U70 (N_70,In_148,In_540);
nand U71 (N_71,In_220,In_28);
and U72 (N_72,In_619,In_35);
nand U73 (N_73,In_521,In_95);
nor U74 (N_74,In_694,In_330);
nand U75 (N_75,In_364,In_647);
nand U76 (N_76,In_55,In_665);
and U77 (N_77,In_159,In_469);
or U78 (N_78,In_583,In_528);
and U79 (N_79,In_181,In_531);
and U80 (N_80,In_199,In_354);
xnor U81 (N_81,In_737,In_532);
nor U82 (N_82,In_123,In_313);
or U83 (N_83,In_553,In_308);
and U84 (N_84,In_356,In_353);
nor U85 (N_85,In_404,In_284);
and U86 (N_86,In_192,In_288);
nor U87 (N_87,In_485,In_156);
nand U88 (N_88,In_617,In_219);
and U89 (N_89,In_376,In_115);
and U90 (N_90,In_341,In_213);
and U91 (N_91,In_390,In_582);
and U92 (N_92,In_215,In_541);
nand U93 (N_93,In_536,In_741);
and U94 (N_94,In_299,In_695);
nor U95 (N_95,In_547,In_559);
nand U96 (N_96,In_656,In_197);
or U97 (N_97,In_489,In_176);
or U98 (N_98,In_701,In_409);
and U99 (N_99,In_342,In_301);
or U100 (N_100,In_177,In_67);
and U101 (N_101,In_90,In_691);
or U102 (N_102,In_666,In_120);
and U103 (N_103,In_114,In_518);
and U104 (N_104,In_608,In_236);
nor U105 (N_105,In_729,In_317);
or U106 (N_106,In_440,In_351);
nor U107 (N_107,In_662,In_33);
nand U108 (N_108,In_422,In_590);
nor U109 (N_109,In_508,In_615);
or U110 (N_110,In_170,In_26);
nor U111 (N_111,In_246,In_491);
and U112 (N_112,In_189,In_252);
nor U113 (N_113,In_498,In_430);
nand U114 (N_114,In_245,In_587);
nor U115 (N_115,In_164,In_681);
or U116 (N_116,In_453,In_130);
nand U117 (N_117,In_514,In_222);
and U118 (N_118,In_628,In_85);
and U119 (N_119,In_452,In_477);
and U120 (N_120,In_746,In_602);
or U121 (N_121,In_605,In_524);
nand U122 (N_122,In_478,In_93);
and U123 (N_123,In_160,In_402);
or U124 (N_124,In_292,In_519);
nor U125 (N_125,In_611,In_125);
nor U126 (N_126,In_178,In_92);
nor U127 (N_127,In_70,In_37);
or U128 (N_128,In_713,In_371);
and U129 (N_129,In_241,In_229);
nand U130 (N_130,In_564,In_248);
nor U131 (N_131,In_463,In_389);
nand U132 (N_132,In_275,In_297);
or U133 (N_133,In_266,In_233);
nor U134 (N_134,In_486,In_459);
and U135 (N_135,In_207,In_109);
or U136 (N_136,In_450,In_370);
or U137 (N_137,In_10,In_355);
and U138 (N_138,In_306,In_327);
nor U139 (N_139,In_742,In_432);
xor U140 (N_140,In_60,In_576);
nor U141 (N_141,In_368,In_102);
and U142 (N_142,In_250,In_13);
nor U143 (N_143,In_426,In_405);
nand U144 (N_144,In_584,In_17);
nor U145 (N_145,In_460,In_614);
nand U146 (N_146,In_431,In_12);
nor U147 (N_147,In_117,In_448);
and U148 (N_148,In_442,In_45);
nand U149 (N_149,In_719,In_40);
nand U150 (N_150,In_449,In_146);
or U151 (N_151,In_290,In_558);
nor U152 (N_152,In_581,In_629);
nand U153 (N_153,In_30,In_62);
nand U154 (N_154,In_569,In_551);
or U155 (N_155,In_417,In_63);
and U156 (N_156,In_255,In_137);
nand U157 (N_157,In_577,In_185);
nand U158 (N_158,In_527,In_572);
nand U159 (N_159,In_435,In_259);
or U160 (N_160,In_247,In_84);
nor U161 (N_161,In_539,In_3);
or U162 (N_162,In_573,In_663);
and U163 (N_163,In_633,In_565);
nor U164 (N_164,In_328,In_393);
or U165 (N_165,In_401,In_142);
and U166 (N_166,In_387,In_443);
and U167 (N_167,In_507,In_692);
or U168 (N_168,In_421,In_671);
and U169 (N_169,In_664,In_151);
and U170 (N_170,In_697,In_339);
nor U171 (N_171,In_623,In_75);
nor U172 (N_172,In_499,In_451);
nor U173 (N_173,In_264,In_140);
and U174 (N_174,In_53,In_490);
and U175 (N_175,In_513,In_231);
and U176 (N_176,In_526,In_338);
or U177 (N_177,In_112,In_155);
and U178 (N_178,In_333,In_319);
nor U179 (N_179,In_228,In_735);
nand U180 (N_180,In_141,In_731);
nand U181 (N_181,In_672,In_162);
nand U182 (N_182,In_696,In_682);
or U183 (N_183,In_429,In_598);
nor U184 (N_184,In_323,In_533);
nor U185 (N_185,In_658,In_274);
and U186 (N_186,In_661,In_172);
and U187 (N_187,In_174,In_4);
nor U188 (N_188,In_626,In_8);
nor U189 (N_189,In_104,In_126);
nand U190 (N_190,In_171,In_352);
and U191 (N_191,In_686,In_362);
nand U192 (N_192,In_745,In_258);
and U193 (N_193,In_272,In_471);
and U194 (N_194,In_221,In_99);
or U195 (N_195,In_747,In_588);
and U196 (N_196,In_161,In_723);
nor U197 (N_197,In_510,In_711);
nor U198 (N_198,In_382,In_110);
nand U199 (N_199,In_594,In_648);
and U200 (N_200,In_708,In_1);
and U201 (N_201,In_455,In_34);
nand U202 (N_202,In_73,In_496);
nand U203 (N_203,In_205,In_413);
nand U204 (N_204,In_6,In_42);
or U205 (N_205,In_309,In_101);
and U206 (N_206,In_621,In_216);
nand U207 (N_207,In_677,In_96);
nor U208 (N_208,In_652,In_302);
and U209 (N_209,In_78,In_14);
and U210 (N_210,In_670,In_585);
or U211 (N_211,In_194,In_307);
and U212 (N_212,In_374,In_253);
nor U213 (N_213,In_706,In_484);
and U214 (N_214,In_260,In_391);
nor U215 (N_215,In_168,In_689);
nor U216 (N_216,In_270,In_481);
or U217 (N_217,In_667,In_654);
nand U218 (N_218,In_204,In_242);
nand U219 (N_219,In_561,In_482);
nand U220 (N_220,In_235,In_116);
or U221 (N_221,In_562,In_720);
nor U222 (N_222,In_441,In_278);
and U223 (N_223,In_97,In_622);
or U224 (N_224,In_135,In_226);
and U225 (N_225,In_145,In_578);
and U226 (N_226,In_304,In_312);
nand U227 (N_227,In_439,In_427);
or U228 (N_228,In_196,In_153);
or U229 (N_229,In_227,In_487);
and U230 (N_230,In_552,In_152);
and U231 (N_231,In_494,In_314);
nor U232 (N_232,In_129,In_320);
and U233 (N_233,In_332,In_467);
and U234 (N_234,In_298,In_715);
or U235 (N_235,In_380,In_678);
nand U236 (N_236,In_311,In_133);
or U237 (N_237,In_415,In_377);
and U238 (N_238,In_113,In_604);
nor U239 (N_239,In_163,In_636);
or U240 (N_240,In_606,In_384);
nor U241 (N_241,In_39,In_420);
xor U242 (N_242,In_416,In_592);
nand U243 (N_243,In_296,In_433);
nand U244 (N_244,In_509,In_631);
nor U245 (N_245,In_361,In_49);
and U246 (N_246,In_653,In_388);
or U247 (N_247,In_76,In_249);
nor U248 (N_248,In_517,In_27);
nand U249 (N_249,In_497,In_411);
nand U250 (N_250,In_166,In_428);
or U251 (N_251,In_91,In_295);
and U252 (N_252,In_61,In_303);
and U253 (N_253,In_645,In_625);
and U254 (N_254,In_639,In_105);
nor U255 (N_255,In_680,In_51);
and U256 (N_256,In_424,In_118);
nand U257 (N_257,In_365,In_512);
nor U258 (N_258,In_712,In_243);
nand U259 (N_259,In_357,In_144);
nor U260 (N_260,In_240,In_378);
and U261 (N_261,In_36,In_121);
nand U262 (N_262,In_86,In_685);
or U263 (N_263,In_520,In_651);
and U264 (N_264,In_25,In_704);
and U265 (N_265,In_412,In_403);
nor U266 (N_266,In_688,In_214);
nor U267 (N_267,In_395,In_728);
nor U268 (N_268,In_748,In_457);
nor U269 (N_269,In_425,In_740);
or U270 (N_270,In_345,In_473);
nor U271 (N_271,In_699,In_472);
or U272 (N_272,In_550,In_149);
nor U273 (N_273,In_632,In_610);
or U274 (N_274,In_225,In_337);
nand U275 (N_275,In_122,In_568);
nor U276 (N_276,In_165,In_646);
or U277 (N_277,In_89,In_265);
or U278 (N_278,In_158,In_71);
nor U279 (N_279,In_535,In_283);
and U280 (N_280,In_276,In_522);
or U281 (N_281,In_749,In_725);
and U282 (N_282,In_285,In_324);
nand U283 (N_283,In_635,In_210);
nand U284 (N_284,In_479,In_212);
nand U285 (N_285,In_251,In_399);
nor U286 (N_286,In_143,In_282);
nand U287 (N_287,In_254,In_191);
or U288 (N_288,In_690,In_209);
nor U289 (N_289,In_150,In_538);
or U290 (N_290,In_279,In_492);
nand U291 (N_291,In_234,In_59);
and U292 (N_292,In_423,In_136);
and U293 (N_293,In_595,In_616);
nor U294 (N_294,In_659,In_325);
or U295 (N_295,In_15,In_444);
or U296 (N_296,In_643,In_406);
and U297 (N_297,In_256,In_657);
nor U298 (N_298,In_673,In_738);
nand U299 (N_299,In_718,In_730);
or U300 (N_300,In_642,In_396);
and U301 (N_301,In_74,In_206);
xor U302 (N_302,In_201,In_599);
xnor U303 (N_303,In_687,In_488);
or U304 (N_304,In_650,In_458);
and U305 (N_305,In_318,In_72);
nand U306 (N_306,In_601,In_556);
nand U307 (N_307,In_321,In_732);
and U308 (N_308,In_263,In_575);
or U309 (N_309,In_230,In_20);
or U310 (N_310,In_57,In_52);
or U311 (N_311,In_593,In_397);
and U312 (N_312,In_269,In_305);
and U313 (N_313,In_208,In_437);
nor U314 (N_314,In_56,In_69);
nand U315 (N_315,In_407,In_77);
and U316 (N_316,In_445,In_224);
or U317 (N_317,In_446,In_683);
or U318 (N_318,In_100,In_175);
and U319 (N_319,In_19,In_127);
or U320 (N_320,In_398,In_271);
and U321 (N_321,In_81,In_358);
nand U322 (N_322,In_523,In_436);
or U323 (N_323,In_310,In_198);
or U324 (N_324,In_88,In_470);
nor U325 (N_325,In_649,In_637);
nor U326 (N_326,In_24,In_394);
nor U327 (N_327,In_58,In_500);
and U328 (N_328,In_280,In_203);
nor U329 (N_329,In_698,In_373);
and U330 (N_330,In_173,In_529);
nand U331 (N_331,In_385,In_131);
or U332 (N_332,In_139,In_468);
or U333 (N_333,In_554,In_43);
and U334 (N_334,In_640,In_379);
or U335 (N_335,In_383,In_286);
nand U336 (N_336,In_48,In_660);
nor U337 (N_337,In_709,In_447);
nor U338 (N_338,In_349,In_438);
nor U339 (N_339,In_476,In_66);
nor U340 (N_340,In_267,In_21);
nor U341 (N_341,In_516,In_54);
nor U342 (N_342,In_530,In_736);
nand U343 (N_343,In_570,In_367);
or U344 (N_344,In_555,In_32);
and U345 (N_345,In_111,In_727);
nor U346 (N_346,In_503,In_702);
and U347 (N_347,In_273,In_360);
or U348 (N_348,In_495,In_22);
or U349 (N_349,In_676,In_315);
nand U350 (N_350,In_674,In_31);
and U351 (N_351,In_107,In_344);
nand U352 (N_352,In_475,In_329);
nand U353 (N_353,In_348,In_620);
nand U354 (N_354,In_322,In_597);
nor U355 (N_355,In_624,In_343);
nand U356 (N_356,In_80,In_493);
nor U357 (N_357,In_261,In_334);
nand U358 (N_358,In_589,In_722);
nor U359 (N_359,In_668,In_434);
or U360 (N_360,In_183,In_184);
nand U361 (N_361,In_138,In_47);
nand U362 (N_362,In_188,In_287);
and U363 (N_363,In_23,In_134);
nand U364 (N_364,In_217,In_132);
nand U365 (N_365,In_0,In_410);
nor U366 (N_366,In_239,In_644);
or U367 (N_367,In_542,In_268);
nand U368 (N_368,In_534,In_716);
nand U369 (N_369,In_187,In_515);
nor U370 (N_370,In_634,In_414);
and U371 (N_371,In_44,In_462);
and U372 (N_372,In_375,In_18);
or U373 (N_373,In_600,In_693);
nor U374 (N_374,In_546,In_232);
and U375 (N_375,In_329,In_123);
nor U376 (N_376,In_742,In_567);
or U377 (N_377,In_344,In_52);
or U378 (N_378,In_339,In_39);
and U379 (N_379,In_0,In_504);
or U380 (N_380,In_685,In_125);
xor U381 (N_381,In_492,In_46);
and U382 (N_382,In_101,In_328);
nor U383 (N_383,In_258,In_321);
nor U384 (N_384,In_81,In_207);
or U385 (N_385,In_264,In_571);
nor U386 (N_386,In_149,In_42);
and U387 (N_387,In_309,In_728);
or U388 (N_388,In_450,In_81);
or U389 (N_389,In_399,In_662);
nor U390 (N_390,In_133,In_302);
nand U391 (N_391,In_461,In_537);
and U392 (N_392,In_317,In_601);
nand U393 (N_393,In_284,In_143);
nand U394 (N_394,In_211,In_226);
or U395 (N_395,In_262,In_73);
nand U396 (N_396,In_468,In_503);
xor U397 (N_397,In_454,In_564);
and U398 (N_398,In_595,In_96);
and U399 (N_399,In_404,In_162);
nand U400 (N_400,In_237,In_243);
nor U401 (N_401,In_593,In_441);
or U402 (N_402,In_23,In_536);
nand U403 (N_403,In_151,In_734);
nand U404 (N_404,In_430,In_120);
nor U405 (N_405,In_314,In_675);
nand U406 (N_406,In_195,In_581);
and U407 (N_407,In_562,In_206);
nand U408 (N_408,In_593,In_391);
nand U409 (N_409,In_207,In_252);
nand U410 (N_410,In_313,In_154);
nand U411 (N_411,In_497,In_744);
and U412 (N_412,In_716,In_582);
nand U413 (N_413,In_347,In_618);
nand U414 (N_414,In_523,In_399);
and U415 (N_415,In_234,In_632);
nor U416 (N_416,In_120,In_83);
and U417 (N_417,In_78,In_136);
and U418 (N_418,In_395,In_393);
nor U419 (N_419,In_107,In_174);
and U420 (N_420,In_507,In_2);
or U421 (N_421,In_515,In_474);
nand U422 (N_422,In_531,In_346);
or U423 (N_423,In_480,In_563);
or U424 (N_424,In_85,In_156);
or U425 (N_425,In_206,In_8);
nor U426 (N_426,In_15,In_49);
and U427 (N_427,In_381,In_667);
or U428 (N_428,In_581,In_21);
and U429 (N_429,In_712,In_308);
and U430 (N_430,In_449,In_424);
nor U431 (N_431,In_368,In_588);
nor U432 (N_432,In_653,In_379);
nor U433 (N_433,In_370,In_600);
and U434 (N_434,In_375,In_21);
nor U435 (N_435,In_277,In_173);
nand U436 (N_436,In_569,In_573);
nand U437 (N_437,In_293,In_383);
nand U438 (N_438,In_719,In_351);
and U439 (N_439,In_64,In_300);
and U440 (N_440,In_591,In_143);
nand U441 (N_441,In_548,In_142);
nand U442 (N_442,In_515,In_217);
nor U443 (N_443,In_396,In_300);
nor U444 (N_444,In_138,In_142);
nor U445 (N_445,In_718,In_18);
nor U446 (N_446,In_8,In_247);
nor U447 (N_447,In_604,In_462);
and U448 (N_448,In_745,In_511);
and U449 (N_449,In_405,In_688);
or U450 (N_450,In_683,In_739);
and U451 (N_451,In_3,In_32);
nor U452 (N_452,In_585,In_372);
or U453 (N_453,In_251,In_699);
nand U454 (N_454,In_480,In_500);
nand U455 (N_455,In_9,In_653);
nor U456 (N_456,In_151,In_645);
and U457 (N_457,In_463,In_190);
nand U458 (N_458,In_525,In_688);
and U459 (N_459,In_249,In_570);
nor U460 (N_460,In_37,In_691);
nor U461 (N_461,In_303,In_700);
or U462 (N_462,In_716,In_512);
and U463 (N_463,In_253,In_336);
nand U464 (N_464,In_586,In_225);
and U465 (N_465,In_326,In_379);
and U466 (N_466,In_578,In_533);
and U467 (N_467,In_175,In_240);
or U468 (N_468,In_533,In_538);
nor U469 (N_469,In_450,In_670);
or U470 (N_470,In_529,In_430);
and U471 (N_471,In_508,In_458);
and U472 (N_472,In_418,In_236);
nand U473 (N_473,In_606,In_412);
and U474 (N_474,In_169,In_129);
or U475 (N_475,In_734,In_422);
nand U476 (N_476,In_173,In_473);
or U477 (N_477,In_427,In_101);
and U478 (N_478,In_139,In_363);
or U479 (N_479,In_51,In_623);
nor U480 (N_480,In_109,In_51);
nand U481 (N_481,In_502,In_401);
or U482 (N_482,In_711,In_533);
nand U483 (N_483,In_397,In_439);
and U484 (N_484,In_591,In_63);
nand U485 (N_485,In_151,In_7);
nor U486 (N_486,In_732,In_159);
nor U487 (N_487,In_155,In_573);
nor U488 (N_488,In_267,In_746);
nor U489 (N_489,In_279,In_307);
nand U490 (N_490,In_150,In_493);
or U491 (N_491,In_148,In_269);
and U492 (N_492,In_192,In_734);
and U493 (N_493,In_609,In_570);
nand U494 (N_494,In_431,In_273);
or U495 (N_495,In_66,In_582);
nor U496 (N_496,In_340,In_277);
or U497 (N_497,In_64,In_511);
or U498 (N_498,In_328,In_718);
nand U499 (N_499,In_412,In_437);
and U500 (N_500,In_98,In_55);
nor U501 (N_501,In_426,In_309);
nand U502 (N_502,In_547,In_393);
and U503 (N_503,In_487,In_39);
and U504 (N_504,In_290,In_264);
nand U505 (N_505,In_331,In_619);
and U506 (N_506,In_11,In_143);
and U507 (N_507,In_279,In_572);
nor U508 (N_508,In_512,In_269);
or U509 (N_509,In_216,In_117);
nand U510 (N_510,In_439,In_133);
nor U511 (N_511,In_336,In_63);
and U512 (N_512,In_355,In_28);
nand U513 (N_513,In_748,In_522);
or U514 (N_514,In_603,In_25);
and U515 (N_515,In_517,In_523);
nand U516 (N_516,In_50,In_383);
and U517 (N_517,In_57,In_219);
and U518 (N_518,In_240,In_318);
or U519 (N_519,In_381,In_231);
nor U520 (N_520,In_101,In_4);
or U521 (N_521,In_584,In_579);
nor U522 (N_522,In_389,In_479);
and U523 (N_523,In_301,In_529);
nor U524 (N_524,In_211,In_131);
nor U525 (N_525,In_495,In_664);
nor U526 (N_526,In_224,In_743);
or U527 (N_527,In_745,In_440);
and U528 (N_528,In_735,In_408);
or U529 (N_529,In_539,In_415);
nor U530 (N_530,In_285,In_638);
nor U531 (N_531,In_317,In_359);
or U532 (N_532,In_174,In_291);
nor U533 (N_533,In_593,In_552);
and U534 (N_534,In_537,In_404);
nand U535 (N_535,In_501,In_93);
nor U536 (N_536,In_681,In_669);
nand U537 (N_537,In_566,In_214);
nor U538 (N_538,In_642,In_208);
and U539 (N_539,In_35,In_262);
nand U540 (N_540,In_532,In_109);
and U541 (N_541,In_365,In_385);
and U542 (N_542,In_647,In_616);
or U543 (N_543,In_678,In_364);
or U544 (N_544,In_707,In_403);
nand U545 (N_545,In_690,In_476);
nand U546 (N_546,In_159,In_530);
or U547 (N_547,In_647,In_449);
nand U548 (N_548,In_64,In_237);
or U549 (N_549,In_613,In_53);
nand U550 (N_550,In_242,In_682);
nand U551 (N_551,In_255,In_458);
and U552 (N_552,In_296,In_274);
nand U553 (N_553,In_124,In_30);
and U554 (N_554,In_641,In_698);
and U555 (N_555,In_129,In_57);
or U556 (N_556,In_263,In_189);
and U557 (N_557,In_434,In_359);
or U558 (N_558,In_418,In_134);
and U559 (N_559,In_697,In_695);
nand U560 (N_560,In_332,In_567);
nand U561 (N_561,In_46,In_747);
nor U562 (N_562,In_454,In_64);
nor U563 (N_563,In_284,In_726);
or U564 (N_564,In_262,In_612);
nor U565 (N_565,In_711,In_425);
and U566 (N_566,In_586,In_537);
and U567 (N_567,In_199,In_20);
or U568 (N_568,In_140,In_703);
nand U569 (N_569,In_455,In_83);
or U570 (N_570,In_429,In_254);
nand U571 (N_571,In_589,In_31);
nor U572 (N_572,In_263,In_357);
or U573 (N_573,In_290,In_440);
nand U574 (N_574,In_205,In_673);
or U575 (N_575,In_85,In_530);
or U576 (N_576,In_483,In_58);
and U577 (N_577,In_668,In_153);
nor U578 (N_578,In_455,In_407);
nand U579 (N_579,In_105,In_549);
or U580 (N_580,In_553,In_605);
nand U581 (N_581,In_570,In_722);
or U582 (N_582,In_620,In_75);
nand U583 (N_583,In_735,In_419);
or U584 (N_584,In_153,In_15);
xnor U585 (N_585,In_502,In_598);
nand U586 (N_586,In_442,In_471);
nand U587 (N_587,In_490,In_737);
nor U588 (N_588,In_430,In_260);
nand U589 (N_589,In_613,In_649);
nand U590 (N_590,In_193,In_608);
and U591 (N_591,In_166,In_652);
nand U592 (N_592,In_240,In_714);
and U593 (N_593,In_594,In_295);
nand U594 (N_594,In_618,In_584);
nor U595 (N_595,In_301,In_659);
nor U596 (N_596,In_376,In_629);
nand U597 (N_597,In_628,In_333);
or U598 (N_598,In_189,In_429);
nand U599 (N_599,In_235,In_516);
xnor U600 (N_600,In_675,In_626);
nand U601 (N_601,In_163,In_717);
and U602 (N_602,In_41,In_218);
or U603 (N_603,In_157,In_133);
nor U604 (N_604,In_129,In_664);
and U605 (N_605,In_705,In_511);
and U606 (N_606,In_65,In_120);
nor U607 (N_607,In_514,In_13);
or U608 (N_608,In_3,In_431);
and U609 (N_609,In_26,In_234);
or U610 (N_610,In_429,In_591);
or U611 (N_611,In_232,In_468);
or U612 (N_612,In_429,In_570);
nand U613 (N_613,In_459,In_95);
or U614 (N_614,In_261,In_100);
nand U615 (N_615,In_731,In_505);
nand U616 (N_616,In_255,In_713);
nor U617 (N_617,In_180,In_592);
nand U618 (N_618,In_133,In_522);
or U619 (N_619,In_601,In_344);
xor U620 (N_620,In_128,In_88);
or U621 (N_621,In_219,In_492);
and U622 (N_622,In_531,In_133);
or U623 (N_623,In_535,In_736);
and U624 (N_624,In_512,In_94);
and U625 (N_625,In_142,In_495);
nor U626 (N_626,In_283,In_733);
nor U627 (N_627,In_694,In_447);
and U628 (N_628,In_105,In_35);
nand U629 (N_629,In_400,In_228);
or U630 (N_630,In_665,In_400);
nor U631 (N_631,In_37,In_238);
nor U632 (N_632,In_465,In_366);
or U633 (N_633,In_388,In_671);
or U634 (N_634,In_301,In_107);
nor U635 (N_635,In_125,In_99);
nor U636 (N_636,In_339,In_85);
nor U637 (N_637,In_121,In_246);
and U638 (N_638,In_264,In_403);
nand U639 (N_639,In_30,In_726);
nor U640 (N_640,In_84,In_155);
and U641 (N_641,In_25,In_406);
nor U642 (N_642,In_300,In_220);
nor U643 (N_643,In_137,In_483);
xor U644 (N_644,In_3,In_362);
and U645 (N_645,In_615,In_316);
or U646 (N_646,In_600,In_131);
and U647 (N_647,In_606,In_323);
or U648 (N_648,In_16,In_290);
or U649 (N_649,In_249,In_282);
and U650 (N_650,In_515,In_60);
or U651 (N_651,In_423,In_124);
and U652 (N_652,In_473,In_699);
and U653 (N_653,In_251,In_434);
or U654 (N_654,In_34,In_166);
nand U655 (N_655,In_327,In_58);
xor U656 (N_656,In_191,In_483);
or U657 (N_657,In_279,In_654);
nor U658 (N_658,In_685,In_500);
and U659 (N_659,In_706,In_409);
and U660 (N_660,In_255,In_268);
nand U661 (N_661,In_474,In_664);
or U662 (N_662,In_13,In_498);
and U663 (N_663,In_90,In_628);
nor U664 (N_664,In_375,In_442);
nor U665 (N_665,In_527,In_385);
or U666 (N_666,In_388,In_709);
nor U667 (N_667,In_646,In_251);
nand U668 (N_668,In_409,In_483);
and U669 (N_669,In_746,In_195);
nor U670 (N_670,In_495,In_276);
nor U671 (N_671,In_47,In_567);
nand U672 (N_672,In_284,In_344);
nor U673 (N_673,In_55,In_22);
nand U674 (N_674,In_218,In_524);
nor U675 (N_675,In_81,In_422);
nand U676 (N_676,In_650,In_153);
and U677 (N_677,In_93,In_530);
nor U678 (N_678,In_462,In_241);
and U679 (N_679,In_746,In_341);
nor U680 (N_680,In_390,In_468);
nor U681 (N_681,In_574,In_489);
nand U682 (N_682,In_102,In_724);
nand U683 (N_683,In_398,In_144);
nor U684 (N_684,In_88,In_255);
xnor U685 (N_685,In_49,In_330);
nor U686 (N_686,In_258,In_336);
nor U687 (N_687,In_678,In_14);
nand U688 (N_688,In_294,In_455);
nor U689 (N_689,In_264,In_167);
nor U690 (N_690,In_341,In_8);
nand U691 (N_691,In_24,In_655);
nor U692 (N_692,In_582,In_606);
and U693 (N_693,In_602,In_188);
and U694 (N_694,In_101,In_440);
and U695 (N_695,In_91,In_177);
or U696 (N_696,In_414,In_351);
and U697 (N_697,In_369,In_427);
or U698 (N_698,In_375,In_7);
or U699 (N_699,In_277,In_273);
and U700 (N_700,In_448,In_254);
xor U701 (N_701,In_302,In_647);
and U702 (N_702,In_688,In_194);
or U703 (N_703,In_464,In_393);
and U704 (N_704,In_278,In_130);
and U705 (N_705,In_387,In_686);
and U706 (N_706,In_279,In_207);
or U707 (N_707,In_369,In_564);
or U708 (N_708,In_515,In_119);
or U709 (N_709,In_513,In_251);
nand U710 (N_710,In_273,In_425);
and U711 (N_711,In_105,In_715);
nand U712 (N_712,In_617,In_453);
or U713 (N_713,In_85,In_724);
nor U714 (N_714,In_694,In_610);
nor U715 (N_715,In_332,In_40);
or U716 (N_716,In_676,In_107);
or U717 (N_717,In_223,In_171);
nand U718 (N_718,In_133,In_287);
nor U719 (N_719,In_329,In_308);
nor U720 (N_720,In_598,In_131);
or U721 (N_721,In_728,In_250);
nor U722 (N_722,In_391,In_489);
nor U723 (N_723,In_230,In_209);
or U724 (N_724,In_48,In_50);
and U725 (N_725,In_118,In_191);
or U726 (N_726,In_659,In_132);
nor U727 (N_727,In_263,In_696);
nor U728 (N_728,In_322,In_598);
nor U729 (N_729,In_25,In_744);
and U730 (N_730,In_470,In_141);
nor U731 (N_731,In_516,In_191);
and U732 (N_732,In_369,In_448);
nor U733 (N_733,In_267,In_475);
and U734 (N_734,In_6,In_392);
or U735 (N_735,In_148,In_689);
nor U736 (N_736,In_261,In_29);
nand U737 (N_737,In_54,In_633);
nor U738 (N_738,In_533,In_404);
and U739 (N_739,In_344,In_402);
and U740 (N_740,In_77,In_667);
or U741 (N_741,In_667,In_636);
nor U742 (N_742,In_734,In_111);
nor U743 (N_743,In_478,In_449);
nor U744 (N_744,In_22,In_95);
nand U745 (N_745,In_93,In_406);
and U746 (N_746,In_266,In_434);
nand U747 (N_747,In_28,In_431);
or U748 (N_748,In_107,In_489);
nor U749 (N_749,In_9,In_691);
and U750 (N_750,In_3,In_401);
or U751 (N_751,In_187,In_424);
or U752 (N_752,In_220,In_30);
or U753 (N_753,In_554,In_264);
nor U754 (N_754,In_40,In_643);
nor U755 (N_755,In_67,In_645);
nand U756 (N_756,In_481,In_320);
nand U757 (N_757,In_721,In_182);
and U758 (N_758,In_718,In_644);
nand U759 (N_759,In_274,In_102);
or U760 (N_760,In_424,In_176);
or U761 (N_761,In_359,In_524);
nand U762 (N_762,In_330,In_480);
nor U763 (N_763,In_117,In_253);
xnor U764 (N_764,In_113,In_28);
nand U765 (N_765,In_31,In_428);
nand U766 (N_766,In_292,In_392);
nor U767 (N_767,In_324,In_659);
or U768 (N_768,In_607,In_13);
or U769 (N_769,In_647,In_52);
xnor U770 (N_770,In_192,In_593);
and U771 (N_771,In_462,In_212);
or U772 (N_772,In_357,In_251);
or U773 (N_773,In_694,In_738);
or U774 (N_774,In_377,In_24);
or U775 (N_775,In_566,In_114);
and U776 (N_776,In_501,In_482);
nor U777 (N_777,In_96,In_314);
nor U778 (N_778,In_448,In_619);
nor U779 (N_779,In_196,In_546);
nand U780 (N_780,In_346,In_8);
and U781 (N_781,In_317,In_694);
nand U782 (N_782,In_736,In_47);
nor U783 (N_783,In_409,In_113);
nand U784 (N_784,In_300,In_536);
nand U785 (N_785,In_708,In_16);
and U786 (N_786,In_588,In_545);
or U787 (N_787,In_663,In_718);
and U788 (N_788,In_293,In_504);
nand U789 (N_789,In_338,In_252);
nor U790 (N_790,In_658,In_69);
nor U791 (N_791,In_360,In_748);
nand U792 (N_792,In_331,In_168);
nand U793 (N_793,In_499,In_38);
or U794 (N_794,In_665,In_137);
and U795 (N_795,In_259,In_158);
or U796 (N_796,In_157,In_219);
and U797 (N_797,In_312,In_117);
nand U798 (N_798,In_651,In_118);
and U799 (N_799,In_321,In_356);
nor U800 (N_800,In_201,In_82);
nor U801 (N_801,In_324,In_232);
and U802 (N_802,In_507,In_262);
nor U803 (N_803,In_342,In_66);
nor U804 (N_804,In_490,In_316);
or U805 (N_805,In_584,In_251);
nor U806 (N_806,In_680,In_278);
or U807 (N_807,In_563,In_442);
nand U808 (N_808,In_714,In_481);
nand U809 (N_809,In_88,In_628);
nor U810 (N_810,In_515,In_546);
and U811 (N_811,In_90,In_684);
nand U812 (N_812,In_258,In_312);
and U813 (N_813,In_215,In_686);
nand U814 (N_814,In_387,In_75);
and U815 (N_815,In_313,In_509);
and U816 (N_816,In_465,In_107);
nand U817 (N_817,In_624,In_86);
nor U818 (N_818,In_264,In_524);
nand U819 (N_819,In_730,In_652);
nor U820 (N_820,In_702,In_660);
nand U821 (N_821,In_368,In_36);
nand U822 (N_822,In_367,In_223);
nand U823 (N_823,In_691,In_521);
and U824 (N_824,In_13,In_634);
and U825 (N_825,In_377,In_395);
and U826 (N_826,In_81,In_283);
or U827 (N_827,In_652,In_317);
nor U828 (N_828,In_132,In_727);
or U829 (N_829,In_258,In_152);
nor U830 (N_830,In_245,In_274);
nor U831 (N_831,In_382,In_713);
and U832 (N_832,In_271,In_274);
nor U833 (N_833,In_200,In_256);
and U834 (N_834,In_457,In_103);
or U835 (N_835,In_746,In_712);
nor U836 (N_836,In_487,In_534);
nand U837 (N_837,In_15,In_462);
or U838 (N_838,In_415,In_264);
nand U839 (N_839,In_656,In_216);
and U840 (N_840,In_227,In_600);
or U841 (N_841,In_561,In_120);
or U842 (N_842,In_330,In_733);
nand U843 (N_843,In_421,In_166);
or U844 (N_844,In_83,In_423);
nor U845 (N_845,In_115,In_711);
and U846 (N_846,In_491,In_690);
or U847 (N_847,In_674,In_281);
nand U848 (N_848,In_374,In_321);
and U849 (N_849,In_668,In_10);
and U850 (N_850,In_309,In_638);
nand U851 (N_851,In_23,In_447);
nand U852 (N_852,In_633,In_120);
or U853 (N_853,In_554,In_409);
nor U854 (N_854,In_153,In_736);
nor U855 (N_855,In_612,In_86);
nor U856 (N_856,In_717,In_168);
nand U857 (N_857,In_472,In_697);
and U858 (N_858,In_315,In_589);
nand U859 (N_859,In_692,In_76);
nor U860 (N_860,In_505,In_265);
nor U861 (N_861,In_370,In_297);
nand U862 (N_862,In_377,In_687);
and U863 (N_863,In_182,In_552);
nand U864 (N_864,In_598,In_48);
or U865 (N_865,In_609,In_440);
nand U866 (N_866,In_141,In_697);
nand U867 (N_867,In_494,In_502);
nand U868 (N_868,In_221,In_745);
and U869 (N_869,In_169,In_230);
nand U870 (N_870,In_396,In_441);
nand U871 (N_871,In_631,In_516);
or U872 (N_872,In_41,In_177);
nor U873 (N_873,In_660,In_41);
and U874 (N_874,In_619,In_9);
nand U875 (N_875,In_189,In_411);
nor U876 (N_876,In_198,In_408);
nand U877 (N_877,In_461,In_231);
nand U878 (N_878,In_274,In_418);
or U879 (N_879,In_468,In_54);
nand U880 (N_880,In_215,In_629);
nand U881 (N_881,In_695,In_276);
nor U882 (N_882,In_34,In_113);
nand U883 (N_883,In_260,In_109);
nor U884 (N_884,In_367,In_263);
nor U885 (N_885,In_491,In_559);
and U886 (N_886,In_161,In_627);
nor U887 (N_887,In_120,In_218);
nor U888 (N_888,In_316,In_609);
nand U889 (N_889,In_509,In_616);
and U890 (N_890,In_157,In_357);
and U891 (N_891,In_553,In_677);
and U892 (N_892,In_531,In_621);
nand U893 (N_893,In_318,In_97);
or U894 (N_894,In_273,In_190);
nor U895 (N_895,In_298,In_123);
nand U896 (N_896,In_124,In_694);
and U897 (N_897,In_669,In_153);
nand U898 (N_898,In_4,In_168);
nand U899 (N_899,In_524,In_58);
nand U900 (N_900,In_743,In_114);
nand U901 (N_901,In_604,In_453);
nand U902 (N_902,In_604,In_458);
and U903 (N_903,In_0,In_706);
or U904 (N_904,In_237,In_715);
xnor U905 (N_905,In_551,In_110);
or U906 (N_906,In_80,In_127);
nor U907 (N_907,In_518,In_63);
nand U908 (N_908,In_355,In_638);
and U909 (N_909,In_453,In_532);
nor U910 (N_910,In_681,In_228);
nand U911 (N_911,In_371,In_236);
nand U912 (N_912,In_10,In_741);
nor U913 (N_913,In_179,In_21);
nand U914 (N_914,In_667,In_429);
nor U915 (N_915,In_465,In_8);
nor U916 (N_916,In_176,In_23);
nor U917 (N_917,In_167,In_500);
nor U918 (N_918,In_59,In_172);
nor U919 (N_919,In_527,In_509);
xor U920 (N_920,In_134,In_274);
nand U921 (N_921,In_205,In_79);
nand U922 (N_922,In_589,In_573);
nand U923 (N_923,In_233,In_50);
nand U924 (N_924,In_571,In_422);
nor U925 (N_925,In_475,In_381);
nand U926 (N_926,In_630,In_242);
nor U927 (N_927,In_361,In_244);
or U928 (N_928,In_113,In_438);
xor U929 (N_929,In_267,In_378);
and U930 (N_930,In_340,In_667);
and U931 (N_931,In_437,In_88);
and U932 (N_932,In_187,In_178);
and U933 (N_933,In_228,In_193);
or U934 (N_934,In_571,In_743);
and U935 (N_935,In_600,In_465);
and U936 (N_936,In_307,In_344);
nand U937 (N_937,In_274,In_337);
and U938 (N_938,In_702,In_547);
nor U939 (N_939,In_248,In_91);
and U940 (N_940,In_537,In_48);
and U941 (N_941,In_245,In_585);
and U942 (N_942,In_188,In_460);
or U943 (N_943,In_16,In_271);
and U944 (N_944,In_115,In_506);
and U945 (N_945,In_466,In_208);
and U946 (N_946,In_693,In_248);
nand U947 (N_947,In_581,In_569);
and U948 (N_948,In_680,In_344);
nor U949 (N_949,In_737,In_110);
or U950 (N_950,In_729,In_582);
nor U951 (N_951,In_642,In_185);
or U952 (N_952,In_21,In_499);
or U953 (N_953,In_337,In_606);
or U954 (N_954,In_47,In_265);
and U955 (N_955,In_337,In_492);
or U956 (N_956,In_699,In_62);
nand U957 (N_957,In_107,In_166);
or U958 (N_958,In_467,In_539);
and U959 (N_959,In_677,In_706);
or U960 (N_960,In_730,In_182);
nor U961 (N_961,In_483,In_599);
xnor U962 (N_962,In_428,In_371);
or U963 (N_963,In_89,In_363);
and U964 (N_964,In_359,In_657);
xnor U965 (N_965,In_435,In_322);
and U966 (N_966,In_149,In_277);
nor U967 (N_967,In_665,In_401);
nand U968 (N_968,In_727,In_383);
and U969 (N_969,In_168,In_609);
nand U970 (N_970,In_576,In_475);
nor U971 (N_971,In_728,In_547);
nor U972 (N_972,In_88,In_526);
or U973 (N_973,In_695,In_599);
and U974 (N_974,In_247,In_494);
xnor U975 (N_975,In_471,In_566);
nand U976 (N_976,In_573,In_309);
and U977 (N_977,In_256,In_357);
or U978 (N_978,In_137,In_401);
nand U979 (N_979,In_642,In_71);
or U980 (N_980,In_655,In_455);
and U981 (N_981,In_129,In_179);
nor U982 (N_982,In_399,In_536);
or U983 (N_983,In_421,In_74);
or U984 (N_984,In_209,In_49);
nand U985 (N_985,In_425,In_678);
and U986 (N_986,In_50,In_627);
nor U987 (N_987,In_734,In_117);
and U988 (N_988,In_531,In_685);
or U989 (N_989,In_179,In_62);
nor U990 (N_990,In_226,In_575);
or U991 (N_991,In_398,In_258);
nor U992 (N_992,In_162,In_729);
nand U993 (N_993,In_215,In_608);
and U994 (N_994,In_638,In_358);
nor U995 (N_995,In_699,In_717);
or U996 (N_996,In_515,In_566);
and U997 (N_997,In_425,In_515);
nand U998 (N_998,In_114,In_274);
or U999 (N_999,In_335,In_215);
and U1000 (N_1000,N_528,N_122);
and U1001 (N_1001,N_55,N_870);
and U1002 (N_1002,N_23,N_495);
nor U1003 (N_1003,N_9,N_754);
nor U1004 (N_1004,N_626,N_649);
and U1005 (N_1005,N_401,N_133);
or U1006 (N_1006,N_197,N_670);
or U1007 (N_1007,N_935,N_387);
nor U1008 (N_1008,N_169,N_116);
nand U1009 (N_1009,N_609,N_155);
nor U1010 (N_1010,N_255,N_981);
nand U1011 (N_1011,N_10,N_687);
and U1012 (N_1012,N_764,N_202);
nor U1013 (N_1013,N_132,N_845);
nand U1014 (N_1014,N_758,N_983);
nor U1015 (N_1015,N_120,N_170);
nand U1016 (N_1016,N_59,N_13);
or U1017 (N_1017,N_242,N_529);
or U1018 (N_1018,N_767,N_549);
and U1019 (N_1019,N_479,N_324);
and U1020 (N_1020,N_821,N_444);
and U1021 (N_1021,N_0,N_276);
nand U1022 (N_1022,N_641,N_838);
nor U1023 (N_1023,N_511,N_623);
nor U1024 (N_1024,N_866,N_857);
nor U1025 (N_1025,N_141,N_910);
nand U1026 (N_1026,N_289,N_553);
xor U1027 (N_1027,N_299,N_968);
nand U1028 (N_1028,N_512,N_157);
or U1029 (N_1029,N_265,N_320);
nor U1030 (N_1030,N_628,N_582);
nor U1031 (N_1031,N_616,N_663);
nand U1032 (N_1032,N_347,N_83);
or U1033 (N_1033,N_538,N_505);
nor U1034 (N_1034,N_638,N_946);
xnor U1035 (N_1035,N_219,N_806);
and U1036 (N_1036,N_636,N_35);
nand U1037 (N_1037,N_251,N_514);
nand U1038 (N_1038,N_556,N_913);
and U1039 (N_1039,N_633,N_621);
nand U1040 (N_1040,N_858,N_301);
nand U1041 (N_1041,N_568,N_381);
or U1042 (N_1042,N_292,N_229);
nor U1043 (N_1043,N_379,N_642);
nor U1044 (N_1044,N_708,N_924);
nor U1045 (N_1045,N_147,N_646);
nor U1046 (N_1046,N_489,N_90);
nand U1047 (N_1047,N_368,N_397);
or U1048 (N_1048,N_825,N_341);
nor U1049 (N_1049,N_565,N_519);
and U1050 (N_1050,N_839,N_305);
or U1051 (N_1051,N_833,N_909);
or U1052 (N_1052,N_793,N_214);
and U1053 (N_1053,N_830,N_238);
nor U1054 (N_1054,N_21,N_541);
nor U1055 (N_1055,N_149,N_325);
nor U1056 (N_1056,N_940,N_989);
nand U1057 (N_1057,N_225,N_603);
or U1058 (N_1058,N_5,N_901);
or U1059 (N_1059,N_645,N_490);
and U1060 (N_1060,N_578,N_705);
or U1061 (N_1061,N_82,N_745);
and U1062 (N_1062,N_486,N_861);
nand U1063 (N_1063,N_716,N_810);
or U1064 (N_1064,N_683,N_611);
and U1065 (N_1065,N_483,N_769);
and U1066 (N_1066,N_762,N_117);
or U1067 (N_1067,N_634,N_900);
or U1068 (N_1068,N_832,N_28);
nor U1069 (N_1069,N_664,N_25);
nand U1070 (N_1070,N_159,N_156);
nand U1071 (N_1071,N_482,N_759);
or U1072 (N_1072,N_58,N_692);
or U1073 (N_1073,N_354,N_186);
and U1074 (N_1074,N_322,N_308);
or U1075 (N_1075,N_882,N_414);
nor U1076 (N_1076,N_163,N_856);
nor U1077 (N_1077,N_213,N_853);
or U1078 (N_1078,N_481,N_784);
nand U1079 (N_1079,N_698,N_417);
nor U1080 (N_1080,N_485,N_287);
nand U1081 (N_1081,N_198,N_343);
and U1082 (N_1082,N_441,N_91);
or U1083 (N_1083,N_96,N_463);
or U1084 (N_1084,N_370,N_721);
and U1085 (N_1085,N_302,N_624);
or U1086 (N_1086,N_46,N_979);
nand U1087 (N_1087,N_748,N_209);
and U1088 (N_1088,N_392,N_936);
and U1089 (N_1089,N_886,N_877);
nor U1090 (N_1090,N_523,N_190);
nand U1091 (N_1091,N_399,N_334);
nor U1092 (N_1092,N_434,N_798);
nand U1093 (N_1093,N_563,N_988);
nor U1094 (N_1094,N_797,N_904);
nand U1095 (N_1095,N_799,N_164);
or U1096 (N_1096,N_182,N_244);
or U1097 (N_1097,N_588,N_267);
or U1098 (N_1098,N_171,N_312);
nand U1099 (N_1099,N_637,N_760);
or U1100 (N_1100,N_390,N_786);
and U1101 (N_1101,N_977,N_696);
xor U1102 (N_1102,N_498,N_232);
or U1103 (N_1103,N_307,N_504);
nand U1104 (N_1104,N_879,N_569);
and U1105 (N_1105,N_819,N_377);
nor U1106 (N_1106,N_772,N_816);
or U1107 (N_1107,N_871,N_233);
nand U1108 (N_1108,N_775,N_329);
nand U1109 (N_1109,N_540,N_718);
or U1110 (N_1110,N_506,N_752);
nor U1111 (N_1111,N_831,N_420);
or U1112 (N_1112,N_321,N_52);
nand U1113 (N_1113,N_532,N_67);
nand U1114 (N_1114,N_261,N_84);
nor U1115 (N_1115,N_773,N_252);
nor U1116 (N_1116,N_63,N_491);
nand U1117 (N_1117,N_531,N_827);
and U1118 (N_1118,N_181,N_820);
nand U1119 (N_1119,N_185,N_126);
or U1120 (N_1120,N_749,N_560);
nor U1121 (N_1121,N_855,N_310);
or U1122 (N_1122,N_515,N_756);
nor U1123 (N_1123,N_602,N_211);
and U1124 (N_1124,N_223,N_475);
xnor U1125 (N_1125,N_7,N_939);
and U1126 (N_1126,N_509,N_889);
or U1127 (N_1127,N_594,N_34);
or U1128 (N_1128,N_258,N_689);
or U1129 (N_1129,N_525,N_818);
nand U1130 (N_1130,N_778,N_448);
and U1131 (N_1131,N_407,N_81);
or U1132 (N_1132,N_524,N_427);
and U1133 (N_1133,N_520,N_224);
nand U1134 (N_1134,N_597,N_707);
nand U1135 (N_1135,N_610,N_927);
and U1136 (N_1136,N_631,N_595);
nor U1137 (N_1137,N_694,N_45);
or U1138 (N_1138,N_26,N_837);
or U1139 (N_1139,N_559,N_766);
or U1140 (N_1140,N_235,N_207);
and U1141 (N_1141,N_279,N_393);
nand U1142 (N_1142,N_576,N_192);
nor U1143 (N_1143,N_620,N_899);
or U1144 (N_1144,N_761,N_554);
nor U1145 (N_1145,N_739,N_323);
or U1146 (N_1146,N_517,N_421);
or U1147 (N_1147,N_194,N_57);
nor U1148 (N_1148,N_848,N_375);
xnor U1149 (N_1149,N_829,N_791);
and U1150 (N_1150,N_906,N_105);
nor U1151 (N_1151,N_885,N_629);
nand U1152 (N_1152,N_562,N_311);
and U1153 (N_1153,N_187,N_389);
nand U1154 (N_1154,N_932,N_89);
and U1155 (N_1155,N_632,N_271);
nand U1156 (N_1156,N_945,N_102);
nand U1157 (N_1157,N_947,N_622);
nor U1158 (N_1158,N_286,N_403);
nor U1159 (N_1159,N_44,N_521);
and U1160 (N_1160,N_706,N_774);
nor U1161 (N_1161,N_39,N_558);
or U1162 (N_1162,N_66,N_297);
and U1163 (N_1163,N_342,N_776);
or U1164 (N_1164,N_815,N_24);
or U1165 (N_1165,N_914,N_113);
nand U1166 (N_1166,N_435,N_476);
or U1167 (N_1167,N_571,N_550);
or U1168 (N_1168,N_250,N_941);
nor U1169 (N_1169,N_513,N_22);
and U1170 (N_1170,N_348,N_350);
and U1171 (N_1171,N_934,N_11);
and U1172 (N_1172,N_919,N_166);
xor U1173 (N_1173,N_564,N_872);
or U1174 (N_1174,N_733,N_240);
nand U1175 (N_1175,N_655,N_743);
nand U1176 (N_1176,N_823,N_65);
and U1177 (N_1177,N_445,N_15);
and U1178 (N_1178,N_953,N_875);
and U1179 (N_1179,N_691,N_777);
and U1180 (N_1180,N_916,N_443);
or U1181 (N_1181,N_152,N_811);
or U1182 (N_1182,N_148,N_253);
or U1183 (N_1183,N_805,N_896);
nand U1184 (N_1184,N_405,N_813);
nor U1185 (N_1185,N_165,N_129);
or U1186 (N_1186,N_690,N_577);
or U1187 (N_1187,N_724,N_902);
nand U1188 (N_1188,N_416,N_175);
or U1189 (N_1189,N_168,N_471);
and U1190 (N_1190,N_836,N_503);
nand U1191 (N_1191,N_959,N_822);
nand U1192 (N_1192,N_136,N_215);
and U1193 (N_1193,N_455,N_138);
or U1194 (N_1194,N_230,N_787);
nand U1195 (N_1195,N_309,N_440);
and U1196 (N_1196,N_100,N_867);
and U1197 (N_1197,N_33,N_684);
nand U1198 (N_1198,N_300,N_682);
nand U1199 (N_1199,N_993,N_627);
or U1200 (N_1200,N_876,N_472);
and U1201 (N_1201,N_336,N_804);
nand U1202 (N_1202,N_709,N_20);
or U1203 (N_1203,N_411,N_931);
nor U1204 (N_1204,N_770,N_176);
nor U1205 (N_1205,N_618,N_703);
or U1206 (N_1206,N_742,N_651);
and U1207 (N_1207,N_842,N_704);
or U1208 (N_1208,N_720,N_677);
and U1209 (N_1209,N_31,N_353);
and U1210 (N_1210,N_468,N_281);
nor U1211 (N_1211,N_275,N_231);
nor U1212 (N_1212,N_142,N_254);
nor U1213 (N_1213,N_847,N_359);
nand U1214 (N_1214,N_154,N_277);
nand U1215 (N_1215,N_178,N_542);
and U1216 (N_1216,N_296,N_710);
nand U1217 (N_1217,N_917,N_41);
and U1218 (N_1218,N_543,N_51);
and U1219 (N_1219,N_747,N_883);
or U1220 (N_1220,N_949,N_119);
nor U1221 (N_1221,N_501,N_608);
nor U1222 (N_1222,N_3,N_60);
or U1223 (N_1223,N_734,N_903);
and U1224 (N_1224,N_54,N_714);
or U1225 (N_1225,N_458,N_400);
and U1226 (N_1226,N_386,N_954);
nand U1227 (N_1227,N_32,N_75);
nand U1228 (N_1228,N_413,N_922);
and U1229 (N_1229,N_408,N_685);
or U1230 (N_1230,N_526,N_966);
and U1231 (N_1231,N_62,N_357);
or U1232 (N_1232,N_881,N_817);
nand U1233 (N_1233,N_278,N_313);
and U1234 (N_1234,N_380,N_730);
nand U1235 (N_1235,N_671,N_680);
or U1236 (N_1236,N_371,N_728);
nand U1237 (N_1237,N_107,N_644);
nor U1238 (N_1238,N_237,N_80);
and U1239 (N_1239,N_969,N_601);
nor U1240 (N_1240,N_667,N_264);
or U1241 (N_1241,N_199,N_139);
nor U1242 (N_1242,N_890,N_109);
nand U1243 (N_1243,N_162,N_183);
nand U1244 (N_1244,N_454,N_161);
or U1245 (N_1245,N_256,N_587);
xnor U1246 (N_1246,N_315,N_702);
nor U1247 (N_1247,N_121,N_727);
or U1248 (N_1248,N_128,N_469);
nand U1249 (N_1249,N_658,N_226);
or U1250 (N_1250,N_803,N_738);
nor U1251 (N_1251,N_318,N_473);
or U1252 (N_1252,N_42,N_790);
or U1253 (N_1253,N_920,N_339);
and U1254 (N_1254,N_561,N_729);
nor U1255 (N_1255,N_335,N_928);
nor U1256 (N_1256,N_755,N_284);
or U1257 (N_1257,N_111,N_585);
nor U1258 (N_1258,N_78,N_765);
and U1259 (N_1259,N_763,N_669);
nor U1260 (N_1260,N_85,N_688);
nand U1261 (N_1261,N_404,N_656);
nor U1262 (N_1262,N_964,N_502);
nand U1263 (N_1263,N_146,N_27);
nand U1264 (N_1264,N_884,N_452);
nor U1265 (N_1265,N_184,N_895);
nor U1266 (N_1266,N_768,N_840);
and U1267 (N_1267,N_952,N_195);
or U1268 (N_1268,N_358,N_783);
or U1269 (N_1269,N_650,N_589);
and U1270 (N_1270,N_852,N_665);
nand U1271 (N_1271,N_480,N_317);
nand U1272 (N_1272,N_746,N_863);
nand U1273 (N_1273,N_662,N_868);
nor U1274 (N_1274,N_672,N_555);
nand U1275 (N_1275,N_807,N_534);
or U1276 (N_1276,N_432,N_835);
and U1277 (N_1277,N_1,N_474);
and U1278 (N_1278,N_639,N_544);
nor U1279 (N_1279,N_779,N_998);
nor U1280 (N_1280,N_77,N_206);
nor U1281 (N_1281,N_911,N_590);
and U1282 (N_1282,N_484,N_94);
nor U1283 (N_1283,N_994,N_826);
nor U1284 (N_1284,N_851,N_374);
or U1285 (N_1285,N_530,N_573);
nor U1286 (N_1286,N_812,N_4);
nand U1287 (N_1287,N_869,N_640);
nor U1288 (N_1288,N_795,N_99);
and U1289 (N_1289,N_189,N_196);
nor U1290 (N_1290,N_48,N_316);
nand U1291 (N_1291,N_70,N_127);
nor U1292 (N_1292,N_566,N_864);
or U1293 (N_1293,N_293,N_272);
and U1294 (N_1294,N_905,N_686);
nor U1295 (N_1295,N_216,N_666);
and U1296 (N_1296,N_438,N_955);
and U1297 (N_1297,N_364,N_948);
nor U1298 (N_1298,N_137,N_679);
and U1299 (N_1299,N_282,N_700);
and U1300 (N_1300,N_970,N_892);
nor U1301 (N_1301,N_647,N_598);
or U1302 (N_1302,N_878,N_101);
xor U1303 (N_1303,N_918,N_2);
nand U1304 (N_1304,N_247,N_228);
and U1305 (N_1305,N_56,N_249);
nand U1306 (N_1306,N_736,N_973);
and U1307 (N_1307,N_453,N_956);
nor U1308 (N_1308,N_151,N_982);
and U1309 (N_1309,N_372,N_987);
and U1310 (N_1310,N_789,N_923);
nor U1311 (N_1311,N_103,N_681);
xor U1312 (N_1312,N_160,N_410);
and U1313 (N_1313,N_391,N_723);
nand U1314 (N_1314,N_263,N_652);
and U1315 (N_1315,N_464,N_290);
or U1316 (N_1316,N_140,N_897);
or U1317 (N_1317,N_725,N_356);
or U1318 (N_1318,N_697,N_114);
or U1319 (N_1319,N_6,N_280);
nand U1320 (N_1320,N_430,N_257);
xor U1321 (N_1321,N_18,N_925);
nand U1322 (N_1322,N_97,N_780);
nor U1323 (N_1323,N_201,N_893);
nand U1324 (N_1324,N_958,N_446);
nor U1325 (N_1325,N_50,N_536);
nand U1326 (N_1326,N_986,N_337);
nor U1327 (N_1327,N_492,N_266);
nand U1328 (N_1328,N_625,N_614);
nand U1329 (N_1329,N_737,N_960);
nand U1330 (N_1330,N_596,N_442);
and U1331 (N_1331,N_447,N_731);
nand U1332 (N_1332,N_217,N_367);
nor U1333 (N_1333,N_615,N_500);
nand U1334 (N_1334,N_303,N_732);
nand U1335 (N_1335,N_288,N_929);
nor U1336 (N_1336,N_507,N_788);
nor U1337 (N_1337,N_873,N_285);
and U1338 (N_1338,N_385,N_539);
xor U1339 (N_1339,N_771,N_841);
or U1340 (N_1340,N_314,N_30);
and U1341 (N_1341,N_584,N_131);
and U1342 (N_1342,N_488,N_984);
nand U1343 (N_1343,N_753,N_557);
or U1344 (N_1344,N_346,N_355);
or U1345 (N_1345,N_674,N_294);
or U1346 (N_1346,N_497,N_980);
and U1347 (N_1347,N_974,N_188);
and U1348 (N_1348,N_996,N_369);
nand U1349 (N_1349,N_978,N_824);
nand U1350 (N_1350,N_715,N_106);
nor U1351 (N_1351,N_844,N_951);
nand U1352 (N_1352,N_802,N_49);
or U1353 (N_1353,N_880,N_834);
or U1354 (N_1354,N_466,N_657);
nor U1355 (N_1355,N_874,N_792);
nand U1356 (N_1356,N_363,N_398);
and U1357 (N_1357,N_961,N_963);
and U1358 (N_1358,N_362,N_349);
nand U1359 (N_1359,N_361,N_428);
nor U1360 (N_1360,N_548,N_533);
and U1361 (N_1361,N_319,N_814);
nand U1362 (N_1362,N_220,N_332);
or U1363 (N_1363,N_551,N_248);
or U1364 (N_1364,N_699,N_93);
nor U1365 (N_1365,N_124,N_545);
and U1366 (N_1366,N_173,N_957);
and U1367 (N_1367,N_383,N_193);
nand U1368 (N_1368,N_575,N_415);
or U1369 (N_1369,N_930,N_887);
nand U1370 (N_1370,N_236,N_972);
nor U1371 (N_1371,N_908,N_260);
and U1372 (N_1372,N_72,N_579);
nand U1373 (N_1373,N_567,N_604);
nor U1374 (N_1374,N_376,N_304);
and U1375 (N_1375,N_693,N_351);
nand U1376 (N_1376,N_907,N_172);
or U1377 (N_1377,N_912,N_535);
nor U1378 (N_1378,N_995,N_145);
nor U1379 (N_1379,N_123,N_843);
nor U1380 (N_1380,N_613,N_808);
or U1381 (N_1381,N_246,N_331);
nor U1382 (N_1382,N_108,N_241);
or U1383 (N_1383,N_200,N_478);
or U1384 (N_1384,N_378,N_898);
or U1385 (N_1385,N_751,N_850);
nand U1386 (N_1386,N_68,N_713);
and U1387 (N_1387,N_177,N_991);
or U1388 (N_1388,N_16,N_104);
and U1389 (N_1389,N_586,N_467);
or U1390 (N_1390,N_926,N_673);
nor U1391 (N_1391,N_326,N_888);
nand U1392 (N_1392,N_43,N_298);
nor U1393 (N_1393,N_654,N_150);
nand U1394 (N_1394,N_431,N_205);
and U1395 (N_1395,N_419,N_274);
or U1396 (N_1396,N_962,N_345);
nor U1397 (N_1397,N_678,N_8);
nand U1398 (N_1398,N_426,N_118);
nand U1399 (N_1399,N_865,N_143);
nor U1400 (N_1400,N_394,N_422);
nand U1401 (N_1401,N_459,N_429);
nor U1402 (N_1402,N_17,N_659);
nand U1403 (N_1403,N_412,N_239);
or U1404 (N_1404,N_617,N_997);
or U1405 (N_1405,N_360,N_757);
and U1406 (N_1406,N_268,N_809);
nor U1407 (N_1407,N_675,N_894);
or U1408 (N_1408,N_915,N_950);
nor U1409 (N_1409,N_406,N_933);
nor U1410 (N_1410,N_270,N_781);
and U1411 (N_1411,N_262,N_676);
nand U1412 (N_1412,N_942,N_717);
nor U1413 (N_1413,N_701,N_508);
xor U1414 (N_1414,N_741,N_36);
nand U1415 (N_1415,N_660,N_88);
and U1416 (N_1416,N_552,N_418);
and U1417 (N_1417,N_937,N_53);
and U1418 (N_1418,N_547,N_846);
nor U1419 (N_1419,N_179,N_330);
and U1420 (N_1420,N_599,N_158);
and U1421 (N_1421,N_273,N_643);
or U1422 (N_1422,N_487,N_366);
and U1423 (N_1423,N_985,N_86);
nand U1424 (N_1424,N_40,N_47);
or U1425 (N_1425,N_465,N_327);
nand U1426 (N_1426,N_135,N_352);
xor U1427 (N_1427,N_648,N_395);
nor U1428 (N_1428,N_891,N_944);
nand U1429 (N_1429,N_19,N_74);
or U1430 (N_1430,N_607,N_295);
xnor U1431 (N_1431,N_965,N_37);
nor U1432 (N_1432,N_462,N_456);
nor U1433 (N_1433,N_494,N_661);
or U1434 (N_1434,N_967,N_735);
nor U1435 (N_1435,N_130,N_695);
nor U1436 (N_1436,N_782,N_69);
nand U1437 (N_1437,N_451,N_457);
or U1438 (N_1438,N_581,N_328);
or U1439 (N_1439,N_191,N_990);
or U1440 (N_1440,N_437,N_800);
nand U1441 (N_1441,N_794,N_570);
nand U1442 (N_1442,N_291,N_860);
nor U1443 (N_1443,N_971,N_134);
and U1444 (N_1444,N_98,N_854);
nand U1445 (N_1445,N_493,N_516);
nor U1446 (N_1446,N_245,N_499);
nand U1447 (N_1447,N_227,N_976);
and U1448 (N_1448,N_71,N_269);
nand U1449 (N_1449,N_388,N_859);
nor U1450 (N_1450,N_344,N_938);
or U1451 (N_1451,N_180,N_439);
and U1452 (N_1452,N_630,N_999);
and U1453 (N_1453,N_653,N_712);
nor U1454 (N_1454,N_174,N_283);
or U1455 (N_1455,N_744,N_112);
xor U1456 (N_1456,N_384,N_64);
nor U1457 (N_1457,N_975,N_340);
nand U1458 (N_1458,N_306,N_450);
or U1459 (N_1459,N_522,N_409);
and U1460 (N_1460,N_76,N_591);
nand U1461 (N_1461,N_203,N_110);
nand U1462 (N_1462,N_612,N_750);
or U1463 (N_1463,N_605,N_259);
nand U1464 (N_1464,N_719,N_92);
or U1465 (N_1465,N_580,N_992);
or U1466 (N_1466,N_204,N_510);
nor U1467 (N_1467,N_449,N_365);
nand U1468 (N_1468,N_221,N_153);
nor U1469 (N_1469,N_338,N_12);
and U1470 (N_1470,N_95,N_14);
nand U1471 (N_1471,N_600,N_496);
nand U1472 (N_1472,N_740,N_583);
nor U1473 (N_1473,N_210,N_218);
and U1474 (N_1474,N_593,N_635);
and U1475 (N_1475,N_785,N_828);
and U1476 (N_1476,N_73,N_396);
nand U1477 (N_1477,N_796,N_862);
nor U1478 (N_1478,N_222,N_115);
nor U1479 (N_1479,N_574,N_243);
nor U1480 (N_1480,N_38,N_433);
nor U1481 (N_1481,N_425,N_79);
nor U1482 (N_1482,N_592,N_572);
or U1483 (N_1483,N_424,N_382);
or U1484 (N_1484,N_402,N_619);
nor U1485 (N_1485,N_668,N_208);
and U1486 (N_1486,N_537,N_527);
and U1487 (N_1487,N_801,N_726);
nor U1488 (N_1488,N_373,N_921);
nor U1489 (N_1489,N_87,N_212);
nor U1490 (N_1490,N_711,N_477);
and U1491 (N_1491,N_460,N_125);
or U1492 (N_1492,N_333,N_29);
nor U1493 (N_1493,N_144,N_518);
nand U1494 (N_1494,N_461,N_61);
or U1495 (N_1495,N_234,N_470);
or U1496 (N_1496,N_423,N_167);
nor U1497 (N_1497,N_849,N_546);
or U1498 (N_1498,N_943,N_722);
or U1499 (N_1499,N_606,N_436);
or U1500 (N_1500,N_862,N_187);
xor U1501 (N_1501,N_887,N_142);
and U1502 (N_1502,N_970,N_500);
or U1503 (N_1503,N_179,N_601);
and U1504 (N_1504,N_563,N_427);
nand U1505 (N_1505,N_973,N_945);
and U1506 (N_1506,N_275,N_585);
and U1507 (N_1507,N_984,N_784);
nor U1508 (N_1508,N_451,N_93);
nor U1509 (N_1509,N_622,N_127);
or U1510 (N_1510,N_401,N_14);
and U1511 (N_1511,N_657,N_925);
or U1512 (N_1512,N_861,N_291);
and U1513 (N_1513,N_485,N_224);
nand U1514 (N_1514,N_334,N_552);
or U1515 (N_1515,N_269,N_666);
nor U1516 (N_1516,N_925,N_266);
or U1517 (N_1517,N_411,N_849);
and U1518 (N_1518,N_887,N_714);
nand U1519 (N_1519,N_40,N_400);
nor U1520 (N_1520,N_681,N_516);
and U1521 (N_1521,N_857,N_438);
nand U1522 (N_1522,N_742,N_519);
xnor U1523 (N_1523,N_653,N_382);
nand U1524 (N_1524,N_739,N_480);
and U1525 (N_1525,N_787,N_656);
nor U1526 (N_1526,N_571,N_433);
nor U1527 (N_1527,N_706,N_470);
nand U1528 (N_1528,N_869,N_307);
nor U1529 (N_1529,N_755,N_592);
nand U1530 (N_1530,N_486,N_883);
xor U1531 (N_1531,N_882,N_963);
xor U1532 (N_1532,N_188,N_228);
nand U1533 (N_1533,N_355,N_528);
nand U1534 (N_1534,N_476,N_567);
xnor U1535 (N_1535,N_239,N_392);
or U1536 (N_1536,N_736,N_329);
nor U1537 (N_1537,N_717,N_989);
or U1538 (N_1538,N_279,N_529);
nand U1539 (N_1539,N_876,N_323);
or U1540 (N_1540,N_361,N_717);
or U1541 (N_1541,N_917,N_598);
nand U1542 (N_1542,N_795,N_681);
and U1543 (N_1543,N_88,N_70);
and U1544 (N_1544,N_626,N_258);
nor U1545 (N_1545,N_558,N_935);
xor U1546 (N_1546,N_379,N_112);
nor U1547 (N_1547,N_617,N_416);
and U1548 (N_1548,N_872,N_96);
nand U1549 (N_1549,N_688,N_294);
and U1550 (N_1550,N_443,N_886);
and U1551 (N_1551,N_126,N_325);
nor U1552 (N_1552,N_896,N_160);
nand U1553 (N_1553,N_798,N_694);
nor U1554 (N_1554,N_213,N_802);
nand U1555 (N_1555,N_11,N_45);
nor U1556 (N_1556,N_730,N_715);
nor U1557 (N_1557,N_227,N_532);
nor U1558 (N_1558,N_259,N_979);
xor U1559 (N_1559,N_466,N_582);
nand U1560 (N_1560,N_890,N_763);
nor U1561 (N_1561,N_15,N_475);
or U1562 (N_1562,N_862,N_402);
or U1563 (N_1563,N_479,N_88);
and U1564 (N_1564,N_823,N_109);
and U1565 (N_1565,N_758,N_426);
and U1566 (N_1566,N_733,N_543);
nand U1567 (N_1567,N_200,N_848);
and U1568 (N_1568,N_378,N_337);
or U1569 (N_1569,N_378,N_20);
nor U1570 (N_1570,N_399,N_60);
and U1571 (N_1571,N_445,N_824);
xnor U1572 (N_1572,N_871,N_32);
and U1573 (N_1573,N_812,N_415);
nor U1574 (N_1574,N_223,N_533);
nor U1575 (N_1575,N_728,N_955);
and U1576 (N_1576,N_690,N_147);
nor U1577 (N_1577,N_613,N_691);
or U1578 (N_1578,N_651,N_91);
nand U1579 (N_1579,N_460,N_398);
nand U1580 (N_1580,N_189,N_424);
nor U1581 (N_1581,N_998,N_754);
xor U1582 (N_1582,N_250,N_947);
nor U1583 (N_1583,N_966,N_139);
nor U1584 (N_1584,N_906,N_852);
nor U1585 (N_1585,N_789,N_551);
and U1586 (N_1586,N_242,N_645);
nor U1587 (N_1587,N_826,N_920);
or U1588 (N_1588,N_163,N_523);
nor U1589 (N_1589,N_521,N_953);
nand U1590 (N_1590,N_244,N_208);
xor U1591 (N_1591,N_324,N_914);
and U1592 (N_1592,N_732,N_222);
or U1593 (N_1593,N_316,N_788);
nor U1594 (N_1594,N_773,N_924);
nand U1595 (N_1595,N_762,N_793);
nand U1596 (N_1596,N_305,N_932);
nand U1597 (N_1597,N_830,N_734);
nand U1598 (N_1598,N_821,N_232);
and U1599 (N_1599,N_889,N_374);
or U1600 (N_1600,N_799,N_319);
or U1601 (N_1601,N_235,N_557);
or U1602 (N_1602,N_491,N_49);
nand U1603 (N_1603,N_85,N_79);
or U1604 (N_1604,N_795,N_984);
and U1605 (N_1605,N_761,N_222);
nor U1606 (N_1606,N_523,N_243);
and U1607 (N_1607,N_421,N_945);
and U1608 (N_1608,N_846,N_702);
or U1609 (N_1609,N_656,N_566);
or U1610 (N_1610,N_999,N_482);
nand U1611 (N_1611,N_40,N_348);
nor U1612 (N_1612,N_185,N_841);
nand U1613 (N_1613,N_876,N_952);
nand U1614 (N_1614,N_110,N_602);
and U1615 (N_1615,N_478,N_973);
or U1616 (N_1616,N_674,N_887);
and U1617 (N_1617,N_44,N_653);
or U1618 (N_1618,N_498,N_364);
or U1619 (N_1619,N_575,N_906);
nand U1620 (N_1620,N_627,N_388);
and U1621 (N_1621,N_133,N_717);
nor U1622 (N_1622,N_723,N_782);
and U1623 (N_1623,N_660,N_477);
nor U1624 (N_1624,N_573,N_286);
nand U1625 (N_1625,N_18,N_662);
nand U1626 (N_1626,N_790,N_331);
nand U1627 (N_1627,N_352,N_574);
or U1628 (N_1628,N_604,N_917);
nor U1629 (N_1629,N_833,N_973);
and U1630 (N_1630,N_662,N_273);
and U1631 (N_1631,N_82,N_80);
or U1632 (N_1632,N_729,N_560);
nand U1633 (N_1633,N_80,N_78);
or U1634 (N_1634,N_819,N_146);
nor U1635 (N_1635,N_258,N_727);
nor U1636 (N_1636,N_460,N_856);
nand U1637 (N_1637,N_868,N_545);
and U1638 (N_1638,N_663,N_530);
nor U1639 (N_1639,N_91,N_969);
nand U1640 (N_1640,N_575,N_467);
or U1641 (N_1641,N_331,N_934);
or U1642 (N_1642,N_953,N_986);
and U1643 (N_1643,N_49,N_591);
or U1644 (N_1644,N_477,N_803);
or U1645 (N_1645,N_698,N_463);
nand U1646 (N_1646,N_852,N_803);
nor U1647 (N_1647,N_472,N_372);
nor U1648 (N_1648,N_556,N_152);
nor U1649 (N_1649,N_837,N_292);
nand U1650 (N_1650,N_468,N_698);
nor U1651 (N_1651,N_266,N_130);
nor U1652 (N_1652,N_159,N_165);
or U1653 (N_1653,N_31,N_686);
and U1654 (N_1654,N_111,N_915);
and U1655 (N_1655,N_160,N_150);
or U1656 (N_1656,N_238,N_354);
and U1657 (N_1657,N_866,N_569);
and U1658 (N_1658,N_322,N_538);
nor U1659 (N_1659,N_121,N_458);
nand U1660 (N_1660,N_344,N_469);
and U1661 (N_1661,N_390,N_588);
nand U1662 (N_1662,N_63,N_9);
and U1663 (N_1663,N_596,N_766);
or U1664 (N_1664,N_109,N_516);
and U1665 (N_1665,N_725,N_810);
nor U1666 (N_1666,N_378,N_112);
and U1667 (N_1667,N_729,N_429);
nor U1668 (N_1668,N_885,N_782);
and U1669 (N_1669,N_246,N_956);
nand U1670 (N_1670,N_882,N_582);
or U1671 (N_1671,N_792,N_284);
and U1672 (N_1672,N_907,N_749);
and U1673 (N_1673,N_487,N_492);
nor U1674 (N_1674,N_73,N_766);
nor U1675 (N_1675,N_560,N_467);
or U1676 (N_1676,N_625,N_556);
and U1677 (N_1677,N_559,N_107);
nor U1678 (N_1678,N_668,N_109);
or U1679 (N_1679,N_505,N_982);
and U1680 (N_1680,N_176,N_630);
nand U1681 (N_1681,N_803,N_16);
nand U1682 (N_1682,N_372,N_174);
or U1683 (N_1683,N_526,N_185);
nor U1684 (N_1684,N_269,N_12);
or U1685 (N_1685,N_143,N_733);
nand U1686 (N_1686,N_717,N_415);
nand U1687 (N_1687,N_934,N_747);
nand U1688 (N_1688,N_508,N_425);
nand U1689 (N_1689,N_587,N_15);
nand U1690 (N_1690,N_616,N_121);
and U1691 (N_1691,N_82,N_649);
nand U1692 (N_1692,N_252,N_928);
nand U1693 (N_1693,N_991,N_632);
nor U1694 (N_1694,N_570,N_16);
or U1695 (N_1695,N_208,N_788);
and U1696 (N_1696,N_505,N_273);
or U1697 (N_1697,N_990,N_202);
or U1698 (N_1698,N_781,N_97);
or U1699 (N_1699,N_200,N_255);
and U1700 (N_1700,N_347,N_481);
or U1701 (N_1701,N_768,N_452);
or U1702 (N_1702,N_586,N_43);
xnor U1703 (N_1703,N_802,N_979);
or U1704 (N_1704,N_298,N_865);
nor U1705 (N_1705,N_340,N_598);
nor U1706 (N_1706,N_51,N_695);
or U1707 (N_1707,N_402,N_636);
nand U1708 (N_1708,N_820,N_213);
nor U1709 (N_1709,N_536,N_438);
nor U1710 (N_1710,N_351,N_981);
or U1711 (N_1711,N_414,N_779);
nand U1712 (N_1712,N_930,N_702);
nand U1713 (N_1713,N_355,N_152);
or U1714 (N_1714,N_96,N_465);
and U1715 (N_1715,N_659,N_918);
nand U1716 (N_1716,N_255,N_772);
and U1717 (N_1717,N_65,N_727);
nor U1718 (N_1718,N_579,N_856);
or U1719 (N_1719,N_816,N_888);
nor U1720 (N_1720,N_976,N_839);
or U1721 (N_1721,N_893,N_352);
and U1722 (N_1722,N_794,N_506);
and U1723 (N_1723,N_697,N_66);
nor U1724 (N_1724,N_412,N_228);
nor U1725 (N_1725,N_221,N_112);
nor U1726 (N_1726,N_525,N_507);
and U1727 (N_1727,N_169,N_273);
nor U1728 (N_1728,N_279,N_72);
or U1729 (N_1729,N_58,N_960);
nand U1730 (N_1730,N_365,N_547);
or U1731 (N_1731,N_495,N_566);
or U1732 (N_1732,N_430,N_252);
nand U1733 (N_1733,N_642,N_625);
or U1734 (N_1734,N_178,N_27);
and U1735 (N_1735,N_11,N_131);
or U1736 (N_1736,N_572,N_618);
nor U1737 (N_1737,N_681,N_950);
nand U1738 (N_1738,N_364,N_164);
nor U1739 (N_1739,N_804,N_875);
nand U1740 (N_1740,N_794,N_921);
and U1741 (N_1741,N_271,N_678);
and U1742 (N_1742,N_32,N_169);
nand U1743 (N_1743,N_613,N_219);
or U1744 (N_1744,N_653,N_1);
nor U1745 (N_1745,N_374,N_612);
and U1746 (N_1746,N_489,N_930);
and U1747 (N_1747,N_88,N_161);
nand U1748 (N_1748,N_343,N_437);
and U1749 (N_1749,N_950,N_843);
or U1750 (N_1750,N_497,N_231);
nand U1751 (N_1751,N_113,N_457);
nor U1752 (N_1752,N_157,N_342);
and U1753 (N_1753,N_356,N_205);
nand U1754 (N_1754,N_916,N_810);
nor U1755 (N_1755,N_95,N_471);
nor U1756 (N_1756,N_805,N_404);
nor U1757 (N_1757,N_151,N_751);
nor U1758 (N_1758,N_68,N_407);
or U1759 (N_1759,N_257,N_333);
or U1760 (N_1760,N_864,N_340);
and U1761 (N_1761,N_621,N_876);
or U1762 (N_1762,N_600,N_723);
and U1763 (N_1763,N_898,N_204);
nor U1764 (N_1764,N_168,N_193);
nand U1765 (N_1765,N_118,N_300);
or U1766 (N_1766,N_59,N_322);
and U1767 (N_1767,N_560,N_788);
and U1768 (N_1768,N_650,N_254);
nand U1769 (N_1769,N_828,N_767);
and U1770 (N_1770,N_43,N_832);
and U1771 (N_1771,N_609,N_992);
nand U1772 (N_1772,N_89,N_141);
or U1773 (N_1773,N_303,N_790);
or U1774 (N_1774,N_514,N_836);
or U1775 (N_1775,N_992,N_251);
or U1776 (N_1776,N_783,N_95);
nor U1777 (N_1777,N_311,N_827);
and U1778 (N_1778,N_323,N_735);
nand U1779 (N_1779,N_141,N_475);
xor U1780 (N_1780,N_669,N_199);
or U1781 (N_1781,N_160,N_764);
and U1782 (N_1782,N_914,N_41);
nand U1783 (N_1783,N_952,N_440);
xnor U1784 (N_1784,N_279,N_854);
and U1785 (N_1785,N_892,N_86);
nand U1786 (N_1786,N_731,N_433);
and U1787 (N_1787,N_932,N_407);
nor U1788 (N_1788,N_944,N_912);
or U1789 (N_1789,N_944,N_660);
nor U1790 (N_1790,N_549,N_798);
or U1791 (N_1791,N_135,N_394);
and U1792 (N_1792,N_767,N_152);
and U1793 (N_1793,N_862,N_449);
and U1794 (N_1794,N_353,N_27);
and U1795 (N_1795,N_669,N_42);
nor U1796 (N_1796,N_871,N_838);
or U1797 (N_1797,N_952,N_939);
or U1798 (N_1798,N_366,N_395);
and U1799 (N_1799,N_428,N_46);
and U1800 (N_1800,N_725,N_657);
nand U1801 (N_1801,N_420,N_619);
nor U1802 (N_1802,N_149,N_914);
xnor U1803 (N_1803,N_280,N_808);
nor U1804 (N_1804,N_189,N_236);
nor U1805 (N_1805,N_648,N_408);
or U1806 (N_1806,N_383,N_167);
nand U1807 (N_1807,N_41,N_326);
and U1808 (N_1808,N_285,N_916);
or U1809 (N_1809,N_844,N_730);
nand U1810 (N_1810,N_856,N_326);
nand U1811 (N_1811,N_884,N_546);
nand U1812 (N_1812,N_729,N_991);
nand U1813 (N_1813,N_512,N_218);
nor U1814 (N_1814,N_114,N_325);
nor U1815 (N_1815,N_618,N_323);
nor U1816 (N_1816,N_7,N_298);
and U1817 (N_1817,N_90,N_525);
or U1818 (N_1818,N_173,N_982);
nor U1819 (N_1819,N_213,N_150);
or U1820 (N_1820,N_874,N_677);
nor U1821 (N_1821,N_210,N_274);
and U1822 (N_1822,N_765,N_665);
nand U1823 (N_1823,N_109,N_176);
nand U1824 (N_1824,N_477,N_273);
nor U1825 (N_1825,N_764,N_925);
nor U1826 (N_1826,N_177,N_440);
or U1827 (N_1827,N_820,N_272);
and U1828 (N_1828,N_842,N_654);
and U1829 (N_1829,N_635,N_408);
nor U1830 (N_1830,N_17,N_534);
and U1831 (N_1831,N_379,N_524);
and U1832 (N_1832,N_933,N_234);
nand U1833 (N_1833,N_484,N_746);
nand U1834 (N_1834,N_735,N_994);
nor U1835 (N_1835,N_965,N_959);
and U1836 (N_1836,N_595,N_798);
nand U1837 (N_1837,N_845,N_202);
or U1838 (N_1838,N_951,N_978);
nor U1839 (N_1839,N_791,N_650);
nor U1840 (N_1840,N_395,N_716);
and U1841 (N_1841,N_827,N_39);
and U1842 (N_1842,N_937,N_928);
or U1843 (N_1843,N_451,N_386);
or U1844 (N_1844,N_643,N_214);
nand U1845 (N_1845,N_351,N_780);
nand U1846 (N_1846,N_225,N_746);
nor U1847 (N_1847,N_638,N_481);
nor U1848 (N_1848,N_623,N_326);
nand U1849 (N_1849,N_800,N_699);
nor U1850 (N_1850,N_238,N_90);
nor U1851 (N_1851,N_496,N_233);
or U1852 (N_1852,N_361,N_588);
and U1853 (N_1853,N_611,N_702);
nand U1854 (N_1854,N_594,N_924);
and U1855 (N_1855,N_576,N_334);
or U1856 (N_1856,N_136,N_715);
nand U1857 (N_1857,N_986,N_865);
nor U1858 (N_1858,N_470,N_903);
nor U1859 (N_1859,N_275,N_958);
nand U1860 (N_1860,N_635,N_410);
and U1861 (N_1861,N_195,N_313);
or U1862 (N_1862,N_777,N_373);
nand U1863 (N_1863,N_0,N_585);
and U1864 (N_1864,N_987,N_643);
and U1865 (N_1865,N_558,N_394);
nor U1866 (N_1866,N_125,N_764);
nand U1867 (N_1867,N_149,N_989);
or U1868 (N_1868,N_234,N_61);
or U1869 (N_1869,N_935,N_532);
nand U1870 (N_1870,N_670,N_719);
nor U1871 (N_1871,N_877,N_885);
nand U1872 (N_1872,N_142,N_153);
nand U1873 (N_1873,N_484,N_789);
nand U1874 (N_1874,N_919,N_529);
and U1875 (N_1875,N_915,N_817);
xor U1876 (N_1876,N_452,N_675);
nor U1877 (N_1877,N_55,N_557);
or U1878 (N_1878,N_529,N_208);
nor U1879 (N_1879,N_616,N_327);
nor U1880 (N_1880,N_605,N_975);
nor U1881 (N_1881,N_98,N_996);
and U1882 (N_1882,N_384,N_562);
nand U1883 (N_1883,N_75,N_977);
or U1884 (N_1884,N_751,N_173);
and U1885 (N_1885,N_294,N_968);
nand U1886 (N_1886,N_516,N_931);
and U1887 (N_1887,N_47,N_115);
nor U1888 (N_1888,N_744,N_833);
or U1889 (N_1889,N_659,N_853);
or U1890 (N_1890,N_300,N_632);
nor U1891 (N_1891,N_156,N_592);
nor U1892 (N_1892,N_662,N_51);
nor U1893 (N_1893,N_510,N_825);
or U1894 (N_1894,N_371,N_171);
nor U1895 (N_1895,N_598,N_971);
nand U1896 (N_1896,N_553,N_814);
nor U1897 (N_1897,N_769,N_193);
nor U1898 (N_1898,N_535,N_461);
nand U1899 (N_1899,N_102,N_325);
nor U1900 (N_1900,N_523,N_503);
nor U1901 (N_1901,N_216,N_406);
nor U1902 (N_1902,N_53,N_273);
and U1903 (N_1903,N_958,N_27);
nand U1904 (N_1904,N_791,N_638);
or U1905 (N_1905,N_636,N_479);
nor U1906 (N_1906,N_425,N_238);
nand U1907 (N_1907,N_924,N_633);
and U1908 (N_1908,N_583,N_164);
and U1909 (N_1909,N_427,N_887);
and U1910 (N_1910,N_504,N_707);
and U1911 (N_1911,N_410,N_807);
and U1912 (N_1912,N_780,N_386);
nor U1913 (N_1913,N_655,N_929);
and U1914 (N_1914,N_113,N_201);
nand U1915 (N_1915,N_199,N_870);
nand U1916 (N_1916,N_208,N_639);
nor U1917 (N_1917,N_415,N_964);
nand U1918 (N_1918,N_617,N_897);
and U1919 (N_1919,N_651,N_438);
and U1920 (N_1920,N_984,N_611);
nand U1921 (N_1921,N_42,N_851);
and U1922 (N_1922,N_446,N_398);
and U1923 (N_1923,N_412,N_874);
nor U1924 (N_1924,N_484,N_737);
nand U1925 (N_1925,N_956,N_41);
nor U1926 (N_1926,N_698,N_432);
or U1927 (N_1927,N_36,N_127);
nor U1928 (N_1928,N_735,N_98);
nor U1929 (N_1929,N_572,N_502);
nand U1930 (N_1930,N_666,N_647);
and U1931 (N_1931,N_748,N_913);
or U1932 (N_1932,N_955,N_180);
and U1933 (N_1933,N_607,N_157);
nand U1934 (N_1934,N_864,N_487);
or U1935 (N_1935,N_334,N_838);
nor U1936 (N_1936,N_863,N_563);
nor U1937 (N_1937,N_883,N_971);
nand U1938 (N_1938,N_553,N_204);
nor U1939 (N_1939,N_739,N_85);
nor U1940 (N_1940,N_567,N_382);
nor U1941 (N_1941,N_702,N_164);
nand U1942 (N_1942,N_509,N_595);
nor U1943 (N_1943,N_476,N_601);
nand U1944 (N_1944,N_167,N_523);
nand U1945 (N_1945,N_70,N_400);
or U1946 (N_1946,N_640,N_528);
xor U1947 (N_1947,N_801,N_838);
and U1948 (N_1948,N_817,N_818);
nand U1949 (N_1949,N_467,N_0);
nor U1950 (N_1950,N_812,N_15);
or U1951 (N_1951,N_287,N_574);
nor U1952 (N_1952,N_931,N_222);
or U1953 (N_1953,N_288,N_398);
nand U1954 (N_1954,N_713,N_696);
nand U1955 (N_1955,N_508,N_51);
or U1956 (N_1956,N_133,N_468);
nor U1957 (N_1957,N_287,N_528);
or U1958 (N_1958,N_33,N_975);
nor U1959 (N_1959,N_644,N_204);
or U1960 (N_1960,N_680,N_11);
and U1961 (N_1961,N_382,N_153);
and U1962 (N_1962,N_67,N_593);
or U1963 (N_1963,N_448,N_611);
nor U1964 (N_1964,N_230,N_164);
or U1965 (N_1965,N_496,N_615);
nor U1966 (N_1966,N_484,N_844);
nand U1967 (N_1967,N_837,N_196);
and U1968 (N_1968,N_516,N_866);
or U1969 (N_1969,N_591,N_933);
or U1970 (N_1970,N_130,N_823);
nor U1971 (N_1971,N_753,N_74);
nand U1972 (N_1972,N_377,N_148);
nand U1973 (N_1973,N_985,N_254);
or U1974 (N_1974,N_275,N_963);
nand U1975 (N_1975,N_728,N_983);
xnor U1976 (N_1976,N_24,N_17);
or U1977 (N_1977,N_972,N_560);
and U1978 (N_1978,N_711,N_844);
or U1979 (N_1979,N_925,N_747);
and U1980 (N_1980,N_539,N_41);
nand U1981 (N_1981,N_841,N_505);
or U1982 (N_1982,N_953,N_435);
or U1983 (N_1983,N_6,N_111);
or U1984 (N_1984,N_3,N_275);
and U1985 (N_1985,N_306,N_460);
and U1986 (N_1986,N_615,N_373);
nor U1987 (N_1987,N_944,N_166);
and U1988 (N_1988,N_0,N_515);
and U1989 (N_1989,N_506,N_821);
and U1990 (N_1990,N_532,N_557);
and U1991 (N_1991,N_976,N_39);
or U1992 (N_1992,N_513,N_177);
nor U1993 (N_1993,N_489,N_708);
nor U1994 (N_1994,N_669,N_738);
nor U1995 (N_1995,N_101,N_722);
or U1996 (N_1996,N_596,N_617);
or U1997 (N_1997,N_488,N_975);
and U1998 (N_1998,N_178,N_293);
and U1999 (N_1999,N_214,N_285);
xor U2000 (N_2000,N_1114,N_1612);
or U2001 (N_2001,N_1601,N_1337);
nor U2002 (N_2002,N_1435,N_1905);
nand U2003 (N_2003,N_1231,N_1668);
and U2004 (N_2004,N_1441,N_1851);
xor U2005 (N_2005,N_1780,N_1691);
nand U2006 (N_2006,N_1627,N_1932);
and U2007 (N_2007,N_1699,N_1823);
and U2008 (N_2008,N_1232,N_1297);
or U2009 (N_2009,N_1426,N_1777);
nor U2010 (N_2010,N_1855,N_1975);
and U2011 (N_2011,N_1792,N_1207);
or U2012 (N_2012,N_1951,N_1999);
and U2013 (N_2013,N_1985,N_1968);
or U2014 (N_2014,N_1836,N_1588);
or U2015 (N_2015,N_1863,N_1814);
nand U2016 (N_2016,N_1468,N_1853);
nand U2017 (N_2017,N_1872,N_1533);
nor U2018 (N_2018,N_1950,N_1742);
or U2019 (N_2019,N_1779,N_1642);
nor U2020 (N_2020,N_1751,N_1469);
nand U2021 (N_2021,N_1040,N_1037);
nand U2022 (N_2022,N_1952,N_1555);
and U2023 (N_2023,N_1586,N_1173);
nand U2024 (N_2024,N_1894,N_1963);
and U2025 (N_2025,N_1225,N_1419);
and U2026 (N_2026,N_1665,N_1883);
and U2027 (N_2027,N_1778,N_1875);
and U2028 (N_2028,N_1375,N_1511);
or U2029 (N_2029,N_1697,N_1657);
nand U2030 (N_2030,N_1947,N_1614);
or U2031 (N_2031,N_1721,N_1577);
or U2032 (N_2032,N_1408,N_1113);
or U2033 (N_2033,N_1867,N_1443);
and U2034 (N_2034,N_1766,N_1467);
nor U2035 (N_2035,N_1007,N_1756);
nand U2036 (N_2036,N_1729,N_1128);
and U2037 (N_2037,N_1322,N_1103);
and U2038 (N_2038,N_1724,N_1786);
or U2039 (N_2039,N_1401,N_1092);
nand U2040 (N_2040,N_1138,N_1366);
nor U2041 (N_2041,N_1785,N_1791);
nand U2042 (N_2042,N_1743,N_1255);
nand U2043 (N_2043,N_1915,N_1198);
nor U2044 (N_2044,N_1827,N_1545);
or U2045 (N_2045,N_1172,N_1871);
nand U2046 (N_2046,N_1678,N_1118);
or U2047 (N_2047,N_1296,N_1439);
nand U2048 (N_2048,N_1147,N_1378);
nor U2049 (N_2049,N_1129,N_1196);
or U2050 (N_2050,N_1325,N_1881);
nor U2051 (N_2051,N_1587,N_1150);
nor U2052 (N_2052,N_1212,N_1796);
and U2053 (N_2053,N_1893,N_1694);
or U2054 (N_2054,N_1794,N_1531);
xor U2055 (N_2055,N_1406,N_1495);
nor U2056 (N_2056,N_1824,N_1575);
or U2057 (N_2057,N_1527,N_1395);
nor U2058 (N_2058,N_1219,N_1059);
and U2059 (N_2059,N_1015,N_1480);
nand U2060 (N_2060,N_1866,N_1681);
nand U2061 (N_2061,N_1611,N_1625);
or U2062 (N_2062,N_1083,N_1935);
or U2063 (N_2063,N_1084,N_1264);
nand U2064 (N_2064,N_1068,N_1978);
and U2065 (N_2065,N_1502,N_1206);
and U2066 (N_2066,N_1943,N_1290);
and U2067 (N_2067,N_1318,N_1649);
nand U2068 (N_2068,N_1339,N_1095);
nor U2069 (N_2069,N_1541,N_1159);
nand U2070 (N_2070,N_1116,N_1921);
nor U2071 (N_2071,N_1217,N_1433);
and U2072 (N_2072,N_1331,N_1201);
nor U2073 (N_2073,N_1885,N_1715);
xnor U2074 (N_2074,N_1271,N_1088);
or U2075 (N_2075,N_1091,N_1039);
nand U2076 (N_2076,N_1817,N_1042);
or U2077 (N_2077,N_1834,N_1631);
or U2078 (N_2078,N_1880,N_1804);
nand U2079 (N_2079,N_1209,N_1122);
or U2080 (N_2080,N_1720,N_1690);
nand U2081 (N_2081,N_1282,N_1162);
or U2082 (N_2082,N_1214,N_1400);
xor U2083 (N_2083,N_1187,N_1598);
nor U2084 (N_2084,N_1213,N_1898);
nor U2085 (N_2085,N_1486,N_1224);
nor U2086 (N_2086,N_1765,N_1987);
nor U2087 (N_2087,N_1416,N_1578);
and U2088 (N_2088,N_1360,N_1491);
nor U2089 (N_2089,N_1452,N_1537);
nand U2090 (N_2090,N_1549,N_1035);
nor U2091 (N_2091,N_1910,N_1284);
or U2092 (N_2092,N_1576,N_1662);
nand U2093 (N_2093,N_1041,N_1470);
or U2094 (N_2094,N_1144,N_1516);
nand U2095 (N_2095,N_1613,N_1574);
nand U2096 (N_2096,N_1350,N_1816);
nor U2097 (N_2097,N_1936,N_1859);
or U2098 (N_2098,N_1292,N_1746);
nor U2099 (N_2099,N_1566,N_1161);
or U2100 (N_2100,N_1979,N_1542);
or U2101 (N_2101,N_1903,N_1228);
or U2102 (N_2102,N_1908,N_1781);
nor U2103 (N_2103,N_1425,N_1391);
or U2104 (N_2104,N_1009,N_1655);
nor U2105 (N_2105,N_1539,N_1496);
or U2106 (N_2106,N_1688,N_1807);
or U2107 (N_2107,N_1929,N_1683);
xnor U2108 (N_2108,N_1772,N_1267);
nor U2109 (N_2109,N_1820,N_1553);
and U2110 (N_2110,N_1479,N_1356);
or U2111 (N_2111,N_1359,N_1074);
nor U2112 (N_2112,N_1775,N_1347);
or U2113 (N_2113,N_1221,N_1078);
and U2114 (N_2114,N_1503,N_1131);
or U2115 (N_2115,N_1167,N_1476);
nand U2116 (N_2116,N_1051,N_1719);
and U2117 (N_2117,N_1022,N_1410);
nand U2118 (N_2118,N_1671,N_1014);
and U2119 (N_2119,N_1760,N_1434);
xnor U2120 (N_2120,N_1517,N_1702);
nor U2121 (N_2121,N_1818,N_1660);
nor U2122 (N_2122,N_1460,N_1392);
and U2123 (N_2123,N_1199,N_1646);
nor U2124 (N_2124,N_1044,N_1973);
and U2125 (N_2125,N_1876,N_1504);
and U2126 (N_2126,N_1399,N_1329);
or U2127 (N_2127,N_1146,N_1530);
or U2128 (N_2128,N_1847,N_1016);
or U2129 (N_2129,N_1311,N_1819);
or U2130 (N_2130,N_1062,N_1269);
nor U2131 (N_2131,N_1286,N_1970);
nand U2132 (N_2132,N_1618,N_1226);
and U2133 (N_2133,N_1349,N_1327);
and U2134 (N_2134,N_1251,N_1056);
nor U2135 (N_2135,N_1080,N_1104);
and U2136 (N_2136,N_1011,N_1250);
and U2137 (N_2137,N_1003,N_1108);
nand U2138 (N_2138,N_1239,N_1698);
or U2139 (N_2139,N_1802,N_1376);
and U2140 (N_2140,N_1237,N_1430);
or U2141 (N_2141,N_1557,N_1570);
and U2142 (N_2142,N_1965,N_1183);
nand U2143 (N_2143,N_1572,N_1732);
nand U2144 (N_2144,N_1205,N_1386);
nand U2145 (N_2145,N_1764,N_1933);
nor U2146 (N_2146,N_1632,N_1143);
or U2147 (N_2147,N_1809,N_1073);
and U2148 (N_2148,N_1909,N_1379);
nor U2149 (N_2149,N_1033,N_1106);
nand U2150 (N_2150,N_1606,N_1730);
or U2151 (N_2151,N_1523,N_1076);
or U2152 (N_2152,N_1639,N_1925);
or U2153 (N_2153,N_1256,N_1299);
or U2154 (N_2154,N_1004,N_1774);
and U2155 (N_2155,N_1930,N_1208);
or U2156 (N_2156,N_1650,N_1442);
xnor U2157 (N_2157,N_1998,N_1628);
nand U2158 (N_2158,N_1494,N_1195);
nor U2159 (N_2159,N_1302,N_1918);
nand U2160 (N_2160,N_1216,N_1077);
nor U2161 (N_2161,N_1609,N_1808);
and U2162 (N_2162,N_1457,N_1990);
and U2163 (N_2163,N_1253,N_1543);
or U2164 (N_2164,N_1850,N_1669);
nor U2165 (N_2165,N_1873,N_1380);
nand U2166 (N_2166,N_1954,N_1584);
nor U2167 (N_2167,N_1300,N_1920);
nor U2168 (N_2168,N_1127,N_1418);
nand U2169 (N_2169,N_1244,N_1787);
or U2170 (N_2170,N_1320,N_1538);
and U2171 (N_2171,N_1346,N_1994);
or U2172 (N_2172,N_1899,N_1629);
or U2173 (N_2173,N_1110,N_1450);
nand U2174 (N_2174,N_1126,N_1397);
and U2175 (N_2175,N_1718,N_1362);
or U2176 (N_2176,N_1653,N_1617);
or U2177 (N_2177,N_1101,N_1886);
nor U2178 (N_2178,N_1884,N_1837);
nor U2179 (N_2179,N_1483,N_1953);
or U2180 (N_2180,N_1013,N_1634);
and U2181 (N_2181,N_1770,N_1102);
and U2182 (N_2182,N_1831,N_1864);
nor U2183 (N_2183,N_1343,N_1687);
and U2184 (N_2184,N_1069,N_1274);
or U2185 (N_2185,N_1050,N_1197);
and U2186 (N_2186,N_1500,N_1165);
and U2187 (N_2187,N_1365,N_1674);
nor U2188 (N_2188,N_1497,N_1142);
nand U2189 (N_2189,N_1405,N_1090);
nor U2190 (N_2190,N_1957,N_1473);
and U2191 (N_2191,N_1793,N_1803);
and U2192 (N_2192,N_1860,N_1471);
nor U2193 (N_2193,N_1745,N_1123);
nand U2194 (N_2194,N_1508,N_1693);
or U2195 (N_2195,N_1506,N_1229);
nor U2196 (N_2196,N_1558,N_1633);
nand U2197 (N_2197,N_1524,N_1319);
and U2198 (N_2198,N_1623,N_1352);
or U2199 (N_2199,N_1171,N_1821);
or U2200 (N_2200,N_1755,N_1326);
or U2201 (N_2201,N_1348,N_1654);
and U2202 (N_2202,N_1342,N_1249);
nor U2203 (N_2203,N_1067,N_1374);
nor U2204 (N_2204,N_1891,N_1499);
and U2205 (N_2205,N_1806,N_1321);
and U2206 (N_2206,N_1676,N_1590);
nand U2207 (N_2207,N_1045,N_1283);
nand U2208 (N_2208,N_1227,N_1130);
or U2209 (N_2209,N_1600,N_1436);
or U2210 (N_2210,N_1140,N_1521);
nand U2211 (N_2211,N_1338,N_1928);
or U2212 (N_2212,N_1712,N_1157);
nand U2213 (N_2213,N_1595,N_1801);
or U2214 (N_2214,N_1394,N_1281);
or U2215 (N_2215,N_1409,N_1310);
and U2216 (N_2216,N_1423,N_1520);
nor U2217 (N_2217,N_1309,N_1235);
and U2218 (N_2218,N_1757,N_1661);
nand U2219 (N_2219,N_1429,N_1017);
and U2220 (N_2220,N_1547,N_1275);
nor U2221 (N_2221,N_1179,N_1843);
nor U2222 (N_2222,N_1288,N_1163);
nand U2223 (N_2223,N_1710,N_1064);
nor U2224 (N_2224,N_1189,N_1752);
nor U2225 (N_2225,N_1663,N_1308);
or U2226 (N_2226,N_1381,N_1939);
and U2227 (N_2227,N_1519,N_1768);
and U2228 (N_2228,N_1484,N_1204);
nand U2229 (N_2229,N_1548,N_1581);
and U2230 (N_2230,N_1280,N_1602);
or U2231 (N_2231,N_1301,N_1658);
and U2232 (N_2232,N_1030,N_1941);
and U2233 (N_2233,N_1677,N_1830);
nor U2234 (N_2234,N_1278,N_1420);
and U2235 (N_2235,N_1166,N_1304);
or U2236 (N_2236,N_1048,N_1431);
nand U2237 (N_2237,N_1713,N_1825);
nor U2238 (N_2238,N_1052,N_1098);
and U2239 (N_2239,N_1822,N_1544);
nor U2240 (N_2240,N_1703,N_1701);
nand U2241 (N_2241,N_1265,N_1367);
and U2242 (N_2242,N_1481,N_1262);
or U2243 (N_2243,N_1324,N_1858);
or U2244 (N_2244,N_1323,N_1332);
nand U2245 (N_2245,N_1466,N_1313);
or U2246 (N_2246,N_1733,N_1285);
or U2247 (N_2247,N_1705,N_1276);
nand U2248 (N_2248,N_1983,N_1513);
nand U2249 (N_2249,N_1370,N_1879);
nand U2250 (N_2250,N_1507,N_1134);
nand U2251 (N_2251,N_1238,N_1967);
nor U2252 (N_2252,N_1289,N_1389);
or U2253 (N_2253,N_1946,N_1961);
and U2254 (N_2254,N_1622,N_1877);
or U2255 (N_2255,N_1222,N_1053);
nor U2256 (N_2256,N_1620,N_1248);
nor U2257 (N_2257,N_1695,N_1707);
nand U2258 (N_2258,N_1252,N_1782);
or U2259 (N_2259,N_1826,N_1445);
or U2260 (N_2260,N_1031,N_1449);
nand U2261 (N_2261,N_1741,N_1036);
or U2262 (N_2262,N_1767,N_1972);
and U2263 (N_2263,N_1372,N_1734);
nor U2264 (N_2264,N_1635,N_1268);
nor U2265 (N_2265,N_1330,N_1675);
nand U2266 (N_2266,N_1021,N_1956);
nand U2267 (N_2267,N_1902,N_1177);
and U2268 (N_2268,N_1192,N_1759);
or U2269 (N_2269,N_1552,N_1740);
nand U2270 (N_2270,N_1242,N_1852);
and U2271 (N_2271,N_1096,N_1156);
nor U2272 (N_2272,N_1846,N_1363);
or U2273 (N_2273,N_1125,N_1492);
nand U2274 (N_2274,N_1763,N_1986);
nand U2275 (N_2275,N_1266,N_1058);
nor U2276 (N_2276,N_1636,N_1498);
and U2277 (N_2277,N_1916,N_1462);
or U2278 (N_2278,N_1841,N_1605);
and U2279 (N_2279,N_1582,N_1413);
or U2280 (N_2280,N_1505,N_1085);
or U2281 (N_2281,N_1133,N_1341);
nor U2282 (N_2282,N_1753,N_1132);
and U2283 (N_2283,N_1805,N_1453);
nand U2284 (N_2284,N_1458,N_1455);
nand U2285 (N_2285,N_1291,N_1569);
and U2286 (N_2286,N_1861,N_1148);
nor U2287 (N_2287,N_1120,N_1888);
and U2288 (N_2288,N_1383,N_1783);
and U2289 (N_2289,N_1551,N_1568);
or U2290 (N_2290,N_1529,N_1263);
or U2291 (N_2291,N_1038,N_1155);
nand U2292 (N_2292,N_1336,N_1949);
nand U2293 (N_2293,N_1560,N_1641);
nor U2294 (N_2294,N_1023,N_1561);
xnor U2295 (N_2295,N_1440,N_1964);
or U2296 (N_2296,N_1727,N_1119);
nor U2297 (N_2297,N_1996,N_1942);
and U2298 (N_2298,N_1739,N_1333);
or U2299 (N_2299,N_1000,N_1488);
nor U2300 (N_2300,N_1184,N_1554);
nor U2301 (N_2301,N_1682,N_1234);
nor U2302 (N_2302,N_1046,N_1984);
nand U2303 (N_2303,N_1997,N_1514);
or U2304 (N_2304,N_1960,N_1644);
or U2305 (N_2305,N_1738,N_1924);
nor U2306 (N_2306,N_1482,N_1896);
and U2307 (N_2307,N_1354,N_1684);
nand U2308 (N_2308,N_1556,N_1927);
nand U2309 (N_2309,N_1828,N_1233);
or U2310 (N_2310,N_1246,N_1857);
nor U2311 (N_2311,N_1082,N_1432);
nand U2312 (N_2312,N_1917,N_1788);
and U2313 (N_2313,N_1061,N_1874);
nand U2314 (N_2314,N_1215,N_1428);
nor U2315 (N_2315,N_1567,N_1312);
nand U2316 (N_2316,N_1931,N_1240);
nand U2317 (N_2317,N_1414,N_1573);
nor U2318 (N_2318,N_1382,N_1464);
and U2319 (N_2319,N_1594,N_1049);
and U2320 (N_2320,N_1670,N_1758);
nand U2321 (N_2321,N_1451,N_1427);
and U2322 (N_2322,N_1008,N_1737);
xnor U2323 (N_2323,N_1944,N_1616);
and U2324 (N_2324,N_1700,N_1535);
nor U2325 (N_2325,N_1328,N_1865);
nor U2326 (N_2326,N_1396,N_1948);
nor U2327 (N_2327,N_1735,N_1995);
and U2328 (N_2328,N_1136,N_1223);
and U2329 (N_2329,N_1200,N_1878);
or U2330 (N_2330,N_1368,N_1769);
and U2331 (N_2331,N_1316,N_1579);
nand U2332 (N_2332,N_1066,N_1991);
nor U2333 (N_2333,N_1461,N_1006);
or U2334 (N_2334,N_1174,N_1728);
nor U2335 (N_2335,N_1647,N_1518);
and U2336 (N_2336,N_1603,N_1478);
nand U2337 (N_2337,N_1487,N_1923);
nor U2338 (N_2338,N_1937,N_1868);
nand U2339 (N_2339,N_1247,N_1640);
and U2340 (N_2340,N_1314,N_1388);
or U2341 (N_2341,N_1387,N_1357);
nor U2342 (N_2342,N_1364,N_1977);
nand U2343 (N_2343,N_1797,N_1904);
nand U2344 (N_2344,N_1043,N_1417);
nor U2345 (N_2345,N_1010,N_1257);
nor U2346 (N_2346,N_1532,N_1709);
nand U2347 (N_2347,N_1412,N_1648);
xor U2348 (N_2348,N_1254,N_1562);
and U2349 (N_2349,N_1093,N_1107);
or U2350 (N_2350,N_1914,N_1369);
nand U2351 (N_2351,N_1024,N_1344);
nand U2352 (N_2352,N_1186,N_1835);
or U2353 (N_2353,N_1444,N_1351);
and U2354 (N_2354,N_1610,N_1962);
and U2355 (N_2355,N_1597,N_1164);
or U2356 (N_2356,N_1559,N_1969);
nand U2357 (N_2357,N_1465,N_1815);
and U2358 (N_2358,N_1811,N_1832);
and U2359 (N_2359,N_1459,N_1563);
or U2360 (N_2360,N_1355,N_1564);
and U2361 (N_2361,N_1111,N_1725);
or U2362 (N_2362,N_1722,N_1882);
and U2363 (N_2363,N_1001,N_1190);
or U2364 (N_2364,N_1895,N_1749);
or U2365 (N_2365,N_1900,N_1075);
or U2366 (N_2366,N_1202,N_1989);
nand U2367 (N_2367,N_1672,N_1976);
and U2368 (N_2368,N_1591,N_1870);
or U2369 (N_2369,N_1153,N_1345);
or U2370 (N_2370,N_1272,N_1081);
and U2371 (N_2371,N_1447,N_1813);
and U2372 (N_2372,N_1180,N_1060);
and U2373 (N_2373,N_1993,N_1773);
or U2374 (N_2374,N_1515,N_1536);
or U2375 (N_2375,N_1057,N_1334);
and U2376 (N_2376,N_1974,N_1005);
nor U2377 (N_2377,N_1901,N_1844);
nor U2378 (N_2378,N_1711,N_1958);
nor U2379 (N_2379,N_1454,N_1176);
or U2380 (N_2380,N_1175,N_1747);
or U2381 (N_2381,N_1981,N_1079);
or U2382 (N_2382,N_1070,N_1135);
and U2383 (N_2383,N_1938,N_1437);
or U2384 (N_2384,N_1714,N_1404);
or U2385 (N_2385,N_1708,N_1696);
nand U2386 (N_2386,N_1589,N_1643);
or U2387 (N_2387,N_1784,N_1615);
nor U2388 (N_2388,N_1795,N_1160);
nor U2389 (N_2389,N_1913,N_1790);
nor U2390 (N_2390,N_1762,N_1115);
or U2391 (N_2391,N_1194,N_1121);
nand U2392 (N_2392,N_1446,N_1854);
nor U2393 (N_2393,N_1055,N_1522);
xor U2394 (N_2394,N_1424,N_1361);
and U2395 (N_2395,N_1243,N_1018);
and U2396 (N_2396,N_1306,N_1407);
or U2397 (N_2397,N_1034,N_1210);
nor U2398 (N_2398,N_1384,N_1472);
nor U2399 (N_2399,N_1029,N_1385);
and U2400 (N_2400,N_1869,N_1493);
nor U2401 (N_2401,N_1652,N_1020);
nor U2402 (N_2402,N_1621,N_1945);
and U2403 (N_2403,N_1245,N_1151);
nand U2404 (N_2404,N_1393,N_1731);
nand U2405 (N_2405,N_1897,N_1754);
nor U2406 (N_2406,N_1580,N_1203);
nand U2407 (N_2407,N_1664,N_1086);
nand U2408 (N_2408,N_1220,N_1087);
and U2409 (N_2409,N_1028,N_1812);
xnor U2410 (N_2410,N_1012,N_1181);
nor U2411 (N_2411,N_1099,N_1071);
nand U2412 (N_2412,N_1659,N_1550);
nand U2413 (N_2413,N_1421,N_1889);
and U2414 (N_2414,N_1353,N_1525);
or U2415 (N_2415,N_1630,N_1260);
nand U2416 (N_2416,N_1706,N_1565);
or U2417 (N_2417,N_1112,N_1032);
or U2418 (N_2418,N_1117,N_1526);
nor U2419 (N_2419,N_1475,N_1840);
nor U2420 (N_2420,N_1571,N_1377);
nor U2421 (N_2421,N_1211,N_1298);
nand U2422 (N_2422,N_1152,N_1448);
and U2423 (N_2423,N_1154,N_1856);
nand U2424 (N_2424,N_1054,N_1063);
nor U2425 (N_2425,N_1604,N_1089);
nand U2426 (N_2426,N_1411,N_1849);
nor U2427 (N_2427,N_1340,N_1839);
nor U2428 (N_2428,N_1922,N_1149);
nor U2429 (N_2429,N_1025,N_1185);
nor U2430 (N_2430,N_1065,N_1277);
nor U2431 (N_2431,N_1358,N_1403);
and U2432 (N_2432,N_1887,N_1259);
nor U2433 (N_2433,N_1188,N_1907);
and U2434 (N_2434,N_1477,N_1305);
and U2435 (N_2435,N_1295,N_1637);
nand U2436 (N_2436,N_1270,N_1799);
and U2437 (N_2437,N_1145,N_1940);
nand U2438 (N_2438,N_1287,N_1842);
and U2439 (N_2439,N_1002,N_1170);
nor U2440 (N_2440,N_1982,N_1988);
and U2441 (N_2441,N_1667,N_1047);
nand U2442 (N_2442,N_1726,N_1638);
nor U2443 (N_2443,N_1934,N_1456);
and U2444 (N_2444,N_1438,N_1335);
nand U2445 (N_2445,N_1137,N_1800);
nand U2446 (N_2446,N_1890,N_1748);
and U2447 (N_2447,N_1510,N_1651);
or U2448 (N_2448,N_1191,N_1810);
or U2449 (N_2449,N_1097,N_1390);
nor U2450 (N_2450,N_1303,N_1273);
and U2451 (N_2451,N_1169,N_1026);
or U2452 (N_2452,N_1489,N_1178);
nor U2453 (N_2453,N_1307,N_1463);
or U2454 (N_2454,N_1966,N_1750);
or U2455 (N_2455,N_1656,N_1789);
and U2456 (N_2456,N_1230,N_1723);
and U2457 (N_2457,N_1680,N_1992);
nand U2458 (N_2458,N_1980,N_1892);
nand U2459 (N_2459,N_1534,N_1139);
and U2460 (N_2460,N_1607,N_1624);
nor U2461 (N_2461,N_1485,N_1838);
or U2462 (N_2462,N_1124,N_1645);
nor U2463 (N_2463,N_1704,N_1906);
nand U2464 (N_2464,N_1919,N_1258);
nor U2465 (N_2465,N_1158,N_1744);
or U2466 (N_2466,N_1736,N_1692);
xor U2467 (N_2467,N_1241,N_1862);
nor U2468 (N_2468,N_1402,N_1168);
nand U2469 (N_2469,N_1182,N_1072);
and U2470 (N_2470,N_1685,N_1105);
or U2471 (N_2471,N_1501,N_1761);
nand U2472 (N_2472,N_1679,N_1673);
and U2473 (N_2473,N_1512,N_1422);
nand U2474 (N_2474,N_1771,N_1717);
nor U2475 (N_2475,N_1592,N_1619);
nor U2476 (N_2476,N_1798,N_1596);
nor U2477 (N_2477,N_1094,N_1261);
nand U2478 (N_2478,N_1315,N_1141);
nand U2479 (N_2479,N_1279,N_1911);
nor U2480 (N_2480,N_1218,N_1626);
nor U2481 (N_2481,N_1528,N_1509);
nor U2482 (N_2482,N_1608,N_1912);
and U2483 (N_2483,N_1415,N_1474);
nand U2484 (N_2484,N_1686,N_1716);
or U2485 (N_2485,N_1845,N_1317);
nand U2486 (N_2486,N_1593,N_1546);
nand U2487 (N_2487,N_1585,N_1583);
nand U2488 (N_2488,N_1236,N_1193);
nor U2489 (N_2489,N_1100,N_1829);
nor U2490 (N_2490,N_1689,N_1833);
and U2491 (N_2491,N_1540,N_1027);
and U2492 (N_2492,N_1848,N_1373);
or U2493 (N_2493,N_1955,N_1971);
nand U2494 (N_2494,N_1371,N_1926);
and U2495 (N_2495,N_1666,N_1490);
or U2496 (N_2496,N_1959,N_1293);
nand U2497 (N_2497,N_1294,N_1109);
and U2498 (N_2498,N_1019,N_1599);
nand U2499 (N_2499,N_1776,N_1398);
nand U2500 (N_2500,N_1832,N_1953);
and U2501 (N_2501,N_1586,N_1064);
or U2502 (N_2502,N_1768,N_1161);
or U2503 (N_2503,N_1785,N_1763);
nand U2504 (N_2504,N_1081,N_1222);
or U2505 (N_2505,N_1917,N_1119);
or U2506 (N_2506,N_1316,N_1733);
nand U2507 (N_2507,N_1546,N_1556);
and U2508 (N_2508,N_1162,N_1713);
nor U2509 (N_2509,N_1777,N_1601);
nand U2510 (N_2510,N_1640,N_1900);
nand U2511 (N_2511,N_1010,N_1119);
nand U2512 (N_2512,N_1673,N_1036);
and U2513 (N_2513,N_1055,N_1007);
nor U2514 (N_2514,N_1228,N_1581);
nand U2515 (N_2515,N_1577,N_1181);
or U2516 (N_2516,N_1143,N_1982);
and U2517 (N_2517,N_1372,N_1443);
nor U2518 (N_2518,N_1280,N_1053);
and U2519 (N_2519,N_1950,N_1576);
or U2520 (N_2520,N_1237,N_1667);
or U2521 (N_2521,N_1688,N_1076);
nand U2522 (N_2522,N_1542,N_1279);
and U2523 (N_2523,N_1284,N_1166);
and U2524 (N_2524,N_1558,N_1234);
or U2525 (N_2525,N_1635,N_1869);
and U2526 (N_2526,N_1140,N_1703);
and U2527 (N_2527,N_1343,N_1721);
nand U2528 (N_2528,N_1547,N_1610);
nor U2529 (N_2529,N_1307,N_1727);
and U2530 (N_2530,N_1379,N_1645);
or U2531 (N_2531,N_1662,N_1422);
nor U2532 (N_2532,N_1123,N_1553);
or U2533 (N_2533,N_1688,N_1279);
nor U2534 (N_2534,N_1194,N_1711);
and U2535 (N_2535,N_1009,N_1777);
or U2536 (N_2536,N_1064,N_1013);
nor U2537 (N_2537,N_1488,N_1436);
or U2538 (N_2538,N_1442,N_1032);
and U2539 (N_2539,N_1324,N_1191);
nor U2540 (N_2540,N_1897,N_1243);
nand U2541 (N_2541,N_1023,N_1551);
and U2542 (N_2542,N_1171,N_1303);
nand U2543 (N_2543,N_1308,N_1883);
nor U2544 (N_2544,N_1349,N_1223);
nand U2545 (N_2545,N_1124,N_1753);
or U2546 (N_2546,N_1286,N_1249);
and U2547 (N_2547,N_1767,N_1768);
and U2548 (N_2548,N_1818,N_1601);
and U2549 (N_2549,N_1874,N_1677);
and U2550 (N_2550,N_1887,N_1894);
or U2551 (N_2551,N_1066,N_1235);
nor U2552 (N_2552,N_1715,N_1801);
nand U2553 (N_2553,N_1807,N_1003);
or U2554 (N_2554,N_1292,N_1583);
and U2555 (N_2555,N_1490,N_1259);
or U2556 (N_2556,N_1038,N_1817);
and U2557 (N_2557,N_1105,N_1194);
nor U2558 (N_2558,N_1731,N_1788);
and U2559 (N_2559,N_1686,N_1693);
or U2560 (N_2560,N_1191,N_1600);
nand U2561 (N_2561,N_1341,N_1689);
xor U2562 (N_2562,N_1618,N_1927);
nand U2563 (N_2563,N_1050,N_1154);
and U2564 (N_2564,N_1415,N_1977);
nand U2565 (N_2565,N_1743,N_1338);
nor U2566 (N_2566,N_1548,N_1041);
nand U2567 (N_2567,N_1635,N_1066);
nand U2568 (N_2568,N_1630,N_1311);
nor U2569 (N_2569,N_1478,N_1175);
and U2570 (N_2570,N_1448,N_1386);
or U2571 (N_2571,N_1299,N_1661);
nor U2572 (N_2572,N_1053,N_1872);
nand U2573 (N_2573,N_1965,N_1999);
and U2574 (N_2574,N_1988,N_1085);
nand U2575 (N_2575,N_1006,N_1800);
nand U2576 (N_2576,N_1534,N_1747);
nor U2577 (N_2577,N_1905,N_1743);
nor U2578 (N_2578,N_1982,N_1839);
or U2579 (N_2579,N_1873,N_1541);
nand U2580 (N_2580,N_1768,N_1081);
and U2581 (N_2581,N_1603,N_1789);
nor U2582 (N_2582,N_1351,N_1067);
or U2583 (N_2583,N_1411,N_1183);
and U2584 (N_2584,N_1084,N_1667);
and U2585 (N_2585,N_1437,N_1289);
and U2586 (N_2586,N_1563,N_1002);
and U2587 (N_2587,N_1112,N_1930);
nand U2588 (N_2588,N_1042,N_1613);
and U2589 (N_2589,N_1452,N_1636);
or U2590 (N_2590,N_1488,N_1175);
and U2591 (N_2591,N_1645,N_1727);
nor U2592 (N_2592,N_1967,N_1448);
nand U2593 (N_2593,N_1785,N_1792);
nand U2594 (N_2594,N_1068,N_1966);
and U2595 (N_2595,N_1065,N_1652);
and U2596 (N_2596,N_1877,N_1608);
or U2597 (N_2597,N_1558,N_1999);
or U2598 (N_2598,N_1756,N_1003);
nor U2599 (N_2599,N_1215,N_1058);
and U2600 (N_2600,N_1529,N_1362);
nor U2601 (N_2601,N_1958,N_1020);
nand U2602 (N_2602,N_1537,N_1908);
or U2603 (N_2603,N_1379,N_1957);
or U2604 (N_2604,N_1938,N_1469);
and U2605 (N_2605,N_1272,N_1403);
or U2606 (N_2606,N_1759,N_1807);
nor U2607 (N_2607,N_1277,N_1409);
nand U2608 (N_2608,N_1074,N_1307);
nor U2609 (N_2609,N_1674,N_1837);
or U2610 (N_2610,N_1318,N_1292);
or U2611 (N_2611,N_1787,N_1495);
or U2612 (N_2612,N_1385,N_1602);
or U2613 (N_2613,N_1227,N_1635);
or U2614 (N_2614,N_1245,N_1681);
nand U2615 (N_2615,N_1733,N_1290);
nand U2616 (N_2616,N_1396,N_1573);
nor U2617 (N_2617,N_1514,N_1327);
nand U2618 (N_2618,N_1179,N_1055);
nand U2619 (N_2619,N_1522,N_1610);
or U2620 (N_2620,N_1614,N_1517);
and U2621 (N_2621,N_1216,N_1092);
nor U2622 (N_2622,N_1183,N_1896);
or U2623 (N_2623,N_1446,N_1028);
and U2624 (N_2624,N_1395,N_1467);
nand U2625 (N_2625,N_1379,N_1500);
nor U2626 (N_2626,N_1278,N_1140);
nand U2627 (N_2627,N_1678,N_1720);
nor U2628 (N_2628,N_1215,N_1124);
and U2629 (N_2629,N_1674,N_1392);
nand U2630 (N_2630,N_1493,N_1879);
nor U2631 (N_2631,N_1943,N_1389);
xor U2632 (N_2632,N_1766,N_1744);
or U2633 (N_2633,N_1673,N_1360);
and U2634 (N_2634,N_1488,N_1969);
or U2635 (N_2635,N_1119,N_1334);
and U2636 (N_2636,N_1614,N_1705);
nor U2637 (N_2637,N_1082,N_1918);
nand U2638 (N_2638,N_1739,N_1565);
and U2639 (N_2639,N_1547,N_1860);
nor U2640 (N_2640,N_1002,N_1355);
and U2641 (N_2641,N_1218,N_1616);
or U2642 (N_2642,N_1876,N_1473);
nand U2643 (N_2643,N_1961,N_1891);
nand U2644 (N_2644,N_1041,N_1326);
or U2645 (N_2645,N_1102,N_1211);
or U2646 (N_2646,N_1146,N_1961);
nand U2647 (N_2647,N_1061,N_1405);
or U2648 (N_2648,N_1082,N_1455);
or U2649 (N_2649,N_1833,N_1811);
or U2650 (N_2650,N_1719,N_1874);
and U2651 (N_2651,N_1099,N_1542);
and U2652 (N_2652,N_1000,N_1659);
or U2653 (N_2653,N_1754,N_1025);
and U2654 (N_2654,N_1033,N_1306);
and U2655 (N_2655,N_1312,N_1957);
or U2656 (N_2656,N_1448,N_1413);
nor U2657 (N_2657,N_1917,N_1612);
and U2658 (N_2658,N_1642,N_1386);
nor U2659 (N_2659,N_1810,N_1724);
nand U2660 (N_2660,N_1427,N_1129);
and U2661 (N_2661,N_1103,N_1848);
nand U2662 (N_2662,N_1525,N_1161);
nand U2663 (N_2663,N_1166,N_1823);
nand U2664 (N_2664,N_1153,N_1629);
and U2665 (N_2665,N_1687,N_1228);
nor U2666 (N_2666,N_1310,N_1283);
xor U2667 (N_2667,N_1971,N_1559);
and U2668 (N_2668,N_1317,N_1739);
and U2669 (N_2669,N_1388,N_1327);
or U2670 (N_2670,N_1326,N_1982);
and U2671 (N_2671,N_1590,N_1374);
nand U2672 (N_2672,N_1931,N_1983);
and U2673 (N_2673,N_1318,N_1687);
and U2674 (N_2674,N_1272,N_1638);
nand U2675 (N_2675,N_1020,N_1031);
nand U2676 (N_2676,N_1157,N_1524);
or U2677 (N_2677,N_1918,N_1107);
nor U2678 (N_2678,N_1915,N_1944);
or U2679 (N_2679,N_1048,N_1251);
and U2680 (N_2680,N_1501,N_1799);
nor U2681 (N_2681,N_1832,N_1094);
or U2682 (N_2682,N_1733,N_1709);
and U2683 (N_2683,N_1558,N_1405);
or U2684 (N_2684,N_1372,N_1477);
nand U2685 (N_2685,N_1046,N_1225);
nor U2686 (N_2686,N_1465,N_1613);
nor U2687 (N_2687,N_1784,N_1476);
or U2688 (N_2688,N_1546,N_1552);
and U2689 (N_2689,N_1869,N_1592);
nand U2690 (N_2690,N_1404,N_1959);
nor U2691 (N_2691,N_1260,N_1126);
nand U2692 (N_2692,N_1690,N_1512);
nor U2693 (N_2693,N_1452,N_1590);
and U2694 (N_2694,N_1270,N_1844);
or U2695 (N_2695,N_1374,N_1466);
nand U2696 (N_2696,N_1001,N_1228);
nor U2697 (N_2697,N_1609,N_1701);
or U2698 (N_2698,N_1487,N_1511);
or U2699 (N_2699,N_1132,N_1907);
nor U2700 (N_2700,N_1406,N_1444);
nand U2701 (N_2701,N_1362,N_1107);
and U2702 (N_2702,N_1476,N_1817);
nor U2703 (N_2703,N_1315,N_1022);
nand U2704 (N_2704,N_1460,N_1046);
nor U2705 (N_2705,N_1607,N_1978);
and U2706 (N_2706,N_1732,N_1124);
nor U2707 (N_2707,N_1853,N_1264);
and U2708 (N_2708,N_1303,N_1525);
and U2709 (N_2709,N_1938,N_1319);
and U2710 (N_2710,N_1910,N_1209);
nand U2711 (N_2711,N_1835,N_1913);
nor U2712 (N_2712,N_1754,N_1978);
nand U2713 (N_2713,N_1885,N_1928);
or U2714 (N_2714,N_1615,N_1166);
and U2715 (N_2715,N_1656,N_1139);
and U2716 (N_2716,N_1555,N_1194);
nand U2717 (N_2717,N_1516,N_1782);
nand U2718 (N_2718,N_1076,N_1800);
nor U2719 (N_2719,N_1557,N_1907);
or U2720 (N_2720,N_1391,N_1599);
or U2721 (N_2721,N_1771,N_1720);
nor U2722 (N_2722,N_1230,N_1630);
or U2723 (N_2723,N_1768,N_1528);
nor U2724 (N_2724,N_1908,N_1772);
nand U2725 (N_2725,N_1902,N_1529);
or U2726 (N_2726,N_1494,N_1539);
nand U2727 (N_2727,N_1591,N_1574);
nor U2728 (N_2728,N_1568,N_1275);
nor U2729 (N_2729,N_1664,N_1125);
nand U2730 (N_2730,N_1735,N_1956);
nand U2731 (N_2731,N_1838,N_1154);
nand U2732 (N_2732,N_1953,N_1140);
and U2733 (N_2733,N_1748,N_1069);
or U2734 (N_2734,N_1322,N_1663);
nor U2735 (N_2735,N_1344,N_1192);
nor U2736 (N_2736,N_1366,N_1026);
nand U2737 (N_2737,N_1562,N_1012);
or U2738 (N_2738,N_1706,N_1698);
nor U2739 (N_2739,N_1508,N_1503);
or U2740 (N_2740,N_1383,N_1198);
and U2741 (N_2741,N_1317,N_1406);
or U2742 (N_2742,N_1624,N_1271);
or U2743 (N_2743,N_1328,N_1491);
nand U2744 (N_2744,N_1795,N_1229);
and U2745 (N_2745,N_1087,N_1453);
nand U2746 (N_2746,N_1421,N_1667);
or U2747 (N_2747,N_1719,N_1958);
or U2748 (N_2748,N_1209,N_1435);
nand U2749 (N_2749,N_1233,N_1766);
nand U2750 (N_2750,N_1109,N_1108);
nor U2751 (N_2751,N_1398,N_1156);
nand U2752 (N_2752,N_1846,N_1825);
nor U2753 (N_2753,N_1619,N_1148);
xnor U2754 (N_2754,N_1517,N_1476);
and U2755 (N_2755,N_1808,N_1920);
or U2756 (N_2756,N_1409,N_1919);
nor U2757 (N_2757,N_1427,N_1204);
or U2758 (N_2758,N_1257,N_1022);
nand U2759 (N_2759,N_1049,N_1997);
or U2760 (N_2760,N_1546,N_1243);
and U2761 (N_2761,N_1926,N_1088);
or U2762 (N_2762,N_1460,N_1230);
nand U2763 (N_2763,N_1928,N_1462);
and U2764 (N_2764,N_1874,N_1205);
nand U2765 (N_2765,N_1097,N_1063);
and U2766 (N_2766,N_1160,N_1876);
and U2767 (N_2767,N_1060,N_1016);
or U2768 (N_2768,N_1797,N_1981);
nor U2769 (N_2769,N_1588,N_1978);
nand U2770 (N_2770,N_1697,N_1037);
or U2771 (N_2771,N_1084,N_1251);
and U2772 (N_2772,N_1710,N_1547);
nor U2773 (N_2773,N_1725,N_1822);
nor U2774 (N_2774,N_1034,N_1504);
nor U2775 (N_2775,N_1995,N_1798);
nand U2776 (N_2776,N_1511,N_1042);
nor U2777 (N_2777,N_1846,N_1142);
nand U2778 (N_2778,N_1191,N_1799);
nand U2779 (N_2779,N_1254,N_1383);
nor U2780 (N_2780,N_1264,N_1832);
nand U2781 (N_2781,N_1131,N_1445);
and U2782 (N_2782,N_1609,N_1126);
and U2783 (N_2783,N_1857,N_1099);
nor U2784 (N_2784,N_1162,N_1755);
or U2785 (N_2785,N_1276,N_1982);
nor U2786 (N_2786,N_1411,N_1619);
nand U2787 (N_2787,N_1502,N_1085);
and U2788 (N_2788,N_1307,N_1719);
or U2789 (N_2789,N_1705,N_1202);
nor U2790 (N_2790,N_1974,N_1355);
or U2791 (N_2791,N_1390,N_1748);
or U2792 (N_2792,N_1829,N_1649);
xnor U2793 (N_2793,N_1685,N_1028);
nor U2794 (N_2794,N_1178,N_1531);
nand U2795 (N_2795,N_1090,N_1908);
nor U2796 (N_2796,N_1540,N_1094);
nor U2797 (N_2797,N_1580,N_1653);
and U2798 (N_2798,N_1995,N_1625);
and U2799 (N_2799,N_1370,N_1158);
or U2800 (N_2800,N_1788,N_1796);
nor U2801 (N_2801,N_1514,N_1127);
nand U2802 (N_2802,N_1302,N_1671);
and U2803 (N_2803,N_1851,N_1572);
or U2804 (N_2804,N_1730,N_1138);
and U2805 (N_2805,N_1762,N_1990);
or U2806 (N_2806,N_1753,N_1260);
nor U2807 (N_2807,N_1755,N_1796);
and U2808 (N_2808,N_1070,N_1542);
nor U2809 (N_2809,N_1313,N_1954);
or U2810 (N_2810,N_1486,N_1741);
nor U2811 (N_2811,N_1744,N_1135);
and U2812 (N_2812,N_1055,N_1407);
or U2813 (N_2813,N_1183,N_1621);
nand U2814 (N_2814,N_1751,N_1054);
and U2815 (N_2815,N_1325,N_1661);
nor U2816 (N_2816,N_1507,N_1564);
nor U2817 (N_2817,N_1375,N_1379);
nor U2818 (N_2818,N_1718,N_1321);
nor U2819 (N_2819,N_1838,N_1321);
nand U2820 (N_2820,N_1758,N_1250);
or U2821 (N_2821,N_1030,N_1298);
nand U2822 (N_2822,N_1757,N_1466);
or U2823 (N_2823,N_1128,N_1018);
xnor U2824 (N_2824,N_1023,N_1595);
nand U2825 (N_2825,N_1559,N_1453);
or U2826 (N_2826,N_1180,N_1070);
or U2827 (N_2827,N_1040,N_1099);
and U2828 (N_2828,N_1239,N_1553);
or U2829 (N_2829,N_1797,N_1628);
xor U2830 (N_2830,N_1544,N_1884);
or U2831 (N_2831,N_1772,N_1623);
nor U2832 (N_2832,N_1608,N_1682);
nand U2833 (N_2833,N_1606,N_1309);
nand U2834 (N_2834,N_1515,N_1853);
or U2835 (N_2835,N_1186,N_1443);
or U2836 (N_2836,N_1592,N_1339);
nand U2837 (N_2837,N_1532,N_1012);
or U2838 (N_2838,N_1785,N_1227);
nand U2839 (N_2839,N_1003,N_1674);
or U2840 (N_2840,N_1382,N_1257);
and U2841 (N_2841,N_1342,N_1966);
and U2842 (N_2842,N_1837,N_1960);
nand U2843 (N_2843,N_1389,N_1992);
nand U2844 (N_2844,N_1190,N_1881);
or U2845 (N_2845,N_1180,N_1528);
or U2846 (N_2846,N_1124,N_1435);
nand U2847 (N_2847,N_1716,N_1329);
nand U2848 (N_2848,N_1749,N_1217);
nand U2849 (N_2849,N_1691,N_1617);
and U2850 (N_2850,N_1654,N_1640);
and U2851 (N_2851,N_1831,N_1165);
or U2852 (N_2852,N_1473,N_1637);
nor U2853 (N_2853,N_1952,N_1371);
and U2854 (N_2854,N_1164,N_1905);
nand U2855 (N_2855,N_1035,N_1362);
or U2856 (N_2856,N_1764,N_1264);
xnor U2857 (N_2857,N_1927,N_1680);
nand U2858 (N_2858,N_1568,N_1513);
nor U2859 (N_2859,N_1302,N_1091);
nand U2860 (N_2860,N_1623,N_1938);
nand U2861 (N_2861,N_1871,N_1094);
and U2862 (N_2862,N_1633,N_1606);
nor U2863 (N_2863,N_1938,N_1738);
nor U2864 (N_2864,N_1311,N_1872);
nand U2865 (N_2865,N_1972,N_1100);
nor U2866 (N_2866,N_1820,N_1003);
or U2867 (N_2867,N_1383,N_1672);
nand U2868 (N_2868,N_1365,N_1886);
or U2869 (N_2869,N_1211,N_1117);
and U2870 (N_2870,N_1873,N_1773);
nor U2871 (N_2871,N_1672,N_1845);
nand U2872 (N_2872,N_1574,N_1344);
and U2873 (N_2873,N_1559,N_1635);
and U2874 (N_2874,N_1511,N_1092);
nand U2875 (N_2875,N_1535,N_1508);
nand U2876 (N_2876,N_1422,N_1090);
and U2877 (N_2877,N_1851,N_1351);
nor U2878 (N_2878,N_1723,N_1943);
nand U2879 (N_2879,N_1710,N_1050);
nor U2880 (N_2880,N_1691,N_1084);
and U2881 (N_2881,N_1145,N_1294);
or U2882 (N_2882,N_1800,N_1900);
xor U2883 (N_2883,N_1109,N_1474);
nor U2884 (N_2884,N_1506,N_1638);
nand U2885 (N_2885,N_1798,N_1578);
nor U2886 (N_2886,N_1121,N_1552);
nor U2887 (N_2887,N_1679,N_1812);
nor U2888 (N_2888,N_1497,N_1563);
nand U2889 (N_2889,N_1010,N_1825);
nand U2890 (N_2890,N_1556,N_1435);
nand U2891 (N_2891,N_1974,N_1094);
and U2892 (N_2892,N_1979,N_1722);
and U2893 (N_2893,N_1781,N_1734);
or U2894 (N_2894,N_1751,N_1615);
and U2895 (N_2895,N_1806,N_1713);
or U2896 (N_2896,N_1898,N_1668);
nand U2897 (N_2897,N_1508,N_1541);
or U2898 (N_2898,N_1889,N_1761);
nand U2899 (N_2899,N_1617,N_1643);
and U2900 (N_2900,N_1927,N_1395);
and U2901 (N_2901,N_1565,N_1529);
and U2902 (N_2902,N_1280,N_1342);
or U2903 (N_2903,N_1164,N_1126);
and U2904 (N_2904,N_1922,N_1025);
or U2905 (N_2905,N_1421,N_1167);
nor U2906 (N_2906,N_1565,N_1259);
or U2907 (N_2907,N_1881,N_1581);
and U2908 (N_2908,N_1068,N_1270);
nand U2909 (N_2909,N_1799,N_1139);
nand U2910 (N_2910,N_1468,N_1758);
or U2911 (N_2911,N_1194,N_1922);
or U2912 (N_2912,N_1515,N_1996);
nor U2913 (N_2913,N_1064,N_1654);
nand U2914 (N_2914,N_1883,N_1768);
and U2915 (N_2915,N_1722,N_1281);
or U2916 (N_2916,N_1214,N_1481);
or U2917 (N_2917,N_1256,N_1109);
and U2918 (N_2918,N_1668,N_1359);
and U2919 (N_2919,N_1989,N_1217);
nand U2920 (N_2920,N_1254,N_1095);
xor U2921 (N_2921,N_1130,N_1236);
and U2922 (N_2922,N_1372,N_1434);
nand U2923 (N_2923,N_1462,N_1985);
or U2924 (N_2924,N_1722,N_1917);
and U2925 (N_2925,N_1166,N_1753);
or U2926 (N_2926,N_1098,N_1217);
and U2927 (N_2927,N_1944,N_1598);
or U2928 (N_2928,N_1060,N_1556);
nand U2929 (N_2929,N_1404,N_1193);
nor U2930 (N_2930,N_1339,N_1240);
nor U2931 (N_2931,N_1562,N_1255);
nor U2932 (N_2932,N_1729,N_1981);
and U2933 (N_2933,N_1621,N_1780);
xor U2934 (N_2934,N_1891,N_1000);
and U2935 (N_2935,N_1050,N_1708);
or U2936 (N_2936,N_1847,N_1830);
and U2937 (N_2937,N_1212,N_1637);
nor U2938 (N_2938,N_1651,N_1908);
or U2939 (N_2939,N_1201,N_1029);
and U2940 (N_2940,N_1096,N_1663);
nor U2941 (N_2941,N_1341,N_1330);
nor U2942 (N_2942,N_1639,N_1088);
and U2943 (N_2943,N_1727,N_1051);
or U2944 (N_2944,N_1284,N_1515);
nand U2945 (N_2945,N_1982,N_1473);
or U2946 (N_2946,N_1801,N_1441);
nor U2947 (N_2947,N_1619,N_1217);
nand U2948 (N_2948,N_1045,N_1026);
nor U2949 (N_2949,N_1706,N_1058);
nor U2950 (N_2950,N_1796,N_1256);
nor U2951 (N_2951,N_1840,N_1581);
nor U2952 (N_2952,N_1875,N_1838);
and U2953 (N_2953,N_1267,N_1542);
and U2954 (N_2954,N_1278,N_1690);
nor U2955 (N_2955,N_1251,N_1756);
or U2956 (N_2956,N_1476,N_1401);
nor U2957 (N_2957,N_1943,N_1006);
or U2958 (N_2958,N_1541,N_1103);
xnor U2959 (N_2959,N_1111,N_1782);
or U2960 (N_2960,N_1841,N_1505);
nor U2961 (N_2961,N_1897,N_1578);
or U2962 (N_2962,N_1463,N_1043);
or U2963 (N_2963,N_1249,N_1315);
or U2964 (N_2964,N_1572,N_1198);
or U2965 (N_2965,N_1851,N_1004);
or U2966 (N_2966,N_1381,N_1576);
nor U2967 (N_2967,N_1036,N_1624);
or U2968 (N_2968,N_1966,N_1088);
nand U2969 (N_2969,N_1043,N_1798);
nand U2970 (N_2970,N_1818,N_1083);
or U2971 (N_2971,N_1913,N_1387);
nor U2972 (N_2972,N_1942,N_1532);
or U2973 (N_2973,N_1248,N_1574);
nand U2974 (N_2974,N_1839,N_1786);
and U2975 (N_2975,N_1234,N_1457);
nand U2976 (N_2976,N_1875,N_1391);
nor U2977 (N_2977,N_1246,N_1364);
or U2978 (N_2978,N_1461,N_1154);
or U2979 (N_2979,N_1431,N_1230);
and U2980 (N_2980,N_1849,N_1468);
and U2981 (N_2981,N_1592,N_1264);
and U2982 (N_2982,N_1871,N_1593);
nand U2983 (N_2983,N_1909,N_1589);
nand U2984 (N_2984,N_1605,N_1254);
nand U2985 (N_2985,N_1216,N_1204);
nand U2986 (N_2986,N_1065,N_1776);
nand U2987 (N_2987,N_1120,N_1213);
or U2988 (N_2988,N_1494,N_1381);
and U2989 (N_2989,N_1019,N_1699);
or U2990 (N_2990,N_1638,N_1362);
or U2991 (N_2991,N_1977,N_1832);
or U2992 (N_2992,N_1472,N_1860);
or U2993 (N_2993,N_1512,N_1663);
nor U2994 (N_2994,N_1875,N_1345);
and U2995 (N_2995,N_1867,N_1700);
and U2996 (N_2996,N_1179,N_1568);
xor U2997 (N_2997,N_1913,N_1139);
nand U2998 (N_2998,N_1067,N_1981);
nor U2999 (N_2999,N_1954,N_1697);
and U3000 (N_3000,N_2327,N_2734);
and U3001 (N_3001,N_2821,N_2118);
nand U3002 (N_3002,N_2162,N_2378);
and U3003 (N_3003,N_2782,N_2564);
nand U3004 (N_3004,N_2780,N_2167);
nand U3005 (N_3005,N_2326,N_2595);
or U3006 (N_3006,N_2049,N_2055);
or U3007 (N_3007,N_2028,N_2153);
nor U3008 (N_3008,N_2507,N_2877);
and U3009 (N_3009,N_2580,N_2294);
or U3010 (N_3010,N_2749,N_2302);
or U3011 (N_3011,N_2590,N_2976);
nand U3012 (N_3012,N_2943,N_2885);
and U3013 (N_3013,N_2374,N_2731);
or U3014 (N_3014,N_2910,N_2841);
nor U3015 (N_3015,N_2983,N_2081);
nor U3016 (N_3016,N_2756,N_2346);
and U3017 (N_3017,N_2314,N_2155);
or U3018 (N_3018,N_2690,N_2770);
nand U3019 (N_3019,N_2565,N_2515);
or U3020 (N_3020,N_2435,N_2000);
nand U3021 (N_3021,N_2644,N_2508);
nand U3022 (N_3022,N_2802,N_2450);
or U3023 (N_3023,N_2546,N_2427);
and U3024 (N_3024,N_2170,N_2874);
or U3025 (N_3025,N_2204,N_2186);
nand U3026 (N_3026,N_2233,N_2177);
and U3027 (N_3027,N_2964,N_2205);
or U3028 (N_3028,N_2924,N_2859);
or U3029 (N_3029,N_2568,N_2274);
nand U3030 (N_3030,N_2742,N_2539);
nand U3031 (N_3031,N_2748,N_2295);
nand U3032 (N_3032,N_2329,N_2847);
nand U3033 (N_3033,N_2579,N_2182);
nor U3034 (N_3034,N_2717,N_2684);
nand U3035 (N_3035,N_2262,N_2797);
or U3036 (N_3036,N_2328,N_2649);
and U3037 (N_3037,N_2862,N_2525);
and U3038 (N_3038,N_2098,N_2111);
nand U3039 (N_3039,N_2234,N_2566);
nor U3040 (N_3040,N_2471,N_2834);
or U3041 (N_3041,N_2975,N_2725);
nand U3042 (N_3042,N_2596,N_2735);
and U3043 (N_3043,N_2809,N_2597);
or U3044 (N_3044,N_2371,N_2033);
or U3045 (N_3045,N_2855,N_2154);
or U3046 (N_3046,N_2345,N_2157);
or U3047 (N_3047,N_2899,N_2465);
nor U3048 (N_3048,N_2627,N_2038);
nand U3049 (N_3049,N_2978,N_2608);
and U3050 (N_3050,N_2617,N_2338);
and U3051 (N_3051,N_2752,N_2444);
and U3052 (N_3052,N_2680,N_2385);
nand U3053 (N_3053,N_2881,N_2810);
or U3054 (N_3054,N_2784,N_2613);
or U3055 (N_3055,N_2016,N_2099);
nor U3056 (N_3056,N_2309,N_2093);
nor U3057 (N_3057,N_2576,N_2535);
nor U3058 (N_3058,N_2626,N_2942);
nand U3059 (N_3059,N_2252,N_2358);
or U3060 (N_3060,N_2168,N_2831);
or U3061 (N_3061,N_2119,N_2330);
or U3062 (N_3062,N_2022,N_2116);
nand U3063 (N_3063,N_2366,N_2823);
nand U3064 (N_3064,N_2029,N_2282);
and U3065 (N_3065,N_2714,N_2072);
and U3066 (N_3066,N_2872,N_2127);
nor U3067 (N_3067,N_2980,N_2082);
nor U3068 (N_3068,N_2667,N_2011);
or U3069 (N_3069,N_2506,N_2880);
nor U3070 (N_3070,N_2422,N_2504);
nor U3071 (N_3071,N_2661,N_2280);
nor U3072 (N_3072,N_2020,N_2962);
nor U3073 (N_3073,N_2973,N_2256);
or U3074 (N_3074,N_2587,N_2307);
or U3075 (N_3075,N_2025,N_2376);
nand U3076 (N_3076,N_2017,N_2904);
nor U3077 (N_3077,N_2032,N_2887);
and U3078 (N_3078,N_2100,N_2778);
nor U3079 (N_3079,N_2863,N_2795);
nand U3080 (N_3080,N_2505,N_2946);
or U3081 (N_3081,N_2551,N_2816);
nand U3082 (N_3082,N_2045,N_2296);
or U3083 (N_3083,N_2929,N_2369);
and U3084 (N_3084,N_2889,N_2960);
or U3085 (N_3085,N_2927,N_2707);
nor U3086 (N_3086,N_2455,N_2287);
nor U3087 (N_3087,N_2041,N_2244);
nand U3088 (N_3088,N_2226,N_2390);
nor U3089 (N_3089,N_2940,N_2763);
or U3090 (N_3090,N_2569,N_2266);
and U3091 (N_3091,N_2901,N_2658);
nand U3092 (N_3092,N_2854,N_2335);
nor U3093 (N_3093,N_2185,N_2736);
and U3094 (N_3094,N_2811,N_2830);
nand U3095 (N_3095,N_2715,N_2024);
or U3096 (N_3096,N_2729,N_2285);
nand U3097 (N_3097,N_2557,N_2298);
or U3098 (N_3098,N_2837,N_2228);
nor U3099 (N_3099,N_2351,N_2728);
nand U3100 (N_3100,N_2651,N_2112);
or U3101 (N_3101,N_2304,N_2395);
nor U3102 (N_3102,N_2951,N_2800);
and U3103 (N_3103,N_2408,N_2674);
and U3104 (N_3104,N_2637,N_2516);
and U3105 (N_3105,N_2340,N_2462);
nor U3106 (N_3106,N_2883,N_2056);
nand U3107 (N_3107,N_2563,N_2473);
nand U3108 (N_3108,N_2105,N_2132);
nor U3109 (N_3109,N_2074,N_2379);
and U3110 (N_3110,N_2218,N_2848);
nand U3111 (N_3111,N_2373,N_2187);
nor U3112 (N_3112,N_2997,N_2085);
or U3113 (N_3113,N_2466,N_2197);
nor U3114 (N_3114,N_2993,N_2347);
nor U3115 (N_3115,N_2625,N_2518);
nand U3116 (N_3116,N_2490,N_2584);
or U3117 (N_3117,N_2048,N_2896);
or U3118 (N_3118,N_2760,N_2487);
nor U3119 (N_3119,N_2148,N_2759);
and U3120 (N_3120,N_2601,N_2433);
nand U3121 (N_3121,N_2727,N_2747);
and U3122 (N_3122,N_2772,N_2381);
or U3123 (N_3123,N_2192,N_2886);
nand U3124 (N_3124,N_2701,N_2143);
and U3125 (N_3125,N_2069,N_2977);
or U3126 (N_3126,N_2773,N_2312);
and U3127 (N_3127,N_2722,N_2189);
or U3128 (N_3128,N_2918,N_2336);
nor U3129 (N_3129,N_2503,N_2656);
or U3130 (N_3130,N_2428,N_2913);
or U3131 (N_3131,N_2719,N_2136);
and U3132 (N_3132,N_2210,N_2398);
nor U3133 (N_3133,N_2589,N_2195);
nand U3134 (N_3134,N_2320,N_2783);
nand U3135 (N_3135,N_2938,N_2190);
and U3136 (N_3136,N_2125,N_2781);
or U3137 (N_3137,N_2540,N_2603);
and U3138 (N_3138,N_2982,N_2765);
and U3139 (N_3139,N_2861,N_2066);
nand U3140 (N_3140,N_2869,N_2893);
nand U3141 (N_3141,N_2392,N_2483);
or U3142 (N_3142,N_2552,N_2219);
or U3143 (N_3143,N_2776,N_2994);
or U3144 (N_3144,N_2633,N_2026);
or U3145 (N_3145,N_2092,N_2009);
and U3146 (N_3146,N_2064,N_2888);
and U3147 (N_3147,N_2316,N_2367);
and U3148 (N_3148,N_2194,N_2002);
and U3149 (N_3149,N_2801,N_2458);
nor U3150 (N_3150,N_2259,N_2394);
nor U3151 (N_3151,N_2995,N_2905);
and U3152 (N_3152,N_2891,N_2249);
nand U3153 (N_3153,N_2057,N_2915);
nor U3154 (N_3154,N_2835,N_2604);
nor U3155 (N_3155,N_2543,N_2434);
nor U3156 (N_3156,N_2819,N_2400);
or U3157 (N_3157,N_2334,N_2971);
nand U3158 (N_3158,N_2686,N_2225);
and U3159 (N_3159,N_2275,N_2716);
nor U3160 (N_3160,N_2332,N_2247);
and U3161 (N_3161,N_2992,N_2598);
and U3162 (N_3162,N_2386,N_2142);
or U3163 (N_3163,N_2426,N_2501);
or U3164 (N_3164,N_2849,N_2704);
nor U3165 (N_3165,N_2549,N_2542);
and U3166 (N_3166,N_2538,N_2526);
nor U3167 (N_3167,N_2903,N_2387);
nand U3168 (N_3168,N_2532,N_2939);
or U3169 (N_3169,N_2771,N_2986);
nand U3170 (N_3170,N_2529,N_2536);
nor U3171 (N_3171,N_2873,N_2870);
nand U3172 (N_3172,N_2289,N_2530);
or U3173 (N_3173,N_2303,N_2948);
nand U3174 (N_3174,N_2969,N_2574);
or U3175 (N_3175,N_2078,N_2953);
and U3176 (N_3176,N_2814,N_2325);
and U3177 (N_3177,N_2678,N_2628);
nor U3178 (N_3178,N_2246,N_2966);
and U3179 (N_3179,N_2003,N_2619);
and U3180 (N_3180,N_2944,N_2703);
nor U3181 (N_3181,N_2528,N_2682);
nor U3182 (N_3182,N_2695,N_2653);
nand U3183 (N_3183,N_2933,N_2646);
or U3184 (N_3184,N_2215,N_2791);
or U3185 (N_3185,N_2413,N_2494);
or U3186 (N_3186,N_2562,N_2990);
or U3187 (N_3187,N_2726,N_2318);
nand U3188 (N_3188,N_2076,N_2527);
nor U3189 (N_3189,N_2464,N_2161);
and U3190 (N_3190,N_2622,N_2169);
nand U3191 (N_3191,N_2101,N_2133);
nor U3192 (N_3192,N_2276,N_2263);
and U3193 (N_3193,N_2900,N_2631);
or U3194 (N_3194,N_2040,N_2806);
nand U3195 (N_3195,N_2470,N_2916);
nand U3196 (N_3196,N_2524,N_2609);
or U3197 (N_3197,N_2865,N_2592);
nand U3198 (N_3198,N_2988,N_2283);
and U3199 (N_3199,N_2547,N_2710);
or U3200 (N_3200,N_2659,N_2123);
or U3201 (N_3201,N_2001,N_2599);
and U3202 (N_3202,N_2152,N_2071);
and U3203 (N_3203,N_2388,N_2702);
xnor U3204 (N_3204,N_2397,N_2838);
nor U3205 (N_3205,N_2050,N_2203);
nor U3206 (N_3206,N_2815,N_2958);
nor U3207 (N_3207,N_2908,N_2229);
and U3208 (N_3208,N_2461,N_2544);
nand U3209 (N_3209,N_2895,N_2805);
or U3210 (N_3210,N_2130,N_2474);
nor U3211 (N_3211,N_2672,N_2406);
and U3212 (N_3212,N_2096,N_2581);
and U3213 (N_3213,N_2110,N_2764);
nor U3214 (N_3214,N_2804,N_2825);
nor U3215 (N_3215,N_2931,N_2774);
or U3216 (N_3216,N_2083,N_2404);
nand U3217 (N_3217,N_2477,N_2956);
or U3218 (N_3218,N_2065,N_2789);
nor U3219 (N_3219,N_2932,N_2242);
nand U3220 (N_3220,N_2221,N_2060);
nor U3221 (N_3221,N_2443,N_2419);
nand U3222 (N_3222,N_2241,N_2984);
or U3223 (N_3223,N_2621,N_2150);
nand U3224 (N_3224,N_2300,N_2585);
nand U3225 (N_3225,N_2531,N_2866);
or U3226 (N_3226,N_2359,N_2632);
and U3227 (N_3227,N_2106,N_2200);
nand U3228 (N_3228,N_2808,N_2522);
or U3229 (N_3229,N_2495,N_2115);
or U3230 (N_3230,N_2253,N_2344);
nor U3231 (N_3231,N_2324,N_2753);
and U3232 (N_3232,N_2441,N_2689);
or U3233 (N_3233,N_2243,N_2793);
nor U3234 (N_3234,N_2094,N_2593);
nor U3235 (N_3235,N_2673,N_2824);
nand U3236 (N_3236,N_2864,N_2537);
nand U3237 (N_3237,N_2623,N_2922);
or U3238 (N_3238,N_2149,N_2794);
or U3239 (N_3239,N_2087,N_2607);
nor U3240 (N_3240,N_2396,N_2213);
nor U3241 (N_3241,N_2250,N_2383);
and U3242 (N_3242,N_2489,N_2757);
or U3243 (N_3243,N_2758,N_2676);
nor U3244 (N_3244,N_2654,N_2139);
or U3245 (N_3245,N_2928,N_2176);
or U3246 (N_3246,N_2493,N_2708);
and U3247 (N_3247,N_2255,N_2611);
nand U3248 (N_3248,N_2140,N_2500);
and U3249 (N_3249,N_2846,N_2217);
xnor U3250 (N_3250,N_2812,N_2239);
and U3251 (N_3251,N_2237,N_2310);
nor U3252 (N_3252,N_2446,N_2286);
or U3253 (N_3253,N_2425,N_2588);
nand U3254 (N_3254,N_2231,N_2655);
nor U3255 (N_3255,N_2251,N_2860);
and U3256 (N_3256,N_2876,N_2311);
nand U3257 (N_3257,N_2448,N_2438);
nor U3258 (N_3258,N_2832,N_2878);
or U3259 (N_3259,N_2699,N_2292);
nor U3260 (N_3260,N_2550,N_2620);
nand U3261 (N_3261,N_2451,N_2754);
nand U3262 (N_3262,N_2365,N_2947);
and U3263 (N_3263,N_2496,N_2792);
nor U3264 (N_3264,N_2479,N_2269);
and U3265 (N_3265,N_2375,N_2468);
nor U3266 (N_3266,N_2052,N_2059);
and U3267 (N_3267,N_2453,N_2919);
and U3268 (N_3268,N_2897,N_2750);
nor U3269 (N_3269,N_2912,N_2817);
nor U3270 (N_3270,N_2670,N_2514);
nand U3271 (N_3271,N_2333,N_2432);
or U3272 (N_3272,N_2521,N_2989);
nor U3273 (N_3273,N_2222,N_2264);
nand U3274 (N_3274,N_2063,N_2355);
and U3275 (N_3275,N_2183,N_2921);
or U3276 (N_3276,N_2488,N_2600);
nand U3277 (N_3277,N_2440,N_2996);
nand U3278 (N_3278,N_2457,N_2520);
or U3279 (N_3279,N_2679,N_2353);
nor U3280 (N_3280,N_2271,N_2401);
or U3281 (N_3281,N_2840,N_2415);
and U3282 (N_3282,N_2934,N_2721);
and U3283 (N_3283,N_2305,N_2454);
or U3284 (N_3284,N_2519,N_2196);
or U3285 (N_3285,N_2165,N_2700);
or U3286 (N_3286,N_2512,N_2023);
nand U3287 (N_3287,N_2662,N_2013);
or U3288 (N_3288,N_2349,N_2743);
or U3289 (N_3289,N_2498,N_2151);
or U3290 (N_3290,N_2724,N_2128);
nor U3291 (N_3291,N_2021,N_2739);
or U3292 (N_3292,N_2265,N_2720);
nand U3293 (N_3293,N_2178,N_2945);
nand U3294 (N_3294,N_2614,N_2987);
or U3295 (N_3295,N_2560,N_2999);
nand U3296 (N_3296,N_2469,N_2472);
and U3297 (N_3297,N_2833,N_2985);
nand U3298 (N_3298,N_2798,N_2718);
nand U3299 (N_3299,N_2012,N_2787);
or U3300 (N_3300,N_2572,N_2019);
or U3301 (N_3301,N_2852,N_2578);
and U3302 (N_3302,N_2027,N_2911);
nand U3303 (N_3303,N_2769,N_2380);
nor U3304 (N_3304,N_2641,N_2267);
nor U3305 (N_3305,N_2967,N_2278);
nand U3306 (N_3306,N_2207,N_2972);
and U3307 (N_3307,N_2981,N_2051);
nor U3308 (N_3308,N_2343,N_2270);
or U3309 (N_3309,N_2301,N_2416);
xnor U3310 (N_3310,N_2652,N_2618);
nor U3311 (N_3311,N_2370,N_2047);
nor U3312 (N_3312,N_2058,N_2350);
nor U3313 (N_3313,N_2126,N_2117);
nand U3314 (N_3314,N_2491,N_2820);
or U3315 (N_3315,N_2171,N_2160);
nor U3316 (N_3316,N_2348,N_2067);
or U3317 (N_3317,N_2744,N_2436);
nand U3318 (N_3318,N_2577,N_2635);
and U3319 (N_3319,N_2372,N_2418);
nor U3320 (N_3320,N_2610,N_2460);
nor U3321 (N_3321,N_2368,N_2675);
or U3322 (N_3322,N_2054,N_2297);
or U3323 (N_3323,N_2232,N_2240);
and U3324 (N_3324,N_2147,N_2467);
and U3325 (N_3325,N_2914,N_2868);
or U3326 (N_3326,N_2583,N_2688);
or U3327 (N_3327,N_2409,N_2144);
and U3328 (N_3328,N_2979,N_2486);
and U3329 (N_3329,N_2008,N_2894);
nor U3330 (N_3330,N_2042,N_2254);
or U3331 (N_3331,N_2363,N_2737);
and U3332 (N_3332,N_2779,N_2902);
nor U3333 (N_3333,N_2073,N_2712);
or U3334 (N_3334,N_2882,N_2687);
nand U3335 (N_3335,N_2634,N_2352);
nor U3336 (N_3336,N_2268,N_2698);
or U3337 (N_3337,N_2236,N_2829);
nand U3338 (N_3338,N_2696,N_2079);
and U3339 (N_3339,N_2998,N_2665);
nor U3340 (N_3340,N_2691,N_2697);
nor U3341 (N_3341,N_2035,N_2786);
nor U3342 (N_3342,N_2173,N_2129);
nor U3343 (N_3343,N_2208,N_2497);
nand U3344 (N_3344,N_2006,N_2850);
or U3345 (N_3345,N_2517,N_2559);
nand U3346 (N_3346,N_2492,N_2181);
nand U3347 (N_3347,N_2965,N_2478);
nor U3348 (N_3348,N_2039,N_2669);
nor U3349 (N_3349,N_2745,N_2260);
and U3350 (N_3350,N_2954,N_2807);
nand U3351 (N_3351,N_2211,N_2313);
and U3352 (N_3352,N_2857,N_2230);
nand U3353 (N_3353,N_2723,N_2636);
nand U3354 (N_3354,N_2818,N_2163);
nand U3355 (N_3355,N_2567,N_2423);
nand U3356 (N_3356,N_2108,N_2879);
and U3357 (N_3357,N_2602,N_2091);
nor U3358 (N_3358,N_2261,N_2452);
nor U3359 (N_3359,N_2164,N_2293);
nand U3360 (N_3360,N_2037,N_2935);
or U3361 (N_3361,N_2509,N_2141);
nand U3362 (N_3362,N_2137,N_2920);
nor U3363 (N_3363,N_2768,N_2867);
nor U3364 (N_3364,N_2323,N_2671);
and U3365 (N_3365,N_2766,N_2582);
nand U3366 (N_3366,N_2523,N_2339);
and U3367 (N_3367,N_2871,N_2445);
nand U3368 (N_3368,N_2061,N_2476);
and U3369 (N_3369,N_2612,N_2828);
nor U3370 (N_3370,N_2796,N_2694);
or U3371 (N_3371,N_2212,N_2273);
nand U3372 (N_3372,N_2959,N_2842);
and U3373 (N_3373,N_2510,N_2319);
nand U3374 (N_3374,N_2555,N_2660);
nor U3375 (N_3375,N_2909,N_2402);
nand U3376 (N_3376,N_2382,N_2412);
nor U3377 (N_3377,N_2179,N_2075);
and U3378 (N_3378,N_2845,N_2088);
nor U3379 (N_3379,N_2227,N_2638);
and U3380 (N_3380,N_2875,N_2031);
xnor U3381 (N_3381,N_2175,N_2356);
and U3382 (N_3382,N_2102,N_2648);
nand U3383 (N_3383,N_2963,N_2214);
nor U3384 (N_3384,N_2591,N_2643);
nor U3385 (N_3385,N_2534,N_2777);
and U3386 (N_3386,N_2044,N_2561);
nor U3387 (N_3387,N_2898,N_2272);
or U3388 (N_3388,N_2799,N_2545);
nand U3389 (N_3389,N_2968,N_2015);
or U3390 (N_3390,N_2640,N_2159);
or U3391 (N_3391,N_2188,N_2384);
nand U3392 (N_3392,N_2755,N_2354);
nand U3393 (N_3393,N_2481,N_2198);
nor U3394 (N_3394,N_2556,N_2166);
nand U3395 (N_3395,N_2104,N_2606);
or U3396 (N_3396,N_2456,N_2482);
and U3397 (N_3397,N_2279,N_2925);
and U3398 (N_3398,N_2693,N_2107);
nor U3399 (N_3399,N_2331,N_2711);
nor U3400 (N_3400,N_2223,N_2357);
nand U3401 (N_3401,N_2172,N_2124);
or U3402 (N_3402,N_2420,N_2018);
or U3403 (N_3403,N_2629,N_2575);
or U3404 (N_3404,N_2930,N_2650);
nor U3405 (N_3405,N_2341,N_2647);
nor U3406 (N_3406,N_2449,N_2321);
and U3407 (N_3407,N_2403,N_2220);
or U3408 (N_3408,N_2389,N_2235);
and U3409 (N_3409,N_2417,N_2014);
nand U3410 (N_3410,N_2068,N_2813);
or U3411 (N_3411,N_2616,N_2974);
nand U3412 (N_3412,N_2853,N_2666);
nor U3413 (N_3413,N_2258,N_2917);
nor U3414 (N_3414,N_2277,N_2030);
nor U3415 (N_3415,N_2706,N_2475);
or U3416 (N_3416,N_2856,N_2843);
nor U3417 (N_3417,N_2089,N_2991);
or U3418 (N_3418,N_2553,N_2424);
or U3419 (N_3419,N_2554,N_2122);
and U3420 (N_3420,N_2109,N_2664);
nor U3421 (N_3421,N_2114,N_2890);
or U3422 (N_3422,N_2746,N_2836);
or U3423 (N_3423,N_2955,N_2624);
nand U3424 (N_3424,N_2892,N_2513);
nand U3425 (N_3425,N_2005,N_2248);
or U3426 (N_3426,N_2570,N_2683);
nand U3427 (N_3427,N_2290,N_2393);
and U3428 (N_3428,N_2216,N_2411);
nor U3429 (N_3429,N_2224,N_2391);
nand U3430 (N_3430,N_2377,N_2437);
and U3431 (N_3431,N_2043,N_2605);
nand U3432 (N_3432,N_2281,N_2086);
or U3433 (N_3433,N_2858,N_2131);
or U3434 (N_3434,N_2010,N_2080);
and U3435 (N_3435,N_2135,N_2439);
nor U3436 (N_3436,N_2209,N_2399);
and U3437 (N_3437,N_2738,N_2070);
nor U3438 (N_3438,N_2788,N_2548);
nor U3439 (N_3439,N_2360,N_2822);
nor U3440 (N_3440,N_2145,N_2034);
and U3441 (N_3441,N_2421,N_2767);
or U3442 (N_3442,N_2180,N_2826);
and U3443 (N_3443,N_2036,N_2558);
nand U3444 (N_3444,N_2484,N_2677);
or U3445 (N_3445,N_2571,N_2362);
and U3446 (N_3446,N_2120,N_2681);
nand U3447 (N_3447,N_2299,N_2923);
or U3448 (N_3448,N_2790,N_2541);
and U3449 (N_3449,N_2447,N_2193);
or U3450 (N_3450,N_2184,N_2095);
nor U3451 (N_3451,N_2630,N_2709);
nor U3452 (N_3452,N_2761,N_2502);
or U3453 (N_3453,N_2084,N_2046);
nor U3454 (N_3454,N_2199,N_2414);
and U3455 (N_3455,N_2844,N_2202);
and U3456 (N_3456,N_2685,N_2315);
and U3457 (N_3457,N_2121,N_2499);
and U3458 (N_3458,N_2586,N_2317);
or U3459 (N_3459,N_2257,N_2663);
nor U3460 (N_3460,N_2713,N_2463);
nand U3461 (N_3461,N_2740,N_2906);
nor U3462 (N_3462,N_2245,N_2615);
and U3463 (N_3463,N_2533,N_2642);
nor U3464 (N_3464,N_2364,N_2952);
nor U3465 (N_3465,N_2803,N_2639);
and U3466 (N_3466,N_2004,N_2113);
and U3467 (N_3467,N_2077,N_2949);
nor U3468 (N_3468,N_2322,N_2884);
nand U3469 (N_3469,N_2097,N_2645);
nand U3470 (N_3470,N_2284,N_2839);
or U3471 (N_3471,N_2134,N_2146);
and U3472 (N_3472,N_2657,N_2741);
and U3473 (N_3473,N_2692,N_2970);
and U3474 (N_3474,N_2007,N_2361);
nor U3475 (N_3475,N_2337,N_2429);
and U3476 (N_3476,N_2926,N_2405);
and U3477 (N_3477,N_2827,N_2431);
nand U3478 (N_3478,N_2410,N_2442);
nor U3479 (N_3479,N_2288,N_2936);
or U3480 (N_3480,N_2306,N_2957);
and U3481 (N_3481,N_2174,N_2775);
nand U3482 (N_3482,N_2785,N_2308);
nand U3483 (N_3483,N_2062,N_2594);
or U3484 (N_3484,N_2459,N_2156);
nand U3485 (N_3485,N_2201,N_2291);
or U3486 (N_3486,N_2751,N_2053);
or U3487 (N_3487,N_2941,N_2138);
and U3488 (N_3488,N_2950,N_2090);
nor U3489 (N_3489,N_2485,N_2730);
nor U3490 (N_3490,N_2342,N_2206);
nand U3491 (N_3491,N_2937,N_2511);
nand U3492 (N_3492,N_2103,N_2407);
and U3493 (N_3493,N_2851,N_2158);
or U3494 (N_3494,N_2705,N_2907);
nand U3495 (N_3495,N_2961,N_2238);
and U3496 (N_3496,N_2573,N_2732);
nand U3497 (N_3497,N_2430,N_2762);
and U3498 (N_3498,N_2668,N_2191);
nand U3499 (N_3499,N_2480,N_2733);
and U3500 (N_3500,N_2674,N_2703);
and U3501 (N_3501,N_2776,N_2779);
and U3502 (N_3502,N_2650,N_2690);
or U3503 (N_3503,N_2694,N_2512);
nand U3504 (N_3504,N_2745,N_2065);
nor U3505 (N_3505,N_2718,N_2347);
xnor U3506 (N_3506,N_2322,N_2440);
nor U3507 (N_3507,N_2358,N_2045);
or U3508 (N_3508,N_2336,N_2826);
and U3509 (N_3509,N_2847,N_2381);
or U3510 (N_3510,N_2725,N_2463);
or U3511 (N_3511,N_2192,N_2401);
nor U3512 (N_3512,N_2469,N_2428);
nand U3513 (N_3513,N_2219,N_2058);
or U3514 (N_3514,N_2995,N_2977);
nand U3515 (N_3515,N_2444,N_2373);
or U3516 (N_3516,N_2481,N_2183);
nor U3517 (N_3517,N_2602,N_2865);
nor U3518 (N_3518,N_2015,N_2900);
and U3519 (N_3519,N_2214,N_2424);
nor U3520 (N_3520,N_2223,N_2991);
nor U3521 (N_3521,N_2290,N_2228);
nand U3522 (N_3522,N_2125,N_2580);
or U3523 (N_3523,N_2418,N_2412);
nand U3524 (N_3524,N_2162,N_2641);
nor U3525 (N_3525,N_2092,N_2454);
nand U3526 (N_3526,N_2284,N_2184);
nand U3527 (N_3527,N_2359,N_2306);
nor U3528 (N_3528,N_2784,N_2196);
and U3529 (N_3529,N_2489,N_2816);
and U3530 (N_3530,N_2630,N_2225);
and U3531 (N_3531,N_2000,N_2609);
nor U3532 (N_3532,N_2409,N_2712);
nand U3533 (N_3533,N_2291,N_2849);
and U3534 (N_3534,N_2805,N_2856);
and U3535 (N_3535,N_2396,N_2428);
and U3536 (N_3536,N_2272,N_2662);
and U3537 (N_3537,N_2100,N_2852);
and U3538 (N_3538,N_2255,N_2406);
nand U3539 (N_3539,N_2736,N_2438);
and U3540 (N_3540,N_2907,N_2377);
nand U3541 (N_3541,N_2170,N_2442);
and U3542 (N_3542,N_2104,N_2050);
nor U3543 (N_3543,N_2418,N_2081);
nor U3544 (N_3544,N_2638,N_2937);
or U3545 (N_3545,N_2677,N_2067);
nand U3546 (N_3546,N_2668,N_2909);
nand U3547 (N_3547,N_2180,N_2110);
and U3548 (N_3548,N_2579,N_2769);
or U3549 (N_3549,N_2477,N_2585);
and U3550 (N_3550,N_2525,N_2898);
or U3551 (N_3551,N_2572,N_2031);
and U3552 (N_3552,N_2658,N_2847);
nor U3553 (N_3553,N_2842,N_2116);
nor U3554 (N_3554,N_2381,N_2160);
and U3555 (N_3555,N_2205,N_2369);
nand U3556 (N_3556,N_2218,N_2233);
and U3557 (N_3557,N_2424,N_2659);
or U3558 (N_3558,N_2483,N_2488);
or U3559 (N_3559,N_2395,N_2986);
nor U3560 (N_3560,N_2041,N_2069);
nand U3561 (N_3561,N_2717,N_2834);
nand U3562 (N_3562,N_2916,N_2650);
or U3563 (N_3563,N_2548,N_2764);
nand U3564 (N_3564,N_2738,N_2198);
nor U3565 (N_3565,N_2012,N_2297);
nand U3566 (N_3566,N_2085,N_2668);
and U3567 (N_3567,N_2285,N_2684);
or U3568 (N_3568,N_2690,N_2991);
nor U3569 (N_3569,N_2578,N_2380);
nand U3570 (N_3570,N_2520,N_2888);
and U3571 (N_3571,N_2751,N_2397);
nand U3572 (N_3572,N_2390,N_2783);
or U3573 (N_3573,N_2533,N_2749);
nor U3574 (N_3574,N_2181,N_2197);
nand U3575 (N_3575,N_2214,N_2929);
and U3576 (N_3576,N_2781,N_2217);
nor U3577 (N_3577,N_2881,N_2422);
nor U3578 (N_3578,N_2454,N_2063);
or U3579 (N_3579,N_2225,N_2803);
nor U3580 (N_3580,N_2440,N_2968);
or U3581 (N_3581,N_2027,N_2139);
nand U3582 (N_3582,N_2561,N_2041);
and U3583 (N_3583,N_2791,N_2440);
nand U3584 (N_3584,N_2630,N_2040);
nor U3585 (N_3585,N_2836,N_2362);
and U3586 (N_3586,N_2372,N_2391);
nor U3587 (N_3587,N_2330,N_2575);
nor U3588 (N_3588,N_2460,N_2660);
nand U3589 (N_3589,N_2054,N_2367);
or U3590 (N_3590,N_2513,N_2351);
or U3591 (N_3591,N_2674,N_2832);
nor U3592 (N_3592,N_2423,N_2997);
and U3593 (N_3593,N_2371,N_2055);
nand U3594 (N_3594,N_2964,N_2494);
and U3595 (N_3595,N_2195,N_2773);
nand U3596 (N_3596,N_2925,N_2137);
nand U3597 (N_3597,N_2626,N_2898);
or U3598 (N_3598,N_2556,N_2093);
or U3599 (N_3599,N_2679,N_2197);
nor U3600 (N_3600,N_2745,N_2737);
or U3601 (N_3601,N_2947,N_2883);
and U3602 (N_3602,N_2443,N_2023);
or U3603 (N_3603,N_2539,N_2314);
nand U3604 (N_3604,N_2644,N_2052);
and U3605 (N_3605,N_2746,N_2020);
or U3606 (N_3606,N_2245,N_2031);
nand U3607 (N_3607,N_2031,N_2634);
nor U3608 (N_3608,N_2979,N_2905);
nand U3609 (N_3609,N_2436,N_2009);
nor U3610 (N_3610,N_2773,N_2923);
and U3611 (N_3611,N_2346,N_2658);
or U3612 (N_3612,N_2197,N_2898);
nand U3613 (N_3613,N_2611,N_2391);
and U3614 (N_3614,N_2557,N_2881);
or U3615 (N_3615,N_2119,N_2486);
xor U3616 (N_3616,N_2099,N_2118);
and U3617 (N_3617,N_2963,N_2686);
nor U3618 (N_3618,N_2587,N_2704);
nand U3619 (N_3619,N_2971,N_2404);
or U3620 (N_3620,N_2851,N_2889);
or U3621 (N_3621,N_2993,N_2136);
and U3622 (N_3622,N_2892,N_2699);
nor U3623 (N_3623,N_2510,N_2110);
nor U3624 (N_3624,N_2841,N_2623);
or U3625 (N_3625,N_2088,N_2792);
nor U3626 (N_3626,N_2055,N_2646);
and U3627 (N_3627,N_2495,N_2054);
nand U3628 (N_3628,N_2510,N_2474);
nand U3629 (N_3629,N_2449,N_2383);
and U3630 (N_3630,N_2908,N_2555);
and U3631 (N_3631,N_2931,N_2282);
or U3632 (N_3632,N_2993,N_2511);
or U3633 (N_3633,N_2911,N_2549);
nand U3634 (N_3634,N_2264,N_2292);
nand U3635 (N_3635,N_2244,N_2610);
nand U3636 (N_3636,N_2126,N_2145);
or U3637 (N_3637,N_2501,N_2304);
and U3638 (N_3638,N_2467,N_2132);
and U3639 (N_3639,N_2146,N_2307);
nor U3640 (N_3640,N_2577,N_2909);
or U3641 (N_3641,N_2610,N_2730);
nor U3642 (N_3642,N_2866,N_2001);
nand U3643 (N_3643,N_2903,N_2639);
or U3644 (N_3644,N_2387,N_2595);
or U3645 (N_3645,N_2757,N_2198);
or U3646 (N_3646,N_2644,N_2095);
nor U3647 (N_3647,N_2354,N_2153);
nand U3648 (N_3648,N_2386,N_2481);
nand U3649 (N_3649,N_2630,N_2995);
nor U3650 (N_3650,N_2334,N_2757);
or U3651 (N_3651,N_2603,N_2435);
nand U3652 (N_3652,N_2800,N_2544);
nor U3653 (N_3653,N_2411,N_2599);
and U3654 (N_3654,N_2419,N_2045);
nor U3655 (N_3655,N_2367,N_2817);
nor U3656 (N_3656,N_2409,N_2173);
or U3657 (N_3657,N_2433,N_2379);
nor U3658 (N_3658,N_2149,N_2854);
or U3659 (N_3659,N_2629,N_2282);
and U3660 (N_3660,N_2592,N_2438);
and U3661 (N_3661,N_2935,N_2342);
and U3662 (N_3662,N_2325,N_2761);
nand U3663 (N_3663,N_2388,N_2481);
nand U3664 (N_3664,N_2158,N_2665);
or U3665 (N_3665,N_2851,N_2111);
nand U3666 (N_3666,N_2159,N_2817);
nand U3667 (N_3667,N_2182,N_2672);
and U3668 (N_3668,N_2000,N_2710);
or U3669 (N_3669,N_2399,N_2298);
nand U3670 (N_3670,N_2366,N_2265);
and U3671 (N_3671,N_2915,N_2558);
or U3672 (N_3672,N_2018,N_2766);
or U3673 (N_3673,N_2975,N_2571);
nand U3674 (N_3674,N_2287,N_2158);
nand U3675 (N_3675,N_2165,N_2923);
or U3676 (N_3676,N_2119,N_2846);
nand U3677 (N_3677,N_2093,N_2441);
or U3678 (N_3678,N_2656,N_2906);
or U3679 (N_3679,N_2993,N_2239);
and U3680 (N_3680,N_2129,N_2916);
nor U3681 (N_3681,N_2049,N_2982);
or U3682 (N_3682,N_2534,N_2370);
nand U3683 (N_3683,N_2936,N_2105);
or U3684 (N_3684,N_2780,N_2106);
xor U3685 (N_3685,N_2040,N_2122);
nor U3686 (N_3686,N_2997,N_2421);
or U3687 (N_3687,N_2534,N_2369);
nor U3688 (N_3688,N_2819,N_2062);
nor U3689 (N_3689,N_2105,N_2897);
nor U3690 (N_3690,N_2318,N_2633);
nor U3691 (N_3691,N_2174,N_2539);
nand U3692 (N_3692,N_2620,N_2989);
nand U3693 (N_3693,N_2313,N_2195);
and U3694 (N_3694,N_2686,N_2604);
nor U3695 (N_3695,N_2264,N_2221);
nand U3696 (N_3696,N_2320,N_2982);
nand U3697 (N_3697,N_2069,N_2954);
nand U3698 (N_3698,N_2905,N_2604);
nand U3699 (N_3699,N_2798,N_2490);
nand U3700 (N_3700,N_2451,N_2943);
nand U3701 (N_3701,N_2660,N_2960);
nand U3702 (N_3702,N_2623,N_2975);
and U3703 (N_3703,N_2864,N_2194);
or U3704 (N_3704,N_2252,N_2689);
and U3705 (N_3705,N_2454,N_2512);
and U3706 (N_3706,N_2186,N_2766);
nand U3707 (N_3707,N_2720,N_2589);
and U3708 (N_3708,N_2595,N_2565);
and U3709 (N_3709,N_2487,N_2345);
nand U3710 (N_3710,N_2820,N_2081);
nor U3711 (N_3711,N_2518,N_2611);
nor U3712 (N_3712,N_2745,N_2954);
or U3713 (N_3713,N_2607,N_2000);
and U3714 (N_3714,N_2073,N_2200);
nor U3715 (N_3715,N_2126,N_2653);
and U3716 (N_3716,N_2756,N_2356);
and U3717 (N_3717,N_2980,N_2607);
or U3718 (N_3718,N_2052,N_2712);
nor U3719 (N_3719,N_2017,N_2544);
nor U3720 (N_3720,N_2046,N_2251);
or U3721 (N_3721,N_2771,N_2901);
nand U3722 (N_3722,N_2978,N_2800);
and U3723 (N_3723,N_2515,N_2073);
nor U3724 (N_3724,N_2946,N_2864);
or U3725 (N_3725,N_2852,N_2354);
nand U3726 (N_3726,N_2961,N_2662);
nand U3727 (N_3727,N_2949,N_2169);
nand U3728 (N_3728,N_2638,N_2744);
nor U3729 (N_3729,N_2821,N_2645);
and U3730 (N_3730,N_2112,N_2435);
or U3731 (N_3731,N_2130,N_2178);
nor U3732 (N_3732,N_2598,N_2437);
nor U3733 (N_3733,N_2036,N_2443);
nand U3734 (N_3734,N_2164,N_2530);
nand U3735 (N_3735,N_2265,N_2355);
nor U3736 (N_3736,N_2879,N_2650);
or U3737 (N_3737,N_2351,N_2447);
and U3738 (N_3738,N_2649,N_2058);
nand U3739 (N_3739,N_2906,N_2183);
nor U3740 (N_3740,N_2657,N_2661);
nor U3741 (N_3741,N_2049,N_2815);
nand U3742 (N_3742,N_2788,N_2123);
xnor U3743 (N_3743,N_2434,N_2723);
nor U3744 (N_3744,N_2539,N_2793);
nand U3745 (N_3745,N_2271,N_2116);
and U3746 (N_3746,N_2412,N_2639);
and U3747 (N_3747,N_2630,N_2632);
and U3748 (N_3748,N_2518,N_2202);
and U3749 (N_3749,N_2753,N_2119);
nor U3750 (N_3750,N_2863,N_2221);
nand U3751 (N_3751,N_2554,N_2016);
nor U3752 (N_3752,N_2467,N_2624);
and U3753 (N_3753,N_2165,N_2427);
nor U3754 (N_3754,N_2979,N_2572);
nor U3755 (N_3755,N_2635,N_2591);
nor U3756 (N_3756,N_2438,N_2250);
nand U3757 (N_3757,N_2418,N_2114);
nand U3758 (N_3758,N_2147,N_2515);
nand U3759 (N_3759,N_2549,N_2767);
or U3760 (N_3760,N_2301,N_2149);
and U3761 (N_3761,N_2225,N_2298);
or U3762 (N_3762,N_2319,N_2083);
nand U3763 (N_3763,N_2433,N_2997);
nor U3764 (N_3764,N_2288,N_2364);
xor U3765 (N_3765,N_2555,N_2528);
nand U3766 (N_3766,N_2336,N_2349);
nand U3767 (N_3767,N_2695,N_2620);
and U3768 (N_3768,N_2489,N_2975);
nand U3769 (N_3769,N_2482,N_2859);
and U3770 (N_3770,N_2656,N_2179);
nor U3771 (N_3771,N_2092,N_2899);
or U3772 (N_3772,N_2503,N_2434);
nor U3773 (N_3773,N_2359,N_2870);
and U3774 (N_3774,N_2000,N_2605);
nand U3775 (N_3775,N_2886,N_2245);
or U3776 (N_3776,N_2115,N_2677);
nor U3777 (N_3777,N_2148,N_2885);
or U3778 (N_3778,N_2206,N_2082);
nand U3779 (N_3779,N_2889,N_2613);
nand U3780 (N_3780,N_2110,N_2588);
and U3781 (N_3781,N_2955,N_2634);
nor U3782 (N_3782,N_2145,N_2035);
nand U3783 (N_3783,N_2999,N_2029);
or U3784 (N_3784,N_2184,N_2978);
nand U3785 (N_3785,N_2425,N_2838);
or U3786 (N_3786,N_2607,N_2203);
nand U3787 (N_3787,N_2522,N_2658);
nand U3788 (N_3788,N_2108,N_2228);
nand U3789 (N_3789,N_2821,N_2479);
or U3790 (N_3790,N_2508,N_2665);
or U3791 (N_3791,N_2626,N_2292);
and U3792 (N_3792,N_2494,N_2070);
and U3793 (N_3793,N_2323,N_2893);
nor U3794 (N_3794,N_2271,N_2508);
and U3795 (N_3795,N_2770,N_2489);
nand U3796 (N_3796,N_2242,N_2320);
nand U3797 (N_3797,N_2349,N_2877);
nor U3798 (N_3798,N_2122,N_2692);
and U3799 (N_3799,N_2440,N_2166);
or U3800 (N_3800,N_2086,N_2625);
nand U3801 (N_3801,N_2632,N_2145);
and U3802 (N_3802,N_2942,N_2019);
nor U3803 (N_3803,N_2329,N_2374);
or U3804 (N_3804,N_2902,N_2150);
and U3805 (N_3805,N_2204,N_2349);
nand U3806 (N_3806,N_2228,N_2494);
nand U3807 (N_3807,N_2697,N_2821);
nor U3808 (N_3808,N_2141,N_2015);
nor U3809 (N_3809,N_2711,N_2080);
nor U3810 (N_3810,N_2123,N_2516);
nand U3811 (N_3811,N_2049,N_2750);
nor U3812 (N_3812,N_2301,N_2142);
nor U3813 (N_3813,N_2954,N_2519);
nand U3814 (N_3814,N_2222,N_2901);
or U3815 (N_3815,N_2690,N_2317);
and U3816 (N_3816,N_2278,N_2218);
nand U3817 (N_3817,N_2069,N_2134);
nand U3818 (N_3818,N_2639,N_2027);
nand U3819 (N_3819,N_2256,N_2981);
and U3820 (N_3820,N_2678,N_2199);
nor U3821 (N_3821,N_2693,N_2527);
or U3822 (N_3822,N_2372,N_2380);
nand U3823 (N_3823,N_2313,N_2570);
or U3824 (N_3824,N_2575,N_2225);
and U3825 (N_3825,N_2754,N_2904);
nor U3826 (N_3826,N_2034,N_2228);
nand U3827 (N_3827,N_2813,N_2511);
or U3828 (N_3828,N_2728,N_2112);
nor U3829 (N_3829,N_2671,N_2443);
or U3830 (N_3830,N_2566,N_2519);
or U3831 (N_3831,N_2275,N_2107);
nor U3832 (N_3832,N_2995,N_2649);
or U3833 (N_3833,N_2533,N_2643);
nor U3834 (N_3834,N_2219,N_2280);
or U3835 (N_3835,N_2458,N_2247);
or U3836 (N_3836,N_2736,N_2592);
or U3837 (N_3837,N_2327,N_2387);
nand U3838 (N_3838,N_2870,N_2924);
and U3839 (N_3839,N_2846,N_2853);
or U3840 (N_3840,N_2549,N_2788);
and U3841 (N_3841,N_2529,N_2715);
and U3842 (N_3842,N_2059,N_2619);
nor U3843 (N_3843,N_2558,N_2419);
nand U3844 (N_3844,N_2899,N_2020);
nand U3845 (N_3845,N_2977,N_2539);
nand U3846 (N_3846,N_2660,N_2549);
and U3847 (N_3847,N_2472,N_2052);
xnor U3848 (N_3848,N_2185,N_2468);
or U3849 (N_3849,N_2238,N_2300);
or U3850 (N_3850,N_2697,N_2013);
nor U3851 (N_3851,N_2034,N_2419);
nand U3852 (N_3852,N_2956,N_2084);
or U3853 (N_3853,N_2989,N_2766);
and U3854 (N_3854,N_2344,N_2189);
nand U3855 (N_3855,N_2832,N_2758);
xnor U3856 (N_3856,N_2481,N_2510);
nor U3857 (N_3857,N_2272,N_2388);
nor U3858 (N_3858,N_2111,N_2780);
or U3859 (N_3859,N_2075,N_2515);
and U3860 (N_3860,N_2632,N_2243);
nor U3861 (N_3861,N_2987,N_2274);
nor U3862 (N_3862,N_2149,N_2859);
nand U3863 (N_3863,N_2677,N_2112);
nand U3864 (N_3864,N_2344,N_2631);
nand U3865 (N_3865,N_2715,N_2386);
nor U3866 (N_3866,N_2864,N_2790);
or U3867 (N_3867,N_2816,N_2852);
and U3868 (N_3868,N_2796,N_2242);
or U3869 (N_3869,N_2814,N_2350);
nor U3870 (N_3870,N_2212,N_2415);
and U3871 (N_3871,N_2286,N_2332);
nand U3872 (N_3872,N_2502,N_2021);
and U3873 (N_3873,N_2371,N_2841);
or U3874 (N_3874,N_2944,N_2874);
or U3875 (N_3875,N_2939,N_2794);
and U3876 (N_3876,N_2593,N_2008);
nor U3877 (N_3877,N_2944,N_2466);
or U3878 (N_3878,N_2323,N_2226);
nor U3879 (N_3879,N_2292,N_2985);
nor U3880 (N_3880,N_2201,N_2165);
nor U3881 (N_3881,N_2683,N_2380);
nand U3882 (N_3882,N_2613,N_2587);
nand U3883 (N_3883,N_2253,N_2219);
and U3884 (N_3884,N_2767,N_2536);
nand U3885 (N_3885,N_2386,N_2075);
and U3886 (N_3886,N_2042,N_2838);
and U3887 (N_3887,N_2835,N_2443);
and U3888 (N_3888,N_2123,N_2481);
nand U3889 (N_3889,N_2177,N_2445);
nor U3890 (N_3890,N_2144,N_2899);
nand U3891 (N_3891,N_2412,N_2889);
nor U3892 (N_3892,N_2037,N_2361);
nand U3893 (N_3893,N_2792,N_2876);
nand U3894 (N_3894,N_2089,N_2447);
or U3895 (N_3895,N_2531,N_2075);
or U3896 (N_3896,N_2528,N_2688);
nor U3897 (N_3897,N_2508,N_2819);
or U3898 (N_3898,N_2052,N_2758);
nor U3899 (N_3899,N_2021,N_2677);
nor U3900 (N_3900,N_2014,N_2778);
nand U3901 (N_3901,N_2447,N_2276);
and U3902 (N_3902,N_2579,N_2028);
or U3903 (N_3903,N_2268,N_2832);
or U3904 (N_3904,N_2847,N_2484);
nand U3905 (N_3905,N_2483,N_2041);
and U3906 (N_3906,N_2420,N_2221);
nor U3907 (N_3907,N_2575,N_2375);
or U3908 (N_3908,N_2153,N_2130);
nand U3909 (N_3909,N_2459,N_2592);
and U3910 (N_3910,N_2566,N_2256);
nand U3911 (N_3911,N_2405,N_2526);
nand U3912 (N_3912,N_2464,N_2898);
nor U3913 (N_3913,N_2368,N_2806);
nor U3914 (N_3914,N_2443,N_2405);
nand U3915 (N_3915,N_2940,N_2446);
and U3916 (N_3916,N_2085,N_2122);
and U3917 (N_3917,N_2238,N_2974);
nor U3918 (N_3918,N_2906,N_2689);
nand U3919 (N_3919,N_2510,N_2151);
and U3920 (N_3920,N_2524,N_2988);
nand U3921 (N_3921,N_2249,N_2550);
and U3922 (N_3922,N_2663,N_2050);
or U3923 (N_3923,N_2370,N_2284);
and U3924 (N_3924,N_2984,N_2521);
or U3925 (N_3925,N_2914,N_2995);
nand U3926 (N_3926,N_2782,N_2681);
and U3927 (N_3927,N_2810,N_2761);
nand U3928 (N_3928,N_2182,N_2204);
nor U3929 (N_3929,N_2859,N_2714);
or U3930 (N_3930,N_2729,N_2742);
nand U3931 (N_3931,N_2554,N_2511);
or U3932 (N_3932,N_2783,N_2601);
nand U3933 (N_3933,N_2007,N_2278);
or U3934 (N_3934,N_2758,N_2143);
nor U3935 (N_3935,N_2622,N_2636);
nor U3936 (N_3936,N_2842,N_2213);
nor U3937 (N_3937,N_2932,N_2048);
nor U3938 (N_3938,N_2710,N_2295);
and U3939 (N_3939,N_2079,N_2285);
nor U3940 (N_3940,N_2580,N_2813);
nand U3941 (N_3941,N_2278,N_2412);
or U3942 (N_3942,N_2155,N_2963);
and U3943 (N_3943,N_2628,N_2634);
nor U3944 (N_3944,N_2165,N_2931);
or U3945 (N_3945,N_2530,N_2588);
nand U3946 (N_3946,N_2286,N_2799);
nand U3947 (N_3947,N_2202,N_2423);
or U3948 (N_3948,N_2068,N_2416);
nor U3949 (N_3949,N_2883,N_2521);
and U3950 (N_3950,N_2864,N_2344);
nor U3951 (N_3951,N_2540,N_2160);
nor U3952 (N_3952,N_2449,N_2056);
and U3953 (N_3953,N_2870,N_2695);
and U3954 (N_3954,N_2299,N_2064);
nand U3955 (N_3955,N_2553,N_2868);
nand U3956 (N_3956,N_2695,N_2673);
or U3957 (N_3957,N_2645,N_2340);
and U3958 (N_3958,N_2600,N_2594);
or U3959 (N_3959,N_2844,N_2895);
nand U3960 (N_3960,N_2692,N_2944);
and U3961 (N_3961,N_2044,N_2999);
nand U3962 (N_3962,N_2681,N_2509);
nand U3963 (N_3963,N_2965,N_2883);
nand U3964 (N_3964,N_2382,N_2429);
nand U3965 (N_3965,N_2005,N_2077);
or U3966 (N_3966,N_2096,N_2937);
and U3967 (N_3967,N_2369,N_2364);
nor U3968 (N_3968,N_2669,N_2876);
or U3969 (N_3969,N_2452,N_2100);
nor U3970 (N_3970,N_2406,N_2643);
and U3971 (N_3971,N_2207,N_2144);
and U3972 (N_3972,N_2252,N_2562);
nor U3973 (N_3973,N_2415,N_2247);
and U3974 (N_3974,N_2396,N_2142);
and U3975 (N_3975,N_2044,N_2164);
or U3976 (N_3976,N_2262,N_2790);
nand U3977 (N_3977,N_2926,N_2504);
nor U3978 (N_3978,N_2913,N_2797);
nand U3979 (N_3979,N_2088,N_2884);
or U3980 (N_3980,N_2264,N_2007);
nor U3981 (N_3981,N_2660,N_2011);
and U3982 (N_3982,N_2501,N_2884);
and U3983 (N_3983,N_2293,N_2299);
nand U3984 (N_3984,N_2744,N_2528);
nand U3985 (N_3985,N_2342,N_2248);
nand U3986 (N_3986,N_2222,N_2838);
nor U3987 (N_3987,N_2629,N_2907);
nand U3988 (N_3988,N_2717,N_2255);
nand U3989 (N_3989,N_2663,N_2206);
nor U3990 (N_3990,N_2724,N_2595);
nor U3991 (N_3991,N_2200,N_2725);
or U3992 (N_3992,N_2487,N_2396);
or U3993 (N_3993,N_2947,N_2394);
nor U3994 (N_3994,N_2954,N_2904);
nand U3995 (N_3995,N_2937,N_2374);
nor U3996 (N_3996,N_2671,N_2824);
and U3997 (N_3997,N_2960,N_2755);
nand U3998 (N_3998,N_2279,N_2869);
nor U3999 (N_3999,N_2335,N_2381);
nand U4000 (N_4000,N_3148,N_3874);
or U4001 (N_4001,N_3089,N_3550);
nor U4002 (N_4002,N_3633,N_3185);
nor U4003 (N_4003,N_3377,N_3733);
or U4004 (N_4004,N_3743,N_3246);
or U4005 (N_4005,N_3953,N_3435);
or U4006 (N_4006,N_3513,N_3034);
nand U4007 (N_4007,N_3121,N_3329);
or U4008 (N_4008,N_3855,N_3910);
and U4009 (N_4009,N_3208,N_3059);
nor U4010 (N_4010,N_3761,N_3697);
nand U4011 (N_4011,N_3860,N_3285);
or U4012 (N_4012,N_3713,N_3505);
and U4013 (N_4013,N_3151,N_3294);
nor U4014 (N_4014,N_3729,N_3959);
nor U4015 (N_4015,N_3841,N_3451);
nand U4016 (N_4016,N_3095,N_3493);
and U4017 (N_4017,N_3683,N_3191);
nor U4018 (N_4018,N_3409,N_3654);
or U4019 (N_4019,N_3621,N_3284);
nand U4020 (N_4020,N_3782,N_3990);
and U4021 (N_4021,N_3081,N_3873);
nor U4022 (N_4022,N_3085,N_3827);
nor U4023 (N_4023,N_3199,N_3460);
and U4024 (N_4024,N_3617,N_3615);
and U4025 (N_4025,N_3047,N_3354);
nor U4026 (N_4026,N_3883,N_3002);
and U4027 (N_4027,N_3023,N_3394);
or U4028 (N_4028,N_3964,N_3630);
nand U4029 (N_4029,N_3719,N_3061);
nand U4030 (N_4030,N_3082,N_3176);
or U4031 (N_4031,N_3888,N_3305);
nand U4032 (N_4032,N_3138,N_3295);
nand U4033 (N_4033,N_3826,N_3171);
and U4034 (N_4034,N_3359,N_3289);
nor U4035 (N_4035,N_3187,N_3226);
or U4036 (N_4036,N_3909,N_3484);
or U4037 (N_4037,N_3033,N_3932);
nand U4038 (N_4038,N_3935,N_3398);
and U4039 (N_4039,N_3358,N_3155);
nor U4040 (N_4040,N_3542,N_3991);
or U4041 (N_4041,N_3929,N_3227);
and U4042 (N_4042,N_3843,N_3390);
nand U4043 (N_4043,N_3598,N_3574);
or U4044 (N_4044,N_3596,N_3576);
or U4045 (N_4045,N_3606,N_3177);
nand U4046 (N_4046,N_3020,N_3983);
nand U4047 (N_4047,N_3568,N_3828);
and U4048 (N_4048,N_3316,N_3547);
nor U4049 (N_4049,N_3342,N_3648);
and U4050 (N_4050,N_3103,N_3355);
nand U4051 (N_4051,N_3425,N_3567);
xor U4052 (N_4052,N_3265,N_3679);
and U4053 (N_4053,N_3360,N_3677);
nor U4054 (N_4054,N_3288,N_3872);
or U4055 (N_4055,N_3689,N_3999);
nand U4056 (N_4056,N_3501,N_3702);
nor U4057 (N_4057,N_3015,N_3337);
nand U4058 (N_4058,N_3789,N_3835);
or U4059 (N_4059,N_3714,N_3041);
or U4060 (N_4060,N_3659,N_3397);
and U4061 (N_4061,N_3544,N_3796);
or U4062 (N_4062,N_3663,N_3507);
nand U4063 (N_4063,N_3192,N_3902);
and U4064 (N_4064,N_3370,N_3647);
or U4065 (N_4065,N_3092,N_3245);
nand U4066 (N_4066,N_3357,N_3980);
or U4067 (N_4067,N_3190,N_3705);
nor U4068 (N_4068,N_3086,N_3043);
nand U4069 (N_4069,N_3688,N_3462);
nor U4070 (N_4070,N_3459,N_3911);
and U4071 (N_4071,N_3139,N_3159);
nand U4072 (N_4072,N_3248,N_3477);
nor U4073 (N_4073,N_3084,N_3514);
and U4074 (N_4074,N_3637,N_3879);
or U4075 (N_4075,N_3340,N_3664);
or U4076 (N_4076,N_3896,N_3449);
or U4077 (N_4077,N_3261,N_3077);
and U4078 (N_4078,N_3282,N_3699);
nand U4079 (N_4079,N_3941,N_3299);
nor U4080 (N_4080,N_3853,N_3848);
nand U4081 (N_4081,N_3231,N_3430);
and U4082 (N_4082,N_3625,N_3816);
or U4083 (N_4083,N_3427,N_3587);
or U4084 (N_4084,N_3785,N_3160);
nor U4085 (N_4085,N_3921,N_3952);
or U4086 (N_4086,N_3846,N_3384);
nor U4087 (N_4087,N_3283,N_3476);
nor U4088 (N_4088,N_3586,N_3483);
nand U4089 (N_4089,N_3150,N_3751);
nor U4090 (N_4090,N_3209,N_3157);
nor U4091 (N_4091,N_3399,N_3642);
and U4092 (N_4092,N_3413,N_3000);
or U4093 (N_4093,N_3831,N_3161);
nor U4094 (N_4094,N_3410,N_3250);
nor U4095 (N_4095,N_3037,N_3017);
and U4096 (N_4096,N_3611,N_3931);
and U4097 (N_4097,N_3525,N_3099);
or U4098 (N_4098,N_3812,N_3717);
or U4099 (N_4099,N_3808,N_3680);
and U4100 (N_4100,N_3762,N_3656);
nor U4101 (N_4101,N_3984,N_3318);
nor U4102 (N_4102,N_3535,N_3122);
and U4103 (N_4103,N_3727,N_3442);
nand U4104 (N_4104,N_3135,N_3113);
and U4105 (N_4105,N_3035,N_3987);
nand U4106 (N_4106,N_3403,N_3842);
nand U4107 (N_4107,N_3876,N_3572);
or U4108 (N_4108,N_3523,N_3710);
nor U4109 (N_4109,N_3806,N_3054);
or U4110 (N_4110,N_3118,N_3040);
nor U4111 (N_4111,N_3454,N_3251);
or U4112 (N_4112,N_3492,N_3439);
and U4113 (N_4113,N_3036,N_3373);
nand U4114 (N_4114,N_3752,N_3830);
or U4115 (N_4115,N_3406,N_3453);
xor U4116 (N_4116,N_3346,N_3850);
nand U4117 (N_4117,N_3924,N_3787);
or U4118 (N_4118,N_3629,N_3276);
and U4119 (N_4119,N_3693,N_3686);
or U4120 (N_4120,N_3700,N_3788);
and U4121 (N_4121,N_3331,N_3851);
and U4122 (N_4122,N_3549,N_3087);
nand U4123 (N_4123,N_3708,N_3170);
and U4124 (N_4124,N_3319,N_3109);
and U4125 (N_4125,N_3973,N_3458);
nor U4126 (N_4126,N_3298,N_3774);
and U4127 (N_4127,N_3821,N_3076);
and U4128 (N_4128,N_3858,N_3676);
or U4129 (N_4129,N_3703,N_3071);
nor U4130 (N_4130,N_3731,N_3420);
nor U4131 (N_4131,N_3770,N_3213);
and U4132 (N_4132,N_3039,N_3595);
or U4133 (N_4133,N_3589,N_3438);
nor U4134 (N_4134,N_3134,N_3417);
nor U4135 (N_4135,N_3739,N_3506);
or U4136 (N_4136,N_3508,N_3375);
nand U4137 (N_4137,N_3877,N_3936);
or U4138 (N_4138,N_3829,N_3105);
nor U4139 (N_4139,N_3728,N_3019);
nand U4140 (N_4140,N_3402,N_3067);
nor U4141 (N_4141,N_3181,N_3328);
nand U4142 (N_4142,N_3669,N_3950);
nor U4143 (N_4143,N_3602,N_3186);
and U4144 (N_4144,N_3674,N_3125);
nand U4145 (N_4145,N_3008,N_3075);
or U4146 (N_4146,N_3107,N_3562);
and U4147 (N_4147,N_3856,N_3545);
nand U4148 (N_4148,N_3579,N_3238);
nor U4149 (N_4149,N_3901,N_3379);
or U4150 (N_4150,N_3783,N_3098);
nor U4151 (N_4151,N_3519,N_3638);
or U4152 (N_4152,N_3396,N_3775);
and U4153 (N_4153,N_3893,N_3264);
and U4154 (N_4154,N_3124,N_3303);
or U4155 (N_4155,N_3204,N_3599);
and U4156 (N_4156,N_3297,N_3322);
and U4157 (N_4157,N_3947,N_3368);
nand U4158 (N_4158,N_3694,N_3600);
nor U4159 (N_4159,N_3978,N_3854);
nor U4160 (N_4160,N_3259,N_3912);
nand U4161 (N_4161,N_3960,N_3064);
nor U4162 (N_4162,N_3369,N_3534);
nor U4163 (N_4163,N_3045,N_3010);
nor U4164 (N_4164,N_3429,N_3012);
nand U4165 (N_4165,N_3018,N_3715);
nand U4166 (N_4166,N_3169,N_3175);
nand U4167 (N_4167,N_3044,N_3604);
or U4168 (N_4168,N_3051,N_3293);
nand U4169 (N_4169,N_3003,N_3217);
nand U4170 (N_4170,N_3884,N_3287);
or U4171 (N_4171,N_3096,N_3024);
nand U4172 (N_4172,N_3543,N_3053);
nand U4173 (N_4173,N_3378,N_3117);
nand U4174 (N_4174,N_3777,N_3533);
nand U4175 (N_4175,N_3132,N_3334);
and U4176 (N_4176,N_3652,N_3823);
or U4177 (N_4177,N_3274,N_3339);
or U4178 (N_4178,N_3363,N_3026);
nor U4179 (N_4179,N_3661,N_3471);
and U4180 (N_4180,N_3690,N_3495);
or U4181 (N_4181,N_3641,N_3174);
nor U4182 (N_4182,N_3895,N_3233);
or U4183 (N_4183,N_3401,N_3809);
and U4184 (N_4184,N_3223,N_3740);
nor U4185 (N_4185,N_3021,N_3046);
nor U4186 (N_4186,N_3219,N_3620);
or U4187 (N_4187,N_3701,N_3852);
and U4188 (N_4188,N_3296,N_3867);
nor U4189 (N_4189,N_3336,N_3210);
nor U4190 (N_4190,N_3166,N_3063);
and U4191 (N_4191,N_3509,N_3801);
or U4192 (N_4192,N_3865,N_3381);
nand U4193 (N_4193,N_3200,N_3335);
and U4194 (N_4194,N_3490,N_3531);
nand U4195 (N_4195,N_3738,N_3685);
nand U4196 (N_4196,N_3764,N_3382);
nand U4197 (N_4197,N_3315,N_3927);
or U4198 (N_4198,N_3861,N_3609);
nand U4199 (N_4199,N_3093,N_3147);
or U4200 (N_4200,N_3455,N_3466);
and U4201 (N_4201,N_3309,N_3206);
nor U4202 (N_4202,N_3112,N_3943);
or U4203 (N_4203,N_3262,N_3247);
or U4204 (N_4204,N_3726,N_3388);
nor U4205 (N_4205,N_3120,N_3280);
or U4206 (N_4206,N_3904,N_3243);
and U4207 (N_4207,N_3769,N_3807);
or U4208 (N_4208,N_3108,N_3193);
and U4209 (N_4209,N_3349,N_3997);
or U4210 (N_4210,N_3446,N_3716);
nand U4211 (N_4211,N_3474,N_3958);
or U4212 (N_4212,N_3326,N_3042);
nor U4213 (N_4213,N_3825,N_3392);
nor U4214 (N_4214,N_3797,N_3682);
and U4215 (N_4215,N_3452,N_3144);
or U4216 (N_4216,N_3754,N_3269);
or U4217 (N_4217,N_3167,N_3836);
and U4218 (N_4218,N_3189,N_3838);
or U4219 (N_4219,N_3324,N_3989);
and U4220 (N_4220,N_3591,N_3091);
nand U4221 (N_4221,N_3753,N_3998);
or U4222 (N_4222,N_3773,N_3344);
and U4223 (N_4223,N_3750,N_3308);
nor U4224 (N_4224,N_3635,N_3944);
or U4225 (N_4225,N_3969,N_3919);
and U4226 (N_4226,N_3651,N_3485);
or U4227 (N_4227,N_3814,N_3639);
nor U4228 (N_4228,N_3057,N_3445);
and U4229 (N_4229,N_3131,N_3317);
and U4230 (N_4230,N_3657,N_3619);
nor U4231 (N_4231,N_3428,N_3553);
nor U4232 (N_4232,N_3992,N_3746);
nor U4233 (N_4233,N_3300,N_3491);
or U4234 (N_4234,N_3631,N_3526);
or U4235 (N_4235,N_3291,N_3791);
nand U4236 (N_4236,N_3815,N_3073);
or U4237 (N_4237,N_3468,N_3756);
nor U4238 (N_4238,N_3271,N_3563);
nand U4239 (N_4239,N_3302,N_3456);
nand U4240 (N_4240,N_3128,N_3594);
and U4241 (N_4241,N_3424,N_3049);
and U4242 (N_4242,N_3031,N_3870);
or U4243 (N_4243,N_3882,N_3421);
nor U4244 (N_4244,N_3802,N_3312);
nand U4245 (N_4245,N_3025,N_3266);
xnor U4246 (N_4246,N_3470,N_3301);
or U4247 (N_4247,N_3878,N_3152);
or U4248 (N_4248,N_3951,N_3643);
nor U4249 (N_4249,N_3706,N_3644);
or U4250 (N_4250,N_3779,N_3325);
nand U4251 (N_4251,N_3433,N_3062);
xnor U4252 (N_4252,N_3432,N_3130);
nor U4253 (N_4253,N_3320,N_3937);
or U4254 (N_4254,N_3968,N_3862);
nand U4255 (N_4255,N_3938,N_3803);
or U4256 (N_4256,N_3709,N_3903);
and U4257 (N_4257,N_3163,N_3899);
or U4258 (N_4258,N_3994,N_3955);
nor U4259 (N_4259,N_3793,N_3143);
nand U4260 (N_4260,N_3240,N_3646);
or U4261 (N_4261,N_3055,N_3725);
and U4262 (N_4262,N_3934,N_3536);
or U4263 (N_4263,N_3292,N_3556);
and U4264 (N_4264,N_3886,N_3624);
or U4265 (N_4265,N_3168,N_3497);
and U4266 (N_4266,N_3343,N_3281);
and U4267 (N_4267,N_3707,N_3612);
nand U4268 (N_4268,N_3634,N_3418);
or U4269 (N_4269,N_3006,N_3141);
and U4270 (N_4270,N_3557,N_3173);
and U4271 (N_4271,N_3792,N_3083);
nand U4272 (N_4272,N_3088,N_3555);
nand U4273 (N_4273,N_3172,N_3583);
nor U4274 (N_4274,N_3577,N_3404);
or U4275 (N_4275,N_3016,N_3214);
nor U4276 (N_4276,N_3887,N_3444);
nand U4277 (N_4277,N_3760,N_3662);
nor U4278 (N_4278,N_3972,N_3195);
and U4279 (N_4279,N_3653,N_3772);
nor U4280 (N_4280,N_3183,N_3440);
nand U4281 (N_4281,N_3804,N_3154);
and U4282 (N_4282,N_3528,N_3580);
or U4283 (N_4283,N_3673,N_3670);
or U4284 (N_4284,N_3718,N_3957);
nand U4285 (N_4285,N_3352,N_3530);
nand U4286 (N_4286,N_3178,N_3573);
nand U4287 (N_4287,N_3126,N_3748);
xor U4288 (N_4288,N_3962,N_3362);
nor U4289 (N_4289,N_3211,N_3857);
nand U4290 (N_4290,N_3529,N_3672);
nand U4291 (N_4291,N_3977,N_3660);
nand U4292 (N_4292,N_3832,N_3948);
or U4293 (N_4293,N_3307,N_3869);
and U4294 (N_4294,N_3868,N_3153);
nor U4295 (N_4295,N_3228,N_3982);
nand U4296 (N_4296,N_3696,N_3817);
or U4297 (N_4297,N_3052,N_3711);
nand U4298 (N_4298,N_3845,N_3389);
or U4299 (N_4299,N_3133,N_3350);
or U4300 (N_4300,N_3640,N_3256);
nor U4301 (N_4301,N_3464,N_3614);
nand U4302 (N_4302,N_3314,N_3482);
or U4303 (N_4303,N_3945,N_3400);
nor U4304 (N_4304,N_3005,N_3813);
nor U4305 (N_4305,N_3747,N_3881);
and U4306 (N_4306,N_3837,N_3116);
or U4307 (N_4307,N_3844,N_3437);
or U4308 (N_4308,N_3889,N_3221);
nor U4309 (N_4309,N_3100,N_3201);
xnor U4310 (N_4310,N_3759,N_3111);
nor U4311 (N_4311,N_3188,N_3650);
nor U4312 (N_4312,N_3165,N_3922);
or U4313 (N_4313,N_3078,N_3794);
nor U4314 (N_4314,N_3559,N_3203);
or U4315 (N_4315,N_3423,N_3028);
or U4316 (N_4316,N_3007,N_3665);
nor U4317 (N_4317,N_3578,N_3541);
or U4318 (N_4318,N_3918,N_3601);
or U4319 (N_4319,N_3494,N_3613);
and U4320 (N_4320,N_3949,N_3561);
and U4321 (N_4321,N_3330,N_3074);
nand U4322 (N_4322,N_3741,N_3839);
and U4323 (N_4323,N_3332,N_3110);
nor U4324 (N_4324,N_3383,N_3610);
or U4325 (N_4325,N_3900,N_3875);
or U4326 (N_4326,N_3755,N_3765);
nor U4327 (N_4327,N_3940,N_3441);
nor U4328 (N_4328,N_3487,N_3894);
and U4329 (N_4329,N_3811,N_3942);
nor U4330 (N_4330,N_3871,N_3735);
nor U4331 (N_4331,N_3162,N_3058);
xor U4332 (N_4332,N_3372,N_3627);
nand U4333 (N_4333,N_3515,N_3333);
or U4334 (N_4334,N_3304,N_3926);
nand U4335 (N_4335,N_3197,N_3608);
nor U4336 (N_4336,N_3554,N_3684);
nand U4337 (N_4337,N_3510,N_3222);
nand U4338 (N_4338,N_3119,N_3560);
or U4339 (N_4339,N_3179,N_3207);
nor U4340 (N_4340,N_3503,N_3618);
or U4341 (N_4341,N_3564,N_3478);
or U4342 (N_4342,N_3890,N_3205);
nor U4343 (N_4343,N_3180,N_3498);
or U4344 (N_4344,N_3475,N_3695);
and U4345 (N_4345,N_3575,N_3986);
nor U4346 (N_4346,N_3450,N_3742);
and U4347 (N_4347,N_3405,N_3101);
nand U4348 (N_4348,N_3414,N_3824);
and U4349 (N_4349,N_3338,N_3744);
nor U4350 (N_4350,N_3249,N_3781);
nand U4351 (N_4351,N_3834,N_3353);
and U4352 (N_4352,N_3242,N_3898);
or U4353 (N_4353,N_3778,N_3540);
nand U4354 (N_4354,N_3009,N_3011);
or U4355 (N_4355,N_3897,N_3798);
or U4356 (N_4356,N_3473,N_3720);
and U4357 (N_4357,N_3571,N_3066);
nand U4358 (N_4358,N_3780,N_3833);
nand U4359 (N_4359,N_3230,N_3645);
or U4360 (N_4360,N_3202,N_3232);
nor U4361 (N_4361,N_3916,N_3480);
nand U4362 (N_4362,N_3253,N_3102);
nand U4363 (N_4363,N_3056,N_3521);
or U4364 (N_4364,N_3115,N_3094);
and U4365 (N_4365,N_3146,N_3722);
nor U4366 (N_4366,N_3810,N_3415);
or U4367 (N_4367,N_3757,N_3065);
and U4368 (N_4368,N_3907,N_3422);
nor U4369 (N_4369,N_3395,N_3588);
or U4370 (N_4370,N_3649,N_3374);
and U4371 (N_4371,N_3979,N_3391);
nand U4372 (N_4372,N_3582,N_3022);
nor U4373 (N_4373,N_3784,N_3849);
and U4374 (N_4374,N_3447,N_3551);
or U4375 (N_4375,N_3323,N_3668);
or U4376 (N_4376,N_3981,N_3114);
and U4377 (N_4377,N_3408,N_3412);
or U4378 (N_4378,N_3182,N_3196);
and U4379 (N_4379,N_3623,N_3140);
and U4380 (N_4380,N_3767,N_3723);
and U4381 (N_4381,N_3229,N_3255);
and U4382 (N_4382,N_3822,N_3286);
nor U4383 (N_4383,N_3995,N_3516);
and U4384 (N_4384,N_3149,N_3988);
nand U4385 (N_4385,N_3434,N_3671);
nand U4386 (N_4386,N_3463,N_3527);
nor U4387 (N_4387,N_3268,N_3393);
nand U4388 (N_4388,N_3137,N_3260);
nor U4389 (N_4389,N_3306,N_3499);
and U4390 (N_4390,N_3345,N_3520);
nand U4391 (N_4391,N_3080,N_3616);
and U4392 (N_4392,N_3361,N_3687);
or U4393 (N_4393,N_3467,N_3603);
or U4394 (N_4394,N_3001,N_3419);
and U4395 (N_4395,N_3313,N_3275);
or U4396 (N_4396,N_3819,N_3164);
nand U4397 (N_4397,N_3636,N_3489);
and U4398 (N_4398,N_3277,N_3786);
nor U4399 (N_4399,N_3795,N_3736);
nand U4400 (N_4400,N_3348,N_3917);
or U4401 (N_4401,N_3675,N_3776);
nor U4402 (N_4402,N_3258,N_3704);
nor U4403 (N_4403,N_3538,N_3605);
nor U4404 (N_4404,N_3771,N_3698);
or U4405 (N_4405,N_3431,N_3129);
nand U4406 (N_4406,N_3278,N_3517);
and U4407 (N_4407,N_3481,N_3993);
or U4408 (N_4408,N_3558,N_3939);
nor U4409 (N_4409,N_3267,N_3273);
nor U4410 (N_4410,N_3050,N_3593);
and U4411 (N_4411,N_3892,N_3351);
or U4412 (N_4412,N_3224,N_3436);
and U4413 (N_4413,N_3263,N_3946);
nand U4414 (N_4414,N_3570,N_3970);
or U4415 (N_4415,N_3565,N_3607);
nor U4416 (N_4416,N_3090,N_3626);
or U4417 (N_4417,N_3681,N_3691);
or U4418 (N_4418,N_3236,N_3863);
nor U4419 (N_4419,N_3965,N_3472);
nor U4420 (N_4420,N_3145,N_3749);
and U4421 (N_4421,N_3581,N_3371);
and U4422 (N_4422,N_3511,N_3321);
and U4423 (N_4423,N_3522,N_3766);
or U4424 (N_4424,N_3244,N_3730);
nor U4425 (N_4425,N_3678,N_3539);
nand U4426 (N_4426,N_3241,N_3237);
nand U4427 (N_4427,N_3079,N_3257);
nor U4428 (N_4428,N_3272,N_3628);
and U4429 (N_4429,N_3225,N_3212);
nor U4430 (N_4430,N_3859,N_3566);
and U4431 (N_4431,N_3768,N_3504);
or U4432 (N_4432,N_3500,N_3805);
nor U4433 (N_4433,N_3127,N_3818);
nor U4434 (N_4434,N_3961,N_3584);
nand U4435 (N_4435,N_3448,N_3758);
and U4436 (N_4436,N_3518,N_3254);
or U4437 (N_4437,N_3915,N_3104);
nand U4438 (N_4438,N_3880,N_3465);
or U4439 (N_4439,N_3763,N_3032);
or U4440 (N_4440,N_3956,N_3799);
or U4441 (N_4441,N_3158,N_3097);
nand U4442 (N_4442,N_3597,N_3220);
nor U4443 (N_4443,N_3908,N_3667);
and U4444 (N_4444,N_3732,N_3411);
nor U4445 (N_4445,N_3790,N_3341);
nor U4446 (N_4446,N_3386,N_3234);
or U4447 (N_4447,N_3712,N_3347);
or U4448 (N_4448,N_3933,N_3745);
or U4449 (N_4449,N_3479,N_3840);
nand U4450 (N_4450,N_3928,N_3996);
nor U4451 (N_4451,N_3367,N_3443);
nor U4452 (N_4452,N_3038,N_3048);
and U4453 (N_4453,N_3914,N_3971);
nand U4454 (N_4454,N_3800,N_3327);
nor U4455 (N_4455,N_3366,N_3954);
nand U4456 (N_4456,N_3885,N_3569);
nor U4457 (N_4457,N_3029,N_3235);
or U4458 (N_4458,N_3546,N_3537);
nor U4459 (N_4459,N_3365,N_3820);
or U4460 (N_4460,N_3734,N_3486);
nand U4461 (N_4461,N_3279,N_3974);
and U4462 (N_4462,N_3311,N_3461);
nor U4463 (N_4463,N_3385,N_3290);
and U4464 (N_4464,N_3407,N_3585);
nor U4465 (N_4465,N_3512,N_3905);
and U4466 (N_4466,N_3496,N_3072);
and U4467 (N_4467,N_3364,N_3976);
nand U4468 (N_4468,N_3724,N_3218);
and U4469 (N_4469,N_3142,N_3030);
nor U4470 (N_4470,N_3975,N_3060);
nand U4471 (N_4471,N_3963,N_3488);
or U4472 (N_4472,N_3069,N_3891);
nand U4473 (N_4473,N_3070,N_3913);
or U4474 (N_4474,N_3156,N_3966);
or U4475 (N_4475,N_3590,N_3270);
and U4476 (N_4476,N_3906,N_3136);
nor U4477 (N_4477,N_3387,N_3502);
nand U4478 (N_4478,N_3655,N_3721);
or U4479 (N_4479,N_3923,N_3524);
nand U4480 (N_4480,N_3457,N_3622);
or U4481 (N_4481,N_3239,N_3198);
nor U4482 (N_4482,N_3215,N_3310);
and U4483 (N_4483,N_3632,N_3666);
or U4484 (N_4484,N_3967,N_3548);
nand U4485 (N_4485,N_3737,N_3004);
or U4486 (N_4486,N_3106,N_3985);
nor U4487 (N_4487,N_3068,N_3184);
and U4488 (N_4488,N_3426,N_3864);
nand U4489 (N_4489,N_3925,N_3552);
nand U4490 (N_4490,N_3252,N_3356);
nor U4491 (N_4491,N_3920,N_3692);
nand U4492 (N_4492,N_3014,N_3123);
nor U4493 (N_4493,N_3376,N_3866);
and U4494 (N_4494,N_3216,N_3469);
or U4495 (N_4495,N_3380,N_3658);
nand U4496 (N_4496,N_3532,N_3416);
nor U4497 (N_4497,N_3194,N_3013);
and U4498 (N_4498,N_3930,N_3847);
or U4499 (N_4499,N_3592,N_3027);
nand U4500 (N_4500,N_3894,N_3745);
nor U4501 (N_4501,N_3358,N_3798);
nand U4502 (N_4502,N_3040,N_3513);
or U4503 (N_4503,N_3227,N_3947);
and U4504 (N_4504,N_3667,N_3755);
nor U4505 (N_4505,N_3396,N_3002);
and U4506 (N_4506,N_3574,N_3298);
and U4507 (N_4507,N_3594,N_3873);
and U4508 (N_4508,N_3199,N_3431);
nor U4509 (N_4509,N_3049,N_3865);
or U4510 (N_4510,N_3654,N_3562);
nand U4511 (N_4511,N_3880,N_3138);
nor U4512 (N_4512,N_3325,N_3079);
nand U4513 (N_4513,N_3177,N_3599);
nor U4514 (N_4514,N_3211,N_3699);
or U4515 (N_4515,N_3530,N_3273);
nand U4516 (N_4516,N_3547,N_3886);
and U4517 (N_4517,N_3251,N_3162);
nor U4518 (N_4518,N_3259,N_3955);
and U4519 (N_4519,N_3084,N_3451);
and U4520 (N_4520,N_3948,N_3258);
or U4521 (N_4521,N_3330,N_3284);
nor U4522 (N_4522,N_3660,N_3104);
or U4523 (N_4523,N_3233,N_3556);
nand U4524 (N_4524,N_3490,N_3680);
and U4525 (N_4525,N_3453,N_3991);
or U4526 (N_4526,N_3944,N_3267);
nor U4527 (N_4527,N_3384,N_3316);
and U4528 (N_4528,N_3803,N_3997);
nor U4529 (N_4529,N_3597,N_3630);
or U4530 (N_4530,N_3443,N_3126);
nand U4531 (N_4531,N_3900,N_3812);
and U4532 (N_4532,N_3346,N_3322);
nand U4533 (N_4533,N_3223,N_3574);
and U4534 (N_4534,N_3725,N_3810);
or U4535 (N_4535,N_3794,N_3870);
nand U4536 (N_4536,N_3151,N_3694);
and U4537 (N_4537,N_3080,N_3499);
nand U4538 (N_4538,N_3782,N_3351);
or U4539 (N_4539,N_3164,N_3003);
nor U4540 (N_4540,N_3366,N_3837);
nor U4541 (N_4541,N_3226,N_3902);
nand U4542 (N_4542,N_3296,N_3975);
and U4543 (N_4543,N_3523,N_3554);
or U4544 (N_4544,N_3700,N_3828);
nor U4545 (N_4545,N_3532,N_3474);
and U4546 (N_4546,N_3062,N_3244);
nor U4547 (N_4547,N_3302,N_3473);
nand U4548 (N_4548,N_3052,N_3462);
or U4549 (N_4549,N_3905,N_3837);
nand U4550 (N_4550,N_3520,N_3148);
nor U4551 (N_4551,N_3097,N_3175);
nand U4552 (N_4552,N_3935,N_3644);
nor U4553 (N_4553,N_3267,N_3556);
nand U4554 (N_4554,N_3626,N_3173);
nand U4555 (N_4555,N_3086,N_3180);
and U4556 (N_4556,N_3350,N_3561);
or U4557 (N_4557,N_3641,N_3674);
and U4558 (N_4558,N_3898,N_3393);
and U4559 (N_4559,N_3295,N_3475);
and U4560 (N_4560,N_3284,N_3837);
nor U4561 (N_4561,N_3586,N_3822);
or U4562 (N_4562,N_3365,N_3770);
or U4563 (N_4563,N_3759,N_3344);
nor U4564 (N_4564,N_3049,N_3257);
or U4565 (N_4565,N_3096,N_3135);
and U4566 (N_4566,N_3255,N_3614);
nor U4567 (N_4567,N_3264,N_3107);
or U4568 (N_4568,N_3710,N_3588);
nand U4569 (N_4569,N_3191,N_3034);
nor U4570 (N_4570,N_3853,N_3009);
or U4571 (N_4571,N_3410,N_3302);
or U4572 (N_4572,N_3545,N_3531);
or U4573 (N_4573,N_3610,N_3709);
and U4574 (N_4574,N_3522,N_3017);
or U4575 (N_4575,N_3005,N_3458);
nor U4576 (N_4576,N_3516,N_3129);
nand U4577 (N_4577,N_3909,N_3443);
and U4578 (N_4578,N_3006,N_3425);
or U4579 (N_4579,N_3050,N_3679);
or U4580 (N_4580,N_3716,N_3096);
nand U4581 (N_4581,N_3852,N_3142);
nand U4582 (N_4582,N_3502,N_3461);
nand U4583 (N_4583,N_3823,N_3534);
nor U4584 (N_4584,N_3344,N_3139);
nand U4585 (N_4585,N_3925,N_3015);
nand U4586 (N_4586,N_3340,N_3778);
or U4587 (N_4587,N_3429,N_3538);
and U4588 (N_4588,N_3616,N_3421);
or U4589 (N_4589,N_3108,N_3855);
nand U4590 (N_4590,N_3506,N_3578);
or U4591 (N_4591,N_3838,N_3869);
nand U4592 (N_4592,N_3306,N_3646);
nor U4593 (N_4593,N_3940,N_3261);
xor U4594 (N_4594,N_3282,N_3875);
nor U4595 (N_4595,N_3147,N_3699);
and U4596 (N_4596,N_3600,N_3588);
and U4597 (N_4597,N_3172,N_3610);
and U4598 (N_4598,N_3771,N_3438);
nand U4599 (N_4599,N_3145,N_3192);
nand U4600 (N_4600,N_3995,N_3082);
and U4601 (N_4601,N_3448,N_3747);
or U4602 (N_4602,N_3050,N_3834);
nand U4603 (N_4603,N_3363,N_3284);
nand U4604 (N_4604,N_3307,N_3320);
nand U4605 (N_4605,N_3798,N_3002);
and U4606 (N_4606,N_3609,N_3221);
and U4607 (N_4607,N_3125,N_3325);
or U4608 (N_4608,N_3610,N_3826);
and U4609 (N_4609,N_3067,N_3276);
nand U4610 (N_4610,N_3889,N_3576);
nand U4611 (N_4611,N_3207,N_3966);
and U4612 (N_4612,N_3239,N_3921);
nor U4613 (N_4613,N_3121,N_3071);
nand U4614 (N_4614,N_3311,N_3157);
nand U4615 (N_4615,N_3153,N_3407);
nand U4616 (N_4616,N_3732,N_3927);
nand U4617 (N_4617,N_3786,N_3677);
nand U4618 (N_4618,N_3316,N_3430);
and U4619 (N_4619,N_3640,N_3989);
or U4620 (N_4620,N_3733,N_3254);
nor U4621 (N_4621,N_3307,N_3922);
or U4622 (N_4622,N_3900,N_3016);
or U4623 (N_4623,N_3045,N_3336);
and U4624 (N_4624,N_3018,N_3220);
or U4625 (N_4625,N_3941,N_3105);
and U4626 (N_4626,N_3468,N_3758);
and U4627 (N_4627,N_3336,N_3496);
and U4628 (N_4628,N_3765,N_3313);
nand U4629 (N_4629,N_3586,N_3882);
nor U4630 (N_4630,N_3392,N_3086);
and U4631 (N_4631,N_3696,N_3478);
nor U4632 (N_4632,N_3036,N_3298);
nor U4633 (N_4633,N_3088,N_3992);
or U4634 (N_4634,N_3758,N_3387);
xnor U4635 (N_4635,N_3651,N_3901);
nand U4636 (N_4636,N_3472,N_3637);
and U4637 (N_4637,N_3927,N_3004);
and U4638 (N_4638,N_3196,N_3060);
xor U4639 (N_4639,N_3151,N_3308);
nor U4640 (N_4640,N_3011,N_3879);
nor U4641 (N_4641,N_3666,N_3612);
and U4642 (N_4642,N_3554,N_3113);
nor U4643 (N_4643,N_3018,N_3060);
or U4644 (N_4644,N_3049,N_3061);
nor U4645 (N_4645,N_3133,N_3972);
nor U4646 (N_4646,N_3884,N_3861);
nor U4647 (N_4647,N_3740,N_3019);
and U4648 (N_4648,N_3387,N_3192);
and U4649 (N_4649,N_3111,N_3477);
and U4650 (N_4650,N_3714,N_3264);
nand U4651 (N_4651,N_3013,N_3719);
nand U4652 (N_4652,N_3533,N_3998);
or U4653 (N_4653,N_3060,N_3809);
or U4654 (N_4654,N_3299,N_3187);
nand U4655 (N_4655,N_3277,N_3446);
and U4656 (N_4656,N_3421,N_3643);
nor U4657 (N_4657,N_3902,N_3420);
and U4658 (N_4658,N_3881,N_3584);
or U4659 (N_4659,N_3904,N_3675);
and U4660 (N_4660,N_3388,N_3555);
and U4661 (N_4661,N_3779,N_3202);
nand U4662 (N_4662,N_3747,N_3007);
and U4663 (N_4663,N_3397,N_3561);
nand U4664 (N_4664,N_3554,N_3685);
nor U4665 (N_4665,N_3091,N_3965);
or U4666 (N_4666,N_3318,N_3780);
and U4667 (N_4667,N_3164,N_3288);
nor U4668 (N_4668,N_3472,N_3080);
nor U4669 (N_4669,N_3572,N_3357);
nand U4670 (N_4670,N_3051,N_3829);
or U4671 (N_4671,N_3875,N_3446);
and U4672 (N_4672,N_3802,N_3773);
and U4673 (N_4673,N_3300,N_3380);
nor U4674 (N_4674,N_3665,N_3921);
or U4675 (N_4675,N_3988,N_3991);
and U4676 (N_4676,N_3611,N_3229);
and U4677 (N_4677,N_3414,N_3403);
nor U4678 (N_4678,N_3481,N_3063);
nand U4679 (N_4679,N_3760,N_3201);
nor U4680 (N_4680,N_3235,N_3748);
nand U4681 (N_4681,N_3791,N_3230);
nand U4682 (N_4682,N_3665,N_3331);
or U4683 (N_4683,N_3613,N_3826);
nor U4684 (N_4684,N_3117,N_3040);
nor U4685 (N_4685,N_3836,N_3372);
nand U4686 (N_4686,N_3444,N_3216);
or U4687 (N_4687,N_3996,N_3027);
nor U4688 (N_4688,N_3386,N_3491);
nor U4689 (N_4689,N_3600,N_3890);
nand U4690 (N_4690,N_3723,N_3274);
nor U4691 (N_4691,N_3478,N_3866);
nor U4692 (N_4692,N_3973,N_3165);
nand U4693 (N_4693,N_3696,N_3561);
or U4694 (N_4694,N_3537,N_3805);
nand U4695 (N_4695,N_3423,N_3311);
nor U4696 (N_4696,N_3570,N_3416);
nor U4697 (N_4697,N_3257,N_3205);
nand U4698 (N_4698,N_3462,N_3977);
or U4699 (N_4699,N_3935,N_3622);
or U4700 (N_4700,N_3887,N_3214);
xor U4701 (N_4701,N_3240,N_3377);
and U4702 (N_4702,N_3938,N_3278);
nand U4703 (N_4703,N_3318,N_3268);
or U4704 (N_4704,N_3583,N_3392);
nor U4705 (N_4705,N_3777,N_3486);
nand U4706 (N_4706,N_3095,N_3715);
nand U4707 (N_4707,N_3132,N_3556);
or U4708 (N_4708,N_3356,N_3803);
or U4709 (N_4709,N_3884,N_3799);
xor U4710 (N_4710,N_3487,N_3742);
nor U4711 (N_4711,N_3529,N_3105);
or U4712 (N_4712,N_3985,N_3716);
nor U4713 (N_4713,N_3848,N_3836);
or U4714 (N_4714,N_3757,N_3419);
nand U4715 (N_4715,N_3750,N_3289);
nor U4716 (N_4716,N_3872,N_3159);
nand U4717 (N_4717,N_3713,N_3997);
nand U4718 (N_4718,N_3334,N_3711);
and U4719 (N_4719,N_3269,N_3222);
and U4720 (N_4720,N_3400,N_3099);
or U4721 (N_4721,N_3954,N_3175);
or U4722 (N_4722,N_3403,N_3549);
nand U4723 (N_4723,N_3667,N_3693);
nand U4724 (N_4724,N_3551,N_3400);
or U4725 (N_4725,N_3495,N_3171);
or U4726 (N_4726,N_3493,N_3082);
and U4727 (N_4727,N_3566,N_3953);
and U4728 (N_4728,N_3489,N_3979);
nand U4729 (N_4729,N_3141,N_3285);
or U4730 (N_4730,N_3669,N_3077);
nand U4731 (N_4731,N_3790,N_3147);
xor U4732 (N_4732,N_3850,N_3521);
or U4733 (N_4733,N_3366,N_3746);
or U4734 (N_4734,N_3533,N_3627);
and U4735 (N_4735,N_3774,N_3731);
nor U4736 (N_4736,N_3229,N_3591);
nor U4737 (N_4737,N_3180,N_3523);
and U4738 (N_4738,N_3305,N_3041);
nand U4739 (N_4739,N_3165,N_3279);
or U4740 (N_4740,N_3744,N_3750);
nand U4741 (N_4741,N_3624,N_3638);
or U4742 (N_4742,N_3551,N_3850);
nor U4743 (N_4743,N_3375,N_3422);
or U4744 (N_4744,N_3219,N_3439);
and U4745 (N_4745,N_3089,N_3519);
or U4746 (N_4746,N_3641,N_3952);
or U4747 (N_4747,N_3506,N_3323);
nor U4748 (N_4748,N_3017,N_3176);
or U4749 (N_4749,N_3460,N_3844);
or U4750 (N_4750,N_3934,N_3115);
and U4751 (N_4751,N_3293,N_3182);
nand U4752 (N_4752,N_3444,N_3150);
xnor U4753 (N_4753,N_3788,N_3689);
nor U4754 (N_4754,N_3107,N_3145);
nor U4755 (N_4755,N_3409,N_3038);
nand U4756 (N_4756,N_3958,N_3026);
or U4757 (N_4757,N_3165,N_3240);
and U4758 (N_4758,N_3329,N_3968);
or U4759 (N_4759,N_3674,N_3717);
or U4760 (N_4760,N_3494,N_3188);
nand U4761 (N_4761,N_3869,N_3393);
or U4762 (N_4762,N_3205,N_3789);
nand U4763 (N_4763,N_3316,N_3579);
nor U4764 (N_4764,N_3690,N_3888);
and U4765 (N_4765,N_3731,N_3456);
nor U4766 (N_4766,N_3036,N_3141);
nor U4767 (N_4767,N_3801,N_3035);
or U4768 (N_4768,N_3185,N_3852);
or U4769 (N_4769,N_3562,N_3006);
and U4770 (N_4770,N_3669,N_3640);
nand U4771 (N_4771,N_3753,N_3449);
nand U4772 (N_4772,N_3599,N_3396);
nand U4773 (N_4773,N_3962,N_3536);
or U4774 (N_4774,N_3168,N_3387);
nand U4775 (N_4775,N_3459,N_3252);
nand U4776 (N_4776,N_3948,N_3072);
and U4777 (N_4777,N_3642,N_3978);
and U4778 (N_4778,N_3468,N_3783);
or U4779 (N_4779,N_3354,N_3315);
or U4780 (N_4780,N_3522,N_3883);
nand U4781 (N_4781,N_3119,N_3860);
nor U4782 (N_4782,N_3142,N_3542);
nor U4783 (N_4783,N_3519,N_3410);
or U4784 (N_4784,N_3376,N_3771);
or U4785 (N_4785,N_3311,N_3613);
or U4786 (N_4786,N_3329,N_3576);
or U4787 (N_4787,N_3960,N_3663);
nor U4788 (N_4788,N_3838,N_3760);
and U4789 (N_4789,N_3475,N_3638);
nand U4790 (N_4790,N_3725,N_3398);
or U4791 (N_4791,N_3942,N_3460);
and U4792 (N_4792,N_3657,N_3379);
and U4793 (N_4793,N_3092,N_3369);
and U4794 (N_4794,N_3005,N_3309);
or U4795 (N_4795,N_3093,N_3668);
nor U4796 (N_4796,N_3583,N_3813);
nor U4797 (N_4797,N_3597,N_3663);
nand U4798 (N_4798,N_3075,N_3491);
nand U4799 (N_4799,N_3777,N_3572);
or U4800 (N_4800,N_3212,N_3062);
or U4801 (N_4801,N_3416,N_3990);
nand U4802 (N_4802,N_3146,N_3842);
or U4803 (N_4803,N_3723,N_3597);
or U4804 (N_4804,N_3923,N_3424);
xnor U4805 (N_4805,N_3473,N_3882);
or U4806 (N_4806,N_3561,N_3308);
nor U4807 (N_4807,N_3702,N_3155);
and U4808 (N_4808,N_3451,N_3401);
and U4809 (N_4809,N_3718,N_3634);
nand U4810 (N_4810,N_3144,N_3718);
and U4811 (N_4811,N_3052,N_3965);
nand U4812 (N_4812,N_3384,N_3776);
or U4813 (N_4813,N_3312,N_3298);
or U4814 (N_4814,N_3558,N_3702);
nand U4815 (N_4815,N_3563,N_3416);
and U4816 (N_4816,N_3131,N_3412);
nor U4817 (N_4817,N_3194,N_3650);
nor U4818 (N_4818,N_3340,N_3797);
or U4819 (N_4819,N_3796,N_3440);
nor U4820 (N_4820,N_3683,N_3911);
nand U4821 (N_4821,N_3346,N_3500);
nand U4822 (N_4822,N_3777,N_3862);
and U4823 (N_4823,N_3566,N_3525);
and U4824 (N_4824,N_3646,N_3559);
and U4825 (N_4825,N_3132,N_3391);
and U4826 (N_4826,N_3653,N_3508);
nand U4827 (N_4827,N_3942,N_3814);
nand U4828 (N_4828,N_3647,N_3743);
or U4829 (N_4829,N_3408,N_3861);
nand U4830 (N_4830,N_3938,N_3894);
or U4831 (N_4831,N_3155,N_3341);
nand U4832 (N_4832,N_3875,N_3878);
and U4833 (N_4833,N_3354,N_3390);
nand U4834 (N_4834,N_3376,N_3514);
nor U4835 (N_4835,N_3963,N_3717);
nor U4836 (N_4836,N_3966,N_3180);
and U4837 (N_4837,N_3821,N_3521);
nand U4838 (N_4838,N_3477,N_3977);
and U4839 (N_4839,N_3511,N_3473);
nand U4840 (N_4840,N_3844,N_3291);
nand U4841 (N_4841,N_3740,N_3144);
or U4842 (N_4842,N_3941,N_3520);
nor U4843 (N_4843,N_3495,N_3972);
nand U4844 (N_4844,N_3672,N_3886);
nand U4845 (N_4845,N_3224,N_3675);
nand U4846 (N_4846,N_3118,N_3786);
and U4847 (N_4847,N_3086,N_3050);
or U4848 (N_4848,N_3653,N_3475);
and U4849 (N_4849,N_3162,N_3663);
nor U4850 (N_4850,N_3719,N_3239);
nand U4851 (N_4851,N_3640,N_3070);
and U4852 (N_4852,N_3752,N_3848);
nor U4853 (N_4853,N_3531,N_3726);
nand U4854 (N_4854,N_3148,N_3708);
nand U4855 (N_4855,N_3697,N_3828);
and U4856 (N_4856,N_3342,N_3360);
nor U4857 (N_4857,N_3109,N_3679);
or U4858 (N_4858,N_3793,N_3950);
nor U4859 (N_4859,N_3871,N_3304);
nor U4860 (N_4860,N_3792,N_3572);
nor U4861 (N_4861,N_3530,N_3925);
or U4862 (N_4862,N_3069,N_3787);
nand U4863 (N_4863,N_3203,N_3821);
and U4864 (N_4864,N_3156,N_3124);
nand U4865 (N_4865,N_3047,N_3575);
nand U4866 (N_4866,N_3687,N_3786);
nand U4867 (N_4867,N_3544,N_3123);
nor U4868 (N_4868,N_3672,N_3732);
nand U4869 (N_4869,N_3556,N_3990);
nor U4870 (N_4870,N_3785,N_3790);
nor U4871 (N_4871,N_3596,N_3203);
and U4872 (N_4872,N_3148,N_3426);
and U4873 (N_4873,N_3301,N_3812);
and U4874 (N_4874,N_3453,N_3274);
and U4875 (N_4875,N_3670,N_3154);
nor U4876 (N_4876,N_3817,N_3575);
and U4877 (N_4877,N_3673,N_3290);
or U4878 (N_4878,N_3553,N_3508);
nand U4879 (N_4879,N_3487,N_3878);
or U4880 (N_4880,N_3939,N_3949);
or U4881 (N_4881,N_3267,N_3580);
nor U4882 (N_4882,N_3393,N_3763);
or U4883 (N_4883,N_3609,N_3433);
and U4884 (N_4884,N_3284,N_3554);
nand U4885 (N_4885,N_3643,N_3254);
nand U4886 (N_4886,N_3222,N_3188);
or U4887 (N_4887,N_3799,N_3184);
nor U4888 (N_4888,N_3327,N_3322);
nor U4889 (N_4889,N_3289,N_3627);
or U4890 (N_4890,N_3492,N_3985);
or U4891 (N_4891,N_3678,N_3145);
nand U4892 (N_4892,N_3758,N_3438);
xor U4893 (N_4893,N_3340,N_3016);
xnor U4894 (N_4894,N_3768,N_3136);
nor U4895 (N_4895,N_3349,N_3578);
nand U4896 (N_4896,N_3398,N_3564);
nor U4897 (N_4897,N_3871,N_3555);
and U4898 (N_4898,N_3578,N_3516);
xnor U4899 (N_4899,N_3642,N_3626);
nor U4900 (N_4900,N_3192,N_3162);
nor U4901 (N_4901,N_3396,N_3347);
nand U4902 (N_4902,N_3765,N_3941);
or U4903 (N_4903,N_3443,N_3793);
or U4904 (N_4904,N_3429,N_3539);
nor U4905 (N_4905,N_3287,N_3509);
or U4906 (N_4906,N_3532,N_3799);
xor U4907 (N_4907,N_3316,N_3646);
or U4908 (N_4908,N_3165,N_3660);
nand U4909 (N_4909,N_3859,N_3170);
nor U4910 (N_4910,N_3295,N_3027);
nand U4911 (N_4911,N_3665,N_3139);
and U4912 (N_4912,N_3514,N_3048);
nor U4913 (N_4913,N_3742,N_3995);
nand U4914 (N_4914,N_3987,N_3298);
or U4915 (N_4915,N_3583,N_3601);
or U4916 (N_4916,N_3934,N_3628);
nand U4917 (N_4917,N_3254,N_3761);
nand U4918 (N_4918,N_3453,N_3736);
nor U4919 (N_4919,N_3323,N_3120);
or U4920 (N_4920,N_3651,N_3282);
nor U4921 (N_4921,N_3085,N_3366);
or U4922 (N_4922,N_3299,N_3455);
and U4923 (N_4923,N_3175,N_3987);
and U4924 (N_4924,N_3743,N_3376);
nor U4925 (N_4925,N_3959,N_3888);
or U4926 (N_4926,N_3002,N_3862);
nand U4927 (N_4927,N_3498,N_3407);
nand U4928 (N_4928,N_3601,N_3501);
or U4929 (N_4929,N_3173,N_3659);
and U4930 (N_4930,N_3042,N_3109);
and U4931 (N_4931,N_3282,N_3343);
and U4932 (N_4932,N_3751,N_3437);
and U4933 (N_4933,N_3149,N_3591);
nor U4934 (N_4934,N_3406,N_3090);
and U4935 (N_4935,N_3576,N_3719);
and U4936 (N_4936,N_3386,N_3860);
nand U4937 (N_4937,N_3885,N_3822);
or U4938 (N_4938,N_3331,N_3217);
or U4939 (N_4939,N_3855,N_3675);
or U4940 (N_4940,N_3885,N_3534);
and U4941 (N_4941,N_3815,N_3499);
and U4942 (N_4942,N_3022,N_3657);
nor U4943 (N_4943,N_3273,N_3705);
nor U4944 (N_4944,N_3847,N_3901);
or U4945 (N_4945,N_3035,N_3392);
nor U4946 (N_4946,N_3782,N_3213);
nor U4947 (N_4947,N_3129,N_3746);
nand U4948 (N_4948,N_3129,N_3001);
and U4949 (N_4949,N_3150,N_3140);
nand U4950 (N_4950,N_3757,N_3644);
nor U4951 (N_4951,N_3515,N_3520);
or U4952 (N_4952,N_3817,N_3632);
nor U4953 (N_4953,N_3142,N_3445);
or U4954 (N_4954,N_3477,N_3808);
and U4955 (N_4955,N_3468,N_3183);
nand U4956 (N_4956,N_3350,N_3920);
and U4957 (N_4957,N_3342,N_3737);
nand U4958 (N_4958,N_3155,N_3752);
nand U4959 (N_4959,N_3928,N_3340);
nand U4960 (N_4960,N_3345,N_3403);
or U4961 (N_4961,N_3582,N_3306);
nor U4962 (N_4962,N_3409,N_3948);
or U4963 (N_4963,N_3094,N_3905);
and U4964 (N_4964,N_3662,N_3232);
or U4965 (N_4965,N_3824,N_3270);
nor U4966 (N_4966,N_3339,N_3373);
and U4967 (N_4967,N_3607,N_3770);
nand U4968 (N_4968,N_3787,N_3865);
nor U4969 (N_4969,N_3597,N_3424);
nand U4970 (N_4970,N_3324,N_3728);
nand U4971 (N_4971,N_3697,N_3485);
or U4972 (N_4972,N_3931,N_3367);
nand U4973 (N_4973,N_3977,N_3741);
or U4974 (N_4974,N_3099,N_3923);
nand U4975 (N_4975,N_3884,N_3216);
or U4976 (N_4976,N_3042,N_3617);
or U4977 (N_4977,N_3470,N_3752);
or U4978 (N_4978,N_3462,N_3155);
or U4979 (N_4979,N_3956,N_3119);
nor U4980 (N_4980,N_3555,N_3176);
or U4981 (N_4981,N_3122,N_3031);
nand U4982 (N_4982,N_3053,N_3267);
nor U4983 (N_4983,N_3690,N_3736);
nor U4984 (N_4984,N_3925,N_3364);
nand U4985 (N_4985,N_3943,N_3186);
or U4986 (N_4986,N_3212,N_3769);
nand U4987 (N_4987,N_3486,N_3104);
or U4988 (N_4988,N_3496,N_3168);
nand U4989 (N_4989,N_3546,N_3049);
nor U4990 (N_4990,N_3563,N_3182);
and U4991 (N_4991,N_3915,N_3133);
nor U4992 (N_4992,N_3144,N_3457);
and U4993 (N_4993,N_3952,N_3022);
and U4994 (N_4994,N_3831,N_3693);
nand U4995 (N_4995,N_3086,N_3331);
nor U4996 (N_4996,N_3151,N_3196);
nor U4997 (N_4997,N_3357,N_3207);
nor U4998 (N_4998,N_3367,N_3803);
or U4999 (N_4999,N_3335,N_3722);
or UO_0 (O_0,N_4901,N_4253);
nand UO_1 (O_1,N_4468,N_4850);
or UO_2 (O_2,N_4416,N_4554);
or UO_3 (O_3,N_4923,N_4004);
nand UO_4 (O_4,N_4002,N_4685);
nand UO_5 (O_5,N_4789,N_4121);
nand UO_6 (O_6,N_4433,N_4087);
nor UO_7 (O_7,N_4930,N_4039);
nand UO_8 (O_8,N_4546,N_4318);
nand UO_9 (O_9,N_4677,N_4198);
and UO_10 (O_10,N_4085,N_4952);
and UO_11 (O_11,N_4893,N_4719);
nand UO_12 (O_12,N_4831,N_4907);
and UO_13 (O_13,N_4038,N_4337);
and UO_14 (O_14,N_4683,N_4608);
or UO_15 (O_15,N_4784,N_4163);
or UO_16 (O_16,N_4955,N_4650);
nor UO_17 (O_17,N_4679,N_4682);
or UO_18 (O_18,N_4880,N_4017);
or UO_19 (O_19,N_4667,N_4480);
nand UO_20 (O_20,N_4265,N_4585);
or UO_21 (O_21,N_4094,N_4985);
nor UO_22 (O_22,N_4963,N_4582);
or UO_23 (O_23,N_4579,N_4353);
and UO_24 (O_24,N_4828,N_4453);
nor UO_25 (O_25,N_4603,N_4047);
nor UO_26 (O_26,N_4500,N_4083);
or UO_27 (O_27,N_4390,N_4474);
nor UO_28 (O_28,N_4544,N_4309);
nor UO_29 (O_29,N_4890,N_4242);
xnor UO_30 (O_30,N_4736,N_4120);
nand UO_31 (O_31,N_4153,N_4558);
and UO_32 (O_32,N_4926,N_4568);
nand UO_33 (O_33,N_4729,N_4670);
or UO_34 (O_34,N_4959,N_4666);
nand UO_35 (O_35,N_4056,N_4340);
and UO_36 (O_36,N_4680,N_4644);
nand UO_37 (O_37,N_4200,N_4075);
nand UO_38 (O_38,N_4999,N_4082);
or UO_39 (O_39,N_4132,N_4431);
xnor UO_40 (O_40,N_4587,N_4933);
or UO_41 (O_41,N_4442,N_4669);
or UO_42 (O_42,N_4098,N_4825);
nand UO_43 (O_43,N_4781,N_4502);
and UO_44 (O_44,N_4172,N_4965);
and UO_45 (O_45,N_4145,N_4175);
and UO_46 (O_46,N_4570,N_4146);
nand UO_47 (O_47,N_4526,N_4355);
or UO_48 (O_48,N_4642,N_4627);
nand UO_49 (O_49,N_4203,N_4081);
nor UO_50 (O_50,N_4223,N_4402);
and UO_51 (O_51,N_4845,N_4698);
nand UO_52 (O_52,N_4283,N_4209);
nor UO_53 (O_53,N_4754,N_4798);
or UO_54 (O_54,N_4564,N_4055);
nor UO_55 (O_55,N_4884,N_4492);
or UO_56 (O_56,N_4243,N_4815);
nand UO_57 (O_57,N_4584,N_4881);
and UO_58 (O_58,N_4425,N_4036);
and UO_59 (O_59,N_4906,N_4541);
nand UO_60 (O_60,N_4673,N_4366);
nor UO_61 (O_61,N_4197,N_4462);
nor UO_62 (O_62,N_4556,N_4772);
and UO_63 (O_63,N_4134,N_4841);
nand UO_64 (O_64,N_4177,N_4596);
nor UO_65 (O_65,N_4836,N_4046);
and UO_66 (O_66,N_4505,N_4634);
and UO_67 (O_67,N_4256,N_4135);
and UO_68 (O_68,N_4948,N_4446);
or UO_69 (O_69,N_4523,N_4941);
nand UO_70 (O_70,N_4591,N_4728);
nand UO_71 (O_71,N_4843,N_4624);
nand UO_72 (O_72,N_4614,N_4143);
or UO_73 (O_73,N_4237,N_4710);
or UO_74 (O_74,N_4069,N_4879);
nor UO_75 (O_75,N_4856,N_4967);
or UO_76 (O_76,N_4645,N_4263);
nor UO_77 (O_77,N_4195,N_4535);
or UO_78 (O_78,N_4168,N_4116);
nand UO_79 (O_79,N_4551,N_4336);
nand UO_80 (O_80,N_4092,N_4285);
and UO_81 (O_81,N_4621,N_4643);
nor UO_82 (O_82,N_4583,N_4981);
or UO_83 (O_83,N_4138,N_4616);
or UO_84 (O_84,N_4157,N_4571);
and UO_85 (O_85,N_4284,N_4771);
and UO_86 (O_86,N_4148,N_4575);
and UO_87 (O_87,N_4574,N_4545);
or UO_88 (O_88,N_4061,N_4258);
nor UO_89 (O_89,N_4808,N_4550);
nor UO_90 (O_90,N_4324,N_4747);
nor UO_91 (O_91,N_4688,N_4302);
nor UO_92 (O_92,N_4974,N_4954);
or UO_93 (O_93,N_4973,N_4569);
nand UO_94 (O_94,N_4025,N_4744);
and UO_95 (O_95,N_4033,N_4429);
and UO_96 (O_96,N_4975,N_4498);
nand UO_97 (O_97,N_4597,N_4212);
nor UO_98 (O_98,N_4900,N_4162);
nand UO_99 (O_99,N_4012,N_4876);
and UO_100 (O_100,N_4536,N_4045);
nand UO_101 (O_101,N_4916,N_4408);
nor UO_102 (O_102,N_4457,N_4581);
nand UO_103 (O_103,N_4181,N_4411);
or UO_104 (O_104,N_4658,N_4717);
nor UO_105 (O_105,N_4185,N_4914);
and UO_106 (O_106,N_4222,N_4803);
or UO_107 (O_107,N_4530,N_4042);
or UO_108 (O_108,N_4481,N_4851);
nor UO_109 (O_109,N_4205,N_4601);
or UO_110 (O_110,N_4816,N_4488);
nor UO_111 (O_111,N_4588,N_4282);
or UO_112 (O_112,N_4348,N_4170);
nor UO_113 (O_113,N_4657,N_4295);
nor UO_114 (O_114,N_4228,N_4761);
and UO_115 (O_115,N_4837,N_4493);
and UO_116 (O_116,N_4130,N_4418);
and UO_117 (O_117,N_4296,N_4066);
and UO_118 (O_118,N_4128,N_4067);
or UO_119 (O_119,N_4547,N_4393);
or UO_120 (O_120,N_4133,N_4427);
xnor UO_121 (O_121,N_4533,N_4392);
or UO_122 (O_122,N_4245,N_4857);
and UO_123 (O_123,N_4312,N_4793);
nor UO_124 (O_124,N_4982,N_4199);
nand UO_125 (O_125,N_4054,N_4885);
or UO_126 (O_126,N_4173,N_4626);
nor UO_127 (O_127,N_4593,N_4994);
nand UO_128 (O_128,N_4641,N_4272);
nand UO_129 (O_129,N_4794,N_4276);
nand UO_130 (O_130,N_4678,N_4328);
and UO_131 (O_131,N_4635,N_4639);
nor UO_132 (O_132,N_4555,N_4167);
and UO_133 (O_133,N_4219,N_4630);
nand UO_134 (O_134,N_4008,N_4315);
and UO_135 (O_135,N_4439,N_4354);
or UO_136 (O_136,N_4022,N_4158);
or UO_137 (O_137,N_4735,N_4229);
and UO_138 (O_138,N_4358,N_4232);
and UO_139 (O_139,N_4420,N_4962);
or UO_140 (O_140,N_4730,N_4227);
nor UO_141 (O_141,N_4592,N_4178);
or UO_142 (O_142,N_4712,N_4938);
nor UO_143 (O_143,N_4001,N_4549);
nand UO_144 (O_144,N_4449,N_4407);
or UO_145 (O_145,N_4822,N_4918);
and UO_146 (O_146,N_4578,N_4006);
nor UO_147 (O_147,N_4726,N_4868);
nor UO_148 (O_148,N_4434,N_4921);
or UO_149 (O_149,N_4887,N_4510);
nand UO_150 (O_150,N_4651,N_4628);
nand UO_151 (O_151,N_4159,N_4350);
and UO_152 (O_152,N_4920,N_4319);
nand UO_153 (O_153,N_4041,N_4059);
nor UO_154 (O_154,N_4231,N_4720);
nor UO_155 (O_155,N_4882,N_4049);
nand UO_156 (O_156,N_4703,N_4196);
and UO_157 (O_157,N_4909,N_4910);
nand UO_158 (O_158,N_4637,N_4649);
nand UO_159 (O_159,N_4180,N_4383);
nand UO_160 (O_160,N_4987,N_4619);
nand UO_161 (O_161,N_4088,N_4942);
nand UO_162 (O_162,N_4104,N_4823);
nand UO_163 (O_163,N_4971,N_4925);
and UO_164 (O_164,N_4102,N_4765);
or UO_165 (O_165,N_4939,N_4397);
nand UO_166 (O_166,N_4832,N_4208);
nand UO_167 (O_167,N_4552,N_4469);
nor UO_168 (O_168,N_4991,N_4993);
or UO_169 (O_169,N_4424,N_4345);
nand UO_170 (O_170,N_4528,N_4950);
and UO_171 (O_171,N_4370,N_4154);
and UO_172 (O_172,N_4463,N_4264);
and UO_173 (O_173,N_4838,N_4112);
or UO_174 (O_174,N_4452,N_4812);
nand UO_175 (O_175,N_4940,N_4511);
or UO_176 (O_176,N_4929,N_4040);
nor UO_177 (O_177,N_4902,N_4438);
nor UO_178 (O_178,N_4935,N_4271);
nand UO_179 (O_179,N_4847,N_4905);
or UO_180 (O_180,N_4129,N_4848);
or UO_181 (O_181,N_4292,N_4738);
nor UO_182 (O_182,N_4386,N_4648);
and UO_183 (O_183,N_4335,N_4969);
or UO_184 (O_184,N_4301,N_4103);
nand UO_185 (O_185,N_4951,N_4695);
nand UO_186 (O_186,N_4853,N_4410);
nand UO_187 (O_187,N_4202,N_4734);
nand UO_188 (O_188,N_4437,N_4108);
and UO_189 (O_189,N_4525,N_4136);
or UO_190 (O_190,N_4507,N_4251);
or UO_191 (O_191,N_4762,N_4293);
nand UO_192 (O_192,N_4382,N_4477);
nand UO_193 (O_193,N_4321,N_4756);
or UO_194 (O_194,N_4891,N_4646);
nor UO_195 (O_195,N_4101,N_4702);
or UO_196 (O_196,N_4466,N_4269);
and UO_197 (O_197,N_4990,N_4095);
nand UO_198 (O_198,N_4846,N_4152);
nor UO_199 (O_199,N_4927,N_4931);
or UO_200 (O_200,N_4028,N_4026);
or UO_201 (O_201,N_4998,N_4977);
or UO_202 (O_202,N_4412,N_4191);
nand UO_203 (O_203,N_4788,N_4300);
nand UO_204 (O_204,N_4878,N_4560);
nor UO_205 (O_205,N_4694,N_4709);
or UO_206 (O_206,N_4377,N_4903);
nand UO_207 (O_207,N_4010,N_4553);
and UO_208 (O_208,N_4946,N_4707);
and UO_209 (O_209,N_4811,N_4141);
or UO_210 (O_210,N_4704,N_4790);
or UO_211 (O_211,N_4338,N_4052);
and UO_212 (O_212,N_4773,N_4883);
or UO_213 (O_213,N_4749,N_4044);
nor UO_214 (O_214,N_4668,N_4443);
or UO_215 (O_215,N_4557,N_4326);
nand UO_216 (O_216,N_4655,N_4661);
nor UO_217 (O_217,N_4415,N_4516);
nor UO_218 (O_218,N_4599,N_4467);
and UO_219 (O_219,N_4612,N_4629);
and UO_220 (O_220,N_4509,N_4632);
or UO_221 (O_221,N_4915,N_4323);
or UO_222 (O_222,N_4779,N_4996);
nand UO_223 (O_223,N_4334,N_4904);
or UO_224 (O_224,N_4381,N_4691);
nand UO_225 (O_225,N_4249,N_4186);
or UO_226 (O_226,N_4015,N_4344);
xnor UO_227 (O_227,N_4675,N_4016);
and UO_228 (O_228,N_4423,N_4944);
nand UO_229 (O_229,N_4123,N_4144);
or UO_230 (O_230,N_4299,N_4693);
or UO_231 (O_231,N_4527,N_4078);
or UO_232 (O_232,N_4428,N_4294);
or UO_233 (O_233,N_4259,N_4214);
nor UO_234 (O_234,N_4986,N_4960);
or UO_235 (O_235,N_4869,N_4610);
or UO_236 (O_236,N_4586,N_4086);
nor UO_237 (O_237,N_4739,N_4031);
or UO_238 (O_238,N_4471,N_4757);
and UO_239 (O_239,N_4606,N_4470);
nor UO_240 (O_240,N_4540,N_4341);
nor UO_241 (O_241,N_4817,N_4529);
nor UO_242 (O_242,N_4864,N_4697);
nor UO_243 (O_243,N_4576,N_4769);
and UO_244 (O_244,N_4852,N_4659);
or UO_245 (O_245,N_4156,N_4786);
nand UO_246 (O_246,N_4791,N_4385);
or UO_247 (O_247,N_4947,N_4182);
nor UO_248 (O_248,N_4352,N_4722);
or UO_249 (O_249,N_4089,N_4833);
nand UO_250 (O_250,N_4745,N_4215);
and UO_251 (O_251,N_4705,N_4567);
nor UO_252 (O_252,N_4631,N_4958);
and UO_253 (O_253,N_4013,N_4161);
or UO_254 (O_254,N_4403,N_4618);
nand UO_255 (O_255,N_4113,N_4444);
and UO_256 (O_256,N_4356,N_4164);
nor UO_257 (O_257,N_4989,N_4458);
and UO_258 (O_258,N_4594,N_4287);
nor UO_259 (O_259,N_4924,N_4665);
and UO_260 (O_260,N_4819,N_4638);
and UO_261 (O_261,N_4672,N_4401);
nand UO_262 (O_262,N_4363,N_4043);
or UO_263 (O_263,N_4539,N_4122);
or UO_264 (O_264,N_4517,N_4814);
or UO_265 (O_265,N_4494,N_4640);
nand UO_266 (O_266,N_4778,N_4413);
nor UO_267 (O_267,N_4241,N_4740);
nand UO_268 (O_268,N_4306,N_4257);
nor UO_269 (O_269,N_4389,N_4867);
or UO_270 (O_270,N_4252,N_4080);
or UO_271 (O_271,N_4827,N_4325);
and UO_272 (O_272,N_4834,N_4731);
nor UO_273 (O_273,N_4213,N_4071);
and UO_274 (O_274,N_4548,N_4187);
nand UO_275 (O_275,N_4795,N_4005);
or UO_276 (O_276,N_4074,N_4274);
nand UO_277 (O_277,N_4713,N_4034);
and UO_278 (O_278,N_4065,N_4331);
or UO_279 (O_279,N_4479,N_4782);
and UO_280 (O_280,N_4435,N_4524);
and UO_281 (O_281,N_4270,N_4978);
nor UO_282 (O_282,N_4204,N_4297);
and UO_283 (O_283,N_4368,N_4715);
nand UO_284 (O_284,N_4035,N_4096);
or UO_285 (O_285,N_4800,N_4422);
and UO_286 (O_286,N_4131,N_4866);
nor UO_287 (O_287,N_4051,N_4486);
or UO_288 (O_288,N_4030,N_4805);
or UO_289 (O_289,N_4724,N_4733);
nor UO_290 (O_290,N_4399,N_4937);
nand UO_291 (O_291,N_4796,N_4362);
nor UO_292 (O_292,N_4000,N_4378);
and UO_293 (O_293,N_4854,N_4647);
xor UO_294 (O_294,N_4023,N_4077);
or UO_295 (O_295,N_4426,N_4577);
or UO_296 (O_296,N_4084,N_4911);
nor UO_297 (O_297,N_4858,N_4859);
nand UO_298 (O_298,N_4995,N_4741);
nor UO_299 (O_299,N_4254,N_4820);
or UO_300 (O_300,N_4060,N_4922);
nand UO_301 (O_301,N_4750,N_4174);
nand UO_302 (O_302,N_4860,N_4919);
nor UO_303 (O_303,N_4322,N_4980);
or UO_304 (O_304,N_4472,N_4656);
and UO_305 (O_305,N_4037,N_4559);
nand UO_306 (O_306,N_4830,N_4395);
and UO_307 (O_307,N_4091,N_4842);
and UO_308 (O_308,N_4244,N_4275);
and UO_309 (O_309,N_4755,N_4976);
or UO_310 (O_310,N_4380,N_4127);
and UO_311 (O_311,N_4785,N_4260);
or UO_312 (O_312,N_4291,N_4775);
nand UO_313 (O_313,N_4388,N_4844);
nor UO_314 (O_314,N_4417,N_4217);
and UO_315 (O_315,N_4347,N_4364);
and UO_316 (O_316,N_4763,N_4166);
nand UO_317 (O_317,N_4063,N_4376);
nand UO_318 (O_318,N_4273,N_4687);
nor UO_319 (O_319,N_4753,N_4288);
nand UO_320 (O_320,N_4405,N_4818);
or UO_321 (O_321,N_4870,N_4058);
nand UO_322 (O_322,N_4032,N_4476);
and UO_323 (O_323,N_4313,N_4169);
nor UO_324 (O_324,N_4473,N_4414);
and UO_325 (O_325,N_4506,N_4877);
and UO_326 (O_326,N_4111,N_4752);
or UO_327 (O_327,N_4686,N_4070);
nor UO_328 (O_328,N_4460,N_4316);
xor UO_329 (O_329,N_4807,N_4100);
nor UO_330 (O_330,N_4743,N_4676);
nor UO_331 (O_331,N_4357,N_4792);
nand UO_332 (O_332,N_4371,N_4247);
or UO_333 (O_333,N_4124,N_4183);
nand UO_334 (O_334,N_4454,N_4018);
or UO_335 (O_335,N_4150,N_4660);
or UO_336 (O_336,N_4620,N_4718);
nand UO_337 (O_337,N_4235,N_4305);
nand UO_338 (O_338,N_4409,N_4598);
nor UO_339 (O_339,N_4727,N_4019);
or UO_340 (O_340,N_4671,N_4165);
or UO_341 (O_341,N_4992,N_4447);
and UO_342 (O_342,N_4107,N_4824);
and UO_343 (O_343,N_4501,N_4106);
nor UO_344 (O_344,N_4320,N_4532);
and UO_345 (O_345,N_4908,N_4459);
nor UO_346 (O_346,N_4953,N_4117);
or UO_347 (O_347,N_4406,N_4465);
or UO_348 (O_348,N_4611,N_4068);
nand UO_349 (O_349,N_4062,N_4384);
nand UO_350 (O_350,N_4455,N_4543);
and UO_351 (O_351,N_4806,N_4277);
or UO_352 (O_352,N_4684,N_4663);
nand UO_353 (O_353,N_4490,N_4246);
nand UO_354 (O_354,N_4396,N_4562);
nand UO_355 (O_355,N_4192,N_4311);
nand UO_356 (O_356,N_4988,N_4072);
and UO_357 (O_357,N_4307,N_4607);
or UO_358 (O_358,N_4531,N_4280);
or UO_359 (O_359,N_4934,N_4139);
and UO_360 (O_360,N_4268,N_4983);
nor UO_361 (O_361,N_4303,N_4142);
nor UO_362 (O_362,N_4286,N_4190);
or UO_363 (O_363,N_4027,N_4105);
nand UO_364 (O_364,N_4349,N_4020);
or UO_365 (O_365,N_4625,N_4188);
or UO_366 (O_366,N_4097,N_4888);
nor UO_367 (O_367,N_4330,N_4398);
or UO_368 (O_368,N_4029,N_4699);
and UO_369 (O_369,N_4700,N_4495);
nor UO_370 (O_370,N_4861,N_4343);
and UO_371 (O_371,N_4821,N_4839);
nor UO_372 (O_372,N_4372,N_4513);
nand UO_373 (O_373,N_4367,N_4871);
and UO_374 (O_374,N_4895,N_4964);
and UO_375 (O_375,N_4913,N_4966);
nor UO_376 (O_376,N_4419,N_4211);
nor UO_377 (O_377,N_4829,N_4563);
nor UO_378 (O_378,N_4514,N_4768);
and UO_379 (O_379,N_4184,N_4011);
nor UO_380 (O_380,N_4725,N_4746);
nor UO_381 (O_381,N_4342,N_4826);
or UO_382 (O_382,N_4478,N_4748);
nand UO_383 (O_383,N_4742,N_4248);
nand UO_384 (O_384,N_4580,N_4804);
nand UO_385 (O_385,N_4233,N_4430);
nand UO_386 (O_386,N_4622,N_4968);
or UO_387 (O_387,N_4674,N_4898);
or UO_388 (O_388,N_4767,N_4053);
and UO_389 (O_389,N_4118,N_4099);
nand UO_390 (O_390,N_4957,N_4445);
nor UO_391 (O_391,N_4997,N_4956);
nand UO_392 (O_392,N_4194,N_4003);
or UO_393 (O_393,N_4522,N_4889);
nand UO_394 (O_394,N_4064,N_4290);
nand UO_395 (O_395,N_4373,N_4394);
nor UO_396 (O_396,N_4664,N_4737);
nand UO_397 (O_397,N_4160,N_4654);
or UO_398 (O_398,N_4261,N_4538);
nor UO_399 (O_399,N_4432,N_4281);
xor UO_400 (O_400,N_4810,N_4266);
or UO_401 (O_401,N_4007,N_4125);
and UO_402 (O_402,N_4332,N_4573);
nor UO_403 (O_403,N_4126,N_4706);
or UO_404 (O_404,N_4482,N_4696);
nor UO_405 (O_405,N_4333,N_4456);
xnor UO_406 (O_406,N_4137,N_4801);
nand UO_407 (O_407,N_4783,N_4797);
xnor UO_408 (O_408,N_4809,N_4542);
nor UO_409 (O_409,N_4210,N_4110);
nand UO_410 (O_410,N_4840,N_4970);
nor UO_411 (O_411,N_4267,N_4206);
and UO_412 (O_412,N_4484,N_4021);
nand UO_413 (O_413,N_4503,N_4572);
and UO_414 (O_414,N_4387,N_4984);
nor UO_415 (O_415,N_4421,N_4865);
nand UO_416 (O_416,N_4653,N_4932);
nand UO_417 (O_417,N_4714,N_4774);
nor UO_418 (O_418,N_4379,N_4849);
and UO_419 (O_419,N_4339,N_4359);
and UO_420 (O_420,N_4140,N_4949);
nand UO_421 (O_421,N_4894,N_4298);
or UO_422 (O_422,N_4566,N_4873);
nor UO_423 (O_423,N_4220,N_4076);
or UO_424 (O_424,N_4681,N_4262);
and UO_425 (O_425,N_4936,N_4499);
and UO_426 (O_426,N_4109,N_4400);
nand UO_427 (O_427,N_4777,N_4689);
and UO_428 (O_428,N_4226,N_4436);
or UO_429 (O_429,N_4732,N_4609);
nor UO_430 (O_430,N_4723,N_4604);
nor UO_431 (O_431,N_4216,N_4751);
and UO_432 (O_432,N_4050,N_4304);
and UO_433 (O_433,N_4721,N_4014);
and UO_434 (O_434,N_4308,N_4279);
or UO_435 (O_435,N_4862,N_4602);
nor UO_436 (O_436,N_4928,N_4508);
nor UO_437 (O_437,N_4515,N_4489);
nor UO_438 (O_438,N_4079,N_4440);
or UO_439 (O_439,N_4369,N_4238);
nor UO_440 (O_440,N_4692,N_4605);
and UO_441 (O_441,N_4617,N_4149);
or UO_442 (O_442,N_4491,N_4497);
nor UO_443 (O_443,N_4221,N_4147);
nor UO_444 (O_444,N_4764,N_4759);
and UO_445 (O_445,N_4314,N_4813);
nand UO_446 (O_446,N_4207,N_4613);
and UO_447 (O_447,N_4835,N_4519);
or UO_448 (O_448,N_4863,N_4701);
and UO_449 (O_449,N_4652,N_4289);
nand UO_450 (O_450,N_4201,N_4776);
and UO_451 (O_451,N_4057,N_4441);
and UO_452 (O_452,N_4375,N_4636);
nor UO_453 (O_453,N_4475,N_4329);
and UO_454 (O_454,N_4189,N_4899);
nor UO_455 (O_455,N_4615,N_4346);
and UO_456 (O_456,N_4151,N_4912);
nand UO_457 (O_457,N_4521,N_4708);
and UO_458 (O_458,N_4799,N_4448);
nor UO_459 (O_459,N_4802,N_4896);
nor UO_460 (O_460,N_4875,N_4351);
and UO_461 (O_461,N_4114,N_4787);
nor UO_462 (O_462,N_4633,N_4716);
nand UO_463 (O_463,N_4115,N_4917);
or UO_464 (O_464,N_4230,N_4758);
nand UO_465 (O_465,N_4193,N_4770);
nand UO_466 (O_466,N_4520,N_4374);
and UO_467 (O_467,N_4589,N_4317);
and UO_468 (O_468,N_4662,N_4690);
nor UO_469 (O_469,N_4225,N_4483);
nand UO_470 (O_470,N_4537,N_4090);
nor UO_471 (O_471,N_4361,N_4365);
nor UO_472 (O_472,N_4278,N_4234);
or UO_473 (O_473,N_4600,N_4961);
or UO_474 (O_474,N_4024,N_4464);
and UO_475 (O_475,N_4512,N_4485);
or UO_476 (O_476,N_4874,N_4250);
nand UO_477 (O_477,N_4872,N_4760);
nor UO_478 (O_478,N_4240,N_4766);
nand UO_479 (O_479,N_4073,N_4236);
nor UO_480 (O_480,N_4119,N_4534);
nor UO_481 (O_481,N_4239,N_4048);
or UO_482 (O_482,N_4224,N_4179);
nor UO_483 (O_483,N_4451,N_4487);
and UO_484 (O_484,N_4310,N_4780);
nor UO_485 (O_485,N_4979,N_4155);
nor UO_486 (O_486,N_4623,N_4972);
nand UO_487 (O_487,N_4504,N_4496);
nand UO_488 (O_488,N_4461,N_4565);
and UO_489 (O_489,N_4711,N_4360);
and UO_490 (O_490,N_4218,N_4897);
nand UO_491 (O_491,N_4327,N_4391);
and UO_492 (O_492,N_4590,N_4886);
nand UO_493 (O_493,N_4255,N_4518);
nor UO_494 (O_494,N_4595,N_4450);
nor UO_495 (O_495,N_4009,N_4404);
and UO_496 (O_496,N_4561,N_4945);
or UO_497 (O_497,N_4855,N_4093);
and UO_498 (O_498,N_4176,N_4171);
nor UO_499 (O_499,N_4892,N_4943);
or UO_500 (O_500,N_4837,N_4094);
or UO_501 (O_501,N_4888,N_4783);
nand UO_502 (O_502,N_4689,N_4014);
and UO_503 (O_503,N_4787,N_4839);
nand UO_504 (O_504,N_4914,N_4765);
nand UO_505 (O_505,N_4700,N_4030);
nand UO_506 (O_506,N_4035,N_4680);
nor UO_507 (O_507,N_4322,N_4223);
nor UO_508 (O_508,N_4729,N_4612);
or UO_509 (O_509,N_4112,N_4321);
and UO_510 (O_510,N_4020,N_4885);
and UO_511 (O_511,N_4405,N_4286);
or UO_512 (O_512,N_4192,N_4469);
nand UO_513 (O_513,N_4761,N_4917);
and UO_514 (O_514,N_4193,N_4070);
or UO_515 (O_515,N_4872,N_4990);
or UO_516 (O_516,N_4035,N_4951);
and UO_517 (O_517,N_4665,N_4125);
or UO_518 (O_518,N_4811,N_4646);
or UO_519 (O_519,N_4041,N_4735);
nor UO_520 (O_520,N_4983,N_4903);
nor UO_521 (O_521,N_4707,N_4519);
or UO_522 (O_522,N_4291,N_4238);
or UO_523 (O_523,N_4819,N_4690);
nor UO_524 (O_524,N_4836,N_4394);
nor UO_525 (O_525,N_4124,N_4940);
nor UO_526 (O_526,N_4029,N_4017);
nor UO_527 (O_527,N_4317,N_4225);
nand UO_528 (O_528,N_4700,N_4254);
nor UO_529 (O_529,N_4352,N_4466);
and UO_530 (O_530,N_4762,N_4188);
and UO_531 (O_531,N_4662,N_4557);
or UO_532 (O_532,N_4120,N_4437);
nand UO_533 (O_533,N_4189,N_4563);
and UO_534 (O_534,N_4168,N_4744);
and UO_535 (O_535,N_4376,N_4716);
nor UO_536 (O_536,N_4256,N_4604);
or UO_537 (O_537,N_4859,N_4098);
nand UO_538 (O_538,N_4657,N_4146);
nand UO_539 (O_539,N_4282,N_4781);
nand UO_540 (O_540,N_4046,N_4736);
nor UO_541 (O_541,N_4310,N_4904);
or UO_542 (O_542,N_4880,N_4252);
or UO_543 (O_543,N_4996,N_4134);
or UO_544 (O_544,N_4879,N_4591);
or UO_545 (O_545,N_4360,N_4469);
or UO_546 (O_546,N_4609,N_4581);
and UO_547 (O_547,N_4794,N_4397);
nor UO_548 (O_548,N_4767,N_4360);
nand UO_549 (O_549,N_4628,N_4639);
nor UO_550 (O_550,N_4375,N_4213);
or UO_551 (O_551,N_4978,N_4190);
and UO_552 (O_552,N_4271,N_4229);
or UO_553 (O_553,N_4919,N_4925);
or UO_554 (O_554,N_4601,N_4618);
or UO_555 (O_555,N_4790,N_4230);
and UO_556 (O_556,N_4400,N_4087);
and UO_557 (O_557,N_4397,N_4523);
nor UO_558 (O_558,N_4229,N_4759);
nand UO_559 (O_559,N_4891,N_4848);
nand UO_560 (O_560,N_4983,N_4026);
and UO_561 (O_561,N_4300,N_4140);
or UO_562 (O_562,N_4656,N_4287);
or UO_563 (O_563,N_4812,N_4863);
nor UO_564 (O_564,N_4471,N_4225);
xor UO_565 (O_565,N_4866,N_4659);
and UO_566 (O_566,N_4264,N_4053);
and UO_567 (O_567,N_4547,N_4227);
and UO_568 (O_568,N_4701,N_4158);
nand UO_569 (O_569,N_4988,N_4480);
nor UO_570 (O_570,N_4318,N_4038);
and UO_571 (O_571,N_4717,N_4904);
and UO_572 (O_572,N_4100,N_4259);
and UO_573 (O_573,N_4429,N_4040);
nand UO_574 (O_574,N_4643,N_4898);
nor UO_575 (O_575,N_4484,N_4283);
or UO_576 (O_576,N_4999,N_4178);
and UO_577 (O_577,N_4445,N_4362);
or UO_578 (O_578,N_4125,N_4788);
nor UO_579 (O_579,N_4556,N_4815);
nor UO_580 (O_580,N_4841,N_4635);
xor UO_581 (O_581,N_4656,N_4038);
nand UO_582 (O_582,N_4460,N_4819);
nor UO_583 (O_583,N_4105,N_4950);
xor UO_584 (O_584,N_4055,N_4417);
or UO_585 (O_585,N_4309,N_4096);
nor UO_586 (O_586,N_4130,N_4789);
nand UO_587 (O_587,N_4873,N_4213);
and UO_588 (O_588,N_4012,N_4450);
nand UO_589 (O_589,N_4004,N_4725);
and UO_590 (O_590,N_4873,N_4906);
and UO_591 (O_591,N_4485,N_4308);
and UO_592 (O_592,N_4574,N_4523);
or UO_593 (O_593,N_4551,N_4357);
or UO_594 (O_594,N_4078,N_4514);
nand UO_595 (O_595,N_4122,N_4785);
nand UO_596 (O_596,N_4636,N_4411);
nand UO_597 (O_597,N_4678,N_4603);
and UO_598 (O_598,N_4294,N_4311);
or UO_599 (O_599,N_4589,N_4886);
nor UO_600 (O_600,N_4596,N_4793);
nor UO_601 (O_601,N_4804,N_4189);
nand UO_602 (O_602,N_4008,N_4535);
and UO_603 (O_603,N_4198,N_4657);
or UO_604 (O_604,N_4556,N_4303);
or UO_605 (O_605,N_4739,N_4446);
nand UO_606 (O_606,N_4012,N_4295);
or UO_607 (O_607,N_4705,N_4964);
or UO_608 (O_608,N_4505,N_4545);
nand UO_609 (O_609,N_4526,N_4015);
nand UO_610 (O_610,N_4519,N_4378);
nor UO_611 (O_611,N_4134,N_4256);
nand UO_612 (O_612,N_4962,N_4232);
or UO_613 (O_613,N_4481,N_4268);
nand UO_614 (O_614,N_4151,N_4439);
or UO_615 (O_615,N_4023,N_4106);
nor UO_616 (O_616,N_4700,N_4300);
and UO_617 (O_617,N_4117,N_4429);
nand UO_618 (O_618,N_4411,N_4650);
or UO_619 (O_619,N_4762,N_4919);
and UO_620 (O_620,N_4916,N_4522);
or UO_621 (O_621,N_4238,N_4865);
nand UO_622 (O_622,N_4416,N_4560);
xnor UO_623 (O_623,N_4277,N_4888);
and UO_624 (O_624,N_4233,N_4345);
and UO_625 (O_625,N_4520,N_4842);
and UO_626 (O_626,N_4721,N_4687);
nor UO_627 (O_627,N_4620,N_4223);
nor UO_628 (O_628,N_4364,N_4545);
nor UO_629 (O_629,N_4598,N_4905);
and UO_630 (O_630,N_4507,N_4740);
nand UO_631 (O_631,N_4404,N_4426);
or UO_632 (O_632,N_4565,N_4648);
nand UO_633 (O_633,N_4644,N_4868);
or UO_634 (O_634,N_4820,N_4904);
nand UO_635 (O_635,N_4031,N_4476);
nor UO_636 (O_636,N_4280,N_4632);
nand UO_637 (O_637,N_4856,N_4819);
xor UO_638 (O_638,N_4737,N_4459);
and UO_639 (O_639,N_4737,N_4821);
nand UO_640 (O_640,N_4977,N_4790);
or UO_641 (O_641,N_4094,N_4065);
nand UO_642 (O_642,N_4474,N_4654);
or UO_643 (O_643,N_4970,N_4555);
nor UO_644 (O_644,N_4659,N_4847);
and UO_645 (O_645,N_4905,N_4589);
and UO_646 (O_646,N_4589,N_4032);
and UO_647 (O_647,N_4091,N_4391);
nand UO_648 (O_648,N_4345,N_4639);
nand UO_649 (O_649,N_4650,N_4245);
nor UO_650 (O_650,N_4863,N_4371);
nor UO_651 (O_651,N_4731,N_4347);
or UO_652 (O_652,N_4571,N_4665);
nor UO_653 (O_653,N_4830,N_4238);
and UO_654 (O_654,N_4113,N_4958);
nor UO_655 (O_655,N_4239,N_4147);
nand UO_656 (O_656,N_4692,N_4997);
nand UO_657 (O_657,N_4554,N_4576);
and UO_658 (O_658,N_4438,N_4652);
nor UO_659 (O_659,N_4419,N_4193);
nor UO_660 (O_660,N_4952,N_4183);
and UO_661 (O_661,N_4617,N_4508);
nor UO_662 (O_662,N_4943,N_4460);
nand UO_663 (O_663,N_4230,N_4558);
or UO_664 (O_664,N_4158,N_4969);
or UO_665 (O_665,N_4158,N_4264);
nor UO_666 (O_666,N_4632,N_4462);
and UO_667 (O_667,N_4528,N_4817);
or UO_668 (O_668,N_4496,N_4298);
and UO_669 (O_669,N_4990,N_4720);
and UO_670 (O_670,N_4280,N_4532);
nor UO_671 (O_671,N_4365,N_4726);
nor UO_672 (O_672,N_4484,N_4834);
nor UO_673 (O_673,N_4729,N_4310);
nand UO_674 (O_674,N_4784,N_4919);
nor UO_675 (O_675,N_4914,N_4249);
xnor UO_676 (O_676,N_4234,N_4684);
nor UO_677 (O_677,N_4738,N_4010);
and UO_678 (O_678,N_4370,N_4354);
or UO_679 (O_679,N_4686,N_4805);
or UO_680 (O_680,N_4268,N_4546);
nand UO_681 (O_681,N_4347,N_4035);
and UO_682 (O_682,N_4880,N_4829);
or UO_683 (O_683,N_4038,N_4181);
or UO_684 (O_684,N_4558,N_4286);
nor UO_685 (O_685,N_4516,N_4098);
or UO_686 (O_686,N_4347,N_4820);
nand UO_687 (O_687,N_4696,N_4201);
or UO_688 (O_688,N_4399,N_4845);
nand UO_689 (O_689,N_4828,N_4999);
nor UO_690 (O_690,N_4347,N_4415);
or UO_691 (O_691,N_4614,N_4829);
or UO_692 (O_692,N_4812,N_4732);
nor UO_693 (O_693,N_4975,N_4473);
or UO_694 (O_694,N_4020,N_4067);
nor UO_695 (O_695,N_4132,N_4331);
nand UO_696 (O_696,N_4528,N_4273);
or UO_697 (O_697,N_4671,N_4186);
nand UO_698 (O_698,N_4521,N_4805);
nand UO_699 (O_699,N_4144,N_4884);
nor UO_700 (O_700,N_4942,N_4212);
and UO_701 (O_701,N_4101,N_4164);
nor UO_702 (O_702,N_4928,N_4155);
and UO_703 (O_703,N_4322,N_4825);
or UO_704 (O_704,N_4675,N_4543);
nor UO_705 (O_705,N_4694,N_4748);
and UO_706 (O_706,N_4509,N_4819);
or UO_707 (O_707,N_4379,N_4727);
or UO_708 (O_708,N_4797,N_4448);
nor UO_709 (O_709,N_4708,N_4742);
nor UO_710 (O_710,N_4863,N_4563);
nor UO_711 (O_711,N_4111,N_4428);
or UO_712 (O_712,N_4723,N_4443);
nor UO_713 (O_713,N_4229,N_4512);
nand UO_714 (O_714,N_4917,N_4076);
nor UO_715 (O_715,N_4253,N_4026);
and UO_716 (O_716,N_4983,N_4732);
nand UO_717 (O_717,N_4873,N_4020);
or UO_718 (O_718,N_4235,N_4619);
nor UO_719 (O_719,N_4440,N_4606);
nand UO_720 (O_720,N_4659,N_4235);
nand UO_721 (O_721,N_4559,N_4171);
nand UO_722 (O_722,N_4052,N_4237);
and UO_723 (O_723,N_4204,N_4026);
or UO_724 (O_724,N_4355,N_4111);
or UO_725 (O_725,N_4766,N_4219);
nand UO_726 (O_726,N_4090,N_4709);
or UO_727 (O_727,N_4283,N_4486);
nand UO_728 (O_728,N_4578,N_4506);
nor UO_729 (O_729,N_4115,N_4920);
or UO_730 (O_730,N_4437,N_4553);
nand UO_731 (O_731,N_4727,N_4396);
nor UO_732 (O_732,N_4427,N_4057);
and UO_733 (O_733,N_4274,N_4260);
nor UO_734 (O_734,N_4637,N_4297);
and UO_735 (O_735,N_4292,N_4604);
or UO_736 (O_736,N_4036,N_4070);
nor UO_737 (O_737,N_4381,N_4067);
or UO_738 (O_738,N_4215,N_4511);
or UO_739 (O_739,N_4991,N_4065);
and UO_740 (O_740,N_4984,N_4351);
and UO_741 (O_741,N_4227,N_4237);
nor UO_742 (O_742,N_4055,N_4204);
and UO_743 (O_743,N_4776,N_4740);
nor UO_744 (O_744,N_4333,N_4026);
nand UO_745 (O_745,N_4983,N_4547);
nand UO_746 (O_746,N_4428,N_4794);
and UO_747 (O_747,N_4878,N_4875);
or UO_748 (O_748,N_4519,N_4102);
nand UO_749 (O_749,N_4158,N_4866);
nand UO_750 (O_750,N_4720,N_4182);
nor UO_751 (O_751,N_4568,N_4600);
or UO_752 (O_752,N_4419,N_4405);
and UO_753 (O_753,N_4965,N_4901);
or UO_754 (O_754,N_4895,N_4577);
or UO_755 (O_755,N_4416,N_4198);
nor UO_756 (O_756,N_4089,N_4486);
nor UO_757 (O_757,N_4253,N_4187);
nand UO_758 (O_758,N_4411,N_4149);
and UO_759 (O_759,N_4730,N_4337);
or UO_760 (O_760,N_4964,N_4027);
nor UO_761 (O_761,N_4120,N_4906);
and UO_762 (O_762,N_4420,N_4430);
or UO_763 (O_763,N_4668,N_4178);
nand UO_764 (O_764,N_4220,N_4205);
or UO_765 (O_765,N_4930,N_4858);
and UO_766 (O_766,N_4075,N_4047);
nand UO_767 (O_767,N_4752,N_4060);
and UO_768 (O_768,N_4722,N_4381);
or UO_769 (O_769,N_4395,N_4964);
and UO_770 (O_770,N_4419,N_4751);
nor UO_771 (O_771,N_4117,N_4316);
and UO_772 (O_772,N_4173,N_4422);
nand UO_773 (O_773,N_4431,N_4836);
nand UO_774 (O_774,N_4310,N_4961);
and UO_775 (O_775,N_4721,N_4053);
nand UO_776 (O_776,N_4445,N_4484);
nand UO_777 (O_777,N_4547,N_4582);
nor UO_778 (O_778,N_4603,N_4376);
xnor UO_779 (O_779,N_4843,N_4712);
and UO_780 (O_780,N_4669,N_4165);
and UO_781 (O_781,N_4136,N_4539);
nand UO_782 (O_782,N_4565,N_4727);
nand UO_783 (O_783,N_4492,N_4417);
or UO_784 (O_784,N_4695,N_4742);
and UO_785 (O_785,N_4559,N_4354);
nand UO_786 (O_786,N_4437,N_4951);
or UO_787 (O_787,N_4426,N_4539);
nand UO_788 (O_788,N_4632,N_4790);
and UO_789 (O_789,N_4622,N_4448);
nand UO_790 (O_790,N_4563,N_4115);
xor UO_791 (O_791,N_4684,N_4604);
and UO_792 (O_792,N_4778,N_4968);
nand UO_793 (O_793,N_4126,N_4149);
nand UO_794 (O_794,N_4988,N_4853);
and UO_795 (O_795,N_4169,N_4436);
nor UO_796 (O_796,N_4478,N_4323);
and UO_797 (O_797,N_4995,N_4739);
or UO_798 (O_798,N_4950,N_4979);
nor UO_799 (O_799,N_4798,N_4040);
nor UO_800 (O_800,N_4115,N_4847);
nand UO_801 (O_801,N_4856,N_4609);
nand UO_802 (O_802,N_4510,N_4862);
nand UO_803 (O_803,N_4139,N_4841);
nor UO_804 (O_804,N_4307,N_4721);
or UO_805 (O_805,N_4529,N_4222);
or UO_806 (O_806,N_4537,N_4165);
nand UO_807 (O_807,N_4207,N_4081);
nor UO_808 (O_808,N_4968,N_4020);
nor UO_809 (O_809,N_4403,N_4701);
and UO_810 (O_810,N_4788,N_4059);
or UO_811 (O_811,N_4989,N_4948);
nor UO_812 (O_812,N_4399,N_4776);
xor UO_813 (O_813,N_4921,N_4245);
xnor UO_814 (O_814,N_4370,N_4271);
and UO_815 (O_815,N_4225,N_4711);
or UO_816 (O_816,N_4359,N_4619);
and UO_817 (O_817,N_4035,N_4844);
and UO_818 (O_818,N_4889,N_4101);
and UO_819 (O_819,N_4139,N_4948);
or UO_820 (O_820,N_4790,N_4776);
and UO_821 (O_821,N_4519,N_4891);
or UO_822 (O_822,N_4068,N_4346);
nor UO_823 (O_823,N_4759,N_4606);
and UO_824 (O_824,N_4405,N_4199);
and UO_825 (O_825,N_4081,N_4960);
or UO_826 (O_826,N_4434,N_4436);
nor UO_827 (O_827,N_4118,N_4353);
nand UO_828 (O_828,N_4467,N_4076);
or UO_829 (O_829,N_4327,N_4378);
nand UO_830 (O_830,N_4796,N_4181);
or UO_831 (O_831,N_4346,N_4466);
nor UO_832 (O_832,N_4611,N_4764);
nor UO_833 (O_833,N_4804,N_4011);
nand UO_834 (O_834,N_4841,N_4047);
or UO_835 (O_835,N_4759,N_4915);
and UO_836 (O_836,N_4452,N_4170);
nand UO_837 (O_837,N_4241,N_4058);
nand UO_838 (O_838,N_4889,N_4484);
nand UO_839 (O_839,N_4210,N_4931);
or UO_840 (O_840,N_4249,N_4759);
or UO_841 (O_841,N_4885,N_4930);
nor UO_842 (O_842,N_4405,N_4745);
nor UO_843 (O_843,N_4079,N_4748);
nand UO_844 (O_844,N_4614,N_4059);
nor UO_845 (O_845,N_4223,N_4228);
and UO_846 (O_846,N_4819,N_4029);
or UO_847 (O_847,N_4657,N_4132);
nor UO_848 (O_848,N_4659,N_4900);
or UO_849 (O_849,N_4701,N_4483);
or UO_850 (O_850,N_4564,N_4207);
or UO_851 (O_851,N_4802,N_4427);
nor UO_852 (O_852,N_4606,N_4453);
and UO_853 (O_853,N_4245,N_4238);
nand UO_854 (O_854,N_4835,N_4977);
nand UO_855 (O_855,N_4854,N_4616);
nand UO_856 (O_856,N_4604,N_4965);
nor UO_857 (O_857,N_4811,N_4274);
nor UO_858 (O_858,N_4956,N_4804);
and UO_859 (O_859,N_4029,N_4380);
nand UO_860 (O_860,N_4787,N_4541);
or UO_861 (O_861,N_4634,N_4936);
nand UO_862 (O_862,N_4303,N_4790);
and UO_863 (O_863,N_4524,N_4185);
or UO_864 (O_864,N_4383,N_4910);
or UO_865 (O_865,N_4696,N_4519);
and UO_866 (O_866,N_4700,N_4379);
and UO_867 (O_867,N_4989,N_4276);
and UO_868 (O_868,N_4619,N_4078);
nand UO_869 (O_869,N_4211,N_4675);
or UO_870 (O_870,N_4358,N_4326);
nor UO_871 (O_871,N_4976,N_4414);
and UO_872 (O_872,N_4698,N_4491);
nor UO_873 (O_873,N_4866,N_4310);
and UO_874 (O_874,N_4213,N_4053);
nand UO_875 (O_875,N_4832,N_4683);
or UO_876 (O_876,N_4083,N_4320);
nand UO_877 (O_877,N_4526,N_4563);
nor UO_878 (O_878,N_4505,N_4380);
nand UO_879 (O_879,N_4586,N_4621);
or UO_880 (O_880,N_4762,N_4985);
or UO_881 (O_881,N_4226,N_4311);
nor UO_882 (O_882,N_4095,N_4620);
nor UO_883 (O_883,N_4711,N_4231);
and UO_884 (O_884,N_4350,N_4388);
and UO_885 (O_885,N_4769,N_4621);
and UO_886 (O_886,N_4022,N_4808);
and UO_887 (O_887,N_4877,N_4651);
and UO_888 (O_888,N_4757,N_4740);
and UO_889 (O_889,N_4463,N_4293);
and UO_890 (O_890,N_4922,N_4609);
or UO_891 (O_891,N_4664,N_4355);
or UO_892 (O_892,N_4990,N_4535);
nor UO_893 (O_893,N_4260,N_4635);
or UO_894 (O_894,N_4463,N_4667);
or UO_895 (O_895,N_4675,N_4616);
and UO_896 (O_896,N_4365,N_4401);
and UO_897 (O_897,N_4600,N_4374);
nand UO_898 (O_898,N_4089,N_4543);
or UO_899 (O_899,N_4669,N_4832);
and UO_900 (O_900,N_4144,N_4570);
nand UO_901 (O_901,N_4340,N_4953);
nand UO_902 (O_902,N_4024,N_4077);
and UO_903 (O_903,N_4061,N_4761);
nor UO_904 (O_904,N_4011,N_4230);
and UO_905 (O_905,N_4981,N_4707);
nor UO_906 (O_906,N_4170,N_4687);
nand UO_907 (O_907,N_4834,N_4827);
nor UO_908 (O_908,N_4997,N_4045);
nand UO_909 (O_909,N_4701,N_4551);
nor UO_910 (O_910,N_4475,N_4237);
or UO_911 (O_911,N_4358,N_4590);
or UO_912 (O_912,N_4362,N_4236);
or UO_913 (O_913,N_4029,N_4062);
or UO_914 (O_914,N_4844,N_4572);
or UO_915 (O_915,N_4664,N_4178);
nor UO_916 (O_916,N_4668,N_4776);
xnor UO_917 (O_917,N_4595,N_4039);
nor UO_918 (O_918,N_4627,N_4749);
and UO_919 (O_919,N_4293,N_4308);
or UO_920 (O_920,N_4996,N_4375);
or UO_921 (O_921,N_4617,N_4299);
nor UO_922 (O_922,N_4531,N_4092);
and UO_923 (O_923,N_4290,N_4502);
nor UO_924 (O_924,N_4988,N_4142);
nor UO_925 (O_925,N_4599,N_4957);
or UO_926 (O_926,N_4560,N_4222);
or UO_927 (O_927,N_4234,N_4049);
nor UO_928 (O_928,N_4464,N_4611);
nand UO_929 (O_929,N_4691,N_4478);
or UO_930 (O_930,N_4555,N_4470);
and UO_931 (O_931,N_4557,N_4643);
or UO_932 (O_932,N_4291,N_4869);
nor UO_933 (O_933,N_4522,N_4281);
nand UO_934 (O_934,N_4286,N_4551);
and UO_935 (O_935,N_4862,N_4464);
or UO_936 (O_936,N_4355,N_4799);
nand UO_937 (O_937,N_4396,N_4343);
or UO_938 (O_938,N_4430,N_4115);
nor UO_939 (O_939,N_4388,N_4946);
or UO_940 (O_940,N_4423,N_4545);
or UO_941 (O_941,N_4010,N_4617);
nand UO_942 (O_942,N_4315,N_4678);
and UO_943 (O_943,N_4437,N_4468);
or UO_944 (O_944,N_4380,N_4314);
nor UO_945 (O_945,N_4509,N_4491);
nand UO_946 (O_946,N_4774,N_4041);
xor UO_947 (O_947,N_4532,N_4763);
and UO_948 (O_948,N_4346,N_4837);
nand UO_949 (O_949,N_4368,N_4763);
nor UO_950 (O_950,N_4317,N_4415);
and UO_951 (O_951,N_4366,N_4502);
nor UO_952 (O_952,N_4200,N_4326);
or UO_953 (O_953,N_4479,N_4769);
and UO_954 (O_954,N_4581,N_4623);
nor UO_955 (O_955,N_4034,N_4220);
nor UO_956 (O_956,N_4742,N_4234);
nand UO_957 (O_957,N_4176,N_4454);
nor UO_958 (O_958,N_4813,N_4099);
and UO_959 (O_959,N_4246,N_4138);
and UO_960 (O_960,N_4986,N_4088);
or UO_961 (O_961,N_4212,N_4861);
nor UO_962 (O_962,N_4053,N_4717);
or UO_963 (O_963,N_4688,N_4607);
nor UO_964 (O_964,N_4089,N_4481);
or UO_965 (O_965,N_4508,N_4336);
nand UO_966 (O_966,N_4126,N_4386);
or UO_967 (O_967,N_4891,N_4588);
nand UO_968 (O_968,N_4111,N_4612);
or UO_969 (O_969,N_4393,N_4317);
nor UO_970 (O_970,N_4884,N_4375);
or UO_971 (O_971,N_4345,N_4382);
or UO_972 (O_972,N_4206,N_4884);
nor UO_973 (O_973,N_4106,N_4424);
nand UO_974 (O_974,N_4516,N_4728);
nor UO_975 (O_975,N_4514,N_4326);
or UO_976 (O_976,N_4860,N_4585);
or UO_977 (O_977,N_4973,N_4492);
nor UO_978 (O_978,N_4306,N_4099);
or UO_979 (O_979,N_4423,N_4592);
and UO_980 (O_980,N_4830,N_4956);
nor UO_981 (O_981,N_4154,N_4981);
and UO_982 (O_982,N_4035,N_4990);
or UO_983 (O_983,N_4543,N_4939);
and UO_984 (O_984,N_4754,N_4806);
nand UO_985 (O_985,N_4814,N_4626);
nand UO_986 (O_986,N_4865,N_4354);
or UO_987 (O_987,N_4406,N_4483);
and UO_988 (O_988,N_4727,N_4240);
and UO_989 (O_989,N_4707,N_4961);
nand UO_990 (O_990,N_4116,N_4653);
nor UO_991 (O_991,N_4248,N_4093);
or UO_992 (O_992,N_4749,N_4909);
nor UO_993 (O_993,N_4168,N_4089);
and UO_994 (O_994,N_4925,N_4346);
and UO_995 (O_995,N_4487,N_4337);
nand UO_996 (O_996,N_4631,N_4521);
nor UO_997 (O_997,N_4270,N_4701);
and UO_998 (O_998,N_4225,N_4281);
and UO_999 (O_999,N_4760,N_4247);
endmodule