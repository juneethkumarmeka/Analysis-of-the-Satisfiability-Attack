module basic_500_3000_500_50_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_117,In_291);
nand U1 (N_1,In_472,In_358);
xor U2 (N_2,In_442,In_407);
nor U3 (N_3,In_342,In_46);
or U4 (N_4,In_238,In_137);
nor U5 (N_5,In_32,In_98);
and U6 (N_6,In_90,In_272);
nand U7 (N_7,In_255,In_419);
or U8 (N_8,In_270,In_11);
or U9 (N_9,In_355,In_375);
nand U10 (N_10,In_313,In_421);
nand U11 (N_11,In_391,In_86);
xnor U12 (N_12,In_151,In_16);
nor U13 (N_13,In_241,In_447);
nand U14 (N_14,In_3,In_108);
or U15 (N_15,In_463,In_274);
or U16 (N_16,In_148,In_326);
xnor U17 (N_17,In_247,In_252);
and U18 (N_18,In_393,In_167);
and U19 (N_19,In_55,In_27);
nor U20 (N_20,In_115,In_344);
xnor U21 (N_21,In_495,In_23);
or U22 (N_22,In_100,In_131);
xor U23 (N_23,In_277,In_488);
nor U24 (N_24,In_94,In_244);
and U25 (N_25,In_194,In_411);
nand U26 (N_26,In_417,In_73);
and U27 (N_27,In_302,In_481);
and U28 (N_28,In_233,In_26);
or U29 (N_29,In_65,In_307);
and U30 (N_30,In_434,In_410);
nand U31 (N_31,In_125,In_455);
nand U32 (N_32,In_394,In_497);
nand U33 (N_33,In_44,In_459);
or U34 (N_34,In_210,In_287);
xor U35 (N_35,In_61,In_234);
nor U36 (N_36,In_118,In_266);
and U37 (N_37,In_8,In_378);
or U38 (N_38,In_352,In_193);
nand U39 (N_39,In_365,In_286);
and U40 (N_40,In_328,In_105);
xnor U41 (N_41,In_418,In_113);
nor U42 (N_42,In_133,In_398);
xor U43 (N_43,In_53,In_437);
nor U44 (N_44,In_412,In_308);
and U45 (N_45,In_17,In_45);
nor U46 (N_46,In_297,In_279);
nor U47 (N_47,In_70,In_168);
or U48 (N_48,In_155,In_35);
and U49 (N_49,In_261,In_310);
or U50 (N_50,In_205,In_356);
or U51 (N_51,In_165,In_329);
and U52 (N_52,In_14,In_119);
nand U53 (N_53,In_350,In_385);
nand U54 (N_54,In_116,In_305);
nor U55 (N_55,In_379,In_346);
nand U56 (N_56,In_106,In_92);
xnor U57 (N_57,In_217,In_34);
nor U58 (N_58,In_7,In_80);
and U59 (N_59,In_317,In_271);
or U60 (N_60,N_25,In_134);
xor U61 (N_61,In_409,In_77);
or U62 (N_62,In_213,In_207);
or U63 (N_63,In_284,In_337);
xnor U64 (N_64,In_36,N_37);
or U65 (N_65,N_52,In_20);
and U66 (N_66,In_62,In_95);
and U67 (N_67,N_19,In_243);
xor U68 (N_68,In_333,In_477);
nand U69 (N_69,In_450,In_97);
xnor U70 (N_70,In_303,In_202);
or U71 (N_71,In_367,In_354);
or U72 (N_72,N_57,N_44);
or U73 (N_73,In_192,In_292);
nor U74 (N_74,In_465,In_248);
and U75 (N_75,In_401,In_179);
nor U76 (N_76,In_327,In_109);
nand U77 (N_77,In_246,In_38);
nor U78 (N_78,In_178,N_32);
xnor U79 (N_79,In_309,In_84);
nand U80 (N_80,In_479,In_404);
nor U81 (N_81,In_147,N_39);
or U82 (N_82,In_226,In_107);
xnor U83 (N_83,In_196,N_13);
nand U84 (N_84,In_439,In_216);
and U85 (N_85,In_275,In_81);
or U86 (N_86,In_458,In_225);
xor U87 (N_87,N_56,In_332);
nor U88 (N_88,In_149,In_273);
and U89 (N_89,In_473,In_215);
nor U90 (N_90,In_397,In_158);
and U91 (N_91,In_175,In_129);
nand U92 (N_92,In_183,In_199);
and U93 (N_93,In_184,In_316);
and U94 (N_94,N_33,In_232);
xnor U95 (N_95,In_114,In_452);
nor U96 (N_96,In_67,In_6);
or U97 (N_97,In_209,In_185);
xnor U98 (N_98,In_290,In_257);
xnor U99 (N_99,In_28,In_264);
and U100 (N_100,In_460,In_161);
nor U101 (N_101,In_164,In_445);
nand U102 (N_102,In_312,N_8);
nor U103 (N_103,In_176,N_18);
nand U104 (N_104,In_403,In_338);
and U105 (N_105,In_120,In_415);
nor U106 (N_106,In_366,In_4);
or U107 (N_107,In_221,In_295);
xnor U108 (N_108,In_75,In_111);
and U109 (N_109,In_282,In_469);
nor U110 (N_110,In_369,In_363);
xnor U111 (N_111,In_123,In_474);
nand U112 (N_112,In_9,In_103);
and U113 (N_113,In_211,In_467);
or U114 (N_114,In_150,In_408);
or U115 (N_115,In_440,N_47);
or U116 (N_116,In_66,In_396);
and U117 (N_117,In_466,In_159);
nand U118 (N_118,In_195,In_222);
and U119 (N_119,In_143,In_174);
xnor U120 (N_120,In_145,In_132);
or U121 (N_121,In_364,In_444);
or U122 (N_122,N_119,In_42);
or U123 (N_123,In_0,In_60);
or U124 (N_124,In_99,In_163);
nor U125 (N_125,In_347,In_349);
xnor U126 (N_126,In_156,N_100);
nor U127 (N_127,In_484,N_92);
nor U128 (N_128,In_37,In_471);
nor U129 (N_129,In_300,In_424);
nand U130 (N_130,N_10,In_334);
nor U131 (N_131,N_86,In_496);
nor U132 (N_132,In_24,N_78);
or U133 (N_133,In_498,In_457);
nor U134 (N_134,In_283,In_443);
nand U135 (N_135,In_227,In_402);
or U136 (N_136,N_21,In_218);
nor U137 (N_137,In_79,In_15);
nor U138 (N_138,In_493,In_50);
xor U139 (N_139,In_235,In_1);
nor U140 (N_140,N_23,In_486);
nand U141 (N_141,In_47,In_262);
xnor U142 (N_142,In_376,In_315);
or U143 (N_143,N_75,In_276);
or U144 (N_144,In_335,In_220);
or U145 (N_145,In_438,In_51);
nor U146 (N_146,In_399,In_370);
or U147 (N_147,In_198,In_30);
and U148 (N_148,N_38,In_476);
or U149 (N_149,In_188,In_311);
nor U150 (N_150,In_426,In_478);
nor U151 (N_151,In_435,In_166);
nor U152 (N_152,N_72,In_231);
or U153 (N_153,In_433,N_85);
nor U154 (N_154,In_322,In_331);
and U155 (N_155,In_13,In_395);
nor U156 (N_156,N_80,In_280);
or U157 (N_157,N_1,In_456);
xnor U158 (N_158,N_104,In_360);
or U159 (N_159,In_281,In_406);
nor U160 (N_160,In_223,In_386);
nor U161 (N_161,In_138,In_212);
nor U162 (N_162,N_101,In_362);
xnor U163 (N_163,In_96,In_206);
nor U164 (N_164,In_160,N_110);
or U165 (N_165,In_173,In_208);
nand U166 (N_166,In_74,In_441);
nand U167 (N_167,N_34,In_368);
and U168 (N_168,In_240,In_197);
nor U169 (N_169,N_31,N_114);
nor U170 (N_170,N_79,N_49);
or U171 (N_171,In_490,In_63);
xor U172 (N_172,N_83,In_239);
nand U173 (N_173,N_40,In_373);
or U174 (N_174,In_269,In_321);
or U175 (N_175,In_285,N_60);
or U176 (N_176,In_374,In_71);
xnor U177 (N_177,In_201,In_122);
nor U178 (N_178,N_111,In_136);
or U179 (N_179,In_323,In_189);
nor U180 (N_180,N_24,N_71);
and U181 (N_181,In_304,In_72);
xor U182 (N_182,In_325,In_449);
and U183 (N_183,N_143,In_22);
and U184 (N_184,N_127,In_88);
or U185 (N_185,In_170,N_68);
xnor U186 (N_186,N_9,In_91);
and U187 (N_187,In_489,In_341);
xnor U188 (N_188,N_162,In_104);
and U189 (N_189,N_16,N_76);
or U190 (N_190,In_339,N_123);
xor U191 (N_191,In_324,N_43);
nor U192 (N_192,N_14,N_84);
nand U193 (N_193,N_168,N_98);
or U194 (N_194,In_390,In_392);
nor U195 (N_195,N_102,In_40);
or U196 (N_196,In_31,In_461);
xnor U197 (N_197,In_144,N_126);
xnor U198 (N_198,In_253,In_237);
and U199 (N_199,N_146,N_165);
nor U200 (N_200,In_33,In_351);
xor U201 (N_201,N_154,In_83);
and U202 (N_202,In_127,N_0);
xnor U203 (N_203,In_318,N_130);
nand U204 (N_204,N_6,N_29);
and U205 (N_205,In_250,In_68);
xor U206 (N_206,N_4,In_470);
or U207 (N_207,In_112,In_432);
nand U208 (N_208,In_357,N_109);
nor U209 (N_209,In_359,In_87);
or U210 (N_210,N_164,N_62);
nor U211 (N_211,N_73,N_145);
xnor U212 (N_212,In_128,N_61);
or U213 (N_213,N_118,N_12);
nand U214 (N_214,In_5,In_177);
or U215 (N_215,In_414,N_26);
or U216 (N_216,N_2,In_25);
and U217 (N_217,In_380,In_361);
or U218 (N_218,N_161,In_330);
and U219 (N_219,N_135,In_59);
and U220 (N_220,In_454,In_485);
xnor U221 (N_221,N_129,N_170);
xor U222 (N_222,In_482,N_113);
and U223 (N_223,N_107,N_42);
nand U224 (N_224,N_103,In_182);
nand U225 (N_225,N_173,N_176);
xnor U226 (N_226,N_88,N_87);
nand U227 (N_227,In_340,N_148);
or U228 (N_228,N_17,N_155);
or U229 (N_229,N_137,N_133);
and U230 (N_230,In_29,In_85);
and U231 (N_231,N_69,N_59);
xnor U232 (N_232,In_19,N_144);
nor U233 (N_233,In_377,N_58);
and U234 (N_234,In_314,In_288);
xor U235 (N_235,N_48,N_3);
nand U236 (N_236,In_256,In_43);
or U237 (N_237,N_160,N_151);
nor U238 (N_238,N_117,N_63);
nand U239 (N_239,In_251,In_260);
nand U240 (N_240,In_371,N_55);
and U241 (N_241,N_219,In_422);
or U242 (N_242,N_184,N_15);
xor U243 (N_243,N_28,In_446);
and U244 (N_244,In_180,N_167);
xor U245 (N_245,N_136,In_203);
nand U246 (N_246,N_97,N_233);
and U247 (N_247,In_157,N_152);
nand U248 (N_248,N_35,In_135);
and U249 (N_249,N_197,In_453);
nor U250 (N_250,N_231,N_64);
nor U251 (N_251,In_427,N_27);
or U252 (N_252,In_56,N_190);
xor U253 (N_253,N_226,In_480);
or U254 (N_254,In_18,In_187);
xnor U255 (N_255,In_265,N_220);
and U256 (N_256,N_112,In_296);
xnor U257 (N_257,In_10,N_189);
nor U258 (N_258,N_178,In_468);
or U259 (N_259,N_149,In_153);
xor U260 (N_260,In_228,N_191);
or U261 (N_261,N_66,In_124);
or U262 (N_262,N_138,N_169);
xnor U263 (N_263,N_131,N_185);
or U264 (N_264,N_91,In_289);
nor U265 (N_265,N_194,N_208);
nand U266 (N_266,N_225,In_384);
nor U267 (N_267,N_134,In_383);
nor U268 (N_268,In_353,In_430);
nor U269 (N_269,In_121,N_53);
nand U270 (N_270,N_90,N_214);
nor U271 (N_271,In_82,In_89);
xnor U272 (N_272,In_451,In_487);
and U273 (N_273,In_78,N_94);
nor U274 (N_274,In_425,In_214);
nand U275 (N_275,N_36,N_210);
xor U276 (N_276,In_464,In_110);
and U277 (N_277,N_209,In_278);
or U278 (N_278,In_499,In_268);
and U279 (N_279,N_65,In_49);
xor U280 (N_280,In_242,N_236);
xnor U281 (N_281,N_95,In_249);
xor U282 (N_282,N_188,N_116);
nor U283 (N_283,N_46,N_142);
or U284 (N_284,N_181,In_293);
or U285 (N_285,N_41,In_93);
xnor U286 (N_286,In_429,In_301);
nor U287 (N_287,N_166,N_141);
xor U288 (N_288,N_93,In_320);
or U289 (N_289,N_177,In_388);
nor U290 (N_290,N_212,N_234);
xor U291 (N_291,N_195,N_22);
xor U292 (N_292,In_382,In_413);
nor U293 (N_293,N_207,N_193);
or U294 (N_294,N_45,In_428);
nor U295 (N_295,In_389,N_150);
or U296 (N_296,In_319,In_306);
nor U297 (N_297,In_200,In_141);
xnor U298 (N_298,In_54,N_174);
and U299 (N_299,N_235,N_115);
nor U300 (N_300,N_279,N_289);
nand U301 (N_301,N_241,In_423);
or U302 (N_302,N_280,N_179);
nand U303 (N_303,In_142,In_219);
nor U304 (N_304,N_269,N_5);
nor U305 (N_305,In_236,N_221);
or U306 (N_306,In_21,N_54);
nand U307 (N_307,In_191,In_405);
nor U308 (N_308,In_336,In_172);
nor U309 (N_309,In_267,In_39);
nor U310 (N_310,N_296,N_240);
nor U311 (N_311,In_372,N_77);
xnor U312 (N_312,In_416,In_57);
nor U313 (N_313,N_252,N_82);
or U314 (N_314,In_169,In_58);
xor U315 (N_315,N_256,In_139);
nor U316 (N_316,In_345,N_261);
xor U317 (N_317,N_213,N_51);
nand U318 (N_318,In_126,In_76);
xor U319 (N_319,N_278,N_198);
nor U320 (N_320,N_106,N_259);
xnor U321 (N_321,N_224,In_431);
nor U322 (N_322,In_69,N_294);
nor U323 (N_323,In_420,In_387);
nor U324 (N_324,N_211,N_120);
and U325 (N_325,N_132,In_64);
nand U326 (N_326,N_175,N_140);
xnor U327 (N_327,In_462,N_253);
nand U328 (N_328,N_257,N_270);
and U329 (N_329,N_200,N_215);
nand U330 (N_330,N_254,N_237);
and U331 (N_331,N_288,N_159);
and U332 (N_332,N_182,In_101);
or U333 (N_333,N_216,N_265);
nor U334 (N_334,N_203,N_285);
nor U335 (N_335,N_271,N_283);
nor U336 (N_336,N_122,N_81);
nand U337 (N_337,N_290,In_258);
xnor U338 (N_338,In_298,N_202);
xnor U339 (N_339,In_259,In_181);
xnor U340 (N_340,In_294,N_273);
xor U341 (N_341,N_217,N_196);
xor U342 (N_342,N_239,N_96);
and U343 (N_343,N_186,N_287);
nor U344 (N_344,N_299,N_244);
or U345 (N_345,N_105,N_99);
nor U346 (N_346,In_492,N_297);
and U347 (N_347,N_156,In_12);
or U348 (N_348,In_245,N_50);
nand U349 (N_349,N_121,In_152);
nand U350 (N_350,N_205,N_293);
nand U351 (N_351,N_229,N_251);
or U352 (N_352,In_171,N_258);
xnor U353 (N_353,N_255,N_20);
nand U354 (N_354,N_201,N_277);
nor U355 (N_355,In_190,In_204);
nor U356 (N_356,In_230,In_140);
xnor U357 (N_357,In_263,N_223);
xor U358 (N_358,N_248,N_74);
xor U359 (N_359,N_157,N_183);
xnor U360 (N_360,In_494,N_349);
and U361 (N_361,N_242,In_475);
nor U362 (N_362,N_347,In_2);
and U363 (N_363,N_67,N_355);
xor U364 (N_364,N_308,N_322);
and U365 (N_365,In_102,N_330);
and U366 (N_366,N_192,N_320);
xnor U367 (N_367,N_351,N_337);
or U368 (N_368,N_321,N_313);
and U369 (N_369,N_295,N_335);
nor U370 (N_370,In_343,N_250);
xor U371 (N_371,N_353,N_89);
xor U372 (N_372,In_491,N_262);
xor U373 (N_373,N_307,N_218);
nor U374 (N_374,N_260,N_206);
nand U375 (N_375,N_147,N_312);
xor U376 (N_376,N_243,N_204);
or U377 (N_377,N_315,N_323);
nor U378 (N_378,N_305,N_329);
and U379 (N_379,N_359,N_222);
nor U380 (N_380,N_344,N_227);
nor U381 (N_381,N_272,N_286);
nand U382 (N_382,N_325,N_350);
or U383 (N_383,N_199,N_291);
nand U384 (N_384,In_52,N_187);
xnor U385 (N_385,N_266,In_146);
xor U386 (N_386,N_336,N_70);
xor U387 (N_387,N_342,N_139);
and U388 (N_388,N_303,N_318);
nor U389 (N_389,N_301,N_354);
xor U390 (N_390,N_317,N_232);
nand U391 (N_391,N_309,N_298);
nor U392 (N_392,In_130,N_332);
or U393 (N_393,In_162,N_275);
xnor U394 (N_394,N_274,N_358);
xor U395 (N_395,In_48,N_339);
xor U396 (N_396,N_249,N_292);
nor U397 (N_397,N_246,N_300);
and U398 (N_398,N_352,In_448);
nand U399 (N_399,N_108,N_245);
or U400 (N_400,In_348,N_324);
nor U401 (N_401,N_125,N_333);
and U402 (N_402,N_327,In_254);
and U403 (N_403,N_302,In_186);
xor U404 (N_404,N_11,N_281);
and U405 (N_405,N_171,N_341);
nand U406 (N_406,N_172,N_180);
or U407 (N_407,In_483,N_310);
nand U408 (N_408,N_282,N_340);
nor U409 (N_409,N_228,N_345);
nand U410 (N_410,N_314,N_346);
xnor U411 (N_411,N_163,N_264);
nor U412 (N_412,N_247,In_299);
and U413 (N_413,N_356,In_436);
nor U414 (N_414,N_306,In_154);
xnor U415 (N_415,N_7,N_338);
or U416 (N_416,N_311,In_400);
and U417 (N_417,N_304,N_230);
nand U418 (N_418,N_158,In_229);
and U419 (N_419,N_328,In_41);
xor U420 (N_420,N_402,N_357);
xnor U421 (N_421,N_390,N_416);
xnor U422 (N_422,N_375,N_396);
xnor U423 (N_423,N_378,N_380);
nand U424 (N_424,N_319,N_364);
or U425 (N_425,N_367,N_394);
and U426 (N_426,N_267,N_382);
xor U427 (N_427,N_404,N_418);
nor U428 (N_428,N_401,N_276);
and U429 (N_429,N_374,N_403);
xnor U430 (N_430,N_348,N_369);
nand U431 (N_431,N_371,N_361);
nor U432 (N_432,N_331,N_377);
and U433 (N_433,N_365,N_366);
and U434 (N_434,N_238,N_372);
nor U435 (N_435,N_268,N_379);
nand U436 (N_436,N_334,N_412);
and U437 (N_437,N_343,N_376);
or U438 (N_438,N_384,N_388);
nor U439 (N_439,In_381,N_398);
xor U440 (N_440,N_263,N_399);
nor U441 (N_441,N_362,N_363);
or U442 (N_442,N_410,N_316);
xnor U443 (N_443,N_360,N_417);
or U444 (N_444,N_406,N_370);
xor U445 (N_445,N_381,N_415);
xor U446 (N_446,N_373,N_383);
nor U447 (N_447,N_153,N_385);
nand U448 (N_448,N_124,N_368);
xor U449 (N_449,N_284,N_400);
xnor U450 (N_450,N_387,N_30);
or U451 (N_451,N_391,N_411);
xor U452 (N_452,N_419,In_224);
or U453 (N_453,N_413,N_408);
xor U454 (N_454,N_386,N_407);
and U455 (N_455,N_393,N_414);
xnor U456 (N_456,N_326,N_395);
and U457 (N_457,N_405,N_389);
and U458 (N_458,N_128,N_392);
or U459 (N_459,N_397,N_409);
or U460 (N_460,N_364,N_371);
and U461 (N_461,N_128,N_408);
or U462 (N_462,N_263,N_400);
nand U463 (N_463,In_381,N_391);
and U464 (N_464,N_383,N_403);
nand U465 (N_465,N_383,N_276);
and U466 (N_466,N_409,N_392);
and U467 (N_467,N_267,N_413);
and U468 (N_468,N_334,N_376);
nand U469 (N_469,N_377,N_365);
nand U470 (N_470,N_385,N_415);
or U471 (N_471,N_368,N_334);
and U472 (N_472,N_369,N_407);
xnor U473 (N_473,N_343,N_400);
and U474 (N_474,N_410,N_375);
nand U475 (N_475,N_371,N_405);
nand U476 (N_476,N_415,N_395);
nand U477 (N_477,N_401,N_395);
nor U478 (N_478,N_386,N_403);
xnor U479 (N_479,N_30,N_392);
nor U480 (N_480,N_422,N_456);
nand U481 (N_481,N_478,N_464);
nand U482 (N_482,N_455,N_445);
or U483 (N_483,N_470,N_442);
nor U484 (N_484,N_457,N_469);
xor U485 (N_485,N_420,N_447);
nand U486 (N_486,N_463,N_452);
nand U487 (N_487,N_429,N_448);
nand U488 (N_488,N_454,N_468);
or U489 (N_489,N_438,N_428);
xor U490 (N_490,N_421,N_451);
nand U491 (N_491,N_424,N_462);
nand U492 (N_492,N_434,N_465);
nor U493 (N_493,N_432,N_435);
nand U494 (N_494,N_427,N_436);
nand U495 (N_495,N_440,N_430);
nand U496 (N_496,N_444,N_426);
and U497 (N_497,N_476,N_443);
nand U498 (N_498,N_433,N_466);
nor U499 (N_499,N_467,N_453);
xor U500 (N_500,N_458,N_449);
nor U501 (N_501,N_471,N_473);
or U502 (N_502,N_460,N_479);
nand U503 (N_503,N_475,N_461);
or U504 (N_504,N_450,N_446);
nand U505 (N_505,N_459,N_477);
nor U506 (N_506,N_431,N_423);
or U507 (N_507,N_437,N_474);
xnor U508 (N_508,N_439,N_425);
nor U509 (N_509,N_441,N_472);
nor U510 (N_510,N_438,N_456);
and U511 (N_511,N_453,N_455);
xor U512 (N_512,N_479,N_470);
or U513 (N_513,N_440,N_474);
nand U514 (N_514,N_462,N_432);
or U515 (N_515,N_429,N_431);
and U516 (N_516,N_460,N_452);
nor U517 (N_517,N_424,N_426);
and U518 (N_518,N_472,N_467);
or U519 (N_519,N_448,N_453);
nand U520 (N_520,N_457,N_447);
and U521 (N_521,N_473,N_425);
nor U522 (N_522,N_425,N_476);
or U523 (N_523,N_466,N_426);
xnor U524 (N_524,N_464,N_426);
nor U525 (N_525,N_427,N_472);
or U526 (N_526,N_430,N_446);
xnor U527 (N_527,N_456,N_446);
nor U528 (N_528,N_423,N_456);
nor U529 (N_529,N_460,N_468);
nand U530 (N_530,N_433,N_462);
or U531 (N_531,N_468,N_436);
nand U532 (N_532,N_473,N_474);
or U533 (N_533,N_440,N_478);
xor U534 (N_534,N_461,N_421);
xnor U535 (N_535,N_468,N_444);
nor U536 (N_536,N_473,N_439);
xnor U537 (N_537,N_445,N_426);
and U538 (N_538,N_451,N_437);
nand U539 (N_539,N_426,N_458);
and U540 (N_540,N_481,N_536);
or U541 (N_541,N_498,N_488);
xnor U542 (N_542,N_486,N_483);
nor U543 (N_543,N_505,N_504);
and U544 (N_544,N_516,N_526);
nand U545 (N_545,N_503,N_506);
nor U546 (N_546,N_518,N_533);
nor U547 (N_547,N_517,N_484);
and U548 (N_548,N_485,N_508);
or U549 (N_549,N_521,N_491);
or U550 (N_550,N_482,N_514);
nand U551 (N_551,N_496,N_501);
nand U552 (N_552,N_513,N_500);
nand U553 (N_553,N_530,N_520);
xor U554 (N_554,N_507,N_492);
nor U555 (N_555,N_490,N_528);
xnor U556 (N_556,N_524,N_525);
or U557 (N_557,N_480,N_531);
xnor U558 (N_558,N_487,N_499);
nor U559 (N_559,N_489,N_522);
or U560 (N_560,N_493,N_539);
nand U561 (N_561,N_512,N_502);
or U562 (N_562,N_523,N_519);
or U563 (N_563,N_494,N_529);
xor U564 (N_564,N_527,N_511);
and U565 (N_565,N_497,N_537);
xor U566 (N_566,N_509,N_535);
xnor U567 (N_567,N_538,N_495);
nand U568 (N_568,N_532,N_515);
or U569 (N_569,N_534,N_510);
nor U570 (N_570,N_538,N_525);
nand U571 (N_571,N_517,N_485);
nor U572 (N_572,N_491,N_507);
nand U573 (N_573,N_536,N_484);
or U574 (N_574,N_482,N_481);
nor U575 (N_575,N_531,N_535);
nor U576 (N_576,N_512,N_498);
xnor U577 (N_577,N_523,N_482);
nand U578 (N_578,N_513,N_520);
nand U579 (N_579,N_517,N_539);
and U580 (N_580,N_483,N_522);
nand U581 (N_581,N_530,N_502);
or U582 (N_582,N_521,N_527);
xor U583 (N_583,N_529,N_509);
and U584 (N_584,N_499,N_490);
or U585 (N_585,N_497,N_501);
and U586 (N_586,N_519,N_535);
nand U587 (N_587,N_488,N_507);
or U588 (N_588,N_494,N_526);
or U589 (N_589,N_517,N_498);
nand U590 (N_590,N_496,N_516);
or U591 (N_591,N_509,N_502);
and U592 (N_592,N_501,N_528);
nand U593 (N_593,N_532,N_490);
nand U594 (N_594,N_538,N_481);
nand U595 (N_595,N_539,N_514);
nor U596 (N_596,N_496,N_493);
nand U597 (N_597,N_538,N_515);
nor U598 (N_598,N_527,N_526);
xor U599 (N_599,N_481,N_537);
and U600 (N_600,N_558,N_576);
xor U601 (N_601,N_567,N_579);
xor U602 (N_602,N_578,N_599);
nand U603 (N_603,N_596,N_565);
or U604 (N_604,N_548,N_586);
or U605 (N_605,N_542,N_540);
or U606 (N_606,N_577,N_580);
or U607 (N_607,N_561,N_553);
or U608 (N_608,N_588,N_571);
and U609 (N_609,N_562,N_564);
nand U610 (N_610,N_566,N_590);
xor U611 (N_611,N_585,N_549);
nand U612 (N_612,N_598,N_556);
and U613 (N_613,N_568,N_581);
nand U614 (N_614,N_554,N_552);
nand U615 (N_615,N_595,N_587);
and U616 (N_616,N_559,N_574);
nor U617 (N_617,N_569,N_584);
nand U618 (N_618,N_597,N_570);
or U619 (N_619,N_550,N_583);
nor U620 (N_620,N_551,N_582);
xor U621 (N_621,N_563,N_591);
nand U622 (N_622,N_572,N_544);
nor U623 (N_623,N_589,N_546);
nor U624 (N_624,N_541,N_545);
nand U625 (N_625,N_593,N_555);
and U626 (N_626,N_594,N_547);
xor U627 (N_627,N_543,N_557);
xor U628 (N_628,N_560,N_592);
nand U629 (N_629,N_573,N_575);
or U630 (N_630,N_561,N_542);
nand U631 (N_631,N_566,N_547);
xor U632 (N_632,N_574,N_598);
nand U633 (N_633,N_543,N_573);
or U634 (N_634,N_584,N_566);
xor U635 (N_635,N_569,N_548);
nor U636 (N_636,N_546,N_547);
xor U637 (N_637,N_570,N_581);
and U638 (N_638,N_542,N_578);
nand U639 (N_639,N_543,N_545);
xor U640 (N_640,N_540,N_543);
or U641 (N_641,N_599,N_540);
nand U642 (N_642,N_563,N_565);
or U643 (N_643,N_561,N_563);
or U644 (N_644,N_575,N_567);
nand U645 (N_645,N_584,N_548);
or U646 (N_646,N_550,N_570);
xor U647 (N_647,N_558,N_578);
nand U648 (N_648,N_595,N_562);
and U649 (N_649,N_574,N_565);
and U650 (N_650,N_560,N_546);
nand U651 (N_651,N_570,N_542);
or U652 (N_652,N_593,N_543);
xnor U653 (N_653,N_570,N_563);
nand U654 (N_654,N_557,N_544);
xnor U655 (N_655,N_552,N_546);
xnor U656 (N_656,N_564,N_542);
xor U657 (N_657,N_576,N_548);
and U658 (N_658,N_567,N_595);
nand U659 (N_659,N_571,N_553);
nand U660 (N_660,N_617,N_603);
or U661 (N_661,N_646,N_659);
xor U662 (N_662,N_655,N_654);
nand U663 (N_663,N_639,N_602);
nand U664 (N_664,N_634,N_622);
nor U665 (N_665,N_652,N_633);
or U666 (N_666,N_653,N_635);
and U667 (N_667,N_615,N_632);
or U668 (N_668,N_657,N_645);
nor U669 (N_669,N_651,N_637);
xnor U670 (N_670,N_647,N_601);
xor U671 (N_671,N_640,N_620);
nand U672 (N_672,N_608,N_619);
nor U673 (N_673,N_628,N_636);
and U674 (N_674,N_621,N_611);
nor U675 (N_675,N_623,N_627);
and U676 (N_676,N_643,N_618);
and U677 (N_677,N_609,N_626);
xor U678 (N_678,N_656,N_604);
and U679 (N_679,N_629,N_658);
nand U680 (N_680,N_605,N_641);
or U681 (N_681,N_614,N_630);
nand U682 (N_682,N_610,N_616);
nor U683 (N_683,N_642,N_613);
nor U684 (N_684,N_644,N_624);
nand U685 (N_685,N_600,N_631);
and U686 (N_686,N_638,N_649);
nand U687 (N_687,N_612,N_648);
nor U688 (N_688,N_650,N_607);
nor U689 (N_689,N_625,N_606);
nand U690 (N_690,N_635,N_633);
nand U691 (N_691,N_650,N_639);
xor U692 (N_692,N_645,N_654);
and U693 (N_693,N_606,N_610);
nor U694 (N_694,N_614,N_627);
xnor U695 (N_695,N_626,N_617);
and U696 (N_696,N_654,N_607);
xor U697 (N_697,N_642,N_611);
and U698 (N_698,N_646,N_645);
and U699 (N_699,N_601,N_618);
or U700 (N_700,N_619,N_647);
or U701 (N_701,N_643,N_650);
xor U702 (N_702,N_657,N_633);
and U703 (N_703,N_627,N_630);
or U704 (N_704,N_627,N_629);
nand U705 (N_705,N_602,N_606);
nor U706 (N_706,N_641,N_647);
nor U707 (N_707,N_635,N_636);
nor U708 (N_708,N_617,N_618);
and U709 (N_709,N_627,N_646);
or U710 (N_710,N_622,N_659);
nor U711 (N_711,N_622,N_647);
xnor U712 (N_712,N_653,N_650);
nor U713 (N_713,N_641,N_600);
or U714 (N_714,N_607,N_608);
nand U715 (N_715,N_658,N_623);
and U716 (N_716,N_649,N_659);
nand U717 (N_717,N_615,N_622);
nand U718 (N_718,N_614,N_615);
nand U719 (N_719,N_611,N_656);
nor U720 (N_720,N_713,N_663);
xor U721 (N_721,N_711,N_660);
nor U722 (N_722,N_671,N_703);
or U723 (N_723,N_694,N_690);
or U724 (N_724,N_683,N_665);
or U725 (N_725,N_708,N_696);
or U726 (N_726,N_684,N_688);
or U727 (N_727,N_662,N_679);
and U728 (N_728,N_673,N_701);
xor U729 (N_729,N_704,N_707);
xor U730 (N_730,N_668,N_706);
nor U731 (N_731,N_692,N_664);
xor U732 (N_732,N_666,N_670);
and U733 (N_733,N_681,N_674);
nand U734 (N_734,N_669,N_685);
nor U735 (N_735,N_695,N_718);
xnor U736 (N_736,N_667,N_710);
xor U737 (N_737,N_716,N_705);
and U738 (N_738,N_682,N_715);
and U739 (N_739,N_689,N_700);
nor U740 (N_740,N_661,N_699);
or U741 (N_741,N_672,N_712);
nand U742 (N_742,N_709,N_697);
nor U743 (N_743,N_677,N_686);
nor U744 (N_744,N_698,N_693);
xnor U745 (N_745,N_678,N_714);
and U746 (N_746,N_691,N_687);
nor U747 (N_747,N_680,N_717);
nor U748 (N_748,N_675,N_676);
and U749 (N_749,N_719,N_702);
nand U750 (N_750,N_690,N_673);
or U751 (N_751,N_677,N_711);
nor U752 (N_752,N_667,N_711);
nor U753 (N_753,N_711,N_680);
nor U754 (N_754,N_687,N_673);
or U755 (N_755,N_688,N_702);
nand U756 (N_756,N_692,N_695);
and U757 (N_757,N_662,N_715);
or U758 (N_758,N_717,N_698);
nor U759 (N_759,N_695,N_661);
or U760 (N_760,N_675,N_712);
and U761 (N_761,N_679,N_688);
and U762 (N_762,N_660,N_681);
xor U763 (N_763,N_696,N_695);
and U764 (N_764,N_681,N_661);
nor U765 (N_765,N_702,N_713);
or U766 (N_766,N_715,N_688);
xor U767 (N_767,N_676,N_688);
nor U768 (N_768,N_704,N_715);
xnor U769 (N_769,N_698,N_711);
and U770 (N_770,N_687,N_714);
and U771 (N_771,N_706,N_676);
and U772 (N_772,N_703,N_685);
nor U773 (N_773,N_670,N_685);
and U774 (N_774,N_696,N_690);
and U775 (N_775,N_678,N_716);
nor U776 (N_776,N_689,N_696);
nand U777 (N_777,N_694,N_702);
nand U778 (N_778,N_682,N_662);
nand U779 (N_779,N_714,N_660);
or U780 (N_780,N_738,N_776);
or U781 (N_781,N_735,N_773);
or U782 (N_782,N_745,N_732);
xnor U783 (N_783,N_758,N_753);
and U784 (N_784,N_731,N_748);
xor U785 (N_785,N_755,N_763);
nor U786 (N_786,N_723,N_724);
xnor U787 (N_787,N_757,N_771);
xor U788 (N_788,N_750,N_729);
nor U789 (N_789,N_761,N_768);
or U790 (N_790,N_739,N_759);
xor U791 (N_791,N_767,N_778);
xnor U792 (N_792,N_743,N_751);
and U793 (N_793,N_737,N_742);
and U794 (N_794,N_741,N_730);
or U795 (N_795,N_728,N_721);
nand U796 (N_796,N_774,N_762);
nor U797 (N_797,N_726,N_756);
xor U798 (N_798,N_766,N_725);
and U799 (N_799,N_764,N_736);
and U800 (N_800,N_765,N_749);
nor U801 (N_801,N_744,N_746);
and U802 (N_802,N_733,N_747);
nor U803 (N_803,N_734,N_775);
and U804 (N_804,N_779,N_770);
nand U805 (N_805,N_752,N_772);
xnor U806 (N_806,N_754,N_720);
nand U807 (N_807,N_777,N_740);
nor U808 (N_808,N_760,N_722);
nor U809 (N_809,N_727,N_769);
nand U810 (N_810,N_722,N_766);
or U811 (N_811,N_733,N_751);
nand U812 (N_812,N_744,N_729);
nor U813 (N_813,N_753,N_748);
xor U814 (N_814,N_737,N_723);
or U815 (N_815,N_754,N_721);
and U816 (N_816,N_739,N_778);
xnor U817 (N_817,N_768,N_752);
nor U818 (N_818,N_768,N_751);
xnor U819 (N_819,N_752,N_769);
or U820 (N_820,N_769,N_760);
or U821 (N_821,N_755,N_771);
and U822 (N_822,N_763,N_730);
nand U823 (N_823,N_759,N_767);
xnor U824 (N_824,N_740,N_726);
nor U825 (N_825,N_771,N_753);
xor U826 (N_826,N_758,N_765);
and U827 (N_827,N_722,N_761);
nand U828 (N_828,N_743,N_752);
and U829 (N_829,N_760,N_768);
nor U830 (N_830,N_771,N_728);
and U831 (N_831,N_757,N_747);
or U832 (N_832,N_761,N_758);
xor U833 (N_833,N_764,N_750);
or U834 (N_834,N_768,N_749);
xnor U835 (N_835,N_730,N_775);
nor U836 (N_836,N_726,N_746);
and U837 (N_837,N_723,N_727);
nand U838 (N_838,N_726,N_725);
or U839 (N_839,N_753,N_737);
or U840 (N_840,N_818,N_799);
nor U841 (N_841,N_832,N_780);
nor U842 (N_842,N_794,N_813);
xnor U843 (N_843,N_835,N_812);
and U844 (N_844,N_795,N_807);
nand U845 (N_845,N_788,N_820);
and U846 (N_846,N_808,N_816);
or U847 (N_847,N_836,N_833);
nor U848 (N_848,N_783,N_786);
or U849 (N_849,N_798,N_784);
and U850 (N_850,N_809,N_831);
or U851 (N_851,N_796,N_829);
nor U852 (N_852,N_785,N_810);
nor U853 (N_853,N_793,N_782);
and U854 (N_854,N_811,N_826);
nor U855 (N_855,N_823,N_824);
xnor U856 (N_856,N_815,N_839);
xnor U857 (N_857,N_828,N_792);
nor U858 (N_858,N_817,N_803);
xor U859 (N_859,N_838,N_822);
xor U860 (N_860,N_837,N_814);
or U861 (N_861,N_787,N_827);
nand U862 (N_862,N_821,N_791);
nand U863 (N_863,N_825,N_830);
nand U864 (N_864,N_790,N_819);
nor U865 (N_865,N_781,N_789);
and U866 (N_866,N_797,N_800);
nand U867 (N_867,N_801,N_804);
and U868 (N_868,N_834,N_806);
nor U869 (N_869,N_805,N_802);
and U870 (N_870,N_808,N_819);
nand U871 (N_871,N_823,N_834);
and U872 (N_872,N_821,N_799);
nor U873 (N_873,N_817,N_808);
xnor U874 (N_874,N_809,N_822);
nor U875 (N_875,N_784,N_789);
or U876 (N_876,N_790,N_801);
or U877 (N_877,N_794,N_789);
or U878 (N_878,N_819,N_798);
nor U879 (N_879,N_786,N_801);
nand U880 (N_880,N_810,N_839);
and U881 (N_881,N_822,N_811);
nand U882 (N_882,N_809,N_806);
nand U883 (N_883,N_834,N_788);
nor U884 (N_884,N_803,N_801);
and U885 (N_885,N_801,N_784);
or U886 (N_886,N_785,N_815);
xnor U887 (N_887,N_826,N_788);
xor U888 (N_888,N_833,N_832);
xor U889 (N_889,N_833,N_838);
nand U890 (N_890,N_780,N_837);
nand U891 (N_891,N_789,N_827);
or U892 (N_892,N_811,N_782);
xor U893 (N_893,N_787,N_835);
xor U894 (N_894,N_827,N_813);
and U895 (N_895,N_797,N_796);
or U896 (N_896,N_803,N_837);
nand U897 (N_897,N_812,N_797);
and U898 (N_898,N_839,N_787);
or U899 (N_899,N_808,N_828);
xor U900 (N_900,N_891,N_843);
or U901 (N_901,N_846,N_880);
and U902 (N_902,N_890,N_848);
xnor U903 (N_903,N_898,N_871);
nand U904 (N_904,N_842,N_896);
xor U905 (N_905,N_852,N_867);
or U906 (N_906,N_856,N_894);
xnor U907 (N_907,N_899,N_855);
and U908 (N_908,N_864,N_874);
nor U909 (N_909,N_887,N_859);
nand U910 (N_910,N_892,N_897);
or U911 (N_911,N_876,N_851);
or U912 (N_912,N_878,N_888);
xor U913 (N_913,N_847,N_886);
or U914 (N_914,N_882,N_883);
and U915 (N_915,N_857,N_862);
nand U916 (N_916,N_875,N_879);
and U917 (N_917,N_895,N_870);
nand U918 (N_918,N_869,N_844);
xor U919 (N_919,N_849,N_868);
and U920 (N_920,N_872,N_877);
or U921 (N_921,N_854,N_860);
xor U922 (N_922,N_863,N_889);
xor U923 (N_923,N_845,N_873);
nor U924 (N_924,N_865,N_853);
nor U925 (N_925,N_881,N_850);
and U926 (N_926,N_858,N_840);
and U927 (N_927,N_841,N_884);
or U928 (N_928,N_893,N_885);
nand U929 (N_929,N_866,N_861);
xnor U930 (N_930,N_875,N_868);
nor U931 (N_931,N_841,N_851);
nand U932 (N_932,N_884,N_860);
xor U933 (N_933,N_850,N_895);
xor U934 (N_934,N_860,N_877);
nor U935 (N_935,N_886,N_852);
nand U936 (N_936,N_864,N_855);
and U937 (N_937,N_869,N_872);
or U938 (N_938,N_895,N_884);
xnor U939 (N_939,N_846,N_889);
or U940 (N_940,N_898,N_849);
or U941 (N_941,N_866,N_867);
or U942 (N_942,N_884,N_899);
and U943 (N_943,N_881,N_844);
or U944 (N_944,N_844,N_855);
and U945 (N_945,N_881,N_864);
nor U946 (N_946,N_855,N_871);
nor U947 (N_947,N_845,N_856);
and U948 (N_948,N_863,N_877);
and U949 (N_949,N_852,N_883);
nand U950 (N_950,N_859,N_840);
xor U951 (N_951,N_887,N_874);
nor U952 (N_952,N_853,N_851);
or U953 (N_953,N_852,N_879);
nand U954 (N_954,N_845,N_891);
xnor U955 (N_955,N_899,N_861);
nor U956 (N_956,N_861,N_854);
and U957 (N_957,N_893,N_883);
nand U958 (N_958,N_858,N_842);
xnor U959 (N_959,N_892,N_874);
nand U960 (N_960,N_956,N_935);
nor U961 (N_961,N_912,N_941);
and U962 (N_962,N_922,N_918);
or U963 (N_963,N_959,N_905);
and U964 (N_964,N_958,N_915);
nor U965 (N_965,N_917,N_907);
nor U966 (N_966,N_955,N_927);
or U967 (N_967,N_942,N_951);
xnor U968 (N_968,N_937,N_929);
and U969 (N_969,N_909,N_932);
nor U970 (N_970,N_945,N_930);
nand U971 (N_971,N_924,N_908);
nor U972 (N_972,N_940,N_934);
xor U973 (N_973,N_914,N_903);
and U974 (N_974,N_954,N_950);
or U975 (N_975,N_904,N_900);
nor U976 (N_976,N_939,N_928);
and U977 (N_977,N_901,N_936);
nor U978 (N_978,N_947,N_952);
xor U979 (N_979,N_910,N_919);
and U980 (N_980,N_921,N_933);
nand U981 (N_981,N_902,N_906);
nor U982 (N_982,N_957,N_948);
nor U983 (N_983,N_923,N_911);
nor U984 (N_984,N_943,N_949);
nand U985 (N_985,N_926,N_938);
xor U986 (N_986,N_920,N_925);
nand U987 (N_987,N_913,N_931);
nor U988 (N_988,N_944,N_953);
nor U989 (N_989,N_916,N_946);
nor U990 (N_990,N_914,N_918);
or U991 (N_991,N_910,N_936);
nand U992 (N_992,N_944,N_935);
and U993 (N_993,N_948,N_908);
or U994 (N_994,N_901,N_904);
nand U995 (N_995,N_952,N_912);
or U996 (N_996,N_913,N_925);
nand U997 (N_997,N_913,N_924);
nor U998 (N_998,N_959,N_931);
xnor U999 (N_999,N_916,N_947);
and U1000 (N_1000,N_919,N_925);
or U1001 (N_1001,N_945,N_941);
or U1002 (N_1002,N_946,N_938);
xor U1003 (N_1003,N_921,N_925);
and U1004 (N_1004,N_946,N_931);
and U1005 (N_1005,N_931,N_938);
and U1006 (N_1006,N_906,N_953);
and U1007 (N_1007,N_915,N_941);
nand U1008 (N_1008,N_953,N_957);
or U1009 (N_1009,N_933,N_951);
xor U1010 (N_1010,N_944,N_934);
xnor U1011 (N_1011,N_953,N_919);
xnor U1012 (N_1012,N_940,N_929);
nor U1013 (N_1013,N_918,N_951);
xnor U1014 (N_1014,N_916,N_925);
xnor U1015 (N_1015,N_932,N_903);
or U1016 (N_1016,N_912,N_934);
and U1017 (N_1017,N_903,N_959);
or U1018 (N_1018,N_949,N_920);
xor U1019 (N_1019,N_909,N_953);
nor U1020 (N_1020,N_996,N_1013);
nor U1021 (N_1021,N_1003,N_1004);
nand U1022 (N_1022,N_960,N_1017);
or U1023 (N_1023,N_1015,N_993);
nor U1024 (N_1024,N_962,N_986);
and U1025 (N_1025,N_1014,N_981);
nor U1026 (N_1026,N_1009,N_990);
nor U1027 (N_1027,N_995,N_964);
or U1028 (N_1028,N_983,N_988);
nor U1029 (N_1029,N_963,N_987);
xnor U1030 (N_1030,N_1016,N_971);
and U1031 (N_1031,N_976,N_970);
xnor U1032 (N_1032,N_978,N_1008);
nand U1033 (N_1033,N_966,N_1001);
xor U1034 (N_1034,N_992,N_1007);
or U1035 (N_1035,N_979,N_980);
nand U1036 (N_1036,N_972,N_974);
nand U1037 (N_1037,N_973,N_1012);
and U1038 (N_1038,N_975,N_969);
nand U1039 (N_1039,N_968,N_999);
nor U1040 (N_1040,N_1000,N_1019);
nor U1041 (N_1041,N_1002,N_997);
nand U1042 (N_1042,N_967,N_998);
or U1043 (N_1043,N_965,N_985);
and U1044 (N_1044,N_991,N_1006);
or U1045 (N_1045,N_1018,N_984);
and U1046 (N_1046,N_1011,N_977);
xor U1047 (N_1047,N_1005,N_994);
xnor U1048 (N_1048,N_982,N_1010);
nand U1049 (N_1049,N_961,N_989);
and U1050 (N_1050,N_965,N_962);
xor U1051 (N_1051,N_1008,N_1015);
nand U1052 (N_1052,N_1004,N_1017);
and U1053 (N_1053,N_984,N_1012);
or U1054 (N_1054,N_997,N_993);
nand U1055 (N_1055,N_966,N_1011);
and U1056 (N_1056,N_978,N_997);
or U1057 (N_1057,N_963,N_997);
nor U1058 (N_1058,N_1009,N_995);
or U1059 (N_1059,N_988,N_1016);
xnor U1060 (N_1060,N_964,N_969);
nand U1061 (N_1061,N_1017,N_1016);
xnor U1062 (N_1062,N_990,N_961);
xnor U1063 (N_1063,N_1014,N_1000);
xnor U1064 (N_1064,N_1011,N_961);
or U1065 (N_1065,N_1001,N_1016);
nand U1066 (N_1066,N_974,N_973);
xnor U1067 (N_1067,N_974,N_991);
xor U1068 (N_1068,N_964,N_985);
nand U1069 (N_1069,N_980,N_986);
and U1070 (N_1070,N_1018,N_988);
nor U1071 (N_1071,N_983,N_981);
or U1072 (N_1072,N_1017,N_982);
or U1073 (N_1073,N_979,N_960);
and U1074 (N_1074,N_972,N_1013);
or U1075 (N_1075,N_1019,N_993);
nand U1076 (N_1076,N_960,N_980);
nand U1077 (N_1077,N_991,N_1019);
and U1078 (N_1078,N_1002,N_1005);
or U1079 (N_1079,N_967,N_976);
nor U1080 (N_1080,N_1057,N_1041);
nand U1081 (N_1081,N_1032,N_1037);
or U1082 (N_1082,N_1045,N_1065);
nor U1083 (N_1083,N_1075,N_1072);
nor U1084 (N_1084,N_1020,N_1055);
nand U1085 (N_1085,N_1047,N_1074);
xnor U1086 (N_1086,N_1040,N_1053);
or U1087 (N_1087,N_1073,N_1063);
or U1088 (N_1088,N_1076,N_1054);
xor U1089 (N_1089,N_1077,N_1078);
nor U1090 (N_1090,N_1028,N_1050);
nor U1091 (N_1091,N_1069,N_1033);
nand U1092 (N_1092,N_1070,N_1067);
nand U1093 (N_1093,N_1046,N_1036);
or U1094 (N_1094,N_1060,N_1024);
or U1095 (N_1095,N_1034,N_1030);
nor U1096 (N_1096,N_1052,N_1029);
and U1097 (N_1097,N_1059,N_1027);
nand U1098 (N_1098,N_1038,N_1064);
or U1099 (N_1099,N_1051,N_1026);
xor U1100 (N_1100,N_1071,N_1049);
and U1101 (N_1101,N_1025,N_1079);
xnor U1102 (N_1102,N_1062,N_1035);
nor U1103 (N_1103,N_1068,N_1044);
nand U1104 (N_1104,N_1021,N_1056);
or U1105 (N_1105,N_1022,N_1042);
nor U1106 (N_1106,N_1023,N_1048);
and U1107 (N_1107,N_1031,N_1043);
and U1108 (N_1108,N_1061,N_1066);
xor U1109 (N_1109,N_1039,N_1058);
nand U1110 (N_1110,N_1066,N_1036);
xnor U1111 (N_1111,N_1043,N_1036);
xnor U1112 (N_1112,N_1045,N_1077);
nor U1113 (N_1113,N_1023,N_1052);
nand U1114 (N_1114,N_1078,N_1036);
or U1115 (N_1115,N_1056,N_1066);
or U1116 (N_1116,N_1060,N_1055);
and U1117 (N_1117,N_1031,N_1022);
nor U1118 (N_1118,N_1028,N_1048);
and U1119 (N_1119,N_1033,N_1052);
and U1120 (N_1120,N_1020,N_1036);
or U1121 (N_1121,N_1044,N_1073);
nand U1122 (N_1122,N_1046,N_1067);
nand U1123 (N_1123,N_1078,N_1051);
xnor U1124 (N_1124,N_1058,N_1040);
xor U1125 (N_1125,N_1048,N_1030);
nor U1126 (N_1126,N_1035,N_1036);
xnor U1127 (N_1127,N_1045,N_1059);
nand U1128 (N_1128,N_1041,N_1076);
or U1129 (N_1129,N_1071,N_1038);
nand U1130 (N_1130,N_1074,N_1065);
or U1131 (N_1131,N_1036,N_1061);
xnor U1132 (N_1132,N_1027,N_1023);
nor U1133 (N_1133,N_1024,N_1064);
and U1134 (N_1134,N_1038,N_1051);
nor U1135 (N_1135,N_1044,N_1047);
and U1136 (N_1136,N_1020,N_1073);
and U1137 (N_1137,N_1029,N_1044);
xor U1138 (N_1138,N_1047,N_1050);
nor U1139 (N_1139,N_1063,N_1071);
or U1140 (N_1140,N_1086,N_1113);
and U1141 (N_1141,N_1132,N_1085);
xor U1142 (N_1142,N_1116,N_1124);
nor U1143 (N_1143,N_1100,N_1097);
or U1144 (N_1144,N_1099,N_1117);
nand U1145 (N_1145,N_1121,N_1114);
xnor U1146 (N_1146,N_1093,N_1138);
nand U1147 (N_1147,N_1125,N_1120);
or U1148 (N_1148,N_1105,N_1137);
xnor U1149 (N_1149,N_1104,N_1096);
nand U1150 (N_1150,N_1081,N_1082);
nand U1151 (N_1151,N_1080,N_1091);
xor U1152 (N_1152,N_1106,N_1110);
or U1153 (N_1153,N_1134,N_1128);
nand U1154 (N_1154,N_1090,N_1133);
xnor U1155 (N_1155,N_1098,N_1119);
and U1156 (N_1156,N_1101,N_1136);
nand U1157 (N_1157,N_1108,N_1139);
or U1158 (N_1158,N_1115,N_1109);
nand U1159 (N_1159,N_1088,N_1092);
nor U1160 (N_1160,N_1087,N_1131);
nand U1161 (N_1161,N_1135,N_1095);
xor U1162 (N_1162,N_1122,N_1102);
and U1163 (N_1163,N_1130,N_1112);
nor U1164 (N_1164,N_1126,N_1103);
and U1165 (N_1165,N_1107,N_1111);
nor U1166 (N_1166,N_1089,N_1127);
nand U1167 (N_1167,N_1129,N_1094);
nor U1168 (N_1168,N_1083,N_1118);
and U1169 (N_1169,N_1084,N_1123);
xnor U1170 (N_1170,N_1098,N_1121);
nand U1171 (N_1171,N_1091,N_1083);
or U1172 (N_1172,N_1094,N_1112);
nor U1173 (N_1173,N_1088,N_1115);
nor U1174 (N_1174,N_1114,N_1096);
nand U1175 (N_1175,N_1113,N_1135);
nor U1176 (N_1176,N_1135,N_1122);
xnor U1177 (N_1177,N_1114,N_1134);
or U1178 (N_1178,N_1090,N_1117);
and U1179 (N_1179,N_1137,N_1099);
or U1180 (N_1180,N_1082,N_1131);
nand U1181 (N_1181,N_1118,N_1084);
nand U1182 (N_1182,N_1114,N_1119);
or U1183 (N_1183,N_1114,N_1127);
and U1184 (N_1184,N_1115,N_1132);
nor U1185 (N_1185,N_1098,N_1106);
and U1186 (N_1186,N_1125,N_1119);
and U1187 (N_1187,N_1101,N_1081);
or U1188 (N_1188,N_1092,N_1086);
nor U1189 (N_1189,N_1134,N_1095);
nand U1190 (N_1190,N_1123,N_1086);
or U1191 (N_1191,N_1130,N_1087);
nand U1192 (N_1192,N_1117,N_1103);
nand U1193 (N_1193,N_1104,N_1135);
nand U1194 (N_1194,N_1101,N_1138);
and U1195 (N_1195,N_1116,N_1112);
xor U1196 (N_1196,N_1139,N_1135);
nor U1197 (N_1197,N_1116,N_1134);
nor U1198 (N_1198,N_1080,N_1121);
and U1199 (N_1199,N_1099,N_1103);
nor U1200 (N_1200,N_1196,N_1160);
and U1201 (N_1201,N_1197,N_1154);
or U1202 (N_1202,N_1177,N_1152);
and U1203 (N_1203,N_1140,N_1143);
nor U1204 (N_1204,N_1185,N_1198);
and U1205 (N_1205,N_1195,N_1183);
and U1206 (N_1206,N_1141,N_1189);
and U1207 (N_1207,N_1150,N_1190);
or U1208 (N_1208,N_1168,N_1157);
or U1209 (N_1209,N_1181,N_1176);
xnor U1210 (N_1210,N_1194,N_1171);
xor U1211 (N_1211,N_1170,N_1155);
nand U1212 (N_1212,N_1164,N_1159);
nor U1213 (N_1213,N_1188,N_1158);
nand U1214 (N_1214,N_1175,N_1163);
nand U1215 (N_1215,N_1186,N_1182);
and U1216 (N_1216,N_1142,N_1146);
xor U1217 (N_1217,N_1179,N_1165);
or U1218 (N_1218,N_1145,N_1153);
xnor U1219 (N_1219,N_1172,N_1149);
or U1220 (N_1220,N_1199,N_1192);
nor U1221 (N_1221,N_1147,N_1144);
nand U1222 (N_1222,N_1151,N_1180);
and U1223 (N_1223,N_1162,N_1166);
nand U1224 (N_1224,N_1187,N_1156);
xor U1225 (N_1225,N_1191,N_1178);
or U1226 (N_1226,N_1148,N_1169);
xnor U1227 (N_1227,N_1161,N_1167);
nand U1228 (N_1228,N_1174,N_1193);
xor U1229 (N_1229,N_1173,N_1184);
or U1230 (N_1230,N_1178,N_1165);
and U1231 (N_1231,N_1143,N_1179);
xor U1232 (N_1232,N_1194,N_1175);
xor U1233 (N_1233,N_1193,N_1161);
nand U1234 (N_1234,N_1176,N_1158);
and U1235 (N_1235,N_1147,N_1148);
nor U1236 (N_1236,N_1155,N_1183);
xor U1237 (N_1237,N_1165,N_1160);
or U1238 (N_1238,N_1152,N_1185);
or U1239 (N_1239,N_1183,N_1143);
xnor U1240 (N_1240,N_1146,N_1160);
and U1241 (N_1241,N_1179,N_1164);
xnor U1242 (N_1242,N_1195,N_1147);
xor U1243 (N_1243,N_1191,N_1149);
and U1244 (N_1244,N_1159,N_1186);
or U1245 (N_1245,N_1148,N_1183);
or U1246 (N_1246,N_1146,N_1159);
nand U1247 (N_1247,N_1174,N_1185);
xor U1248 (N_1248,N_1168,N_1185);
or U1249 (N_1249,N_1178,N_1158);
xor U1250 (N_1250,N_1154,N_1152);
xor U1251 (N_1251,N_1156,N_1175);
nand U1252 (N_1252,N_1150,N_1192);
and U1253 (N_1253,N_1163,N_1160);
nor U1254 (N_1254,N_1169,N_1141);
xnor U1255 (N_1255,N_1147,N_1191);
or U1256 (N_1256,N_1172,N_1182);
and U1257 (N_1257,N_1195,N_1141);
xnor U1258 (N_1258,N_1194,N_1163);
nor U1259 (N_1259,N_1161,N_1142);
nor U1260 (N_1260,N_1235,N_1247);
or U1261 (N_1261,N_1248,N_1251);
xor U1262 (N_1262,N_1225,N_1241);
or U1263 (N_1263,N_1217,N_1207);
xnor U1264 (N_1264,N_1219,N_1236);
and U1265 (N_1265,N_1232,N_1237);
nor U1266 (N_1266,N_1202,N_1239);
or U1267 (N_1267,N_1256,N_1246);
nand U1268 (N_1268,N_1212,N_1210);
nor U1269 (N_1269,N_1230,N_1242);
nand U1270 (N_1270,N_1258,N_1206);
xnor U1271 (N_1271,N_1249,N_1254);
nor U1272 (N_1272,N_1250,N_1257);
nand U1273 (N_1273,N_1253,N_1222);
nor U1274 (N_1274,N_1226,N_1234);
and U1275 (N_1275,N_1221,N_1218);
or U1276 (N_1276,N_1203,N_1216);
nor U1277 (N_1277,N_1211,N_1255);
xor U1278 (N_1278,N_1209,N_1240);
nand U1279 (N_1279,N_1205,N_1220);
or U1280 (N_1280,N_1229,N_1223);
nor U1281 (N_1281,N_1233,N_1228);
xor U1282 (N_1282,N_1231,N_1204);
and U1283 (N_1283,N_1252,N_1215);
nor U1284 (N_1284,N_1227,N_1208);
or U1285 (N_1285,N_1243,N_1259);
nor U1286 (N_1286,N_1245,N_1213);
or U1287 (N_1287,N_1201,N_1238);
nor U1288 (N_1288,N_1200,N_1244);
xnor U1289 (N_1289,N_1224,N_1214);
and U1290 (N_1290,N_1242,N_1235);
and U1291 (N_1291,N_1248,N_1212);
or U1292 (N_1292,N_1254,N_1248);
nor U1293 (N_1293,N_1245,N_1208);
xnor U1294 (N_1294,N_1239,N_1208);
or U1295 (N_1295,N_1249,N_1214);
nor U1296 (N_1296,N_1214,N_1259);
or U1297 (N_1297,N_1248,N_1238);
and U1298 (N_1298,N_1251,N_1208);
nand U1299 (N_1299,N_1250,N_1204);
and U1300 (N_1300,N_1223,N_1205);
and U1301 (N_1301,N_1207,N_1210);
xnor U1302 (N_1302,N_1254,N_1238);
or U1303 (N_1303,N_1244,N_1205);
nand U1304 (N_1304,N_1251,N_1239);
nand U1305 (N_1305,N_1232,N_1211);
nor U1306 (N_1306,N_1224,N_1255);
and U1307 (N_1307,N_1201,N_1236);
and U1308 (N_1308,N_1241,N_1223);
or U1309 (N_1309,N_1225,N_1200);
nand U1310 (N_1310,N_1215,N_1225);
nor U1311 (N_1311,N_1230,N_1202);
nor U1312 (N_1312,N_1203,N_1226);
and U1313 (N_1313,N_1229,N_1255);
nor U1314 (N_1314,N_1230,N_1212);
nor U1315 (N_1315,N_1204,N_1222);
and U1316 (N_1316,N_1200,N_1217);
xnor U1317 (N_1317,N_1229,N_1222);
nand U1318 (N_1318,N_1200,N_1245);
nor U1319 (N_1319,N_1220,N_1209);
xnor U1320 (N_1320,N_1278,N_1312);
xnor U1321 (N_1321,N_1268,N_1280);
nor U1322 (N_1322,N_1304,N_1262);
and U1323 (N_1323,N_1305,N_1292);
nor U1324 (N_1324,N_1298,N_1296);
xnor U1325 (N_1325,N_1274,N_1301);
or U1326 (N_1326,N_1270,N_1302);
xor U1327 (N_1327,N_1295,N_1291);
nor U1328 (N_1328,N_1311,N_1273);
nor U1329 (N_1329,N_1264,N_1285);
xnor U1330 (N_1330,N_1286,N_1315);
nor U1331 (N_1331,N_1277,N_1299);
or U1332 (N_1332,N_1290,N_1263);
xnor U1333 (N_1333,N_1306,N_1281);
nor U1334 (N_1334,N_1282,N_1272);
or U1335 (N_1335,N_1293,N_1269);
nor U1336 (N_1336,N_1318,N_1307);
nand U1337 (N_1337,N_1309,N_1271);
xor U1338 (N_1338,N_1317,N_1316);
nor U1339 (N_1339,N_1310,N_1303);
nand U1340 (N_1340,N_1294,N_1279);
nand U1341 (N_1341,N_1260,N_1267);
and U1342 (N_1342,N_1288,N_1275);
nand U1343 (N_1343,N_1308,N_1300);
nand U1344 (N_1344,N_1297,N_1276);
nand U1345 (N_1345,N_1266,N_1283);
or U1346 (N_1346,N_1265,N_1313);
xnor U1347 (N_1347,N_1284,N_1289);
nor U1348 (N_1348,N_1261,N_1319);
xnor U1349 (N_1349,N_1314,N_1287);
nand U1350 (N_1350,N_1295,N_1283);
nand U1351 (N_1351,N_1284,N_1297);
and U1352 (N_1352,N_1280,N_1290);
and U1353 (N_1353,N_1261,N_1297);
nand U1354 (N_1354,N_1287,N_1312);
or U1355 (N_1355,N_1316,N_1290);
nand U1356 (N_1356,N_1292,N_1303);
and U1357 (N_1357,N_1272,N_1267);
and U1358 (N_1358,N_1268,N_1290);
nand U1359 (N_1359,N_1309,N_1287);
nor U1360 (N_1360,N_1261,N_1260);
nand U1361 (N_1361,N_1260,N_1289);
xor U1362 (N_1362,N_1316,N_1273);
nor U1363 (N_1363,N_1305,N_1289);
or U1364 (N_1364,N_1291,N_1287);
nand U1365 (N_1365,N_1282,N_1293);
or U1366 (N_1366,N_1279,N_1311);
nor U1367 (N_1367,N_1272,N_1301);
nand U1368 (N_1368,N_1316,N_1294);
nand U1369 (N_1369,N_1306,N_1308);
and U1370 (N_1370,N_1262,N_1300);
or U1371 (N_1371,N_1272,N_1274);
xnor U1372 (N_1372,N_1273,N_1266);
or U1373 (N_1373,N_1274,N_1319);
and U1374 (N_1374,N_1318,N_1278);
nand U1375 (N_1375,N_1284,N_1281);
xnor U1376 (N_1376,N_1279,N_1293);
and U1377 (N_1377,N_1303,N_1279);
nand U1378 (N_1378,N_1269,N_1317);
and U1379 (N_1379,N_1283,N_1285);
or U1380 (N_1380,N_1353,N_1359);
and U1381 (N_1381,N_1320,N_1335);
nor U1382 (N_1382,N_1352,N_1337);
and U1383 (N_1383,N_1366,N_1341);
nand U1384 (N_1384,N_1345,N_1378);
xnor U1385 (N_1385,N_1338,N_1375);
nand U1386 (N_1386,N_1334,N_1365);
or U1387 (N_1387,N_1324,N_1351);
or U1388 (N_1388,N_1356,N_1323);
xnor U1389 (N_1389,N_1362,N_1371);
nand U1390 (N_1390,N_1330,N_1343);
or U1391 (N_1391,N_1364,N_1361);
nor U1392 (N_1392,N_1358,N_1369);
and U1393 (N_1393,N_1350,N_1344);
nand U1394 (N_1394,N_1340,N_1348);
or U1395 (N_1395,N_1367,N_1325);
nand U1396 (N_1396,N_1372,N_1327);
and U1397 (N_1397,N_1347,N_1376);
nor U1398 (N_1398,N_1355,N_1336);
nand U1399 (N_1399,N_1377,N_1363);
xnor U1400 (N_1400,N_1373,N_1328);
and U1401 (N_1401,N_1332,N_1379);
nand U1402 (N_1402,N_1321,N_1322);
and U1403 (N_1403,N_1326,N_1374);
nand U1404 (N_1404,N_1360,N_1357);
nor U1405 (N_1405,N_1368,N_1339);
nor U1406 (N_1406,N_1329,N_1333);
or U1407 (N_1407,N_1370,N_1342);
or U1408 (N_1408,N_1349,N_1354);
or U1409 (N_1409,N_1346,N_1331);
nor U1410 (N_1410,N_1339,N_1332);
nand U1411 (N_1411,N_1364,N_1350);
or U1412 (N_1412,N_1330,N_1366);
xnor U1413 (N_1413,N_1359,N_1333);
xor U1414 (N_1414,N_1365,N_1341);
nor U1415 (N_1415,N_1341,N_1356);
nand U1416 (N_1416,N_1338,N_1328);
nor U1417 (N_1417,N_1336,N_1333);
xnor U1418 (N_1418,N_1360,N_1375);
nor U1419 (N_1419,N_1373,N_1325);
and U1420 (N_1420,N_1378,N_1357);
nor U1421 (N_1421,N_1368,N_1370);
nor U1422 (N_1422,N_1344,N_1359);
and U1423 (N_1423,N_1337,N_1365);
or U1424 (N_1424,N_1332,N_1357);
or U1425 (N_1425,N_1356,N_1368);
xnor U1426 (N_1426,N_1335,N_1378);
or U1427 (N_1427,N_1376,N_1369);
xor U1428 (N_1428,N_1328,N_1378);
or U1429 (N_1429,N_1325,N_1375);
nand U1430 (N_1430,N_1379,N_1351);
or U1431 (N_1431,N_1354,N_1320);
nand U1432 (N_1432,N_1370,N_1322);
and U1433 (N_1433,N_1353,N_1327);
xnor U1434 (N_1434,N_1373,N_1341);
or U1435 (N_1435,N_1320,N_1326);
nand U1436 (N_1436,N_1323,N_1336);
nand U1437 (N_1437,N_1353,N_1326);
and U1438 (N_1438,N_1346,N_1329);
xnor U1439 (N_1439,N_1338,N_1364);
nand U1440 (N_1440,N_1399,N_1409);
xor U1441 (N_1441,N_1404,N_1390);
or U1442 (N_1442,N_1436,N_1406);
and U1443 (N_1443,N_1417,N_1432);
nor U1444 (N_1444,N_1414,N_1425);
or U1445 (N_1445,N_1385,N_1388);
nand U1446 (N_1446,N_1437,N_1391);
and U1447 (N_1447,N_1395,N_1383);
and U1448 (N_1448,N_1387,N_1415);
nand U1449 (N_1449,N_1396,N_1410);
or U1450 (N_1450,N_1398,N_1434);
nand U1451 (N_1451,N_1403,N_1424);
xor U1452 (N_1452,N_1400,N_1426);
or U1453 (N_1453,N_1382,N_1429);
nor U1454 (N_1454,N_1380,N_1439);
and U1455 (N_1455,N_1427,N_1405);
and U1456 (N_1456,N_1418,N_1419);
nand U1457 (N_1457,N_1416,N_1421);
xor U1458 (N_1458,N_1423,N_1411);
xor U1459 (N_1459,N_1407,N_1420);
or U1460 (N_1460,N_1389,N_1392);
nor U1461 (N_1461,N_1428,N_1384);
or U1462 (N_1462,N_1438,N_1393);
nor U1463 (N_1463,N_1381,N_1435);
nand U1464 (N_1464,N_1412,N_1413);
nand U1465 (N_1465,N_1408,N_1431);
nor U1466 (N_1466,N_1397,N_1430);
nor U1467 (N_1467,N_1386,N_1433);
or U1468 (N_1468,N_1402,N_1401);
or U1469 (N_1469,N_1422,N_1394);
or U1470 (N_1470,N_1414,N_1413);
xnor U1471 (N_1471,N_1395,N_1414);
and U1472 (N_1472,N_1433,N_1397);
nor U1473 (N_1473,N_1412,N_1421);
and U1474 (N_1474,N_1432,N_1431);
and U1475 (N_1475,N_1426,N_1427);
nand U1476 (N_1476,N_1419,N_1397);
and U1477 (N_1477,N_1432,N_1403);
xor U1478 (N_1478,N_1425,N_1384);
nand U1479 (N_1479,N_1411,N_1421);
nand U1480 (N_1480,N_1423,N_1385);
nand U1481 (N_1481,N_1432,N_1427);
nor U1482 (N_1482,N_1419,N_1439);
xnor U1483 (N_1483,N_1398,N_1394);
or U1484 (N_1484,N_1427,N_1415);
xnor U1485 (N_1485,N_1424,N_1397);
xnor U1486 (N_1486,N_1390,N_1431);
or U1487 (N_1487,N_1418,N_1405);
nand U1488 (N_1488,N_1381,N_1389);
nand U1489 (N_1489,N_1393,N_1394);
nor U1490 (N_1490,N_1431,N_1392);
nor U1491 (N_1491,N_1381,N_1412);
xor U1492 (N_1492,N_1432,N_1430);
nand U1493 (N_1493,N_1411,N_1392);
xnor U1494 (N_1494,N_1413,N_1400);
xnor U1495 (N_1495,N_1437,N_1431);
xnor U1496 (N_1496,N_1410,N_1404);
and U1497 (N_1497,N_1405,N_1399);
nand U1498 (N_1498,N_1396,N_1427);
nand U1499 (N_1499,N_1414,N_1415);
and U1500 (N_1500,N_1462,N_1485);
nor U1501 (N_1501,N_1468,N_1451);
nand U1502 (N_1502,N_1498,N_1489);
or U1503 (N_1503,N_1461,N_1452);
xnor U1504 (N_1504,N_1447,N_1490);
and U1505 (N_1505,N_1497,N_1494);
or U1506 (N_1506,N_1467,N_1495);
and U1507 (N_1507,N_1464,N_1458);
nor U1508 (N_1508,N_1472,N_1486);
xor U1509 (N_1509,N_1460,N_1499);
nand U1510 (N_1510,N_1454,N_1459);
xor U1511 (N_1511,N_1474,N_1475);
xor U1512 (N_1512,N_1483,N_1477);
nand U1513 (N_1513,N_1450,N_1479);
xnor U1514 (N_1514,N_1482,N_1442);
or U1515 (N_1515,N_1492,N_1473);
xnor U1516 (N_1516,N_1441,N_1481);
or U1517 (N_1517,N_1470,N_1440);
nand U1518 (N_1518,N_1463,N_1456);
nor U1519 (N_1519,N_1444,N_1448);
nor U1520 (N_1520,N_1493,N_1466);
nand U1521 (N_1521,N_1478,N_1455);
xor U1522 (N_1522,N_1471,N_1443);
and U1523 (N_1523,N_1465,N_1496);
or U1524 (N_1524,N_1487,N_1446);
and U1525 (N_1525,N_1480,N_1453);
xor U1526 (N_1526,N_1476,N_1484);
and U1527 (N_1527,N_1491,N_1445);
nor U1528 (N_1528,N_1449,N_1488);
xor U1529 (N_1529,N_1457,N_1469);
nand U1530 (N_1530,N_1447,N_1468);
or U1531 (N_1531,N_1485,N_1475);
nand U1532 (N_1532,N_1497,N_1498);
or U1533 (N_1533,N_1452,N_1472);
or U1534 (N_1534,N_1459,N_1497);
or U1535 (N_1535,N_1477,N_1459);
or U1536 (N_1536,N_1456,N_1441);
nand U1537 (N_1537,N_1489,N_1448);
or U1538 (N_1538,N_1496,N_1487);
nor U1539 (N_1539,N_1485,N_1486);
or U1540 (N_1540,N_1458,N_1443);
nand U1541 (N_1541,N_1452,N_1469);
nand U1542 (N_1542,N_1466,N_1447);
xor U1543 (N_1543,N_1474,N_1463);
xor U1544 (N_1544,N_1496,N_1488);
nand U1545 (N_1545,N_1471,N_1493);
nand U1546 (N_1546,N_1477,N_1450);
and U1547 (N_1547,N_1494,N_1476);
and U1548 (N_1548,N_1494,N_1464);
and U1549 (N_1549,N_1476,N_1479);
or U1550 (N_1550,N_1481,N_1453);
nand U1551 (N_1551,N_1460,N_1488);
nor U1552 (N_1552,N_1452,N_1499);
or U1553 (N_1553,N_1474,N_1460);
nand U1554 (N_1554,N_1486,N_1454);
xor U1555 (N_1555,N_1492,N_1476);
or U1556 (N_1556,N_1486,N_1460);
and U1557 (N_1557,N_1496,N_1476);
nand U1558 (N_1558,N_1477,N_1447);
nand U1559 (N_1559,N_1442,N_1493);
nand U1560 (N_1560,N_1551,N_1530);
or U1561 (N_1561,N_1534,N_1540);
xor U1562 (N_1562,N_1531,N_1529);
nand U1563 (N_1563,N_1546,N_1544);
and U1564 (N_1564,N_1518,N_1536);
nor U1565 (N_1565,N_1513,N_1558);
nor U1566 (N_1566,N_1538,N_1510);
and U1567 (N_1567,N_1528,N_1515);
xnor U1568 (N_1568,N_1549,N_1541);
nor U1569 (N_1569,N_1508,N_1537);
nand U1570 (N_1570,N_1535,N_1547);
and U1571 (N_1571,N_1505,N_1527);
or U1572 (N_1572,N_1501,N_1502);
or U1573 (N_1573,N_1503,N_1526);
xor U1574 (N_1574,N_1552,N_1517);
or U1575 (N_1575,N_1553,N_1504);
and U1576 (N_1576,N_1523,N_1532);
xor U1577 (N_1577,N_1557,N_1507);
nand U1578 (N_1578,N_1525,N_1539);
nand U1579 (N_1579,N_1548,N_1555);
or U1580 (N_1580,N_1500,N_1550);
or U1581 (N_1581,N_1516,N_1554);
nand U1582 (N_1582,N_1519,N_1522);
xnor U1583 (N_1583,N_1543,N_1559);
and U1584 (N_1584,N_1520,N_1509);
nor U1585 (N_1585,N_1524,N_1545);
or U1586 (N_1586,N_1511,N_1533);
nand U1587 (N_1587,N_1542,N_1512);
or U1588 (N_1588,N_1514,N_1506);
and U1589 (N_1589,N_1556,N_1521);
or U1590 (N_1590,N_1535,N_1558);
or U1591 (N_1591,N_1548,N_1557);
nand U1592 (N_1592,N_1515,N_1509);
nand U1593 (N_1593,N_1544,N_1520);
xnor U1594 (N_1594,N_1526,N_1539);
and U1595 (N_1595,N_1519,N_1510);
xnor U1596 (N_1596,N_1557,N_1533);
nor U1597 (N_1597,N_1554,N_1537);
nand U1598 (N_1598,N_1507,N_1520);
and U1599 (N_1599,N_1526,N_1524);
and U1600 (N_1600,N_1557,N_1550);
or U1601 (N_1601,N_1511,N_1521);
nand U1602 (N_1602,N_1534,N_1511);
nor U1603 (N_1603,N_1537,N_1507);
and U1604 (N_1604,N_1502,N_1505);
nor U1605 (N_1605,N_1508,N_1510);
nor U1606 (N_1606,N_1545,N_1534);
and U1607 (N_1607,N_1513,N_1511);
nand U1608 (N_1608,N_1535,N_1516);
nand U1609 (N_1609,N_1510,N_1517);
nand U1610 (N_1610,N_1539,N_1500);
nand U1611 (N_1611,N_1518,N_1526);
nand U1612 (N_1612,N_1543,N_1552);
or U1613 (N_1613,N_1542,N_1522);
and U1614 (N_1614,N_1532,N_1535);
or U1615 (N_1615,N_1558,N_1534);
xor U1616 (N_1616,N_1504,N_1515);
nor U1617 (N_1617,N_1529,N_1508);
and U1618 (N_1618,N_1523,N_1540);
xnor U1619 (N_1619,N_1526,N_1512);
nor U1620 (N_1620,N_1564,N_1581);
and U1621 (N_1621,N_1570,N_1591);
nand U1622 (N_1622,N_1563,N_1586);
and U1623 (N_1623,N_1560,N_1585);
nand U1624 (N_1624,N_1616,N_1610);
nor U1625 (N_1625,N_1587,N_1598);
xnor U1626 (N_1626,N_1588,N_1583);
xnor U1627 (N_1627,N_1568,N_1597);
xor U1628 (N_1628,N_1571,N_1601);
nand U1629 (N_1629,N_1599,N_1602);
and U1630 (N_1630,N_1606,N_1590);
nor U1631 (N_1631,N_1592,N_1608);
or U1632 (N_1632,N_1607,N_1589);
and U1633 (N_1633,N_1566,N_1613);
nand U1634 (N_1634,N_1578,N_1582);
and U1635 (N_1635,N_1596,N_1577);
nand U1636 (N_1636,N_1605,N_1600);
and U1637 (N_1637,N_1561,N_1567);
nand U1638 (N_1638,N_1593,N_1580);
nor U1639 (N_1639,N_1574,N_1619);
and U1640 (N_1640,N_1584,N_1611);
xor U1641 (N_1641,N_1562,N_1617);
or U1642 (N_1642,N_1604,N_1603);
xor U1643 (N_1643,N_1565,N_1569);
or U1644 (N_1644,N_1575,N_1594);
or U1645 (N_1645,N_1573,N_1614);
or U1646 (N_1646,N_1576,N_1615);
and U1647 (N_1647,N_1609,N_1572);
nor U1648 (N_1648,N_1612,N_1595);
or U1649 (N_1649,N_1579,N_1618);
nand U1650 (N_1650,N_1595,N_1563);
nor U1651 (N_1651,N_1605,N_1575);
xnor U1652 (N_1652,N_1614,N_1599);
nand U1653 (N_1653,N_1611,N_1613);
and U1654 (N_1654,N_1590,N_1592);
nor U1655 (N_1655,N_1601,N_1596);
or U1656 (N_1656,N_1581,N_1597);
nand U1657 (N_1657,N_1590,N_1610);
nand U1658 (N_1658,N_1604,N_1586);
nor U1659 (N_1659,N_1576,N_1565);
nand U1660 (N_1660,N_1599,N_1571);
nand U1661 (N_1661,N_1572,N_1577);
nor U1662 (N_1662,N_1606,N_1580);
xnor U1663 (N_1663,N_1604,N_1569);
xor U1664 (N_1664,N_1609,N_1602);
or U1665 (N_1665,N_1604,N_1576);
nand U1666 (N_1666,N_1582,N_1567);
nand U1667 (N_1667,N_1617,N_1595);
nand U1668 (N_1668,N_1595,N_1590);
xor U1669 (N_1669,N_1612,N_1570);
xor U1670 (N_1670,N_1571,N_1586);
nand U1671 (N_1671,N_1573,N_1581);
nand U1672 (N_1672,N_1598,N_1571);
and U1673 (N_1673,N_1592,N_1570);
nor U1674 (N_1674,N_1566,N_1602);
xor U1675 (N_1675,N_1584,N_1600);
or U1676 (N_1676,N_1576,N_1594);
nor U1677 (N_1677,N_1598,N_1565);
nand U1678 (N_1678,N_1594,N_1583);
nor U1679 (N_1679,N_1578,N_1590);
and U1680 (N_1680,N_1659,N_1641);
nor U1681 (N_1681,N_1623,N_1630);
nor U1682 (N_1682,N_1661,N_1670);
and U1683 (N_1683,N_1663,N_1674);
xor U1684 (N_1684,N_1666,N_1648);
and U1685 (N_1685,N_1636,N_1632);
or U1686 (N_1686,N_1676,N_1643);
nor U1687 (N_1687,N_1667,N_1622);
xor U1688 (N_1688,N_1631,N_1627);
nor U1689 (N_1689,N_1678,N_1654);
nand U1690 (N_1690,N_1635,N_1634);
or U1691 (N_1691,N_1660,N_1633);
nor U1692 (N_1692,N_1644,N_1665);
and U1693 (N_1693,N_1620,N_1649);
nor U1694 (N_1694,N_1642,N_1668);
xor U1695 (N_1695,N_1647,N_1646);
nand U1696 (N_1696,N_1662,N_1645);
or U1697 (N_1697,N_1679,N_1638);
or U1698 (N_1698,N_1640,N_1655);
nand U1699 (N_1699,N_1637,N_1652);
nand U1700 (N_1700,N_1664,N_1673);
xnor U1701 (N_1701,N_1672,N_1624);
nor U1702 (N_1702,N_1625,N_1675);
nand U1703 (N_1703,N_1669,N_1671);
nand U1704 (N_1704,N_1650,N_1626);
and U1705 (N_1705,N_1658,N_1621);
xor U1706 (N_1706,N_1628,N_1639);
xnor U1707 (N_1707,N_1651,N_1656);
xor U1708 (N_1708,N_1677,N_1629);
nand U1709 (N_1709,N_1657,N_1653);
nand U1710 (N_1710,N_1625,N_1635);
and U1711 (N_1711,N_1640,N_1674);
nand U1712 (N_1712,N_1632,N_1635);
nand U1713 (N_1713,N_1641,N_1627);
nand U1714 (N_1714,N_1658,N_1626);
xor U1715 (N_1715,N_1665,N_1651);
and U1716 (N_1716,N_1643,N_1667);
nand U1717 (N_1717,N_1654,N_1642);
or U1718 (N_1718,N_1662,N_1658);
xor U1719 (N_1719,N_1677,N_1626);
or U1720 (N_1720,N_1646,N_1667);
nand U1721 (N_1721,N_1644,N_1625);
and U1722 (N_1722,N_1672,N_1644);
nand U1723 (N_1723,N_1640,N_1641);
nand U1724 (N_1724,N_1633,N_1627);
and U1725 (N_1725,N_1625,N_1645);
xor U1726 (N_1726,N_1621,N_1625);
nand U1727 (N_1727,N_1641,N_1652);
xnor U1728 (N_1728,N_1631,N_1637);
xor U1729 (N_1729,N_1648,N_1632);
and U1730 (N_1730,N_1651,N_1622);
and U1731 (N_1731,N_1662,N_1641);
xor U1732 (N_1732,N_1631,N_1676);
or U1733 (N_1733,N_1637,N_1646);
and U1734 (N_1734,N_1669,N_1626);
and U1735 (N_1735,N_1670,N_1625);
or U1736 (N_1736,N_1652,N_1639);
nand U1737 (N_1737,N_1638,N_1634);
xor U1738 (N_1738,N_1626,N_1670);
nand U1739 (N_1739,N_1656,N_1675);
and U1740 (N_1740,N_1704,N_1700);
nor U1741 (N_1741,N_1681,N_1730);
nor U1742 (N_1742,N_1702,N_1709);
and U1743 (N_1743,N_1697,N_1715);
xor U1744 (N_1744,N_1680,N_1693);
nand U1745 (N_1745,N_1687,N_1694);
and U1746 (N_1746,N_1705,N_1729);
and U1747 (N_1747,N_1722,N_1708);
and U1748 (N_1748,N_1707,N_1720);
or U1749 (N_1749,N_1684,N_1734);
nor U1750 (N_1750,N_1686,N_1739);
and U1751 (N_1751,N_1690,N_1692);
nand U1752 (N_1752,N_1685,N_1717);
nor U1753 (N_1753,N_1726,N_1696);
nand U1754 (N_1754,N_1723,N_1716);
xor U1755 (N_1755,N_1711,N_1719);
xor U1756 (N_1756,N_1727,N_1732);
xor U1757 (N_1757,N_1703,N_1695);
nor U1758 (N_1758,N_1688,N_1735);
nor U1759 (N_1759,N_1698,N_1736);
and U1760 (N_1760,N_1689,N_1714);
or U1761 (N_1761,N_1713,N_1718);
or U1762 (N_1762,N_1710,N_1731);
or U1763 (N_1763,N_1733,N_1682);
or U1764 (N_1764,N_1724,N_1683);
and U1765 (N_1765,N_1699,N_1738);
or U1766 (N_1766,N_1706,N_1712);
and U1767 (N_1767,N_1691,N_1725);
or U1768 (N_1768,N_1701,N_1737);
nor U1769 (N_1769,N_1721,N_1728);
and U1770 (N_1770,N_1706,N_1700);
nand U1771 (N_1771,N_1692,N_1702);
nand U1772 (N_1772,N_1707,N_1708);
xnor U1773 (N_1773,N_1728,N_1716);
xnor U1774 (N_1774,N_1720,N_1716);
nand U1775 (N_1775,N_1691,N_1721);
and U1776 (N_1776,N_1710,N_1724);
nand U1777 (N_1777,N_1722,N_1717);
nand U1778 (N_1778,N_1723,N_1707);
nand U1779 (N_1779,N_1686,N_1719);
xnor U1780 (N_1780,N_1704,N_1737);
and U1781 (N_1781,N_1735,N_1720);
and U1782 (N_1782,N_1731,N_1713);
nand U1783 (N_1783,N_1699,N_1715);
and U1784 (N_1784,N_1731,N_1735);
nand U1785 (N_1785,N_1730,N_1689);
nand U1786 (N_1786,N_1739,N_1680);
xor U1787 (N_1787,N_1694,N_1709);
or U1788 (N_1788,N_1737,N_1680);
or U1789 (N_1789,N_1726,N_1736);
nor U1790 (N_1790,N_1735,N_1718);
nor U1791 (N_1791,N_1706,N_1695);
nand U1792 (N_1792,N_1681,N_1698);
xnor U1793 (N_1793,N_1720,N_1715);
xnor U1794 (N_1794,N_1700,N_1715);
nand U1795 (N_1795,N_1726,N_1702);
or U1796 (N_1796,N_1698,N_1680);
or U1797 (N_1797,N_1731,N_1719);
and U1798 (N_1798,N_1689,N_1700);
nand U1799 (N_1799,N_1729,N_1688);
and U1800 (N_1800,N_1799,N_1746);
nor U1801 (N_1801,N_1747,N_1749);
or U1802 (N_1802,N_1753,N_1789);
and U1803 (N_1803,N_1754,N_1767);
nand U1804 (N_1804,N_1773,N_1796);
nor U1805 (N_1805,N_1795,N_1775);
xnor U1806 (N_1806,N_1762,N_1771);
or U1807 (N_1807,N_1752,N_1745);
and U1808 (N_1808,N_1742,N_1755);
nand U1809 (N_1809,N_1778,N_1788);
nor U1810 (N_1810,N_1768,N_1751);
nand U1811 (N_1811,N_1783,N_1759);
nand U1812 (N_1812,N_1791,N_1740);
xnor U1813 (N_1813,N_1794,N_1793);
xor U1814 (N_1814,N_1756,N_1777);
nor U1815 (N_1815,N_1763,N_1779);
xor U1816 (N_1816,N_1782,N_1741);
xnor U1817 (N_1817,N_1781,N_1743);
nand U1818 (N_1818,N_1744,N_1792);
xnor U1819 (N_1819,N_1758,N_1780);
nor U1820 (N_1820,N_1765,N_1785);
xor U1821 (N_1821,N_1766,N_1757);
xnor U1822 (N_1822,N_1750,N_1772);
and U1823 (N_1823,N_1776,N_1797);
or U1824 (N_1824,N_1769,N_1760);
nand U1825 (N_1825,N_1748,N_1774);
nand U1826 (N_1826,N_1784,N_1761);
or U1827 (N_1827,N_1790,N_1798);
or U1828 (N_1828,N_1786,N_1787);
and U1829 (N_1829,N_1764,N_1770);
nor U1830 (N_1830,N_1763,N_1756);
xor U1831 (N_1831,N_1747,N_1744);
xor U1832 (N_1832,N_1780,N_1744);
xnor U1833 (N_1833,N_1754,N_1795);
xor U1834 (N_1834,N_1767,N_1760);
or U1835 (N_1835,N_1795,N_1770);
nand U1836 (N_1836,N_1765,N_1761);
and U1837 (N_1837,N_1780,N_1784);
nand U1838 (N_1838,N_1789,N_1791);
nand U1839 (N_1839,N_1743,N_1770);
nand U1840 (N_1840,N_1762,N_1748);
nor U1841 (N_1841,N_1744,N_1746);
xnor U1842 (N_1842,N_1763,N_1767);
or U1843 (N_1843,N_1772,N_1777);
xor U1844 (N_1844,N_1766,N_1759);
nor U1845 (N_1845,N_1743,N_1750);
or U1846 (N_1846,N_1788,N_1774);
nand U1847 (N_1847,N_1754,N_1759);
nor U1848 (N_1848,N_1777,N_1768);
nor U1849 (N_1849,N_1797,N_1742);
nand U1850 (N_1850,N_1764,N_1743);
nor U1851 (N_1851,N_1764,N_1772);
nor U1852 (N_1852,N_1740,N_1779);
or U1853 (N_1853,N_1782,N_1790);
nand U1854 (N_1854,N_1789,N_1765);
or U1855 (N_1855,N_1790,N_1749);
nand U1856 (N_1856,N_1795,N_1783);
nand U1857 (N_1857,N_1752,N_1787);
or U1858 (N_1858,N_1761,N_1746);
nand U1859 (N_1859,N_1741,N_1762);
and U1860 (N_1860,N_1819,N_1837);
and U1861 (N_1861,N_1815,N_1808);
nor U1862 (N_1862,N_1814,N_1848);
and U1863 (N_1863,N_1852,N_1801);
nor U1864 (N_1864,N_1825,N_1824);
xor U1865 (N_1865,N_1818,N_1817);
nor U1866 (N_1866,N_1847,N_1813);
xnor U1867 (N_1867,N_1840,N_1849);
nand U1868 (N_1868,N_1846,N_1839);
or U1869 (N_1869,N_1844,N_1811);
xnor U1870 (N_1870,N_1800,N_1802);
or U1871 (N_1871,N_1831,N_1855);
nand U1872 (N_1872,N_1810,N_1838);
nand U1873 (N_1873,N_1816,N_1842);
and U1874 (N_1874,N_1828,N_1820);
and U1875 (N_1875,N_1805,N_1850);
nand U1876 (N_1876,N_1834,N_1841);
and U1877 (N_1877,N_1836,N_1803);
or U1878 (N_1878,N_1827,N_1821);
nor U1879 (N_1879,N_1857,N_1829);
nand U1880 (N_1880,N_1854,N_1826);
and U1881 (N_1881,N_1807,N_1804);
xnor U1882 (N_1882,N_1812,N_1832);
or U1883 (N_1883,N_1822,N_1823);
or U1884 (N_1884,N_1853,N_1859);
and U1885 (N_1885,N_1835,N_1845);
nor U1886 (N_1886,N_1856,N_1809);
xnor U1887 (N_1887,N_1830,N_1858);
nor U1888 (N_1888,N_1833,N_1851);
or U1889 (N_1889,N_1843,N_1806);
and U1890 (N_1890,N_1851,N_1826);
xor U1891 (N_1891,N_1844,N_1829);
xnor U1892 (N_1892,N_1853,N_1818);
or U1893 (N_1893,N_1819,N_1807);
and U1894 (N_1894,N_1843,N_1811);
and U1895 (N_1895,N_1809,N_1831);
nor U1896 (N_1896,N_1848,N_1805);
nand U1897 (N_1897,N_1843,N_1849);
and U1898 (N_1898,N_1838,N_1833);
nor U1899 (N_1899,N_1814,N_1855);
nor U1900 (N_1900,N_1821,N_1824);
and U1901 (N_1901,N_1836,N_1854);
xor U1902 (N_1902,N_1830,N_1838);
and U1903 (N_1903,N_1834,N_1825);
and U1904 (N_1904,N_1822,N_1800);
xor U1905 (N_1905,N_1804,N_1821);
nor U1906 (N_1906,N_1845,N_1834);
nand U1907 (N_1907,N_1836,N_1832);
and U1908 (N_1908,N_1830,N_1850);
nor U1909 (N_1909,N_1812,N_1856);
nor U1910 (N_1910,N_1814,N_1836);
or U1911 (N_1911,N_1818,N_1823);
nand U1912 (N_1912,N_1843,N_1808);
nor U1913 (N_1913,N_1842,N_1834);
or U1914 (N_1914,N_1836,N_1825);
nand U1915 (N_1915,N_1842,N_1814);
or U1916 (N_1916,N_1803,N_1802);
nor U1917 (N_1917,N_1854,N_1835);
nand U1918 (N_1918,N_1840,N_1827);
nor U1919 (N_1919,N_1856,N_1849);
or U1920 (N_1920,N_1915,N_1916);
nor U1921 (N_1921,N_1886,N_1897);
nor U1922 (N_1922,N_1878,N_1903);
nand U1923 (N_1923,N_1873,N_1872);
nand U1924 (N_1924,N_1895,N_1876);
or U1925 (N_1925,N_1871,N_1866);
nand U1926 (N_1926,N_1906,N_1912);
nor U1927 (N_1927,N_1887,N_1870);
nand U1928 (N_1928,N_1904,N_1891);
nand U1929 (N_1929,N_1918,N_1874);
nand U1930 (N_1930,N_1884,N_1900);
and U1931 (N_1931,N_1883,N_1864);
and U1932 (N_1932,N_1889,N_1894);
nand U1933 (N_1933,N_1902,N_1898);
nor U1934 (N_1934,N_1893,N_1888);
nor U1935 (N_1935,N_1917,N_1905);
or U1936 (N_1936,N_1919,N_1860);
nand U1937 (N_1937,N_1892,N_1901);
and U1938 (N_1938,N_1861,N_1863);
xor U1939 (N_1939,N_1877,N_1862);
or U1940 (N_1940,N_1882,N_1867);
and U1941 (N_1941,N_1911,N_1913);
xor U1942 (N_1942,N_1907,N_1865);
nand U1943 (N_1943,N_1910,N_1868);
nor U1944 (N_1944,N_1869,N_1880);
nor U1945 (N_1945,N_1890,N_1881);
nand U1946 (N_1946,N_1879,N_1885);
nand U1947 (N_1947,N_1875,N_1914);
nand U1948 (N_1948,N_1899,N_1896);
and U1949 (N_1949,N_1909,N_1908);
nor U1950 (N_1950,N_1909,N_1910);
nand U1951 (N_1951,N_1860,N_1881);
xor U1952 (N_1952,N_1885,N_1895);
nand U1953 (N_1953,N_1891,N_1878);
nand U1954 (N_1954,N_1902,N_1907);
xnor U1955 (N_1955,N_1898,N_1918);
and U1956 (N_1956,N_1910,N_1916);
nor U1957 (N_1957,N_1898,N_1895);
nand U1958 (N_1958,N_1913,N_1916);
nand U1959 (N_1959,N_1861,N_1914);
nand U1960 (N_1960,N_1892,N_1886);
or U1961 (N_1961,N_1893,N_1908);
nor U1962 (N_1962,N_1904,N_1861);
xor U1963 (N_1963,N_1863,N_1908);
nand U1964 (N_1964,N_1905,N_1918);
or U1965 (N_1965,N_1886,N_1874);
nand U1966 (N_1966,N_1867,N_1902);
nor U1967 (N_1967,N_1912,N_1918);
nor U1968 (N_1968,N_1898,N_1860);
and U1969 (N_1969,N_1895,N_1880);
nor U1970 (N_1970,N_1915,N_1888);
and U1971 (N_1971,N_1908,N_1910);
nor U1972 (N_1972,N_1894,N_1863);
nor U1973 (N_1973,N_1881,N_1912);
or U1974 (N_1974,N_1867,N_1907);
nand U1975 (N_1975,N_1888,N_1885);
nor U1976 (N_1976,N_1911,N_1888);
or U1977 (N_1977,N_1899,N_1913);
nor U1978 (N_1978,N_1863,N_1867);
nor U1979 (N_1979,N_1895,N_1886);
xor U1980 (N_1980,N_1937,N_1933);
and U1981 (N_1981,N_1961,N_1960);
nand U1982 (N_1982,N_1923,N_1966);
nand U1983 (N_1983,N_1931,N_1926);
xor U1984 (N_1984,N_1924,N_1930);
nand U1985 (N_1985,N_1947,N_1945);
or U1986 (N_1986,N_1954,N_1921);
and U1987 (N_1987,N_1963,N_1955);
nand U1988 (N_1988,N_1936,N_1949);
nor U1989 (N_1989,N_1946,N_1935);
nor U1990 (N_1990,N_1972,N_1943);
nor U1991 (N_1991,N_1964,N_1976);
nand U1992 (N_1992,N_1956,N_1971);
and U1993 (N_1993,N_1941,N_1973);
nand U1994 (N_1994,N_1968,N_1969);
xnor U1995 (N_1995,N_1965,N_1957);
xor U1996 (N_1996,N_1978,N_1928);
nor U1997 (N_1997,N_1979,N_1953);
or U1998 (N_1998,N_1939,N_1940);
or U1999 (N_1999,N_1962,N_1934);
nand U2000 (N_2000,N_1970,N_1920);
and U2001 (N_2001,N_1950,N_1951);
and U2002 (N_2002,N_1944,N_1952);
xor U2003 (N_2003,N_1948,N_1977);
and U2004 (N_2004,N_1922,N_1975);
xnor U2005 (N_2005,N_1967,N_1974);
nand U2006 (N_2006,N_1927,N_1959);
nor U2007 (N_2007,N_1925,N_1932);
or U2008 (N_2008,N_1938,N_1942);
xor U2009 (N_2009,N_1958,N_1929);
xnor U2010 (N_2010,N_1973,N_1974);
nand U2011 (N_2011,N_1940,N_1965);
or U2012 (N_2012,N_1946,N_1968);
and U2013 (N_2013,N_1978,N_1946);
nand U2014 (N_2014,N_1934,N_1977);
and U2015 (N_2015,N_1963,N_1975);
xor U2016 (N_2016,N_1933,N_1924);
or U2017 (N_2017,N_1954,N_1960);
nand U2018 (N_2018,N_1978,N_1967);
xor U2019 (N_2019,N_1923,N_1929);
or U2020 (N_2020,N_1964,N_1924);
nand U2021 (N_2021,N_1969,N_1966);
and U2022 (N_2022,N_1932,N_1944);
or U2023 (N_2023,N_1922,N_1948);
xnor U2024 (N_2024,N_1960,N_1923);
xor U2025 (N_2025,N_1945,N_1956);
nor U2026 (N_2026,N_1949,N_1939);
nand U2027 (N_2027,N_1945,N_1944);
nor U2028 (N_2028,N_1921,N_1973);
and U2029 (N_2029,N_1973,N_1944);
nor U2030 (N_2030,N_1975,N_1979);
nand U2031 (N_2031,N_1942,N_1958);
xor U2032 (N_2032,N_1934,N_1955);
or U2033 (N_2033,N_1945,N_1964);
or U2034 (N_2034,N_1977,N_1949);
nand U2035 (N_2035,N_1951,N_1920);
nor U2036 (N_2036,N_1971,N_1952);
xor U2037 (N_2037,N_1953,N_1959);
or U2038 (N_2038,N_1949,N_1937);
xor U2039 (N_2039,N_1971,N_1970);
nor U2040 (N_2040,N_2023,N_2024);
or U2041 (N_2041,N_2016,N_1986);
xnor U2042 (N_2042,N_2032,N_1994);
nand U2043 (N_2043,N_1995,N_2038);
nor U2044 (N_2044,N_2022,N_1990);
and U2045 (N_2045,N_1987,N_2019);
and U2046 (N_2046,N_2025,N_2011);
and U2047 (N_2047,N_2000,N_1985);
xnor U2048 (N_2048,N_2004,N_2031);
nand U2049 (N_2049,N_1998,N_2027);
or U2050 (N_2050,N_2020,N_2037);
xnor U2051 (N_2051,N_2018,N_2010);
and U2052 (N_2052,N_2009,N_2012);
or U2053 (N_2053,N_2001,N_2006);
or U2054 (N_2054,N_2026,N_2028);
or U2055 (N_2055,N_2007,N_2008);
and U2056 (N_2056,N_1983,N_2017);
xor U2057 (N_2057,N_1981,N_2034);
xnor U2058 (N_2058,N_2033,N_1984);
and U2059 (N_2059,N_2039,N_1993);
or U2060 (N_2060,N_2014,N_2036);
nor U2061 (N_2061,N_2035,N_1982);
or U2062 (N_2062,N_2003,N_2005);
nor U2063 (N_2063,N_2021,N_1991);
nand U2064 (N_2064,N_1997,N_2013);
nand U2065 (N_2065,N_2015,N_1988);
and U2066 (N_2066,N_2029,N_1992);
nand U2067 (N_2067,N_2002,N_2030);
nor U2068 (N_2068,N_1996,N_1989);
xnor U2069 (N_2069,N_1999,N_1980);
nor U2070 (N_2070,N_2005,N_1988);
and U2071 (N_2071,N_1991,N_1981);
nor U2072 (N_2072,N_2011,N_1985);
and U2073 (N_2073,N_1999,N_2035);
nor U2074 (N_2074,N_2031,N_1992);
and U2075 (N_2075,N_2004,N_2020);
nor U2076 (N_2076,N_1991,N_1990);
and U2077 (N_2077,N_1992,N_1994);
or U2078 (N_2078,N_2004,N_2017);
or U2079 (N_2079,N_1992,N_2003);
xor U2080 (N_2080,N_2035,N_1994);
nand U2081 (N_2081,N_1995,N_1999);
or U2082 (N_2082,N_1985,N_2026);
nand U2083 (N_2083,N_2033,N_2011);
nand U2084 (N_2084,N_1984,N_2028);
and U2085 (N_2085,N_1980,N_1991);
and U2086 (N_2086,N_2001,N_2024);
nand U2087 (N_2087,N_2008,N_2005);
xor U2088 (N_2088,N_2013,N_1990);
nand U2089 (N_2089,N_1996,N_1998);
and U2090 (N_2090,N_1998,N_2013);
xor U2091 (N_2091,N_2012,N_2016);
and U2092 (N_2092,N_2009,N_1980);
xor U2093 (N_2093,N_2022,N_1994);
and U2094 (N_2094,N_1991,N_2015);
nor U2095 (N_2095,N_2024,N_2003);
or U2096 (N_2096,N_1989,N_1992);
xor U2097 (N_2097,N_2022,N_2035);
nand U2098 (N_2098,N_2012,N_2032);
nand U2099 (N_2099,N_2021,N_1984);
xor U2100 (N_2100,N_2047,N_2080);
or U2101 (N_2101,N_2066,N_2057);
or U2102 (N_2102,N_2087,N_2051);
and U2103 (N_2103,N_2060,N_2048);
xnor U2104 (N_2104,N_2073,N_2045);
and U2105 (N_2105,N_2054,N_2055);
nand U2106 (N_2106,N_2040,N_2098);
xnor U2107 (N_2107,N_2059,N_2041);
and U2108 (N_2108,N_2078,N_2049);
nor U2109 (N_2109,N_2079,N_2050);
or U2110 (N_2110,N_2062,N_2097);
xor U2111 (N_2111,N_2083,N_2082);
xor U2112 (N_2112,N_2075,N_2056);
and U2113 (N_2113,N_2065,N_2068);
nand U2114 (N_2114,N_2063,N_2064);
or U2115 (N_2115,N_2086,N_2088);
nand U2116 (N_2116,N_2044,N_2058);
and U2117 (N_2117,N_2099,N_2071);
or U2118 (N_2118,N_2046,N_2096);
or U2119 (N_2119,N_2069,N_2043);
and U2120 (N_2120,N_2053,N_2094);
or U2121 (N_2121,N_2085,N_2093);
or U2122 (N_2122,N_2067,N_2042);
and U2123 (N_2123,N_2089,N_2095);
xnor U2124 (N_2124,N_2074,N_2070);
or U2125 (N_2125,N_2091,N_2061);
nand U2126 (N_2126,N_2081,N_2052);
or U2127 (N_2127,N_2092,N_2076);
xor U2128 (N_2128,N_2090,N_2077);
and U2129 (N_2129,N_2072,N_2084);
and U2130 (N_2130,N_2058,N_2082);
xnor U2131 (N_2131,N_2062,N_2040);
nand U2132 (N_2132,N_2082,N_2045);
nor U2133 (N_2133,N_2092,N_2083);
xor U2134 (N_2134,N_2064,N_2041);
nand U2135 (N_2135,N_2071,N_2083);
and U2136 (N_2136,N_2078,N_2052);
nand U2137 (N_2137,N_2088,N_2053);
or U2138 (N_2138,N_2049,N_2043);
and U2139 (N_2139,N_2049,N_2097);
nor U2140 (N_2140,N_2074,N_2085);
or U2141 (N_2141,N_2094,N_2087);
nor U2142 (N_2142,N_2097,N_2076);
xor U2143 (N_2143,N_2064,N_2048);
nand U2144 (N_2144,N_2099,N_2068);
xnor U2145 (N_2145,N_2076,N_2063);
xor U2146 (N_2146,N_2052,N_2070);
nand U2147 (N_2147,N_2092,N_2080);
nand U2148 (N_2148,N_2061,N_2096);
nand U2149 (N_2149,N_2055,N_2098);
or U2150 (N_2150,N_2094,N_2083);
and U2151 (N_2151,N_2090,N_2097);
and U2152 (N_2152,N_2082,N_2072);
xor U2153 (N_2153,N_2084,N_2090);
nor U2154 (N_2154,N_2082,N_2056);
xor U2155 (N_2155,N_2040,N_2060);
nor U2156 (N_2156,N_2070,N_2062);
xnor U2157 (N_2157,N_2061,N_2043);
xnor U2158 (N_2158,N_2083,N_2078);
nand U2159 (N_2159,N_2058,N_2083);
and U2160 (N_2160,N_2109,N_2158);
and U2161 (N_2161,N_2122,N_2152);
and U2162 (N_2162,N_2102,N_2115);
and U2163 (N_2163,N_2126,N_2139);
xnor U2164 (N_2164,N_2141,N_2155);
nand U2165 (N_2165,N_2150,N_2100);
nor U2166 (N_2166,N_2125,N_2118);
nor U2167 (N_2167,N_2121,N_2156);
or U2168 (N_2168,N_2142,N_2147);
and U2169 (N_2169,N_2104,N_2134);
xor U2170 (N_2170,N_2107,N_2153);
and U2171 (N_2171,N_2135,N_2114);
and U2172 (N_2172,N_2127,N_2128);
xor U2173 (N_2173,N_2124,N_2148);
nand U2174 (N_2174,N_2113,N_2116);
and U2175 (N_2175,N_2108,N_2106);
and U2176 (N_2176,N_2112,N_2138);
nor U2177 (N_2177,N_2131,N_2105);
xnor U2178 (N_2178,N_2130,N_2119);
xnor U2179 (N_2179,N_2154,N_2143);
nor U2180 (N_2180,N_2144,N_2129);
or U2181 (N_2181,N_2123,N_2140);
and U2182 (N_2182,N_2159,N_2120);
nor U2183 (N_2183,N_2101,N_2133);
and U2184 (N_2184,N_2146,N_2132);
xnor U2185 (N_2185,N_2117,N_2149);
xor U2186 (N_2186,N_2151,N_2111);
and U2187 (N_2187,N_2110,N_2157);
xor U2188 (N_2188,N_2145,N_2103);
nand U2189 (N_2189,N_2137,N_2136);
or U2190 (N_2190,N_2125,N_2147);
or U2191 (N_2191,N_2128,N_2113);
or U2192 (N_2192,N_2111,N_2129);
xnor U2193 (N_2193,N_2130,N_2152);
and U2194 (N_2194,N_2153,N_2149);
or U2195 (N_2195,N_2144,N_2139);
and U2196 (N_2196,N_2132,N_2115);
nor U2197 (N_2197,N_2137,N_2110);
nor U2198 (N_2198,N_2154,N_2159);
nand U2199 (N_2199,N_2115,N_2122);
or U2200 (N_2200,N_2118,N_2147);
xnor U2201 (N_2201,N_2151,N_2108);
nor U2202 (N_2202,N_2115,N_2131);
and U2203 (N_2203,N_2133,N_2157);
or U2204 (N_2204,N_2136,N_2138);
nand U2205 (N_2205,N_2117,N_2100);
or U2206 (N_2206,N_2146,N_2140);
xnor U2207 (N_2207,N_2119,N_2126);
nor U2208 (N_2208,N_2137,N_2131);
or U2209 (N_2209,N_2158,N_2137);
or U2210 (N_2210,N_2119,N_2122);
nor U2211 (N_2211,N_2133,N_2144);
xnor U2212 (N_2212,N_2114,N_2129);
xnor U2213 (N_2213,N_2134,N_2157);
or U2214 (N_2214,N_2109,N_2153);
or U2215 (N_2215,N_2155,N_2146);
xor U2216 (N_2216,N_2111,N_2139);
and U2217 (N_2217,N_2115,N_2123);
or U2218 (N_2218,N_2120,N_2153);
and U2219 (N_2219,N_2146,N_2122);
or U2220 (N_2220,N_2168,N_2202);
nor U2221 (N_2221,N_2190,N_2216);
xor U2222 (N_2222,N_2201,N_2204);
or U2223 (N_2223,N_2160,N_2188);
nor U2224 (N_2224,N_2186,N_2174);
and U2225 (N_2225,N_2184,N_2171);
nor U2226 (N_2226,N_2207,N_2214);
nand U2227 (N_2227,N_2164,N_2189);
and U2228 (N_2228,N_2178,N_2173);
nand U2229 (N_2229,N_2215,N_2210);
nor U2230 (N_2230,N_2162,N_2199);
nand U2231 (N_2231,N_2187,N_2175);
xor U2232 (N_2232,N_2208,N_2177);
and U2233 (N_2233,N_2195,N_2218);
or U2234 (N_2234,N_2198,N_2209);
xor U2235 (N_2235,N_2161,N_2205);
or U2236 (N_2236,N_2217,N_2166);
xnor U2237 (N_2237,N_2212,N_2182);
nor U2238 (N_2238,N_2181,N_2213);
nand U2239 (N_2239,N_2167,N_2194);
or U2240 (N_2240,N_2206,N_2196);
nand U2241 (N_2241,N_2211,N_2172);
xnor U2242 (N_2242,N_2197,N_2185);
nand U2243 (N_2243,N_2179,N_2170);
xnor U2244 (N_2244,N_2192,N_2203);
and U2245 (N_2245,N_2191,N_2183);
xnor U2246 (N_2246,N_2180,N_2169);
xnor U2247 (N_2247,N_2165,N_2193);
and U2248 (N_2248,N_2200,N_2176);
or U2249 (N_2249,N_2163,N_2219);
nor U2250 (N_2250,N_2199,N_2167);
nor U2251 (N_2251,N_2217,N_2194);
or U2252 (N_2252,N_2181,N_2160);
nand U2253 (N_2253,N_2165,N_2208);
or U2254 (N_2254,N_2200,N_2216);
or U2255 (N_2255,N_2189,N_2198);
nand U2256 (N_2256,N_2214,N_2204);
xnor U2257 (N_2257,N_2185,N_2195);
nand U2258 (N_2258,N_2192,N_2185);
xnor U2259 (N_2259,N_2197,N_2172);
nor U2260 (N_2260,N_2207,N_2174);
and U2261 (N_2261,N_2184,N_2181);
and U2262 (N_2262,N_2162,N_2179);
nand U2263 (N_2263,N_2176,N_2172);
nor U2264 (N_2264,N_2199,N_2213);
nor U2265 (N_2265,N_2207,N_2198);
or U2266 (N_2266,N_2176,N_2208);
nand U2267 (N_2267,N_2188,N_2177);
and U2268 (N_2268,N_2176,N_2190);
nor U2269 (N_2269,N_2171,N_2200);
nor U2270 (N_2270,N_2217,N_2163);
xor U2271 (N_2271,N_2171,N_2209);
xnor U2272 (N_2272,N_2212,N_2217);
nor U2273 (N_2273,N_2205,N_2211);
and U2274 (N_2274,N_2174,N_2162);
or U2275 (N_2275,N_2201,N_2219);
nor U2276 (N_2276,N_2207,N_2188);
and U2277 (N_2277,N_2160,N_2214);
or U2278 (N_2278,N_2193,N_2219);
and U2279 (N_2279,N_2162,N_2217);
xnor U2280 (N_2280,N_2248,N_2230);
or U2281 (N_2281,N_2263,N_2251);
nor U2282 (N_2282,N_2240,N_2229);
nor U2283 (N_2283,N_2225,N_2272);
nand U2284 (N_2284,N_2239,N_2255);
nand U2285 (N_2285,N_2242,N_2220);
nor U2286 (N_2286,N_2277,N_2236);
and U2287 (N_2287,N_2245,N_2265);
xnor U2288 (N_2288,N_2224,N_2270);
and U2289 (N_2289,N_2275,N_2233);
nor U2290 (N_2290,N_2228,N_2264);
nand U2291 (N_2291,N_2223,N_2249);
or U2292 (N_2292,N_2237,N_2246);
nor U2293 (N_2293,N_2244,N_2269);
nand U2294 (N_2294,N_2226,N_2274);
and U2295 (N_2295,N_2222,N_2267);
and U2296 (N_2296,N_2261,N_2238);
nor U2297 (N_2297,N_2268,N_2235);
and U2298 (N_2298,N_2227,N_2231);
or U2299 (N_2299,N_2273,N_2276);
nor U2300 (N_2300,N_2259,N_2257);
or U2301 (N_2301,N_2258,N_2271);
nor U2302 (N_2302,N_2256,N_2279);
or U2303 (N_2303,N_2247,N_2262);
nor U2304 (N_2304,N_2260,N_2234);
and U2305 (N_2305,N_2266,N_2252);
nor U2306 (N_2306,N_2221,N_2232);
nor U2307 (N_2307,N_2254,N_2253);
and U2308 (N_2308,N_2241,N_2250);
nor U2309 (N_2309,N_2243,N_2278);
and U2310 (N_2310,N_2235,N_2222);
nor U2311 (N_2311,N_2245,N_2270);
nand U2312 (N_2312,N_2249,N_2273);
or U2313 (N_2313,N_2255,N_2233);
nor U2314 (N_2314,N_2275,N_2262);
nor U2315 (N_2315,N_2230,N_2226);
nor U2316 (N_2316,N_2227,N_2269);
and U2317 (N_2317,N_2246,N_2226);
or U2318 (N_2318,N_2271,N_2278);
or U2319 (N_2319,N_2277,N_2224);
nor U2320 (N_2320,N_2269,N_2278);
and U2321 (N_2321,N_2265,N_2271);
nor U2322 (N_2322,N_2239,N_2244);
nor U2323 (N_2323,N_2267,N_2260);
or U2324 (N_2324,N_2252,N_2251);
nor U2325 (N_2325,N_2278,N_2274);
nand U2326 (N_2326,N_2224,N_2234);
or U2327 (N_2327,N_2237,N_2265);
nand U2328 (N_2328,N_2278,N_2277);
or U2329 (N_2329,N_2275,N_2273);
nand U2330 (N_2330,N_2279,N_2263);
and U2331 (N_2331,N_2273,N_2229);
nor U2332 (N_2332,N_2240,N_2238);
and U2333 (N_2333,N_2246,N_2250);
nor U2334 (N_2334,N_2221,N_2220);
nor U2335 (N_2335,N_2232,N_2267);
xor U2336 (N_2336,N_2265,N_2259);
nand U2337 (N_2337,N_2222,N_2253);
or U2338 (N_2338,N_2252,N_2237);
nor U2339 (N_2339,N_2256,N_2269);
nor U2340 (N_2340,N_2295,N_2285);
xnor U2341 (N_2341,N_2339,N_2331);
and U2342 (N_2342,N_2309,N_2306);
nand U2343 (N_2343,N_2286,N_2317);
nand U2344 (N_2344,N_2316,N_2305);
xor U2345 (N_2345,N_2313,N_2303);
or U2346 (N_2346,N_2289,N_2315);
nand U2347 (N_2347,N_2290,N_2333);
nor U2348 (N_2348,N_2292,N_2319);
nand U2349 (N_2349,N_2320,N_2307);
nor U2350 (N_2350,N_2281,N_2294);
nand U2351 (N_2351,N_2284,N_2296);
nor U2352 (N_2352,N_2337,N_2336);
nor U2353 (N_2353,N_2335,N_2327);
nor U2354 (N_2354,N_2288,N_2326);
or U2355 (N_2355,N_2334,N_2328);
or U2356 (N_2356,N_2293,N_2325);
nor U2357 (N_2357,N_2282,N_2300);
nor U2358 (N_2358,N_2310,N_2302);
or U2359 (N_2359,N_2304,N_2287);
xnor U2360 (N_2360,N_2332,N_2321);
nor U2361 (N_2361,N_2283,N_2318);
and U2362 (N_2362,N_2322,N_2314);
and U2363 (N_2363,N_2338,N_2308);
nand U2364 (N_2364,N_2280,N_2298);
xnor U2365 (N_2365,N_2311,N_2329);
xnor U2366 (N_2366,N_2291,N_2312);
nor U2367 (N_2367,N_2330,N_2301);
xor U2368 (N_2368,N_2299,N_2297);
and U2369 (N_2369,N_2324,N_2323);
xnor U2370 (N_2370,N_2289,N_2299);
nand U2371 (N_2371,N_2289,N_2285);
nand U2372 (N_2372,N_2323,N_2309);
or U2373 (N_2373,N_2281,N_2316);
and U2374 (N_2374,N_2308,N_2313);
nand U2375 (N_2375,N_2291,N_2337);
nand U2376 (N_2376,N_2298,N_2338);
or U2377 (N_2377,N_2301,N_2283);
or U2378 (N_2378,N_2288,N_2299);
nor U2379 (N_2379,N_2312,N_2307);
and U2380 (N_2380,N_2330,N_2335);
or U2381 (N_2381,N_2316,N_2320);
or U2382 (N_2382,N_2317,N_2312);
or U2383 (N_2383,N_2302,N_2307);
or U2384 (N_2384,N_2334,N_2339);
and U2385 (N_2385,N_2282,N_2299);
or U2386 (N_2386,N_2311,N_2334);
nor U2387 (N_2387,N_2311,N_2322);
or U2388 (N_2388,N_2322,N_2285);
xnor U2389 (N_2389,N_2287,N_2301);
xor U2390 (N_2390,N_2290,N_2305);
or U2391 (N_2391,N_2296,N_2324);
xor U2392 (N_2392,N_2338,N_2325);
and U2393 (N_2393,N_2284,N_2289);
or U2394 (N_2394,N_2309,N_2336);
or U2395 (N_2395,N_2325,N_2297);
nand U2396 (N_2396,N_2332,N_2314);
nand U2397 (N_2397,N_2319,N_2333);
or U2398 (N_2398,N_2336,N_2324);
and U2399 (N_2399,N_2318,N_2308);
nor U2400 (N_2400,N_2362,N_2388);
or U2401 (N_2401,N_2341,N_2369);
nand U2402 (N_2402,N_2384,N_2349);
nand U2403 (N_2403,N_2354,N_2381);
or U2404 (N_2404,N_2399,N_2355);
or U2405 (N_2405,N_2345,N_2394);
nand U2406 (N_2406,N_2375,N_2385);
or U2407 (N_2407,N_2376,N_2395);
or U2408 (N_2408,N_2387,N_2391);
and U2409 (N_2409,N_2348,N_2380);
and U2410 (N_2410,N_2396,N_2366);
and U2411 (N_2411,N_2378,N_2363);
nor U2412 (N_2412,N_2353,N_2379);
xnor U2413 (N_2413,N_2360,N_2342);
or U2414 (N_2414,N_2364,N_2377);
and U2415 (N_2415,N_2367,N_2389);
and U2416 (N_2416,N_2340,N_2356);
and U2417 (N_2417,N_2371,N_2368);
or U2418 (N_2418,N_2393,N_2346);
xnor U2419 (N_2419,N_2359,N_2365);
nor U2420 (N_2420,N_2351,N_2373);
xor U2421 (N_2421,N_2397,N_2374);
xnor U2422 (N_2422,N_2347,N_2386);
nor U2423 (N_2423,N_2352,N_2344);
nand U2424 (N_2424,N_2398,N_2390);
or U2425 (N_2425,N_2357,N_2392);
and U2426 (N_2426,N_2350,N_2343);
or U2427 (N_2427,N_2361,N_2372);
xor U2428 (N_2428,N_2370,N_2383);
xor U2429 (N_2429,N_2358,N_2382);
nand U2430 (N_2430,N_2352,N_2378);
or U2431 (N_2431,N_2388,N_2372);
nand U2432 (N_2432,N_2390,N_2387);
and U2433 (N_2433,N_2341,N_2398);
nand U2434 (N_2434,N_2392,N_2354);
nor U2435 (N_2435,N_2364,N_2376);
nor U2436 (N_2436,N_2392,N_2360);
xor U2437 (N_2437,N_2361,N_2376);
nor U2438 (N_2438,N_2396,N_2385);
and U2439 (N_2439,N_2354,N_2376);
nand U2440 (N_2440,N_2379,N_2376);
nor U2441 (N_2441,N_2377,N_2359);
xor U2442 (N_2442,N_2375,N_2393);
nor U2443 (N_2443,N_2358,N_2369);
nand U2444 (N_2444,N_2368,N_2398);
or U2445 (N_2445,N_2356,N_2378);
xnor U2446 (N_2446,N_2374,N_2368);
and U2447 (N_2447,N_2343,N_2391);
or U2448 (N_2448,N_2358,N_2366);
nor U2449 (N_2449,N_2373,N_2345);
nor U2450 (N_2450,N_2356,N_2357);
or U2451 (N_2451,N_2374,N_2344);
nor U2452 (N_2452,N_2377,N_2362);
xor U2453 (N_2453,N_2396,N_2377);
or U2454 (N_2454,N_2358,N_2389);
nor U2455 (N_2455,N_2377,N_2369);
nor U2456 (N_2456,N_2380,N_2354);
and U2457 (N_2457,N_2375,N_2376);
xnor U2458 (N_2458,N_2398,N_2388);
and U2459 (N_2459,N_2357,N_2345);
xor U2460 (N_2460,N_2455,N_2405);
nand U2461 (N_2461,N_2400,N_2416);
and U2462 (N_2462,N_2401,N_2403);
nor U2463 (N_2463,N_2430,N_2427);
xor U2464 (N_2464,N_2426,N_2428);
or U2465 (N_2465,N_2425,N_2421);
and U2466 (N_2466,N_2402,N_2444);
nand U2467 (N_2467,N_2448,N_2441);
xnor U2468 (N_2468,N_2446,N_2423);
nor U2469 (N_2469,N_2412,N_2406);
and U2470 (N_2470,N_2407,N_2422);
xnor U2471 (N_2471,N_2431,N_2437);
xnor U2472 (N_2472,N_2439,N_2457);
nor U2473 (N_2473,N_2418,N_2409);
xor U2474 (N_2474,N_2436,N_2417);
or U2475 (N_2475,N_2442,N_2433);
nor U2476 (N_2476,N_2404,N_2419);
and U2477 (N_2477,N_2435,N_2451);
nor U2478 (N_2478,N_2413,N_2408);
nand U2479 (N_2479,N_2443,N_2415);
nor U2480 (N_2480,N_2458,N_2434);
or U2481 (N_2481,N_2420,N_2445);
and U2482 (N_2482,N_2432,N_2459);
xnor U2483 (N_2483,N_2450,N_2411);
nand U2484 (N_2484,N_2424,N_2414);
xor U2485 (N_2485,N_2454,N_2452);
xnor U2486 (N_2486,N_2440,N_2429);
or U2487 (N_2487,N_2447,N_2453);
and U2488 (N_2488,N_2449,N_2456);
xor U2489 (N_2489,N_2438,N_2410);
nand U2490 (N_2490,N_2438,N_2445);
and U2491 (N_2491,N_2440,N_2448);
nand U2492 (N_2492,N_2433,N_2440);
xnor U2493 (N_2493,N_2455,N_2414);
nor U2494 (N_2494,N_2415,N_2442);
xor U2495 (N_2495,N_2418,N_2439);
nand U2496 (N_2496,N_2457,N_2443);
and U2497 (N_2497,N_2400,N_2448);
nand U2498 (N_2498,N_2420,N_2423);
nand U2499 (N_2499,N_2404,N_2444);
nand U2500 (N_2500,N_2411,N_2432);
xnor U2501 (N_2501,N_2457,N_2452);
and U2502 (N_2502,N_2424,N_2402);
and U2503 (N_2503,N_2427,N_2453);
nor U2504 (N_2504,N_2441,N_2402);
nand U2505 (N_2505,N_2446,N_2445);
nand U2506 (N_2506,N_2448,N_2422);
nor U2507 (N_2507,N_2437,N_2409);
and U2508 (N_2508,N_2442,N_2452);
nor U2509 (N_2509,N_2419,N_2436);
nand U2510 (N_2510,N_2426,N_2414);
and U2511 (N_2511,N_2447,N_2424);
nor U2512 (N_2512,N_2435,N_2436);
nand U2513 (N_2513,N_2454,N_2450);
nand U2514 (N_2514,N_2427,N_2448);
and U2515 (N_2515,N_2431,N_2405);
xnor U2516 (N_2516,N_2443,N_2401);
or U2517 (N_2517,N_2456,N_2428);
or U2518 (N_2518,N_2404,N_2401);
or U2519 (N_2519,N_2458,N_2402);
xnor U2520 (N_2520,N_2476,N_2518);
or U2521 (N_2521,N_2510,N_2493);
and U2522 (N_2522,N_2482,N_2460);
or U2523 (N_2523,N_2500,N_2472);
and U2524 (N_2524,N_2513,N_2468);
or U2525 (N_2525,N_2470,N_2488);
xor U2526 (N_2526,N_2487,N_2506);
xnor U2527 (N_2527,N_2465,N_2490);
nand U2528 (N_2528,N_2497,N_2463);
or U2529 (N_2529,N_2517,N_2496);
and U2530 (N_2530,N_2502,N_2509);
xor U2531 (N_2531,N_2466,N_2512);
or U2532 (N_2532,N_2477,N_2486);
or U2533 (N_2533,N_2484,N_2489);
and U2534 (N_2534,N_2464,N_2480);
nand U2535 (N_2535,N_2479,N_2461);
xor U2536 (N_2536,N_2519,N_2474);
xor U2537 (N_2537,N_2462,N_2508);
nor U2538 (N_2538,N_2498,N_2483);
xnor U2539 (N_2539,N_2516,N_2494);
nor U2540 (N_2540,N_2492,N_2515);
nor U2541 (N_2541,N_2485,N_2504);
nor U2542 (N_2542,N_2481,N_2495);
and U2543 (N_2543,N_2507,N_2471);
and U2544 (N_2544,N_2511,N_2467);
nor U2545 (N_2545,N_2501,N_2475);
nand U2546 (N_2546,N_2505,N_2491);
xnor U2547 (N_2547,N_2503,N_2473);
nand U2548 (N_2548,N_2478,N_2499);
and U2549 (N_2549,N_2469,N_2514);
and U2550 (N_2550,N_2464,N_2510);
nor U2551 (N_2551,N_2484,N_2512);
or U2552 (N_2552,N_2485,N_2465);
nor U2553 (N_2553,N_2505,N_2495);
nor U2554 (N_2554,N_2468,N_2475);
nor U2555 (N_2555,N_2480,N_2482);
xnor U2556 (N_2556,N_2498,N_2501);
nand U2557 (N_2557,N_2486,N_2488);
nand U2558 (N_2558,N_2483,N_2492);
nand U2559 (N_2559,N_2478,N_2497);
nand U2560 (N_2560,N_2502,N_2514);
and U2561 (N_2561,N_2498,N_2486);
xor U2562 (N_2562,N_2473,N_2519);
and U2563 (N_2563,N_2495,N_2512);
xor U2564 (N_2564,N_2490,N_2500);
xor U2565 (N_2565,N_2519,N_2481);
or U2566 (N_2566,N_2493,N_2506);
and U2567 (N_2567,N_2477,N_2473);
and U2568 (N_2568,N_2466,N_2484);
and U2569 (N_2569,N_2480,N_2516);
nand U2570 (N_2570,N_2461,N_2467);
nand U2571 (N_2571,N_2504,N_2463);
nand U2572 (N_2572,N_2509,N_2475);
nor U2573 (N_2573,N_2517,N_2518);
xor U2574 (N_2574,N_2498,N_2491);
nor U2575 (N_2575,N_2468,N_2470);
nand U2576 (N_2576,N_2483,N_2517);
nor U2577 (N_2577,N_2462,N_2467);
nand U2578 (N_2578,N_2504,N_2465);
and U2579 (N_2579,N_2498,N_2472);
or U2580 (N_2580,N_2526,N_2559);
nor U2581 (N_2581,N_2546,N_2552);
or U2582 (N_2582,N_2553,N_2536);
or U2583 (N_2583,N_2578,N_2527);
and U2584 (N_2584,N_2548,N_2547);
or U2585 (N_2585,N_2533,N_2524);
nor U2586 (N_2586,N_2544,N_2534);
nor U2587 (N_2587,N_2542,N_2523);
nor U2588 (N_2588,N_2564,N_2577);
and U2589 (N_2589,N_2576,N_2573);
and U2590 (N_2590,N_2570,N_2561);
xnor U2591 (N_2591,N_2558,N_2528);
nor U2592 (N_2592,N_2571,N_2545);
and U2593 (N_2593,N_2568,N_2560);
and U2594 (N_2594,N_2557,N_2531);
xnor U2595 (N_2595,N_2540,N_2520);
or U2596 (N_2596,N_2551,N_2538);
xor U2597 (N_2597,N_2549,N_2529);
and U2598 (N_2598,N_2543,N_2525);
or U2599 (N_2599,N_2554,N_2530);
nand U2600 (N_2600,N_2521,N_2535);
and U2601 (N_2601,N_2532,N_2572);
or U2602 (N_2602,N_2562,N_2522);
or U2603 (N_2603,N_2574,N_2550);
or U2604 (N_2604,N_2579,N_2555);
nand U2605 (N_2605,N_2537,N_2556);
or U2606 (N_2606,N_2541,N_2565);
xor U2607 (N_2607,N_2575,N_2567);
or U2608 (N_2608,N_2566,N_2563);
nor U2609 (N_2609,N_2539,N_2569);
xor U2610 (N_2610,N_2571,N_2531);
and U2611 (N_2611,N_2523,N_2567);
xor U2612 (N_2612,N_2577,N_2547);
or U2613 (N_2613,N_2527,N_2547);
or U2614 (N_2614,N_2549,N_2577);
or U2615 (N_2615,N_2533,N_2553);
nand U2616 (N_2616,N_2538,N_2572);
or U2617 (N_2617,N_2526,N_2562);
and U2618 (N_2618,N_2553,N_2558);
or U2619 (N_2619,N_2552,N_2561);
and U2620 (N_2620,N_2548,N_2528);
xor U2621 (N_2621,N_2530,N_2556);
xnor U2622 (N_2622,N_2544,N_2576);
or U2623 (N_2623,N_2525,N_2548);
and U2624 (N_2624,N_2566,N_2524);
nand U2625 (N_2625,N_2573,N_2564);
or U2626 (N_2626,N_2543,N_2524);
xnor U2627 (N_2627,N_2541,N_2533);
nand U2628 (N_2628,N_2542,N_2546);
nand U2629 (N_2629,N_2561,N_2548);
nor U2630 (N_2630,N_2568,N_2564);
nor U2631 (N_2631,N_2578,N_2567);
nor U2632 (N_2632,N_2565,N_2542);
xnor U2633 (N_2633,N_2546,N_2575);
nand U2634 (N_2634,N_2567,N_2541);
or U2635 (N_2635,N_2561,N_2572);
and U2636 (N_2636,N_2529,N_2544);
or U2637 (N_2637,N_2551,N_2542);
nor U2638 (N_2638,N_2520,N_2573);
xnor U2639 (N_2639,N_2536,N_2531);
nor U2640 (N_2640,N_2609,N_2613);
nand U2641 (N_2641,N_2584,N_2628);
or U2642 (N_2642,N_2582,N_2638);
and U2643 (N_2643,N_2603,N_2580);
or U2644 (N_2644,N_2630,N_2618);
and U2645 (N_2645,N_2622,N_2631);
xnor U2646 (N_2646,N_2624,N_2588);
or U2647 (N_2647,N_2601,N_2633);
and U2648 (N_2648,N_2608,N_2611);
nor U2649 (N_2649,N_2637,N_2626);
and U2650 (N_2650,N_2587,N_2607);
nor U2651 (N_2651,N_2610,N_2592);
xor U2652 (N_2652,N_2606,N_2639);
nor U2653 (N_2653,N_2586,N_2617);
nor U2654 (N_2654,N_2604,N_2600);
and U2655 (N_2655,N_2620,N_2589);
or U2656 (N_2656,N_2623,N_2585);
xnor U2657 (N_2657,N_2583,N_2621);
nor U2658 (N_2658,N_2634,N_2636);
nor U2659 (N_2659,N_2616,N_2594);
xor U2660 (N_2660,N_2612,N_2635);
and U2661 (N_2661,N_2581,N_2627);
xnor U2662 (N_2662,N_2615,N_2590);
and U2663 (N_2663,N_2597,N_2596);
xor U2664 (N_2664,N_2602,N_2614);
xor U2665 (N_2665,N_2598,N_2632);
and U2666 (N_2666,N_2595,N_2625);
and U2667 (N_2667,N_2591,N_2605);
nor U2668 (N_2668,N_2619,N_2593);
and U2669 (N_2669,N_2629,N_2599);
nor U2670 (N_2670,N_2609,N_2604);
and U2671 (N_2671,N_2596,N_2608);
nand U2672 (N_2672,N_2581,N_2606);
xor U2673 (N_2673,N_2596,N_2601);
or U2674 (N_2674,N_2586,N_2611);
nor U2675 (N_2675,N_2632,N_2588);
and U2676 (N_2676,N_2623,N_2600);
and U2677 (N_2677,N_2599,N_2632);
xnor U2678 (N_2678,N_2584,N_2638);
and U2679 (N_2679,N_2582,N_2624);
nand U2680 (N_2680,N_2585,N_2622);
or U2681 (N_2681,N_2586,N_2599);
nand U2682 (N_2682,N_2616,N_2607);
nand U2683 (N_2683,N_2621,N_2600);
nand U2684 (N_2684,N_2584,N_2592);
nor U2685 (N_2685,N_2597,N_2607);
or U2686 (N_2686,N_2606,N_2621);
or U2687 (N_2687,N_2601,N_2630);
nor U2688 (N_2688,N_2592,N_2615);
nor U2689 (N_2689,N_2636,N_2587);
and U2690 (N_2690,N_2618,N_2623);
and U2691 (N_2691,N_2596,N_2628);
xor U2692 (N_2692,N_2637,N_2587);
xnor U2693 (N_2693,N_2581,N_2607);
nand U2694 (N_2694,N_2628,N_2624);
and U2695 (N_2695,N_2619,N_2610);
xnor U2696 (N_2696,N_2623,N_2625);
nand U2697 (N_2697,N_2587,N_2622);
or U2698 (N_2698,N_2606,N_2605);
and U2699 (N_2699,N_2597,N_2595);
nand U2700 (N_2700,N_2646,N_2650);
xor U2701 (N_2701,N_2684,N_2651);
nand U2702 (N_2702,N_2662,N_2663);
or U2703 (N_2703,N_2690,N_2656);
or U2704 (N_2704,N_2643,N_2694);
or U2705 (N_2705,N_2641,N_2654);
nor U2706 (N_2706,N_2676,N_2687);
and U2707 (N_2707,N_2679,N_2649);
nand U2708 (N_2708,N_2647,N_2665);
and U2709 (N_2709,N_2695,N_2668);
and U2710 (N_2710,N_2652,N_2677);
and U2711 (N_2711,N_2657,N_2692);
and U2712 (N_2712,N_2689,N_2669);
or U2713 (N_2713,N_2660,N_2671);
xnor U2714 (N_2714,N_2672,N_2699);
or U2715 (N_2715,N_2680,N_2683);
nand U2716 (N_2716,N_2658,N_2681);
nor U2717 (N_2717,N_2640,N_2655);
or U2718 (N_2718,N_2667,N_2686);
and U2719 (N_2719,N_2659,N_2678);
and U2720 (N_2720,N_2697,N_2653);
xnor U2721 (N_2721,N_2693,N_2648);
xor U2722 (N_2722,N_2675,N_2698);
xnor U2723 (N_2723,N_2644,N_2661);
xor U2724 (N_2724,N_2682,N_2696);
nor U2725 (N_2725,N_2664,N_2645);
and U2726 (N_2726,N_2688,N_2642);
nor U2727 (N_2727,N_2673,N_2666);
nand U2728 (N_2728,N_2691,N_2674);
nand U2729 (N_2729,N_2685,N_2670);
and U2730 (N_2730,N_2676,N_2699);
or U2731 (N_2731,N_2694,N_2688);
or U2732 (N_2732,N_2690,N_2650);
nand U2733 (N_2733,N_2646,N_2657);
or U2734 (N_2734,N_2696,N_2681);
nand U2735 (N_2735,N_2693,N_2691);
nor U2736 (N_2736,N_2672,N_2673);
nand U2737 (N_2737,N_2676,N_2671);
xor U2738 (N_2738,N_2656,N_2655);
and U2739 (N_2739,N_2643,N_2655);
or U2740 (N_2740,N_2687,N_2691);
xor U2741 (N_2741,N_2676,N_2681);
and U2742 (N_2742,N_2675,N_2679);
xnor U2743 (N_2743,N_2693,N_2661);
xnor U2744 (N_2744,N_2682,N_2667);
or U2745 (N_2745,N_2646,N_2640);
xor U2746 (N_2746,N_2650,N_2657);
and U2747 (N_2747,N_2682,N_2688);
or U2748 (N_2748,N_2649,N_2652);
nand U2749 (N_2749,N_2668,N_2667);
and U2750 (N_2750,N_2683,N_2686);
or U2751 (N_2751,N_2674,N_2667);
nor U2752 (N_2752,N_2648,N_2688);
or U2753 (N_2753,N_2659,N_2656);
or U2754 (N_2754,N_2645,N_2656);
nor U2755 (N_2755,N_2647,N_2691);
and U2756 (N_2756,N_2682,N_2642);
nand U2757 (N_2757,N_2653,N_2671);
nand U2758 (N_2758,N_2657,N_2648);
and U2759 (N_2759,N_2685,N_2681);
nand U2760 (N_2760,N_2730,N_2713);
nand U2761 (N_2761,N_2741,N_2719);
and U2762 (N_2762,N_2710,N_2718);
and U2763 (N_2763,N_2708,N_2747);
or U2764 (N_2764,N_2704,N_2723);
xnor U2765 (N_2765,N_2736,N_2716);
nand U2766 (N_2766,N_2750,N_2739);
xor U2767 (N_2767,N_2758,N_2700);
xnor U2768 (N_2768,N_2720,N_2717);
nand U2769 (N_2769,N_2743,N_2721);
or U2770 (N_2770,N_2722,N_2748);
xnor U2771 (N_2771,N_2755,N_2749);
and U2772 (N_2772,N_2754,N_2746);
or U2773 (N_2773,N_2701,N_2727);
nand U2774 (N_2774,N_2738,N_2705);
or U2775 (N_2775,N_2732,N_2734);
nand U2776 (N_2776,N_2702,N_2715);
and U2777 (N_2777,N_2744,N_2703);
nand U2778 (N_2778,N_2731,N_2726);
and U2779 (N_2779,N_2714,N_2733);
and U2780 (N_2780,N_2742,N_2728);
nor U2781 (N_2781,N_2752,N_2706);
or U2782 (N_2782,N_2759,N_2712);
xor U2783 (N_2783,N_2753,N_2711);
and U2784 (N_2784,N_2709,N_2740);
and U2785 (N_2785,N_2724,N_2737);
and U2786 (N_2786,N_2729,N_2745);
and U2787 (N_2787,N_2757,N_2751);
nand U2788 (N_2788,N_2756,N_2735);
nand U2789 (N_2789,N_2707,N_2725);
xor U2790 (N_2790,N_2732,N_2733);
nand U2791 (N_2791,N_2744,N_2722);
xor U2792 (N_2792,N_2753,N_2755);
nor U2793 (N_2793,N_2751,N_2725);
xnor U2794 (N_2794,N_2732,N_2719);
nand U2795 (N_2795,N_2754,N_2750);
nor U2796 (N_2796,N_2729,N_2710);
and U2797 (N_2797,N_2719,N_2755);
xor U2798 (N_2798,N_2751,N_2726);
nor U2799 (N_2799,N_2710,N_2719);
nand U2800 (N_2800,N_2730,N_2717);
and U2801 (N_2801,N_2733,N_2705);
nand U2802 (N_2802,N_2718,N_2728);
or U2803 (N_2803,N_2738,N_2749);
nor U2804 (N_2804,N_2734,N_2708);
nor U2805 (N_2805,N_2728,N_2736);
nor U2806 (N_2806,N_2750,N_2716);
and U2807 (N_2807,N_2706,N_2712);
and U2808 (N_2808,N_2734,N_2740);
and U2809 (N_2809,N_2726,N_2706);
or U2810 (N_2810,N_2743,N_2702);
and U2811 (N_2811,N_2714,N_2704);
and U2812 (N_2812,N_2726,N_2710);
and U2813 (N_2813,N_2715,N_2738);
and U2814 (N_2814,N_2724,N_2727);
or U2815 (N_2815,N_2736,N_2749);
nand U2816 (N_2816,N_2709,N_2730);
nand U2817 (N_2817,N_2727,N_2711);
xnor U2818 (N_2818,N_2703,N_2728);
nand U2819 (N_2819,N_2726,N_2700);
and U2820 (N_2820,N_2771,N_2791);
and U2821 (N_2821,N_2808,N_2780);
and U2822 (N_2822,N_2775,N_2793);
and U2823 (N_2823,N_2786,N_2807);
and U2824 (N_2824,N_2781,N_2815);
nand U2825 (N_2825,N_2765,N_2800);
xnor U2826 (N_2826,N_2810,N_2777);
nand U2827 (N_2827,N_2763,N_2785);
nor U2828 (N_2828,N_2792,N_2761);
xnor U2829 (N_2829,N_2795,N_2799);
and U2830 (N_2830,N_2764,N_2760);
xor U2831 (N_2831,N_2788,N_2783);
and U2832 (N_2832,N_2802,N_2797);
nor U2833 (N_2833,N_2803,N_2787);
or U2834 (N_2834,N_2798,N_2778);
xor U2835 (N_2835,N_2768,N_2813);
nand U2836 (N_2836,N_2784,N_2814);
and U2837 (N_2837,N_2762,N_2767);
xor U2838 (N_2838,N_2818,N_2769);
nand U2839 (N_2839,N_2796,N_2772);
nor U2840 (N_2840,N_2766,N_2817);
xor U2841 (N_2841,N_2819,N_2782);
nand U2842 (N_2842,N_2790,N_2773);
nand U2843 (N_2843,N_2816,N_2806);
nor U2844 (N_2844,N_2774,N_2805);
xnor U2845 (N_2845,N_2779,N_2776);
or U2846 (N_2846,N_2789,N_2809);
nand U2847 (N_2847,N_2770,N_2812);
nand U2848 (N_2848,N_2794,N_2801);
xor U2849 (N_2849,N_2804,N_2811);
and U2850 (N_2850,N_2805,N_2803);
and U2851 (N_2851,N_2772,N_2794);
xnor U2852 (N_2852,N_2778,N_2797);
and U2853 (N_2853,N_2799,N_2798);
xor U2854 (N_2854,N_2788,N_2804);
or U2855 (N_2855,N_2771,N_2800);
xor U2856 (N_2856,N_2783,N_2789);
and U2857 (N_2857,N_2800,N_2807);
nor U2858 (N_2858,N_2760,N_2801);
or U2859 (N_2859,N_2802,N_2801);
nor U2860 (N_2860,N_2819,N_2767);
or U2861 (N_2861,N_2802,N_2789);
nor U2862 (N_2862,N_2780,N_2785);
xor U2863 (N_2863,N_2812,N_2796);
or U2864 (N_2864,N_2810,N_2807);
nor U2865 (N_2865,N_2783,N_2813);
or U2866 (N_2866,N_2765,N_2762);
or U2867 (N_2867,N_2792,N_2763);
nand U2868 (N_2868,N_2784,N_2782);
nor U2869 (N_2869,N_2802,N_2815);
nand U2870 (N_2870,N_2764,N_2799);
nor U2871 (N_2871,N_2763,N_2789);
and U2872 (N_2872,N_2768,N_2783);
xnor U2873 (N_2873,N_2791,N_2773);
nand U2874 (N_2874,N_2783,N_2801);
or U2875 (N_2875,N_2816,N_2797);
nor U2876 (N_2876,N_2760,N_2784);
and U2877 (N_2877,N_2792,N_2782);
nor U2878 (N_2878,N_2816,N_2795);
nor U2879 (N_2879,N_2773,N_2811);
and U2880 (N_2880,N_2857,N_2875);
and U2881 (N_2881,N_2842,N_2863);
nand U2882 (N_2882,N_2858,N_2850);
and U2883 (N_2883,N_2820,N_2864);
nor U2884 (N_2884,N_2832,N_2862);
or U2885 (N_2885,N_2821,N_2877);
nand U2886 (N_2886,N_2853,N_2855);
nand U2887 (N_2887,N_2823,N_2840);
and U2888 (N_2888,N_2865,N_2848);
xnor U2889 (N_2889,N_2871,N_2868);
or U2890 (N_2890,N_2867,N_2860);
or U2891 (N_2891,N_2849,N_2839);
xor U2892 (N_2892,N_2831,N_2835);
nor U2893 (N_2893,N_2845,N_2829);
and U2894 (N_2894,N_2879,N_2834);
or U2895 (N_2895,N_2836,N_2870);
nor U2896 (N_2896,N_2861,N_2843);
or U2897 (N_2897,N_2824,N_2869);
or U2898 (N_2898,N_2846,N_2866);
and U2899 (N_2899,N_2825,N_2852);
and U2900 (N_2900,N_2833,N_2830);
nand U2901 (N_2901,N_2851,N_2874);
nand U2902 (N_2902,N_2859,N_2872);
and U2903 (N_2903,N_2822,N_2856);
nor U2904 (N_2904,N_2873,N_2854);
or U2905 (N_2905,N_2826,N_2837);
or U2906 (N_2906,N_2838,N_2847);
or U2907 (N_2907,N_2841,N_2828);
nand U2908 (N_2908,N_2876,N_2878);
nor U2909 (N_2909,N_2827,N_2844);
or U2910 (N_2910,N_2863,N_2822);
xnor U2911 (N_2911,N_2830,N_2837);
and U2912 (N_2912,N_2869,N_2850);
nand U2913 (N_2913,N_2847,N_2844);
nand U2914 (N_2914,N_2879,N_2876);
nand U2915 (N_2915,N_2863,N_2869);
nand U2916 (N_2916,N_2875,N_2876);
or U2917 (N_2917,N_2825,N_2831);
and U2918 (N_2918,N_2857,N_2867);
or U2919 (N_2919,N_2848,N_2862);
xnor U2920 (N_2920,N_2850,N_2833);
nor U2921 (N_2921,N_2870,N_2852);
xnor U2922 (N_2922,N_2879,N_2854);
nor U2923 (N_2923,N_2856,N_2851);
nor U2924 (N_2924,N_2853,N_2844);
nor U2925 (N_2925,N_2871,N_2842);
or U2926 (N_2926,N_2851,N_2870);
nand U2927 (N_2927,N_2863,N_2835);
or U2928 (N_2928,N_2845,N_2839);
nor U2929 (N_2929,N_2826,N_2850);
and U2930 (N_2930,N_2876,N_2855);
and U2931 (N_2931,N_2853,N_2837);
or U2932 (N_2932,N_2877,N_2837);
xor U2933 (N_2933,N_2842,N_2827);
nor U2934 (N_2934,N_2865,N_2870);
and U2935 (N_2935,N_2821,N_2827);
nor U2936 (N_2936,N_2820,N_2875);
and U2937 (N_2937,N_2875,N_2873);
nand U2938 (N_2938,N_2846,N_2860);
nand U2939 (N_2939,N_2863,N_2866);
xnor U2940 (N_2940,N_2891,N_2924);
nor U2941 (N_2941,N_2911,N_2914);
xor U2942 (N_2942,N_2921,N_2884);
or U2943 (N_2943,N_2913,N_2912);
xnor U2944 (N_2944,N_2920,N_2935);
nand U2945 (N_2945,N_2904,N_2929);
and U2946 (N_2946,N_2918,N_2881);
nor U2947 (N_2947,N_2932,N_2909);
xnor U2948 (N_2948,N_2936,N_2925);
or U2949 (N_2949,N_2926,N_2907);
or U2950 (N_2950,N_2880,N_2903);
xor U2951 (N_2951,N_2886,N_2922);
and U2952 (N_2952,N_2899,N_2895);
or U2953 (N_2953,N_2908,N_2923);
or U2954 (N_2954,N_2892,N_2893);
and U2955 (N_2955,N_2930,N_2902);
or U2956 (N_2956,N_2896,N_2939);
nor U2957 (N_2957,N_2917,N_2938);
nor U2958 (N_2958,N_2900,N_2905);
and U2959 (N_2959,N_2937,N_2933);
or U2960 (N_2960,N_2916,N_2897);
or U2961 (N_2961,N_2919,N_2894);
or U2962 (N_2962,N_2885,N_2898);
nand U2963 (N_2963,N_2934,N_2927);
or U2964 (N_2964,N_2906,N_2910);
nand U2965 (N_2965,N_2928,N_2888);
and U2966 (N_2966,N_2890,N_2915);
and U2967 (N_2967,N_2882,N_2901);
nor U2968 (N_2968,N_2889,N_2931);
xnor U2969 (N_2969,N_2887,N_2883);
nand U2970 (N_2970,N_2928,N_2931);
and U2971 (N_2971,N_2900,N_2889);
xnor U2972 (N_2972,N_2910,N_2909);
xnor U2973 (N_2973,N_2919,N_2937);
nand U2974 (N_2974,N_2928,N_2897);
xnor U2975 (N_2975,N_2939,N_2892);
and U2976 (N_2976,N_2886,N_2907);
or U2977 (N_2977,N_2937,N_2917);
and U2978 (N_2978,N_2908,N_2933);
nand U2979 (N_2979,N_2884,N_2898);
nor U2980 (N_2980,N_2884,N_2937);
nor U2981 (N_2981,N_2912,N_2899);
nor U2982 (N_2982,N_2929,N_2907);
or U2983 (N_2983,N_2924,N_2925);
xnor U2984 (N_2984,N_2898,N_2909);
and U2985 (N_2985,N_2904,N_2901);
or U2986 (N_2986,N_2883,N_2896);
and U2987 (N_2987,N_2891,N_2884);
nand U2988 (N_2988,N_2922,N_2895);
nor U2989 (N_2989,N_2900,N_2880);
nor U2990 (N_2990,N_2891,N_2935);
xnor U2991 (N_2991,N_2904,N_2895);
nand U2992 (N_2992,N_2924,N_2928);
and U2993 (N_2993,N_2920,N_2938);
nor U2994 (N_2994,N_2923,N_2939);
xor U2995 (N_2995,N_2908,N_2935);
nand U2996 (N_2996,N_2904,N_2905);
or U2997 (N_2997,N_2886,N_2935);
nand U2998 (N_2998,N_2895,N_2928);
and U2999 (N_2999,N_2912,N_2886);
or UO_0 (O_0,N_2966,N_2979);
nor UO_1 (O_1,N_2950,N_2991);
xor UO_2 (O_2,N_2975,N_2952);
nand UO_3 (O_3,N_2980,N_2972);
or UO_4 (O_4,N_2948,N_2993);
and UO_5 (O_5,N_2974,N_2996);
and UO_6 (O_6,N_2946,N_2963);
or UO_7 (O_7,N_2973,N_2970);
and UO_8 (O_8,N_2951,N_2978);
or UO_9 (O_9,N_2997,N_2988);
xnor UO_10 (O_10,N_2940,N_2945);
nor UO_11 (O_11,N_2985,N_2986);
and UO_12 (O_12,N_2990,N_2943);
nor UO_13 (O_13,N_2983,N_2965);
and UO_14 (O_14,N_2969,N_2954);
nand UO_15 (O_15,N_2994,N_2962);
and UO_16 (O_16,N_2949,N_2998);
or UO_17 (O_17,N_2959,N_2956);
nor UO_18 (O_18,N_2942,N_2968);
nor UO_19 (O_19,N_2989,N_2995);
and UO_20 (O_20,N_2941,N_2967);
xor UO_21 (O_21,N_2984,N_2947);
xnor UO_22 (O_22,N_2960,N_2999);
and UO_23 (O_23,N_2992,N_2961);
xnor UO_24 (O_24,N_2987,N_2981);
xnor UO_25 (O_25,N_2955,N_2958);
or UO_26 (O_26,N_2976,N_2977);
or UO_27 (O_27,N_2982,N_2964);
xor UO_28 (O_28,N_2971,N_2957);
and UO_29 (O_29,N_2953,N_2944);
xnor UO_30 (O_30,N_2959,N_2980);
and UO_31 (O_31,N_2943,N_2997);
and UO_32 (O_32,N_2994,N_2945);
or UO_33 (O_33,N_2991,N_2993);
nor UO_34 (O_34,N_2973,N_2948);
nor UO_35 (O_35,N_2977,N_2983);
xnor UO_36 (O_36,N_2965,N_2981);
nand UO_37 (O_37,N_2979,N_2957);
nand UO_38 (O_38,N_2960,N_2953);
nand UO_39 (O_39,N_2941,N_2985);
nor UO_40 (O_40,N_2943,N_2963);
and UO_41 (O_41,N_2994,N_2964);
nand UO_42 (O_42,N_2941,N_2953);
xor UO_43 (O_43,N_2987,N_2970);
and UO_44 (O_44,N_2966,N_2965);
and UO_45 (O_45,N_2993,N_2976);
and UO_46 (O_46,N_2948,N_2949);
nor UO_47 (O_47,N_2998,N_2967);
xnor UO_48 (O_48,N_2990,N_2954);
or UO_49 (O_49,N_2964,N_2984);
nand UO_50 (O_50,N_2948,N_2987);
xnor UO_51 (O_51,N_2953,N_2995);
nand UO_52 (O_52,N_2953,N_2959);
xor UO_53 (O_53,N_2987,N_2973);
and UO_54 (O_54,N_2965,N_2984);
nand UO_55 (O_55,N_2992,N_2946);
and UO_56 (O_56,N_2948,N_2990);
nor UO_57 (O_57,N_2957,N_2973);
and UO_58 (O_58,N_2962,N_2989);
and UO_59 (O_59,N_2959,N_2942);
xor UO_60 (O_60,N_2969,N_2985);
and UO_61 (O_61,N_2971,N_2965);
or UO_62 (O_62,N_2940,N_2947);
nand UO_63 (O_63,N_2987,N_2953);
xnor UO_64 (O_64,N_2947,N_2970);
xnor UO_65 (O_65,N_2995,N_2959);
nand UO_66 (O_66,N_2995,N_2963);
xor UO_67 (O_67,N_2967,N_2960);
nand UO_68 (O_68,N_2993,N_2973);
xor UO_69 (O_69,N_2976,N_2957);
or UO_70 (O_70,N_2978,N_2958);
and UO_71 (O_71,N_2988,N_2958);
nand UO_72 (O_72,N_2946,N_2970);
xor UO_73 (O_73,N_2970,N_2949);
and UO_74 (O_74,N_2946,N_2983);
nor UO_75 (O_75,N_2945,N_2965);
nor UO_76 (O_76,N_2961,N_2943);
nand UO_77 (O_77,N_2977,N_2942);
nand UO_78 (O_78,N_2967,N_2976);
nor UO_79 (O_79,N_2958,N_2983);
or UO_80 (O_80,N_2995,N_2988);
or UO_81 (O_81,N_2959,N_2947);
and UO_82 (O_82,N_2952,N_2996);
or UO_83 (O_83,N_2993,N_2975);
nand UO_84 (O_84,N_2947,N_2978);
nor UO_85 (O_85,N_2974,N_2971);
nor UO_86 (O_86,N_2940,N_2965);
or UO_87 (O_87,N_2997,N_2990);
xnor UO_88 (O_88,N_2964,N_2975);
and UO_89 (O_89,N_2943,N_2995);
nor UO_90 (O_90,N_2964,N_2941);
nand UO_91 (O_91,N_2950,N_2960);
nand UO_92 (O_92,N_2990,N_2996);
and UO_93 (O_93,N_2980,N_2955);
nor UO_94 (O_94,N_2995,N_2993);
nand UO_95 (O_95,N_2991,N_2967);
xor UO_96 (O_96,N_2957,N_2972);
or UO_97 (O_97,N_2952,N_2964);
nand UO_98 (O_98,N_2971,N_2949);
nand UO_99 (O_99,N_2995,N_2977);
and UO_100 (O_100,N_2957,N_2962);
and UO_101 (O_101,N_2945,N_2955);
or UO_102 (O_102,N_2992,N_2971);
and UO_103 (O_103,N_2977,N_2965);
xnor UO_104 (O_104,N_2969,N_2997);
and UO_105 (O_105,N_2953,N_2961);
xnor UO_106 (O_106,N_2994,N_2972);
and UO_107 (O_107,N_2966,N_2943);
or UO_108 (O_108,N_2981,N_2972);
or UO_109 (O_109,N_2967,N_2974);
xnor UO_110 (O_110,N_2986,N_2947);
xnor UO_111 (O_111,N_2987,N_2963);
nor UO_112 (O_112,N_2960,N_2972);
nor UO_113 (O_113,N_2949,N_2997);
and UO_114 (O_114,N_2985,N_2954);
xnor UO_115 (O_115,N_2989,N_2966);
nor UO_116 (O_116,N_2976,N_2971);
nor UO_117 (O_117,N_2974,N_2966);
nor UO_118 (O_118,N_2971,N_2993);
or UO_119 (O_119,N_2955,N_2988);
xnor UO_120 (O_120,N_2943,N_2996);
xnor UO_121 (O_121,N_2959,N_2973);
nor UO_122 (O_122,N_2969,N_2996);
nor UO_123 (O_123,N_2948,N_2983);
xor UO_124 (O_124,N_2984,N_2960);
xor UO_125 (O_125,N_2957,N_2994);
and UO_126 (O_126,N_2965,N_2964);
nor UO_127 (O_127,N_2945,N_2954);
and UO_128 (O_128,N_2949,N_2991);
xor UO_129 (O_129,N_2956,N_2980);
xor UO_130 (O_130,N_2950,N_2985);
nand UO_131 (O_131,N_2965,N_2970);
nor UO_132 (O_132,N_2970,N_2971);
and UO_133 (O_133,N_2974,N_2944);
or UO_134 (O_134,N_2944,N_2972);
or UO_135 (O_135,N_2950,N_2975);
nand UO_136 (O_136,N_2980,N_2981);
xor UO_137 (O_137,N_2943,N_2949);
and UO_138 (O_138,N_2996,N_2988);
or UO_139 (O_139,N_2954,N_2956);
nand UO_140 (O_140,N_2963,N_2974);
and UO_141 (O_141,N_2957,N_2980);
and UO_142 (O_142,N_2961,N_2985);
nand UO_143 (O_143,N_2944,N_2995);
nor UO_144 (O_144,N_2967,N_2943);
or UO_145 (O_145,N_2984,N_2978);
nand UO_146 (O_146,N_2949,N_2952);
and UO_147 (O_147,N_2988,N_2950);
nor UO_148 (O_148,N_2999,N_2965);
nor UO_149 (O_149,N_2958,N_2948);
or UO_150 (O_150,N_2975,N_2957);
or UO_151 (O_151,N_2982,N_2978);
or UO_152 (O_152,N_2973,N_2945);
nor UO_153 (O_153,N_2958,N_2968);
xor UO_154 (O_154,N_2986,N_2991);
or UO_155 (O_155,N_2966,N_2975);
and UO_156 (O_156,N_2943,N_2989);
and UO_157 (O_157,N_2981,N_2975);
and UO_158 (O_158,N_2987,N_2956);
nand UO_159 (O_159,N_2982,N_2998);
nand UO_160 (O_160,N_2993,N_2990);
nor UO_161 (O_161,N_2993,N_2957);
xnor UO_162 (O_162,N_2974,N_2993);
nor UO_163 (O_163,N_2972,N_2958);
and UO_164 (O_164,N_2977,N_2982);
xnor UO_165 (O_165,N_2957,N_2968);
nor UO_166 (O_166,N_2964,N_2945);
and UO_167 (O_167,N_2989,N_2967);
or UO_168 (O_168,N_2992,N_2953);
nor UO_169 (O_169,N_2965,N_2972);
nand UO_170 (O_170,N_2965,N_2950);
and UO_171 (O_171,N_2994,N_2970);
nor UO_172 (O_172,N_2964,N_2998);
xnor UO_173 (O_173,N_2990,N_2981);
xnor UO_174 (O_174,N_2951,N_2960);
xnor UO_175 (O_175,N_2958,N_2967);
or UO_176 (O_176,N_2978,N_2945);
nand UO_177 (O_177,N_2941,N_2970);
nand UO_178 (O_178,N_2986,N_2954);
or UO_179 (O_179,N_2941,N_2959);
and UO_180 (O_180,N_2963,N_2965);
nand UO_181 (O_181,N_2979,N_2949);
xor UO_182 (O_182,N_2954,N_2941);
nor UO_183 (O_183,N_2981,N_2950);
and UO_184 (O_184,N_2997,N_2965);
nor UO_185 (O_185,N_2971,N_2981);
xnor UO_186 (O_186,N_2949,N_2974);
xnor UO_187 (O_187,N_2942,N_2955);
and UO_188 (O_188,N_2970,N_2978);
nor UO_189 (O_189,N_2977,N_2957);
and UO_190 (O_190,N_2996,N_2944);
xor UO_191 (O_191,N_2978,N_2967);
and UO_192 (O_192,N_2969,N_2993);
xor UO_193 (O_193,N_2987,N_2960);
xnor UO_194 (O_194,N_2941,N_2980);
or UO_195 (O_195,N_2989,N_2941);
or UO_196 (O_196,N_2959,N_2967);
xor UO_197 (O_197,N_2999,N_2991);
xor UO_198 (O_198,N_2944,N_2988);
nand UO_199 (O_199,N_2993,N_2980);
xor UO_200 (O_200,N_2969,N_2951);
nor UO_201 (O_201,N_2953,N_2967);
and UO_202 (O_202,N_2965,N_2979);
nor UO_203 (O_203,N_2968,N_2999);
or UO_204 (O_204,N_2979,N_2958);
xnor UO_205 (O_205,N_2950,N_2947);
nand UO_206 (O_206,N_2993,N_2950);
and UO_207 (O_207,N_2979,N_2940);
or UO_208 (O_208,N_2967,N_2985);
nand UO_209 (O_209,N_2943,N_2946);
nor UO_210 (O_210,N_2982,N_2970);
nor UO_211 (O_211,N_2968,N_2956);
nor UO_212 (O_212,N_2953,N_2942);
and UO_213 (O_213,N_2964,N_2992);
or UO_214 (O_214,N_2974,N_2961);
and UO_215 (O_215,N_2996,N_2992);
xor UO_216 (O_216,N_2955,N_2975);
nand UO_217 (O_217,N_2971,N_2964);
and UO_218 (O_218,N_2978,N_2957);
or UO_219 (O_219,N_2990,N_2958);
or UO_220 (O_220,N_2958,N_2998);
xnor UO_221 (O_221,N_2944,N_2961);
xor UO_222 (O_222,N_2992,N_2972);
xor UO_223 (O_223,N_2952,N_2970);
and UO_224 (O_224,N_2946,N_2947);
nor UO_225 (O_225,N_2944,N_2945);
xor UO_226 (O_226,N_2966,N_2987);
nor UO_227 (O_227,N_2986,N_2952);
or UO_228 (O_228,N_2993,N_2961);
nor UO_229 (O_229,N_2950,N_2987);
nor UO_230 (O_230,N_2958,N_2999);
xor UO_231 (O_231,N_2990,N_2952);
or UO_232 (O_232,N_2989,N_2954);
xor UO_233 (O_233,N_2961,N_2970);
nor UO_234 (O_234,N_2968,N_2959);
xor UO_235 (O_235,N_2977,N_2985);
and UO_236 (O_236,N_2996,N_2957);
nand UO_237 (O_237,N_2941,N_2948);
xor UO_238 (O_238,N_2973,N_2969);
or UO_239 (O_239,N_2967,N_2949);
or UO_240 (O_240,N_2950,N_2996);
or UO_241 (O_241,N_2968,N_2977);
nor UO_242 (O_242,N_2974,N_2992);
xor UO_243 (O_243,N_2963,N_2942);
xnor UO_244 (O_244,N_2994,N_2981);
nand UO_245 (O_245,N_2975,N_2943);
nor UO_246 (O_246,N_2998,N_2971);
nand UO_247 (O_247,N_2966,N_2951);
and UO_248 (O_248,N_2956,N_2966);
and UO_249 (O_249,N_2971,N_2973);
xnor UO_250 (O_250,N_2982,N_2994);
nand UO_251 (O_251,N_2979,N_2964);
xor UO_252 (O_252,N_2975,N_2960);
nor UO_253 (O_253,N_2953,N_2952);
and UO_254 (O_254,N_2989,N_2958);
nor UO_255 (O_255,N_2980,N_2962);
xnor UO_256 (O_256,N_2962,N_2974);
and UO_257 (O_257,N_2961,N_2979);
nor UO_258 (O_258,N_2969,N_2972);
nand UO_259 (O_259,N_2970,N_2964);
and UO_260 (O_260,N_2969,N_2984);
or UO_261 (O_261,N_2941,N_2950);
xor UO_262 (O_262,N_2959,N_2969);
and UO_263 (O_263,N_2949,N_2960);
xor UO_264 (O_264,N_2954,N_2961);
xor UO_265 (O_265,N_2956,N_2973);
nor UO_266 (O_266,N_2945,N_2966);
and UO_267 (O_267,N_2957,N_2960);
xnor UO_268 (O_268,N_2967,N_2971);
nand UO_269 (O_269,N_2952,N_2984);
and UO_270 (O_270,N_2984,N_2957);
xor UO_271 (O_271,N_2976,N_2984);
or UO_272 (O_272,N_2961,N_2967);
nand UO_273 (O_273,N_2977,N_2959);
xor UO_274 (O_274,N_2999,N_2990);
and UO_275 (O_275,N_2975,N_2980);
nand UO_276 (O_276,N_2961,N_2984);
and UO_277 (O_277,N_2989,N_2940);
nand UO_278 (O_278,N_2967,N_2990);
xor UO_279 (O_279,N_2987,N_2985);
nor UO_280 (O_280,N_2974,N_2964);
nor UO_281 (O_281,N_2995,N_2999);
or UO_282 (O_282,N_2958,N_2942);
nor UO_283 (O_283,N_2946,N_2964);
nand UO_284 (O_284,N_2972,N_2991);
and UO_285 (O_285,N_2993,N_2951);
nand UO_286 (O_286,N_2982,N_2944);
nand UO_287 (O_287,N_2948,N_2978);
or UO_288 (O_288,N_2986,N_2940);
and UO_289 (O_289,N_2949,N_2953);
or UO_290 (O_290,N_2989,N_2993);
and UO_291 (O_291,N_2971,N_2941);
and UO_292 (O_292,N_2950,N_2946);
xnor UO_293 (O_293,N_2944,N_2998);
or UO_294 (O_294,N_2940,N_2943);
nand UO_295 (O_295,N_2957,N_2988);
and UO_296 (O_296,N_2942,N_2971);
or UO_297 (O_297,N_2965,N_2946);
and UO_298 (O_298,N_2969,N_2955);
or UO_299 (O_299,N_2943,N_2980);
nor UO_300 (O_300,N_2940,N_2959);
or UO_301 (O_301,N_2983,N_2996);
or UO_302 (O_302,N_2983,N_2981);
nor UO_303 (O_303,N_2966,N_2995);
nand UO_304 (O_304,N_2954,N_2943);
xnor UO_305 (O_305,N_2947,N_2968);
or UO_306 (O_306,N_2946,N_2941);
nand UO_307 (O_307,N_2966,N_2980);
nand UO_308 (O_308,N_2962,N_2940);
and UO_309 (O_309,N_2974,N_2968);
or UO_310 (O_310,N_2952,N_2980);
nor UO_311 (O_311,N_2954,N_2981);
and UO_312 (O_312,N_2969,N_2987);
xor UO_313 (O_313,N_2987,N_2975);
nor UO_314 (O_314,N_2989,N_2957);
nand UO_315 (O_315,N_2945,N_2983);
or UO_316 (O_316,N_2980,N_2984);
xor UO_317 (O_317,N_2949,N_2947);
nor UO_318 (O_318,N_2982,N_2952);
nand UO_319 (O_319,N_2943,N_2958);
and UO_320 (O_320,N_2943,N_2964);
and UO_321 (O_321,N_2967,N_2977);
nor UO_322 (O_322,N_2940,N_2968);
nand UO_323 (O_323,N_2977,N_2966);
or UO_324 (O_324,N_2955,N_2979);
or UO_325 (O_325,N_2940,N_2958);
xor UO_326 (O_326,N_2954,N_2940);
nand UO_327 (O_327,N_2942,N_2965);
and UO_328 (O_328,N_2959,N_2962);
nor UO_329 (O_329,N_2961,N_2951);
or UO_330 (O_330,N_2948,N_2967);
and UO_331 (O_331,N_2994,N_2953);
nand UO_332 (O_332,N_2995,N_2952);
nor UO_333 (O_333,N_2993,N_2996);
and UO_334 (O_334,N_2988,N_2967);
nor UO_335 (O_335,N_2959,N_2976);
nor UO_336 (O_336,N_2980,N_2958);
nor UO_337 (O_337,N_2990,N_2964);
xor UO_338 (O_338,N_2963,N_2966);
nand UO_339 (O_339,N_2964,N_2940);
or UO_340 (O_340,N_2963,N_2945);
nor UO_341 (O_341,N_2948,N_2988);
or UO_342 (O_342,N_2941,N_2960);
xnor UO_343 (O_343,N_2975,N_2949);
nor UO_344 (O_344,N_2965,N_2953);
or UO_345 (O_345,N_2985,N_2974);
nand UO_346 (O_346,N_2943,N_2981);
and UO_347 (O_347,N_2968,N_2989);
nor UO_348 (O_348,N_2979,N_2941);
or UO_349 (O_349,N_2945,N_2999);
and UO_350 (O_350,N_2958,N_2970);
xnor UO_351 (O_351,N_2999,N_2972);
nand UO_352 (O_352,N_2963,N_2968);
xnor UO_353 (O_353,N_2968,N_2992);
nand UO_354 (O_354,N_2979,N_2944);
xor UO_355 (O_355,N_2969,N_2988);
nor UO_356 (O_356,N_2946,N_2994);
xnor UO_357 (O_357,N_2994,N_2992);
or UO_358 (O_358,N_2974,N_2970);
and UO_359 (O_359,N_2961,N_2980);
nand UO_360 (O_360,N_2967,N_2965);
xnor UO_361 (O_361,N_2976,N_2998);
nor UO_362 (O_362,N_2961,N_2947);
or UO_363 (O_363,N_2991,N_2965);
nand UO_364 (O_364,N_2994,N_2960);
xnor UO_365 (O_365,N_2969,N_2950);
nand UO_366 (O_366,N_2991,N_2946);
nor UO_367 (O_367,N_2945,N_2976);
nand UO_368 (O_368,N_2959,N_2964);
nor UO_369 (O_369,N_2971,N_2963);
and UO_370 (O_370,N_2998,N_2975);
xor UO_371 (O_371,N_2987,N_2943);
xor UO_372 (O_372,N_2947,N_2985);
and UO_373 (O_373,N_2984,N_2945);
nand UO_374 (O_374,N_2991,N_2958);
nor UO_375 (O_375,N_2961,N_2976);
xnor UO_376 (O_376,N_2991,N_2966);
and UO_377 (O_377,N_2946,N_2985);
or UO_378 (O_378,N_2995,N_2978);
nor UO_379 (O_379,N_2980,N_2964);
nand UO_380 (O_380,N_2942,N_2972);
xnor UO_381 (O_381,N_2948,N_2970);
xnor UO_382 (O_382,N_2974,N_2946);
nand UO_383 (O_383,N_2946,N_2945);
and UO_384 (O_384,N_2960,N_2946);
nor UO_385 (O_385,N_2969,N_2999);
or UO_386 (O_386,N_2952,N_2973);
xnor UO_387 (O_387,N_2980,N_2946);
nor UO_388 (O_388,N_2991,N_2977);
nor UO_389 (O_389,N_2957,N_2982);
nand UO_390 (O_390,N_2998,N_2991);
xnor UO_391 (O_391,N_2946,N_2958);
nand UO_392 (O_392,N_2960,N_2995);
or UO_393 (O_393,N_2964,N_2949);
xnor UO_394 (O_394,N_2948,N_2971);
xnor UO_395 (O_395,N_2942,N_2981);
nor UO_396 (O_396,N_2985,N_2942);
and UO_397 (O_397,N_2976,N_2949);
and UO_398 (O_398,N_2977,N_2958);
xor UO_399 (O_399,N_2955,N_2992);
xnor UO_400 (O_400,N_2942,N_2964);
or UO_401 (O_401,N_2956,N_2999);
xor UO_402 (O_402,N_2986,N_2974);
nor UO_403 (O_403,N_2988,N_2946);
xor UO_404 (O_404,N_2997,N_2940);
or UO_405 (O_405,N_2981,N_2969);
nand UO_406 (O_406,N_2970,N_2951);
or UO_407 (O_407,N_2984,N_2944);
and UO_408 (O_408,N_2988,N_2999);
nand UO_409 (O_409,N_2997,N_2977);
or UO_410 (O_410,N_2986,N_2967);
nand UO_411 (O_411,N_2979,N_2995);
xnor UO_412 (O_412,N_2986,N_2944);
nand UO_413 (O_413,N_2946,N_2953);
nand UO_414 (O_414,N_2985,N_2982);
nor UO_415 (O_415,N_2963,N_2976);
or UO_416 (O_416,N_2986,N_2994);
and UO_417 (O_417,N_2979,N_2946);
nand UO_418 (O_418,N_2956,N_2981);
xor UO_419 (O_419,N_2968,N_2948);
xnor UO_420 (O_420,N_2976,N_2991);
and UO_421 (O_421,N_2955,N_2977);
or UO_422 (O_422,N_2952,N_2950);
nand UO_423 (O_423,N_2944,N_2968);
and UO_424 (O_424,N_2967,N_2956);
or UO_425 (O_425,N_2974,N_2995);
or UO_426 (O_426,N_2993,N_2956);
and UO_427 (O_427,N_2953,N_2999);
xor UO_428 (O_428,N_2964,N_2989);
nor UO_429 (O_429,N_2974,N_2942);
nand UO_430 (O_430,N_2948,N_2989);
nor UO_431 (O_431,N_2999,N_2974);
xnor UO_432 (O_432,N_2957,N_2943);
or UO_433 (O_433,N_2949,N_2994);
nand UO_434 (O_434,N_2995,N_2986);
nand UO_435 (O_435,N_2956,N_2952);
nand UO_436 (O_436,N_2987,N_2997);
xor UO_437 (O_437,N_2960,N_2944);
or UO_438 (O_438,N_2979,N_2992);
xor UO_439 (O_439,N_2957,N_2965);
or UO_440 (O_440,N_2982,N_2981);
and UO_441 (O_441,N_2955,N_2989);
nor UO_442 (O_442,N_2956,N_2970);
nor UO_443 (O_443,N_2986,N_2949);
xor UO_444 (O_444,N_2995,N_2996);
and UO_445 (O_445,N_2949,N_2985);
xnor UO_446 (O_446,N_2941,N_2962);
or UO_447 (O_447,N_2973,N_2976);
xor UO_448 (O_448,N_2940,N_2998);
and UO_449 (O_449,N_2982,N_2953);
nor UO_450 (O_450,N_2993,N_2946);
nor UO_451 (O_451,N_2941,N_2978);
nor UO_452 (O_452,N_2975,N_2940);
and UO_453 (O_453,N_2972,N_2964);
or UO_454 (O_454,N_2946,N_2969);
xnor UO_455 (O_455,N_2993,N_2964);
or UO_456 (O_456,N_2989,N_2976);
nand UO_457 (O_457,N_2950,N_2956);
xor UO_458 (O_458,N_2958,N_2953);
or UO_459 (O_459,N_2977,N_2947);
and UO_460 (O_460,N_2954,N_2979);
and UO_461 (O_461,N_2991,N_2997);
or UO_462 (O_462,N_2980,N_2949);
or UO_463 (O_463,N_2977,N_2952);
and UO_464 (O_464,N_2971,N_2956);
nor UO_465 (O_465,N_2960,N_2956);
or UO_466 (O_466,N_2946,N_2967);
nand UO_467 (O_467,N_2949,N_2977);
or UO_468 (O_468,N_2945,N_2952);
nand UO_469 (O_469,N_2954,N_2970);
or UO_470 (O_470,N_2998,N_2984);
and UO_471 (O_471,N_2964,N_2955);
and UO_472 (O_472,N_2997,N_2993);
nor UO_473 (O_473,N_2963,N_2981);
and UO_474 (O_474,N_2969,N_2998);
nand UO_475 (O_475,N_2968,N_2983);
nor UO_476 (O_476,N_2958,N_2954);
or UO_477 (O_477,N_2984,N_2981);
and UO_478 (O_478,N_2982,N_2986);
and UO_479 (O_479,N_2994,N_2995);
nand UO_480 (O_480,N_2945,N_2968);
and UO_481 (O_481,N_2990,N_2969);
nand UO_482 (O_482,N_2966,N_2947);
or UO_483 (O_483,N_2958,N_2960);
and UO_484 (O_484,N_2971,N_2954);
nor UO_485 (O_485,N_2966,N_2959);
xor UO_486 (O_486,N_2972,N_2987);
and UO_487 (O_487,N_2997,N_2944);
nand UO_488 (O_488,N_2990,N_2975);
nor UO_489 (O_489,N_2950,N_2990);
nor UO_490 (O_490,N_2990,N_2991);
xnor UO_491 (O_491,N_2960,N_2969);
and UO_492 (O_492,N_2984,N_2967);
or UO_493 (O_493,N_2963,N_2975);
nand UO_494 (O_494,N_2957,N_2970);
or UO_495 (O_495,N_2974,N_2973);
or UO_496 (O_496,N_2993,N_2992);
nand UO_497 (O_497,N_2959,N_2961);
nand UO_498 (O_498,N_2999,N_2946);
and UO_499 (O_499,N_2950,N_2984);
endmodule