module basic_1500_15000_2000_120_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_1140,In_59);
xor U1 (N_1,In_316,In_170);
or U2 (N_2,In_79,In_738);
nor U3 (N_3,In_551,In_493);
nor U4 (N_4,In_305,In_436);
nand U5 (N_5,In_669,In_1320);
xor U6 (N_6,In_1378,In_652);
nor U7 (N_7,In_573,In_877);
nand U8 (N_8,In_293,In_169);
nand U9 (N_9,In_354,In_654);
nand U10 (N_10,In_905,In_484);
nand U11 (N_11,In_275,In_350);
and U12 (N_12,In_308,In_1168);
or U13 (N_13,In_796,In_158);
and U14 (N_14,In_247,In_1091);
xnor U15 (N_15,In_1055,In_1054);
or U16 (N_16,In_632,In_1072);
nand U17 (N_17,In_506,In_115);
nor U18 (N_18,In_945,In_580);
and U19 (N_19,In_181,In_581);
or U20 (N_20,In_596,In_613);
or U21 (N_21,In_163,In_872);
xnor U22 (N_22,In_427,In_1487);
xor U23 (N_23,In_457,In_1462);
xor U24 (N_24,In_880,In_1275);
nand U25 (N_25,In_698,In_235);
nor U26 (N_26,In_629,In_263);
nor U27 (N_27,In_579,In_1131);
xnor U28 (N_28,In_360,In_385);
and U29 (N_29,In_448,In_672);
and U30 (N_30,In_641,In_783);
xor U31 (N_31,In_98,In_812);
nand U32 (N_32,In_836,In_37);
and U33 (N_33,In_1496,In_352);
or U34 (N_34,In_392,In_219);
nand U35 (N_35,In_1143,In_696);
or U36 (N_36,In_482,In_31);
xnor U37 (N_37,In_110,In_324);
or U38 (N_38,In_1115,In_398);
or U39 (N_39,In_1481,In_97);
and U40 (N_40,In_546,In_1337);
nor U41 (N_41,In_881,In_186);
and U42 (N_42,In_676,In_1263);
or U43 (N_43,In_847,In_1355);
nor U44 (N_44,In_1228,In_931);
and U45 (N_45,In_1004,In_44);
or U46 (N_46,In_524,In_1379);
or U47 (N_47,In_520,In_375);
nor U48 (N_48,In_1293,In_1157);
or U49 (N_49,In_1229,In_96);
xnor U50 (N_50,In_1443,In_148);
xor U51 (N_51,In_887,In_374);
xnor U52 (N_52,In_675,In_1284);
nor U53 (N_53,In_1221,In_401);
nor U54 (N_54,In_825,In_509);
nor U55 (N_55,In_198,In_1136);
or U56 (N_56,In_917,In_902);
and U57 (N_57,In_954,In_1213);
nand U58 (N_58,In_190,In_963);
nand U59 (N_59,In_787,In_239);
or U60 (N_60,In_707,In_1017);
and U61 (N_61,In_600,In_1303);
and U62 (N_62,In_777,In_863);
and U63 (N_63,In_1109,In_793);
and U64 (N_64,In_1094,In_936);
or U65 (N_65,In_1068,In_538);
or U66 (N_66,In_1483,In_1190);
nand U67 (N_67,In_666,In_764);
xnor U68 (N_68,In_145,In_737);
nand U69 (N_69,In_842,In_471);
or U70 (N_70,In_107,In_1311);
and U71 (N_71,In_477,In_1251);
nor U72 (N_72,In_1458,In_495);
and U73 (N_73,In_1286,In_334);
nor U74 (N_74,In_161,In_194);
nor U75 (N_75,In_1291,In_257);
nand U76 (N_76,In_390,In_1063);
or U77 (N_77,In_588,In_333);
nand U78 (N_78,In_1045,In_1051);
nand U79 (N_79,In_655,In_1012);
nor U80 (N_80,In_1093,In_1202);
or U81 (N_81,In_1319,In_1002);
and U82 (N_82,In_1475,In_307);
and U83 (N_83,In_47,In_1267);
nand U84 (N_84,In_775,In_1048);
nand U85 (N_85,In_911,In_95);
and U86 (N_86,In_261,In_1405);
xnor U87 (N_87,In_713,In_41);
or U88 (N_88,In_871,In_1220);
nand U89 (N_89,In_1135,In_1150);
or U90 (N_90,In_590,In_785);
or U91 (N_91,In_1078,In_172);
nor U92 (N_92,In_949,In_970);
or U93 (N_93,In_356,In_941);
nand U94 (N_94,In_802,In_202);
xnor U95 (N_95,In_1359,In_1420);
nor U96 (N_96,In_1246,In_1301);
or U97 (N_97,In_1421,In_1389);
and U98 (N_98,In_1075,In_761);
xnor U99 (N_99,In_743,In_790);
and U100 (N_100,In_922,In_755);
xnor U101 (N_101,In_1008,In_810);
xnor U102 (N_102,In_1398,In_772);
xnor U103 (N_103,In_688,In_1231);
xnor U104 (N_104,In_822,In_187);
nor U105 (N_105,In_921,In_1375);
nor U106 (N_106,In_684,In_742);
or U107 (N_107,In_1428,In_665);
or U108 (N_108,In_497,In_1290);
nor U109 (N_109,In_1488,In_971);
xor U110 (N_110,In_1025,In_725);
or U111 (N_111,In_394,In_109);
or U112 (N_112,In_719,In_301);
or U113 (N_113,In_1167,In_164);
nand U114 (N_114,In_25,In_1262);
xor U115 (N_115,In_824,In_55);
nor U116 (N_116,In_266,In_953);
nand U117 (N_117,In_80,In_1189);
or U118 (N_118,In_204,In_1226);
and U119 (N_119,In_607,In_150);
or U120 (N_120,In_171,In_1088);
or U121 (N_121,In_991,In_965);
nor U122 (N_122,In_1219,In_1384);
or U123 (N_123,In_259,In_1186);
xnor U124 (N_124,In_1036,In_1418);
or U125 (N_125,In_623,In_1181);
and U126 (N_126,In_1423,In_8);
or U127 (N_127,In_69,N_16);
nand U128 (N_128,In_144,In_421);
xor U129 (N_129,In_1438,N_62);
xnor U130 (N_130,In_433,N_77);
nor U131 (N_131,N_122,In_536);
and U132 (N_132,In_1408,N_28);
or U133 (N_133,In_814,In_211);
and U134 (N_134,In_1486,In_1411);
and U135 (N_135,In_18,In_503);
or U136 (N_136,N_17,In_463);
nand U137 (N_137,N_0,In_203);
xnor U138 (N_138,In_856,In_1225);
xor U139 (N_139,In_1372,N_63);
nor U140 (N_140,In_1436,In_693);
and U141 (N_141,In_1125,In_434);
nor U142 (N_142,In_1374,In_156);
nand U143 (N_143,N_7,In_870);
xor U144 (N_144,In_313,In_1138);
or U145 (N_145,In_231,In_347);
nor U146 (N_146,N_114,In_658);
nor U147 (N_147,In_1383,N_33);
and U148 (N_148,In_1322,In_254);
nand U149 (N_149,In_391,In_0);
nand U150 (N_150,In_56,In_1050);
and U151 (N_151,In_1193,In_136);
xnor U152 (N_152,In_48,In_1349);
nand U153 (N_153,In_90,N_109);
nor U154 (N_154,In_748,In_1092);
and U155 (N_155,In_185,In_129);
nor U156 (N_156,In_1159,In_1201);
or U157 (N_157,In_544,In_660);
nor U158 (N_158,In_1027,In_205);
nand U159 (N_159,In_166,In_1172);
or U160 (N_160,In_1010,In_567);
nand U161 (N_161,In_1477,In_253);
and U162 (N_162,In_75,In_319);
or U163 (N_163,In_1195,In_915);
nor U164 (N_164,In_816,N_106);
xnor U165 (N_165,In_232,In_1282);
nor U166 (N_166,In_1313,In_1204);
nor U167 (N_167,In_677,In_889);
and U168 (N_168,In_66,In_680);
nand U169 (N_169,N_96,N_37);
and U170 (N_170,In_657,In_1142);
or U171 (N_171,N_93,In_376);
or U172 (N_172,In_472,In_1234);
and U173 (N_173,In_982,In_966);
and U174 (N_174,In_568,In_387);
and U175 (N_175,In_972,In_1214);
or U176 (N_176,In_592,In_1403);
nand U177 (N_177,N_58,In_20);
xor U178 (N_178,In_828,In_890);
nand U179 (N_179,In_687,In_673);
nand U180 (N_180,In_711,In_282);
and U181 (N_181,In_426,In_1070);
and U182 (N_182,In_106,In_516);
and U183 (N_183,In_769,In_64);
xor U184 (N_184,In_1060,In_786);
xnor U185 (N_185,In_1437,In_357);
xor U186 (N_186,In_28,In_1480);
xnor U187 (N_187,In_1454,In_326);
nor U188 (N_188,In_58,In_310);
and U189 (N_189,N_70,In_1028);
and U190 (N_190,In_771,In_882);
nor U191 (N_191,In_1256,In_746);
nor U192 (N_192,In_380,In_1241);
xor U193 (N_193,In_1067,In_1433);
nand U194 (N_194,In_1400,N_108);
nor U195 (N_195,In_691,In_992);
or U196 (N_196,In_1151,In_1169);
or U197 (N_197,In_1222,N_11);
nand U198 (N_198,In_479,In_303);
xor U199 (N_199,In_542,In_236);
nand U200 (N_200,In_429,In_1430);
or U201 (N_201,In_386,In_1388);
xor U202 (N_202,In_1310,In_33);
nand U203 (N_203,In_1118,In_645);
nand U204 (N_204,In_952,In_238);
and U205 (N_205,In_633,In_206);
or U206 (N_206,In_744,In_1264);
nand U207 (N_207,In_1132,In_1099);
nand U208 (N_208,In_1110,N_15);
nor U209 (N_209,In_900,In_1364);
and U210 (N_210,In_910,In_832);
or U211 (N_211,In_1001,In_1023);
xor U212 (N_212,In_859,In_745);
or U213 (N_213,In_42,In_736);
nand U214 (N_214,In_1120,In_1339);
nand U215 (N_215,In_1268,In_608);
nor U216 (N_216,In_1020,In_1367);
or U217 (N_217,In_138,In_1119);
xnor U218 (N_218,In_620,In_4);
nand U219 (N_219,In_218,In_296);
xor U220 (N_220,N_90,In_445);
xnor U221 (N_221,N_88,In_443);
and U222 (N_222,In_511,In_811);
and U223 (N_223,In_1305,In_1279);
xnor U224 (N_224,In_60,In_1197);
nand U225 (N_225,In_76,In_715);
and U226 (N_226,In_1484,N_56);
xnor U227 (N_227,In_476,N_97);
xnor U228 (N_228,In_1352,In_733);
or U229 (N_229,In_710,In_1258);
xor U230 (N_230,In_1216,In_1343);
nand U231 (N_231,In_605,In_312);
xnor U232 (N_232,In_425,N_103);
or U233 (N_233,In_1183,In_402);
nand U234 (N_234,In_1232,In_930);
and U235 (N_235,In_1162,In_819);
or U236 (N_236,In_656,In_121);
and U237 (N_237,In_1071,In_217);
and U238 (N_238,In_1250,In_286);
xor U239 (N_239,In_378,In_1495);
nor U240 (N_240,In_230,In_1425);
nand U241 (N_241,In_220,In_321);
nor U242 (N_242,In_1356,In_345);
or U243 (N_243,In_529,In_649);
xnor U244 (N_244,In_1331,In_749);
nor U245 (N_245,N_81,In_1327);
or U246 (N_246,N_34,In_679);
nor U247 (N_247,In_182,In_451);
xor U248 (N_248,In_29,In_639);
nand U249 (N_249,In_1106,In_40);
xor U250 (N_250,In_807,N_101);
nand U251 (N_251,In_291,In_740);
nor U252 (N_252,N_203,In_1321);
and U253 (N_253,N_59,In_265);
and U254 (N_254,In_1390,In_88);
nor U255 (N_255,In_420,N_173);
nor U256 (N_256,In_120,In_1435);
xnor U257 (N_257,In_984,In_1179);
nand U258 (N_258,In_726,In_1373);
nand U259 (N_259,N_84,In_770);
or U260 (N_260,N_228,N_66);
or U261 (N_261,N_140,N_112);
nor U262 (N_262,In_1451,In_722);
and U263 (N_263,In_617,In_1165);
nor U264 (N_264,In_1401,In_417);
and U265 (N_265,In_46,In_522);
nor U266 (N_266,N_78,In_1455);
nor U267 (N_267,In_139,N_230);
nor U268 (N_268,In_1368,In_983);
or U269 (N_269,In_1144,In_6);
and U270 (N_270,In_15,In_1399);
nor U271 (N_271,In_1380,In_1358);
xnor U272 (N_272,In_431,In_862);
or U273 (N_273,In_1126,In_974);
or U274 (N_274,In_852,In_1447);
or U275 (N_275,N_126,In_1215);
xor U276 (N_276,In_81,In_112);
nand U277 (N_277,In_188,In_125);
nand U278 (N_278,In_1182,In_1252);
nor U279 (N_279,In_1259,N_248);
xor U280 (N_280,In_835,In_1253);
nor U281 (N_281,In_944,In_450);
xnor U282 (N_282,In_1460,In_507);
or U283 (N_283,In_519,In_1328);
xnor U284 (N_284,In_388,In_967);
xnor U285 (N_285,In_858,N_113);
and U286 (N_286,In_184,In_1113);
or U287 (N_287,In_1049,In_728);
or U288 (N_288,In_716,In_10);
nor U289 (N_289,In_1345,In_874);
xor U290 (N_290,In_1160,In_937);
xor U291 (N_291,In_912,In_94);
nor U292 (N_292,In_885,In_16);
nand U293 (N_293,In_585,In_1471);
nand U294 (N_294,In_116,In_1416);
or U295 (N_295,In_703,In_24);
or U296 (N_296,In_299,In_1422);
nor U297 (N_297,In_845,In_789);
nand U298 (N_298,In_108,In_932);
or U299 (N_299,In_593,In_948);
nand U300 (N_300,N_160,In_651);
nand U301 (N_301,In_549,In_21);
nor U302 (N_302,In_844,In_798);
nor U303 (N_303,N_75,In_343);
or U304 (N_304,In_1090,In_1133);
xnor U305 (N_305,In_1130,In_36);
nand U306 (N_306,In_1344,In_1205);
nor U307 (N_307,N_225,In_1041);
xor U308 (N_308,In_1254,N_115);
nand U309 (N_309,N_170,N_129);
xnor U310 (N_310,In_1244,In_117);
nor U311 (N_311,In_78,In_779);
xnor U312 (N_312,N_169,In_1043);
and U313 (N_313,In_327,In_277);
or U314 (N_314,In_1414,N_190);
or U315 (N_315,In_126,In_1035);
nor U316 (N_316,In_782,In_208);
and U317 (N_317,In_616,In_829);
or U318 (N_318,In_734,In_153);
or U319 (N_319,In_404,In_653);
xnor U320 (N_320,N_57,In_207);
and U321 (N_321,In_504,In_701);
xor U322 (N_322,In_444,In_418);
or U323 (N_323,In_416,N_240);
or U324 (N_324,In_167,In_919);
or U325 (N_325,In_1489,N_164);
and U326 (N_326,In_1469,In_1276);
nand U327 (N_327,In_84,In_988);
and U328 (N_328,In_846,In_1185);
or U329 (N_329,In_1289,N_65);
nand U330 (N_330,In_980,In_256);
nor U331 (N_331,N_131,N_13);
or U332 (N_332,In_35,N_111);
nand U333 (N_333,In_353,In_1270);
nand U334 (N_334,In_997,In_987);
xnor U335 (N_335,In_951,In_712);
xnor U336 (N_336,In_876,In_499);
xor U337 (N_337,In_1209,N_76);
xor U338 (N_338,N_154,N_132);
or U339 (N_339,In_857,In_1314);
xor U340 (N_340,In_640,In_706);
xnor U341 (N_341,N_83,In_1180);
nor U342 (N_342,In_1040,In_827);
nor U343 (N_343,In_323,N_147);
xnor U344 (N_344,N_165,In_1192);
nand U345 (N_345,In_159,In_860);
or U346 (N_346,In_1248,In_280);
xnor U347 (N_347,In_68,In_621);
or U348 (N_348,In_381,In_1281);
xnor U349 (N_349,In_754,In_897);
nand U350 (N_350,In_552,N_245);
xor U351 (N_351,In_947,In_985);
nor U352 (N_352,In_582,In_916);
nand U353 (N_353,In_946,In_510);
nand U354 (N_354,In_234,In_1360);
and U355 (N_355,In_1003,N_124);
xnor U356 (N_356,In_780,In_689);
nand U357 (N_357,In_57,In_854);
xor U358 (N_358,In_1163,In_1274);
and U359 (N_359,In_867,In_584);
xor U360 (N_360,N_130,In_242);
or U361 (N_361,N_44,N_178);
nor U362 (N_362,In_470,In_285);
or U363 (N_363,In_1278,In_705);
nor U364 (N_364,In_1302,In_468);
and U365 (N_365,In_346,In_1312);
nand U366 (N_366,In_17,In_597);
xnor U367 (N_367,In_478,In_441);
nand U368 (N_368,In_309,In_413);
xnor U369 (N_369,In_214,N_208);
or U370 (N_370,In_1061,In_396);
or U371 (N_371,In_1152,In_1129);
xor U372 (N_372,In_1463,In_751);
or U373 (N_373,In_614,In_210);
or U374 (N_374,In_1357,In_1239);
xnor U375 (N_375,In_583,In_225);
or U376 (N_376,In_160,In_674);
nor U377 (N_377,In_270,N_110);
xor U378 (N_378,N_224,In_304);
nor U379 (N_379,N_215,In_704);
or U380 (N_380,In_646,In_1161);
nor U381 (N_381,In_851,In_678);
and U382 (N_382,In_791,In_1493);
or U383 (N_383,In_1304,N_287);
nand U384 (N_384,N_142,In_545);
nand U385 (N_385,In_572,In_1056);
and U386 (N_386,In_528,In_1300);
or U387 (N_387,In_1015,In_1081);
nor U388 (N_388,In_594,In_1194);
or U389 (N_389,In_1431,In_487);
xor U390 (N_390,In_694,N_214);
nor U391 (N_391,In_834,N_175);
and U392 (N_392,N_91,N_279);
nor U393 (N_393,In_759,N_123);
xor U394 (N_394,In_1376,In_795);
or U395 (N_395,In_393,In_1038);
xnor U396 (N_396,In_615,In_873);
or U397 (N_397,In_1086,N_171);
xor U398 (N_398,In_1295,In_473);
and U399 (N_399,N_260,In_561);
and U400 (N_400,N_22,In_27);
nand U401 (N_401,N_27,N_355);
and U402 (N_402,In_399,N_102);
nor U403 (N_403,In_535,In_907);
nand U404 (N_404,In_648,In_525);
nor U405 (N_405,In_661,In_730);
nor U406 (N_406,In_1464,N_237);
and U407 (N_407,In_492,N_273);
and U408 (N_408,In_636,In_363);
xnor U409 (N_409,N_212,In_197);
nor U410 (N_410,In_532,N_241);
xor U411 (N_411,In_395,N_285);
nor U412 (N_412,In_569,N_243);
nand U413 (N_413,N_48,In_1415);
xnor U414 (N_414,In_335,In_1325);
or U415 (N_415,N_369,N_21);
and U416 (N_416,In_447,In_1139);
or U417 (N_417,In_38,In_554);
or U418 (N_418,In_909,In_784);
xnor U419 (N_419,In_149,N_67);
or U420 (N_420,N_278,In_517);
nor U421 (N_421,N_367,In_1108);
nand U422 (N_422,In_630,In_1485);
xnor U423 (N_423,In_223,In_1176);
and U424 (N_424,N_153,In_273);
xnor U425 (N_425,N_326,N_211);
and U426 (N_426,In_142,In_539);
nand U427 (N_427,In_226,In_700);
and U428 (N_428,In_49,In_888);
or U429 (N_429,N_290,In_918);
nand U430 (N_430,In_833,In_864);
or U431 (N_431,In_54,N_182);
nor U432 (N_432,In_295,In_193);
nor U433 (N_433,In_776,N_29);
nor U434 (N_434,N_38,In_1184);
and U435 (N_435,In_818,In_1101);
nor U436 (N_436,N_301,In_837);
or U437 (N_437,N_52,In_1335);
xor U438 (N_438,In_514,In_1233);
and U439 (N_439,In_574,In_717);
nand U440 (N_440,In_475,In_1224);
nand U441 (N_441,N_309,In_955);
and U442 (N_442,In_1394,In_1333);
or U443 (N_443,In_644,In_1392);
and U444 (N_444,In_229,In_183);
or U445 (N_445,In_595,In_465);
xnor U446 (N_446,In_322,In_1297);
nor U447 (N_447,N_319,In_32);
or U448 (N_448,In_1097,In_879);
or U449 (N_449,N_333,In_663);
and U450 (N_450,In_808,In_279);
nor U451 (N_451,N_276,N_330);
nand U452 (N_452,In_367,In_875);
nor U453 (N_453,In_1391,In_1127);
nor U454 (N_454,N_133,In_320);
nand U455 (N_455,In_702,In_927);
nand U456 (N_456,In_70,N_137);
or U457 (N_457,In_1336,N_239);
xor U458 (N_458,N_100,In_1227);
and U459 (N_459,In_690,In_351);
nand U460 (N_460,N_216,N_255);
or U461 (N_461,In_1211,In_578);
xnor U462 (N_462,N_222,In_358);
or U463 (N_463,In_406,N_143);
nor U464 (N_464,In_591,In_865);
and U465 (N_465,N_352,In_709);
and U466 (N_466,In_1461,In_102);
and U467 (N_467,In_1011,In_1191);
nand U468 (N_468,In_1087,In_1217);
xor U469 (N_469,In_11,In_400);
and U470 (N_470,In_1404,In_720);
nor U471 (N_471,In_563,In_294);
and U472 (N_472,N_226,N_104);
or U473 (N_473,N_314,N_263);
and U474 (N_474,In_659,In_577);
or U475 (N_475,N_302,In_289);
nand U476 (N_476,In_603,In_222);
nand U477 (N_477,In_553,In_359);
and U478 (N_478,In_1065,N_292);
or U479 (N_479,In_1292,N_179);
nand U480 (N_480,N_282,In_337);
or U481 (N_481,In_855,In_389);
xor U482 (N_482,N_350,In_1153);
or U483 (N_483,N_189,In_422);
nand U484 (N_484,In_306,In_1188);
nand U485 (N_485,In_1288,N_336);
nand U486 (N_486,In_440,In_260);
nand U487 (N_487,In_276,In_23);
xor U488 (N_488,In_598,In_1257);
nor U489 (N_489,In_609,N_30);
or U490 (N_490,In_901,In_1385);
xor U491 (N_491,In_1069,In_575);
nor U492 (N_492,In_899,In_175);
or U493 (N_493,N_232,In_634);
nand U494 (N_494,N_156,In_372);
and U495 (N_495,N_299,N_151);
or U496 (N_496,In_841,In_799);
xor U497 (N_497,N_363,In_14);
xnor U498 (N_498,In_558,In_556);
and U499 (N_499,In_502,In_898);
nand U500 (N_500,N_328,In_466);
xnor U501 (N_501,N_289,In_1059);
and U502 (N_502,N_148,In_199);
xor U503 (N_503,In_348,N_139);
or U504 (N_504,N_424,N_427);
xnor U505 (N_505,In_1146,In_727);
nor U506 (N_506,N_271,In_43);
xor U507 (N_507,In_515,N_146);
or U508 (N_508,In_1426,N_387);
or U509 (N_509,N_294,N_50);
and U510 (N_510,N_428,In_1318);
or U511 (N_511,In_245,In_1424);
xnor U512 (N_512,In_1000,In_508);
xor U513 (N_513,N_217,In_449);
nor U514 (N_514,N_234,N_85);
nor U515 (N_515,N_196,In_100);
or U516 (N_516,N_341,In_368);
and U517 (N_517,In_39,N_411);
or U518 (N_518,N_9,In_849);
nand U519 (N_519,In_1114,In_438);
and U520 (N_520,In_505,In_1046);
and U521 (N_521,In_604,N_269);
and U522 (N_522,In_805,In_1137);
nand U523 (N_523,In_547,In_1166);
nor U524 (N_524,In_464,In_1442);
and U525 (N_525,N_322,In_1178);
nor U526 (N_526,In_1066,In_62);
and U527 (N_527,In_1448,In_332);
or U528 (N_528,In_1037,In_920);
and U529 (N_529,In_1309,In_1158);
nor U530 (N_530,In_92,N_210);
nor U531 (N_531,In_848,N_391);
nand U532 (N_532,In_494,In_228);
xnor U533 (N_533,In_72,N_24);
or U534 (N_534,N_462,In_248);
nand U535 (N_535,In_555,In_314);
nand U536 (N_536,In_5,N_457);
nand U537 (N_537,N_366,In_1307);
nor U538 (N_538,In_878,In_1174);
xnor U539 (N_539,In_1084,In_414);
or U540 (N_540,In_1402,In_361);
xnor U541 (N_541,N_470,In_1237);
or U542 (N_542,In_311,In_283);
nor U543 (N_543,In_365,N_150);
nand U544 (N_544,In_34,N_253);
nand U545 (N_545,N_445,N_406);
xor U546 (N_546,In_571,N_493);
or U547 (N_547,N_136,In_624);
and U548 (N_548,In_123,In_1468);
nor U549 (N_549,In_589,In_268);
nor U550 (N_550,In_397,In_1039);
or U551 (N_551,In_1315,N_310);
xnor U552 (N_552,In_255,In_1047);
and U553 (N_553,N_155,In_809);
xnor U554 (N_554,In_1124,In_896);
or U555 (N_555,In_140,In_405);
or U556 (N_556,In_1449,In_797);
and U557 (N_557,In_147,In_686);
and U558 (N_558,In_409,In_906);
or U559 (N_559,N_18,In_474);
nand U560 (N_560,In_883,In_1076);
xnor U561 (N_561,In_73,N_403);
nor U562 (N_562,In_1444,In_1338);
and U563 (N_563,N_329,In_959);
nand U564 (N_564,In_325,N_439);
or U565 (N_565,N_107,In_274);
and U566 (N_566,In_747,In_1112);
and U567 (N_567,In_246,N_236);
nand U568 (N_568,N_167,N_220);
and U569 (N_569,N_266,In_1260);
nor U570 (N_570,In_765,In_973);
nand U571 (N_571,In_766,N_256);
nor U572 (N_572,In_903,In_1353);
and U573 (N_573,In_87,In_180);
nor U574 (N_574,N_264,In_278);
nand U575 (N_575,In_1034,In_1294);
nand U576 (N_576,In_1324,In_767);
nor U577 (N_577,In_599,N_98);
and U578 (N_578,N_498,In_637);
xor U579 (N_579,In_272,In_1261);
nand U580 (N_580,N_79,N_473);
xor U581 (N_581,In_344,N_19);
xnor U582 (N_582,In_338,N_162);
xor U583 (N_583,N_413,N_368);
xor U584 (N_584,In_328,In_1243);
nor U585 (N_585,N_323,In_559);
nor U586 (N_586,In_1452,In_469);
xor U587 (N_587,In_2,In_960);
xnor U588 (N_588,In_566,In_1173);
xor U589 (N_589,In_292,N_456);
xnor U590 (N_590,In_1014,In_570);
xnor U591 (N_591,In_1095,In_962);
nand U592 (N_592,N_251,N_291);
or U593 (N_593,In_362,In_1013);
nand U594 (N_594,N_244,N_386);
or U595 (N_595,In_105,N_61);
nor U596 (N_596,In_801,N_334);
nand U597 (N_597,In_131,In_1351);
or U598 (N_598,N_349,N_379);
or U599 (N_599,N_324,N_486);
and U600 (N_600,N_202,N_40);
xor U601 (N_601,In_562,In_103);
nor U602 (N_602,In_77,In_750);
nor U603 (N_603,In_756,In_1033);
nand U604 (N_604,In_1198,In_647);
nor U605 (N_605,N_448,In_998);
nor U606 (N_606,In_412,N_375);
nand U607 (N_607,In_800,N_117);
nand U608 (N_608,In_1016,N_490);
nand U609 (N_609,N_267,In_1042);
xnor U610 (N_610,N_163,N_74);
nand U611 (N_611,In_803,In_1203);
and U612 (N_612,In_1265,N_2);
and U613 (N_613,In_699,In_530);
nor U614 (N_614,N_64,In_866);
xor U615 (N_615,N_1,N_268);
nand U616 (N_616,N_463,In_934);
xnor U617 (N_617,In_480,N_354);
nor U618 (N_618,In_1006,N_347);
or U619 (N_619,In_839,In_1134);
nor U620 (N_620,N_10,In_1235);
and U621 (N_621,N_80,In_1459);
nand U622 (N_622,N_311,N_423);
nor U623 (N_623,In_1240,In_1386);
nor U624 (N_624,In_868,In_155);
and U625 (N_625,N_398,In_667);
nor U626 (N_626,N_509,In_1369);
xnor U627 (N_627,In_1287,In_964);
nand U628 (N_628,In_215,In_1354);
and U629 (N_629,N_339,In_626);
and U630 (N_630,N_118,In_430);
nand U631 (N_631,In_1058,In_521);
nand U632 (N_632,In_462,In_86);
and U633 (N_633,In_224,In_1445);
xnor U634 (N_634,In_500,N_570);
xor U635 (N_635,In_978,N_573);
nor U636 (N_636,N_42,N_525);
nand U637 (N_637,In_284,N_180);
or U638 (N_638,N_53,N_344);
nor U639 (N_639,N_580,N_426);
or U640 (N_640,In_1107,N_152);
and U641 (N_641,N_622,N_261);
and U642 (N_642,In_723,N_316);
or U643 (N_643,In_297,In_1199);
xnor U644 (N_644,N_358,N_68);
xnor U645 (N_645,N_401,In_382);
xor U646 (N_646,In_1074,N_233);
or U647 (N_647,N_149,N_449);
nand U648 (N_648,In_52,In_612);
and U649 (N_649,In_958,In_82);
xnor U650 (N_650,N_589,N_527);
nand U651 (N_651,N_523,N_407);
nand U652 (N_652,N_205,N_177);
nor U653 (N_653,In_830,N_471);
nor U654 (N_654,In_1123,In_26);
and U655 (N_655,N_483,N_192);
nand U656 (N_656,In_1299,In_315);
and U657 (N_657,In_174,In_127);
nand U658 (N_658,N_528,In_1473);
or U659 (N_659,In_1406,In_1187);
and U660 (N_660,N_95,N_588);
nand U661 (N_661,In_113,N_204);
and U662 (N_662,In_773,In_1362);
and U663 (N_663,N_602,N_4);
xor U664 (N_664,In_152,In_735);
or U665 (N_665,N_176,N_599);
and U666 (N_666,N_158,In_134);
and U667 (N_667,In_1249,N_318);
or U668 (N_668,In_565,N_300);
nor U669 (N_669,In_638,N_105);
or U670 (N_670,N_547,N_385);
nor U671 (N_671,N_608,N_71);
nor U672 (N_672,In_586,N_469);
nand U673 (N_673,N_174,N_524);
and U674 (N_674,N_145,In_453);
nand U675 (N_675,In_428,In_1280);
nor U676 (N_676,In_240,N_86);
nand U677 (N_677,N_23,In_821);
nand U678 (N_678,N_331,N_458);
xnor U679 (N_679,In_501,In_695);
nand U680 (N_680,N_574,In_662);
xnor U681 (N_681,In_1341,In_7);
xnor U682 (N_682,N_46,N_561);
or U683 (N_683,N_436,N_560);
nand U684 (N_684,In_124,In_1330);
xnor U685 (N_685,In_891,In_192);
and U686 (N_686,In_1141,In_302);
xor U687 (N_687,In_1236,N_396);
nor U688 (N_688,In_969,In_1350);
xor U689 (N_689,N_418,In_1347);
nand U690 (N_690,N_197,N_194);
or U691 (N_691,In_119,N_519);
or U692 (N_692,In_165,N_348);
xnor U693 (N_693,In_1053,In_1456);
nand U694 (N_694,In_1323,In_895);
nor U695 (N_695,N_200,In_1147);
and U696 (N_696,In_1427,N_479);
xnor U697 (N_697,In_496,In_22);
nor U698 (N_698,N_571,In_377);
nand U699 (N_699,In_1326,In_370);
and U700 (N_700,N_501,N_601);
or U701 (N_701,N_534,In_439);
and U702 (N_702,N_572,In_461);
nand U703 (N_703,N_481,In_383);
nor U704 (N_704,In_1064,N_337);
xor U705 (N_705,In_938,N_468);
and U706 (N_706,In_1029,In_627);
xnor U707 (N_707,In_435,In_50);
or U708 (N_708,In_1170,In_446);
and U709 (N_709,N_549,N_550);
and U710 (N_710,In_714,In_928);
xnor U711 (N_711,N_242,In_741);
xor U712 (N_712,N_134,In_1024);
or U713 (N_713,N_591,In_135);
nor U714 (N_714,N_338,In_1298);
or U715 (N_715,N_356,In_93);
and U716 (N_716,N_451,In_683);
xor U717 (N_717,In_1149,In_1497);
or U718 (N_718,In_459,N_437);
and U719 (N_719,In_287,In_1116);
and U720 (N_720,In_151,N_432);
nand U721 (N_721,In_264,In_1128);
or U722 (N_722,In_1247,N_478);
nor U723 (N_723,N_364,In_1492);
nor U724 (N_724,In_442,In_130);
nor U725 (N_725,In_762,In_1332);
xor U726 (N_726,N_539,In_486);
xnor U727 (N_727,N_515,N_497);
and U728 (N_728,In_45,N_72);
or U729 (N_729,In_990,In_241);
nand U730 (N_730,N_284,In_1210);
and U731 (N_731,N_467,N_536);
or U732 (N_732,In_692,In_622);
and U733 (N_733,N_191,In_806);
and U734 (N_734,N_161,In_512);
nor U735 (N_735,In_1450,N_373);
or U736 (N_736,In_237,N_295);
nor U737 (N_737,N_453,In_752);
xnor U738 (N_738,In_757,N_556);
and U739 (N_739,N_254,N_513);
and U740 (N_740,N_296,N_614);
and U741 (N_741,N_219,In_1271);
and U742 (N_742,In_201,In_1122);
or U743 (N_743,In_1083,N_564);
nor U744 (N_744,In_30,In_610);
and U745 (N_745,In_531,N_293);
xnor U746 (N_746,N_541,N_397);
and U747 (N_747,In_768,In_99);
and U748 (N_748,In_1329,In_935);
xor U749 (N_749,In_606,In_1412);
and U750 (N_750,N_585,N_227);
nand U751 (N_751,N_694,N_737);
and U752 (N_752,N_43,In_995);
xor U753 (N_753,In_989,N_450);
nor U754 (N_754,In_943,N_39);
or U755 (N_755,N_672,N_409);
and U756 (N_756,In_51,In_371);
or U757 (N_757,N_542,N_660);
nand U758 (N_758,In_452,N_740);
and U759 (N_759,In_534,In_1490);
and U760 (N_760,N_736,In_1491);
nand U761 (N_761,In_1218,N_372);
or U762 (N_762,N_701,In_262);
and U763 (N_763,N_616,N_141);
and U764 (N_764,N_669,In_794);
and U765 (N_765,In_342,In_1031);
xnor U766 (N_766,In_850,In_1073);
and U767 (N_767,N_168,In_681);
xnor U768 (N_768,In_61,In_143);
nor U769 (N_769,N_404,In_252);
and U770 (N_770,In_527,In_366);
or U771 (N_771,In_251,N_166);
or U772 (N_772,N_213,In_298);
nor U773 (N_773,In_133,In_1397);
and U774 (N_774,N_712,N_250);
xor U775 (N_775,N_135,N_659);
or U776 (N_776,N_5,N_632);
or U777 (N_777,In_114,N_730);
nor U778 (N_778,In_560,N_327);
and U779 (N_779,In_550,In_1381);
nor U780 (N_780,N_745,In_137);
and U781 (N_781,N_714,N_45);
xnor U782 (N_782,N_392,In_341);
or U783 (N_783,N_383,In_564);
or U784 (N_784,In_1223,N_593);
and U785 (N_785,N_370,N_320);
or U786 (N_786,In_458,N_738);
xnor U787 (N_787,N_340,N_512);
nor U788 (N_788,In_1269,In_437);
nand U789 (N_789,N_429,In_540);
and U790 (N_790,N_454,In_423);
xor U791 (N_791,In_481,In_491);
xor U792 (N_792,N_377,N_518);
nor U793 (N_793,N_452,N_157);
xor U794 (N_794,N_492,N_748);
xnor U795 (N_795,In_330,In_489);
nor U796 (N_796,N_567,In_894);
or U797 (N_797,In_697,N_648);
and U798 (N_798,N_618,N_315);
xor U799 (N_799,N_711,N_384);
nand U800 (N_800,In_249,N_651);
nand U801 (N_801,N_621,In_177);
xor U802 (N_802,N_584,N_625);
or U803 (N_803,N_482,In_1018);
nor U804 (N_804,N_653,In_1111);
or U805 (N_805,N_517,N_569);
and U806 (N_806,In_778,N_609);
xor U807 (N_807,N_606,N_442);
xnor U808 (N_808,In_132,In_216);
or U809 (N_809,In_999,In_1440);
xnor U810 (N_810,In_1245,In_141);
nand U811 (N_811,N_476,N_508);
nand U812 (N_812,In_195,In_1164);
nand U813 (N_813,In_267,In_904);
or U814 (N_814,N_26,In_537);
nand U815 (N_815,In_67,In_913);
and U816 (N_816,N_20,N_277);
nand U817 (N_817,N_719,In_1446);
or U818 (N_818,In_1396,In_227);
nand U819 (N_819,In_63,N_346);
or U820 (N_820,N_31,In_467);
or U821 (N_821,N_87,In_1062);
nand U822 (N_822,In_424,N_529);
and U823 (N_823,In_1032,N_283);
nand U824 (N_824,N_378,N_678);
nor U825 (N_825,N_718,N_382);
or U826 (N_826,In_162,N_746);
nor U827 (N_827,N_193,In_1361);
or U828 (N_828,In_993,N_686);
xnor U829 (N_829,N_345,N_623);
or U830 (N_830,N_610,In_869);
and U831 (N_831,In_1370,In_1409);
nand U832 (N_832,N_388,In_1494);
nor U833 (N_833,In_682,N_272);
nand U834 (N_834,N_195,In_173);
nor U835 (N_835,N_305,N_36);
nor U836 (N_836,In_1200,N_73);
nor U837 (N_837,N_692,N_408);
and U838 (N_838,N_538,In_1196);
nor U839 (N_839,N_727,In_763);
or U840 (N_840,In_432,In_1439);
and U841 (N_841,N_138,N_390);
nand U842 (N_842,N_543,N_521);
nand U843 (N_843,In_1052,N_376);
and U844 (N_844,In_281,In_104);
nand U845 (N_845,In_813,In_221);
nand U846 (N_846,N_725,In_1366);
nand U847 (N_847,In_923,N_607);
xor U848 (N_848,In_884,N_721);
or U849 (N_849,In_1407,In_840);
xnor U850 (N_850,In_1255,In_994);
xnor U851 (N_851,In_1365,N_627);
nand U852 (N_852,In_176,N_420);
nand U853 (N_853,N_3,N_304);
nor U854 (N_854,N_732,N_405);
or U855 (N_855,N_663,In_781);
and U856 (N_856,N_582,N_638);
xnor U857 (N_857,In_1470,N_689);
nor U858 (N_858,In_979,In_178);
or U859 (N_859,N_362,N_645);
nand U860 (N_860,In_101,In_533);
nor U861 (N_861,N_729,N_499);
and U862 (N_862,N_562,N_395);
nor U863 (N_863,In_939,N_281);
nor U864 (N_864,N_658,In_1085);
and U865 (N_865,N_551,In_664);
nand U866 (N_866,N_500,In_576);
and U867 (N_867,N_485,N_274);
nand U868 (N_868,N_431,In_1476);
nor U869 (N_869,N_414,N_465);
and U870 (N_870,In_209,N_235);
xor U871 (N_871,N_6,N_516);
nand U872 (N_872,In_739,In_718);
or U873 (N_873,In_1474,In_1100);
or U874 (N_874,In_498,In_543);
nor U875 (N_875,In_233,In_1117);
or U876 (N_876,N_713,N_417);
nor U877 (N_877,In_168,In_1479);
xnor U878 (N_878,In_1457,N_707);
and U879 (N_879,N_654,In_1266);
and U880 (N_880,N_799,N_520);
xor U881 (N_881,In_685,N_757);
or U882 (N_882,In_1419,N_866);
nor U883 (N_883,In_89,N_581);
and U884 (N_884,N_630,N_836);
xor U885 (N_885,In_1044,In_820);
nor U886 (N_886,In_601,N_844);
xnor U887 (N_887,In_1079,N_837);
xnor U888 (N_888,N_41,N_360);
nor U889 (N_889,In_85,N_706);
nand U890 (N_890,N_187,N_419);
nand U891 (N_891,N_507,In_976);
nand U892 (N_892,In_317,In_853);
nand U893 (N_893,In_408,In_1363);
nor U894 (N_894,N_629,N_814);
or U895 (N_895,N_825,N_553);
nand U896 (N_896,N_773,N_795);
nor U897 (N_897,In_269,N_125);
nand U898 (N_898,In_53,N_834);
nand U899 (N_899,In_1499,N_808);
nand U900 (N_900,N_55,In_1441);
xor U901 (N_901,N_644,N_862);
and U902 (N_902,In_1057,N_733);
nand U903 (N_903,N_357,N_280);
or U904 (N_904,In_191,In_122);
or U905 (N_905,N_677,N_759);
and U906 (N_906,N_780,N_598);
nor U907 (N_907,N_667,In_611);
and U908 (N_908,N_771,N_637);
and U909 (N_909,In_826,In_1171);
nor U910 (N_910,In_1156,N_822);
nor U911 (N_911,In_513,N_696);
nand U912 (N_912,N_752,In_557);
nand U913 (N_913,N_690,In_968);
or U914 (N_914,N_800,In_65);
and U915 (N_915,N_206,N_776);
or U916 (N_916,N_703,N_531);
nand U917 (N_917,N_704,In_1465);
xor U918 (N_918,N_691,N_246);
xnor U919 (N_919,In_1340,N_849);
or U920 (N_920,N_642,In_128);
nand U921 (N_921,N_183,N_446);
or U922 (N_922,N_662,N_494);
and U923 (N_923,In_1212,N_511);
nor U924 (N_924,N_466,N_297);
nor U925 (N_925,In_1019,N_265);
xor U926 (N_926,In_83,N_774);
or U927 (N_927,In_329,N_312);
nor U928 (N_928,In_1,N_491);
nand U929 (N_929,N_811,In_154);
nor U930 (N_930,In_1030,N_699);
nand U931 (N_931,N_765,N_596);
or U932 (N_932,N_259,In_724);
or U933 (N_933,N_433,In_369);
nand U934 (N_934,N_639,N_12);
and U935 (N_935,In_650,N_674);
and U936 (N_936,N_688,In_961);
nand U937 (N_937,N_680,N_850);
nor U938 (N_938,In_1207,N_116);
nand U939 (N_939,N_459,N_734);
nand U940 (N_940,In_977,N_715);
nand U941 (N_941,N_460,N_592);
xor U942 (N_942,In_861,N_749);
or U943 (N_943,N_506,In_1410);
or U944 (N_944,In_635,In_1466);
nand U945 (N_945,In_379,N_846);
or U946 (N_946,N_8,In_942);
nand U947 (N_947,In_419,N_51);
xor U948 (N_948,N_394,N_548);
or U949 (N_949,In_1308,N_873);
xnor U950 (N_950,N_99,N_693);
nand U951 (N_951,In_625,N_600);
or U952 (N_952,N_421,In_213);
xor U953 (N_953,N_308,N_181);
xnor U954 (N_954,N_842,N_835);
and U955 (N_955,N_840,In_643);
xor U956 (N_956,In_1272,N_698);
and U957 (N_957,N_731,In_355);
nor U958 (N_958,N_768,N_619);
nor U959 (N_959,N_535,In_1148);
or U960 (N_960,In_271,N_743);
xnor U961 (N_961,N_252,N_769);
or U962 (N_962,N_683,In_454);
or U963 (N_963,In_415,N_807);
nand U964 (N_964,N_652,In_410);
and U965 (N_965,In_1080,N_565);
nand U966 (N_966,N_647,N_818);
nand U967 (N_967,In_1206,In_1306);
nor U968 (N_968,N_270,In_1005);
nand U969 (N_969,In_384,In_1077);
nand U970 (N_970,N_402,N_624);
or U971 (N_971,In_753,In_1387);
or U972 (N_972,N_209,N_857);
and U973 (N_973,N_313,In_670);
or U974 (N_974,N_741,In_71);
nor U975 (N_975,In_340,N_32);
or U976 (N_976,N_824,In_957);
or U977 (N_977,N_578,N_447);
xor U978 (N_978,In_157,In_336);
nor U979 (N_979,N_636,N_782);
xor U980 (N_980,N_628,In_111);
xor U981 (N_981,N_47,In_13);
nor U982 (N_982,N_586,N_286);
and U983 (N_983,N_590,In_1273);
or U984 (N_984,In_19,N_829);
and U985 (N_985,In_908,N_597);
xor U986 (N_986,In_914,In_244);
nor U987 (N_987,N_783,In_200);
xnor U988 (N_988,In_671,N_342);
nor U989 (N_989,In_1478,N_258);
xor U990 (N_990,N_826,N_412);
and U991 (N_991,N_577,N_303);
and U992 (N_992,N_522,N_231);
or U993 (N_993,N_823,N_92);
or U994 (N_994,In_731,In_488);
or U995 (N_995,N_751,N_640);
and U996 (N_996,N_568,N_440);
nand U997 (N_997,N_472,N_747);
and U998 (N_998,N_587,N_685);
xnor U999 (N_999,N_262,N_775);
and U1000 (N_1000,N_533,N_991);
nor U1001 (N_1001,N_993,N_207);
xnor U1002 (N_1002,N_853,N_861);
nor U1003 (N_1003,N_455,N_909);
and U1004 (N_1004,N_365,In_1155);
nand U1005 (N_1005,N_415,In_1467);
or U1006 (N_1006,N_495,In_760);
or U1007 (N_1007,N_670,N_887);
nand U1008 (N_1008,N_744,N_552);
and U1009 (N_1009,In_1009,N_918);
nor U1010 (N_1010,N_898,N_930);
and U1011 (N_1011,In_774,In_758);
xor U1012 (N_1012,In_933,N_787);
nand U1013 (N_1013,N_199,N_631);
nand U1014 (N_1014,N_665,N_257);
and U1015 (N_1015,N_926,N_756);
and U1016 (N_1016,In_300,N_537);
and U1017 (N_1017,In_74,N_546);
or U1018 (N_1018,N_720,N_868);
nor U1019 (N_1019,N_595,N_188);
or U1020 (N_1020,N_399,N_962);
xnor U1021 (N_1021,N_510,N_943);
and U1022 (N_1022,In_1285,N_247);
and U1023 (N_1023,N_976,N_946);
nor U1024 (N_1024,N_819,N_988);
or U1025 (N_1025,N_505,N_649);
nor U1026 (N_1026,N_477,N_934);
nor U1027 (N_1027,In_483,N_753);
and U1028 (N_1028,N_655,N_874);
xor U1029 (N_1029,N_750,N_978);
or U1030 (N_1030,N_796,N_858);
nand U1031 (N_1031,N_786,N_855);
and U1032 (N_1032,In_526,N_802);
nand U1033 (N_1033,In_618,In_1317);
nand U1034 (N_1034,In_732,In_1104);
or U1035 (N_1035,N_889,N_778);
or U1036 (N_1036,N_758,In_940);
and U1037 (N_1037,In_981,N_475);
or U1038 (N_1038,N_970,N_761);
or U1039 (N_1039,N_901,N_661);
xnor U1040 (N_1040,In_1103,N_959);
nor U1041 (N_1041,In_490,N_504);
xor U1042 (N_1042,In_518,N_990);
or U1043 (N_1043,In_485,In_146);
and U1044 (N_1044,N_950,In_892);
and U1045 (N_1045,N_657,In_1334);
nor U1046 (N_1046,N_931,N_947);
and U1047 (N_1047,N_865,N_815);
xor U1048 (N_1048,N_579,N_673);
xnor U1049 (N_1049,N_119,N_902);
or U1050 (N_1050,N_643,N_992);
nor U1051 (N_1051,N_935,N_351);
xnor U1052 (N_1052,N_679,In_587);
nand U1053 (N_1053,In_1283,N_928);
and U1054 (N_1054,In_1121,N_717);
nor U1055 (N_1055,N_998,In_986);
xor U1056 (N_1056,N_890,N_705);
or U1057 (N_1057,N_764,In_815);
xor U1058 (N_1058,N_545,In_843);
or U1059 (N_1059,N_726,N_306);
and U1060 (N_1060,N_886,In_364);
nor U1061 (N_1061,N_888,N_779);
xor U1062 (N_1062,N_120,N_876);
nor U1063 (N_1063,N_894,N_885);
nand U1064 (N_1064,N_867,N_288);
nand U1065 (N_1065,N_728,N_863);
and U1066 (N_1066,N_332,N_563);
nor U1067 (N_1067,N_666,N_851);
nand U1068 (N_1068,N_833,N_566);
and U1069 (N_1069,N_893,N_435);
nand U1070 (N_1070,N_957,In_886);
and U1071 (N_1071,N_575,In_1453);
and U1072 (N_1072,N_989,N_695);
nor U1073 (N_1073,N_856,In_642);
or U1074 (N_1074,In_1482,N_832);
or U1075 (N_1075,N_410,In_3);
or U1076 (N_1076,In_1498,N_634);
nor U1077 (N_1077,In_541,N_791);
or U1078 (N_1078,In_1022,N_880);
xnor U1079 (N_1079,N_958,In_1021);
nor U1080 (N_1080,N_937,In_708);
nor U1081 (N_1081,In_1277,N_82);
or U1082 (N_1082,N_971,In_1089);
xnor U1083 (N_1083,N_884,In_1371);
xnor U1084 (N_1084,N_766,N_682);
or U1085 (N_1085,In_631,In_403);
xnor U1086 (N_1086,In_407,N_792);
nand U1087 (N_1087,In_956,In_548);
or U1088 (N_1088,N_805,In_339);
and U1089 (N_1089,In_1429,N_892);
nor U1090 (N_1090,In_456,N_684);
nor U1091 (N_1091,N_929,N_961);
xor U1092 (N_1092,N_502,N_975);
nand U1093 (N_1093,N_675,In_349);
nor U1094 (N_1094,N_980,N_532);
xnor U1095 (N_1095,N_700,N_223);
xor U1096 (N_1096,N_724,N_999);
xnor U1097 (N_1097,N_797,N_755);
xor U1098 (N_1098,N_881,In_212);
xor U1099 (N_1099,N_831,In_189);
and U1100 (N_1100,N_891,N_810);
or U1101 (N_1101,N_434,N_813);
and U1102 (N_1102,N_710,In_91);
nand U1103 (N_1103,N_983,N_249);
nor U1104 (N_1104,N_49,N_969);
xnor U1105 (N_1105,In_1296,N_671);
xor U1106 (N_1106,In_1238,In_792);
nor U1107 (N_1107,N_925,N_650);
nor U1108 (N_1108,N_948,N_972);
nor U1109 (N_1109,N_827,N_854);
nor U1110 (N_1110,N_924,N_953);
xnor U1111 (N_1111,N_464,N_951);
or U1112 (N_1112,N_438,N_359);
and U1113 (N_1113,N_557,N_613);
nand U1114 (N_1114,In_523,N_911);
nand U1115 (N_1115,N_604,N_914);
nand U1116 (N_1116,N_900,N_830);
nand U1117 (N_1117,N_952,N_967);
and U1118 (N_1118,N_770,N_430);
xor U1119 (N_1119,N_664,In_1346);
xnor U1120 (N_1120,N_514,N_443);
nor U1121 (N_1121,In_926,N_668);
xor U1122 (N_1122,N_540,N_869);
nand U1123 (N_1123,N_985,N_781);
or U1124 (N_1124,In_817,N_54);
nor U1125 (N_1125,N_933,N_940);
and U1126 (N_1126,N_620,N_594);
nand U1127 (N_1127,N_676,N_809);
nand U1128 (N_1128,N_1075,N_1095);
and U1129 (N_1129,N_954,N_960);
xor U1130 (N_1130,N_907,N_687);
nand U1131 (N_1131,N_544,N_1070);
and U1132 (N_1132,N_803,N_955);
and U1133 (N_1133,N_742,In_1230);
xnor U1134 (N_1134,N_1110,N_1056);
xnor U1135 (N_1135,N_488,N_1046);
or U1136 (N_1136,In_1208,N_656);
nor U1137 (N_1137,N_127,N_1005);
or U1138 (N_1138,N_702,N_938);
xor U1139 (N_1139,N_371,N_1086);
nand U1140 (N_1140,N_968,N_927);
nor U1141 (N_1141,N_878,N_1124);
and U1142 (N_1142,N_1097,N_1120);
nor U1143 (N_1143,N_899,N_966);
nor U1144 (N_1144,In_1102,In_243);
nor U1145 (N_1145,N_1040,N_1061);
and U1146 (N_1146,In_12,N_1034);
and U1147 (N_1147,N_275,N_915);
nor U1148 (N_1148,N_681,N_1094);
nor U1149 (N_1149,N_1084,N_784);
xnor U1150 (N_1150,N_201,N_1001);
nand U1151 (N_1151,N_790,N_860);
nor U1152 (N_1152,In_250,N_1004);
and U1153 (N_1153,In_721,In_619);
nor U1154 (N_1154,In_1026,N_1028);
xor U1155 (N_1155,N_870,In_196);
and U1156 (N_1156,N_1080,N_1027);
nand U1157 (N_1157,N_1102,N_1098);
and U1158 (N_1158,N_944,In_729);
nor U1159 (N_1159,N_794,N_461);
nor U1160 (N_1160,N_558,N_474);
xnor U1161 (N_1161,N_218,N_1099);
nand U1162 (N_1162,In_455,N_919);
xor U1163 (N_1163,N_380,In_1348);
xnor U1164 (N_1164,N_903,N_1113);
nor U1165 (N_1165,N_646,N_963);
nand U1166 (N_1166,N_839,In_1105);
or U1167 (N_1167,N_1054,N_1109);
nor U1168 (N_1168,N_1042,N_895);
xnor U1169 (N_1169,In_838,N_793);
nor U1170 (N_1170,N_94,N_1030);
nand U1171 (N_1171,N_635,N_1052);
nand U1172 (N_1172,N_1033,N_480);
xnor U1173 (N_1173,N_317,In_929);
nor U1174 (N_1174,In_1177,In_924);
and U1175 (N_1175,In_1145,N_941);
nand U1176 (N_1176,In_1432,N_1025);
and U1177 (N_1177,N_1081,N_939);
nand U1178 (N_1178,N_716,N_503);
nand U1179 (N_1179,N_1049,In_1154);
xor U1180 (N_1180,N_828,N_1087);
nand U1181 (N_1181,N_1050,N_820);
or U1182 (N_1182,N_789,N_353);
nor U1183 (N_1183,N_605,N_982);
nand U1184 (N_1184,N_1059,N_307);
or U1185 (N_1185,N_128,N_859);
xor U1186 (N_1186,N_1020,N_821);
or U1187 (N_1187,N_1003,N_1011);
nor U1188 (N_1188,N_936,N_910);
nor U1189 (N_1189,N_1106,N_735);
and U1190 (N_1190,In_996,N_996);
or U1191 (N_1191,N_576,N_772);
or U1192 (N_1192,In_9,In_1082);
nor U1193 (N_1193,N_1112,N_1038);
nor U1194 (N_1194,N_1088,N_184);
nand U1195 (N_1195,N_1103,N_801);
nor U1196 (N_1196,N_1035,N_1101);
nand U1197 (N_1197,In_331,N_1114);
nand U1198 (N_1198,N_1073,N_1058);
xnor U1199 (N_1199,N_977,In_318);
nand U1200 (N_1200,N_1064,N_882);
nor U1201 (N_1201,N_626,N_1022);
and U1202 (N_1202,In_1393,In_373);
nand U1203 (N_1203,N_1077,N_956);
and U1204 (N_1204,N_908,N_1036);
and U1205 (N_1205,N_1066,N_641);
xnor U1206 (N_1206,N_1093,N_838);
or U1207 (N_1207,In_118,N_965);
nand U1208 (N_1208,N_1091,N_484);
or U1209 (N_1209,N_762,N_872);
nand U1210 (N_1210,N_603,N_922);
nor U1211 (N_1211,N_816,N_1115);
or U1212 (N_1212,N_1051,N_1039);
and U1213 (N_1213,N_984,N_444);
and U1214 (N_1214,N_932,N_697);
xor U1215 (N_1215,N_981,N_1010);
nand U1216 (N_1216,N_172,In_788);
nor U1217 (N_1217,In_1382,N_1069);
and U1218 (N_1218,N_1065,N_1014);
and U1219 (N_1219,N_722,N_1000);
and U1220 (N_1220,N_843,N_997);
or U1221 (N_1221,N_949,N_1006);
nand U1222 (N_1222,N_917,N_186);
or U1223 (N_1223,N_877,N_817);
and U1224 (N_1224,N_1089,N_159);
and U1225 (N_1225,N_185,N_1053);
nor U1226 (N_1226,N_852,N_1024);
and U1227 (N_1227,In_925,N_973);
nand U1228 (N_1228,N_760,N_335);
xnor U1229 (N_1229,N_554,N_1100);
or U1230 (N_1230,N_812,N_35);
xnor U1231 (N_1231,N_416,N_238);
nor U1232 (N_1232,N_1032,N_1021);
nor U1233 (N_1233,N_767,N_905);
nand U1234 (N_1234,N_487,N_1067);
or U1235 (N_1235,N_1116,N_883);
xor U1236 (N_1236,N_441,N_381);
nand U1237 (N_1237,N_121,N_198);
nand U1238 (N_1238,N_229,In_1342);
and U1239 (N_1239,N_986,N_1122);
nor U1240 (N_1240,N_1092,In_290);
or U1241 (N_1241,N_913,N_1012);
or U1242 (N_1242,N_777,N_343);
or U1243 (N_1243,N_1085,N_617);
nor U1244 (N_1244,N_979,N_14);
or U1245 (N_1245,In_1316,N_875);
or U1246 (N_1246,In_975,N_389);
or U1247 (N_1247,N_298,N_1008);
and U1248 (N_1248,N_1105,N_144);
or U1249 (N_1249,N_921,N_1083);
and U1250 (N_1250,N_1104,In_1096);
nand U1251 (N_1251,N_1233,N_1180);
nand U1252 (N_1252,N_1218,N_1221);
and U1253 (N_1253,N_1207,N_1170);
and U1254 (N_1254,N_1107,N_754);
and U1255 (N_1255,N_1155,N_1140);
nor U1256 (N_1256,In_668,In_1242);
and U1257 (N_1257,N_1208,N_1019);
xnor U1258 (N_1258,N_1212,N_788);
nor U1259 (N_1259,N_806,N_1241);
and U1260 (N_1260,N_1135,N_1238);
and U1261 (N_1261,N_1063,N_1136);
nand U1262 (N_1262,N_871,N_1211);
or U1263 (N_1263,In_602,In_823);
xor U1264 (N_1264,N_1223,N_1045);
and U1265 (N_1265,In_950,N_798);
nand U1266 (N_1266,N_1074,N_1214);
nand U1267 (N_1267,N_1230,N_974);
and U1268 (N_1268,N_615,N_964);
nand U1269 (N_1269,N_1247,N_1164);
nand U1270 (N_1270,N_879,N_25);
nor U1271 (N_1271,N_1119,N_864);
xor U1272 (N_1272,N_1125,N_1057);
and U1273 (N_1273,N_995,N_400);
nor U1274 (N_1274,N_1123,N_1172);
or U1275 (N_1275,N_1197,N_1231);
nor U1276 (N_1276,N_1137,N_1007);
and U1277 (N_1277,N_1026,N_1127);
xor U1278 (N_1278,N_611,N_1204);
and U1279 (N_1279,N_60,N_526);
or U1280 (N_1280,N_1243,N_1194);
or U1281 (N_1281,In_1472,N_1210);
xnor U1282 (N_1282,N_1206,N_945);
and U1283 (N_1283,In_179,N_1018);
xnor U1284 (N_1284,N_1111,N_496);
or U1285 (N_1285,N_1245,N_1129);
and U1286 (N_1286,N_1190,In_1395);
nor U1287 (N_1287,N_1126,N_1239);
xnor U1288 (N_1288,N_1068,N_1242);
nor U1289 (N_1289,N_1141,N_1217);
or U1290 (N_1290,N_1209,In_893);
nor U1291 (N_1291,N_1178,N_633);
or U1292 (N_1292,N_1156,In_460);
and U1293 (N_1293,N_1072,N_1048);
and U1294 (N_1294,N_1183,In_1098);
xor U1295 (N_1295,In_628,N_1139);
or U1296 (N_1296,In_804,N_1235);
or U1297 (N_1297,N_1133,N_1143);
xnor U1298 (N_1298,N_1216,N_1225);
xor U1299 (N_1299,N_1016,N_1191);
and U1300 (N_1300,N_739,N_1144);
xor U1301 (N_1301,N_1043,N_393);
xor U1302 (N_1302,N_1076,N_1062);
nand U1303 (N_1303,N_1228,In_1434);
xnor U1304 (N_1304,N_1031,N_912);
or U1305 (N_1305,N_1166,N_1108);
nand U1306 (N_1306,N_1060,N_1236);
or U1307 (N_1307,N_1157,N_1229);
nand U1308 (N_1308,N_845,N_1174);
or U1309 (N_1309,In_1175,N_847);
nand U1310 (N_1310,N_1185,N_1186);
and U1311 (N_1311,N_994,N_1219);
nor U1312 (N_1312,N_1082,N_1181);
xnor U1313 (N_1313,N_1079,N_1163);
xor U1314 (N_1314,N_1118,N_1078);
xor U1315 (N_1315,N_723,N_1169);
nor U1316 (N_1316,N_1249,N_1132);
xnor U1317 (N_1317,N_1182,N_1131);
nor U1318 (N_1318,N_1179,N_763);
xor U1319 (N_1319,N_69,N_1017);
xnor U1320 (N_1320,N_1117,N_785);
or U1321 (N_1321,N_1162,N_1215);
and U1322 (N_1322,N_942,N_1226);
and U1323 (N_1323,N_530,N_708);
or U1324 (N_1324,N_1147,N_848);
and U1325 (N_1325,N_1193,N_1189);
xnor U1326 (N_1326,N_1158,N_1037);
xnor U1327 (N_1327,N_1096,N_425);
xor U1328 (N_1328,N_904,N_1196);
xnor U1329 (N_1329,N_1151,N_1002);
xnor U1330 (N_1330,N_422,N_1173);
and U1331 (N_1331,N_1159,N_361);
and U1332 (N_1332,N_1198,N_1234);
nand U1333 (N_1333,N_1227,In_258);
xnor U1334 (N_1334,N_1152,N_1188);
and U1335 (N_1335,N_1013,N_1090);
xor U1336 (N_1336,N_559,N_1130);
xnor U1337 (N_1337,N_1071,N_709);
nand U1338 (N_1338,N_1047,N_1154);
nor U1339 (N_1339,N_1176,N_1232);
nor U1340 (N_1340,N_1168,N_1167);
and U1341 (N_1341,N_906,N_325);
and U1342 (N_1342,N_1248,N_1202);
nor U1343 (N_1343,N_1177,N_1150);
nand U1344 (N_1344,N_1142,N_1200);
nor U1345 (N_1345,N_1192,N_1121);
or U1346 (N_1346,N_1029,N_1184);
or U1347 (N_1347,N_916,N_321);
nand U1348 (N_1348,In_1413,N_1044);
or U1349 (N_1349,N_1224,N_1161);
nand U1350 (N_1350,N_555,N_1148);
nand U1351 (N_1351,N_89,N_1195);
nor U1352 (N_1352,In_1417,N_1237);
and U1353 (N_1353,N_1222,N_221);
and U1354 (N_1354,N_896,N_1149);
and U1355 (N_1355,N_1246,N_1160);
or U1356 (N_1356,N_583,N_1041);
nor U1357 (N_1357,N_1201,N_1220);
and U1358 (N_1358,N_987,In_1377);
nand U1359 (N_1359,N_1153,N_374);
xnor U1360 (N_1360,N_1009,N_1128);
xnor U1361 (N_1361,N_1134,N_1023);
xnor U1362 (N_1362,N_1171,N_923);
xor U1363 (N_1363,N_1015,In_831);
or U1364 (N_1364,N_1203,N_489);
xnor U1365 (N_1365,N_1240,N_1213);
or U1366 (N_1366,N_1145,N_1146);
nand U1367 (N_1367,N_1138,N_1187);
or U1368 (N_1368,N_1175,In_411);
nor U1369 (N_1369,N_1199,N_1244);
or U1370 (N_1370,In_1007,In_288);
or U1371 (N_1371,N_1205,N_920);
or U1372 (N_1372,N_897,N_1055);
and U1373 (N_1373,N_1165,N_841);
or U1374 (N_1374,N_612,N_804);
xnor U1375 (N_1375,N_1261,N_1287);
or U1376 (N_1376,N_1276,N_1330);
xnor U1377 (N_1377,N_1273,N_1313);
or U1378 (N_1378,N_1304,N_1339);
nand U1379 (N_1379,N_1301,N_1346);
xnor U1380 (N_1380,N_1252,N_1325);
and U1381 (N_1381,N_1316,N_1250);
nand U1382 (N_1382,N_1333,N_1259);
and U1383 (N_1383,N_1292,N_1344);
and U1384 (N_1384,N_1326,N_1274);
nor U1385 (N_1385,N_1372,N_1373);
nor U1386 (N_1386,N_1270,N_1295);
nand U1387 (N_1387,N_1343,N_1319);
xnor U1388 (N_1388,N_1257,N_1298);
nand U1389 (N_1389,N_1263,N_1309);
and U1390 (N_1390,N_1268,N_1291);
nand U1391 (N_1391,N_1306,N_1369);
nor U1392 (N_1392,N_1310,N_1266);
xor U1393 (N_1393,N_1328,N_1277);
and U1394 (N_1394,N_1305,N_1285);
nor U1395 (N_1395,N_1324,N_1253);
xnor U1396 (N_1396,N_1359,N_1258);
xnor U1397 (N_1397,N_1307,N_1327);
xnor U1398 (N_1398,N_1323,N_1363);
and U1399 (N_1399,N_1275,N_1288);
nor U1400 (N_1400,N_1368,N_1351);
nor U1401 (N_1401,N_1251,N_1367);
nand U1402 (N_1402,N_1300,N_1338);
nor U1403 (N_1403,N_1284,N_1321);
nand U1404 (N_1404,N_1332,N_1357);
or U1405 (N_1405,N_1254,N_1322);
or U1406 (N_1406,N_1272,N_1342);
or U1407 (N_1407,N_1299,N_1336);
and U1408 (N_1408,N_1364,N_1267);
nand U1409 (N_1409,N_1294,N_1317);
nand U1410 (N_1410,N_1280,N_1335);
or U1411 (N_1411,N_1350,N_1348);
and U1412 (N_1412,N_1308,N_1278);
or U1413 (N_1413,N_1353,N_1293);
and U1414 (N_1414,N_1269,N_1365);
or U1415 (N_1415,N_1352,N_1289);
nor U1416 (N_1416,N_1334,N_1370);
nor U1417 (N_1417,N_1374,N_1360);
nand U1418 (N_1418,N_1312,N_1290);
nand U1419 (N_1419,N_1256,N_1341);
xnor U1420 (N_1420,N_1362,N_1311);
or U1421 (N_1421,N_1303,N_1265);
nor U1422 (N_1422,N_1356,N_1371);
and U1423 (N_1423,N_1320,N_1318);
or U1424 (N_1424,N_1279,N_1314);
and U1425 (N_1425,N_1337,N_1286);
or U1426 (N_1426,N_1329,N_1282);
or U1427 (N_1427,N_1347,N_1260);
and U1428 (N_1428,N_1315,N_1345);
xnor U1429 (N_1429,N_1358,N_1297);
xor U1430 (N_1430,N_1283,N_1281);
xor U1431 (N_1431,N_1302,N_1271);
and U1432 (N_1432,N_1296,N_1354);
xor U1433 (N_1433,N_1262,N_1331);
nand U1434 (N_1434,N_1355,N_1366);
or U1435 (N_1435,N_1361,N_1255);
xnor U1436 (N_1436,N_1340,N_1349);
nor U1437 (N_1437,N_1264,N_1253);
nor U1438 (N_1438,N_1367,N_1263);
nor U1439 (N_1439,N_1347,N_1358);
xnor U1440 (N_1440,N_1324,N_1351);
xor U1441 (N_1441,N_1332,N_1271);
xor U1442 (N_1442,N_1356,N_1277);
and U1443 (N_1443,N_1339,N_1266);
nor U1444 (N_1444,N_1275,N_1348);
xnor U1445 (N_1445,N_1311,N_1353);
nor U1446 (N_1446,N_1354,N_1251);
xnor U1447 (N_1447,N_1350,N_1269);
nor U1448 (N_1448,N_1306,N_1290);
or U1449 (N_1449,N_1263,N_1274);
nand U1450 (N_1450,N_1302,N_1282);
nand U1451 (N_1451,N_1308,N_1327);
or U1452 (N_1452,N_1292,N_1316);
nor U1453 (N_1453,N_1324,N_1295);
nor U1454 (N_1454,N_1284,N_1369);
or U1455 (N_1455,N_1267,N_1332);
xor U1456 (N_1456,N_1370,N_1314);
and U1457 (N_1457,N_1338,N_1311);
or U1458 (N_1458,N_1274,N_1351);
and U1459 (N_1459,N_1252,N_1301);
or U1460 (N_1460,N_1360,N_1258);
nand U1461 (N_1461,N_1274,N_1374);
and U1462 (N_1462,N_1276,N_1264);
nor U1463 (N_1463,N_1308,N_1280);
or U1464 (N_1464,N_1351,N_1279);
nand U1465 (N_1465,N_1360,N_1313);
and U1466 (N_1466,N_1306,N_1307);
or U1467 (N_1467,N_1263,N_1295);
or U1468 (N_1468,N_1321,N_1261);
or U1469 (N_1469,N_1271,N_1293);
nor U1470 (N_1470,N_1305,N_1294);
nand U1471 (N_1471,N_1280,N_1329);
or U1472 (N_1472,N_1334,N_1263);
nand U1473 (N_1473,N_1341,N_1332);
nand U1474 (N_1474,N_1347,N_1346);
xor U1475 (N_1475,N_1306,N_1309);
and U1476 (N_1476,N_1351,N_1260);
nor U1477 (N_1477,N_1363,N_1297);
xnor U1478 (N_1478,N_1359,N_1291);
or U1479 (N_1479,N_1300,N_1280);
nand U1480 (N_1480,N_1328,N_1343);
nand U1481 (N_1481,N_1344,N_1286);
xor U1482 (N_1482,N_1320,N_1252);
or U1483 (N_1483,N_1289,N_1360);
and U1484 (N_1484,N_1321,N_1317);
nand U1485 (N_1485,N_1374,N_1288);
xor U1486 (N_1486,N_1348,N_1335);
nand U1487 (N_1487,N_1360,N_1311);
and U1488 (N_1488,N_1350,N_1354);
nor U1489 (N_1489,N_1251,N_1319);
and U1490 (N_1490,N_1257,N_1369);
and U1491 (N_1491,N_1334,N_1362);
nor U1492 (N_1492,N_1272,N_1274);
nand U1493 (N_1493,N_1274,N_1359);
and U1494 (N_1494,N_1348,N_1314);
and U1495 (N_1495,N_1323,N_1340);
xnor U1496 (N_1496,N_1371,N_1298);
nor U1497 (N_1497,N_1287,N_1303);
and U1498 (N_1498,N_1337,N_1298);
or U1499 (N_1499,N_1353,N_1341);
xnor U1500 (N_1500,N_1486,N_1377);
or U1501 (N_1501,N_1451,N_1424);
nor U1502 (N_1502,N_1493,N_1423);
xnor U1503 (N_1503,N_1452,N_1430);
nand U1504 (N_1504,N_1411,N_1417);
or U1505 (N_1505,N_1383,N_1425);
nand U1506 (N_1506,N_1459,N_1497);
nand U1507 (N_1507,N_1395,N_1433);
or U1508 (N_1508,N_1426,N_1472);
nor U1509 (N_1509,N_1385,N_1470);
nor U1510 (N_1510,N_1456,N_1449);
and U1511 (N_1511,N_1439,N_1415);
xor U1512 (N_1512,N_1488,N_1445);
and U1513 (N_1513,N_1474,N_1460);
xor U1514 (N_1514,N_1406,N_1429);
xor U1515 (N_1515,N_1495,N_1455);
nor U1516 (N_1516,N_1391,N_1480);
nand U1517 (N_1517,N_1487,N_1458);
and U1518 (N_1518,N_1421,N_1483);
xnor U1519 (N_1519,N_1443,N_1477);
or U1520 (N_1520,N_1498,N_1489);
nand U1521 (N_1521,N_1478,N_1410);
and U1522 (N_1522,N_1427,N_1462);
or U1523 (N_1523,N_1393,N_1407);
nand U1524 (N_1524,N_1467,N_1440);
nor U1525 (N_1525,N_1476,N_1446);
nand U1526 (N_1526,N_1418,N_1485);
xnor U1527 (N_1527,N_1380,N_1414);
or U1528 (N_1528,N_1399,N_1475);
xor U1529 (N_1529,N_1379,N_1419);
and U1530 (N_1530,N_1413,N_1389);
nor U1531 (N_1531,N_1457,N_1382);
nor U1532 (N_1532,N_1481,N_1402);
nor U1533 (N_1533,N_1494,N_1499);
or U1534 (N_1534,N_1465,N_1400);
nand U1535 (N_1535,N_1422,N_1386);
nand U1536 (N_1536,N_1412,N_1420);
and U1537 (N_1537,N_1453,N_1431);
and U1538 (N_1538,N_1404,N_1384);
and U1539 (N_1539,N_1461,N_1491);
and U1540 (N_1540,N_1468,N_1438);
xor U1541 (N_1541,N_1463,N_1432);
and U1542 (N_1542,N_1409,N_1447);
nor U1543 (N_1543,N_1403,N_1387);
xor U1544 (N_1544,N_1482,N_1376);
nor U1545 (N_1545,N_1434,N_1496);
nor U1546 (N_1546,N_1466,N_1401);
xor U1547 (N_1547,N_1394,N_1381);
xor U1548 (N_1548,N_1398,N_1388);
xor U1549 (N_1549,N_1469,N_1416);
xor U1550 (N_1550,N_1454,N_1442);
nand U1551 (N_1551,N_1428,N_1484);
xor U1552 (N_1552,N_1492,N_1479);
nor U1553 (N_1553,N_1490,N_1464);
nor U1554 (N_1554,N_1441,N_1397);
and U1555 (N_1555,N_1448,N_1471);
or U1556 (N_1556,N_1396,N_1390);
and U1557 (N_1557,N_1436,N_1375);
and U1558 (N_1558,N_1437,N_1392);
nor U1559 (N_1559,N_1444,N_1435);
nand U1560 (N_1560,N_1450,N_1378);
xor U1561 (N_1561,N_1473,N_1408);
nand U1562 (N_1562,N_1405,N_1468);
nand U1563 (N_1563,N_1453,N_1468);
nand U1564 (N_1564,N_1431,N_1461);
and U1565 (N_1565,N_1389,N_1456);
xnor U1566 (N_1566,N_1453,N_1418);
nor U1567 (N_1567,N_1452,N_1400);
nand U1568 (N_1568,N_1478,N_1466);
xnor U1569 (N_1569,N_1492,N_1446);
xor U1570 (N_1570,N_1440,N_1407);
nor U1571 (N_1571,N_1402,N_1376);
nand U1572 (N_1572,N_1462,N_1435);
xnor U1573 (N_1573,N_1396,N_1394);
xnor U1574 (N_1574,N_1445,N_1487);
and U1575 (N_1575,N_1497,N_1378);
nand U1576 (N_1576,N_1395,N_1410);
or U1577 (N_1577,N_1386,N_1464);
nor U1578 (N_1578,N_1403,N_1454);
or U1579 (N_1579,N_1477,N_1417);
nand U1580 (N_1580,N_1423,N_1381);
xor U1581 (N_1581,N_1458,N_1400);
and U1582 (N_1582,N_1473,N_1464);
nor U1583 (N_1583,N_1414,N_1381);
and U1584 (N_1584,N_1406,N_1446);
nand U1585 (N_1585,N_1436,N_1465);
and U1586 (N_1586,N_1412,N_1398);
or U1587 (N_1587,N_1445,N_1377);
xnor U1588 (N_1588,N_1449,N_1446);
nand U1589 (N_1589,N_1428,N_1432);
nand U1590 (N_1590,N_1381,N_1428);
xor U1591 (N_1591,N_1435,N_1449);
and U1592 (N_1592,N_1471,N_1398);
or U1593 (N_1593,N_1412,N_1383);
or U1594 (N_1594,N_1459,N_1479);
xnor U1595 (N_1595,N_1475,N_1398);
or U1596 (N_1596,N_1438,N_1494);
nand U1597 (N_1597,N_1455,N_1496);
xnor U1598 (N_1598,N_1419,N_1397);
and U1599 (N_1599,N_1450,N_1423);
nand U1600 (N_1600,N_1389,N_1383);
nand U1601 (N_1601,N_1399,N_1428);
nor U1602 (N_1602,N_1469,N_1459);
xor U1603 (N_1603,N_1403,N_1462);
xor U1604 (N_1604,N_1375,N_1396);
nor U1605 (N_1605,N_1499,N_1391);
xor U1606 (N_1606,N_1421,N_1495);
nand U1607 (N_1607,N_1480,N_1419);
or U1608 (N_1608,N_1493,N_1376);
xnor U1609 (N_1609,N_1473,N_1453);
or U1610 (N_1610,N_1461,N_1417);
nand U1611 (N_1611,N_1400,N_1412);
nand U1612 (N_1612,N_1422,N_1444);
or U1613 (N_1613,N_1484,N_1402);
or U1614 (N_1614,N_1462,N_1458);
xnor U1615 (N_1615,N_1483,N_1462);
and U1616 (N_1616,N_1486,N_1437);
or U1617 (N_1617,N_1495,N_1427);
nand U1618 (N_1618,N_1492,N_1497);
and U1619 (N_1619,N_1417,N_1390);
nand U1620 (N_1620,N_1430,N_1396);
or U1621 (N_1621,N_1452,N_1434);
nand U1622 (N_1622,N_1390,N_1399);
or U1623 (N_1623,N_1391,N_1393);
nand U1624 (N_1624,N_1482,N_1461);
xnor U1625 (N_1625,N_1620,N_1554);
or U1626 (N_1626,N_1619,N_1596);
nand U1627 (N_1627,N_1611,N_1539);
xor U1628 (N_1628,N_1517,N_1532);
nor U1629 (N_1629,N_1592,N_1606);
and U1630 (N_1630,N_1541,N_1526);
or U1631 (N_1631,N_1597,N_1577);
nand U1632 (N_1632,N_1614,N_1612);
and U1633 (N_1633,N_1535,N_1585);
or U1634 (N_1634,N_1608,N_1584);
nand U1635 (N_1635,N_1549,N_1505);
and U1636 (N_1636,N_1565,N_1605);
nor U1637 (N_1637,N_1525,N_1502);
and U1638 (N_1638,N_1618,N_1566);
and U1639 (N_1639,N_1530,N_1582);
nand U1640 (N_1640,N_1518,N_1515);
nor U1641 (N_1641,N_1536,N_1602);
nor U1642 (N_1642,N_1531,N_1508);
nor U1643 (N_1643,N_1586,N_1556);
xnor U1644 (N_1644,N_1575,N_1599);
or U1645 (N_1645,N_1519,N_1512);
nand U1646 (N_1646,N_1589,N_1550);
and U1647 (N_1647,N_1583,N_1617);
nand U1648 (N_1648,N_1568,N_1522);
nor U1649 (N_1649,N_1514,N_1609);
or U1650 (N_1650,N_1545,N_1563);
nor U1651 (N_1651,N_1613,N_1615);
nand U1652 (N_1652,N_1521,N_1595);
and U1653 (N_1653,N_1520,N_1580);
xor U1654 (N_1654,N_1607,N_1534);
xor U1655 (N_1655,N_1574,N_1537);
and U1656 (N_1656,N_1572,N_1576);
and U1657 (N_1657,N_1559,N_1513);
or U1658 (N_1658,N_1587,N_1564);
xor U1659 (N_1659,N_1501,N_1540);
xor U1660 (N_1660,N_1593,N_1523);
or U1661 (N_1661,N_1504,N_1555);
nand U1662 (N_1662,N_1578,N_1528);
nor U1663 (N_1663,N_1546,N_1571);
nand U1664 (N_1664,N_1569,N_1529);
or U1665 (N_1665,N_1551,N_1567);
and U1666 (N_1666,N_1538,N_1621);
nand U1667 (N_1667,N_1561,N_1510);
nor U1668 (N_1668,N_1570,N_1524);
nor U1669 (N_1669,N_1624,N_1543);
nor U1670 (N_1670,N_1622,N_1511);
and U1671 (N_1671,N_1600,N_1610);
xor U1672 (N_1672,N_1616,N_1590);
or U1673 (N_1673,N_1579,N_1588);
or U1674 (N_1674,N_1547,N_1553);
xor U1675 (N_1675,N_1500,N_1533);
nand U1676 (N_1676,N_1558,N_1527);
nor U1677 (N_1677,N_1507,N_1581);
xor U1678 (N_1678,N_1516,N_1542);
nor U1679 (N_1679,N_1544,N_1603);
xor U1680 (N_1680,N_1509,N_1623);
xnor U1681 (N_1681,N_1573,N_1594);
nor U1682 (N_1682,N_1557,N_1598);
nand U1683 (N_1683,N_1560,N_1503);
xnor U1684 (N_1684,N_1552,N_1548);
or U1685 (N_1685,N_1591,N_1562);
nand U1686 (N_1686,N_1604,N_1506);
and U1687 (N_1687,N_1601,N_1504);
nand U1688 (N_1688,N_1585,N_1608);
and U1689 (N_1689,N_1508,N_1527);
nand U1690 (N_1690,N_1562,N_1536);
and U1691 (N_1691,N_1548,N_1593);
nand U1692 (N_1692,N_1516,N_1536);
nor U1693 (N_1693,N_1511,N_1615);
nor U1694 (N_1694,N_1606,N_1561);
and U1695 (N_1695,N_1571,N_1590);
nand U1696 (N_1696,N_1600,N_1590);
and U1697 (N_1697,N_1569,N_1533);
or U1698 (N_1698,N_1552,N_1553);
and U1699 (N_1699,N_1591,N_1589);
xor U1700 (N_1700,N_1603,N_1553);
or U1701 (N_1701,N_1511,N_1560);
nand U1702 (N_1702,N_1558,N_1521);
or U1703 (N_1703,N_1508,N_1620);
or U1704 (N_1704,N_1535,N_1594);
and U1705 (N_1705,N_1527,N_1532);
or U1706 (N_1706,N_1624,N_1513);
xnor U1707 (N_1707,N_1555,N_1577);
and U1708 (N_1708,N_1528,N_1529);
or U1709 (N_1709,N_1620,N_1592);
xnor U1710 (N_1710,N_1569,N_1526);
nor U1711 (N_1711,N_1520,N_1559);
xor U1712 (N_1712,N_1506,N_1575);
nor U1713 (N_1713,N_1566,N_1587);
nor U1714 (N_1714,N_1581,N_1548);
nor U1715 (N_1715,N_1532,N_1561);
nor U1716 (N_1716,N_1537,N_1528);
xnor U1717 (N_1717,N_1509,N_1557);
nand U1718 (N_1718,N_1611,N_1614);
and U1719 (N_1719,N_1515,N_1614);
or U1720 (N_1720,N_1581,N_1561);
xor U1721 (N_1721,N_1519,N_1542);
nor U1722 (N_1722,N_1575,N_1609);
nor U1723 (N_1723,N_1553,N_1611);
nor U1724 (N_1724,N_1606,N_1520);
nand U1725 (N_1725,N_1554,N_1572);
xnor U1726 (N_1726,N_1544,N_1614);
nor U1727 (N_1727,N_1543,N_1588);
or U1728 (N_1728,N_1588,N_1623);
or U1729 (N_1729,N_1501,N_1521);
xnor U1730 (N_1730,N_1535,N_1552);
nor U1731 (N_1731,N_1562,N_1569);
xnor U1732 (N_1732,N_1621,N_1558);
nor U1733 (N_1733,N_1508,N_1590);
or U1734 (N_1734,N_1549,N_1597);
nor U1735 (N_1735,N_1620,N_1519);
nor U1736 (N_1736,N_1524,N_1531);
nor U1737 (N_1737,N_1596,N_1534);
nor U1738 (N_1738,N_1614,N_1605);
or U1739 (N_1739,N_1511,N_1592);
nand U1740 (N_1740,N_1566,N_1529);
nand U1741 (N_1741,N_1536,N_1577);
or U1742 (N_1742,N_1586,N_1523);
or U1743 (N_1743,N_1611,N_1530);
and U1744 (N_1744,N_1588,N_1567);
nand U1745 (N_1745,N_1509,N_1622);
xnor U1746 (N_1746,N_1539,N_1594);
or U1747 (N_1747,N_1559,N_1569);
xor U1748 (N_1748,N_1590,N_1592);
and U1749 (N_1749,N_1576,N_1585);
or U1750 (N_1750,N_1665,N_1652);
or U1751 (N_1751,N_1688,N_1659);
nand U1752 (N_1752,N_1731,N_1747);
xor U1753 (N_1753,N_1713,N_1668);
or U1754 (N_1754,N_1630,N_1653);
xor U1755 (N_1755,N_1667,N_1692);
xnor U1756 (N_1756,N_1661,N_1672);
nand U1757 (N_1757,N_1744,N_1631);
and U1758 (N_1758,N_1735,N_1650);
nor U1759 (N_1759,N_1651,N_1682);
nor U1760 (N_1760,N_1640,N_1742);
or U1761 (N_1761,N_1723,N_1629);
nor U1762 (N_1762,N_1626,N_1724);
and U1763 (N_1763,N_1728,N_1647);
and U1764 (N_1764,N_1648,N_1725);
nand U1765 (N_1765,N_1703,N_1686);
and U1766 (N_1766,N_1704,N_1736);
or U1767 (N_1767,N_1680,N_1656);
or U1768 (N_1768,N_1709,N_1637);
and U1769 (N_1769,N_1722,N_1673);
xor U1770 (N_1770,N_1649,N_1628);
xnor U1771 (N_1771,N_1700,N_1732);
nand U1772 (N_1772,N_1730,N_1697);
nor U1773 (N_1773,N_1642,N_1702);
nand U1774 (N_1774,N_1739,N_1726);
xnor U1775 (N_1775,N_1707,N_1727);
nor U1776 (N_1776,N_1664,N_1710);
nand U1777 (N_1777,N_1689,N_1643);
or U1778 (N_1778,N_1729,N_1632);
xnor U1779 (N_1779,N_1641,N_1633);
nor U1780 (N_1780,N_1658,N_1695);
and U1781 (N_1781,N_1654,N_1683);
nor U1782 (N_1782,N_1737,N_1740);
or U1783 (N_1783,N_1693,N_1687);
nor U1784 (N_1784,N_1645,N_1717);
xnor U1785 (N_1785,N_1743,N_1639);
or U1786 (N_1786,N_1663,N_1635);
or U1787 (N_1787,N_1675,N_1699);
nor U1788 (N_1788,N_1734,N_1711);
nor U1789 (N_1789,N_1655,N_1705);
xnor U1790 (N_1790,N_1634,N_1712);
xor U1791 (N_1791,N_1746,N_1636);
nand U1792 (N_1792,N_1627,N_1716);
xor U1793 (N_1793,N_1741,N_1748);
xor U1794 (N_1794,N_1646,N_1715);
or U1795 (N_1795,N_1677,N_1733);
and U1796 (N_1796,N_1660,N_1745);
nor U1797 (N_1797,N_1662,N_1690);
nand U1798 (N_1798,N_1681,N_1684);
or U1799 (N_1799,N_1701,N_1698);
or U1800 (N_1800,N_1670,N_1657);
or U1801 (N_1801,N_1679,N_1676);
nor U1802 (N_1802,N_1738,N_1638);
nor U1803 (N_1803,N_1706,N_1749);
nor U1804 (N_1804,N_1721,N_1671);
nand U1805 (N_1805,N_1708,N_1691);
nand U1806 (N_1806,N_1644,N_1678);
nor U1807 (N_1807,N_1714,N_1696);
or U1808 (N_1808,N_1685,N_1694);
xor U1809 (N_1809,N_1720,N_1666);
xor U1810 (N_1810,N_1625,N_1674);
and U1811 (N_1811,N_1719,N_1718);
and U1812 (N_1812,N_1669,N_1715);
nand U1813 (N_1813,N_1686,N_1712);
nand U1814 (N_1814,N_1654,N_1645);
and U1815 (N_1815,N_1715,N_1736);
xnor U1816 (N_1816,N_1709,N_1711);
nor U1817 (N_1817,N_1732,N_1660);
xor U1818 (N_1818,N_1678,N_1641);
and U1819 (N_1819,N_1696,N_1717);
nand U1820 (N_1820,N_1728,N_1683);
and U1821 (N_1821,N_1645,N_1709);
and U1822 (N_1822,N_1710,N_1679);
nand U1823 (N_1823,N_1739,N_1662);
or U1824 (N_1824,N_1729,N_1658);
nor U1825 (N_1825,N_1674,N_1671);
and U1826 (N_1826,N_1716,N_1719);
nor U1827 (N_1827,N_1672,N_1721);
nor U1828 (N_1828,N_1679,N_1711);
and U1829 (N_1829,N_1646,N_1700);
or U1830 (N_1830,N_1673,N_1743);
nand U1831 (N_1831,N_1735,N_1728);
nor U1832 (N_1832,N_1715,N_1668);
nand U1833 (N_1833,N_1651,N_1649);
xor U1834 (N_1834,N_1681,N_1735);
nor U1835 (N_1835,N_1719,N_1641);
nor U1836 (N_1836,N_1646,N_1748);
xor U1837 (N_1837,N_1714,N_1718);
xnor U1838 (N_1838,N_1745,N_1648);
nand U1839 (N_1839,N_1731,N_1628);
nand U1840 (N_1840,N_1641,N_1716);
nand U1841 (N_1841,N_1718,N_1672);
nor U1842 (N_1842,N_1718,N_1660);
nor U1843 (N_1843,N_1647,N_1635);
xnor U1844 (N_1844,N_1688,N_1654);
nor U1845 (N_1845,N_1680,N_1668);
nor U1846 (N_1846,N_1662,N_1683);
nand U1847 (N_1847,N_1629,N_1727);
and U1848 (N_1848,N_1665,N_1669);
or U1849 (N_1849,N_1637,N_1708);
and U1850 (N_1850,N_1679,N_1745);
nand U1851 (N_1851,N_1661,N_1694);
nand U1852 (N_1852,N_1672,N_1643);
xnor U1853 (N_1853,N_1746,N_1652);
xnor U1854 (N_1854,N_1729,N_1691);
nor U1855 (N_1855,N_1703,N_1732);
nand U1856 (N_1856,N_1712,N_1649);
nor U1857 (N_1857,N_1680,N_1672);
and U1858 (N_1858,N_1698,N_1647);
or U1859 (N_1859,N_1733,N_1634);
nor U1860 (N_1860,N_1685,N_1675);
or U1861 (N_1861,N_1640,N_1701);
xnor U1862 (N_1862,N_1709,N_1655);
xor U1863 (N_1863,N_1646,N_1705);
nand U1864 (N_1864,N_1676,N_1744);
xor U1865 (N_1865,N_1683,N_1631);
xor U1866 (N_1866,N_1738,N_1703);
xnor U1867 (N_1867,N_1706,N_1694);
nor U1868 (N_1868,N_1718,N_1628);
nand U1869 (N_1869,N_1715,N_1657);
xnor U1870 (N_1870,N_1711,N_1704);
xor U1871 (N_1871,N_1661,N_1668);
and U1872 (N_1872,N_1650,N_1744);
xor U1873 (N_1873,N_1631,N_1635);
and U1874 (N_1874,N_1711,N_1628);
nand U1875 (N_1875,N_1817,N_1846);
and U1876 (N_1876,N_1750,N_1804);
nor U1877 (N_1877,N_1873,N_1765);
and U1878 (N_1878,N_1775,N_1823);
and U1879 (N_1879,N_1778,N_1808);
xnor U1880 (N_1880,N_1798,N_1790);
nor U1881 (N_1881,N_1776,N_1868);
nor U1882 (N_1882,N_1760,N_1753);
and U1883 (N_1883,N_1856,N_1828);
xnor U1884 (N_1884,N_1865,N_1872);
nor U1885 (N_1885,N_1763,N_1807);
nor U1886 (N_1886,N_1767,N_1847);
and U1887 (N_1887,N_1841,N_1803);
nand U1888 (N_1888,N_1770,N_1800);
or U1889 (N_1889,N_1801,N_1764);
nand U1890 (N_1890,N_1788,N_1810);
or U1891 (N_1891,N_1758,N_1831);
and U1892 (N_1892,N_1786,N_1777);
nand U1893 (N_1893,N_1843,N_1799);
nand U1894 (N_1894,N_1862,N_1858);
nand U1895 (N_1895,N_1853,N_1867);
nand U1896 (N_1896,N_1866,N_1837);
and U1897 (N_1897,N_1848,N_1791);
nor U1898 (N_1898,N_1755,N_1757);
and U1899 (N_1899,N_1754,N_1797);
xnor U1900 (N_1900,N_1827,N_1871);
nand U1901 (N_1901,N_1766,N_1839);
or U1902 (N_1902,N_1840,N_1849);
nor U1903 (N_1903,N_1864,N_1819);
xor U1904 (N_1904,N_1812,N_1783);
xor U1905 (N_1905,N_1851,N_1814);
nand U1906 (N_1906,N_1785,N_1834);
nor U1907 (N_1907,N_1769,N_1779);
nor U1908 (N_1908,N_1870,N_1838);
nor U1909 (N_1909,N_1772,N_1829);
xor U1910 (N_1910,N_1771,N_1751);
nand U1911 (N_1911,N_1855,N_1822);
nor U1912 (N_1912,N_1759,N_1832);
xor U1913 (N_1913,N_1821,N_1869);
nor U1914 (N_1914,N_1780,N_1860);
nor U1915 (N_1915,N_1802,N_1781);
and U1916 (N_1916,N_1752,N_1813);
nor U1917 (N_1917,N_1805,N_1815);
or U1918 (N_1918,N_1793,N_1784);
nor U1919 (N_1919,N_1773,N_1833);
or U1920 (N_1920,N_1825,N_1842);
and U1921 (N_1921,N_1768,N_1796);
and U1922 (N_1922,N_1835,N_1874);
and U1923 (N_1923,N_1756,N_1854);
nor U1924 (N_1924,N_1850,N_1762);
nor U1925 (N_1925,N_1836,N_1824);
and U1926 (N_1926,N_1818,N_1859);
xnor U1927 (N_1927,N_1844,N_1809);
xor U1928 (N_1928,N_1795,N_1863);
and U1929 (N_1929,N_1789,N_1774);
or U1930 (N_1930,N_1806,N_1852);
xor U1931 (N_1931,N_1816,N_1826);
and U1932 (N_1932,N_1787,N_1811);
nor U1933 (N_1933,N_1782,N_1761);
nand U1934 (N_1934,N_1857,N_1845);
nand U1935 (N_1935,N_1861,N_1820);
nor U1936 (N_1936,N_1794,N_1830);
or U1937 (N_1937,N_1792,N_1839);
or U1938 (N_1938,N_1829,N_1809);
xor U1939 (N_1939,N_1815,N_1863);
nor U1940 (N_1940,N_1789,N_1858);
and U1941 (N_1941,N_1839,N_1824);
nand U1942 (N_1942,N_1790,N_1842);
nor U1943 (N_1943,N_1813,N_1814);
or U1944 (N_1944,N_1816,N_1837);
xor U1945 (N_1945,N_1765,N_1811);
nand U1946 (N_1946,N_1801,N_1840);
xnor U1947 (N_1947,N_1779,N_1861);
or U1948 (N_1948,N_1789,N_1827);
xor U1949 (N_1949,N_1785,N_1820);
nand U1950 (N_1950,N_1863,N_1775);
xnor U1951 (N_1951,N_1814,N_1788);
nor U1952 (N_1952,N_1802,N_1783);
xnor U1953 (N_1953,N_1870,N_1813);
and U1954 (N_1954,N_1835,N_1763);
nand U1955 (N_1955,N_1868,N_1837);
or U1956 (N_1956,N_1776,N_1855);
or U1957 (N_1957,N_1801,N_1796);
or U1958 (N_1958,N_1865,N_1867);
xnor U1959 (N_1959,N_1773,N_1777);
xnor U1960 (N_1960,N_1797,N_1822);
nor U1961 (N_1961,N_1860,N_1762);
nor U1962 (N_1962,N_1820,N_1790);
and U1963 (N_1963,N_1786,N_1767);
and U1964 (N_1964,N_1803,N_1836);
nand U1965 (N_1965,N_1802,N_1778);
and U1966 (N_1966,N_1798,N_1799);
or U1967 (N_1967,N_1843,N_1860);
and U1968 (N_1968,N_1806,N_1828);
nand U1969 (N_1969,N_1811,N_1846);
xnor U1970 (N_1970,N_1759,N_1857);
nand U1971 (N_1971,N_1847,N_1856);
nor U1972 (N_1972,N_1851,N_1839);
xnor U1973 (N_1973,N_1798,N_1826);
xnor U1974 (N_1974,N_1770,N_1813);
nor U1975 (N_1975,N_1768,N_1769);
nor U1976 (N_1976,N_1852,N_1835);
or U1977 (N_1977,N_1862,N_1849);
and U1978 (N_1978,N_1763,N_1770);
nor U1979 (N_1979,N_1810,N_1864);
xnor U1980 (N_1980,N_1775,N_1764);
and U1981 (N_1981,N_1850,N_1857);
xnor U1982 (N_1982,N_1861,N_1818);
or U1983 (N_1983,N_1838,N_1842);
nand U1984 (N_1984,N_1861,N_1784);
nand U1985 (N_1985,N_1856,N_1762);
xor U1986 (N_1986,N_1786,N_1833);
nor U1987 (N_1987,N_1805,N_1829);
or U1988 (N_1988,N_1785,N_1773);
nand U1989 (N_1989,N_1787,N_1784);
nand U1990 (N_1990,N_1825,N_1786);
nor U1991 (N_1991,N_1843,N_1787);
and U1992 (N_1992,N_1821,N_1784);
xnor U1993 (N_1993,N_1790,N_1846);
nand U1994 (N_1994,N_1751,N_1852);
or U1995 (N_1995,N_1779,N_1781);
xor U1996 (N_1996,N_1874,N_1757);
and U1997 (N_1997,N_1826,N_1792);
nand U1998 (N_1998,N_1835,N_1821);
or U1999 (N_1999,N_1790,N_1825);
nor U2000 (N_2000,N_1954,N_1922);
xnor U2001 (N_2001,N_1953,N_1903);
nor U2002 (N_2002,N_1940,N_1885);
or U2003 (N_2003,N_1875,N_1958);
nand U2004 (N_2004,N_1936,N_1967);
or U2005 (N_2005,N_1892,N_1876);
or U2006 (N_2006,N_1999,N_1923);
nor U2007 (N_2007,N_1884,N_1916);
or U2008 (N_2008,N_1906,N_1889);
xor U2009 (N_2009,N_1969,N_1998);
nor U2010 (N_2010,N_1979,N_1900);
nor U2011 (N_2011,N_1995,N_1890);
and U2012 (N_2012,N_1981,N_1960);
nand U2013 (N_2013,N_1882,N_1942);
or U2014 (N_2014,N_1909,N_1878);
nand U2015 (N_2015,N_1930,N_1913);
nor U2016 (N_2016,N_1898,N_1948);
xnor U2017 (N_2017,N_1919,N_1915);
and U2018 (N_2018,N_1937,N_1896);
xnor U2019 (N_2019,N_1944,N_1907);
xor U2020 (N_2020,N_1991,N_1992);
and U2021 (N_2021,N_1963,N_1893);
xor U2022 (N_2022,N_1881,N_1972);
xnor U2023 (N_2023,N_1888,N_1978);
nor U2024 (N_2024,N_1927,N_1973);
nand U2025 (N_2025,N_1957,N_1897);
xor U2026 (N_2026,N_1966,N_1899);
nand U2027 (N_2027,N_1902,N_1920);
nor U2028 (N_2028,N_1887,N_1941);
and U2029 (N_2029,N_1977,N_1968);
nand U2030 (N_2030,N_1910,N_1933);
or U2031 (N_2031,N_1877,N_1971);
xnor U2032 (N_2032,N_1894,N_1952);
xnor U2033 (N_2033,N_1949,N_1880);
and U2034 (N_2034,N_1895,N_1987);
nand U2035 (N_2035,N_1980,N_1939);
nor U2036 (N_2036,N_1989,N_1962);
and U2037 (N_2037,N_1914,N_1988);
or U2038 (N_2038,N_1946,N_1908);
xor U2039 (N_2039,N_1983,N_1886);
xnor U2040 (N_2040,N_1974,N_1955);
nor U2041 (N_2041,N_1996,N_1932);
and U2042 (N_2042,N_1950,N_1929);
or U2043 (N_2043,N_1883,N_1905);
or U2044 (N_2044,N_1943,N_1951);
or U2045 (N_2045,N_1935,N_1994);
or U2046 (N_2046,N_1984,N_1982);
or U2047 (N_2047,N_1964,N_1901);
xor U2048 (N_2048,N_1985,N_1891);
xor U2049 (N_2049,N_1965,N_1947);
nor U2050 (N_2050,N_1912,N_1961);
and U2051 (N_2051,N_1956,N_1879);
or U2052 (N_2052,N_1970,N_1959);
nor U2053 (N_2053,N_1918,N_1925);
and U2054 (N_2054,N_1911,N_1990);
nor U2055 (N_2055,N_1976,N_1938);
nand U2056 (N_2056,N_1997,N_1917);
nor U2057 (N_2057,N_1986,N_1904);
and U2058 (N_2058,N_1934,N_1931);
or U2059 (N_2059,N_1924,N_1928);
nor U2060 (N_2060,N_1975,N_1945);
xnor U2061 (N_2061,N_1993,N_1921);
or U2062 (N_2062,N_1926,N_1996);
nand U2063 (N_2063,N_1878,N_1966);
xnor U2064 (N_2064,N_1893,N_1930);
nor U2065 (N_2065,N_1883,N_1976);
xnor U2066 (N_2066,N_1984,N_1878);
nor U2067 (N_2067,N_1923,N_1876);
or U2068 (N_2068,N_1937,N_1953);
xnor U2069 (N_2069,N_1886,N_1943);
or U2070 (N_2070,N_1923,N_1935);
nand U2071 (N_2071,N_1975,N_1876);
xor U2072 (N_2072,N_1952,N_1916);
and U2073 (N_2073,N_1982,N_1996);
or U2074 (N_2074,N_1909,N_1897);
xnor U2075 (N_2075,N_1969,N_1980);
xor U2076 (N_2076,N_1910,N_1952);
nor U2077 (N_2077,N_1985,N_1944);
and U2078 (N_2078,N_1952,N_1950);
and U2079 (N_2079,N_1875,N_1887);
xnor U2080 (N_2080,N_1980,N_1944);
nand U2081 (N_2081,N_1916,N_1958);
or U2082 (N_2082,N_1959,N_1978);
nand U2083 (N_2083,N_1943,N_1998);
nand U2084 (N_2084,N_1966,N_1997);
xnor U2085 (N_2085,N_1877,N_1939);
or U2086 (N_2086,N_1981,N_1999);
and U2087 (N_2087,N_1972,N_1921);
nand U2088 (N_2088,N_1961,N_1963);
and U2089 (N_2089,N_1907,N_1997);
or U2090 (N_2090,N_1960,N_1956);
xnor U2091 (N_2091,N_1971,N_1884);
and U2092 (N_2092,N_1904,N_1875);
nand U2093 (N_2093,N_1969,N_1943);
or U2094 (N_2094,N_1973,N_1893);
or U2095 (N_2095,N_1886,N_1967);
nand U2096 (N_2096,N_1988,N_1925);
nor U2097 (N_2097,N_1875,N_1895);
nand U2098 (N_2098,N_1885,N_1907);
and U2099 (N_2099,N_1963,N_1878);
and U2100 (N_2100,N_1920,N_1993);
or U2101 (N_2101,N_1982,N_1917);
or U2102 (N_2102,N_1946,N_1895);
nor U2103 (N_2103,N_1924,N_1886);
and U2104 (N_2104,N_1915,N_1963);
nand U2105 (N_2105,N_1896,N_1955);
xor U2106 (N_2106,N_1990,N_1993);
nand U2107 (N_2107,N_1971,N_1908);
or U2108 (N_2108,N_1985,N_1939);
nand U2109 (N_2109,N_1989,N_1911);
and U2110 (N_2110,N_1989,N_1940);
nor U2111 (N_2111,N_1982,N_1876);
and U2112 (N_2112,N_1892,N_1910);
xor U2113 (N_2113,N_1994,N_1951);
nand U2114 (N_2114,N_1875,N_1947);
xnor U2115 (N_2115,N_1961,N_1905);
xor U2116 (N_2116,N_1887,N_1948);
or U2117 (N_2117,N_1982,N_1903);
xor U2118 (N_2118,N_1982,N_1974);
xor U2119 (N_2119,N_1885,N_1917);
nand U2120 (N_2120,N_1994,N_1890);
or U2121 (N_2121,N_1960,N_1927);
nand U2122 (N_2122,N_1902,N_1926);
nor U2123 (N_2123,N_1908,N_1879);
nor U2124 (N_2124,N_1994,N_1906);
nand U2125 (N_2125,N_2106,N_2028);
and U2126 (N_2126,N_2085,N_2030);
or U2127 (N_2127,N_2069,N_2082);
or U2128 (N_2128,N_2032,N_2081);
xor U2129 (N_2129,N_2061,N_2066);
nor U2130 (N_2130,N_2033,N_2056);
and U2131 (N_2131,N_2046,N_2092);
nand U2132 (N_2132,N_2067,N_2100);
nand U2133 (N_2133,N_2059,N_2015);
xor U2134 (N_2134,N_2121,N_2037);
or U2135 (N_2135,N_2044,N_2041);
and U2136 (N_2136,N_2043,N_2002);
or U2137 (N_2137,N_2076,N_2112);
and U2138 (N_2138,N_2047,N_2019);
and U2139 (N_2139,N_2093,N_2083);
or U2140 (N_2140,N_2089,N_2009);
nand U2141 (N_2141,N_2014,N_2001);
nor U2142 (N_2142,N_2107,N_2039);
xor U2143 (N_2143,N_2024,N_2020);
and U2144 (N_2144,N_2096,N_2074);
xnor U2145 (N_2145,N_2110,N_2016);
or U2146 (N_2146,N_2115,N_2091);
xnor U2147 (N_2147,N_2101,N_2031);
or U2148 (N_2148,N_2124,N_2108);
and U2149 (N_2149,N_2042,N_2049);
and U2150 (N_2150,N_2051,N_2058);
nor U2151 (N_2151,N_2021,N_2109);
nand U2152 (N_2152,N_2045,N_2098);
nand U2153 (N_2153,N_2104,N_2075);
or U2154 (N_2154,N_2084,N_2048);
nand U2155 (N_2155,N_2099,N_2095);
nor U2156 (N_2156,N_2063,N_2065);
and U2157 (N_2157,N_2029,N_2079);
and U2158 (N_2158,N_2114,N_2040);
and U2159 (N_2159,N_2086,N_2027);
nor U2160 (N_2160,N_2022,N_2052);
xnor U2161 (N_2161,N_2113,N_2119);
and U2162 (N_2162,N_2017,N_2006);
xor U2163 (N_2163,N_2034,N_2025);
nand U2164 (N_2164,N_2122,N_2102);
or U2165 (N_2165,N_2068,N_2064);
nand U2166 (N_2166,N_2116,N_2118);
nor U2167 (N_2167,N_2077,N_2062);
xnor U2168 (N_2168,N_2011,N_2120);
nand U2169 (N_2169,N_2055,N_2071);
or U2170 (N_2170,N_2005,N_2111);
and U2171 (N_2171,N_2007,N_2018);
or U2172 (N_2172,N_2097,N_2060);
nand U2173 (N_2173,N_2000,N_2057);
and U2174 (N_2174,N_2078,N_2123);
xnor U2175 (N_2175,N_2010,N_2038);
xor U2176 (N_2176,N_2117,N_2054);
xor U2177 (N_2177,N_2008,N_2073);
nor U2178 (N_2178,N_2105,N_2023);
nand U2179 (N_2179,N_2004,N_2003);
xnor U2180 (N_2180,N_2013,N_2050);
nor U2181 (N_2181,N_2012,N_2087);
and U2182 (N_2182,N_2036,N_2103);
nor U2183 (N_2183,N_2088,N_2053);
and U2184 (N_2184,N_2070,N_2035);
or U2185 (N_2185,N_2026,N_2072);
xnor U2186 (N_2186,N_2094,N_2090);
nand U2187 (N_2187,N_2080,N_2102);
xor U2188 (N_2188,N_2024,N_2005);
xor U2189 (N_2189,N_2068,N_2017);
or U2190 (N_2190,N_2035,N_2018);
and U2191 (N_2191,N_2014,N_2117);
or U2192 (N_2192,N_2056,N_2011);
nor U2193 (N_2193,N_2062,N_2052);
or U2194 (N_2194,N_2081,N_2101);
nand U2195 (N_2195,N_2047,N_2053);
xnor U2196 (N_2196,N_2121,N_2042);
nand U2197 (N_2197,N_2081,N_2048);
xor U2198 (N_2198,N_2086,N_2014);
nand U2199 (N_2199,N_2006,N_2076);
nand U2200 (N_2200,N_2057,N_2121);
nor U2201 (N_2201,N_2021,N_2002);
nand U2202 (N_2202,N_2119,N_2085);
and U2203 (N_2203,N_2097,N_2083);
or U2204 (N_2204,N_2105,N_2024);
xor U2205 (N_2205,N_2093,N_2052);
xor U2206 (N_2206,N_2109,N_2024);
nor U2207 (N_2207,N_2021,N_2026);
nand U2208 (N_2208,N_2022,N_2071);
nand U2209 (N_2209,N_2038,N_2015);
xor U2210 (N_2210,N_2107,N_2091);
xor U2211 (N_2211,N_2108,N_2011);
nor U2212 (N_2212,N_2056,N_2078);
nand U2213 (N_2213,N_2085,N_2089);
or U2214 (N_2214,N_2118,N_2081);
xor U2215 (N_2215,N_2039,N_2070);
and U2216 (N_2216,N_2096,N_2036);
or U2217 (N_2217,N_2120,N_2072);
nor U2218 (N_2218,N_2022,N_2043);
xor U2219 (N_2219,N_2120,N_2099);
and U2220 (N_2220,N_2064,N_2080);
nand U2221 (N_2221,N_2101,N_2088);
nand U2222 (N_2222,N_2106,N_2095);
and U2223 (N_2223,N_2103,N_2072);
nand U2224 (N_2224,N_2009,N_2059);
xnor U2225 (N_2225,N_2087,N_2124);
nor U2226 (N_2226,N_2062,N_2089);
xor U2227 (N_2227,N_2041,N_2103);
xor U2228 (N_2228,N_2090,N_2014);
or U2229 (N_2229,N_2062,N_2117);
and U2230 (N_2230,N_2086,N_2115);
xor U2231 (N_2231,N_2030,N_2071);
or U2232 (N_2232,N_2015,N_2056);
xnor U2233 (N_2233,N_2036,N_2086);
xor U2234 (N_2234,N_2081,N_2024);
and U2235 (N_2235,N_2020,N_2060);
nand U2236 (N_2236,N_2065,N_2103);
and U2237 (N_2237,N_2057,N_2045);
or U2238 (N_2238,N_2074,N_2037);
or U2239 (N_2239,N_2064,N_2062);
or U2240 (N_2240,N_2051,N_2003);
nor U2241 (N_2241,N_2064,N_2066);
nor U2242 (N_2242,N_2074,N_2000);
xor U2243 (N_2243,N_2102,N_2065);
and U2244 (N_2244,N_2122,N_2060);
nor U2245 (N_2245,N_2007,N_2044);
and U2246 (N_2246,N_2030,N_2043);
nor U2247 (N_2247,N_2089,N_2081);
nor U2248 (N_2248,N_2101,N_2096);
or U2249 (N_2249,N_2084,N_2057);
xnor U2250 (N_2250,N_2201,N_2151);
or U2251 (N_2251,N_2127,N_2207);
nor U2252 (N_2252,N_2224,N_2187);
nand U2253 (N_2253,N_2248,N_2163);
nor U2254 (N_2254,N_2190,N_2162);
nor U2255 (N_2255,N_2134,N_2225);
or U2256 (N_2256,N_2130,N_2172);
nor U2257 (N_2257,N_2171,N_2176);
or U2258 (N_2258,N_2136,N_2178);
and U2259 (N_2259,N_2161,N_2218);
xnor U2260 (N_2260,N_2236,N_2189);
or U2261 (N_2261,N_2166,N_2245);
and U2262 (N_2262,N_2237,N_2152);
or U2263 (N_2263,N_2234,N_2202);
and U2264 (N_2264,N_2217,N_2243);
xor U2265 (N_2265,N_2200,N_2148);
and U2266 (N_2266,N_2241,N_2131);
xor U2267 (N_2267,N_2203,N_2181);
and U2268 (N_2268,N_2157,N_2229);
nand U2269 (N_2269,N_2137,N_2167);
and U2270 (N_2270,N_2126,N_2182);
xnor U2271 (N_2271,N_2149,N_2185);
and U2272 (N_2272,N_2139,N_2228);
or U2273 (N_2273,N_2221,N_2219);
xnor U2274 (N_2274,N_2186,N_2220);
or U2275 (N_2275,N_2150,N_2183);
and U2276 (N_2276,N_2193,N_2214);
nor U2277 (N_2277,N_2153,N_2240);
nor U2278 (N_2278,N_2198,N_2154);
nor U2279 (N_2279,N_2208,N_2158);
or U2280 (N_2280,N_2192,N_2128);
or U2281 (N_2281,N_2164,N_2249);
nand U2282 (N_2282,N_2232,N_2179);
nor U2283 (N_2283,N_2125,N_2196);
or U2284 (N_2284,N_2246,N_2197);
and U2285 (N_2285,N_2132,N_2177);
xor U2286 (N_2286,N_2146,N_2147);
nor U2287 (N_2287,N_2211,N_2165);
and U2288 (N_2288,N_2194,N_2235);
nor U2289 (N_2289,N_2231,N_2143);
nand U2290 (N_2290,N_2233,N_2180);
nand U2291 (N_2291,N_2141,N_2173);
xnor U2292 (N_2292,N_2242,N_2213);
nand U2293 (N_2293,N_2212,N_2174);
xor U2294 (N_2294,N_2239,N_2168);
and U2295 (N_2295,N_2204,N_2199);
nand U2296 (N_2296,N_2135,N_2223);
xnor U2297 (N_2297,N_2238,N_2227);
nand U2298 (N_2298,N_2195,N_2170);
xor U2299 (N_2299,N_2138,N_2215);
xor U2300 (N_2300,N_2206,N_2247);
nor U2301 (N_2301,N_2159,N_2184);
nand U2302 (N_2302,N_2210,N_2175);
nor U2303 (N_2303,N_2188,N_2133);
xnor U2304 (N_2304,N_2155,N_2191);
or U2305 (N_2305,N_2156,N_2140);
or U2306 (N_2306,N_2169,N_2160);
xnor U2307 (N_2307,N_2145,N_2222);
or U2308 (N_2308,N_2230,N_2205);
nor U2309 (N_2309,N_2129,N_2244);
or U2310 (N_2310,N_2216,N_2226);
xnor U2311 (N_2311,N_2209,N_2144);
nor U2312 (N_2312,N_2142,N_2151);
and U2313 (N_2313,N_2141,N_2224);
and U2314 (N_2314,N_2133,N_2125);
nand U2315 (N_2315,N_2130,N_2234);
xor U2316 (N_2316,N_2209,N_2242);
xor U2317 (N_2317,N_2224,N_2218);
nor U2318 (N_2318,N_2243,N_2183);
nand U2319 (N_2319,N_2170,N_2126);
or U2320 (N_2320,N_2156,N_2185);
or U2321 (N_2321,N_2147,N_2151);
nor U2322 (N_2322,N_2208,N_2200);
xor U2323 (N_2323,N_2214,N_2211);
xor U2324 (N_2324,N_2229,N_2198);
or U2325 (N_2325,N_2160,N_2161);
xor U2326 (N_2326,N_2226,N_2161);
and U2327 (N_2327,N_2162,N_2248);
nor U2328 (N_2328,N_2163,N_2145);
xor U2329 (N_2329,N_2243,N_2246);
xnor U2330 (N_2330,N_2166,N_2169);
or U2331 (N_2331,N_2232,N_2167);
nand U2332 (N_2332,N_2144,N_2237);
and U2333 (N_2333,N_2137,N_2160);
nand U2334 (N_2334,N_2152,N_2211);
xnor U2335 (N_2335,N_2154,N_2125);
xor U2336 (N_2336,N_2241,N_2164);
xnor U2337 (N_2337,N_2133,N_2136);
nor U2338 (N_2338,N_2243,N_2240);
xor U2339 (N_2339,N_2249,N_2161);
or U2340 (N_2340,N_2193,N_2232);
nand U2341 (N_2341,N_2219,N_2146);
or U2342 (N_2342,N_2186,N_2160);
nand U2343 (N_2343,N_2243,N_2147);
nor U2344 (N_2344,N_2203,N_2144);
and U2345 (N_2345,N_2211,N_2134);
nor U2346 (N_2346,N_2224,N_2173);
xor U2347 (N_2347,N_2204,N_2129);
and U2348 (N_2348,N_2195,N_2176);
and U2349 (N_2349,N_2163,N_2146);
nand U2350 (N_2350,N_2165,N_2199);
nand U2351 (N_2351,N_2171,N_2218);
nand U2352 (N_2352,N_2195,N_2197);
or U2353 (N_2353,N_2127,N_2220);
and U2354 (N_2354,N_2131,N_2210);
and U2355 (N_2355,N_2180,N_2249);
xnor U2356 (N_2356,N_2181,N_2193);
or U2357 (N_2357,N_2174,N_2136);
and U2358 (N_2358,N_2182,N_2135);
nor U2359 (N_2359,N_2241,N_2150);
or U2360 (N_2360,N_2199,N_2212);
or U2361 (N_2361,N_2173,N_2236);
nor U2362 (N_2362,N_2139,N_2213);
or U2363 (N_2363,N_2183,N_2160);
xnor U2364 (N_2364,N_2128,N_2172);
nand U2365 (N_2365,N_2213,N_2143);
xnor U2366 (N_2366,N_2138,N_2203);
nand U2367 (N_2367,N_2136,N_2160);
nor U2368 (N_2368,N_2131,N_2159);
nand U2369 (N_2369,N_2227,N_2193);
nor U2370 (N_2370,N_2237,N_2219);
and U2371 (N_2371,N_2204,N_2164);
xnor U2372 (N_2372,N_2235,N_2246);
or U2373 (N_2373,N_2177,N_2236);
or U2374 (N_2374,N_2150,N_2205);
or U2375 (N_2375,N_2358,N_2301);
or U2376 (N_2376,N_2359,N_2370);
or U2377 (N_2377,N_2268,N_2282);
nand U2378 (N_2378,N_2251,N_2250);
and U2379 (N_2379,N_2325,N_2317);
or U2380 (N_2380,N_2351,N_2277);
nand U2381 (N_2381,N_2264,N_2265);
and U2382 (N_2382,N_2321,N_2292);
xor U2383 (N_2383,N_2273,N_2324);
and U2384 (N_2384,N_2255,N_2304);
nor U2385 (N_2385,N_2363,N_2340);
and U2386 (N_2386,N_2295,N_2360);
and U2387 (N_2387,N_2356,N_2322);
nand U2388 (N_2388,N_2323,N_2367);
nor U2389 (N_2389,N_2327,N_2372);
and U2390 (N_2390,N_2300,N_2320);
and U2391 (N_2391,N_2281,N_2289);
xor U2392 (N_2392,N_2298,N_2349);
and U2393 (N_2393,N_2344,N_2280);
or U2394 (N_2394,N_2361,N_2297);
nor U2395 (N_2395,N_2253,N_2318);
or U2396 (N_2396,N_2326,N_2315);
and U2397 (N_2397,N_2328,N_2284);
nor U2398 (N_2398,N_2330,N_2316);
xnor U2399 (N_2399,N_2336,N_2256);
nor U2400 (N_2400,N_2337,N_2369);
xor U2401 (N_2401,N_2314,N_2275);
or U2402 (N_2402,N_2262,N_2364);
and U2403 (N_2403,N_2306,N_2259);
nor U2404 (N_2404,N_2254,N_2341);
nand U2405 (N_2405,N_2354,N_2270);
or U2406 (N_2406,N_2258,N_2371);
or U2407 (N_2407,N_2348,N_2335);
nor U2408 (N_2408,N_2342,N_2290);
xnor U2409 (N_2409,N_2332,N_2261);
or U2410 (N_2410,N_2345,N_2374);
or U2411 (N_2411,N_2307,N_2299);
xor U2412 (N_2412,N_2338,N_2339);
or U2413 (N_2413,N_2308,N_2312);
nand U2414 (N_2414,N_2286,N_2334);
and U2415 (N_2415,N_2287,N_2285);
or U2416 (N_2416,N_2346,N_2350);
nor U2417 (N_2417,N_2352,N_2293);
xor U2418 (N_2418,N_2288,N_2365);
nand U2419 (N_2419,N_2291,N_2303);
xor U2420 (N_2420,N_2357,N_2329);
or U2421 (N_2421,N_2319,N_2294);
nor U2422 (N_2422,N_2310,N_2260);
nor U2423 (N_2423,N_2278,N_2343);
nand U2424 (N_2424,N_2269,N_2302);
nand U2425 (N_2425,N_2274,N_2309);
nand U2426 (N_2426,N_2276,N_2368);
xnor U2427 (N_2427,N_2267,N_2296);
nor U2428 (N_2428,N_2331,N_2311);
xor U2429 (N_2429,N_2366,N_2305);
and U2430 (N_2430,N_2257,N_2266);
xnor U2431 (N_2431,N_2353,N_2347);
or U2432 (N_2432,N_2373,N_2271);
or U2433 (N_2433,N_2263,N_2333);
nand U2434 (N_2434,N_2252,N_2283);
nand U2435 (N_2435,N_2355,N_2362);
nor U2436 (N_2436,N_2313,N_2279);
and U2437 (N_2437,N_2272,N_2299);
nor U2438 (N_2438,N_2315,N_2297);
nor U2439 (N_2439,N_2362,N_2329);
and U2440 (N_2440,N_2360,N_2349);
nor U2441 (N_2441,N_2341,N_2260);
and U2442 (N_2442,N_2276,N_2354);
xor U2443 (N_2443,N_2314,N_2335);
or U2444 (N_2444,N_2314,N_2311);
xnor U2445 (N_2445,N_2312,N_2314);
and U2446 (N_2446,N_2337,N_2299);
nand U2447 (N_2447,N_2311,N_2254);
nand U2448 (N_2448,N_2357,N_2288);
nor U2449 (N_2449,N_2335,N_2255);
or U2450 (N_2450,N_2277,N_2264);
and U2451 (N_2451,N_2300,N_2283);
or U2452 (N_2452,N_2302,N_2324);
and U2453 (N_2453,N_2352,N_2349);
and U2454 (N_2454,N_2317,N_2291);
or U2455 (N_2455,N_2307,N_2334);
or U2456 (N_2456,N_2374,N_2358);
nor U2457 (N_2457,N_2334,N_2305);
nor U2458 (N_2458,N_2366,N_2336);
or U2459 (N_2459,N_2336,N_2339);
and U2460 (N_2460,N_2367,N_2280);
and U2461 (N_2461,N_2307,N_2287);
or U2462 (N_2462,N_2263,N_2364);
nand U2463 (N_2463,N_2271,N_2297);
or U2464 (N_2464,N_2256,N_2272);
or U2465 (N_2465,N_2357,N_2327);
or U2466 (N_2466,N_2258,N_2282);
nor U2467 (N_2467,N_2323,N_2317);
and U2468 (N_2468,N_2319,N_2348);
or U2469 (N_2469,N_2269,N_2266);
nand U2470 (N_2470,N_2282,N_2374);
or U2471 (N_2471,N_2351,N_2294);
nand U2472 (N_2472,N_2271,N_2265);
nand U2473 (N_2473,N_2306,N_2267);
nor U2474 (N_2474,N_2261,N_2277);
or U2475 (N_2475,N_2276,N_2328);
and U2476 (N_2476,N_2366,N_2347);
or U2477 (N_2477,N_2311,N_2266);
or U2478 (N_2478,N_2261,N_2328);
nand U2479 (N_2479,N_2355,N_2265);
nand U2480 (N_2480,N_2266,N_2334);
xnor U2481 (N_2481,N_2301,N_2347);
nand U2482 (N_2482,N_2361,N_2255);
or U2483 (N_2483,N_2276,N_2275);
nand U2484 (N_2484,N_2366,N_2286);
and U2485 (N_2485,N_2264,N_2322);
and U2486 (N_2486,N_2340,N_2374);
or U2487 (N_2487,N_2354,N_2373);
xnor U2488 (N_2488,N_2337,N_2368);
or U2489 (N_2489,N_2286,N_2332);
nand U2490 (N_2490,N_2344,N_2257);
and U2491 (N_2491,N_2261,N_2306);
or U2492 (N_2492,N_2280,N_2270);
nor U2493 (N_2493,N_2259,N_2256);
or U2494 (N_2494,N_2362,N_2327);
or U2495 (N_2495,N_2261,N_2331);
and U2496 (N_2496,N_2330,N_2262);
nor U2497 (N_2497,N_2374,N_2297);
nand U2498 (N_2498,N_2266,N_2284);
nand U2499 (N_2499,N_2342,N_2348);
nor U2500 (N_2500,N_2409,N_2410);
nor U2501 (N_2501,N_2425,N_2403);
nand U2502 (N_2502,N_2464,N_2468);
and U2503 (N_2503,N_2487,N_2417);
xnor U2504 (N_2504,N_2455,N_2498);
or U2505 (N_2505,N_2477,N_2492);
nor U2506 (N_2506,N_2480,N_2382);
and U2507 (N_2507,N_2454,N_2438);
or U2508 (N_2508,N_2448,N_2408);
and U2509 (N_2509,N_2437,N_2489);
or U2510 (N_2510,N_2424,N_2377);
xor U2511 (N_2511,N_2427,N_2385);
nand U2512 (N_2512,N_2460,N_2391);
and U2513 (N_2513,N_2461,N_2444);
and U2514 (N_2514,N_2466,N_2432);
or U2515 (N_2515,N_2490,N_2384);
or U2516 (N_2516,N_2485,N_2423);
nor U2517 (N_2517,N_2411,N_2428);
xnor U2518 (N_2518,N_2493,N_2462);
xor U2519 (N_2519,N_2484,N_2440);
nor U2520 (N_2520,N_2435,N_2415);
or U2521 (N_2521,N_2421,N_2416);
and U2522 (N_2522,N_2482,N_2459);
and U2523 (N_2523,N_2451,N_2407);
nand U2524 (N_2524,N_2447,N_2479);
xor U2525 (N_2525,N_2394,N_2449);
and U2526 (N_2526,N_2426,N_2474);
nor U2527 (N_2527,N_2483,N_2475);
xnor U2528 (N_2528,N_2433,N_2481);
or U2529 (N_2529,N_2496,N_2497);
nor U2530 (N_2530,N_2422,N_2376);
or U2531 (N_2531,N_2388,N_2381);
nor U2532 (N_2532,N_2414,N_2406);
xnor U2533 (N_2533,N_2495,N_2397);
and U2534 (N_2534,N_2456,N_2465);
nor U2535 (N_2535,N_2419,N_2491);
or U2536 (N_2536,N_2445,N_2472);
or U2537 (N_2537,N_2386,N_2418);
or U2538 (N_2538,N_2441,N_2389);
nand U2539 (N_2539,N_2442,N_2458);
nor U2540 (N_2540,N_2393,N_2486);
nor U2541 (N_2541,N_2413,N_2404);
and U2542 (N_2542,N_2446,N_2399);
and U2543 (N_2543,N_2430,N_2434);
nor U2544 (N_2544,N_2379,N_2405);
or U2545 (N_2545,N_2450,N_2471);
nand U2546 (N_2546,N_2443,N_2402);
nand U2547 (N_2547,N_2383,N_2452);
nor U2548 (N_2548,N_2412,N_2436);
xnor U2549 (N_2549,N_2387,N_2453);
nor U2550 (N_2550,N_2398,N_2499);
or U2551 (N_2551,N_2431,N_2478);
xnor U2552 (N_2552,N_2473,N_2457);
nand U2553 (N_2553,N_2395,N_2476);
and U2554 (N_2554,N_2390,N_2469);
xor U2555 (N_2555,N_2396,N_2378);
or U2556 (N_2556,N_2488,N_2401);
xnor U2557 (N_2557,N_2392,N_2439);
xnor U2558 (N_2558,N_2463,N_2470);
and U2559 (N_2559,N_2400,N_2375);
and U2560 (N_2560,N_2420,N_2467);
xnor U2561 (N_2561,N_2429,N_2380);
and U2562 (N_2562,N_2494,N_2462);
or U2563 (N_2563,N_2398,N_2473);
nand U2564 (N_2564,N_2388,N_2489);
or U2565 (N_2565,N_2451,N_2478);
nor U2566 (N_2566,N_2379,N_2486);
nand U2567 (N_2567,N_2413,N_2420);
and U2568 (N_2568,N_2443,N_2445);
or U2569 (N_2569,N_2463,N_2479);
xor U2570 (N_2570,N_2405,N_2486);
nand U2571 (N_2571,N_2484,N_2396);
or U2572 (N_2572,N_2396,N_2454);
xnor U2573 (N_2573,N_2388,N_2494);
xor U2574 (N_2574,N_2414,N_2412);
and U2575 (N_2575,N_2452,N_2407);
nor U2576 (N_2576,N_2377,N_2396);
nand U2577 (N_2577,N_2419,N_2446);
xor U2578 (N_2578,N_2434,N_2493);
xor U2579 (N_2579,N_2452,N_2422);
xnor U2580 (N_2580,N_2444,N_2479);
or U2581 (N_2581,N_2419,N_2461);
and U2582 (N_2582,N_2448,N_2493);
and U2583 (N_2583,N_2470,N_2383);
nor U2584 (N_2584,N_2477,N_2437);
and U2585 (N_2585,N_2474,N_2468);
xor U2586 (N_2586,N_2488,N_2435);
xnor U2587 (N_2587,N_2392,N_2412);
nand U2588 (N_2588,N_2437,N_2404);
or U2589 (N_2589,N_2468,N_2400);
nor U2590 (N_2590,N_2379,N_2420);
xor U2591 (N_2591,N_2377,N_2472);
xnor U2592 (N_2592,N_2377,N_2403);
xnor U2593 (N_2593,N_2479,N_2494);
or U2594 (N_2594,N_2378,N_2492);
xnor U2595 (N_2595,N_2432,N_2423);
and U2596 (N_2596,N_2475,N_2465);
nand U2597 (N_2597,N_2440,N_2489);
nor U2598 (N_2598,N_2485,N_2467);
or U2599 (N_2599,N_2466,N_2447);
xnor U2600 (N_2600,N_2440,N_2486);
xnor U2601 (N_2601,N_2490,N_2493);
and U2602 (N_2602,N_2376,N_2455);
nand U2603 (N_2603,N_2451,N_2385);
and U2604 (N_2604,N_2443,N_2469);
xor U2605 (N_2605,N_2379,N_2438);
and U2606 (N_2606,N_2454,N_2386);
xor U2607 (N_2607,N_2377,N_2406);
or U2608 (N_2608,N_2427,N_2480);
xnor U2609 (N_2609,N_2391,N_2424);
xnor U2610 (N_2610,N_2402,N_2410);
or U2611 (N_2611,N_2386,N_2387);
nand U2612 (N_2612,N_2400,N_2429);
xnor U2613 (N_2613,N_2398,N_2388);
xnor U2614 (N_2614,N_2477,N_2462);
or U2615 (N_2615,N_2398,N_2401);
xnor U2616 (N_2616,N_2446,N_2425);
nand U2617 (N_2617,N_2385,N_2482);
nand U2618 (N_2618,N_2468,N_2495);
xor U2619 (N_2619,N_2471,N_2421);
nand U2620 (N_2620,N_2441,N_2418);
xor U2621 (N_2621,N_2436,N_2483);
xnor U2622 (N_2622,N_2462,N_2482);
nor U2623 (N_2623,N_2455,N_2446);
or U2624 (N_2624,N_2419,N_2441);
or U2625 (N_2625,N_2543,N_2611);
xor U2626 (N_2626,N_2559,N_2605);
nand U2627 (N_2627,N_2554,N_2528);
nand U2628 (N_2628,N_2585,N_2539);
or U2629 (N_2629,N_2575,N_2558);
or U2630 (N_2630,N_2581,N_2566);
xor U2631 (N_2631,N_2522,N_2599);
and U2632 (N_2632,N_2608,N_2572);
nor U2633 (N_2633,N_2580,N_2565);
nor U2634 (N_2634,N_2613,N_2513);
nor U2635 (N_2635,N_2519,N_2541);
and U2636 (N_2636,N_2531,N_2597);
and U2637 (N_2637,N_2560,N_2537);
nand U2638 (N_2638,N_2591,N_2600);
and U2639 (N_2639,N_2576,N_2507);
nor U2640 (N_2640,N_2593,N_2500);
nor U2641 (N_2641,N_2502,N_2587);
and U2642 (N_2642,N_2556,N_2515);
and U2643 (N_2643,N_2508,N_2609);
or U2644 (N_2644,N_2548,N_2529);
or U2645 (N_2645,N_2551,N_2586);
and U2646 (N_2646,N_2540,N_2533);
nor U2647 (N_2647,N_2589,N_2530);
and U2648 (N_2648,N_2544,N_2618);
and U2649 (N_2649,N_2623,N_2506);
nor U2650 (N_2650,N_2567,N_2574);
nor U2651 (N_2651,N_2536,N_2616);
or U2652 (N_2652,N_2619,N_2579);
or U2653 (N_2653,N_2557,N_2620);
or U2654 (N_2654,N_2523,N_2546);
or U2655 (N_2655,N_2521,N_2538);
nand U2656 (N_2656,N_2518,N_2520);
xor U2657 (N_2657,N_2612,N_2516);
xor U2658 (N_2658,N_2511,N_2583);
and U2659 (N_2659,N_2527,N_2514);
nand U2660 (N_2660,N_2562,N_2561);
nand U2661 (N_2661,N_2532,N_2526);
nor U2662 (N_2662,N_2525,N_2582);
nor U2663 (N_2663,N_2553,N_2596);
nor U2664 (N_2664,N_2503,N_2577);
xor U2665 (N_2665,N_2501,N_2555);
xnor U2666 (N_2666,N_2510,N_2590);
xor U2667 (N_2667,N_2598,N_2504);
and U2668 (N_2668,N_2509,N_2517);
or U2669 (N_2669,N_2569,N_2550);
nand U2670 (N_2670,N_2563,N_2601);
nand U2671 (N_2671,N_2622,N_2512);
nor U2672 (N_2672,N_2588,N_2595);
or U2673 (N_2673,N_2602,N_2534);
or U2674 (N_2674,N_2617,N_2624);
or U2675 (N_2675,N_2564,N_2547);
nor U2676 (N_2676,N_2603,N_2535);
or U2677 (N_2677,N_2584,N_2552);
nand U2678 (N_2678,N_2604,N_2505);
or U2679 (N_2679,N_2571,N_2607);
nand U2680 (N_2680,N_2578,N_2606);
nor U2681 (N_2681,N_2524,N_2592);
nand U2682 (N_2682,N_2549,N_2570);
or U2683 (N_2683,N_2615,N_2621);
nor U2684 (N_2684,N_2568,N_2545);
nor U2685 (N_2685,N_2610,N_2542);
xnor U2686 (N_2686,N_2614,N_2594);
nand U2687 (N_2687,N_2573,N_2518);
or U2688 (N_2688,N_2584,N_2588);
and U2689 (N_2689,N_2524,N_2610);
or U2690 (N_2690,N_2578,N_2556);
nor U2691 (N_2691,N_2525,N_2596);
xnor U2692 (N_2692,N_2509,N_2577);
nor U2693 (N_2693,N_2530,N_2537);
nor U2694 (N_2694,N_2528,N_2579);
nand U2695 (N_2695,N_2616,N_2591);
nor U2696 (N_2696,N_2588,N_2580);
or U2697 (N_2697,N_2555,N_2562);
or U2698 (N_2698,N_2537,N_2572);
or U2699 (N_2699,N_2590,N_2543);
or U2700 (N_2700,N_2561,N_2591);
nor U2701 (N_2701,N_2600,N_2508);
xnor U2702 (N_2702,N_2604,N_2615);
and U2703 (N_2703,N_2500,N_2613);
or U2704 (N_2704,N_2555,N_2572);
or U2705 (N_2705,N_2603,N_2541);
or U2706 (N_2706,N_2579,N_2598);
xor U2707 (N_2707,N_2622,N_2563);
or U2708 (N_2708,N_2553,N_2543);
or U2709 (N_2709,N_2531,N_2582);
xor U2710 (N_2710,N_2514,N_2583);
and U2711 (N_2711,N_2551,N_2570);
xor U2712 (N_2712,N_2505,N_2517);
and U2713 (N_2713,N_2618,N_2600);
nand U2714 (N_2714,N_2533,N_2618);
or U2715 (N_2715,N_2588,N_2527);
and U2716 (N_2716,N_2540,N_2591);
nor U2717 (N_2717,N_2610,N_2536);
nand U2718 (N_2718,N_2518,N_2507);
or U2719 (N_2719,N_2607,N_2560);
nand U2720 (N_2720,N_2568,N_2607);
or U2721 (N_2721,N_2521,N_2603);
or U2722 (N_2722,N_2594,N_2572);
or U2723 (N_2723,N_2501,N_2533);
and U2724 (N_2724,N_2598,N_2568);
nand U2725 (N_2725,N_2611,N_2545);
nor U2726 (N_2726,N_2589,N_2515);
xnor U2727 (N_2727,N_2581,N_2500);
and U2728 (N_2728,N_2531,N_2617);
xor U2729 (N_2729,N_2616,N_2542);
or U2730 (N_2730,N_2602,N_2595);
nand U2731 (N_2731,N_2555,N_2545);
or U2732 (N_2732,N_2540,N_2563);
xnor U2733 (N_2733,N_2604,N_2551);
or U2734 (N_2734,N_2537,N_2598);
nand U2735 (N_2735,N_2612,N_2511);
and U2736 (N_2736,N_2574,N_2621);
xor U2737 (N_2737,N_2573,N_2550);
xor U2738 (N_2738,N_2573,N_2540);
nand U2739 (N_2739,N_2506,N_2595);
nor U2740 (N_2740,N_2527,N_2500);
nor U2741 (N_2741,N_2508,N_2598);
nor U2742 (N_2742,N_2545,N_2548);
nor U2743 (N_2743,N_2569,N_2604);
and U2744 (N_2744,N_2576,N_2620);
or U2745 (N_2745,N_2576,N_2565);
and U2746 (N_2746,N_2592,N_2527);
and U2747 (N_2747,N_2509,N_2594);
nand U2748 (N_2748,N_2586,N_2525);
or U2749 (N_2749,N_2617,N_2605);
and U2750 (N_2750,N_2739,N_2734);
xnor U2751 (N_2751,N_2680,N_2670);
and U2752 (N_2752,N_2682,N_2650);
xnor U2753 (N_2753,N_2669,N_2672);
nor U2754 (N_2754,N_2746,N_2658);
and U2755 (N_2755,N_2738,N_2706);
nand U2756 (N_2756,N_2626,N_2635);
nor U2757 (N_2757,N_2664,N_2722);
xor U2758 (N_2758,N_2728,N_2665);
xnor U2759 (N_2759,N_2634,N_2683);
xnor U2760 (N_2760,N_2639,N_2716);
and U2761 (N_2761,N_2733,N_2656);
nor U2762 (N_2762,N_2667,N_2748);
and U2763 (N_2763,N_2740,N_2659);
xor U2764 (N_2764,N_2645,N_2673);
xnor U2765 (N_2765,N_2663,N_2653);
and U2766 (N_2766,N_2689,N_2652);
and U2767 (N_2767,N_2657,N_2671);
nand U2768 (N_2768,N_2717,N_2698);
nand U2769 (N_2769,N_2725,N_2654);
xnor U2770 (N_2770,N_2647,N_2719);
nor U2771 (N_2771,N_2702,N_2629);
xor U2772 (N_2772,N_2735,N_2692);
and U2773 (N_2773,N_2676,N_2732);
nor U2774 (N_2774,N_2684,N_2641);
and U2775 (N_2775,N_2693,N_2749);
or U2776 (N_2776,N_2697,N_2631);
and U2777 (N_2777,N_2660,N_2644);
nor U2778 (N_2778,N_2704,N_2710);
xnor U2779 (N_2779,N_2679,N_2736);
xnor U2780 (N_2780,N_2731,N_2712);
nand U2781 (N_2781,N_2661,N_2638);
nor U2782 (N_2782,N_2723,N_2701);
nor U2783 (N_2783,N_2708,N_2691);
nand U2784 (N_2784,N_2628,N_2687);
xnor U2785 (N_2785,N_2727,N_2632);
and U2786 (N_2786,N_2709,N_2705);
and U2787 (N_2787,N_2713,N_2651);
nand U2788 (N_2788,N_2630,N_2718);
or U2789 (N_2789,N_2677,N_2668);
nand U2790 (N_2790,N_2686,N_2690);
or U2791 (N_2791,N_2649,N_2637);
nor U2792 (N_2792,N_2685,N_2674);
and U2793 (N_2793,N_2627,N_2694);
nor U2794 (N_2794,N_2688,N_2741);
nor U2795 (N_2795,N_2675,N_2703);
nor U2796 (N_2796,N_2666,N_2695);
or U2797 (N_2797,N_2715,N_2730);
and U2798 (N_2798,N_2729,N_2745);
or U2799 (N_2799,N_2724,N_2699);
nand U2800 (N_2800,N_2707,N_2742);
nor U2801 (N_2801,N_2700,N_2696);
nand U2802 (N_2802,N_2636,N_2640);
or U2803 (N_2803,N_2737,N_2662);
nand U2804 (N_2804,N_2743,N_2648);
xor U2805 (N_2805,N_2646,N_2714);
xor U2806 (N_2806,N_2678,N_2747);
and U2807 (N_2807,N_2655,N_2726);
nand U2808 (N_2808,N_2744,N_2720);
nand U2809 (N_2809,N_2642,N_2721);
nor U2810 (N_2810,N_2633,N_2625);
nor U2811 (N_2811,N_2681,N_2711);
or U2812 (N_2812,N_2643,N_2662);
xor U2813 (N_2813,N_2717,N_2687);
and U2814 (N_2814,N_2741,N_2642);
or U2815 (N_2815,N_2712,N_2683);
nor U2816 (N_2816,N_2634,N_2670);
nand U2817 (N_2817,N_2654,N_2719);
and U2818 (N_2818,N_2685,N_2714);
or U2819 (N_2819,N_2637,N_2631);
nand U2820 (N_2820,N_2715,N_2625);
and U2821 (N_2821,N_2679,N_2645);
nor U2822 (N_2822,N_2732,N_2718);
nand U2823 (N_2823,N_2690,N_2626);
and U2824 (N_2824,N_2656,N_2744);
and U2825 (N_2825,N_2636,N_2664);
or U2826 (N_2826,N_2685,N_2692);
xnor U2827 (N_2827,N_2733,N_2731);
nor U2828 (N_2828,N_2665,N_2694);
or U2829 (N_2829,N_2703,N_2700);
nor U2830 (N_2830,N_2713,N_2694);
nor U2831 (N_2831,N_2679,N_2709);
nor U2832 (N_2832,N_2739,N_2635);
or U2833 (N_2833,N_2647,N_2676);
nand U2834 (N_2834,N_2644,N_2747);
or U2835 (N_2835,N_2705,N_2731);
nand U2836 (N_2836,N_2749,N_2739);
and U2837 (N_2837,N_2711,N_2713);
or U2838 (N_2838,N_2700,N_2716);
and U2839 (N_2839,N_2654,N_2689);
nand U2840 (N_2840,N_2727,N_2685);
nor U2841 (N_2841,N_2727,N_2736);
nor U2842 (N_2842,N_2700,N_2733);
and U2843 (N_2843,N_2672,N_2677);
xnor U2844 (N_2844,N_2713,N_2659);
xnor U2845 (N_2845,N_2746,N_2742);
nand U2846 (N_2846,N_2748,N_2683);
xor U2847 (N_2847,N_2679,N_2716);
or U2848 (N_2848,N_2651,N_2645);
nor U2849 (N_2849,N_2730,N_2635);
or U2850 (N_2850,N_2690,N_2631);
nor U2851 (N_2851,N_2744,N_2666);
or U2852 (N_2852,N_2652,N_2672);
nor U2853 (N_2853,N_2662,N_2647);
xnor U2854 (N_2854,N_2680,N_2697);
or U2855 (N_2855,N_2681,N_2697);
and U2856 (N_2856,N_2721,N_2668);
and U2857 (N_2857,N_2684,N_2714);
and U2858 (N_2858,N_2684,N_2626);
nand U2859 (N_2859,N_2696,N_2678);
xnor U2860 (N_2860,N_2646,N_2734);
and U2861 (N_2861,N_2681,N_2649);
nand U2862 (N_2862,N_2685,N_2638);
nand U2863 (N_2863,N_2641,N_2712);
nor U2864 (N_2864,N_2745,N_2643);
nor U2865 (N_2865,N_2641,N_2643);
nand U2866 (N_2866,N_2740,N_2632);
xnor U2867 (N_2867,N_2715,N_2720);
nand U2868 (N_2868,N_2663,N_2651);
or U2869 (N_2869,N_2674,N_2702);
and U2870 (N_2870,N_2706,N_2717);
nor U2871 (N_2871,N_2638,N_2738);
xnor U2872 (N_2872,N_2655,N_2711);
xnor U2873 (N_2873,N_2629,N_2706);
nand U2874 (N_2874,N_2660,N_2695);
xnor U2875 (N_2875,N_2778,N_2867);
nand U2876 (N_2876,N_2837,N_2854);
or U2877 (N_2877,N_2865,N_2850);
nor U2878 (N_2878,N_2871,N_2784);
or U2879 (N_2879,N_2800,N_2752);
nor U2880 (N_2880,N_2814,N_2805);
nor U2881 (N_2881,N_2763,N_2821);
and U2882 (N_2882,N_2864,N_2755);
and U2883 (N_2883,N_2874,N_2790);
xor U2884 (N_2884,N_2858,N_2832);
and U2885 (N_2885,N_2789,N_2857);
nand U2886 (N_2886,N_2840,N_2827);
or U2887 (N_2887,N_2863,N_2833);
or U2888 (N_2888,N_2802,N_2862);
nand U2889 (N_2889,N_2776,N_2797);
or U2890 (N_2890,N_2785,N_2868);
or U2891 (N_2891,N_2774,N_2824);
nand U2892 (N_2892,N_2777,N_2753);
xor U2893 (N_2893,N_2804,N_2793);
nand U2894 (N_2894,N_2751,N_2765);
nor U2895 (N_2895,N_2846,N_2869);
nor U2896 (N_2896,N_2801,N_2835);
or U2897 (N_2897,N_2870,N_2781);
xnor U2898 (N_2898,N_2808,N_2799);
xor U2899 (N_2899,N_2807,N_2779);
nor U2900 (N_2900,N_2754,N_2841);
xnor U2901 (N_2901,N_2770,N_2794);
xor U2902 (N_2902,N_2828,N_2768);
xor U2903 (N_2903,N_2775,N_2758);
nand U2904 (N_2904,N_2829,N_2787);
nor U2905 (N_2905,N_2847,N_2825);
nor U2906 (N_2906,N_2815,N_2816);
nand U2907 (N_2907,N_2836,N_2798);
nor U2908 (N_2908,N_2826,N_2773);
and U2909 (N_2909,N_2757,N_2855);
or U2910 (N_2910,N_2852,N_2760);
and U2911 (N_2911,N_2750,N_2759);
and U2912 (N_2912,N_2803,N_2792);
nor U2913 (N_2913,N_2783,N_2812);
nor U2914 (N_2914,N_2849,N_2842);
xnor U2915 (N_2915,N_2856,N_2845);
nor U2916 (N_2916,N_2796,N_2819);
nor U2917 (N_2917,N_2782,N_2830);
xnor U2918 (N_2918,N_2853,N_2761);
xnor U2919 (N_2919,N_2795,N_2786);
nand U2920 (N_2920,N_2851,N_2844);
nand U2921 (N_2921,N_2766,N_2838);
and U2922 (N_2922,N_2771,N_2823);
nand U2923 (N_2923,N_2813,N_2860);
and U2924 (N_2924,N_2762,N_2756);
or U2925 (N_2925,N_2767,N_2769);
and U2926 (N_2926,N_2859,N_2839);
xor U2927 (N_2927,N_2810,N_2843);
nor U2928 (N_2928,N_2806,N_2872);
xnor U2929 (N_2929,N_2834,N_2791);
nand U2930 (N_2930,N_2788,N_2848);
nor U2931 (N_2931,N_2811,N_2861);
or U2932 (N_2932,N_2772,N_2831);
and U2933 (N_2933,N_2820,N_2822);
and U2934 (N_2934,N_2809,N_2764);
xnor U2935 (N_2935,N_2818,N_2780);
or U2936 (N_2936,N_2866,N_2817);
nand U2937 (N_2937,N_2873,N_2793);
nor U2938 (N_2938,N_2810,N_2799);
or U2939 (N_2939,N_2768,N_2809);
or U2940 (N_2940,N_2842,N_2851);
nor U2941 (N_2941,N_2828,N_2831);
or U2942 (N_2942,N_2807,N_2783);
xor U2943 (N_2943,N_2782,N_2792);
nor U2944 (N_2944,N_2827,N_2848);
nand U2945 (N_2945,N_2823,N_2829);
or U2946 (N_2946,N_2862,N_2815);
nand U2947 (N_2947,N_2818,N_2760);
nand U2948 (N_2948,N_2760,N_2841);
xor U2949 (N_2949,N_2871,N_2840);
or U2950 (N_2950,N_2810,N_2873);
and U2951 (N_2951,N_2861,N_2789);
nand U2952 (N_2952,N_2831,N_2783);
nor U2953 (N_2953,N_2856,N_2769);
or U2954 (N_2954,N_2783,N_2809);
nand U2955 (N_2955,N_2823,N_2865);
and U2956 (N_2956,N_2827,N_2856);
or U2957 (N_2957,N_2777,N_2854);
or U2958 (N_2958,N_2796,N_2770);
xnor U2959 (N_2959,N_2811,N_2808);
and U2960 (N_2960,N_2870,N_2807);
nor U2961 (N_2961,N_2765,N_2787);
nand U2962 (N_2962,N_2796,N_2797);
or U2963 (N_2963,N_2858,N_2853);
nand U2964 (N_2964,N_2761,N_2787);
xnor U2965 (N_2965,N_2784,N_2830);
nor U2966 (N_2966,N_2766,N_2780);
and U2967 (N_2967,N_2872,N_2858);
xnor U2968 (N_2968,N_2812,N_2782);
nor U2969 (N_2969,N_2873,N_2843);
xor U2970 (N_2970,N_2792,N_2790);
nor U2971 (N_2971,N_2828,N_2754);
xnor U2972 (N_2972,N_2848,N_2807);
nor U2973 (N_2973,N_2781,N_2832);
or U2974 (N_2974,N_2831,N_2804);
nor U2975 (N_2975,N_2788,N_2839);
and U2976 (N_2976,N_2754,N_2839);
nor U2977 (N_2977,N_2870,N_2788);
xnor U2978 (N_2978,N_2835,N_2789);
nand U2979 (N_2979,N_2804,N_2863);
nor U2980 (N_2980,N_2787,N_2752);
nand U2981 (N_2981,N_2846,N_2791);
and U2982 (N_2982,N_2787,N_2868);
nor U2983 (N_2983,N_2753,N_2772);
and U2984 (N_2984,N_2857,N_2759);
nand U2985 (N_2985,N_2827,N_2754);
nand U2986 (N_2986,N_2805,N_2861);
nand U2987 (N_2987,N_2854,N_2764);
and U2988 (N_2988,N_2790,N_2856);
xor U2989 (N_2989,N_2856,N_2779);
xor U2990 (N_2990,N_2773,N_2865);
or U2991 (N_2991,N_2783,N_2821);
nor U2992 (N_2992,N_2847,N_2753);
nor U2993 (N_2993,N_2859,N_2790);
xor U2994 (N_2994,N_2862,N_2762);
or U2995 (N_2995,N_2839,N_2829);
and U2996 (N_2996,N_2846,N_2810);
nor U2997 (N_2997,N_2868,N_2756);
xnor U2998 (N_2998,N_2778,N_2855);
nand U2999 (N_2999,N_2840,N_2869);
nor U3000 (N_3000,N_2949,N_2913);
xor U3001 (N_3001,N_2991,N_2989);
or U3002 (N_3002,N_2922,N_2979);
and U3003 (N_3003,N_2980,N_2881);
xor U3004 (N_3004,N_2898,N_2876);
nand U3005 (N_3005,N_2953,N_2901);
or U3006 (N_3006,N_2905,N_2887);
or U3007 (N_3007,N_2946,N_2950);
nand U3008 (N_3008,N_2877,N_2959);
nand U3009 (N_3009,N_2954,N_2948);
nand U3010 (N_3010,N_2994,N_2977);
and U3011 (N_3011,N_2878,N_2970);
xor U3012 (N_3012,N_2918,N_2884);
nor U3013 (N_3013,N_2961,N_2938);
xnor U3014 (N_3014,N_2908,N_2943);
xor U3015 (N_3015,N_2909,N_2886);
and U3016 (N_3016,N_2955,N_2920);
and U3017 (N_3017,N_2911,N_2974);
nor U3018 (N_3018,N_2995,N_2937);
nor U3019 (N_3019,N_2917,N_2968);
or U3020 (N_3020,N_2891,N_2965);
or U3021 (N_3021,N_2964,N_2983);
xor U3022 (N_3022,N_2996,N_2892);
and U3023 (N_3023,N_2986,N_2935);
xor U3024 (N_3024,N_2929,N_2889);
nor U3025 (N_3025,N_2925,N_2879);
and U3026 (N_3026,N_2988,N_2899);
and U3027 (N_3027,N_2941,N_2947);
nor U3028 (N_3028,N_2933,N_2999);
nand U3029 (N_3029,N_2900,N_2934);
or U3030 (N_3030,N_2975,N_2930);
nor U3031 (N_3031,N_2967,N_2992);
and U3032 (N_3032,N_2984,N_2942);
xnor U3033 (N_3033,N_2915,N_2897);
nand U3034 (N_3034,N_2924,N_2904);
xor U3035 (N_3035,N_2957,N_2890);
and U3036 (N_3036,N_2921,N_2875);
nor U3037 (N_3037,N_2973,N_2952);
and U3038 (N_3038,N_2914,N_2981);
nor U3039 (N_3039,N_2976,N_2888);
and U3040 (N_3040,N_2993,N_2907);
xnor U3041 (N_3041,N_2960,N_2894);
nand U3042 (N_3042,N_2883,N_2896);
nand U3043 (N_3043,N_2882,N_2963);
nor U3044 (N_3044,N_2945,N_2962);
and U3045 (N_3045,N_2969,N_2971);
and U3046 (N_3046,N_2940,N_2939);
xnor U3047 (N_3047,N_2987,N_2951);
nand U3048 (N_3048,N_2927,N_2990);
or U3049 (N_3049,N_2936,N_2958);
xor U3050 (N_3050,N_2885,N_2923);
and U3051 (N_3051,N_2985,N_2944);
nor U3052 (N_3052,N_2893,N_2978);
and U3053 (N_3053,N_2902,N_2926);
xnor U3054 (N_3054,N_2910,N_2895);
nor U3055 (N_3055,N_2931,N_2912);
nand U3056 (N_3056,N_2916,N_2906);
and U3057 (N_3057,N_2956,N_2982);
nand U3058 (N_3058,N_2998,N_2903);
or U3059 (N_3059,N_2932,N_2972);
or U3060 (N_3060,N_2997,N_2928);
xnor U3061 (N_3061,N_2966,N_2880);
or U3062 (N_3062,N_2919,N_2910);
or U3063 (N_3063,N_2891,N_2996);
and U3064 (N_3064,N_2937,N_2917);
nor U3065 (N_3065,N_2878,N_2947);
xnor U3066 (N_3066,N_2898,N_2991);
or U3067 (N_3067,N_2939,N_2963);
nand U3068 (N_3068,N_2978,N_2920);
or U3069 (N_3069,N_2985,N_2891);
and U3070 (N_3070,N_2926,N_2977);
nor U3071 (N_3071,N_2992,N_2882);
nand U3072 (N_3072,N_2940,N_2912);
or U3073 (N_3073,N_2880,N_2889);
nor U3074 (N_3074,N_2957,N_2939);
xor U3075 (N_3075,N_2955,N_2954);
xnor U3076 (N_3076,N_2901,N_2920);
or U3077 (N_3077,N_2981,N_2937);
nand U3078 (N_3078,N_2951,N_2978);
or U3079 (N_3079,N_2887,N_2889);
xnor U3080 (N_3080,N_2949,N_2966);
or U3081 (N_3081,N_2934,N_2925);
or U3082 (N_3082,N_2937,N_2906);
nor U3083 (N_3083,N_2959,N_2933);
xnor U3084 (N_3084,N_2891,N_2981);
and U3085 (N_3085,N_2931,N_2929);
xor U3086 (N_3086,N_2924,N_2960);
nor U3087 (N_3087,N_2972,N_2965);
xnor U3088 (N_3088,N_2905,N_2968);
nor U3089 (N_3089,N_2941,N_2969);
xnor U3090 (N_3090,N_2925,N_2917);
nor U3091 (N_3091,N_2913,N_2891);
or U3092 (N_3092,N_2951,N_2982);
and U3093 (N_3093,N_2987,N_2971);
and U3094 (N_3094,N_2948,N_2931);
or U3095 (N_3095,N_2940,N_2992);
nand U3096 (N_3096,N_2954,N_2903);
nand U3097 (N_3097,N_2990,N_2935);
and U3098 (N_3098,N_2968,N_2952);
nand U3099 (N_3099,N_2875,N_2977);
nor U3100 (N_3100,N_2992,N_2994);
nand U3101 (N_3101,N_2946,N_2905);
xnor U3102 (N_3102,N_2975,N_2990);
nor U3103 (N_3103,N_2913,N_2885);
nor U3104 (N_3104,N_2927,N_2905);
and U3105 (N_3105,N_2949,N_2947);
nor U3106 (N_3106,N_2988,N_2951);
nand U3107 (N_3107,N_2913,N_2934);
or U3108 (N_3108,N_2887,N_2882);
or U3109 (N_3109,N_2952,N_2950);
nand U3110 (N_3110,N_2895,N_2936);
nand U3111 (N_3111,N_2931,N_2886);
nor U3112 (N_3112,N_2943,N_2974);
nor U3113 (N_3113,N_2880,N_2877);
nor U3114 (N_3114,N_2960,N_2940);
nor U3115 (N_3115,N_2927,N_2955);
or U3116 (N_3116,N_2892,N_2898);
xor U3117 (N_3117,N_2956,N_2889);
nand U3118 (N_3118,N_2892,N_2896);
xnor U3119 (N_3119,N_2957,N_2895);
or U3120 (N_3120,N_2948,N_2955);
or U3121 (N_3121,N_2965,N_2939);
or U3122 (N_3122,N_2994,N_2971);
nand U3123 (N_3123,N_2880,N_2927);
nor U3124 (N_3124,N_2878,N_2902);
or U3125 (N_3125,N_3051,N_3040);
or U3126 (N_3126,N_3033,N_3061);
nand U3127 (N_3127,N_3060,N_3002);
nor U3128 (N_3128,N_3119,N_3088);
xnor U3129 (N_3129,N_3115,N_3053);
or U3130 (N_3130,N_3123,N_3111);
nor U3131 (N_3131,N_3103,N_3031);
nor U3132 (N_3132,N_3102,N_3015);
nand U3133 (N_3133,N_3078,N_3058);
and U3134 (N_3134,N_3034,N_3025);
or U3135 (N_3135,N_3022,N_3065);
and U3136 (N_3136,N_3029,N_3049);
nor U3137 (N_3137,N_3037,N_3018);
and U3138 (N_3138,N_3059,N_3045);
or U3139 (N_3139,N_3003,N_3116);
or U3140 (N_3140,N_3090,N_3094);
and U3141 (N_3141,N_3124,N_3004);
or U3142 (N_3142,N_3001,N_3036);
and U3143 (N_3143,N_3047,N_3109);
or U3144 (N_3144,N_3106,N_3057);
nor U3145 (N_3145,N_3016,N_3030);
nand U3146 (N_3146,N_3010,N_3120);
nor U3147 (N_3147,N_3114,N_3066);
xnor U3148 (N_3148,N_3099,N_3054);
xor U3149 (N_3149,N_3052,N_3100);
and U3150 (N_3150,N_3113,N_3009);
and U3151 (N_3151,N_3062,N_3077);
or U3152 (N_3152,N_3073,N_3085);
nor U3153 (N_3153,N_3023,N_3007);
or U3154 (N_3154,N_3043,N_3011);
nand U3155 (N_3155,N_3112,N_3008);
nand U3156 (N_3156,N_3035,N_3110);
nand U3157 (N_3157,N_3063,N_3091);
nor U3158 (N_3158,N_3044,N_3075);
and U3159 (N_3159,N_3050,N_3074);
and U3160 (N_3160,N_3081,N_3076);
nand U3161 (N_3161,N_3028,N_3024);
and U3162 (N_3162,N_3042,N_3064);
nand U3163 (N_3163,N_3006,N_3095);
nor U3164 (N_3164,N_3122,N_3032);
xnor U3165 (N_3165,N_3039,N_3084);
xor U3166 (N_3166,N_3072,N_3020);
and U3167 (N_3167,N_3097,N_3019);
or U3168 (N_3168,N_3000,N_3087);
and U3169 (N_3169,N_3079,N_3041);
and U3170 (N_3170,N_3098,N_3012);
xnor U3171 (N_3171,N_3082,N_3101);
xor U3172 (N_3172,N_3093,N_3080);
or U3173 (N_3173,N_3056,N_3048);
nand U3174 (N_3174,N_3021,N_3117);
or U3175 (N_3175,N_3089,N_3104);
nand U3176 (N_3176,N_3046,N_3055);
nand U3177 (N_3177,N_3038,N_3107);
and U3178 (N_3178,N_3096,N_3005);
xor U3179 (N_3179,N_3070,N_3121);
xor U3180 (N_3180,N_3027,N_3069);
xor U3181 (N_3181,N_3108,N_3092);
nand U3182 (N_3182,N_3071,N_3017);
xor U3183 (N_3183,N_3083,N_3014);
xor U3184 (N_3184,N_3105,N_3068);
nor U3185 (N_3185,N_3013,N_3086);
nor U3186 (N_3186,N_3118,N_3026);
xnor U3187 (N_3187,N_3067,N_3017);
nand U3188 (N_3188,N_3065,N_3093);
or U3189 (N_3189,N_3089,N_3006);
nand U3190 (N_3190,N_3016,N_3093);
nor U3191 (N_3191,N_3020,N_3083);
xor U3192 (N_3192,N_3055,N_3097);
xnor U3193 (N_3193,N_3079,N_3043);
nor U3194 (N_3194,N_3091,N_3011);
xnor U3195 (N_3195,N_3071,N_3051);
or U3196 (N_3196,N_3011,N_3120);
nor U3197 (N_3197,N_3122,N_3036);
nor U3198 (N_3198,N_3085,N_3005);
nor U3199 (N_3199,N_3009,N_3095);
and U3200 (N_3200,N_3104,N_3054);
nand U3201 (N_3201,N_3006,N_3016);
nor U3202 (N_3202,N_3042,N_3117);
nor U3203 (N_3203,N_3111,N_3087);
nand U3204 (N_3204,N_3036,N_3047);
nor U3205 (N_3205,N_3077,N_3043);
xor U3206 (N_3206,N_3100,N_3055);
nor U3207 (N_3207,N_3096,N_3084);
and U3208 (N_3208,N_3122,N_3004);
xor U3209 (N_3209,N_3078,N_3092);
nand U3210 (N_3210,N_3027,N_3055);
xor U3211 (N_3211,N_3050,N_3006);
and U3212 (N_3212,N_3106,N_3090);
nor U3213 (N_3213,N_3048,N_3005);
xor U3214 (N_3214,N_3092,N_3002);
xor U3215 (N_3215,N_3073,N_3010);
nor U3216 (N_3216,N_3072,N_3094);
nor U3217 (N_3217,N_3043,N_3105);
xor U3218 (N_3218,N_3008,N_3006);
or U3219 (N_3219,N_3109,N_3124);
and U3220 (N_3220,N_3002,N_3056);
nor U3221 (N_3221,N_3070,N_3001);
nor U3222 (N_3222,N_3051,N_3070);
or U3223 (N_3223,N_3113,N_3022);
xnor U3224 (N_3224,N_3072,N_3040);
nand U3225 (N_3225,N_3109,N_3046);
or U3226 (N_3226,N_3003,N_3042);
and U3227 (N_3227,N_3122,N_3041);
xor U3228 (N_3228,N_3102,N_3096);
nand U3229 (N_3229,N_3004,N_3113);
and U3230 (N_3230,N_3015,N_3020);
nor U3231 (N_3231,N_3016,N_3045);
nand U3232 (N_3232,N_3004,N_3086);
and U3233 (N_3233,N_3052,N_3059);
nand U3234 (N_3234,N_3107,N_3016);
or U3235 (N_3235,N_3015,N_3008);
nor U3236 (N_3236,N_3068,N_3040);
or U3237 (N_3237,N_3000,N_3041);
xor U3238 (N_3238,N_3063,N_3055);
nor U3239 (N_3239,N_3118,N_3022);
nor U3240 (N_3240,N_3112,N_3082);
or U3241 (N_3241,N_3011,N_3073);
xnor U3242 (N_3242,N_3012,N_3096);
xor U3243 (N_3243,N_3061,N_3048);
or U3244 (N_3244,N_3042,N_3018);
or U3245 (N_3245,N_3107,N_3041);
nand U3246 (N_3246,N_3040,N_3108);
xor U3247 (N_3247,N_3003,N_3010);
and U3248 (N_3248,N_3035,N_3001);
nor U3249 (N_3249,N_3072,N_3090);
nand U3250 (N_3250,N_3212,N_3131);
nor U3251 (N_3251,N_3184,N_3125);
xnor U3252 (N_3252,N_3137,N_3230);
nor U3253 (N_3253,N_3240,N_3185);
xnor U3254 (N_3254,N_3203,N_3168);
xor U3255 (N_3255,N_3175,N_3195);
xor U3256 (N_3256,N_3206,N_3219);
xor U3257 (N_3257,N_3221,N_3157);
or U3258 (N_3258,N_3208,N_3214);
nand U3259 (N_3259,N_3162,N_3244);
and U3260 (N_3260,N_3245,N_3128);
or U3261 (N_3261,N_3170,N_3187);
or U3262 (N_3262,N_3163,N_3236);
nand U3263 (N_3263,N_3165,N_3153);
or U3264 (N_3264,N_3151,N_3243);
xnor U3265 (N_3265,N_3136,N_3217);
or U3266 (N_3266,N_3127,N_3130);
or U3267 (N_3267,N_3179,N_3158);
nand U3268 (N_3268,N_3164,N_3148);
xnor U3269 (N_3269,N_3229,N_3237);
xor U3270 (N_3270,N_3149,N_3210);
or U3271 (N_3271,N_3202,N_3235);
nand U3272 (N_3272,N_3216,N_3138);
xor U3273 (N_3273,N_3232,N_3227);
nor U3274 (N_3274,N_3211,N_3248);
nand U3275 (N_3275,N_3132,N_3241);
nor U3276 (N_3276,N_3172,N_3146);
or U3277 (N_3277,N_3171,N_3173);
and U3278 (N_3278,N_3166,N_3133);
or U3279 (N_3279,N_3198,N_3197);
and U3280 (N_3280,N_3182,N_3142);
and U3281 (N_3281,N_3196,N_3190);
or U3282 (N_3282,N_3220,N_3177);
or U3283 (N_3283,N_3186,N_3193);
nor U3284 (N_3284,N_3150,N_3189);
or U3285 (N_3285,N_3215,N_3204);
or U3286 (N_3286,N_3143,N_3200);
or U3287 (N_3287,N_3218,N_3228);
nand U3288 (N_3288,N_3134,N_3161);
nand U3289 (N_3289,N_3222,N_3154);
nor U3290 (N_3290,N_3139,N_3191);
nor U3291 (N_3291,N_3238,N_3145);
nor U3292 (N_3292,N_3226,N_3224);
or U3293 (N_3293,N_3159,N_3156);
and U3294 (N_3294,N_3180,N_3144);
nand U3295 (N_3295,N_3141,N_3234);
nand U3296 (N_3296,N_3205,N_3176);
and U3297 (N_3297,N_3167,N_3242);
nand U3298 (N_3298,N_3199,N_3152);
and U3299 (N_3299,N_3246,N_3178);
nand U3300 (N_3300,N_3181,N_3140);
or U3301 (N_3301,N_3249,N_3155);
and U3302 (N_3302,N_3126,N_3183);
nand U3303 (N_3303,N_3169,N_3223);
nand U3304 (N_3304,N_3174,N_3135);
and U3305 (N_3305,N_3194,N_3213);
xor U3306 (N_3306,N_3129,N_3201);
nand U3307 (N_3307,N_3160,N_3247);
nand U3308 (N_3308,N_3239,N_3188);
xnor U3309 (N_3309,N_3192,N_3225);
xor U3310 (N_3310,N_3233,N_3207);
xor U3311 (N_3311,N_3209,N_3231);
xor U3312 (N_3312,N_3147,N_3212);
xnor U3313 (N_3313,N_3246,N_3190);
or U3314 (N_3314,N_3212,N_3132);
xnor U3315 (N_3315,N_3219,N_3152);
and U3316 (N_3316,N_3167,N_3214);
or U3317 (N_3317,N_3246,N_3141);
and U3318 (N_3318,N_3166,N_3145);
xor U3319 (N_3319,N_3127,N_3147);
xnor U3320 (N_3320,N_3139,N_3146);
xor U3321 (N_3321,N_3207,N_3161);
or U3322 (N_3322,N_3136,N_3222);
or U3323 (N_3323,N_3231,N_3232);
xor U3324 (N_3324,N_3148,N_3191);
and U3325 (N_3325,N_3142,N_3171);
or U3326 (N_3326,N_3153,N_3139);
and U3327 (N_3327,N_3234,N_3203);
or U3328 (N_3328,N_3134,N_3236);
nor U3329 (N_3329,N_3185,N_3225);
or U3330 (N_3330,N_3204,N_3221);
xnor U3331 (N_3331,N_3199,N_3216);
or U3332 (N_3332,N_3128,N_3176);
nor U3333 (N_3333,N_3187,N_3245);
nor U3334 (N_3334,N_3208,N_3246);
xor U3335 (N_3335,N_3162,N_3125);
nor U3336 (N_3336,N_3218,N_3247);
nor U3337 (N_3337,N_3187,N_3175);
nand U3338 (N_3338,N_3178,N_3150);
or U3339 (N_3339,N_3125,N_3221);
and U3340 (N_3340,N_3155,N_3212);
nor U3341 (N_3341,N_3147,N_3200);
or U3342 (N_3342,N_3130,N_3150);
and U3343 (N_3343,N_3148,N_3144);
nor U3344 (N_3344,N_3182,N_3162);
nand U3345 (N_3345,N_3249,N_3241);
nand U3346 (N_3346,N_3136,N_3205);
or U3347 (N_3347,N_3211,N_3223);
xor U3348 (N_3348,N_3159,N_3220);
xnor U3349 (N_3349,N_3211,N_3158);
nand U3350 (N_3350,N_3141,N_3137);
or U3351 (N_3351,N_3168,N_3178);
and U3352 (N_3352,N_3181,N_3175);
xor U3353 (N_3353,N_3183,N_3164);
or U3354 (N_3354,N_3155,N_3223);
nand U3355 (N_3355,N_3161,N_3214);
and U3356 (N_3356,N_3183,N_3158);
nor U3357 (N_3357,N_3130,N_3198);
xnor U3358 (N_3358,N_3225,N_3155);
and U3359 (N_3359,N_3248,N_3249);
nand U3360 (N_3360,N_3237,N_3151);
nor U3361 (N_3361,N_3235,N_3219);
and U3362 (N_3362,N_3237,N_3181);
xnor U3363 (N_3363,N_3233,N_3247);
nand U3364 (N_3364,N_3196,N_3240);
and U3365 (N_3365,N_3188,N_3194);
and U3366 (N_3366,N_3171,N_3216);
or U3367 (N_3367,N_3182,N_3159);
or U3368 (N_3368,N_3187,N_3130);
nand U3369 (N_3369,N_3241,N_3233);
xnor U3370 (N_3370,N_3202,N_3244);
and U3371 (N_3371,N_3133,N_3128);
nand U3372 (N_3372,N_3146,N_3179);
nor U3373 (N_3373,N_3168,N_3166);
or U3374 (N_3374,N_3144,N_3219);
nand U3375 (N_3375,N_3304,N_3333);
xnor U3376 (N_3376,N_3284,N_3286);
or U3377 (N_3377,N_3255,N_3334);
nor U3378 (N_3378,N_3311,N_3279);
or U3379 (N_3379,N_3320,N_3276);
xor U3380 (N_3380,N_3308,N_3314);
and U3381 (N_3381,N_3263,N_3352);
and U3382 (N_3382,N_3296,N_3372);
xor U3383 (N_3383,N_3362,N_3259);
or U3384 (N_3384,N_3294,N_3319);
nand U3385 (N_3385,N_3312,N_3307);
nor U3386 (N_3386,N_3280,N_3250);
or U3387 (N_3387,N_3287,N_3295);
or U3388 (N_3388,N_3373,N_3316);
xor U3389 (N_3389,N_3355,N_3274);
nor U3390 (N_3390,N_3335,N_3283);
nor U3391 (N_3391,N_3328,N_3253);
nand U3392 (N_3392,N_3285,N_3305);
nand U3393 (N_3393,N_3289,N_3336);
nor U3394 (N_3394,N_3266,N_3360);
or U3395 (N_3395,N_3357,N_3254);
nand U3396 (N_3396,N_3356,N_3306);
xnor U3397 (N_3397,N_3337,N_3363);
nand U3398 (N_3398,N_3349,N_3331);
nor U3399 (N_3399,N_3368,N_3277);
and U3400 (N_3400,N_3265,N_3293);
or U3401 (N_3401,N_3270,N_3370);
or U3402 (N_3402,N_3347,N_3325);
xor U3403 (N_3403,N_3339,N_3310);
nor U3404 (N_3404,N_3374,N_3338);
or U3405 (N_3405,N_3344,N_3369);
and U3406 (N_3406,N_3354,N_3343);
nand U3407 (N_3407,N_3299,N_3318);
nand U3408 (N_3408,N_3353,N_3309);
nand U3409 (N_3409,N_3351,N_3261);
nand U3410 (N_3410,N_3340,N_3329);
nor U3411 (N_3411,N_3348,N_3268);
nor U3412 (N_3412,N_3313,N_3345);
nand U3413 (N_3413,N_3346,N_3251);
or U3414 (N_3414,N_3332,N_3361);
or U3415 (N_3415,N_3365,N_3321);
and U3416 (N_3416,N_3282,N_3302);
nand U3417 (N_3417,N_3366,N_3267);
nor U3418 (N_3418,N_3257,N_3297);
nand U3419 (N_3419,N_3350,N_3326);
xnor U3420 (N_3420,N_3291,N_3342);
nand U3421 (N_3421,N_3273,N_3262);
and U3422 (N_3422,N_3264,N_3315);
xnor U3423 (N_3423,N_3290,N_3341);
nand U3424 (N_3424,N_3260,N_3272);
nor U3425 (N_3425,N_3258,N_3256);
xnor U3426 (N_3426,N_3301,N_3322);
nand U3427 (N_3427,N_3292,N_3269);
and U3428 (N_3428,N_3367,N_3359);
or U3429 (N_3429,N_3327,N_3358);
nand U3430 (N_3430,N_3317,N_3281);
nor U3431 (N_3431,N_3371,N_3298);
xnor U3432 (N_3432,N_3271,N_3303);
xnor U3433 (N_3433,N_3275,N_3288);
xor U3434 (N_3434,N_3330,N_3300);
or U3435 (N_3435,N_3278,N_3364);
xor U3436 (N_3436,N_3324,N_3323);
and U3437 (N_3437,N_3252,N_3327);
nor U3438 (N_3438,N_3284,N_3340);
xor U3439 (N_3439,N_3270,N_3316);
and U3440 (N_3440,N_3308,N_3306);
or U3441 (N_3441,N_3355,N_3368);
xor U3442 (N_3442,N_3309,N_3339);
nor U3443 (N_3443,N_3283,N_3342);
and U3444 (N_3444,N_3362,N_3344);
or U3445 (N_3445,N_3289,N_3260);
nor U3446 (N_3446,N_3321,N_3356);
and U3447 (N_3447,N_3275,N_3311);
nand U3448 (N_3448,N_3365,N_3258);
or U3449 (N_3449,N_3305,N_3322);
nand U3450 (N_3450,N_3354,N_3341);
nand U3451 (N_3451,N_3340,N_3300);
and U3452 (N_3452,N_3303,N_3318);
xor U3453 (N_3453,N_3254,N_3260);
xor U3454 (N_3454,N_3374,N_3331);
nand U3455 (N_3455,N_3277,N_3357);
or U3456 (N_3456,N_3361,N_3310);
nor U3457 (N_3457,N_3345,N_3281);
nor U3458 (N_3458,N_3350,N_3309);
or U3459 (N_3459,N_3336,N_3328);
xor U3460 (N_3460,N_3267,N_3335);
nor U3461 (N_3461,N_3269,N_3320);
or U3462 (N_3462,N_3290,N_3308);
nor U3463 (N_3463,N_3308,N_3366);
xnor U3464 (N_3464,N_3269,N_3347);
or U3465 (N_3465,N_3274,N_3335);
nor U3466 (N_3466,N_3290,N_3372);
nand U3467 (N_3467,N_3282,N_3270);
nand U3468 (N_3468,N_3267,N_3341);
and U3469 (N_3469,N_3323,N_3367);
nand U3470 (N_3470,N_3367,N_3291);
xor U3471 (N_3471,N_3281,N_3308);
or U3472 (N_3472,N_3325,N_3358);
xor U3473 (N_3473,N_3258,N_3342);
and U3474 (N_3474,N_3293,N_3304);
xnor U3475 (N_3475,N_3288,N_3305);
or U3476 (N_3476,N_3279,N_3352);
xor U3477 (N_3477,N_3250,N_3266);
nor U3478 (N_3478,N_3291,N_3287);
or U3479 (N_3479,N_3271,N_3321);
and U3480 (N_3480,N_3323,N_3342);
and U3481 (N_3481,N_3360,N_3341);
nand U3482 (N_3482,N_3322,N_3296);
xor U3483 (N_3483,N_3262,N_3346);
nand U3484 (N_3484,N_3321,N_3343);
and U3485 (N_3485,N_3326,N_3254);
or U3486 (N_3486,N_3373,N_3295);
or U3487 (N_3487,N_3272,N_3281);
nor U3488 (N_3488,N_3326,N_3303);
and U3489 (N_3489,N_3372,N_3323);
nor U3490 (N_3490,N_3351,N_3278);
and U3491 (N_3491,N_3266,N_3325);
nor U3492 (N_3492,N_3335,N_3276);
and U3493 (N_3493,N_3292,N_3266);
and U3494 (N_3494,N_3251,N_3324);
nor U3495 (N_3495,N_3251,N_3339);
nand U3496 (N_3496,N_3315,N_3283);
xor U3497 (N_3497,N_3304,N_3325);
and U3498 (N_3498,N_3278,N_3318);
or U3499 (N_3499,N_3316,N_3288);
and U3500 (N_3500,N_3425,N_3429);
nand U3501 (N_3501,N_3460,N_3483);
or U3502 (N_3502,N_3447,N_3481);
xnor U3503 (N_3503,N_3475,N_3385);
nand U3504 (N_3504,N_3487,N_3441);
nand U3505 (N_3505,N_3420,N_3473);
xor U3506 (N_3506,N_3403,N_3484);
nand U3507 (N_3507,N_3470,N_3438);
xnor U3508 (N_3508,N_3471,N_3397);
nor U3509 (N_3509,N_3436,N_3442);
nor U3510 (N_3510,N_3390,N_3409);
nor U3511 (N_3511,N_3392,N_3472);
and U3512 (N_3512,N_3431,N_3380);
xor U3513 (N_3513,N_3389,N_3485);
and U3514 (N_3514,N_3417,N_3494);
nand U3515 (N_3515,N_3378,N_3434);
nor U3516 (N_3516,N_3432,N_3445);
nand U3517 (N_3517,N_3418,N_3427);
nor U3518 (N_3518,N_3444,N_3398);
xor U3519 (N_3519,N_3450,N_3476);
xor U3520 (N_3520,N_3401,N_3486);
xor U3521 (N_3521,N_3413,N_3382);
or U3522 (N_3522,N_3448,N_3394);
nor U3523 (N_3523,N_3455,N_3498);
nand U3524 (N_3524,N_3489,N_3452);
nand U3525 (N_3525,N_3421,N_3446);
nor U3526 (N_3526,N_3400,N_3495);
nor U3527 (N_3527,N_3477,N_3381);
xor U3528 (N_3528,N_3491,N_3488);
and U3529 (N_3529,N_3454,N_3405);
nor U3530 (N_3530,N_3419,N_3404);
xor U3531 (N_3531,N_3459,N_3377);
or U3532 (N_3532,N_3456,N_3435);
xor U3533 (N_3533,N_3383,N_3478);
nor U3534 (N_3534,N_3440,N_3479);
or U3535 (N_3535,N_3393,N_3490);
nor U3536 (N_3536,N_3453,N_3412);
nand U3537 (N_3537,N_3499,N_3424);
nand U3538 (N_3538,N_3462,N_3384);
and U3539 (N_3539,N_3496,N_3449);
xnor U3540 (N_3540,N_3402,N_3411);
nand U3541 (N_3541,N_3388,N_3430);
nand U3542 (N_3542,N_3463,N_3396);
and U3543 (N_3543,N_3387,N_3437);
or U3544 (N_3544,N_3439,N_3410);
xnor U3545 (N_3545,N_3428,N_3433);
xor U3546 (N_3546,N_3466,N_3497);
or U3547 (N_3547,N_3458,N_3416);
nor U3548 (N_3548,N_3407,N_3493);
or U3549 (N_3549,N_3469,N_3391);
nor U3550 (N_3550,N_3492,N_3474);
nand U3551 (N_3551,N_3443,N_3399);
or U3552 (N_3552,N_3414,N_3406);
or U3553 (N_3553,N_3451,N_3482);
xnor U3554 (N_3554,N_3426,N_3395);
nand U3555 (N_3555,N_3480,N_3468);
nand U3556 (N_3556,N_3408,N_3422);
nand U3557 (N_3557,N_3375,N_3465);
nand U3558 (N_3558,N_3461,N_3415);
xor U3559 (N_3559,N_3467,N_3386);
xor U3560 (N_3560,N_3379,N_3423);
and U3561 (N_3561,N_3376,N_3457);
xnor U3562 (N_3562,N_3464,N_3422);
or U3563 (N_3563,N_3378,N_3393);
or U3564 (N_3564,N_3446,N_3490);
nand U3565 (N_3565,N_3493,N_3441);
nand U3566 (N_3566,N_3451,N_3412);
nand U3567 (N_3567,N_3404,N_3417);
and U3568 (N_3568,N_3484,N_3415);
and U3569 (N_3569,N_3409,N_3437);
and U3570 (N_3570,N_3395,N_3441);
and U3571 (N_3571,N_3437,N_3468);
and U3572 (N_3572,N_3443,N_3418);
nand U3573 (N_3573,N_3491,N_3487);
and U3574 (N_3574,N_3489,N_3499);
and U3575 (N_3575,N_3452,N_3486);
nor U3576 (N_3576,N_3493,N_3478);
and U3577 (N_3577,N_3429,N_3376);
or U3578 (N_3578,N_3378,N_3493);
or U3579 (N_3579,N_3420,N_3494);
and U3580 (N_3580,N_3403,N_3448);
or U3581 (N_3581,N_3493,N_3394);
and U3582 (N_3582,N_3448,N_3399);
and U3583 (N_3583,N_3380,N_3466);
and U3584 (N_3584,N_3409,N_3392);
xor U3585 (N_3585,N_3484,N_3472);
nand U3586 (N_3586,N_3486,N_3429);
nor U3587 (N_3587,N_3409,N_3459);
nor U3588 (N_3588,N_3383,N_3432);
xor U3589 (N_3589,N_3461,N_3471);
nand U3590 (N_3590,N_3488,N_3435);
nand U3591 (N_3591,N_3478,N_3414);
or U3592 (N_3592,N_3432,N_3421);
or U3593 (N_3593,N_3465,N_3495);
or U3594 (N_3594,N_3414,N_3391);
and U3595 (N_3595,N_3385,N_3413);
nand U3596 (N_3596,N_3459,N_3463);
or U3597 (N_3597,N_3488,N_3436);
or U3598 (N_3598,N_3452,N_3462);
xnor U3599 (N_3599,N_3463,N_3392);
or U3600 (N_3600,N_3381,N_3383);
nand U3601 (N_3601,N_3489,N_3470);
nor U3602 (N_3602,N_3473,N_3476);
nor U3603 (N_3603,N_3397,N_3378);
or U3604 (N_3604,N_3488,N_3476);
nand U3605 (N_3605,N_3468,N_3395);
xor U3606 (N_3606,N_3425,N_3382);
or U3607 (N_3607,N_3456,N_3465);
and U3608 (N_3608,N_3474,N_3444);
xnor U3609 (N_3609,N_3401,N_3412);
nand U3610 (N_3610,N_3483,N_3444);
or U3611 (N_3611,N_3483,N_3433);
or U3612 (N_3612,N_3422,N_3444);
xnor U3613 (N_3613,N_3400,N_3412);
xor U3614 (N_3614,N_3445,N_3468);
xnor U3615 (N_3615,N_3451,N_3494);
nor U3616 (N_3616,N_3435,N_3463);
nand U3617 (N_3617,N_3462,N_3405);
nand U3618 (N_3618,N_3416,N_3384);
nor U3619 (N_3619,N_3378,N_3375);
and U3620 (N_3620,N_3408,N_3463);
xor U3621 (N_3621,N_3376,N_3430);
nand U3622 (N_3622,N_3470,N_3465);
and U3623 (N_3623,N_3423,N_3428);
or U3624 (N_3624,N_3381,N_3420);
nand U3625 (N_3625,N_3582,N_3556);
nor U3626 (N_3626,N_3511,N_3571);
or U3627 (N_3627,N_3569,N_3595);
or U3628 (N_3628,N_3538,N_3590);
and U3629 (N_3629,N_3617,N_3586);
and U3630 (N_3630,N_3604,N_3605);
nor U3631 (N_3631,N_3516,N_3581);
xor U3632 (N_3632,N_3540,N_3561);
xnor U3633 (N_3633,N_3557,N_3542);
and U3634 (N_3634,N_3544,N_3577);
xnor U3635 (N_3635,N_3530,N_3572);
or U3636 (N_3636,N_3578,N_3521);
xnor U3637 (N_3637,N_3585,N_3619);
xnor U3638 (N_3638,N_3529,N_3547);
nand U3639 (N_3639,N_3580,N_3514);
nor U3640 (N_3640,N_3623,N_3515);
nor U3641 (N_3641,N_3509,N_3524);
xor U3642 (N_3642,N_3512,N_3546);
and U3643 (N_3643,N_3537,N_3600);
xnor U3644 (N_3644,N_3549,N_3555);
nor U3645 (N_3645,N_3618,N_3596);
or U3646 (N_3646,N_3612,N_3584);
or U3647 (N_3647,N_3624,N_3541);
xor U3648 (N_3648,N_3510,N_3599);
xnor U3649 (N_3649,N_3607,N_3506);
nand U3650 (N_3650,N_3568,N_3608);
or U3651 (N_3651,N_3543,N_3566);
xnor U3652 (N_3652,N_3621,N_3552);
or U3653 (N_3653,N_3548,N_3551);
nor U3654 (N_3654,N_3613,N_3560);
xnor U3655 (N_3655,N_3587,N_3533);
or U3656 (N_3656,N_3500,N_3616);
xor U3657 (N_3657,N_3589,N_3563);
and U3658 (N_3658,N_3622,N_3528);
xnor U3659 (N_3659,N_3598,N_3603);
and U3660 (N_3660,N_3597,N_3501);
and U3661 (N_3661,N_3517,N_3606);
or U3662 (N_3662,N_3525,N_3601);
nor U3663 (N_3663,N_3610,N_3531);
nor U3664 (N_3664,N_3523,N_3575);
and U3665 (N_3665,N_3527,N_3508);
or U3666 (N_3666,N_3574,N_3522);
nor U3667 (N_3667,N_3553,N_3545);
or U3668 (N_3668,N_3564,N_3554);
nand U3669 (N_3669,N_3579,N_3573);
xnor U3670 (N_3670,N_3593,N_3615);
nor U3671 (N_3671,N_3558,N_3559);
xnor U3672 (N_3672,N_3518,N_3614);
nor U3673 (N_3673,N_3532,N_3576);
nand U3674 (N_3674,N_3588,N_3609);
or U3675 (N_3675,N_3539,N_3567);
nor U3676 (N_3676,N_3550,N_3602);
nand U3677 (N_3677,N_3611,N_3620);
nor U3678 (N_3678,N_3520,N_3565);
xor U3679 (N_3679,N_3570,N_3526);
nand U3680 (N_3680,N_3507,N_3513);
nand U3681 (N_3681,N_3502,N_3594);
nand U3682 (N_3682,N_3534,N_3592);
nand U3683 (N_3683,N_3562,N_3503);
xnor U3684 (N_3684,N_3583,N_3591);
nand U3685 (N_3685,N_3505,N_3535);
nand U3686 (N_3686,N_3519,N_3536);
nand U3687 (N_3687,N_3504,N_3597);
nand U3688 (N_3688,N_3516,N_3554);
or U3689 (N_3689,N_3609,N_3585);
nor U3690 (N_3690,N_3624,N_3535);
xor U3691 (N_3691,N_3569,N_3575);
and U3692 (N_3692,N_3577,N_3575);
and U3693 (N_3693,N_3594,N_3513);
xnor U3694 (N_3694,N_3553,N_3572);
nor U3695 (N_3695,N_3544,N_3562);
or U3696 (N_3696,N_3547,N_3555);
nand U3697 (N_3697,N_3590,N_3551);
nor U3698 (N_3698,N_3516,N_3574);
and U3699 (N_3699,N_3538,N_3620);
nor U3700 (N_3700,N_3615,N_3568);
nor U3701 (N_3701,N_3506,N_3567);
and U3702 (N_3702,N_3600,N_3571);
nor U3703 (N_3703,N_3619,N_3590);
or U3704 (N_3704,N_3568,N_3585);
or U3705 (N_3705,N_3501,N_3504);
nor U3706 (N_3706,N_3623,N_3511);
nor U3707 (N_3707,N_3617,N_3563);
and U3708 (N_3708,N_3524,N_3609);
and U3709 (N_3709,N_3603,N_3548);
or U3710 (N_3710,N_3571,N_3546);
nor U3711 (N_3711,N_3505,N_3529);
nand U3712 (N_3712,N_3548,N_3606);
nand U3713 (N_3713,N_3611,N_3564);
xor U3714 (N_3714,N_3508,N_3502);
and U3715 (N_3715,N_3572,N_3511);
nand U3716 (N_3716,N_3527,N_3598);
xor U3717 (N_3717,N_3531,N_3575);
nand U3718 (N_3718,N_3583,N_3568);
xnor U3719 (N_3719,N_3579,N_3504);
nor U3720 (N_3720,N_3518,N_3565);
and U3721 (N_3721,N_3611,N_3613);
and U3722 (N_3722,N_3520,N_3506);
or U3723 (N_3723,N_3583,N_3566);
xor U3724 (N_3724,N_3557,N_3553);
and U3725 (N_3725,N_3501,N_3529);
xnor U3726 (N_3726,N_3619,N_3559);
nand U3727 (N_3727,N_3578,N_3538);
nand U3728 (N_3728,N_3535,N_3589);
xor U3729 (N_3729,N_3614,N_3580);
nand U3730 (N_3730,N_3525,N_3562);
and U3731 (N_3731,N_3561,N_3524);
or U3732 (N_3732,N_3502,N_3580);
and U3733 (N_3733,N_3610,N_3553);
or U3734 (N_3734,N_3511,N_3603);
nand U3735 (N_3735,N_3528,N_3585);
nor U3736 (N_3736,N_3538,N_3529);
nand U3737 (N_3737,N_3591,N_3584);
and U3738 (N_3738,N_3549,N_3619);
and U3739 (N_3739,N_3611,N_3569);
nor U3740 (N_3740,N_3599,N_3570);
xor U3741 (N_3741,N_3511,N_3568);
nor U3742 (N_3742,N_3617,N_3604);
nor U3743 (N_3743,N_3557,N_3522);
and U3744 (N_3744,N_3588,N_3574);
nor U3745 (N_3745,N_3595,N_3554);
nor U3746 (N_3746,N_3613,N_3619);
or U3747 (N_3747,N_3614,N_3513);
nand U3748 (N_3748,N_3541,N_3591);
xnor U3749 (N_3749,N_3580,N_3548);
or U3750 (N_3750,N_3691,N_3748);
and U3751 (N_3751,N_3687,N_3717);
or U3752 (N_3752,N_3669,N_3629);
and U3753 (N_3753,N_3644,N_3654);
or U3754 (N_3754,N_3689,N_3722);
nor U3755 (N_3755,N_3706,N_3649);
xnor U3756 (N_3756,N_3699,N_3678);
and U3757 (N_3757,N_3676,N_3725);
and U3758 (N_3758,N_3633,N_3695);
and U3759 (N_3759,N_3635,N_3696);
xor U3760 (N_3760,N_3651,N_3673);
nand U3761 (N_3761,N_3704,N_3749);
xnor U3762 (N_3762,N_3666,N_3718);
nand U3763 (N_3763,N_3652,N_3632);
and U3764 (N_3764,N_3744,N_3721);
nor U3765 (N_3765,N_3720,N_3734);
nand U3766 (N_3766,N_3715,N_3684);
or U3767 (N_3767,N_3692,N_3735);
or U3768 (N_3768,N_3727,N_3733);
or U3769 (N_3769,N_3668,N_3698);
xor U3770 (N_3770,N_3627,N_3739);
nor U3771 (N_3771,N_3670,N_3642);
or U3772 (N_3772,N_3630,N_3643);
or U3773 (N_3773,N_3626,N_3640);
and U3774 (N_3774,N_3697,N_3660);
and U3775 (N_3775,N_3657,N_3667);
or U3776 (N_3776,N_3634,N_3679);
nor U3777 (N_3777,N_3707,N_3710);
xnor U3778 (N_3778,N_3740,N_3701);
nor U3779 (N_3779,N_3631,N_3653);
nand U3780 (N_3780,N_3694,N_3746);
xor U3781 (N_3781,N_3646,N_3636);
nor U3782 (N_3782,N_3724,N_3705);
nand U3783 (N_3783,N_3714,N_3731);
nand U3784 (N_3784,N_3650,N_3716);
or U3785 (N_3785,N_3637,N_3662);
nand U3786 (N_3786,N_3664,N_3728);
or U3787 (N_3787,N_3639,N_3690);
and U3788 (N_3788,N_3647,N_3713);
or U3789 (N_3789,N_3745,N_3625);
nand U3790 (N_3790,N_3702,N_3719);
xor U3791 (N_3791,N_3675,N_3729);
xor U3792 (N_3792,N_3747,N_3665);
xnor U3793 (N_3793,N_3685,N_3737);
or U3794 (N_3794,N_3742,N_3663);
nand U3795 (N_3795,N_3743,N_3656);
nor U3796 (N_3796,N_3655,N_3658);
nand U3797 (N_3797,N_3645,N_3681);
nand U3798 (N_3798,N_3674,N_3732);
nor U3799 (N_3799,N_3682,N_3672);
and U3800 (N_3800,N_3680,N_3736);
xnor U3801 (N_3801,N_3628,N_3686);
xor U3802 (N_3802,N_3741,N_3638);
xor U3803 (N_3803,N_3661,N_3730);
or U3804 (N_3804,N_3671,N_3648);
and U3805 (N_3805,N_3641,N_3726);
or U3806 (N_3806,N_3683,N_3708);
and U3807 (N_3807,N_3659,N_3693);
nand U3808 (N_3808,N_3703,N_3677);
xor U3809 (N_3809,N_3723,N_3688);
xnor U3810 (N_3810,N_3712,N_3700);
and U3811 (N_3811,N_3709,N_3711);
or U3812 (N_3812,N_3738,N_3688);
xor U3813 (N_3813,N_3739,N_3727);
xor U3814 (N_3814,N_3700,N_3722);
or U3815 (N_3815,N_3650,N_3678);
and U3816 (N_3816,N_3649,N_3697);
xor U3817 (N_3817,N_3739,N_3696);
xor U3818 (N_3818,N_3690,N_3741);
xor U3819 (N_3819,N_3642,N_3644);
nand U3820 (N_3820,N_3695,N_3647);
xnor U3821 (N_3821,N_3733,N_3676);
nand U3822 (N_3822,N_3649,N_3659);
and U3823 (N_3823,N_3748,N_3654);
xor U3824 (N_3824,N_3745,N_3748);
nand U3825 (N_3825,N_3667,N_3626);
and U3826 (N_3826,N_3683,N_3630);
or U3827 (N_3827,N_3662,N_3642);
nor U3828 (N_3828,N_3740,N_3714);
nor U3829 (N_3829,N_3743,N_3740);
or U3830 (N_3830,N_3723,N_3654);
xnor U3831 (N_3831,N_3672,N_3649);
nand U3832 (N_3832,N_3722,N_3674);
nand U3833 (N_3833,N_3706,N_3712);
or U3834 (N_3834,N_3708,N_3718);
nor U3835 (N_3835,N_3732,N_3676);
nand U3836 (N_3836,N_3740,N_3657);
or U3837 (N_3837,N_3627,N_3707);
nor U3838 (N_3838,N_3699,N_3704);
nand U3839 (N_3839,N_3649,N_3732);
xnor U3840 (N_3840,N_3652,N_3705);
nand U3841 (N_3841,N_3719,N_3688);
xnor U3842 (N_3842,N_3659,N_3661);
and U3843 (N_3843,N_3676,N_3632);
or U3844 (N_3844,N_3736,N_3729);
or U3845 (N_3845,N_3715,N_3739);
xnor U3846 (N_3846,N_3694,N_3666);
nor U3847 (N_3847,N_3660,N_3629);
nand U3848 (N_3848,N_3746,N_3696);
nor U3849 (N_3849,N_3643,N_3707);
nor U3850 (N_3850,N_3628,N_3747);
or U3851 (N_3851,N_3692,N_3627);
nand U3852 (N_3852,N_3702,N_3668);
and U3853 (N_3853,N_3732,N_3650);
xnor U3854 (N_3854,N_3694,N_3719);
and U3855 (N_3855,N_3713,N_3638);
nand U3856 (N_3856,N_3727,N_3712);
nand U3857 (N_3857,N_3661,N_3710);
xnor U3858 (N_3858,N_3697,N_3700);
nand U3859 (N_3859,N_3686,N_3659);
nand U3860 (N_3860,N_3739,N_3704);
or U3861 (N_3861,N_3684,N_3662);
and U3862 (N_3862,N_3634,N_3677);
nor U3863 (N_3863,N_3640,N_3659);
xnor U3864 (N_3864,N_3633,N_3661);
nand U3865 (N_3865,N_3740,N_3674);
or U3866 (N_3866,N_3681,N_3650);
xnor U3867 (N_3867,N_3719,N_3675);
and U3868 (N_3868,N_3675,N_3651);
nand U3869 (N_3869,N_3629,N_3662);
nor U3870 (N_3870,N_3697,N_3672);
and U3871 (N_3871,N_3727,N_3655);
or U3872 (N_3872,N_3741,N_3705);
or U3873 (N_3873,N_3637,N_3636);
xnor U3874 (N_3874,N_3723,N_3738);
and U3875 (N_3875,N_3806,N_3831);
and U3876 (N_3876,N_3857,N_3847);
nand U3877 (N_3877,N_3768,N_3789);
nor U3878 (N_3878,N_3792,N_3824);
xnor U3879 (N_3879,N_3849,N_3767);
xor U3880 (N_3880,N_3870,N_3828);
or U3881 (N_3881,N_3859,N_3769);
and U3882 (N_3882,N_3811,N_3752);
xor U3883 (N_3883,N_3843,N_3809);
and U3884 (N_3884,N_3755,N_3835);
nand U3885 (N_3885,N_3830,N_3786);
nor U3886 (N_3886,N_3842,N_3819);
and U3887 (N_3887,N_3832,N_3800);
or U3888 (N_3888,N_3815,N_3782);
xor U3889 (N_3889,N_3802,N_3783);
nand U3890 (N_3890,N_3814,N_3820);
nand U3891 (N_3891,N_3762,N_3764);
and U3892 (N_3892,N_3780,N_3827);
xnor U3893 (N_3893,N_3804,N_3777);
or U3894 (N_3894,N_3866,N_3781);
nand U3895 (N_3895,N_3773,N_3869);
xnor U3896 (N_3896,N_3791,N_3841);
or U3897 (N_3897,N_3779,N_3864);
xor U3898 (N_3898,N_3821,N_3837);
nor U3899 (N_3899,N_3839,N_3816);
nand U3900 (N_3900,N_3872,N_3756);
nor U3901 (N_3901,N_3860,N_3778);
nand U3902 (N_3902,N_3754,N_3763);
nor U3903 (N_3903,N_3852,N_3774);
or U3904 (N_3904,N_3868,N_3854);
or U3905 (N_3905,N_3785,N_3840);
or U3906 (N_3906,N_3797,N_3829);
nor U3907 (N_3907,N_3751,N_3784);
and U3908 (N_3908,N_3874,N_3817);
nor U3909 (N_3909,N_3848,N_3838);
nor U3910 (N_3910,N_3753,N_3836);
nor U3911 (N_3911,N_3760,N_3790);
or U3912 (N_3912,N_3787,N_3873);
or U3913 (N_3913,N_3750,N_3851);
nor U3914 (N_3914,N_3825,N_3858);
and U3915 (N_3915,N_3862,N_3776);
or U3916 (N_3916,N_3812,N_3770);
or U3917 (N_3917,N_3765,N_3865);
or U3918 (N_3918,N_3799,N_3771);
nor U3919 (N_3919,N_3833,N_3813);
nor U3920 (N_3920,N_3810,N_3823);
nor U3921 (N_3921,N_3803,N_3801);
and U3922 (N_3922,N_3805,N_3850);
or U3923 (N_3923,N_3796,N_3867);
xnor U3924 (N_3924,N_3871,N_3772);
xor U3925 (N_3925,N_3853,N_3759);
nand U3926 (N_3926,N_3758,N_3846);
and U3927 (N_3927,N_3795,N_3761);
xnor U3928 (N_3928,N_3788,N_3834);
nor U3929 (N_3929,N_3845,N_3775);
nand U3930 (N_3930,N_3766,N_3856);
nand U3931 (N_3931,N_3861,N_3794);
nor U3932 (N_3932,N_3822,N_3807);
nand U3933 (N_3933,N_3863,N_3826);
xnor U3934 (N_3934,N_3844,N_3798);
nor U3935 (N_3935,N_3793,N_3818);
or U3936 (N_3936,N_3808,N_3757);
nand U3937 (N_3937,N_3855,N_3846);
or U3938 (N_3938,N_3832,N_3764);
nand U3939 (N_3939,N_3857,N_3854);
or U3940 (N_3940,N_3799,N_3862);
and U3941 (N_3941,N_3834,N_3820);
nand U3942 (N_3942,N_3792,N_3844);
or U3943 (N_3943,N_3785,N_3849);
or U3944 (N_3944,N_3789,N_3868);
nor U3945 (N_3945,N_3790,N_3797);
xor U3946 (N_3946,N_3796,N_3778);
nand U3947 (N_3947,N_3868,N_3795);
nand U3948 (N_3948,N_3860,N_3815);
or U3949 (N_3949,N_3861,N_3782);
or U3950 (N_3950,N_3839,N_3873);
nand U3951 (N_3951,N_3867,N_3799);
nand U3952 (N_3952,N_3840,N_3771);
xor U3953 (N_3953,N_3755,N_3767);
and U3954 (N_3954,N_3838,N_3751);
xor U3955 (N_3955,N_3843,N_3804);
nor U3956 (N_3956,N_3827,N_3758);
xor U3957 (N_3957,N_3810,N_3763);
xnor U3958 (N_3958,N_3799,N_3825);
or U3959 (N_3959,N_3844,N_3851);
and U3960 (N_3960,N_3771,N_3854);
nor U3961 (N_3961,N_3831,N_3766);
nor U3962 (N_3962,N_3766,N_3848);
nor U3963 (N_3963,N_3765,N_3813);
and U3964 (N_3964,N_3826,N_3801);
and U3965 (N_3965,N_3813,N_3787);
nand U3966 (N_3966,N_3869,N_3846);
or U3967 (N_3967,N_3844,N_3867);
and U3968 (N_3968,N_3823,N_3859);
xor U3969 (N_3969,N_3861,N_3789);
nor U3970 (N_3970,N_3767,N_3811);
nor U3971 (N_3971,N_3857,N_3826);
nor U3972 (N_3972,N_3785,N_3872);
nand U3973 (N_3973,N_3821,N_3756);
or U3974 (N_3974,N_3872,N_3806);
nor U3975 (N_3975,N_3804,N_3819);
nor U3976 (N_3976,N_3811,N_3833);
or U3977 (N_3977,N_3865,N_3874);
and U3978 (N_3978,N_3840,N_3867);
xor U3979 (N_3979,N_3863,N_3823);
xnor U3980 (N_3980,N_3820,N_3851);
or U3981 (N_3981,N_3762,N_3780);
and U3982 (N_3982,N_3799,N_3764);
nor U3983 (N_3983,N_3848,N_3830);
nor U3984 (N_3984,N_3869,N_3790);
and U3985 (N_3985,N_3763,N_3823);
nor U3986 (N_3986,N_3834,N_3842);
and U3987 (N_3987,N_3773,N_3785);
nand U3988 (N_3988,N_3792,N_3754);
or U3989 (N_3989,N_3794,N_3843);
or U3990 (N_3990,N_3791,N_3829);
nand U3991 (N_3991,N_3802,N_3826);
nand U3992 (N_3992,N_3788,N_3762);
nor U3993 (N_3993,N_3760,N_3751);
nand U3994 (N_3994,N_3809,N_3856);
or U3995 (N_3995,N_3783,N_3773);
and U3996 (N_3996,N_3808,N_3825);
nor U3997 (N_3997,N_3800,N_3756);
or U3998 (N_3998,N_3820,N_3772);
nand U3999 (N_3999,N_3783,N_3860);
or U4000 (N_4000,N_3906,N_3989);
nor U4001 (N_4001,N_3986,N_3933);
and U4002 (N_4002,N_3974,N_3919);
xor U4003 (N_4003,N_3975,N_3963);
or U4004 (N_4004,N_3969,N_3927);
or U4005 (N_4005,N_3924,N_3903);
nand U4006 (N_4006,N_3920,N_3971);
nor U4007 (N_4007,N_3943,N_3931);
or U4008 (N_4008,N_3939,N_3904);
nand U4009 (N_4009,N_3957,N_3911);
nor U4010 (N_4010,N_3944,N_3973);
xnor U4011 (N_4011,N_3886,N_3949);
nor U4012 (N_4012,N_3896,N_3916);
nand U4013 (N_4013,N_3994,N_3895);
xor U4014 (N_4014,N_3995,N_3992);
xor U4015 (N_4015,N_3999,N_3953);
and U4016 (N_4016,N_3898,N_3936);
nor U4017 (N_4017,N_3976,N_3908);
nand U4018 (N_4018,N_3978,N_3991);
nor U4019 (N_4019,N_3954,N_3902);
nand U4020 (N_4020,N_3942,N_3889);
or U4021 (N_4021,N_3948,N_3882);
nand U4022 (N_4022,N_3941,N_3979);
or U4023 (N_4023,N_3985,N_3909);
or U4024 (N_4024,N_3968,N_3937);
nand U4025 (N_4025,N_3959,N_3929);
or U4026 (N_4026,N_3984,N_3901);
or U4027 (N_4027,N_3878,N_3952);
xnor U4028 (N_4028,N_3883,N_3890);
and U4029 (N_4029,N_3900,N_3998);
and U4030 (N_4030,N_3996,N_3893);
or U4031 (N_4031,N_3956,N_3928);
and U4032 (N_4032,N_3932,N_3977);
xnor U4033 (N_4033,N_3970,N_3938);
and U4034 (N_4034,N_3972,N_3881);
or U4035 (N_4035,N_3982,N_3988);
xor U4036 (N_4036,N_3987,N_3950);
nand U4037 (N_4037,N_3915,N_3934);
nor U4038 (N_4038,N_3997,N_3923);
xnor U4039 (N_4039,N_3892,N_3981);
xor U4040 (N_4040,N_3940,N_3912);
nand U4041 (N_4041,N_3885,N_3897);
nand U4042 (N_4042,N_3990,N_3913);
or U4043 (N_4043,N_3961,N_3879);
and U4044 (N_4044,N_3960,N_3930);
or U4045 (N_4045,N_3955,N_3917);
nor U4046 (N_4046,N_3910,N_3921);
nand U4047 (N_4047,N_3891,N_3980);
nor U4048 (N_4048,N_3967,N_3899);
nand U4049 (N_4049,N_3884,N_3945);
nand U4050 (N_4050,N_3965,N_3946);
xnor U4051 (N_4051,N_3983,N_3926);
xor U4052 (N_4052,N_3887,N_3962);
nor U4053 (N_4053,N_3966,N_3958);
xor U4054 (N_4054,N_3876,N_3888);
and U4055 (N_4055,N_3935,N_3905);
xnor U4056 (N_4056,N_3907,N_3914);
nor U4057 (N_4057,N_3993,N_3877);
nor U4058 (N_4058,N_3925,N_3918);
and U4059 (N_4059,N_3947,N_3951);
and U4060 (N_4060,N_3875,N_3894);
or U4061 (N_4061,N_3880,N_3964);
nor U4062 (N_4062,N_3922,N_3905);
nor U4063 (N_4063,N_3973,N_3877);
nor U4064 (N_4064,N_3948,N_3935);
nand U4065 (N_4065,N_3943,N_3994);
nand U4066 (N_4066,N_3909,N_3924);
xor U4067 (N_4067,N_3983,N_3912);
nand U4068 (N_4068,N_3928,N_3955);
and U4069 (N_4069,N_3879,N_3892);
and U4070 (N_4070,N_3969,N_3950);
or U4071 (N_4071,N_3951,N_3925);
xor U4072 (N_4072,N_3967,N_3897);
nor U4073 (N_4073,N_3952,N_3877);
nor U4074 (N_4074,N_3921,N_3988);
xnor U4075 (N_4075,N_3883,N_3879);
nand U4076 (N_4076,N_3945,N_3938);
and U4077 (N_4077,N_3931,N_3885);
nand U4078 (N_4078,N_3970,N_3896);
or U4079 (N_4079,N_3992,N_3922);
nand U4080 (N_4080,N_3995,N_3970);
nor U4081 (N_4081,N_3977,N_3970);
nor U4082 (N_4082,N_3905,N_3964);
and U4083 (N_4083,N_3875,N_3889);
xnor U4084 (N_4084,N_3905,N_3875);
and U4085 (N_4085,N_3966,N_3981);
xnor U4086 (N_4086,N_3897,N_3988);
nor U4087 (N_4087,N_3918,N_3910);
nand U4088 (N_4088,N_3925,N_3961);
and U4089 (N_4089,N_3893,N_3897);
and U4090 (N_4090,N_3928,N_3876);
nor U4091 (N_4091,N_3921,N_3936);
xor U4092 (N_4092,N_3983,N_3940);
nor U4093 (N_4093,N_3991,N_3890);
nand U4094 (N_4094,N_3909,N_3923);
nand U4095 (N_4095,N_3904,N_3950);
xor U4096 (N_4096,N_3996,N_3902);
nor U4097 (N_4097,N_3881,N_3894);
xor U4098 (N_4098,N_3979,N_3997);
or U4099 (N_4099,N_3963,N_3978);
nor U4100 (N_4100,N_3943,N_3988);
xor U4101 (N_4101,N_3958,N_3889);
nand U4102 (N_4102,N_3976,N_3941);
or U4103 (N_4103,N_3902,N_3913);
and U4104 (N_4104,N_3941,N_3890);
or U4105 (N_4105,N_3983,N_3903);
and U4106 (N_4106,N_3890,N_3936);
xor U4107 (N_4107,N_3881,N_3909);
xor U4108 (N_4108,N_3984,N_3916);
xnor U4109 (N_4109,N_3927,N_3971);
nor U4110 (N_4110,N_3891,N_3949);
or U4111 (N_4111,N_3883,N_3994);
or U4112 (N_4112,N_3945,N_3919);
nand U4113 (N_4113,N_3904,N_3962);
or U4114 (N_4114,N_3900,N_3940);
xnor U4115 (N_4115,N_3955,N_3974);
and U4116 (N_4116,N_3921,N_3908);
nor U4117 (N_4117,N_3956,N_3909);
nor U4118 (N_4118,N_3995,N_3914);
nor U4119 (N_4119,N_3968,N_3974);
and U4120 (N_4120,N_3890,N_3998);
or U4121 (N_4121,N_3886,N_3979);
nand U4122 (N_4122,N_3981,N_3934);
nor U4123 (N_4123,N_3947,N_3962);
and U4124 (N_4124,N_3920,N_3933);
nor U4125 (N_4125,N_4019,N_4037);
or U4126 (N_4126,N_4026,N_4007);
nand U4127 (N_4127,N_4120,N_4067);
nand U4128 (N_4128,N_4122,N_4113);
or U4129 (N_4129,N_4069,N_4017);
xor U4130 (N_4130,N_4048,N_4039);
nor U4131 (N_4131,N_4032,N_4095);
xor U4132 (N_4132,N_4035,N_4005);
and U4133 (N_4133,N_4055,N_4022);
nand U4134 (N_4134,N_4118,N_4042);
nand U4135 (N_4135,N_4115,N_4104);
nand U4136 (N_4136,N_4066,N_4085);
nand U4137 (N_4137,N_4068,N_4056);
nor U4138 (N_4138,N_4082,N_4029);
or U4139 (N_4139,N_4094,N_4077);
and U4140 (N_4140,N_4053,N_4052);
nand U4141 (N_4141,N_4074,N_4083);
nand U4142 (N_4142,N_4025,N_4065);
and U4143 (N_4143,N_4008,N_4112);
nand U4144 (N_4144,N_4090,N_4108);
and U4145 (N_4145,N_4121,N_4107);
xor U4146 (N_4146,N_4078,N_4038);
and U4147 (N_4147,N_4089,N_4073);
xor U4148 (N_4148,N_4111,N_4041);
and U4149 (N_4149,N_4015,N_4043);
and U4150 (N_4150,N_4109,N_4002);
and U4151 (N_4151,N_4106,N_4098);
nand U4152 (N_4152,N_4027,N_4096);
and U4153 (N_4153,N_4004,N_4000);
xnor U4154 (N_4154,N_4014,N_4088);
or U4155 (N_4155,N_4024,N_4110);
nor U4156 (N_4156,N_4086,N_4080);
nor U4157 (N_4157,N_4058,N_4105);
or U4158 (N_4158,N_4040,N_4051);
xor U4159 (N_4159,N_4020,N_4023);
xnor U4160 (N_4160,N_4124,N_4079);
nor U4161 (N_4161,N_4030,N_4063);
nand U4162 (N_4162,N_4009,N_4123);
nor U4163 (N_4163,N_4054,N_4100);
nand U4164 (N_4164,N_4046,N_4116);
xnor U4165 (N_4165,N_4033,N_4064);
nand U4166 (N_4166,N_4018,N_4091);
nor U4167 (N_4167,N_4001,N_4031);
nor U4168 (N_4168,N_4013,N_4117);
and U4169 (N_4169,N_4102,N_4072);
xor U4170 (N_4170,N_4061,N_4070);
nor U4171 (N_4171,N_4003,N_4101);
or U4172 (N_4172,N_4087,N_4049);
and U4173 (N_4173,N_4010,N_4092);
and U4174 (N_4174,N_4034,N_4012);
xnor U4175 (N_4175,N_4071,N_4097);
nor U4176 (N_4176,N_4011,N_4021);
nor U4177 (N_4177,N_4016,N_4084);
and U4178 (N_4178,N_4036,N_4075);
xor U4179 (N_4179,N_4057,N_4103);
nor U4180 (N_4180,N_4114,N_4081);
nor U4181 (N_4181,N_4028,N_4044);
and U4182 (N_4182,N_4076,N_4050);
nand U4183 (N_4183,N_4062,N_4093);
nor U4184 (N_4184,N_4045,N_4060);
nand U4185 (N_4185,N_4119,N_4047);
nor U4186 (N_4186,N_4099,N_4059);
and U4187 (N_4187,N_4006,N_4115);
nor U4188 (N_4188,N_4102,N_4006);
or U4189 (N_4189,N_4016,N_4110);
or U4190 (N_4190,N_4049,N_4104);
xnor U4191 (N_4191,N_4076,N_4038);
nand U4192 (N_4192,N_4112,N_4046);
and U4193 (N_4193,N_4067,N_4030);
or U4194 (N_4194,N_4002,N_4104);
or U4195 (N_4195,N_4045,N_4017);
and U4196 (N_4196,N_4017,N_4060);
and U4197 (N_4197,N_4119,N_4002);
xor U4198 (N_4198,N_4076,N_4012);
nor U4199 (N_4199,N_4017,N_4117);
and U4200 (N_4200,N_4089,N_4011);
and U4201 (N_4201,N_4031,N_4067);
nand U4202 (N_4202,N_4118,N_4081);
xnor U4203 (N_4203,N_4117,N_4076);
and U4204 (N_4204,N_4088,N_4009);
and U4205 (N_4205,N_4008,N_4051);
and U4206 (N_4206,N_4043,N_4020);
nor U4207 (N_4207,N_4025,N_4004);
nand U4208 (N_4208,N_4060,N_4072);
or U4209 (N_4209,N_4074,N_4080);
nand U4210 (N_4210,N_4062,N_4016);
nand U4211 (N_4211,N_4103,N_4115);
nand U4212 (N_4212,N_4078,N_4069);
and U4213 (N_4213,N_4043,N_4071);
nand U4214 (N_4214,N_4043,N_4051);
nor U4215 (N_4215,N_4052,N_4098);
or U4216 (N_4216,N_4057,N_4065);
nor U4217 (N_4217,N_4062,N_4117);
nor U4218 (N_4218,N_4023,N_4056);
xor U4219 (N_4219,N_4056,N_4031);
nor U4220 (N_4220,N_4119,N_4082);
nand U4221 (N_4221,N_4058,N_4047);
xnor U4222 (N_4222,N_4099,N_4004);
and U4223 (N_4223,N_4084,N_4052);
or U4224 (N_4224,N_4076,N_4068);
and U4225 (N_4225,N_4016,N_4113);
and U4226 (N_4226,N_4096,N_4118);
and U4227 (N_4227,N_4014,N_4033);
or U4228 (N_4228,N_4005,N_4078);
nor U4229 (N_4229,N_4037,N_4047);
xnor U4230 (N_4230,N_4088,N_4076);
nor U4231 (N_4231,N_4065,N_4000);
or U4232 (N_4232,N_4092,N_4029);
and U4233 (N_4233,N_4061,N_4114);
or U4234 (N_4234,N_4037,N_4041);
nand U4235 (N_4235,N_4015,N_4108);
nor U4236 (N_4236,N_4048,N_4115);
and U4237 (N_4237,N_4001,N_4108);
and U4238 (N_4238,N_4025,N_4015);
and U4239 (N_4239,N_4111,N_4042);
and U4240 (N_4240,N_4106,N_4075);
nand U4241 (N_4241,N_4024,N_4116);
nor U4242 (N_4242,N_4048,N_4037);
nand U4243 (N_4243,N_4112,N_4061);
nor U4244 (N_4244,N_4054,N_4079);
or U4245 (N_4245,N_4055,N_4052);
and U4246 (N_4246,N_4000,N_4119);
xor U4247 (N_4247,N_4043,N_4055);
or U4248 (N_4248,N_4089,N_4065);
and U4249 (N_4249,N_4038,N_4018);
xor U4250 (N_4250,N_4133,N_4245);
or U4251 (N_4251,N_4129,N_4209);
nor U4252 (N_4252,N_4130,N_4193);
and U4253 (N_4253,N_4192,N_4226);
nand U4254 (N_4254,N_4221,N_4240);
xor U4255 (N_4255,N_4212,N_4153);
nor U4256 (N_4256,N_4154,N_4249);
nor U4257 (N_4257,N_4207,N_4224);
nor U4258 (N_4258,N_4196,N_4143);
nand U4259 (N_4259,N_4204,N_4148);
nand U4260 (N_4260,N_4201,N_4132);
or U4261 (N_4261,N_4195,N_4203);
and U4262 (N_4262,N_4131,N_4223);
xor U4263 (N_4263,N_4210,N_4172);
or U4264 (N_4264,N_4231,N_4241);
nand U4265 (N_4265,N_4137,N_4167);
nor U4266 (N_4266,N_4228,N_4141);
nand U4267 (N_4267,N_4181,N_4227);
xor U4268 (N_4268,N_4162,N_4235);
or U4269 (N_4269,N_4238,N_4244);
and U4270 (N_4270,N_4215,N_4247);
and U4271 (N_4271,N_4177,N_4179);
or U4272 (N_4272,N_4234,N_4222);
and U4273 (N_4273,N_4173,N_4211);
nor U4274 (N_4274,N_4145,N_4152);
or U4275 (N_4275,N_4135,N_4164);
xor U4276 (N_4276,N_4242,N_4134);
nand U4277 (N_4277,N_4155,N_4198);
nor U4278 (N_4278,N_4197,N_4170);
or U4279 (N_4279,N_4166,N_4205);
xor U4280 (N_4280,N_4237,N_4146);
or U4281 (N_4281,N_4208,N_4144);
and U4282 (N_4282,N_4230,N_4220);
and U4283 (N_4283,N_4236,N_4246);
nor U4284 (N_4284,N_4126,N_4142);
nand U4285 (N_4285,N_4199,N_4190);
and U4286 (N_4286,N_4157,N_4171);
nor U4287 (N_4287,N_4229,N_4186);
nand U4288 (N_4288,N_4139,N_4185);
nand U4289 (N_4289,N_4183,N_4176);
nor U4290 (N_4290,N_4213,N_4202);
nor U4291 (N_4291,N_4232,N_4169);
xor U4292 (N_4292,N_4165,N_4138);
nand U4293 (N_4293,N_4159,N_4161);
xor U4294 (N_4294,N_4150,N_4200);
or U4295 (N_4295,N_4214,N_4180);
nor U4296 (N_4296,N_4156,N_4216);
or U4297 (N_4297,N_4160,N_4149);
and U4298 (N_4298,N_4248,N_4125);
nor U4299 (N_4299,N_4158,N_4218);
xnor U4300 (N_4300,N_4194,N_4178);
nor U4301 (N_4301,N_4191,N_4243);
nand U4302 (N_4302,N_4187,N_4219);
nor U4303 (N_4303,N_4147,N_4188);
nand U4304 (N_4304,N_4127,N_4233);
nand U4305 (N_4305,N_4225,N_4239);
xor U4306 (N_4306,N_4174,N_4189);
and U4307 (N_4307,N_4182,N_4151);
xor U4308 (N_4308,N_4217,N_4175);
xor U4309 (N_4309,N_4128,N_4168);
nand U4310 (N_4310,N_4184,N_4140);
nor U4311 (N_4311,N_4136,N_4163);
nand U4312 (N_4312,N_4206,N_4239);
or U4313 (N_4313,N_4146,N_4169);
and U4314 (N_4314,N_4176,N_4147);
and U4315 (N_4315,N_4142,N_4170);
nand U4316 (N_4316,N_4139,N_4200);
or U4317 (N_4317,N_4192,N_4133);
nand U4318 (N_4318,N_4144,N_4151);
xnor U4319 (N_4319,N_4223,N_4132);
and U4320 (N_4320,N_4190,N_4230);
nand U4321 (N_4321,N_4125,N_4220);
nor U4322 (N_4322,N_4218,N_4211);
nor U4323 (N_4323,N_4140,N_4233);
or U4324 (N_4324,N_4210,N_4183);
nand U4325 (N_4325,N_4195,N_4213);
or U4326 (N_4326,N_4234,N_4143);
or U4327 (N_4327,N_4205,N_4193);
nand U4328 (N_4328,N_4199,N_4233);
and U4329 (N_4329,N_4170,N_4231);
or U4330 (N_4330,N_4134,N_4244);
nor U4331 (N_4331,N_4185,N_4158);
xnor U4332 (N_4332,N_4154,N_4174);
or U4333 (N_4333,N_4149,N_4182);
or U4334 (N_4334,N_4149,N_4170);
nor U4335 (N_4335,N_4127,N_4205);
and U4336 (N_4336,N_4137,N_4129);
and U4337 (N_4337,N_4188,N_4133);
and U4338 (N_4338,N_4197,N_4225);
or U4339 (N_4339,N_4237,N_4205);
or U4340 (N_4340,N_4160,N_4153);
nand U4341 (N_4341,N_4166,N_4135);
xnor U4342 (N_4342,N_4133,N_4211);
nor U4343 (N_4343,N_4235,N_4131);
xor U4344 (N_4344,N_4224,N_4169);
nor U4345 (N_4345,N_4139,N_4249);
nand U4346 (N_4346,N_4140,N_4195);
nor U4347 (N_4347,N_4126,N_4248);
and U4348 (N_4348,N_4161,N_4190);
nor U4349 (N_4349,N_4180,N_4162);
or U4350 (N_4350,N_4249,N_4159);
and U4351 (N_4351,N_4207,N_4160);
nor U4352 (N_4352,N_4172,N_4166);
or U4353 (N_4353,N_4141,N_4243);
and U4354 (N_4354,N_4200,N_4175);
nor U4355 (N_4355,N_4135,N_4147);
xor U4356 (N_4356,N_4148,N_4145);
nor U4357 (N_4357,N_4197,N_4137);
and U4358 (N_4358,N_4224,N_4130);
nand U4359 (N_4359,N_4223,N_4237);
nand U4360 (N_4360,N_4179,N_4196);
nand U4361 (N_4361,N_4157,N_4239);
or U4362 (N_4362,N_4142,N_4215);
and U4363 (N_4363,N_4163,N_4213);
or U4364 (N_4364,N_4243,N_4205);
and U4365 (N_4365,N_4210,N_4156);
nand U4366 (N_4366,N_4146,N_4210);
or U4367 (N_4367,N_4167,N_4149);
and U4368 (N_4368,N_4235,N_4191);
or U4369 (N_4369,N_4130,N_4173);
xnor U4370 (N_4370,N_4223,N_4169);
xnor U4371 (N_4371,N_4209,N_4240);
xor U4372 (N_4372,N_4201,N_4164);
nor U4373 (N_4373,N_4212,N_4239);
nor U4374 (N_4374,N_4137,N_4242);
nand U4375 (N_4375,N_4263,N_4303);
nand U4376 (N_4376,N_4269,N_4324);
xor U4377 (N_4377,N_4267,N_4316);
nand U4378 (N_4378,N_4308,N_4331);
or U4379 (N_4379,N_4262,N_4306);
and U4380 (N_4380,N_4360,N_4260);
or U4381 (N_4381,N_4334,N_4340);
or U4382 (N_4382,N_4284,N_4250);
or U4383 (N_4383,N_4319,N_4300);
or U4384 (N_4384,N_4295,N_4372);
and U4385 (N_4385,N_4281,N_4365);
xor U4386 (N_4386,N_4325,N_4348);
nor U4387 (N_4387,N_4353,N_4330);
xor U4388 (N_4388,N_4251,N_4302);
nand U4389 (N_4389,N_4321,N_4339);
xnor U4390 (N_4390,N_4282,N_4320);
and U4391 (N_4391,N_4307,N_4374);
nand U4392 (N_4392,N_4350,N_4294);
nor U4393 (N_4393,N_4346,N_4305);
nand U4394 (N_4394,N_4253,N_4332);
or U4395 (N_4395,N_4371,N_4259);
or U4396 (N_4396,N_4264,N_4291);
nor U4397 (N_4397,N_4257,N_4337);
xor U4398 (N_4398,N_4285,N_4347);
nor U4399 (N_4399,N_4317,N_4278);
or U4400 (N_4400,N_4361,N_4256);
xor U4401 (N_4401,N_4275,N_4266);
or U4402 (N_4402,N_4351,N_4280);
or U4403 (N_4403,N_4369,N_4314);
nor U4404 (N_4404,N_4289,N_4363);
nor U4405 (N_4405,N_4318,N_4327);
xor U4406 (N_4406,N_4315,N_4287);
xnor U4407 (N_4407,N_4370,N_4286);
nand U4408 (N_4408,N_4368,N_4310);
or U4409 (N_4409,N_4341,N_4312);
xor U4410 (N_4410,N_4359,N_4254);
and U4411 (N_4411,N_4288,N_4276);
nand U4412 (N_4412,N_4356,N_4342);
and U4413 (N_4413,N_4279,N_4367);
and U4414 (N_4414,N_4358,N_4355);
nand U4415 (N_4415,N_4336,N_4364);
nor U4416 (N_4416,N_4283,N_4373);
xor U4417 (N_4417,N_4338,N_4297);
nor U4418 (N_4418,N_4329,N_4345);
or U4419 (N_4419,N_4270,N_4328);
or U4420 (N_4420,N_4301,N_4296);
nand U4421 (N_4421,N_4357,N_4298);
nand U4422 (N_4422,N_4366,N_4309);
or U4423 (N_4423,N_4326,N_4258);
xnor U4424 (N_4424,N_4349,N_4277);
nand U4425 (N_4425,N_4292,N_4273);
and U4426 (N_4426,N_4343,N_4261);
nor U4427 (N_4427,N_4344,N_4352);
or U4428 (N_4428,N_4333,N_4272);
or U4429 (N_4429,N_4299,N_4354);
and U4430 (N_4430,N_4274,N_4323);
xnor U4431 (N_4431,N_4271,N_4290);
nor U4432 (N_4432,N_4255,N_4335);
and U4433 (N_4433,N_4265,N_4293);
and U4434 (N_4434,N_4311,N_4268);
xnor U4435 (N_4435,N_4322,N_4304);
nor U4436 (N_4436,N_4362,N_4313);
and U4437 (N_4437,N_4252,N_4345);
nor U4438 (N_4438,N_4286,N_4365);
nand U4439 (N_4439,N_4313,N_4355);
xnor U4440 (N_4440,N_4273,N_4333);
xnor U4441 (N_4441,N_4310,N_4373);
and U4442 (N_4442,N_4344,N_4362);
xor U4443 (N_4443,N_4342,N_4264);
and U4444 (N_4444,N_4281,N_4285);
or U4445 (N_4445,N_4327,N_4293);
and U4446 (N_4446,N_4272,N_4365);
or U4447 (N_4447,N_4254,N_4271);
xnor U4448 (N_4448,N_4250,N_4365);
and U4449 (N_4449,N_4368,N_4373);
nand U4450 (N_4450,N_4362,N_4292);
xor U4451 (N_4451,N_4341,N_4360);
and U4452 (N_4452,N_4323,N_4321);
nor U4453 (N_4453,N_4299,N_4350);
xor U4454 (N_4454,N_4313,N_4260);
or U4455 (N_4455,N_4329,N_4343);
nor U4456 (N_4456,N_4273,N_4332);
or U4457 (N_4457,N_4282,N_4368);
and U4458 (N_4458,N_4349,N_4333);
or U4459 (N_4459,N_4282,N_4374);
nor U4460 (N_4460,N_4285,N_4269);
xnor U4461 (N_4461,N_4294,N_4333);
and U4462 (N_4462,N_4260,N_4270);
xor U4463 (N_4463,N_4371,N_4270);
or U4464 (N_4464,N_4299,N_4251);
xor U4465 (N_4465,N_4364,N_4255);
and U4466 (N_4466,N_4348,N_4341);
nor U4467 (N_4467,N_4251,N_4366);
and U4468 (N_4468,N_4287,N_4286);
nand U4469 (N_4469,N_4255,N_4251);
or U4470 (N_4470,N_4366,N_4373);
or U4471 (N_4471,N_4350,N_4331);
and U4472 (N_4472,N_4332,N_4254);
nor U4473 (N_4473,N_4329,N_4330);
or U4474 (N_4474,N_4252,N_4312);
nor U4475 (N_4475,N_4325,N_4284);
or U4476 (N_4476,N_4277,N_4280);
or U4477 (N_4477,N_4266,N_4372);
nand U4478 (N_4478,N_4278,N_4253);
or U4479 (N_4479,N_4267,N_4280);
xor U4480 (N_4480,N_4371,N_4352);
nor U4481 (N_4481,N_4342,N_4315);
nand U4482 (N_4482,N_4277,N_4274);
xor U4483 (N_4483,N_4369,N_4290);
xnor U4484 (N_4484,N_4287,N_4336);
and U4485 (N_4485,N_4343,N_4318);
xnor U4486 (N_4486,N_4363,N_4323);
xor U4487 (N_4487,N_4253,N_4314);
and U4488 (N_4488,N_4340,N_4359);
nand U4489 (N_4489,N_4312,N_4331);
xor U4490 (N_4490,N_4267,N_4270);
nand U4491 (N_4491,N_4309,N_4334);
xnor U4492 (N_4492,N_4266,N_4283);
or U4493 (N_4493,N_4356,N_4363);
nor U4494 (N_4494,N_4327,N_4302);
and U4495 (N_4495,N_4269,N_4360);
xor U4496 (N_4496,N_4266,N_4354);
or U4497 (N_4497,N_4342,N_4365);
or U4498 (N_4498,N_4344,N_4257);
and U4499 (N_4499,N_4354,N_4318);
or U4500 (N_4500,N_4473,N_4492);
nor U4501 (N_4501,N_4445,N_4474);
and U4502 (N_4502,N_4449,N_4465);
nand U4503 (N_4503,N_4427,N_4454);
xor U4504 (N_4504,N_4419,N_4447);
nor U4505 (N_4505,N_4446,N_4420);
and U4506 (N_4506,N_4382,N_4402);
and U4507 (N_4507,N_4455,N_4493);
nor U4508 (N_4508,N_4470,N_4375);
xor U4509 (N_4509,N_4451,N_4387);
xnor U4510 (N_4510,N_4411,N_4464);
xor U4511 (N_4511,N_4389,N_4456);
xor U4512 (N_4512,N_4472,N_4439);
nand U4513 (N_4513,N_4421,N_4378);
and U4514 (N_4514,N_4475,N_4448);
xor U4515 (N_4515,N_4435,N_4380);
nand U4516 (N_4516,N_4488,N_4407);
or U4517 (N_4517,N_4476,N_4499);
nand U4518 (N_4518,N_4482,N_4422);
xor U4519 (N_4519,N_4392,N_4377);
and U4520 (N_4520,N_4381,N_4404);
nand U4521 (N_4521,N_4414,N_4403);
and U4522 (N_4522,N_4415,N_4489);
nand U4523 (N_4523,N_4486,N_4408);
nor U4524 (N_4524,N_4497,N_4494);
or U4525 (N_4525,N_4401,N_4416);
and U4526 (N_4526,N_4491,N_4483);
or U4527 (N_4527,N_4406,N_4394);
nand U4528 (N_4528,N_4490,N_4400);
nand U4529 (N_4529,N_4441,N_4484);
nor U4530 (N_4530,N_4385,N_4399);
xnor U4531 (N_4531,N_4481,N_4405);
and U4532 (N_4532,N_4383,N_4461);
or U4533 (N_4533,N_4477,N_4478);
and U4534 (N_4534,N_4384,N_4452);
and U4535 (N_4535,N_4432,N_4480);
nand U4536 (N_4536,N_4430,N_4424);
or U4537 (N_4537,N_4417,N_4434);
or U4538 (N_4538,N_4467,N_4443);
nand U4539 (N_4539,N_4431,N_4460);
or U4540 (N_4540,N_4463,N_4450);
or U4541 (N_4541,N_4438,N_4457);
nor U4542 (N_4542,N_4388,N_4469);
nor U4543 (N_4543,N_4468,N_4386);
and U4544 (N_4544,N_4413,N_4487);
and U4545 (N_4545,N_4485,N_4410);
and U4546 (N_4546,N_4395,N_4496);
or U4547 (N_4547,N_4390,N_4458);
nor U4548 (N_4548,N_4453,N_4442);
xnor U4549 (N_4549,N_4428,N_4479);
or U4550 (N_4550,N_4379,N_4436);
or U4551 (N_4551,N_4397,N_4471);
xnor U4552 (N_4552,N_4498,N_4433);
and U4553 (N_4553,N_4423,N_4444);
nand U4554 (N_4554,N_4466,N_4391);
nor U4555 (N_4555,N_4412,N_4393);
or U4556 (N_4556,N_4425,N_4495);
nand U4557 (N_4557,N_4418,N_4409);
and U4558 (N_4558,N_4462,N_4426);
xnor U4559 (N_4559,N_4376,N_4398);
or U4560 (N_4560,N_4429,N_4396);
or U4561 (N_4561,N_4440,N_4459);
xor U4562 (N_4562,N_4437,N_4376);
nand U4563 (N_4563,N_4427,N_4440);
xor U4564 (N_4564,N_4453,N_4396);
nor U4565 (N_4565,N_4462,N_4442);
xor U4566 (N_4566,N_4482,N_4391);
or U4567 (N_4567,N_4479,N_4490);
nor U4568 (N_4568,N_4416,N_4409);
nand U4569 (N_4569,N_4446,N_4479);
nand U4570 (N_4570,N_4380,N_4465);
and U4571 (N_4571,N_4485,N_4392);
and U4572 (N_4572,N_4410,N_4399);
nand U4573 (N_4573,N_4434,N_4483);
nor U4574 (N_4574,N_4419,N_4418);
xnor U4575 (N_4575,N_4440,N_4452);
xnor U4576 (N_4576,N_4409,N_4461);
nand U4577 (N_4577,N_4399,N_4463);
nand U4578 (N_4578,N_4442,N_4412);
nor U4579 (N_4579,N_4478,N_4492);
xor U4580 (N_4580,N_4474,N_4405);
or U4581 (N_4581,N_4388,N_4460);
xor U4582 (N_4582,N_4489,N_4492);
or U4583 (N_4583,N_4459,N_4376);
nand U4584 (N_4584,N_4376,N_4395);
nor U4585 (N_4585,N_4476,N_4472);
nor U4586 (N_4586,N_4397,N_4465);
and U4587 (N_4587,N_4490,N_4496);
xnor U4588 (N_4588,N_4468,N_4389);
nand U4589 (N_4589,N_4398,N_4391);
xor U4590 (N_4590,N_4442,N_4483);
or U4591 (N_4591,N_4437,N_4404);
xor U4592 (N_4592,N_4471,N_4473);
and U4593 (N_4593,N_4462,N_4479);
and U4594 (N_4594,N_4439,N_4478);
nor U4595 (N_4595,N_4483,N_4414);
or U4596 (N_4596,N_4463,N_4426);
nor U4597 (N_4597,N_4382,N_4473);
or U4598 (N_4598,N_4490,N_4420);
or U4599 (N_4599,N_4414,N_4465);
nand U4600 (N_4600,N_4430,N_4496);
and U4601 (N_4601,N_4446,N_4495);
nor U4602 (N_4602,N_4431,N_4386);
and U4603 (N_4603,N_4464,N_4397);
nand U4604 (N_4604,N_4494,N_4475);
nor U4605 (N_4605,N_4377,N_4444);
nand U4606 (N_4606,N_4438,N_4420);
or U4607 (N_4607,N_4441,N_4499);
xnor U4608 (N_4608,N_4433,N_4390);
nor U4609 (N_4609,N_4442,N_4394);
nand U4610 (N_4610,N_4409,N_4427);
or U4611 (N_4611,N_4452,N_4434);
and U4612 (N_4612,N_4445,N_4410);
and U4613 (N_4613,N_4417,N_4411);
nor U4614 (N_4614,N_4469,N_4429);
or U4615 (N_4615,N_4383,N_4409);
and U4616 (N_4616,N_4413,N_4486);
nor U4617 (N_4617,N_4392,N_4455);
or U4618 (N_4618,N_4411,N_4484);
nor U4619 (N_4619,N_4412,N_4377);
xor U4620 (N_4620,N_4435,N_4442);
nand U4621 (N_4621,N_4462,N_4390);
nand U4622 (N_4622,N_4467,N_4376);
nand U4623 (N_4623,N_4421,N_4472);
xnor U4624 (N_4624,N_4448,N_4466);
xor U4625 (N_4625,N_4501,N_4568);
xnor U4626 (N_4626,N_4550,N_4586);
or U4627 (N_4627,N_4575,N_4500);
nand U4628 (N_4628,N_4559,N_4606);
xnor U4629 (N_4629,N_4591,N_4552);
and U4630 (N_4630,N_4565,N_4617);
and U4631 (N_4631,N_4554,N_4517);
or U4632 (N_4632,N_4537,N_4514);
nor U4633 (N_4633,N_4557,N_4508);
or U4634 (N_4634,N_4526,N_4515);
nor U4635 (N_4635,N_4562,N_4595);
or U4636 (N_4636,N_4504,N_4556);
nor U4637 (N_4637,N_4536,N_4603);
nor U4638 (N_4638,N_4602,N_4596);
and U4639 (N_4639,N_4605,N_4566);
or U4640 (N_4640,N_4574,N_4618);
xnor U4641 (N_4641,N_4542,N_4553);
and U4642 (N_4642,N_4611,N_4598);
nand U4643 (N_4643,N_4607,N_4583);
and U4644 (N_4644,N_4569,N_4608);
nand U4645 (N_4645,N_4571,N_4532);
or U4646 (N_4646,N_4581,N_4524);
or U4647 (N_4647,N_4534,N_4590);
xor U4648 (N_4648,N_4582,N_4551);
xnor U4649 (N_4649,N_4572,N_4573);
and U4650 (N_4650,N_4513,N_4547);
or U4651 (N_4651,N_4604,N_4588);
or U4652 (N_4652,N_4587,N_4612);
nor U4653 (N_4653,N_4594,N_4577);
nor U4654 (N_4654,N_4580,N_4599);
or U4655 (N_4655,N_4619,N_4576);
and U4656 (N_4656,N_4522,N_4531);
nor U4657 (N_4657,N_4519,N_4613);
nand U4658 (N_4658,N_4541,N_4540);
and U4659 (N_4659,N_4564,N_4518);
xor U4660 (N_4660,N_4616,N_4530);
nor U4661 (N_4661,N_4506,N_4507);
nor U4662 (N_4662,N_4538,N_4528);
or U4663 (N_4663,N_4610,N_4592);
and U4664 (N_4664,N_4614,N_4543);
nand U4665 (N_4665,N_4589,N_4584);
xor U4666 (N_4666,N_4609,N_4563);
nand U4667 (N_4667,N_4621,N_4597);
and U4668 (N_4668,N_4567,N_4624);
xnor U4669 (N_4669,N_4548,N_4600);
nand U4670 (N_4670,N_4525,N_4579);
xor U4671 (N_4671,N_4511,N_4560);
nor U4672 (N_4672,N_4615,N_4502);
nor U4673 (N_4673,N_4510,N_4622);
nand U4674 (N_4674,N_4516,N_4546);
or U4675 (N_4675,N_4512,N_4539);
and U4676 (N_4676,N_4523,N_4620);
or U4677 (N_4677,N_4623,N_4585);
nand U4678 (N_4678,N_4544,N_4533);
or U4679 (N_4679,N_4549,N_4545);
or U4680 (N_4680,N_4509,N_4561);
xnor U4681 (N_4681,N_4520,N_4529);
nor U4682 (N_4682,N_4527,N_4505);
nor U4683 (N_4683,N_4503,N_4578);
xor U4684 (N_4684,N_4558,N_4601);
or U4685 (N_4685,N_4555,N_4535);
xor U4686 (N_4686,N_4593,N_4521);
xor U4687 (N_4687,N_4570,N_4563);
nand U4688 (N_4688,N_4552,N_4556);
and U4689 (N_4689,N_4557,N_4589);
xor U4690 (N_4690,N_4589,N_4516);
or U4691 (N_4691,N_4596,N_4616);
and U4692 (N_4692,N_4563,N_4550);
xor U4693 (N_4693,N_4502,N_4533);
nor U4694 (N_4694,N_4586,N_4582);
nand U4695 (N_4695,N_4601,N_4532);
or U4696 (N_4696,N_4577,N_4587);
xnor U4697 (N_4697,N_4518,N_4592);
nor U4698 (N_4698,N_4511,N_4621);
xnor U4699 (N_4699,N_4596,N_4543);
nand U4700 (N_4700,N_4603,N_4503);
or U4701 (N_4701,N_4510,N_4573);
and U4702 (N_4702,N_4562,N_4556);
xnor U4703 (N_4703,N_4543,N_4530);
nand U4704 (N_4704,N_4528,N_4610);
nor U4705 (N_4705,N_4558,N_4590);
nor U4706 (N_4706,N_4593,N_4621);
and U4707 (N_4707,N_4580,N_4523);
xnor U4708 (N_4708,N_4521,N_4524);
nand U4709 (N_4709,N_4566,N_4546);
nor U4710 (N_4710,N_4549,N_4602);
and U4711 (N_4711,N_4612,N_4506);
and U4712 (N_4712,N_4510,N_4525);
nand U4713 (N_4713,N_4607,N_4569);
and U4714 (N_4714,N_4544,N_4502);
nand U4715 (N_4715,N_4573,N_4514);
nor U4716 (N_4716,N_4506,N_4611);
xnor U4717 (N_4717,N_4546,N_4602);
and U4718 (N_4718,N_4623,N_4592);
and U4719 (N_4719,N_4524,N_4558);
or U4720 (N_4720,N_4517,N_4510);
nor U4721 (N_4721,N_4559,N_4532);
or U4722 (N_4722,N_4520,N_4558);
and U4723 (N_4723,N_4545,N_4505);
nor U4724 (N_4724,N_4551,N_4561);
and U4725 (N_4725,N_4503,N_4574);
nor U4726 (N_4726,N_4540,N_4533);
and U4727 (N_4727,N_4535,N_4515);
nand U4728 (N_4728,N_4571,N_4614);
and U4729 (N_4729,N_4561,N_4520);
and U4730 (N_4730,N_4622,N_4544);
and U4731 (N_4731,N_4586,N_4538);
xnor U4732 (N_4732,N_4596,N_4547);
nand U4733 (N_4733,N_4617,N_4607);
nor U4734 (N_4734,N_4536,N_4512);
xor U4735 (N_4735,N_4534,N_4505);
nand U4736 (N_4736,N_4608,N_4523);
xnor U4737 (N_4737,N_4546,N_4568);
and U4738 (N_4738,N_4544,N_4540);
nor U4739 (N_4739,N_4545,N_4611);
or U4740 (N_4740,N_4560,N_4619);
nand U4741 (N_4741,N_4580,N_4559);
nor U4742 (N_4742,N_4534,N_4540);
or U4743 (N_4743,N_4589,N_4579);
xor U4744 (N_4744,N_4539,N_4573);
xor U4745 (N_4745,N_4606,N_4615);
nor U4746 (N_4746,N_4591,N_4562);
nand U4747 (N_4747,N_4556,N_4540);
nor U4748 (N_4748,N_4557,N_4539);
or U4749 (N_4749,N_4561,N_4505);
nor U4750 (N_4750,N_4682,N_4703);
nor U4751 (N_4751,N_4637,N_4691);
or U4752 (N_4752,N_4668,N_4671);
or U4753 (N_4753,N_4677,N_4734);
nor U4754 (N_4754,N_4735,N_4655);
or U4755 (N_4755,N_4708,N_4749);
nor U4756 (N_4756,N_4643,N_4736);
and U4757 (N_4757,N_4744,N_4636);
nor U4758 (N_4758,N_4707,N_4665);
nand U4759 (N_4759,N_4747,N_4646);
and U4760 (N_4760,N_4645,N_4698);
nand U4761 (N_4761,N_4712,N_4695);
and U4762 (N_4762,N_4675,N_4648);
nand U4763 (N_4763,N_4697,N_4689);
nor U4764 (N_4764,N_4661,N_4639);
xnor U4765 (N_4765,N_4656,N_4629);
and U4766 (N_4766,N_4638,N_4663);
xor U4767 (N_4767,N_4653,N_4699);
or U4768 (N_4768,N_4716,N_4659);
nor U4769 (N_4769,N_4626,N_4741);
nor U4770 (N_4770,N_4679,N_4654);
xor U4771 (N_4771,N_4630,N_4644);
nor U4772 (N_4772,N_4704,N_4721);
nand U4773 (N_4773,N_4700,N_4714);
xor U4774 (N_4774,N_4633,N_4660);
nor U4775 (N_4775,N_4690,N_4628);
nor U4776 (N_4776,N_4672,N_4715);
or U4777 (N_4777,N_4746,N_4739);
xor U4778 (N_4778,N_4676,N_4625);
nand U4779 (N_4779,N_4693,N_4728);
nand U4780 (N_4780,N_4692,N_4627);
xnor U4781 (N_4781,N_4678,N_4680);
or U4782 (N_4782,N_4702,N_4694);
xor U4783 (N_4783,N_4667,N_4642);
or U4784 (N_4784,N_4685,N_4743);
nand U4785 (N_4785,N_4740,N_4673);
xnor U4786 (N_4786,N_4658,N_4725);
and U4787 (N_4787,N_4657,N_4687);
and U4788 (N_4788,N_4720,N_4650);
nor U4789 (N_4789,N_4641,N_4664);
nor U4790 (N_4790,N_4710,N_4737);
and U4791 (N_4791,N_4666,N_4717);
nand U4792 (N_4792,N_4688,N_4701);
or U4793 (N_4793,N_4669,N_4631);
xor U4794 (N_4794,N_4632,N_4726);
nor U4795 (N_4795,N_4696,N_4651);
or U4796 (N_4796,N_4681,N_4647);
or U4797 (N_4797,N_4686,N_4706);
or U4798 (N_4798,N_4729,N_4748);
xor U4799 (N_4799,N_4732,N_4718);
nand U4800 (N_4800,N_4731,N_4730);
and U4801 (N_4801,N_4711,N_4684);
and U4802 (N_4802,N_4745,N_4674);
nand U4803 (N_4803,N_4723,N_4670);
nand U4804 (N_4804,N_4722,N_4724);
nand U4805 (N_4805,N_4640,N_4738);
nand U4806 (N_4806,N_4652,N_4635);
nand U4807 (N_4807,N_4705,N_4713);
and U4808 (N_4808,N_4742,N_4727);
nand U4809 (N_4809,N_4649,N_4634);
nand U4810 (N_4810,N_4709,N_4662);
xor U4811 (N_4811,N_4683,N_4733);
xor U4812 (N_4812,N_4719,N_4665);
nor U4813 (N_4813,N_4654,N_4705);
nand U4814 (N_4814,N_4747,N_4745);
or U4815 (N_4815,N_4707,N_4651);
nor U4816 (N_4816,N_4658,N_4645);
nor U4817 (N_4817,N_4648,N_4744);
xnor U4818 (N_4818,N_4683,N_4713);
xor U4819 (N_4819,N_4746,N_4648);
or U4820 (N_4820,N_4713,N_4625);
nor U4821 (N_4821,N_4657,N_4706);
or U4822 (N_4822,N_4655,N_4656);
nand U4823 (N_4823,N_4669,N_4704);
nor U4824 (N_4824,N_4645,N_4626);
nand U4825 (N_4825,N_4638,N_4674);
xnor U4826 (N_4826,N_4674,N_4685);
and U4827 (N_4827,N_4636,N_4651);
xnor U4828 (N_4828,N_4737,N_4628);
xor U4829 (N_4829,N_4677,N_4638);
or U4830 (N_4830,N_4672,N_4748);
or U4831 (N_4831,N_4746,N_4696);
xnor U4832 (N_4832,N_4719,N_4695);
nand U4833 (N_4833,N_4664,N_4705);
nor U4834 (N_4834,N_4679,N_4699);
xor U4835 (N_4835,N_4657,N_4704);
xor U4836 (N_4836,N_4707,N_4742);
or U4837 (N_4837,N_4726,N_4684);
nor U4838 (N_4838,N_4713,N_4669);
or U4839 (N_4839,N_4746,N_4689);
nand U4840 (N_4840,N_4643,N_4699);
xnor U4841 (N_4841,N_4648,N_4718);
or U4842 (N_4842,N_4727,N_4628);
or U4843 (N_4843,N_4637,N_4656);
nand U4844 (N_4844,N_4675,N_4678);
xnor U4845 (N_4845,N_4742,N_4732);
nor U4846 (N_4846,N_4649,N_4642);
or U4847 (N_4847,N_4707,N_4686);
or U4848 (N_4848,N_4677,N_4673);
xor U4849 (N_4849,N_4698,N_4650);
nor U4850 (N_4850,N_4650,N_4652);
xor U4851 (N_4851,N_4656,N_4697);
xor U4852 (N_4852,N_4638,N_4705);
or U4853 (N_4853,N_4731,N_4642);
and U4854 (N_4854,N_4705,N_4701);
and U4855 (N_4855,N_4714,N_4704);
nand U4856 (N_4856,N_4646,N_4706);
nor U4857 (N_4857,N_4688,N_4637);
nor U4858 (N_4858,N_4695,N_4702);
xnor U4859 (N_4859,N_4695,N_4694);
nor U4860 (N_4860,N_4644,N_4680);
nand U4861 (N_4861,N_4685,N_4689);
xor U4862 (N_4862,N_4652,N_4640);
or U4863 (N_4863,N_4729,N_4665);
xor U4864 (N_4864,N_4718,N_4666);
nand U4865 (N_4865,N_4727,N_4653);
or U4866 (N_4866,N_4698,N_4704);
nand U4867 (N_4867,N_4649,N_4680);
nor U4868 (N_4868,N_4676,N_4651);
nand U4869 (N_4869,N_4722,N_4663);
xor U4870 (N_4870,N_4718,N_4714);
or U4871 (N_4871,N_4740,N_4678);
or U4872 (N_4872,N_4705,N_4656);
and U4873 (N_4873,N_4688,N_4748);
and U4874 (N_4874,N_4668,N_4737);
and U4875 (N_4875,N_4851,N_4827);
and U4876 (N_4876,N_4774,N_4788);
xor U4877 (N_4877,N_4840,N_4803);
xor U4878 (N_4878,N_4819,N_4753);
or U4879 (N_4879,N_4814,N_4842);
or U4880 (N_4880,N_4815,N_4785);
nor U4881 (N_4881,N_4800,N_4775);
xnor U4882 (N_4882,N_4861,N_4850);
xor U4883 (N_4883,N_4873,N_4829);
nand U4884 (N_4884,N_4763,N_4764);
and U4885 (N_4885,N_4762,N_4857);
or U4886 (N_4886,N_4822,N_4801);
xnor U4887 (N_4887,N_4810,N_4849);
and U4888 (N_4888,N_4852,N_4824);
nand U4889 (N_4889,N_4848,N_4821);
nand U4890 (N_4890,N_4863,N_4812);
xor U4891 (N_4891,N_4767,N_4798);
nand U4892 (N_4892,N_4807,N_4792);
nor U4893 (N_4893,N_4765,N_4776);
xnor U4894 (N_4894,N_4811,N_4772);
nand U4895 (N_4895,N_4825,N_4846);
or U4896 (N_4896,N_4797,N_4791);
nand U4897 (N_4897,N_4833,N_4828);
or U4898 (N_4898,N_4808,N_4855);
xnor U4899 (N_4899,N_4860,N_4778);
or U4900 (N_4900,N_4799,N_4847);
or U4901 (N_4901,N_4862,N_4780);
and U4902 (N_4902,N_4750,N_4816);
or U4903 (N_4903,N_4813,N_4872);
or U4904 (N_4904,N_4769,N_4871);
or U4905 (N_4905,N_4856,N_4820);
nand U4906 (N_4906,N_4838,N_4826);
or U4907 (N_4907,N_4874,N_4836);
or U4908 (N_4908,N_4802,N_4817);
and U4909 (N_4909,N_4845,N_4841);
nand U4910 (N_4910,N_4866,N_4787);
xnor U4911 (N_4911,N_4834,N_4752);
nand U4912 (N_4912,N_4756,N_4773);
nand U4913 (N_4913,N_4781,N_4751);
nor U4914 (N_4914,N_4794,N_4831);
or U4915 (N_4915,N_4809,N_4823);
xnor U4916 (N_4916,N_4771,N_4790);
xor U4917 (N_4917,N_4870,N_4830);
nand U4918 (N_4918,N_4760,N_4844);
or U4919 (N_4919,N_4754,N_4868);
nand U4920 (N_4920,N_4786,N_4843);
xor U4921 (N_4921,N_4835,N_4784);
or U4922 (N_4922,N_4869,N_4837);
or U4923 (N_4923,N_4779,N_4806);
or U4924 (N_4924,N_4839,N_4777);
nor U4925 (N_4925,N_4796,N_4805);
and U4926 (N_4926,N_4854,N_4864);
nand U4927 (N_4927,N_4758,N_4782);
nor U4928 (N_4928,N_4793,N_4795);
and U4929 (N_4929,N_4865,N_4761);
nor U4930 (N_4930,N_4804,N_4770);
nor U4931 (N_4931,N_4832,N_4759);
and U4932 (N_4932,N_4867,N_4768);
nand U4933 (N_4933,N_4789,N_4858);
nor U4934 (N_4934,N_4757,N_4766);
and U4935 (N_4935,N_4783,N_4859);
or U4936 (N_4936,N_4853,N_4755);
xor U4937 (N_4937,N_4818,N_4814);
or U4938 (N_4938,N_4807,N_4847);
nor U4939 (N_4939,N_4873,N_4781);
xnor U4940 (N_4940,N_4823,N_4785);
or U4941 (N_4941,N_4850,N_4789);
or U4942 (N_4942,N_4771,N_4782);
and U4943 (N_4943,N_4786,N_4784);
xnor U4944 (N_4944,N_4855,N_4799);
and U4945 (N_4945,N_4830,N_4761);
xnor U4946 (N_4946,N_4831,N_4841);
or U4947 (N_4947,N_4860,N_4850);
and U4948 (N_4948,N_4822,N_4873);
nor U4949 (N_4949,N_4808,N_4798);
nor U4950 (N_4950,N_4767,N_4872);
nand U4951 (N_4951,N_4828,N_4791);
nand U4952 (N_4952,N_4835,N_4768);
and U4953 (N_4953,N_4861,N_4860);
xor U4954 (N_4954,N_4796,N_4785);
or U4955 (N_4955,N_4871,N_4763);
xor U4956 (N_4956,N_4852,N_4870);
nand U4957 (N_4957,N_4823,N_4835);
nand U4958 (N_4958,N_4855,N_4835);
and U4959 (N_4959,N_4775,N_4856);
and U4960 (N_4960,N_4803,N_4856);
xnor U4961 (N_4961,N_4846,N_4774);
nor U4962 (N_4962,N_4785,N_4873);
and U4963 (N_4963,N_4829,N_4867);
and U4964 (N_4964,N_4802,N_4754);
xor U4965 (N_4965,N_4762,N_4816);
and U4966 (N_4966,N_4789,N_4843);
and U4967 (N_4967,N_4803,N_4804);
and U4968 (N_4968,N_4820,N_4848);
xnor U4969 (N_4969,N_4823,N_4763);
nor U4970 (N_4970,N_4754,N_4842);
nor U4971 (N_4971,N_4802,N_4871);
or U4972 (N_4972,N_4870,N_4780);
nor U4973 (N_4973,N_4757,N_4753);
nor U4974 (N_4974,N_4849,N_4817);
nor U4975 (N_4975,N_4848,N_4777);
nand U4976 (N_4976,N_4782,N_4853);
or U4977 (N_4977,N_4768,N_4788);
xnor U4978 (N_4978,N_4806,N_4819);
and U4979 (N_4979,N_4853,N_4846);
and U4980 (N_4980,N_4807,N_4872);
and U4981 (N_4981,N_4843,N_4869);
nor U4982 (N_4982,N_4781,N_4812);
nor U4983 (N_4983,N_4776,N_4865);
xnor U4984 (N_4984,N_4778,N_4840);
and U4985 (N_4985,N_4870,N_4849);
and U4986 (N_4986,N_4854,N_4801);
nand U4987 (N_4987,N_4865,N_4775);
xnor U4988 (N_4988,N_4871,N_4762);
and U4989 (N_4989,N_4866,N_4752);
nor U4990 (N_4990,N_4761,N_4789);
xnor U4991 (N_4991,N_4784,N_4826);
nor U4992 (N_4992,N_4755,N_4859);
xor U4993 (N_4993,N_4841,N_4785);
and U4994 (N_4994,N_4788,N_4812);
nand U4995 (N_4995,N_4860,N_4847);
xor U4996 (N_4996,N_4830,N_4787);
xnor U4997 (N_4997,N_4785,N_4842);
xnor U4998 (N_4998,N_4783,N_4844);
xnor U4999 (N_4999,N_4845,N_4751);
nand U5000 (N_5000,N_4877,N_4897);
xnor U5001 (N_5001,N_4925,N_4984);
or U5002 (N_5002,N_4923,N_4883);
or U5003 (N_5003,N_4888,N_4992);
or U5004 (N_5004,N_4898,N_4902);
nand U5005 (N_5005,N_4971,N_4931);
or U5006 (N_5006,N_4977,N_4903);
nand U5007 (N_5007,N_4935,N_4882);
or U5008 (N_5008,N_4907,N_4928);
nand U5009 (N_5009,N_4948,N_4937);
nand U5010 (N_5010,N_4890,N_4885);
nand U5011 (N_5011,N_4952,N_4983);
and U5012 (N_5012,N_4924,N_4959);
or U5013 (N_5013,N_4887,N_4965);
nor U5014 (N_5014,N_4997,N_4884);
nand U5015 (N_5015,N_4975,N_4981);
or U5016 (N_5016,N_4974,N_4960);
or U5017 (N_5017,N_4916,N_4879);
or U5018 (N_5018,N_4964,N_4911);
nor U5019 (N_5019,N_4982,N_4987);
nor U5020 (N_5020,N_4973,N_4993);
nand U5021 (N_5021,N_4893,N_4979);
and U5022 (N_5022,N_4966,N_4895);
and U5023 (N_5023,N_4968,N_4875);
xnor U5024 (N_5024,N_4953,N_4936);
and U5025 (N_5025,N_4989,N_4891);
xnor U5026 (N_5026,N_4990,N_4942);
or U5027 (N_5027,N_4900,N_4967);
xor U5028 (N_5028,N_4958,N_4886);
nand U5029 (N_5029,N_4932,N_4951);
and U5030 (N_5030,N_4929,N_4878);
nor U5031 (N_5031,N_4947,N_4991);
and U5032 (N_5032,N_4956,N_4933);
xor U5033 (N_5033,N_4892,N_4912);
nand U5034 (N_5034,N_4944,N_4921);
nor U5035 (N_5035,N_4941,N_4998);
and U5036 (N_5036,N_4943,N_4908);
nand U5037 (N_5037,N_4939,N_4896);
nand U5038 (N_5038,N_4876,N_4986);
and U5039 (N_5039,N_4949,N_4978);
or U5040 (N_5040,N_4957,N_4918);
nor U5041 (N_5041,N_4976,N_4920);
xor U5042 (N_5042,N_4940,N_4963);
nand U5043 (N_5043,N_4927,N_4919);
xor U5044 (N_5044,N_4910,N_4985);
and U5045 (N_5045,N_4906,N_4938);
and U5046 (N_5046,N_4934,N_4914);
xnor U5047 (N_5047,N_4889,N_4962);
and U5048 (N_5048,N_4904,N_4917);
nor U5049 (N_5049,N_4930,N_4995);
nand U5050 (N_5050,N_4961,N_4915);
or U5051 (N_5051,N_4980,N_4881);
or U5052 (N_5052,N_4909,N_4954);
nor U5053 (N_5053,N_4894,N_4946);
and U5054 (N_5054,N_4969,N_4899);
xor U5055 (N_5055,N_4996,N_4922);
nor U5056 (N_5056,N_4880,N_4994);
and U5057 (N_5057,N_4945,N_4926);
nand U5058 (N_5058,N_4905,N_4988);
xnor U5059 (N_5059,N_4970,N_4913);
xor U5060 (N_5060,N_4955,N_4950);
xnor U5061 (N_5061,N_4901,N_4972);
nand U5062 (N_5062,N_4999,N_4901);
and U5063 (N_5063,N_4896,N_4919);
nand U5064 (N_5064,N_4904,N_4963);
nand U5065 (N_5065,N_4950,N_4948);
nor U5066 (N_5066,N_4956,N_4989);
nor U5067 (N_5067,N_4968,N_4964);
xnor U5068 (N_5068,N_4907,N_4940);
or U5069 (N_5069,N_4924,N_4925);
nand U5070 (N_5070,N_4882,N_4984);
or U5071 (N_5071,N_4880,N_4898);
and U5072 (N_5072,N_4968,N_4990);
nor U5073 (N_5073,N_4926,N_4881);
nor U5074 (N_5074,N_4899,N_4877);
or U5075 (N_5075,N_4907,N_4892);
nor U5076 (N_5076,N_4892,N_4897);
nand U5077 (N_5077,N_4949,N_4934);
nor U5078 (N_5078,N_4985,N_4995);
nand U5079 (N_5079,N_4993,N_4880);
or U5080 (N_5080,N_4895,N_4925);
and U5081 (N_5081,N_4904,N_4926);
or U5082 (N_5082,N_4882,N_4915);
xnor U5083 (N_5083,N_4947,N_4887);
or U5084 (N_5084,N_4949,N_4882);
nor U5085 (N_5085,N_4910,N_4893);
and U5086 (N_5086,N_4974,N_4977);
or U5087 (N_5087,N_4939,N_4920);
and U5088 (N_5088,N_4890,N_4980);
or U5089 (N_5089,N_4946,N_4991);
nor U5090 (N_5090,N_4941,N_4952);
nor U5091 (N_5091,N_4970,N_4877);
xnor U5092 (N_5092,N_4986,N_4962);
nor U5093 (N_5093,N_4903,N_4902);
nor U5094 (N_5094,N_4991,N_4956);
xnor U5095 (N_5095,N_4880,N_4912);
nand U5096 (N_5096,N_4891,N_4901);
or U5097 (N_5097,N_4917,N_4933);
or U5098 (N_5098,N_4918,N_4891);
nor U5099 (N_5099,N_4905,N_4906);
nand U5100 (N_5100,N_4981,N_4998);
nor U5101 (N_5101,N_4899,N_4932);
nor U5102 (N_5102,N_4899,N_4960);
nand U5103 (N_5103,N_4901,N_4882);
nand U5104 (N_5104,N_4902,N_4967);
or U5105 (N_5105,N_4920,N_4899);
nand U5106 (N_5106,N_4969,N_4972);
or U5107 (N_5107,N_4970,N_4992);
nor U5108 (N_5108,N_4879,N_4990);
xnor U5109 (N_5109,N_4908,N_4991);
and U5110 (N_5110,N_4962,N_4967);
nor U5111 (N_5111,N_4925,N_4953);
and U5112 (N_5112,N_4964,N_4884);
and U5113 (N_5113,N_4955,N_4929);
nor U5114 (N_5114,N_4893,N_4897);
nor U5115 (N_5115,N_4875,N_4946);
nor U5116 (N_5116,N_4965,N_4915);
and U5117 (N_5117,N_4936,N_4949);
or U5118 (N_5118,N_4988,N_4969);
nor U5119 (N_5119,N_4880,N_4970);
nand U5120 (N_5120,N_4976,N_4911);
nand U5121 (N_5121,N_4945,N_4929);
nor U5122 (N_5122,N_4883,N_4943);
or U5123 (N_5123,N_4905,N_4946);
nor U5124 (N_5124,N_4878,N_4920);
nor U5125 (N_5125,N_5123,N_5115);
xnor U5126 (N_5126,N_5060,N_5032);
nor U5127 (N_5127,N_5086,N_5111);
nor U5128 (N_5128,N_5096,N_5108);
nand U5129 (N_5129,N_5001,N_5026);
nand U5130 (N_5130,N_5062,N_5121);
nand U5131 (N_5131,N_5065,N_5112);
nand U5132 (N_5132,N_5047,N_5028);
or U5133 (N_5133,N_5052,N_5013);
nor U5134 (N_5134,N_5041,N_5030);
and U5135 (N_5135,N_5092,N_5005);
nor U5136 (N_5136,N_5098,N_5011);
nand U5137 (N_5137,N_5116,N_5007);
or U5138 (N_5138,N_5019,N_5072);
nand U5139 (N_5139,N_5002,N_5034);
xor U5140 (N_5140,N_5027,N_5021);
and U5141 (N_5141,N_5094,N_5006);
nand U5142 (N_5142,N_5104,N_5122);
nand U5143 (N_5143,N_5120,N_5050);
and U5144 (N_5144,N_5084,N_5015);
or U5145 (N_5145,N_5054,N_5033);
xor U5146 (N_5146,N_5114,N_5066);
nor U5147 (N_5147,N_5024,N_5073);
nor U5148 (N_5148,N_5075,N_5100);
nor U5149 (N_5149,N_5010,N_5124);
nand U5150 (N_5150,N_5035,N_5067);
or U5151 (N_5151,N_5089,N_5105);
xnor U5152 (N_5152,N_5099,N_5031);
and U5153 (N_5153,N_5048,N_5078);
or U5154 (N_5154,N_5009,N_5082);
or U5155 (N_5155,N_5017,N_5076);
and U5156 (N_5156,N_5046,N_5036);
nor U5157 (N_5157,N_5091,N_5040);
and U5158 (N_5158,N_5064,N_5087);
nor U5159 (N_5159,N_5095,N_5042);
and U5160 (N_5160,N_5055,N_5012);
nor U5161 (N_5161,N_5083,N_5109);
nand U5162 (N_5162,N_5057,N_5063);
xnor U5163 (N_5163,N_5008,N_5077);
xor U5164 (N_5164,N_5049,N_5093);
or U5165 (N_5165,N_5029,N_5039);
and U5166 (N_5166,N_5119,N_5107);
nor U5167 (N_5167,N_5102,N_5043);
xor U5168 (N_5168,N_5061,N_5059);
xnor U5169 (N_5169,N_5088,N_5003);
or U5170 (N_5170,N_5038,N_5113);
xnor U5171 (N_5171,N_5020,N_5079);
nand U5172 (N_5172,N_5045,N_5110);
nor U5173 (N_5173,N_5058,N_5117);
and U5174 (N_5174,N_5068,N_5070);
and U5175 (N_5175,N_5000,N_5071);
or U5176 (N_5176,N_5069,N_5025);
nor U5177 (N_5177,N_5081,N_5022);
or U5178 (N_5178,N_5080,N_5051);
or U5179 (N_5179,N_5023,N_5103);
and U5180 (N_5180,N_5118,N_5004);
xor U5181 (N_5181,N_5074,N_5014);
or U5182 (N_5182,N_5106,N_5016);
or U5183 (N_5183,N_5056,N_5053);
nor U5184 (N_5184,N_5090,N_5085);
nor U5185 (N_5185,N_5097,N_5018);
xor U5186 (N_5186,N_5044,N_5037);
nand U5187 (N_5187,N_5101,N_5115);
nor U5188 (N_5188,N_5080,N_5120);
or U5189 (N_5189,N_5027,N_5014);
and U5190 (N_5190,N_5090,N_5107);
and U5191 (N_5191,N_5119,N_5116);
nor U5192 (N_5192,N_5031,N_5061);
xnor U5193 (N_5193,N_5034,N_5116);
xor U5194 (N_5194,N_5115,N_5023);
nor U5195 (N_5195,N_5046,N_5007);
xor U5196 (N_5196,N_5013,N_5099);
nor U5197 (N_5197,N_5081,N_5010);
or U5198 (N_5198,N_5044,N_5049);
and U5199 (N_5199,N_5031,N_5084);
nand U5200 (N_5200,N_5079,N_5001);
nand U5201 (N_5201,N_5028,N_5114);
xor U5202 (N_5202,N_5092,N_5065);
and U5203 (N_5203,N_5016,N_5060);
or U5204 (N_5204,N_5102,N_5065);
nand U5205 (N_5205,N_5052,N_5016);
or U5206 (N_5206,N_5011,N_5026);
nor U5207 (N_5207,N_5120,N_5025);
or U5208 (N_5208,N_5006,N_5007);
nor U5209 (N_5209,N_5025,N_5040);
xor U5210 (N_5210,N_5060,N_5081);
and U5211 (N_5211,N_5046,N_5100);
xor U5212 (N_5212,N_5061,N_5091);
nand U5213 (N_5213,N_5086,N_5007);
and U5214 (N_5214,N_5040,N_5121);
nor U5215 (N_5215,N_5020,N_5052);
nor U5216 (N_5216,N_5101,N_5015);
xnor U5217 (N_5217,N_5059,N_5104);
xor U5218 (N_5218,N_5123,N_5029);
and U5219 (N_5219,N_5007,N_5009);
nor U5220 (N_5220,N_5043,N_5114);
xnor U5221 (N_5221,N_5116,N_5072);
nand U5222 (N_5222,N_5072,N_5074);
or U5223 (N_5223,N_5087,N_5008);
and U5224 (N_5224,N_5003,N_5083);
xor U5225 (N_5225,N_5018,N_5099);
nand U5226 (N_5226,N_5094,N_5062);
xnor U5227 (N_5227,N_5006,N_5037);
and U5228 (N_5228,N_5081,N_5106);
xor U5229 (N_5229,N_5106,N_5072);
nand U5230 (N_5230,N_5009,N_5036);
or U5231 (N_5231,N_5045,N_5119);
xor U5232 (N_5232,N_5092,N_5121);
nand U5233 (N_5233,N_5094,N_5099);
xor U5234 (N_5234,N_5109,N_5055);
and U5235 (N_5235,N_5050,N_5058);
or U5236 (N_5236,N_5032,N_5063);
nand U5237 (N_5237,N_5105,N_5009);
xnor U5238 (N_5238,N_5039,N_5098);
nand U5239 (N_5239,N_5115,N_5056);
nand U5240 (N_5240,N_5096,N_5030);
nor U5241 (N_5241,N_5114,N_5115);
nor U5242 (N_5242,N_5040,N_5050);
nand U5243 (N_5243,N_5045,N_5075);
or U5244 (N_5244,N_5029,N_5064);
xor U5245 (N_5245,N_5090,N_5054);
and U5246 (N_5246,N_5097,N_5014);
and U5247 (N_5247,N_5024,N_5110);
nand U5248 (N_5248,N_5006,N_5017);
and U5249 (N_5249,N_5098,N_5048);
nand U5250 (N_5250,N_5139,N_5206);
nor U5251 (N_5251,N_5165,N_5181);
and U5252 (N_5252,N_5177,N_5130);
xnor U5253 (N_5253,N_5126,N_5207);
and U5254 (N_5254,N_5217,N_5228);
nand U5255 (N_5255,N_5147,N_5218);
and U5256 (N_5256,N_5168,N_5223);
nand U5257 (N_5257,N_5247,N_5162);
nand U5258 (N_5258,N_5140,N_5166);
nor U5259 (N_5259,N_5174,N_5176);
nand U5260 (N_5260,N_5195,N_5208);
xnor U5261 (N_5261,N_5155,N_5158);
and U5262 (N_5262,N_5203,N_5154);
and U5263 (N_5263,N_5143,N_5136);
and U5264 (N_5264,N_5238,N_5185);
xor U5265 (N_5265,N_5156,N_5201);
nand U5266 (N_5266,N_5157,N_5241);
nor U5267 (N_5267,N_5222,N_5146);
xnor U5268 (N_5268,N_5202,N_5213);
or U5269 (N_5269,N_5173,N_5171);
nand U5270 (N_5270,N_5245,N_5179);
xnor U5271 (N_5271,N_5200,N_5129);
xnor U5272 (N_5272,N_5133,N_5233);
nor U5273 (N_5273,N_5239,N_5209);
nor U5274 (N_5274,N_5234,N_5175);
and U5275 (N_5275,N_5249,N_5199);
and U5276 (N_5276,N_5125,N_5127);
xor U5277 (N_5277,N_5230,N_5248);
nand U5278 (N_5278,N_5167,N_5193);
xor U5279 (N_5279,N_5150,N_5178);
xnor U5280 (N_5280,N_5191,N_5145);
nor U5281 (N_5281,N_5132,N_5216);
xor U5282 (N_5282,N_5151,N_5159);
xor U5283 (N_5283,N_5225,N_5212);
nor U5284 (N_5284,N_5231,N_5197);
nand U5285 (N_5285,N_5192,N_5220);
and U5286 (N_5286,N_5153,N_5190);
nand U5287 (N_5287,N_5204,N_5142);
nor U5288 (N_5288,N_5164,N_5131);
xnor U5289 (N_5289,N_5135,N_5243);
and U5290 (N_5290,N_5205,N_5227);
or U5291 (N_5291,N_5138,N_5184);
nor U5292 (N_5292,N_5219,N_5137);
nand U5293 (N_5293,N_5246,N_5186);
nor U5294 (N_5294,N_5163,N_5180);
nor U5295 (N_5295,N_5214,N_5221);
xor U5296 (N_5296,N_5187,N_5141);
or U5297 (N_5297,N_5215,N_5128);
nand U5298 (N_5298,N_5149,N_5183);
or U5299 (N_5299,N_5240,N_5148);
xor U5300 (N_5300,N_5196,N_5236);
nand U5301 (N_5301,N_5169,N_5189);
xor U5302 (N_5302,N_5144,N_5194);
xnor U5303 (N_5303,N_5235,N_5170);
xnor U5304 (N_5304,N_5244,N_5152);
or U5305 (N_5305,N_5237,N_5182);
xnor U5306 (N_5306,N_5188,N_5226);
and U5307 (N_5307,N_5172,N_5211);
xnor U5308 (N_5308,N_5160,N_5134);
xor U5309 (N_5309,N_5210,N_5229);
or U5310 (N_5310,N_5161,N_5224);
xnor U5311 (N_5311,N_5242,N_5232);
nor U5312 (N_5312,N_5198,N_5132);
or U5313 (N_5313,N_5200,N_5154);
xnor U5314 (N_5314,N_5225,N_5164);
and U5315 (N_5315,N_5234,N_5224);
xor U5316 (N_5316,N_5213,N_5204);
nand U5317 (N_5317,N_5169,N_5190);
or U5318 (N_5318,N_5219,N_5160);
nand U5319 (N_5319,N_5166,N_5206);
nand U5320 (N_5320,N_5164,N_5216);
and U5321 (N_5321,N_5190,N_5230);
and U5322 (N_5322,N_5242,N_5167);
nor U5323 (N_5323,N_5175,N_5191);
nand U5324 (N_5324,N_5130,N_5200);
xor U5325 (N_5325,N_5244,N_5133);
or U5326 (N_5326,N_5176,N_5168);
and U5327 (N_5327,N_5192,N_5191);
nand U5328 (N_5328,N_5219,N_5136);
and U5329 (N_5329,N_5125,N_5243);
or U5330 (N_5330,N_5209,N_5236);
xnor U5331 (N_5331,N_5187,N_5142);
or U5332 (N_5332,N_5214,N_5136);
nor U5333 (N_5333,N_5213,N_5165);
nor U5334 (N_5334,N_5184,N_5197);
nand U5335 (N_5335,N_5181,N_5141);
nand U5336 (N_5336,N_5231,N_5240);
nand U5337 (N_5337,N_5154,N_5234);
and U5338 (N_5338,N_5231,N_5189);
xor U5339 (N_5339,N_5139,N_5186);
or U5340 (N_5340,N_5171,N_5181);
nor U5341 (N_5341,N_5200,N_5196);
nor U5342 (N_5342,N_5143,N_5126);
nor U5343 (N_5343,N_5214,N_5206);
xor U5344 (N_5344,N_5133,N_5220);
nand U5345 (N_5345,N_5165,N_5154);
nand U5346 (N_5346,N_5218,N_5133);
and U5347 (N_5347,N_5148,N_5182);
nor U5348 (N_5348,N_5215,N_5136);
nand U5349 (N_5349,N_5199,N_5139);
xor U5350 (N_5350,N_5163,N_5152);
and U5351 (N_5351,N_5212,N_5204);
or U5352 (N_5352,N_5126,N_5228);
nor U5353 (N_5353,N_5207,N_5232);
nand U5354 (N_5354,N_5162,N_5154);
xnor U5355 (N_5355,N_5161,N_5246);
or U5356 (N_5356,N_5181,N_5186);
and U5357 (N_5357,N_5151,N_5209);
xnor U5358 (N_5358,N_5181,N_5206);
xor U5359 (N_5359,N_5207,N_5138);
or U5360 (N_5360,N_5129,N_5233);
nor U5361 (N_5361,N_5184,N_5146);
nand U5362 (N_5362,N_5210,N_5167);
nor U5363 (N_5363,N_5145,N_5207);
xor U5364 (N_5364,N_5229,N_5223);
nand U5365 (N_5365,N_5248,N_5128);
nand U5366 (N_5366,N_5247,N_5165);
and U5367 (N_5367,N_5241,N_5156);
or U5368 (N_5368,N_5167,N_5199);
and U5369 (N_5369,N_5165,N_5150);
nand U5370 (N_5370,N_5182,N_5169);
and U5371 (N_5371,N_5200,N_5222);
or U5372 (N_5372,N_5148,N_5210);
or U5373 (N_5373,N_5231,N_5246);
nand U5374 (N_5374,N_5189,N_5248);
or U5375 (N_5375,N_5302,N_5260);
nor U5376 (N_5376,N_5289,N_5354);
or U5377 (N_5377,N_5374,N_5339);
xor U5378 (N_5378,N_5251,N_5373);
and U5379 (N_5379,N_5352,N_5299);
and U5380 (N_5380,N_5256,N_5361);
xnor U5381 (N_5381,N_5275,N_5318);
nor U5382 (N_5382,N_5346,N_5314);
and U5383 (N_5383,N_5348,N_5283);
xor U5384 (N_5384,N_5284,N_5295);
nor U5385 (N_5385,N_5291,N_5257);
xor U5386 (N_5386,N_5313,N_5349);
or U5387 (N_5387,N_5356,N_5266);
and U5388 (N_5388,N_5368,N_5350);
or U5389 (N_5389,N_5369,N_5370);
nand U5390 (N_5390,N_5269,N_5277);
or U5391 (N_5391,N_5296,N_5357);
or U5392 (N_5392,N_5290,N_5322);
nor U5393 (N_5393,N_5324,N_5273);
and U5394 (N_5394,N_5268,N_5315);
nor U5395 (N_5395,N_5303,N_5336);
xnor U5396 (N_5396,N_5316,N_5331);
xnor U5397 (N_5397,N_5319,N_5308);
nor U5398 (N_5398,N_5367,N_5371);
nor U5399 (N_5399,N_5335,N_5334);
nor U5400 (N_5400,N_5263,N_5342);
nor U5401 (N_5401,N_5366,N_5355);
nor U5402 (N_5402,N_5250,N_5294);
or U5403 (N_5403,N_5292,N_5287);
nand U5404 (N_5404,N_5285,N_5329);
or U5405 (N_5405,N_5317,N_5310);
nor U5406 (N_5406,N_5281,N_5353);
and U5407 (N_5407,N_5305,N_5365);
nor U5408 (N_5408,N_5282,N_5307);
nand U5409 (N_5409,N_5343,N_5255);
xor U5410 (N_5410,N_5274,N_5372);
xor U5411 (N_5411,N_5300,N_5330);
nand U5412 (N_5412,N_5279,N_5262);
and U5413 (N_5413,N_5293,N_5271);
or U5414 (N_5414,N_5345,N_5332);
nand U5415 (N_5415,N_5301,N_5298);
and U5416 (N_5416,N_5264,N_5278);
xor U5417 (N_5417,N_5267,N_5323);
or U5418 (N_5418,N_5362,N_5259);
nor U5419 (N_5419,N_5304,N_5261);
nand U5420 (N_5420,N_5333,N_5320);
and U5421 (N_5421,N_5270,N_5272);
nor U5422 (N_5422,N_5312,N_5258);
nand U5423 (N_5423,N_5364,N_5351);
nand U5424 (N_5424,N_5359,N_5344);
nor U5425 (N_5425,N_5280,N_5309);
and U5426 (N_5426,N_5286,N_5337);
nand U5427 (N_5427,N_5297,N_5325);
nand U5428 (N_5428,N_5252,N_5265);
or U5429 (N_5429,N_5321,N_5288);
nor U5430 (N_5430,N_5338,N_5276);
nand U5431 (N_5431,N_5358,N_5363);
and U5432 (N_5432,N_5360,N_5254);
nand U5433 (N_5433,N_5341,N_5327);
nand U5434 (N_5434,N_5306,N_5328);
nor U5435 (N_5435,N_5347,N_5340);
nand U5436 (N_5436,N_5253,N_5311);
or U5437 (N_5437,N_5326,N_5352);
or U5438 (N_5438,N_5358,N_5312);
and U5439 (N_5439,N_5341,N_5340);
nand U5440 (N_5440,N_5319,N_5317);
nand U5441 (N_5441,N_5266,N_5334);
xor U5442 (N_5442,N_5314,N_5323);
nand U5443 (N_5443,N_5311,N_5346);
xnor U5444 (N_5444,N_5345,N_5365);
and U5445 (N_5445,N_5308,N_5288);
nand U5446 (N_5446,N_5372,N_5320);
and U5447 (N_5447,N_5344,N_5294);
nor U5448 (N_5448,N_5335,N_5310);
nor U5449 (N_5449,N_5295,N_5368);
nor U5450 (N_5450,N_5258,N_5309);
and U5451 (N_5451,N_5326,N_5309);
or U5452 (N_5452,N_5283,N_5285);
xor U5453 (N_5453,N_5344,N_5258);
and U5454 (N_5454,N_5319,N_5366);
xnor U5455 (N_5455,N_5301,N_5338);
xor U5456 (N_5456,N_5345,N_5272);
nand U5457 (N_5457,N_5341,N_5294);
or U5458 (N_5458,N_5286,N_5332);
xnor U5459 (N_5459,N_5323,N_5256);
nand U5460 (N_5460,N_5357,N_5274);
nand U5461 (N_5461,N_5300,N_5342);
nor U5462 (N_5462,N_5303,N_5276);
and U5463 (N_5463,N_5301,N_5331);
and U5464 (N_5464,N_5335,N_5258);
nor U5465 (N_5465,N_5264,N_5357);
nand U5466 (N_5466,N_5369,N_5262);
and U5467 (N_5467,N_5314,N_5287);
nor U5468 (N_5468,N_5293,N_5275);
nor U5469 (N_5469,N_5287,N_5336);
nor U5470 (N_5470,N_5326,N_5287);
and U5471 (N_5471,N_5263,N_5356);
and U5472 (N_5472,N_5350,N_5347);
nand U5473 (N_5473,N_5299,N_5367);
nor U5474 (N_5474,N_5282,N_5354);
or U5475 (N_5475,N_5366,N_5320);
and U5476 (N_5476,N_5264,N_5292);
nand U5477 (N_5477,N_5265,N_5277);
xor U5478 (N_5478,N_5333,N_5359);
nand U5479 (N_5479,N_5325,N_5269);
and U5480 (N_5480,N_5296,N_5271);
nand U5481 (N_5481,N_5266,N_5255);
nor U5482 (N_5482,N_5277,N_5301);
and U5483 (N_5483,N_5302,N_5369);
and U5484 (N_5484,N_5321,N_5260);
nor U5485 (N_5485,N_5354,N_5262);
or U5486 (N_5486,N_5353,N_5344);
nor U5487 (N_5487,N_5296,N_5343);
nand U5488 (N_5488,N_5347,N_5330);
or U5489 (N_5489,N_5284,N_5302);
nand U5490 (N_5490,N_5309,N_5331);
nor U5491 (N_5491,N_5369,N_5354);
and U5492 (N_5492,N_5356,N_5338);
and U5493 (N_5493,N_5269,N_5349);
and U5494 (N_5494,N_5334,N_5316);
nand U5495 (N_5495,N_5351,N_5255);
and U5496 (N_5496,N_5291,N_5337);
or U5497 (N_5497,N_5331,N_5361);
nor U5498 (N_5498,N_5347,N_5296);
and U5499 (N_5499,N_5321,N_5304);
nor U5500 (N_5500,N_5409,N_5442);
nand U5501 (N_5501,N_5479,N_5408);
or U5502 (N_5502,N_5395,N_5434);
nand U5503 (N_5503,N_5407,N_5485);
nor U5504 (N_5504,N_5424,N_5461);
or U5505 (N_5505,N_5383,N_5435);
and U5506 (N_5506,N_5417,N_5437);
xnor U5507 (N_5507,N_5470,N_5441);
nor U5508 (N_5508,N_5410,N_5484);
and U5509 (N_5509,N_5454,N_5448);
xor U5510 (N_5510,N_5480,N_5444);
nand U5511 (N_5511,N_5481,N_5459);
nand U5512 (N_5512,N_5384,N_5419);
xnor U5513 (N_5513,N_5376,N_5496);
nand U5514 (N_5514,N_5426,N_5457);
or U5515 (N_5515,N_5396,N_5456);
nor U5516 (N_5516,N_5446,N_5406);
xnor U5517 (N_5517,N_5433,N_5398);
or U5518 (N_5518,N_5497,N_5445);
or U5519 (N_5519,N_5411,N_5385);
or U5520 (N_5520,N_5449,N_5400);
or U5521 (N_5521,N_5468,N_5462);
and U5522 (N_5522,N_5450,N_5438);
nand U5523 (N_5523,N_5390,N_5403);
or U5524 (N_5524,N_5402,N_5483);
or U5525 (N_5525,N_5386,N_5405);
nand U5526 (N_5526,N_5381,N_5425);
nor U5527 (N_5527,N_5393,N_5375);
or U5528 (N_5528,N_5498,N_5465);
or U5529 (N_5529,N_5472,N_5377);
nor U5530 (N_5530,N_5487,N_5432);
xor U5531 (N_5531,N_5436,N_5430);
and U5532 (N_5532,N_5399,N_5451);
nand U5533 (N_5533,N_5413,N_5466);
nand U5534 (N_5534,N_5471,N_5475);
nand U5535 (N_5535,N_5490,N_5420);
and U5536 (N_5536,N_5412,N_5421);
or U5537 (N_5537,N_5478,N_5404);
and U5538 (N_5538,N_5427,N_5431);
nor U5539 (N_5539,N_5486,N_5476);
xnor U5540 (N_5540,N_5423,N_5452);
or U5541 (N_5541,N_5401,N_5418);
nand U5542 (N_5542,N_5474,N_5387);
or U5543 (N_5543,N_5397,N_5440);
xnor U5544 (N_5544,N_5382,N_5464);
xnor U5545 (N_5545,N_5499,N_5495);
xnor U5546 (N_5546,N_5379,N_5380);
nor U5547 (N_5547,N_5463,N_5467);
and U5548 (N_5548,N_5489,N_5422);
nand U5549 (N_5549,N_5477,N_5455);
or U5550 (N_5550,N_5491,N_5389);
xnor U5551 (N_5551,N_5394,N_5482);
nor U5552 (N_5552,N_5388,N_5443);
nor U5553 (N_5553,N_5494,N_5458);
or U5554 (N_5554,N_5416,N_5460);
and U5555 (N_5555,N_5447,N_5392);
or U5556 (N_5556,N_5473,N_5453);
xnor U5557 (N_5557,N_5492,N_5391);
and U5558 (N_5558,N_5414,N_5493);
nor U5559 (N_5559,N_5429,N_5439);
and U5560 (N_5560,N_5469,N_5488);
nand U5561 (N_5561,N_5428,N_5415);
nand U5562 (N_5562,N_5378,N_5391);
xnor U5563 (N_5563,N_5437,N_5446);
xor U5564 (N_5564,N_5421,N_5417);
nor U5565 (N_5565,N_5414,N_5380);
nand U5566 (N_5566,N_5384,N_5426);
nor U5567 (N_5567,N_5481,N_5463);
nor U5568 (N_5568,N_5468,N_5477);
or U5569 (N_5569,N_5437,N_5380);
nor U5570 (N_5570,N_5397,N_5483);
or U5571 (N_5571,N_5496,N_5389);
nand U5572 (N_5572,N_5383,N_5492);
and U5573 (N_5573,N_5385,N_5478);
xor U5574 (N_5574,N_5479,N_5451);
xnor U5575 (N_5575,N_5499,N_5376);
or U5576 (N_5576,N_5441,N_5484);
or U5577 (N_5577,N_5499,N_5383);
xor U5578 (N_5578,N_5409,N_5387);
or U5579 (N_5579,N_5440,N_5485);
and U5580 (N_5580,N_5420,N_5397);
nand U5581 (N_5581,N_5449,N_5425);
nand U5582 (N_5582,N_5464,N_5465);
or U5583 (N_5583,N_5411,N_5387);
nand U5584 (N_5584,N_5478,N_5480);
xnor U5585 (N_5585,N_5388,N_5405);
nor U5586 (N_5586,N_5490,N_5408);
xor U5587 (N_5587,N_5428,N_5383);
xnor U5588 (N_5588,N_5391,N_5419);
nor U5589 (N_5589,N_5433,N_5443);
nor U5590 (N_5590,N_5487,N_5463);
or U5591 (N_5591,N_5487,N_5489);
and U5592 (N_5592,N_5394,N_5479);
or U5593 (N_5593,N_5398,N_5480);
nor U5594 (N_5594,N_5453,N_5449);
and U5595 (N_5595,N_5400,N_5461);
or U5596 (N_5596,N_5412,N_5403);
and U5597 (N_5597,N_5458,N_5439);
xor U5598 (N_5598,N_5484,N_5455);
nor U5599 (N_5599,N_5388,N_5450);
or U5600 (N_5600,N_5378,N_5495);
xnor U5601 (N_5601,N_5485,N_5414);
xnor U5602 (N_5602,N_5468,N_5444);
or U5603 (N_5603,N_5389,N_5487);
nand U5604 (N_5604,N_5394,N_5426);
xor U5605 (N_5605,N_5381,N_5437);
xor U5606 (N_5606,N_5382,N_5379);
or U5607 (N_5607,N_5413,N_5416);
or U5608 (N_5608,N_5421,N_5430);
xor U5609 (N_5609,N_5475,N_5400);
nand U5610 (N_5610,N_5440,N_5444);
nand U5611 (N_5611,N_5430,N_5451);
nor U5612 (N_5612,N_5397,N_5480);
nand U5613 (N_5613,N_5450,N_5467);
xnor U5614 (N_5614,N_5396,N_5415);
and U5615 (N_5615,N_5388,N_5376);
xor U5616 (N_5616,N_5441,N_5487);
nand U5617 (N_5617,N_5379,N_5494);
or U5618 (N_5618,N_5461,N_5375);
or U5619 (N_5619,N_5437,N_5414);
or U5620 (N_5620,N_5445,N_5424);
and U5621 (N_5621,N_5444,N_5428);
xor U5622 (N_5622,N_5419,N_5427);
nor U5623 (N_5623,N_5462,N_5401);
xnor U5624 (N_5624,N_5406,N_5392);
nand U5625 (N_5625,N_5580,N_5532);
xor U5626 (N_5626,N_5623,N_5517);
nor U5627 (N_5627,N_5583,N_5616);
nor U5628 (N_5628,N_5602,N_5548);
nand U5629 (N_5629,N_5550,N_5614);
and U5630 (N_5630,N_5593,N_5565);
nand U5631 (N_5631,N_5527,N_5554);
nor U5632 (N_5632,N_5621,N_5526);
and U5633 (N_5633,N_5610,N_5609);
nand U5634 (N_5634,N_5539,N_5543);
nand U5635 (N_5635,N_5562,N_5612);
or U5636 (N_5636,N_5589,N_5533);
nor U5637 (N_5637,N_5608,N_5500);
and U5638 (N_5638,N_5592,N_5618);
xnor U5639 (N_5639,N_5513,N_5587);
xnor U5640 (N_5640,N_5509,N_5557);
and U5641 (N_5641,N_5617,N_5505);
and U5642 (N_5642,N_5619,N_5572);
nand U5643 (N_5643,N_5535,N_5512);
nor U5644 (N_5644,N_5624,N_5515);
nand U5645 (N_5645,N_5605,N_5521);
nor U5646 (N_5646,N_5540,N_5560);
nand U5647 (N_5647,N_5520,N_5607);
and U5648 (N_5648,N_5586,N_5516);
xor U5649 (N_5649,N_5551,N_5518);
and U5650 (N_5650,N_5547,N_5567);
nor U5651 (N_5651,N_5504,N_5541);
and U5652 (N_5652,N_5530,N_5581);
and U5653 (N_5653,N_5603,N_5542);
and U5654 (N_5654,N_5552,N_5503);
xor U5655 (N_5655,N_5506,N_5531);
and U5656 (N_5656,N_5555,N_5622);
and U5657 (N_5657,N_5588,N_5613);
and U5658 (N_5658,N_5596,N_5601);
or U5659 (N_5659,N_5615,N_5574);
nand U5660 (N_5660,N_5620,N_5508);
xor U5661 (N_5661,N_5595,N_5546);
and U5662 (N_5662,N_5510,N_5575);
or U5663 (N_5663,N_5570,N_5528);
nand U5664 (N_5664,N_5573,N_5598);
or U5665 (N_5665,N_5523,N_5564);
or U5666 (N_5666,N_5594,N_5600);
nor U5667 (N_5667,N_5604,N_5514);
and U5668 (N_5668,N_5585,N_5534);
nor U5669 (N_5669,N_5599,N_5590);
or U5670 (N_5670,N_5529,N_5569);
xnor U5671 (N_5671,N_5571,N_5566);
xor U5672 (N_5672,N_5502,N_5559);
and U5673 (N_5673,N_5563,N_5579);
xor U5674 (N_5674,N_5578,N_5507);
nand U5675 (N_5675,N_5545,N_5553);
xnor U5676 (N_5676,N_5606,N_5577);
or U5677 (N_5677,N_5519,N_5501);
and U5678 (N_5678,N_5582,N_5544);
xnor U5679 (N_5679,N_5556,N_5538);
and U5680 (N_5680,N_5597,N_5536);
and U5681 (N_5681,N_5522,N_5561);
or U5682 (N_5682,N_5584,N_5549);
nor U5683 (N_5683,N_5611,N_5568);
or U5684 (N_5684,N_5558,N_5511);
xor U5685 (N_5685,N_5591,N_5525);
nor U5686 (N_5686,N_5524,N_5537);
nor U5687 (N_5687,N_5576,N_5522);
nor U5688 (N_5688,N_5618,N_5532);
nor U5689 (N_5689,N_5575,N_5570);
or U5690 (N_5690,N_5542,N_5514);
nor U5691 (N_5691,N_5620,N_5549);
xor U5692 (N_5692,N_5608,N_5579);
nor U5693 (N_5693,N_5608,N_5542);
nor U5694 (N_5694,N_5515,N_5593);
and U5695 (N_5695,N_5546,N_5579);
nor U5696 (N_5696,N_5574,N_5591);
and U5697 (N_5697,N_5581,N_5509);
xor U5698 (N_5698,N_5544,N_5509);
nor U5699 (N_5699,N_5539,N_5522);
nand U5700 (N_5700,N_5508,N_5513);
nor U5701 (N_5701,N_5590,N_5579);
nor U5702 (N_5702,N_5581,N_5534);
and U5703 (N_5703,N_5602,N_5623);
xor U5704 (N_5704,N_5569,N_5581);
nor U5705 (N_5705,N_5514,N_5595);
nor U5706 (N_5706,N_5570,N_5615);
nor U5707 (N_5707,N_5618,N_5522);
xnor U5708 (N_5708,N_5500,N_5581);
or U5709 (N_5709,N_5528,N_5553);
nand U5710 (N_5710,N_5510,N_5609);
or U5711 (N_5711,N_5570,N_5503);
xnor U5712 (N_5712,N_5611,N_5589);
nor U5713 (N_5713,N_5570,N_5608);
or U5714 (N_5714,N_5500,N_5527);
nor U5715 (N_5715,N_5587,N_5592);
or U5716 (N_5716,N_5559,N_5508);
nand U5717 (N_5717,N_5621,N_5564);
nand U5718 (N_5718,N_5582,N_5551);
nand U5719 (N_5719,N_5526,N_5577);
xor U5720 (N_5720,N_5539,N_5587);
and U5721 (N_5721,N_5537,N_5539);
or U5722 (N_5722,N_5543,N_5523);
xor U5723 (N_5723,N_5589,N_5588);
nand U5724 (N_5724,N_5608,N_5566);
nor U5725 (N_5725,N_5593,N_5542);
nand U5726 (N_5726,N_5596,N_5556);
xnor U5727 (N_5727,N_5582,N_5561);
nor U5728 (N_5728,N_5522,N_5540);
xnor U5729 (N_5729,N_5513,N_5620);
nand U5730 (N_5730,N_5522,N_5571);
xnor U5731 (N_5731,N_5595,N_5559);
xnor U5732 (N_5732,N_5514,N_5591);
xor U5733 (N_5733,N_5581,N_5568);
or U5734 (N_5734,N_5527,N_5601);
nor U5735 (N_5735,N_5501,N_5516);
or U5736 (N_5736,N_5539,N_5593);
or U5737 (N_5737,N_5595,N_5574);
or U5738 (N_5738,N_5521,N_5622);
xnor U5739 (N_5739,N_5545,N_5588);
or U5740 (N_5740,N_5583,N_5515);
nand U5741 (N_5741,N_5591,N_5522);
xor U5742 (N_5742,N_5542,N_5565);
and U5743 (N_5743,N_5537,N_5612);
nand U5744 (N_5744,N_5544,N_5534);
nand U5745 (N_5745,N_5616,N_5537);
nor U5746 (N_5746,N_5518,N_5548);
and U5747 (N_5747,N_5617,N_5553);
xnor U5748 (N_5748,N_5542,N_5574);
nor U5749 (N_5749,N_5533,N_5602);
nand U5750 (N_5750,N_5671,N_5711);
xnor U5751 (N_5751,N_5742,N_5692);
xnor U5752 (N_5752,N_5724,N_5647);
xnor U5753 (N_5753,N_5746,N_5687);
or U5754 (N_5754,N_5749,N_5659);
or U5755 (N_5755,N_5676,N_5663);
nand U5756 (N_5756,N_5715,N_5716);
nor U5757 (N_5757,N_5734,N_5726);
and U5758 (N_5758,N_5675,N_5635);
nor U5759 (N_5759,N_5627,N_5737);
nor U5760 (N_5760,N_5643,N_5625);
and U5761 (N_5761,N_5631,N_5740);
or U5762 (N_5762,N_5634,N_5654);
or U5763 (N_5763,N_5697,N_5673);
or U5764 (N_5764,N_5641,N_5668);
and U5765 (N_5765,N_5665,N_5702);
nor U5766 (N_5766,N_5661,N_5704);
xnor U5767 (N_5767,N_5730,N_5728);
and U5768 (N_5768,N_5735,N_5690);
nor U5769 (N_5769,N_5649,N_5679);
and U5770 (N_5770,N_5693,N_5733);
xnor U5771 (N_5771,N_5655,N_5656);
or U5772 (N_5772,N_5664,N_5630);
and U5773 (N_5773,N_5744,N_5718);
nand U5774 (N_5774,N_5695,N_5717);
xor U5775 (N_5775,N_5731,N_5719);
nand U5776 (N_5776,N_5698,N_5644);
xnor U5777 (N_5777,N_5642,N_5651);
nor U5778 (N_5778,N_5712,N_5632);
or U5779 (N_5779,N_5696,N_5710);
nand U5780 (N_5780,N_5729,N_5682);
xor U5781 (N_5781,N_5722,N_5694);
xnor U5782 (N_5782,N_5684,N_5713);
or U5783 (N_5783,N_5677,N_5670);
and U5784 (N_5784,N_5738,N_5640);
or U5785 (N_5785,N_5660,N_5645);
or U5786 (N_5786,N_5736,N_5748);
and U5787 (N_5787,N_5699,N_5741);
xnor U5788 (N_5788,N_5723,N_5666);
xnor U5789 (N_5789,N_5637,N_5688);
and U5790 (N_5790,N_5662,N_5709);
and U5791 (N_5791,N_5629,N_5747);
nand U5792 (N_5792,N_5725,N_5653);
nor U5793 (N_5793,N_5639,N_5674);
nor U5794 (N_5794,N_5628,N_5680);
xnor U5795 (N_5795,N_5727,N_5691);
and U5796 (N_5796,N_5720,N_5650);
or U5797 (N_5797,N_5648,N_5721);
nor U5798 (N_5798,N_5626,N_5700);
xor U5799 (N_5799,N_5705,N_5745);
xor U5800 (N_5800,N_5686,N_5701);
xnor U5801 (N_5801,N_5657,N_5714);
and U5802 (N_5802,N_5732,N_5708);
nand U5803 (N_5803,N_5743,N_5703);
xnor U5804 (N_5804,N_5672,N_5633);
and U5805 (N_5805,N_5683,N_5646);
nand U5806 (N_5806,N_5739,N_5652);
or U5807 (N_5807,N_5681,N_5678);
or U5808 (N_5808,N_5636,N_5685);
xor U5809 (N_5809,N_5689,N_5706);
and U5810 (N_5810,N_5669,N_5658);
or U5811 (N_5811,N_5667,N_5707);
nor U5812 (N_5812,N_5638,N_5700);
nor U5813 (N_5813,N_5655,N_5747);
nor U5814 (N_5814,N_5654,N_5718);
and U5815 (N_5815,N_5643,N_5691);
nor U5816 (N_5816,N_5711,N_5691);
xor U5817 (N_5817,N_5631,N_5654);
xnor U5818 (N_5818,N_5738,N_5703);
nor U5819 (N_5819,N_5683,N_5658);
and U5820 (N_5820,N_5687,N_5642);
or U5821 (N_5821,N_5665,N_5746);
nor U5822 (N_5822,N_5698,N_5681);
xnor U5823 (N_5823,N_5685,N_5720);
nand U5824 (N_5824,N_5705,N_5692);
and U5825 (N_5825,N_5731,N_5748);
or U5826 (N_5826,N_5688,N_5685);
and U5827 (N_5827,N_5667,N_5629);
and U5828 (N_5828,N_5665,N_5669);
and U5829 (N_5829,N_5686,N_5739);
and U5830 (N_5830,N_5732,N_5641);
nor U5831 (N_5831,N_5636,N_5666);
xnor U5832 (N_5832,N_5693,N_5625);
nand U5833 (N_5833,N_5650,N_5715);
nor U5834 (N_5834,N_5745,N_5675);
or U5835 (N_5835,N_5708,N_5681);
or U5836 (N_5836,N_5740,N_5675);
or U5837 (N_5837,N_5703,N_5693);
or U5838 (N_5838,N_5683,N_5647);
or U5839 (N_5839,N_5746,N_5727);
and U5840 (N_5840,N_5705,N_5667);
nor U5841 (N_5841,N_5655,N_5748);
and U5842 (N_5842,N_5628,N_5721);
xnor U5843 (N_5843,N_5679,N_5633);
nand U5844 (N_5844,N_5672,N_5696);
nor U5845 (N_5845,N_5635,N_5686);
or U5846 (N_5846,N_5749,N_5672);
or U5847 (N_5847,N_5658,N_5739);
nand U5848 (N_5848,N_5749,N_5666);
nand U5849 (N_5849,N_5682,N_5636);
nand U5850 (N_5850,N_5702,N_5659);
nor U5851 (N_5851,N_5744,N_5643);
xor U5852 (N_5852,N_5633,N_5691);
or U5853 (N_5853,N_5653,N_5627);
or U5854 (N_5854,N_5667,N_5668);
and U5855 (N_5855,N_5664,N_5665);
or U5856 (N_5856,N_5653,N_5655);
or U5857 (N_5857,N_5688,N_5734);
and U5858 (N_5858,N_5638,N_5637);
nor U5859 (N_5859,N_5640,N_5644);
nand U5860 (N_5860,N_5709,N_5633);
xnor U5861 (N_5861,N_5741,N_5661);
xor U5862 (N_5862,N_5716,N_5682);
and U5863 (N_5863,N_5720,N_5712);
nand U5864 (N_5864,N_5667,N_5649);
xnor U5865 (N_5865,N_5677,N_5628);
nor U5866 (N_5866,N_5721,N_5668);
or U5867 (N_5867,N_5663,N_5747);
and U5868 (N_5868,N_5711,N_5697);
or U5869 (N_5869,N_5637,N_5747);
nor U5870 (N_5870,N_5627,N_5718);
or U5871 (N_5871,N_5647,N_5630);
xor U5872 (N_5872,N_5657,N_5673);
nand U5873 (N_5873,N_5710,N_5720);
or U5874 (N_5874,N_5636,N_5727);
and U5875 (N_5875,N_5799,N_5863);
or U5876 (N_5876,N_5845,N_5834);
and U5877 (N_5877,N_5757,N_5840);
nand U5878 (N_5878,N_5761,N_5788);
xnor U5879 (N_5879,N_5855,N_5812);
nand U5880 (N_5880,N_5820,N_5755);
xnor U5881 (N_5881,N_5803,N_5769);
and U5882 (N_5882,N_5865,N_5821);
and U5883 (N_5883,N_5779,N_5854);
nand U5884 (N_5884,N_5833,N_5817);
or U5885 (N_5885,N_5847,N_5774);
or U5886 (N_5886,N_5866,N_5811);
nor U5887 (N_5887,N_5829,N_5760);
nand U5888 (N_5888,N_5825,N_5835);
xnor U5889 (N_5889,N_5838,N_5782);
and U5890 (N_5890,N_5853,N_5816);
and U5891 (N_5891,N_5780,N_5837);
nor U5892 (N_5892,N_5762,N_5867);
nor U5893 (N_5893,N_5809,N_5787);
or U5894 (N_5894,N_5756,N_5860);
nor U5895 (N_5895,N_5842,N_5831);
xnor U5896 (N_5896,N_5850,N_5818);
and U5897 (N_5897,N_5822,N_5832);
xor U5898 (N_5898,N_5797,N_5870);
nand U5899 (N_5899,N_5794,N_5871);
xnor U5900 (N_5900,N_5868,N_5862);
and U5901 (N_5901,N_5805,N_5751);
nor U5902 (N_5902,N_5857,N_5828);
nor U5903 (N_5903,N_5784,N_5851);
nand U5904 (N_5904,N_5767,N_5802);
nand U5905 (N_5905,N_5792,N_5815);
nor U5906 (N_5906,N_5859,N_5770);
and U5907 (N_5907,N_5848,N_5861);
nor U5908 (N_5908,N_5858,N_5874);
xnor U5909 (N_5909,N_5873,N_5852);
nor U5910 (N_5910,N_5776,N_5785);
nand U5911 (N_5911,N_5795,N_5823);
and U5912 (N_5912,N_5772,N_5786);
nand U5913 (N_5913,N_5778,N_5758);
nor U5914 (N_5914,N_5872,N_5801);
xor U5915 (N_5915,N_5846,N_5798);
nor U5916 (N_5916,N_5819,N_5789);
and U5917 (N_5917,N_5775,N_5777);
and U5918 (N_5918,N_5752,N_5839);
xor U5919 (N_5919,N_5754,N_5808);
nand U5920 (N_5920,N_5759,N_5781);
and U5921 (N_5921,N_5810,N_5826);
or U5922 (N_5922,N_5806,N_5791);
nand U5923 (N_5923,N_5783,N_5836);
or U5924 (N_5924,N_5804,N_5764);
nor U5925 (N_5925,N_5827,N_5793);
xnor U5926 (N_5926,N_5807,N_5841);
nor U5927 (N_5927,N_5814,N_5750);
or U5928 (N_5928,N_5766,N_5864);
xor U5929 (N_5929,N_5790,N_5796);
xnor U5930 (N_5930,N_5768,N_5856);
nor U5931 (N_5931,N_5763,N_5753);
nor U5932 (N_5932,N_5824,N_5800);
nor U5933 (N_5933,N_5765,N_5869);
nand U5934 (N_5934,N_5773,N_5813);
or U5935 (N_5935,N_5771,N_5844);
nand U5936 (N_5936,N_5843,N_5830);
nand U5937 (N_5937,N_5849,N_5842);
nor U5938 (N_5938,N_5870,N_5809);
nand U5939 (N_5939,N_5823,N_5822);
and U5940 (N_5940,N_5772,N_5826);
xor U5941 (N_5941,N_5865,N_5761);
and U5942 (N_5942,N_5871,N_5758);
nand U5943 (N_5943,N_5835,N_5866);
or U5944 (N_5944,N_5831,N_5845);
and U5945 (N_5945,N_5843,N_5868);
xnor U5946 (N_5946,N_5814,N_5787);
or U5947 (N_5947,N_5804,N_5826);
or U5948 (N_5948,N_5802,N_5874);
xor U5949 (N_5949,N_5849,N_5812);
nor U5950 (N_5950,N_5869,N_5764);
or U5951 (N_5951,N_5823,N_5775);
nor U5952 (N_5952,N_5847,N_5816);
nor U5953 (N_5953,N_5766,N_5810);
nand U5954 (N_5954,N_5785,N_5817);
nor U5955 (N_5955,N_5849,N_5796);
or U5956 (N_5956,N_5833,N_5866);
nand U5957 (N_5957,N_5870,N_5754);
and U5958 (N_5958,N_5872,N_5783);
and U5959 (N_5959,N_5782,N_5774);
nand U5960 (N_5960,N_5830,N_5804);
xnor U5961 (N_5961,N_5754,N_5863);
or U5962 (N_5962,N_5856,N_5809);
nor U5963 (N_5963,N_5822,N_5860);
or U5964 (N_5964,N_5821,N_5790);
nand U5965 (N_5965,N_5799,N_5803);
xor U5966 (N_5966,N_5758,N_5867);
nor U5967 (N_5967,N_5863,N_5853);
nand U5968 (N_5968,N_5795,N_5799);
xnor U5969 (N_5969,N_5809,N_5813);
and U5970 (N_5970,N_5785,N_5845);
and U5971 (N_5971,N_5834,N_5766);
and U5972 (N_5972,N_5842,N_5789);
or U5973 (N_5973,N_5829,N_5800);
nor U5974 (N_5974,N_5812,N_5762);
or U5975 (N_5975,N_5786,N_5861);
nor U5976 (N_5976,N_5795,N_5764);
nand U5977 (N_5977,N_5771,N_5757);
and U5978 (N_5978,N_5760,N_5778);
nor U5979 (N_5979,N_5818,N_5757);
and U5980 (N_5980,N_5785,N_5823);
nor U5981 (N_5981,N_5839,N_5818);
nand U5982 (N_5982,N_5784,N_5846);
and U5983 (N_5983,N_5871,N_5775);
xnor U5984 (N_5984,N_5814,N_5872);
xnor U5985 (N_5985,N_5821,N_5845);
or U5986 (N_5986,N_5787,N_5790);
xor U5987 (N_5987,N_5799,N_5839);
xor U5988 (N_5988,N_5758,N_5866);
xor U5989 (N_5989,N_5801,N_5854);
nand U5990 (N_5990,N_5811,N_5851);
or U5991 (N_5991,N_5789,N_5793);
xnor U5992 (N_5992,N_5858,N_5872);
and U5993 (N_5993,N_5819,N_5807);
nor U5994 (N_5994,N_5807,N_5791);
nor U5995 (N_5995,N_5801,N_5835);
xor U5996 (N_5996,N_5784,N_5775);
nand U5997 (N_5997,N_5821,N_5774);
nand U5998 (N_5998,N_5785,N_5810);
or U5999 (N_5999,N_5855,N_5765);
xnor U6000 (N_6000,N_5894,N_5914);
and U6001 (N_6001,N_5942,N_5919);
and U6002 (N_6002,N_5879,N_5975);
xnor U6003 (N_6003,N_5999,N_5916);
nor U6004 (N_6004,N_5949,N_5977);
nand U6005 (N_6005,N_5971,N_5891);
or U6006 (N_6006,N_5944,N_5943);
nor U6007 (N_6007,N_5966,N_5945);
or U6008 (N_6008,N_5970,N_5994);
nand U6009 (N_6009,N_5881,N_5991);
and U6010 (N_6010,N_5963,N_5960);
nand U6011 (N_6011,N_5933,N_5956);
and U6012 (N_6012,N_5954,N_5998);
xor U6013 (N_6013,N_5896,N_5987);
xnor U6014 (N_6014,N_5926,N_5951);
nand U6015 (N_6015,N_5952,N_5899);
nand U6016 (N_6016,N_5875,N_5953);
or U6017 (N_6017,N_5989,N_5969);
xor U6018 (N_6018,N_5887,N_5938);
nand U6019 (N_6019,N_5900,N_5957);
nand U6020 (N_6020,N_5993,N_5934);
nand U6021 (N_6021,N_5984,N_5913);
and U6022 (N_6022,N_5893,N_5990);
nor U6023 (N_6023,N_5904,N_5927);
xnor U6024 (N_6024,N_5915,N_5986);
or U6025 (N_6025,N_5907,N_5895);
or U6026 (N_6026,N_5923,N_5947);
nor U6027 (N_6027,N_5889,N_5892);
nand U6028 (N_6028,N_5978,N_5924);
nand U6029 (N_6029,N_5882,N_5902);
or U6030 (N_6030,N_5906,N_5884);
nor U6031 (N_6031,N_5950,N_5964);
nand U6032 (N_6032,N_5901,N_5905);
and U6033 (N_6033,N_5903,N_5911);
and U6034 (N_6034,N_5929,N_5948);
and U6035 (N_6035,N_5918,N_5910);
xor U6036 (N_6036,N_5932,N_5922);
nor U6037 (N_6037,N_5937,N_5886);
nand U6038 (N_6038,N_5939,N_5968);
nor U6039 (N_6039,N_5885,N_5909);
and U6040 (N_6040,N_5981,N_5976);
nand U6041 (N_6041,N_5931,N_5983);
or U6042 (N_6042,N_5890,N_5912);
nor U6043 (N_6043,N_5941,N_5920);
nand U6044 (N_6044,N_5962,N_5997);
xor U6045 (N_6045,N_5930,N_5974);
or U6046 (N_6046,N_5965,N_5880);
xnor U6047 (N_6047,N_5898,N_5936);
xor U6048 (N_6048,N_5972,N_5946);
xnor U6049 (N_6049,N_5980,N_5973);
nand U6050 (N_6050,N_5995,N_5921);
xor U6051 (N_6051,N_5955,N_5935);
nand U6052 (N_6052,N_5925,N_5917);
xnor U6053 (N_6053,N_5940,N_5996);
nand U6054 (N_6054,N_5992,N_5979);
or U6055 (N_6055,N_5985,N_5988);
nand U6056 (N_6056,N_5878,N_5967);
nand U6057 (N_6057,N_5958,N_5908);
xnor U6058 (N_6058,N_5959,N_5883);
nor U6059 (N_6059,N_5877,N_5876);
nor U6060 (N_6060,N_5961,N_5982);
nor U6061 (N_6061,N_5928,N_5897);
xnor U6062 (N_6062,N_5888,N_5876);
or U6063 (N_6063,N_5967,N_5990);
or U6064 (N_6064,N_5939,N_5982);
xnor U6065 (N_6065,N_5911,N_5950);
nor U6066 (N_6066,N_5999,N_5989);
nand U6067 (N_6067,N_5968,N_5984);
or U6068 (N_6068,N_5911,N_5907);
nand U6069 (N_6069,N_5954,N_5970);
nor U6070 (N_6070,N_5915,N_5882);
and U6071 (N_6071,N_5907,N_5949);
nor U6072 (N_6072,N_5880,N_5979);
xor U6073 (N_6073,N_5939,N_5906);
nand U6074 (N_6074,N_5912,N_5899);
and U6075 (N_6075,N_5909,N_5979);
xor U6076 (N_6076,N_5886,N_5979);
nor U6077 (N_6077,N_5925,N_5926);
and U6078 (N_6078,N_5939,N_5981);
nand U6079 (N_6079,N_5940,N_5882);
and U6080 (N_6080,N_5994,N_5917);
or U6081 (N_6081,N_5924,N_5992);
nand U6082 (N_6082,N_5941,N_5969);
and U6083 (N_6083,N_5957,N_5916);
or U6084 (N_6084,N_5879,N_5912);
or U6085 (N_6085,N_5953,N_5928);
nand U6086 (N_6086,N_5895,N_5927);
and U6087 (N_6087,N_5982,N_5930);
nand U6088 (N_6088,N_5890,N_5892);
nand U6089 (N_6089,N_5880,N_5962);
or U6090 (N_6090,N_5949,N_5915);
nor U6091 (N_6091,N_5953,N_5978);
xnor U6092 (N_6092,N_5956,N_5879);
nor U6093 (N_6093,N_5955,N_5991);
or U6094 (N_6094,N_5966,N_5921);
xnor U6095 (N_6095,N_5966,N_5905);
nand U6096 (N_6096,N_5926,N_5903);
nor U6097 (N_6097,N_5996,N_5908);
nor U6098 (N_6098,N_5931,N_5877);
or U6099 (N_6099,N_5880,N_5998);
nand U6100 (N_6100,N_5974,N_5977);
and U6101 (N_6101,N_5888,N_5952);
or U6102 (N_6102,N_5920,N_5995);
xnor U6103 (N_6103,N_5937,N_5974);
and U6104 (N_6104,N_5964,N_5997);
xnor U6105 (N_6105,N_5952,N_5943);
xor U6106 (N_6106,N_5972,N_5937);
or U6107 (N_6107,N_5991,N_5893);
or U6108 (N_6108,N_5899,N_5905);
xor U6109 (N_6109,N_5956,N_5890);
and U6110 (N_6110,N_5875,N_5929);
or U6111 (N_6111,N_5881,N_5929);
nand U6112 (N_6112,N_5929,N_5957);
xor U6113 (N_6113,N_5918,N_5939);
and U6114 (N_6114,N_5876,N_5950);
xor U6115 (N_6115,N_5932,N_5973);
or U6116 (N_6116,N_5966,N_5903);
nor U6117 (N_6117,N_5922,N_5967);
nor U6118 (N_6118,N_5916,N_5960);
nor U6119 (N_6119,N_5980,N_5928);
nand U6120 (N_6120,N_5959,N_5898);
and U6121 (N_6121,N_5973,N_5927);
and U6122 (N_6122,N_5978,N_5919);
nand U6123 (N_6123,N_5941,N_5976);
nor U6124 (N_6124,N_5892,N_5921);
nor U6125 (N_6125,N_6075,N_6027);
nor U6126 (N_6126,N_6017,N_6080);
xor U6127 (N_6127,N_6042,N_6029);
and U6128 (N_6128,N_6007,N_6022);
xor U6129 (N_6129,N_6054,N_6081);
nand U6130 (N_6130,N_6100,N_6019);
nor U6131 (N_6131,N_6055,N_6111);
nand U6132 (N_6132,N_6059,N_6043);
nor U6133 (N_6133,N_6089,N_6020);
nor U6134 (N_6134,N_6066,N_6032);
xor U6135 (N_6135,N_6114,N_6082);
xor U6136 (N_6136,N_6049,N_6069);
nand U6137 (N_6137,N_6067,N_6098);
and U6138 (N_6138,N_6009,N_6006);
nand U6139 (N_6139,N_6103,N_6086);
or U6140 (N_6140,N_6018,N_6031);
xor U6141 (N_6141,N_6104,N_6025);
and U6142 (N_6142,N_6105,N_6000);
xor U6143 (N_6143,N_6110,N_6002);
and U6144 (N_6144,N_6041,N_6109);
and U6145 (N_6145,N_6078,N_6060);
nor U6146 (N_6146,N_6021,N_6062);
and U6147 (N_6147,N_6063,N_6064);
nand U6148 (N_6148,N_6004,N_6047);
nor U6149 (N_6149,N_6124,N_6011);
xnor U6150 (N_6150,N_6088,N_6096);
nand U6151 (N_6151,N_6106,N_6051);
xnor U6152 (N_6152,N_6123,N_6087);
xor U6153 (N_6153,N_6076,N_6074);
nor U6154 (N_6154,N_6052,N_6099);
nand U6155 (N_6155,N_6003,N_6094);
nor U6156 (N_6156,N_6045,N_6001);
nor U6157 (N_6157,N_6084,N_6048);
xnor U6158 (N_6158,N_6073,N_6065);
nand U6159 (N_6159,N_6097,N_6122);
or U6160 (N_6160,N_6085,N_6046);
nand U6161 (N_6161,N_6068,N_6117);
xnor U6162 (N_6162,N_6077,N_6024);
and U6163 (N_6163,N_6038,N_6058);
xnor U6164 (N_6164,N_6023,N_6108);
xor U6165 (N_6165,N_6013,N_6014);
nor U6166 (N_6166,N_6034,N_6071);
and U6167 (N_6167,N_6118,N_6036);
and U6168 (N_6168,N_6061,N_6070);
nor U6169 (N_6169,N_6056,N_6119);
xnor U6170 (N_6170,N_6016,N_6101);
nand U6171 (N_6171,N_6026,N_6107);
and U6172 (N_6172,N_6095,N_6053);
nor U6173 (N_6173,N_6005,N_6030);
nor U6174 (N_6174,N_6112,N_6028);
or U6175 (N_6175,N_6079,N_6057);
xnor U6176 (N_6176,N_6015,N_6037);
xnor U6177 (N_6177,N_6072,N_6008);
nor U6178 (N_6178,N_6091,N_6092);
xnor U6179 (N_6179,N_6093,N_6116);
or U6180 (N_6180,N_6102,N_6121);
xnor U6181 (N_6181,N_6050,N_6120);
nand U6182 (N_6182,N_6010,N_6113);
and U6183 (N_6183,N_6115,N_6090);
nand U6184 (N_6184,N_6033,N_6044);
or U6185 (N_6185,N_6039,N_6040);
and U6186 (N_6186,N_6083,N_6035);
or U6187 (N_6187,N_6012,N_6043);
xor U6188 (N_6188,N_6040,N_6097);
nand U6189 (N_6189,N_6032,N_6063);
or U6190 (N_6190,N_6049,N_6056);
nand U6191 (N_6191,N_6095,N_6019);
or U6192 (N_6192,N_6095,N_6083);
and U6193 (N_6193,N_6114,N_6116);
and U6194 (N_6194,N_6006,N_6122);
or U6195 (N_6195,N_6090,N_6078);
nand U6196 (N_6196,N_6090,N_6072);
and U6197 (N_6197,N_6119,N_6057);
xor U6198 (N_6198,N_6027,N_6084);
xor U6199 (N_6199,N_6002,N_6008);
xor U6200 (N_6200,N_6080,N_6121);
xnor U6201 (N_6201,N_6116,N_6101);
xor U6202 (N_6202,N_6005,N_6004);
or U6203 (N_6203,N_6046,N_6084);
xnor U6204 (N_6204,N_6018,N_6023);
or U6205 (N_6205,N_6032,N_6107);
xnor U6206 (N_6206,N_6013,N_6034);
and U6207 (N_6207,N_6064,N_6042);
nor U6208 (N_6208,N_6018,N_6102);
nand U6209 (N_6209,N_6033,N_6060);
nand U6210 (N_6210,N_6073,N_6022);
and U6211 (N_6211,N_6072,N_6074);
or U6212 (N_6212,N_6078,N_6100);
xnor U6213 (N_6213,N_6078,N_6097);
nor U6214 (N_6214,N_6123,N_6050);
nor U6215 (N_6215,N_6031,N_6104);
nand U6216 (N_6216,N_6035,N_6098);
and U6217 (N_6217,N_6019,N_6009);
nand U6218 (N_6218,N_6078,N_6119);
or U6219 (N_6219,N_6090,N_6021);
or U6220 (N_6220,N_6087,N_6098);
nand U6221 (N_6221,N_6083,N_6087);
nand U6222 (N_6222,N_6117,N_6073);
nor U6223 (N_6223,N_6093,N_6117);
and U6224 (N_6224,N_6036,N_6058);
nand U6225 (N_6225,N_6088,N_6077);
xor U6226 (N_6226,N_6111,N_6075);
nand U6227 (N_6227,N_6110,N_6050);
xor U6228 (N_6228,N_6124,N_6078);
xor U6229 (N_6229,N_6092,N_6058);
and U6230 (N_6230,N_6083,N_6073);
nor U6231 (N_6231,N_6074,N_6026);
nor U6232 (N_6232,N_6023,N_6097);
nand U6233 (N_6233,N_6063,N_6013);
nand U6234 (N_6234,N_6081,N_6079);
or U6235 (N_6235,N_6035,N_6103);
xnor U6236 (N_6236,N_6097,N_6083);
nand U6237 (N_6237,N_6016,N_6068);
and U6238 (N_6238,N_6108,N_6087);
nor U6239 (N_6239,N_6053,N_6016);
and U6240 (N_6240,N_6113,N_6000);
nor U6241 (N_6241,N_6096,N_6117);
nor U6242 (N_6242,N_6040,N_6025);
and U6243 (N_6243,N_6008,N_6018);
nand U6244 (N_6244,N_6109,N_6124);
nor U6245 (N_6245,N_6023,N_6086);
and U6246 (N_6246,N_6028,N_6011);
nor U6247 (N_6247,N_6063,N_6094);
nand U6248 (N_6248,N_6078,N_6063);
or U6249 (N_6249,N_6113,N_6003);
nor U6250 (N_6250,N_6193,N_6185);
and U6251 (N_6251,N_6151,N_6189);
or U6252 (N_6252,N_6247,N_6128);
nand U6253 (N_6253,N_6212,N_6236);
nand U6254 (N_6254,N_6214,N_6175);
nand U6255 (N_6255,N_6216,N_6130);
xor U6256 (N_6256,N_6177,N_6150);
nand U6257 (N_6257,N_6141,N_6244);
xor U6258 (N_6258,N_6224,N_6181);
nor U6259 (N_6259,N_6184,N_6213);
nand U6260 (N_6260,N_6174,N_6140);
and U6261 (N_6261,N_6204,N_6182);
xnor U6262 (N_6262,N_6142,N_6195);
nand U6263 (N_6263,N_6132,N_6191);
nand U6264 (N_6264,N_6127,N_6183);
xor U6265 (N_6265,N_6240,N_6166);
nand U6266 (N_6266,N_6217,N_6241);
nand U6267 (N_6267,N_6125,N_6155);
nand U6268 (N_6268,N_6215,N_6199);
and U6269 (N_6269,N_6205,N_6176);
and U6270 (N_6270,N_6126,N_6234);
or U6271 (N_6271,N_6196,N_6197);
and U6272 (N_6272,N_6165,N_6163);
and U6273 (N_6273,N_6143,N_6146);
and U6274 (N_6274,N_6220,N_6167);
and U6275 (N_6275,N_6134,N_6190);
or U6276 (N_6276,N_6249,N_6180);
or U6277 (N_6277,N_6209,N_6170);
xor U6278 (N_6278,N_6237,N_6194);
nor U6279 (N_6279,N_6145,N_6242);
xnor U6280 (N_6280,N_6229,N_6172);
nand U6281 (N_6281,N_6248,N_6136);
xnor U6282 (N_6282,N_6187,N_6207);
nor U6283 (N_6283,N_6153,N_6233);
xor U6284 (N_6284,N_6203,N_6178);
and U6285 (N_6285,N_6179,N_6156);
or U6286 (N_6286,N_6202,N_6131);
nor U6287 (N_6287,N_6154,N_6210);
or U6288 (N_6288,N_6157,N_6186);
nand U6289 (N_6289,N_6149,N_6173);
nor U6290 (N_6290,N_6246,N_6171);
nor U6291 (N_6291,N_6168,N_6230);
and U6292 (N_6292,N_6138,N_6208);
nand U6293 (N_6293,N_6147,N_6225);
and U6294 (N_6294,N_6198,N_6152);
xor U6295 (N_6295,N_6211,N_6218);
nand U6296 (N_6296,N_6161,N_6235);
nand U6297 (N_6297,N_6200,N_6226);
nor U6298 (N_6298,N_6129,N_6243);
nand U6299 (N_6299,N_6135,N_6169);
nand U6300 (N_6300,N_6221,N_6144);
xnor U6301 (N_6301,N_6201,N_6222);
nor U6302 (N_6302,N_6239,N_6158);
nand U6303 (N_6303,N_6159,N_6231);
nand U6304 (N_6304,N_6232,N_6148);
or U6305 (N_6305,N_6164,N_6160);
and U6306 (N_6306,N_6162,N_6139);
nand U6307 (N_6307,N_6238,N_6133);
and U6308 (N_6308,N_6219,N_6206);
or U6309 (N_6309,N_6245,N_6188);
nand U6310 (N_6310,N_6227,N_6137);
and U6311 (N_6311,N_6228,N_6192);
xnor U6312 (N_6312,N_6223,N_6156);
xor U6313 (N_6313,N_6224,N_6163);
nand U6314 (N_6314,N_6126,N_6179);
xnor U6315 (N_6315,N_6179,N_6127);
and U6316 (N_6316,N_6157,N_6158);
nor U6317 (N_6317,N_6178,N_6172);
nand U6318 (N_6318,N_6227,N_6165);
or U6319 (N_6319,N_6146,N_6215);
nor U6320 (N_6320,N_6227,N_6125);
nor U6321 (N_6321,N_6147,N_6230);
nor U6322 (N_6322,N_6177,N_6175);
nor U6323 (N_6323,N_6166,N_6152);
nor U6324 (N_6324,N_6212,N_6180);
nand U6325 (N_6325,N_6242,N_6148);
or U6326 (N_6326,N_6159,N_6228);
nand U6327 (N_6327,N_6235,N_6244);
xor U6328 (N_6328,N_6201,N_6148);
nand U6329 (N_6329,N_6201,N_6185);
and U6330 (N_6330,N_6220,N_6170);
nor U6331 (N_6331,N_6144,N_6236);
nand U6332 (N_6332,N_6186,N_6237);
nand U6333 (N_6333,N_6151,N_6201);
and U6334 (N_6334,N_6184,N_6233);
or U6335 (N_6335,N_6182,N_6211);
or U6336 (N_6336,N_6156,N_6152);
nor U6337 (N_6337,N_6221,N_6209);
or U6338 (N_6338,N_6215,N_6198);
nand U6339 (N_6339,N_6241,N_6244);
nand U6340 (N_6340,N_6241,N_6128);
nand U6341 (N_6341,N_6137,N_6135);
or U6342 (N_6342,N_6140,N_6161);
xor U6343 (N_6343,N_6131,N_6193);
nand U6344 (N_6344,N_6142,N_6215);
or U6345 (N_6345,N_6165,N_6226);
and U6346 (N_6346,N_6130,N_6192);
or U6347 (N_6347,N_6148,N_6187);
nand U6348 (N_6348,N_6213,N_6247);
nor U6349 (N_6349,N_6242,N_6195);
or U6350 (N_6350,N_6150,N_6173);
nor U6351 (N_6351,N_6205,N_6153);
and U6352 (N_6352,N_6128,N_6237);
or U6353 (N_6353,N_6219,N_6227);
xor U6354 (N_6354,N_6172,N_6234);
nor U6355 (N_6355,N_6164,N_6197);
or U6356 (N_6356,N_6157,N_6146);
xor U6357 (N_6357,N_6245,N_6244);
and U6358 (N_6358,N_6182,N_6191);
nor U6359 (N_6359,N_6244,N_6201);
and U6360 (N_6360,N_6245,N_6176);
nor U6361 (N_6361,N_6200,N_6247);
nor U6362 (N_6362,N_6159,N_6131);
xor U6363 (N_6363,N_6173,N_6135);
or U6364 (N_6364,N_6227,N_6175);
or U6365 (N_6365,N_6208,N_6172);
nand U6366 (N_6366,N_6168,N_6202);
nor U6367 (N_6367,N_6183,N_6176);
nor U6368 (N_6368,N_6132,N_6180);
xor U6369 (N_6369,N_6140,N_6141);
and U6370 (N_6370,N_6131,N_6137);
and U6371 (N_6371,N_6229,N_6185);
and U6372 (N_6372,N_6141,N_6167);
or U6373 (N_6373,N_6241,N_6181);
and U6374 (N_6374,N_6208,N_6173);
nor U6375 (N_6375,N_6260,N_6344);
nand U6376 (N_6376,N_6345,N_6305);
and U6377 (N_6377,N_6301,N_6274);
nor U6378 (N_6378,N_6291,N_6330);
xor U6379 (N_6379,N_6350,N_6342);
nand U6380 (N_6380,N_6316,N_6261);
xor U6381 (N_6381,N_6292,N_6368);
and U6382 (N_6382,N_6290,N_6329);
nand U6383 (N_6383,N_6252,N_6311);
xor U6384 (N_6384,N_6323,N_6283);
nor U6385 (N_6385,N_6346,N_6349);
xor U6386 (N_6386,N_6262,N_6367);
and U6387 (N_6387,N_6319,N_6271);
xnor U6388 (N_6388,N_6321,N_6334);
or U6389 (N_6389,N_6318,N_6357);
or U6390 (N_6390,N_6270,N_6253);
xor U6391 (N_6391,N_6322,N_6338);
nand U6392 (N_6392,N_6313,N_6364);
or U6393 (N_6393,N_6303,N_6267);
and U6394 (N_6394,N_6273,N_6310);
nor U6395 (N_6395,N_6312,N_6255);
and U6396 (N_6396,N_6333,N_6356);
nand U6397 (N_6397,N_6361,N_6275);
and U6398 (N_6398,N_6337,N_6279);
xor U6399 (N_6399,N_6282,N_6307);
xor U6400 (N_6400,N_6299,N_6363);
or U6401 (N_6401,N_6256,N_6269);
nor U6402 (N_6402,N_6373,N_6293);
xor U6403 (N_6403,N_6298,N_6278);
xnor U6404 (N_6404,N_6365,N_6280);
and U6405 (N_6405,N_6353,N_6296);
and U6406 (N_6406,N_6258,N_6360);
nand U6407 (N_6407,N_6372,N_6352);
xnor U6408 (N_6408,N_6370,N_6281);
or U6409 (N_6409,N_6264,N_6347);
or U6410 (N_6410,N_6371,N_6287);
nand U6411 (N_6411,N_6266,N_6317);
or U6412 (N_6412,N_6263,N_6257);
xor U6413 (N_6413,N_6306,N_6351);
nand U6414 (N_6414,N_6288,N_6362);
or U6415 (N_6415,N_6336,N_6295);
nand U6416 (N_6416,N_6308,N_6325);
xnor U6417 (N_6417,N_6285,N_6339);
xnor U6418 (N_6418,N_6302,N_6374);
and U6419 (N_6419,N_6277,N_6276);
and U6420 (N_6420,N_6254,N_6272);
xnor U6421 (N_6421,N_6335,N_6265);
nor U6422 (N_6422,N_6369,N_6284);
nor U6423 (N_6423,N_6314,N_6289);
and U6424 (N_6424,N_6251,N_6355);
nand U6425 (N_6425,N_6348,N_6327);
nor U6426 (N_6426,N_6366,N_6331);
or U6427 (N_6427,N_6309,N_6268);
nor U6428 (N_6428,N_6354,N_6300);
nand U6429 (N_6429,N_6324,N_6340);
xor U6430 (N_6430,N_6326,N_6315);
nand U6431 (N_6431,N_6286,N_6250);
or U6432 (N_6432,N_6328,N_6294);
and U6433 (N_6433,N_6358,N_6259);
or U6434 (N_6434,N_6304,N_6343);
xnor U6435 (N_6435,N_6320,N_6297);
nor U6436 (N_6436,N_6332,N_6359);
or U6437 (N_6437,N_6341,N_6259);
nor U6438 (N_6438,N_6364,N_6303);
nor U6439 (N_6439,N_6274,N_6339);
nor U6440 (N_6440,N_6275,N_6320);
nor U6441 (N_6441,N_6358,N_6339);
and U6442 (N_6442,N_6286,N_6317);
nor U6443 (N_6443,N_6265,N_6346);
and U6444 (N_6444,N_6347,N_6314);
nand U6445 (N_6445,N_6255,N_6359);
nor U6446 (N_6446,N_6252,N_6257);
and U6447 (N_6447,N_6279,N_6336);
nand U6448 (N_6448,N_6285,N_6367);
nor U6449 (N_6449,N_6355,N_6293);
or U6450 (N_6450,N_6362,N_6251);
nand U6451 (N_6451,N_6269,N_6251);
or U6452 (N_6452,N_6311,N_6324);
or U6453 (N_6453,N_6316,N_6283);
xnor U6454 (N_6454,N_6353,N_6261);
xnor U6455 (N_6455,N_6305,N_6258);
nand U6456 (N_6456,N_6314,N_6313);
xnor U6457 (N_6457,N_6283,N_6358);
or U6458 (N_6458,N_6278,N_6319);
or U6459 (N_6459,N_6250,N_6339);
or U6460 (N_6460,N_6360,N_6312);
xor U6461 (N_6461,N_6350,N_6366);
or U6462 (N_6462,N_6369,N_6362);
xor U6463 (N_6463,N_6359,N_6334);
and U6464 (N_6464,N_6302,N_6341);
nand U6465 (N_6465,N_6273,N_6252);
nand U6466 (N_6466,N_6257,N_6366);
nor U6467 (N_6467,N_6338,N_6371);
or U6468 (N_6468,N_6268,N_6362);
xor U6469 (N_6469,N_6282,N_6369);
nor U6470 (N_6470,N_6332,N_6320);
nor U6471 (N_6471,N_6269,N_6283);
or U6472 (N_6472,N_6302,N_6276);
and U6473 (N_6473,N_6338,N_6363);
xor U6474 (N_6474,N_6320,N_6278);
or U6475 (N_6475,N_6292,N_6296);
nor U6476 (N_6476,N_6251,N_6322);
and U6477 (N_6477,N_6276,N_6252);
nand U6478 (N_6478,N_6274,N_6358);
nor U6479 (N_6479,N_6258,N_6339);
nor U6480 (N_6480,N_6309,N_6356);
or U6481 (N_6481,N_6301,N_6340);
or U6482 (N_6482,N_6343,N_6287);
or U6483 (N_6483,N_6340,N_6323);
nor U6484 (N_6484,N_6252,N_6331);
and U6485 (N_6485,N_6354,N_6345);
nor U6486 (N_6486,N_6328,N_6304);
nand U6487 (N_6487,N_6337,N_6299);
nand U6488 (N_6488,N_6338,N_6306);
or U6489 (N_6489,N_6275,N_6339);
or U6490 (N_6490,N_6298,N_6366);
nand U6491 (N_6491,N_6295,N_6290);
nor U6492 (N_6492,N_6322,N_6333);
nor U6493 (N_6493,N_6308,N_6268);
nand U6494 (N_6494,N_6363,N_6346);
xnor U6495 (N_6495,N_6297,N_6302);
or U6496 (N_6496,N_6343,N_6294);
and U6497 (N_6497,N_6361,N_6370);
xor U6498 (N_6498,N_6301,N_6371);
nand U6499 (N_6499,N_6314,N_6336);
or U6500 (N_6500,N_6474,N_6460);
nand U6501 (N_6501,N_6454,N_6422);
nand U6502 (N_6502,N_6472,N_6485);
nor U6503 (N_6503,N_6420,N_6493);
or U6504 (N_6504,N_6496,N_6428);
nand U6505 (N_6505,N_6494,N_6467);
nor U6506 (N_6506,N_6421,N_6383);
nor U6507 (N_6507,N_6488,N_6405);
xor U6508 (N_6508,N_6430,N_6378);
xnor U6509 (N_6509,N_6436,N_6492);
and U6510 (N_6510,N_6412,N_6448);
xor U6511 (N_6511,N_6487,N_6478);
xor U6512 (N_6512,N_6377,N_6469);
nand U6513 (N_6513,N_6482,N_6431);
nor U6514 (N_6514,N_6416,N_6379);
xnor U6515 (N_6515,N_6388,N_6423);
nand U6516 (N_6516,N_6476,N_6499);
and U6517 (N_6517,N_6429,N_6434);
or U6518 (N_6518,N_6400,N_6380);
nand U6519 (N_6519,N_6425,N_6393);
nand U6520 (N_6520,N_6387,N_6450);
and U6521 (N_6521,N_6444,N_6375);
and U6522 (N_6522,N_6468,N_6435);
and U6523 (N_6523,N_6451,N_6401);
and U6524 (N_6524,N_6403,N_6402);
or U6525 (N_6525,N_6465,N_6437);
xor U6526 (N_6526,N_6470,N_6489);
and U6527 (N_6527,N_6433,N_6479);
and U6528 (N_6528,N_6490,N_6381);
or U6529 (N_6529,N_6376,N_6386);
nor U6530 (N_6530,N_6417,N_6418);
and U6531 (N_6531,N_6458,N_6457);
or U6532 (N_6532,N_6419,N_6447);
nand U6533 (N_6533,N_6453,N_6424);
and U6534 (N_6534,N_6389,N_6473);
or U6535 (N_6535,N_6475,N_6456);
xnor U6536 (N_6536,N_6396,N_6439);
nand U6537 (N_6537,N_6399,N_6446);
or U6538 (N_6538,N_6477,N_6427);
nand U6539 (N_6539,N_6462,N_6440);
nand U6540 (N_6540,N_6449,N_6415);
or U6541 (N_6541,N_6414,N_6394);
or U6542 (N_6542,N_6471,N_6459);
nor U6543 (N_6543,N_6486,N_6407);
nor U6544 (N_6544,N_6455,N_6438);
and U6545 (N_6545,N_6480,N_6398);
and U6546 (N_6546,N_6445,N_6413);
nor U6547 (N_6547,N_6404,N_6411);
nand U6548 (N_6548,N_6481,N_6384);
xor U6549 (N_6549,N_6410,N_6464);
nand U6550 (N_6550,N_6441,N_6391);
or U6551 (N_6551,N_6491,N_6390);
xor U6552 (N_6552,N_6443,N_6409);
nand U6553 (N_6553,N_6483,N_6432);
nor U6554 (N_6554,N_6461,N_6466);
and U6555 (N_6555,N_6463,N_6397);
or U6556 (N_6556,N_6406,N_6484);
nand U6557 (N_6557,N_6382,N_6498);
nand U6558 (N_6558,N_6497,N_6452);
nor U6559 (N_6559,N_6408,N_6442);
and U6560 (N_6560,N_6495,N_6426);
nor U6561 (N_6561,N_6392,N_6395);
xnor U6562 (N_6562,N_6385,N_6401);
nand U6563 (N_6563,N_6461,N_6442);
nand U6564 (N_6564,N_6430,N_6413);
xor U6565 (N_6565,N_6404,N_6481);
xnor U6566 (N_6566,N_6432,N_6454);
or U6567 (N_6567,N_6483,N_6382);
nor U6568 (N_6568,N_6498,N_6474);
xnor U6569 (N_6569,N_6419,N_6448);
and U6570 (N_6570,N_6431,N_6424);
and U6571 (N_6571,N_6436,N_6403);
or U6572 (N_6572,N_6413,N_6401);
xnor U6573 (N_6573,N_6435,N_6445);
nor U6574 (N_6574,N_6459,N_6408);
and U6575 (N_6575,N_6481,N_6458);
nand U6576 (N_6576,N_6484,N_6408);
or U6577 (N_6577,N_6467,N_6403);
xnor U6578 (N_6578,N_6419,N_6486);
xnor U6579 (N_6579,N_6377,N_6430);
nor U6580 (N_6580,N_6384,N_6441);
nor U6581 (N_6581,N_6426,N_6380);
or U6582 (N_6582,N_6410,N_6425);
nor U6583 (N_6583,N_6456,N_6495);
nor U6584 (N_6584,N_6446,N_6493);
nor U6585 (N_6585,N_6391,N_6473);
nor U6586 (N_6586,N_6404,N_6445);
nand U6587 (N_6587,N_6492,N_6386);
or U6588 (N_6588,N_6487,N_6496);
nor U6589 (N_6589,N_6377,N_6387);
or U6590 (N_6590,N_6479,N_6446);
xor U6591 (N_6591,N_6403,N_6445);
nor U6592 (N_6592,N_6401,N_6375);
nand U6593 (N_6593,N_6417,N_6475);
xnor U6594 (N_6594,N_6488,N_6494);
nor U6595 (N_6595,N_6476,N_6415);
xor U6596 (N_6596,N_6404,N_6383);
or U6597 (N_6597,N_6441,N_6419);
xnor U6598 (N_6598,N_6375,N_6450);
nor U6599 (N_6599,N_6386,N_6411);
nand U6600 (N_6600,N_6396,N_6400);
or U6601 (N_6601,N_6402,N_6463);
and U6602 (N_6602,N_6495,N_6465);
nor U6603 (N_6603,N_6464,N_6499);
or U6604 (N_6604,N_6442,N_6472);
xnor U6605 (N_6605,N_6487,N_6493);
nor U6606 (N_6606,N_6390,N_6471);
xor U6607 (N_6607,N_6407,N_6412);
or U6608 (N_6608,N_6402,N_6449);
and U6609 (N_6609,N_6489,N_6464);
nor U6610 (N_6610,N_6441,N_6458);
nor U6611 (N_6611,N_6431,N_6401);
xnor U6612 (N_6612,N_6482,N_6419);
and U6613 (N_6613,N_6479,N_6447);
xor U6614 (N_6614,N_6498,N_6384);
nand U6615 (N_6615,N_6456,N_6410);
and U6616 (N_6616,N_6420,N_6378);
nor U6617 (N_6617,N_6381,N_6477);
and U6618 (N_6618,N_6496,N_6448);
nor U6619 (N_6619,N_6499,N_6483);
nand U6620 (N_6620,N_6391,N_6485);
nand U6621 (N_6621,N_6410,N_6412);
nand U6622 (N_6622,N_6456,N_6402);
and U6623 (N_6623,N_6380,N_6375);
or U6624 (N_6624,N_6391,N_6420);
nand U6625 (N_6625,N_6536,N_6612);
or U6626 (N_6626,N_6556,N_6515);
and U6627 (N_6627,N_6553,N_6604);
and U6628 (N_6628,N_6551,N_6514);
or U6629 (N_6629,N_6535,N_6573);
and U6630 (N_6630,N_6571,N_6577);
xor U6631 (N_6631,N_6575,N_6505);
nor U6632 (N_6632,N_6516,N_6528);
nand U6633 (N_6633,N_6507,N_6506);
xnor U6634 (N_6634,N_6605,N_6579);
xnor U6635 (N_6635,N_6576,N_6592);
or U6636 (N_6636,N_6568,N_6513);
nand U6637 (N_6637,N_6615,N_6623);
or U6638 (N_6638,N_6527,N_6531);
or U6639 (N_6639,N_6508,N_6520);
nor U6640 (N_6640,N_6569,N_6583);
xnor U6641 (N_6641,N_6564,N_6590);
nand U6642 (N_6642,N_6501,N_6606);
and U6643 (N_6643,N_6619,N_6584);
or U6644 (N_6644,N_6522,N_6512);
xor U6645 (N_6645,N_6563,N_6600);
nand U6646 (N_6646,N_6578,N_6610);
xnor U6647 (N_6647,N_6529,N_6599);
or U6648 (N_6648,N_6601,N_6596);
nand U6649 (N_6649,N_6617,N_6549);
and U6650 (N_6650,N_6591,N_6503);
or U6651 (N_6651,N_6609,N_6543);
xnor U6652 (N_6652,N_6521,N_6618);
xnor U6653 (N_6653,N_6539,N_6594);
nand U6654 (N_6654,N_6525,N_6541);
and U6655 (N_6655,N_6552,N_6622);
and U6656 (N_6656,N_6587,N_6544);
and U6657 (N_6657,N_6614,N_6566);
nor U6658 (N_6658,N_6580,N_6585);
and U6659 (N_6659,N_6545,N_6582);
nor U6660 (N_6660,N_6547,N_6616);
nor U6661 (N_6661,N_6524,N_6532);
xnor U6662 (N_6662,N_6546,N_6542);
nand U6663 (N_6663,N_6523,N_6603);
nand U6664 (N_6664,N_6509,N_6562);
nor U6665 (N_6665,N_6519,N_6611);
and U6666 (N_6666,N_6560,N_6565);
nor U6667 (N_6667,N_6602,N_6589);
nand U6668 (N_6668,N_6559,N_6593);
and U6669 (N_6669,N_6561,N_6540);
or U6670 (N_6670,N_6530,N_6624);
or U6671 (N_6671,N_6613,N_6534);
nor U6672 (N_6672,N_6518,N_6554);
or U6673 (N_6673,N_6567,N_6607);
and U6674 (N_6674,N_6500,N_6550);
or U6675 (N_6675,N_6510,N_6511);
or U6676 (N_6676,N_6570,N_6526);
and U6677 (N_6677,N_6574,N_6620);
nor U6678 (N_6678,N_6621,N_6533);
nand U6679 (N_6679,N_6538,N_6588);
and U6680 (N_6680,N_6548,N_6504);
or U6681 (N_6681,N_6555,N_6557);
nor U6682 (N_6682,N_6608,N_6595);
nand U6683 (N_6683,N_6598,N_6597);
xor U6684 (N_6684,N_6517,N_6581);
xor U6685 (N_6685,N_6537,N_6586);
or U6686 (N_6686,N_6558,N_6572);
and U6687 (N_6687,N_6502,N_6612);
nand U6688 (N_6688,N_6577,N_6543);
or U6689 (N_6689,N_6510,N_6503);
xor U6690 (N_6690,N_6514,N_6506);
or U6691 (N_6691,N_6540,N_6520);
xor U6692 (N_6692,N_6506,N_6609);
and U6693 (N_6693,N_6536,N_6590);
and U6694 (N_6694,N_6563,N_6556);
or U6695 (N_6695,N_6588,N_6598);
nand U6696 (N_6696,N_6601,N_6513);
and U6697 (N_6697,N_6504,N_6524);
or U6698 (N_6698,N_6614,N_6617);
or U6699 (N_6699,N_6531,N_6538);
nor U6700 (N_6700,N_6519,N_6501);
and U6701 (N_6701,N_6621,N_6605);
and U6702 (N_6702,N_6548,N_6553);
nor U6703 (N_6703,N_6551,N_6540);
or U6704 (N_6704,N_6507,N_6511);
nor U6705 (N_6705,N_6596,N_6534);
nor U6706 (N_6706,N_6512,N_6620);
nand U6707 (N_6707,N_6589,N_6600);
xnor U6708 (N_6708,N_6609,N_6533);
and U6709 (N_6709,N_6571,N_6582);
nor U6710 (N_6710,N_6566,N_6586);
nand U6711 (N_6711,N_6548,N_6574);
nor U6712 (N_6712,N_6533,N_6618);
nor U6713 (N_6713,N_6592,N_6620);
and U6714 (N_6714,N_6505,N_6601);
nor U6715 (N_6715,N_6589,N_6620);
xnor U6716 (N_6716,N_6550,N_6507);
and U6717 (N_6717,N_6617,N_6575);
and U6718 (N_6718,N_6591,N_6587);
and U6719 (N_6719,N_6502,N_6504);
nor U6720 (N_6720,N_6529,N_6623);
xnor U6721 (N_6721,N_6618,N_6513);
nand U6722 (N_6722,N_6529,N_6541);
xor U6723 (N_6723,N_6609,N_6555);
or U6724 (N_6724,N_6546,N_6596);
or U6725 (N_6725,N_6587,N_6577);
or U6726 (N_6726,N_6622,N_6506);
nand U6727 (N_6727,N_6605,N_6546);
xor U6728 (N_6728,N_6563,N_6502);
nor U6729 (N_6729,N_6507,N_6577);
nand U6730 (N_6730,N_6514,N_6535);
or U6731 (N_6731,N_6605,N_6612);
and U6732 (N_6732,N_6521,N_6611);
nand U6733 (N_6733,N_6576,N_6559);
xor U6734 (N_6734,N_6549,N_6506);
nor U6735 (N_6735,N_6525,N_6551);
xor U6736 (N_6736,N_6516,N_6549);
and U6737 (N_6737,N_6545,N_6565);
nor U6738 (N_6738,N_6562,N_6521);
or U6739 (N_6739,N_6541,N_6600);
nand U6740 (N_6740,N_6546,N_6615);
nand U6741 (N_6741,N_6599,N_6504);
nor U6742 (N_6742,N_6507,N_6501);
nand U6743 (N_6743,N_6605,N_6542);
xor U6744 (N_6744,N_6585,N_6609);
or U6745 (N_6745,N_6609,N_6607);
and U6746 (N_6746,N_6595,N_6611);
and U6747 (N_6747,N_6620,N_6507);
xor U6748 (N_6748,N_6607,N_6528);
xor U6749 (N_6749,N_6580,N_6554);
nor U6750 (N_6750,N_6635,N_6684);
and U6751 (N_6751,N_6652,N_6690);
or U6752 (N_6752,N_6714,N_6749);
nand U6753 (N_6753,N_6718,N_6683);
nor U6754 (N_6754,N_6729,N_6738);
nand U6755 (N_6755,N_6630,N_6726);
xnor U6756 (N_6756,N_6672,N_6703);
and U6757 (N_6757,N_6731,N_6691);
nor U6758 (N_6758,N_6686,N_6737);
or U6759 (N_6759,N_6694,N_6735);
nor U6760 (N_6760,N_6700,N_6657);
nand U6761 (N_6761,N_6695,N_6648);
or U6762 (N_6762,N_6677,N_6634);
or U6763 (N_6763,N_6633,N_6654);
or U6764 (N_6764,N_6734,N_6706);
nand U6765 (N_6765,N_6681,N_6643);
or U6766 (N_6766,N_6650,N_6644);
xnor U6767 (N_6767,N_6716,N_6748);
xor U6768 (N_6768,N_6712,N_6640);
and U6769 (N_6769,N_6745,N_6670);
nor U6770 (N_6770,N_6709,N_6717);
or U6771 (N_6771,N_6708,N_6741);
nor U6772 (N_6772,N_6675,N_6722);
and U6773 (N_6773,N_6639,N_6730);
and U6774 (N_6774,N_6646,N_6636);
nor U6775 (N_6775,N_6711,N_6649);
nand U6776 (N_6776,N_6698,N_6705);
nand U6777 (N_6777,N_6638,N_6732);
xor U6778 (N_6778,N_6723,N_6693);
nor U6779 (N_6779,N_6701,N_6663);
nand U6780 (N_6780,N_6653,N_6673);
xor U6781 (N_6781,N_6727,N_6627);
and U6782 (N_6782,N_6674,N_6728);
and U6783 (N_6783,N_6720,N_6661);
or U6784 (N_6784,N_6721,N_6739);
nand U6785 (N_6785,N_6626,N_6656);
nand U6786 (N_6786,N_6697,N_6687);
or U6787 (N_6787,N_6746,N_6665);
and U6788 (N_6788,N_6733,N_6667);
nor U6789 (N_6789,N_6660,N_6680);
xnor U6790 (N_6790,N_6689,N_6668);
nand U6791 (N_6791,N_6724,N_6664);
or U6792 (N_6792,N_6736,N_6671);
nor U6793 (N_6793,N_6651,N_6628);
xor U6794 (N_6794,N_6744,N_6715);
nor U6795 (N_6795,N_6692,N_6740);
nor U6796 (N_6796,N_6662,N_6713);
or U6797 (N_6797,N_6637,N_6659);
or U6798 (N_6798,N_6647,N_6702);
and U6799 (N_6799,N_6625,N_6696);
or U6800 (N_6800,N_6743,N_6699);
xor U6801 (N_6801,N_6645,N_6704);
xnor U6802 (N_6802,N_6742,N_6629);
and U6803 (N_6803,N_6666,N_6707);
xor U6804 (N_6804,N_6642,N_6679);
xnor U6805 (N_6805,N_6747,N_6719);
or U6806 (N_6806,N_6655,N_6682);
nand U6807 (N_6807,N_6710,N_6631);
or U6808 (N_6808,N_6678,N_6658);
nor U6809 (N_6809,N_6632,N_6676);
xnor U6810 (N_6810,N_6669,N_6685);
and U6811 (N_6811,N_6641,N_6725);
nand U6812 (N_6812,N_6688,N_6717);
or U6813 (N_6813,N_6676,N_6703);
or U6814 (N_6814,N_6712,N_6727);
or U6815 (N_6815,N_6680,N_6645);
or U6816 (N_6816,N_6632,N_6708);
and U6817 (N_6817,N_6743,N_6658);
nor U6818 (N_6818,N_6641,N_6682);
and U6819 (N_6819,N_6745,N_6632);
or U6820 (N_6820,N_6685,N_6645);
and U6821 (N_6821,N_6739,N_6695);
nor U6822 (N_6822,N_6644,N_6721);
and U6823 (N_6823,N_6743,N_6668);
xor U6824 (N_6824,N_6676,N_6662);
and U6825 (N_6825,N_6684,N_6666);
xor U6826 (N_6826,N_6719,N_6746);
nand U6827 (N_6827,N_6731,N_6644);
nor U6828 (N_6828,N_6688,N_6673);
or U6829 (N_6829,N_6651,N_6626);
or U6830 (N_6830,N_6676,N_6712);
or U6831 (N_6831,N_6663,N_6672);
and U6832 (N_6832,N_6684,N_6694);
or U6833 (N_6833,N_6680,N_6714);
nor U6834 (N_6834,N_6662,N_6740);
and U6835 (N_6835,N_6681,N_6653);
or U6836 (N_6836,N_6668,N_6659);
xnor U6837 (N_6837,N_6719,N_6666);
nor U6838 (N_6838,N_6655,N_6727);
or U6839 (N_6839,N_6636,N_6644);
xor U6840 (N_6840,N_6685,N_6663);
xnor U6841 (N_6841,N_6664,N_6635);
or U6842 (N_6842,N_6641,N_6686);
and U6843 (N_6843,N_6649,N_6724);
and U6844 (N_6844,N_6739,N_6669);
or U6845 (N_6845,N_6654,N_6641);
or U6846 (N_6846,N_6732,N_6663);
or U6847 (N_6847,N_6660,N_6626);
nor U6848 (N_6848,N_6726,N_6700);
nand U6849 (N_6849,N_6626,N_6735);
or U6850 (N_6850,N_6719,N_6652);
and U6851 (N_6851,N_6686,N_6716);
nand U6852 (N_6852,N_6712,N_6669);
xnor U6853 (N_6853,N_6682,N_6667);
xor U6854 (N_6854,N_6639,N_6679);
nand U6855 (N_6855,N_6747,N_6636);
and U6856 (N_6856,N_6739,N_6704);
and U6857 (N_6857,N_6666,N_6674);
or U6858 (N_6858,N_6677,N_6741);
or U6859 (N_6859,N_6711,N_6646);
nand U6860 (N_6860,N_6678,N_6661);
xnor U6861 (N_6861,N_6726,N_6665);
nand U6862 (N_6862,N_6695,N_6626);
and U6863 (N_6863,N_6688,N_6719);
and U6864 (N_6864,N_6683,N_6681);
xnor U6865 (N_6865,N_6672,N_6656);
xnor U6866 (N_6866,N_6680,N_6671);
or U6867 (N_6867,N_6682,N_6658);
and U6868 (N_6868,N_6731,N_6687);
nor U6869 (N_6869,N_6652,N_6676);
nand U6870 (N_6870,N_6629,N_6685);
or U6871 (N_6871,N_6679,N_6705);
or U6872 (N_6872,N_6681,N_6742);
nor U6873 (N_6873,N_6700,N_6649);
xnor U6874 (N_6874,N_6682,N_6625);
nor U6875 (N_6875,N_6863,N_6822);
nor U6876 (N_6876,N_6793,N_6859);
and U6877 (N_6877,N_6838,N_6766);
or U6878 (N_6878,N_6765,N_6811);
nor U6879 (N_6879,N_6824,N_6841);
and U6880 (N_6880,N_6812,N_6825);
xor U6881 (N_6881,N_6855,N_6873);
or U6882 (N_6882,N_6817,N_6809);
xor U6883 (N_6883,N_6844,N_6827);
nor U6884 (N_6884,N_6795,N_6796);
nand U6885 (N_6885,N_6770,N_6871);
nor U6886 (N_6886,N_6816,N_6804);
or U6887 (N_6887,N_6759,N_6798);
and U6888 (N_6888,N_6854,N_6790);
and U6889 (N_6889,N_6784,N_6763);
xor U6890 (N_6890,N_6806,N_6828);
and U6891 (N_6891,N_6752,N_6836);
or U6892 (N_6892,N_6820,N_6788);
nand U6893 (N_6893,N_6778,N_6842);
or U6894 (N_6894,N_6857,N_6802);
nor U6895 (N_6895,N_6847,N_6858);
xor U6896 (N_6896,N_6794,N_6768);
nor U6897 (N_6897,N_6799,N_6769);
nand U6898 (N_6898,N_6818,N_6754);
and U6899 (N_6899,N_6755,N_6792);
or U6900 (N_6900,N_6864,N_6753);
and U6901 (N_6901,N_6865,N_6815);
and U6902 (N_6902,N_6803,N_6814);
nand U6903 (N_6903,N_6772,N_6868);
xnor U6904 (N_6904,N_6761,N_6808);
and U6905 (N_6905,N_6779,N_6774);
or U6906 (N_6906,N_6810,N_6830);
nand U6907 (N_6907,N_6800,N_6831);
and U6908 (N_6908,N_6758,N_6805);
xnor U6909 (N_6909,N_6839,N_6807);
and U6910 (N_6910,N_6869,N_6843);
nor U6911 (N_6911,N_6787,N_6776);
xnor U6912 (N_6912,N_6837,N_6849);
and U6913 (N_6913,N_6853,N_6781);
nor U6914 (N_6914,N_6823,N_6777);
nand U6915 (N_6915,N_6835,N_6861);
xnor U6916 (N_6916,N_6832,N_6767);
nor U6917 (N_6917,N_6821,N_6826);
or U6918 (N_6918,N_6860,N_6764);
nand U6919 (N_6919,N_6756,N_6862);
xor U6920 (N_6920,N_6872,N_6780);
and U6921 (N_6921,N_6813,N_6870);
and U6922 (N_6922,N_6782,N_6833);
nor U6923 (N_6923,N_6773,N_6852);
nand U6924 (N_6924,N_6750,N_6845);
or U6925 (N_6925,N_6775,N_6762);
or U6926 (N_6926,N_6829,N_6783);
nand U6927 (N_6927,N_6846,N_6866);
xor U6928 (N_6928,N_6819,N_6840);
xnor U6929 (N_6929,N_6785,N_6789);
xnor U6930 (N_6930,N_6850,N_6851);
and U6931 (N_6931,N_6786,N_6751);
nor U6932 (N_6932,N_6867,N_6757);
nand U6933 (N_6933,N_6791,N_6797);
or U6934 (N_6934,N_6760,N_6801);
nand U6935 (N_6935,N_6771,N_6848);
nor U6936 (N_6936,N_6874,N_6834);
or U6937 (N_6937,N_6856,N_6865);
and U6938 (N_6938,N_6768,N_6868);
and U6939 (N_6939,N_6752,N_6763);
nor U6940 (N_6940,N_6806,N_6764);
and U6941 (N_6941,N_6777,N_6798);
nor U6942 (N_6942,N_6809,N_6833);
xnor U6943 (N_6943,N_6852,N_6842);
xnor U6944 (N_6944,N_6851,N_6825);
nor U6945 (N_6945,N_6833,N_6844);
and U6946 (N_6946,N_6861,N_6752);
nor U6947 (N_6947,N_6786,N_6753);
xnor U6948 (N_6948,N_6868,N_6779);
and U6949 (N_6949,N_6761,N_6804);
nor U6950 (N_6950,N_6772,N_6851);
and U6951 (N_6951,N_6765,N_6827);
nand U6952 (N_6952,N_6806,N_6793);
nor U6953 (N_6953,N_6813,N_6793);
xnor U6954 (N_6954,N_6817,N_6778);
and U6955 (N_6955,N_6860,N_6771);
or U6956 (N_6956,N_6781,N_6796);
or U6957 (N_6957,N_6765,N_6866);
xnor U6958 (N_6958,N_6868,N_6871);
or U6959 (N_6959,N_6752,N_6862);
nand U6960 (N_6960,N_6865,N_6853);
nand U6961 (N_6961,N_6854,N_6850);
xor U6962 (N_6962,N_6799,N_6871);
nor U6963 (N_6963,N_6793,N_6848);
nor U6964 (N_6964,N_6807,N_6833);
or U6965 (N_6965,N_6805,N_6808);
nand U6966 (N_6966,N_6796,N_6841);
xor U6967 (N_6967,N_6837,N_6800);
nor U6968 (N_6968,N_6761,N_6758);
nand U6969 (N_6969,N_6820,N_6850);
or U6970 (N_6970,N_6861,N_6778);
nand U6971 (N_6971,N_6853,N_6822);
xor U6972 (N_6972,N_6797,N_6772);
or U6973 (N_6973,N_6818,N_6761);
nor U6974 (N_6974,N_6812,N_6873);
and U6975 (N_6975,N_6855,N_6825);
nand U6976 (N_6976,N_6862,N_6775);
and U6977 (N_6977,N_6758,N_6830);
and U6978 (N_6978,N_6874,N_6847);
xnor U6979 (N_6979,N_6766,N_6855);
nand U6980 (N_6980,N_6787,N_6826);
nor U6981 (N_6981,N_6788,N_6818);
nor U6982 (N_6982,N_6800,N_6785);
or U6983 (N_6983,N_6762,N_6853);
nor U6984 (N_6984,N_6810,N_6782);
and U6985 (N_6985,N_6822,N_6845);
or U6986 (N_6986,N_6853,N_6830);
or U6987 (N_6987,N_6848,N_6812);
nor U6988 (N_6988,N_6752,N_6799);
and U6989 (N_6989,N_6811,N_6837);
and U6990 (N_6990,N_6790,N_6769);
xnor U6991 (N_6991,N_6826,N_6846);
nor U6992 (N_6992,N_6834,N_6838);
or U6993 (N_6993,N_6837,N_6792);
and U6994 (N_6994,N_6782,N_6859);
or U6995 (N_6995,N_6769,N_6766);
nand U6996 (N_6996,N_6782,N_6808);
and U6997 (N_6997,N_6808,N_6751);
or U6998 (N_6998,N_6855,N_6834);
xor U6999 (N_6999,N_6765,N_6772);
nand U7000 (N_7000,N_6902,N_6962);
or U7001 (N_7001,N_6963,N_6970);
and U7002 (N_7002,N_6882,N_6913);
nor U7003 (N_7003,N_6960,N_6928);
and U7004 (N_7004,N_6938,N_6885);
xor U7005 (N_7005,N_6978,N_6896);
nand U7006 (N_7006,N_6971,N_6922);
nand U7007 (N_7007,N_6966,N_6911);
xor U7008 (N_7008,N_6967,N_6876);
or U7009 (N_7009,N_6988,N_6879);
or U7010 (N_7010,N_6916,N_6976);
and U7011 (N_7011,N_6893,N_6886);
nand U7012 (N_7012,N_6908,N_6969);
xnor U7013 (N_7013,N_6974,N_6888);
xor U7014 (N_7014,N_6891,N_6946);
xnor U7015 (N_7015,N_6989,N_6941);
and U7016 (N_7016,N_6926,N_6880);
or U7017 (N_7017,N_6956,N_6952);
xnor U7018 (N_7018,N_6972,N_6955);
and U7019 (N_7019,N_6982,N_6901);
xor U7020 (N_7020,N_6918,N_6930);
and U7021 (N_7021,N_6954,N_6914);
nor U7022 (N_7022,N_6991,N_6894);
xor U7023 (N_7023,N_6947,N_6986);
nor U7024 (N_7024,N_6987,N_6968);
and U7025 (N_7025,N_6927,N_6973);
and U7026 (N_7026,N_6898,N_6921);
or U7027 (N_7027,N_6899,N_6881);
nor U7028 (N_7028,N_6897,N_6957);
nor U7029 (N_7029,N_6999,N_6985);
nand U7030 (N_7030,N_6895,N_6951);
and U7031 (N_7031,N_6905,N_6917);
xnor U7032 (N_7032,N_6904,N_6981);
nand U7033 (N_7033,N_6934,N_6915);
or U7034 (N_7034,N_6933,N_6984);
nand U7035 (N_7035,N_6920,N_6937);
nand U7036 (N_7036,N_6936,N_6995);
nor U7037 (N_7037,N_6909,N_6959);
and U7038 (N_7038,N_6889,N_6939);
xor U7039 (N_7039,N_6932,N_6950);
xor U7040 (N_7040,N_6878,N_6929);
nand U7041 (N_7041,N_6983,N_6977);
nand U7042 (N_7042,N_6925,N_6912);
nor U7043 (N_7043,N_6924,N_6900);
or U7044 (N_7044,N_6953,N_6919);
nor U7045 (N_7045,N_6884,N_6883);
nand U7046 (N_7046,N_6980,N_6945);
xor U7047 (N_7047,N_6875,N_6993);
or U7048 (N_7048,N_6958,N_6990);
nand U7049 (N_7049,N_6979,N_6890);
nand U7050 (N_7050,N_6877,N_6910);
or U7051 (N_7051,N_6903,N_6994);
nor U7052 (N_7052,N_6949,N_6923);
or U7053 (N_7053,N_6998,N_6943);
and U7054 (N_7054,N_6948,N_6935);
or U7055 (N_7055,N_6906,N_6940);
nor U7056 (N_7056,N_6964,N_6975);
nor U7057 (N_7057,N_6944,N_6992);
nand U7058 (N_7058,N_6965,N_6997);
and U7059 (N_7059,N_6907,N_6892);
nor U7060 (N_7060,N_6887,N_6942);
xnor U7061 (N_7061,N_6961,N_6931);
and U7062 (N_7062,N_6996,N_6961);
nor U7063 (N_7063,N_6884,N_6926);
nand U7064 (N_7064,N_6912,N_6884);
nand U7065 (N_7065,N_6941,N_6878);
nand U7066 (N_7066,N_6889,N_6975);
nor U7067 (N_7067,N_6909,N_6897);
nand U7068 (N_7068,N_6956,N_6881);
or U7069 (N_7069,N_6979,N_6959);
nor U7070 (N_7070,N_6880,N_6894);
or U7071 (N_7071,N_6900,N_6943);
xnor U7072 (N_7072,N_6991,N_6967);
nand U7073 (N_7073,N_6880,N_6955);
and U7074 (N_7074,N_6885,N_6928);
and U7075 (N_7075,N_6949,N_6957);
and U7076 (N_7076,N_6985,N_6933);
nor U7077 (N_7077,N_6875,N_6907);
or U7078 (N_7078,N_6887,N_6926);
or U7079 (N_7079,N_6977,N_6978);
or U7080 (N_7080,N_6882,N_6943);
and U7081 (N_7081,N_6936,N_6978);
nor U7082 (N_7082,N_6961,N_6904);
and U7083 (N_7083,N_6958,N_6968);
nand U7084 (N_7084,N_6928,N_6917);
and U7085 (N_7085,N_6907,N_6978);
xnor U7086 (N_7086,N_6885,N_6994);
and U7087 (N_7087,N_6897,N_6898);
nand U7088 (N_7088,N_6958,N_6890);
nor U7089 (N_7089,N_6905,N_6947);
xor U7090 (N_7090,N_6974,N_6909);
and U7091 (N_7091,N_6931,N_6963);
nor U7092 (N_7092,N_6921,N_6935);
nand U7093 (N_7093,N_6933,N_6960);
nor U7094 (N_7094,N_6985,N_6908);
nand U7095 (N_7095,N_6915,N_6931);
nand U7096 (N_7096,N_6880,N_6899);
or U7097 (N_7097,N_6929,N_6995);
nand U7098 (N_7098,N_6979,N_6926);
and U7099 (N_7099,N_6946,N_6950);
and U7100 (N_7100,N_6908,N_6934);
or U7101 (N_7101,N_6935,N_6950);
or U7102 (N_7102,N_6919,N_6880);
xor U7103 (N_7103,N_6888,N_6928);
nor U7104 (N_7104,N_6952,N_6887);
nor U7105 (N_7105,N_6913,N_6991);
or U7106 (N_7106,N_6929,N_6899);
nand U7107 (N_7107,N_6990,N_6995);
nor U7108 (N_7108,N_6938,N_6918);
and U7109 (N_7109,N_6972,N_6943);
xnor U7110 (N_7110,N_6888,N_6953);
nor U7111 (N_7111,N_6890,N_6906);
nor U7112 (N_7112,N_6945,N_6904);
nor U7113 (N_7113,N_6968,N_6879);
or U7114 (N_7114,N_6995,N_6967);
and U7115 (N_7115,N_6947,N_6998);
nor U7116 (N_7116,N_6923,N_6996);
nor U7117 (N_7117,N_6938,N_6990);
and U7118 (N_7118,N_6958,N_6942);
xor U7119 (N_7119,N_6912,N_6992);
nand U7120 (N_7120,N_6963,N_6992);
xor U7121 (N_7121,N_6994,N_6894);
xnor U7122 (N_7122,N_6996,N_6998);
and U7123 (N_7123,N_6902,N_6994);
nand U7124 (N_7124,N_6998,N_6904);
or U7125 (N_7125,N_7022,N_7015);
xnor U7126 (N_7126,N_7045,N_7097);
nor U7127 (N_7127,N_7079,N_7041);
and U7128 (N_7128,N_7069,N_7007);
nand U7129 (N_7129,N_7013,N_7046);
nor U7130 (N_7130,N_7080,N_7032);
nand U7131 (N_7131,N_7093,N_7063);
nor U7132 (N_7132,N_7017,N_7123);
or U7133 (N_7133,N_7028,N_7116);
or U7134 (N_7134,N_7121,N_7065);
or U7135 (N_7135,N_7039,N_7003);
nor U7136 (N_7136,N_7082,N_7095);
and U7137 (N_7137,N_7010,N_7107);
nand U7138 (N_7138,N_7112,N_7070);
nor U7139 (N_7139,N_7076,N_7056);
nand U7140 (N_7140,N_7077,N_7086);
or U7141 (N_7141,N_7072,N_7040);
nand U7142 (N_7142,N_7043,N_7057);
xnor U7143 (N_7143,N_7081,N_7052);
and U7144 (N_7144,N_7011,N_7026);
and U7145 (N_7145,N_7088,N_7113);
xnor U7146 (N_7146,N_7025,N_7060);
xnor U7147 (N_7147,N_7005,N_7037);
nand U7148 (N_7148,N_7050,N_7034);
nand U7149 (N_7149,N_7085,N_7038);
xor U7150 (N_7150,N_7094,N_7006);
or U7151 (N_7151,N_7104,N_7115);
nor U7152 (N_7152,N_7118,N_7018);
nand U7153 (N_7153,N_7103,N_7000);
nand U7154 (N_7154,N_7117,N_7049);
and U7155 (N_7155,N_7111,N_7058);
nor U7156 (N_7156,N_7098,N_7092);
nand U7157 (N_7157,N_7091,N_7089);
or U7158 (N_7158,N_7024,N_7055);
xnor U7159 (N_7159,N_7108,N_7071);
nand U7160 (N_7160,N_7009,N_7023);
nand U7161 (N_7161,N_7110,N_7067);
and U7162 (N_7162,N_7062,N_7096);
nor U7163 (N_7163,N_7073,N_7090);
and U7164 (N_7164,N_7083,N_7031);
nor U7165 (N_7165,N_7099,N_7106);
or U7166 (N_7166,N_7033,N_7059);
or U7167 (N_7167,N_7048,N_7087);
nor U7168 (N_7168,N_7102,N_7074);
nand U7169 (N_7169,N_7044,N_7029);
or U7170 (N_7170,N_7051,N_7066);
nand U7171 (N_7171,N_7068,N_7109);
nor U7172 (N_7172,N_7035,N_7054);
or U7173 (N_7173,N_7001,N_7061);
and U7174 (N_7174,N_7019,N_7030);
or U7175 (N_7175,N_7027,N_7053);
xor U7176 (N_7176,N_7084,N_7014);
and U7177 (N_7177,N_7075,N_7002);
and U7178 (N_7178,N_7122,N_7047);
or U7179 (N_7179,N_7119,N_7016);
xor U7180 (N_7180,N_7004,N_7021);
nand U7181 (N_7181,N_7078,N_7120);
xor U7182 (N_7182,N_7008,N_7124);
nand U7183 (N_7183,N_7114,N_7100);
nor U7184 (N_7184,N_7064,N_7012);
xor U7185 (N_7185,N_7020,N_7042);
or U7186 (N_7186,N_7101,N_7036);
or U7187 (N_7187,N_7105,N_7010);
xor U7188 (N_7188,N_7025,N_7107);
nor U7189 (N_7189,N_7005,N_7050);
nor U7190 (N_7190,N_7067,N_7022);
or U7191 (N_7191,N_7055,N_7067);
nand U7192 (N_7192,N_7103,N_7112);
and U7193 (N_7193,N_7087,N_7091);
and U7194 (N_7194,N_7062,N_7031);
nor U7195 (N_7195,N_7038,N_7089);
or U7196 (N_7196,N_7025,N_7023);
nor U7197 (N_7197,N_7065,N_7037);
nor U7198 (N_7198,N_7079,N_7050);
xnor U7199 (N_7199,N_7044,N_7051);
or U7200 (N_7200,N_7016,N_7070);
and U7201 (N_7201,N_7046,N_7030);
and U7202 (N_7202,N_7036,N_7075);
xnor U7203 (N_7203,N_7047,N_7048);
xor U7204 (N_7204,N_7092,N_7107);
nor U7205 (N_7205,N_7100,N_7095);
or U7206 (N_7206,N_7101,N_7118);
nor U7207 (N_7207,N_7115,N_7022);
nand U7208 (N_7208,N_7083,N_7038);
and U7209 (N_7209,N_7090,N_7092);
and U7210 (N_7210,N_7018,N_7012);
or U7211 (N_7211,N_7005,N_7122);
or U7212 (N_7212,N_7021,N_7082);
and U7213 (N_7213,N_7055,N_7105);
nand U7214 (N_7214,N_7094,N_7039);
nand U7215 (N_7215,N_7109,N_7037);
and U7216 (N_7216,N_7117,N_7011);
xnor U7217 (N_7217,N_7103,N_7089);
nor U7218 (N_7218,N_7102,N_7113);
and U7219 (N_7219,N_7101,N_7057);
nand U7220 (N_7220,N_7060,N_7016);
nand U7221 (N_7221,N_7070,N_7017);
and U7222 (N_7222,N_7048,N_7058);
xnor U7223 (N_7223,N_7029,N_7080);
nand U7224 (N_7224,N_7055,N_7023);
nor U7225 (N_7225,N_7052,N_7007);
and U7226 (N_7226,N_7111,N_7078);
and U7227 (N_7227,N_7008,N_7020);
nor U7228 (N_7228,N_7096,N_7030);
or U7229 (N_7229,N_7021,N_7049);
nand U7230 (N_7230,N_7005,N_7027);
or U7231 (N_7231,N_7105,N_7046);
and U7232 (N_7232,N_7101,N_7102);
nand U7233 (N_7233,N_7050,N_7071);
nor U7234 (N_7234,N_7004,N_7069);
or U7235 (N_7235,N_7040,N_7001);
and U7236 (N_7236,N_7034,N_7096);
or U7237 (N_7237,N_7090,N_7046);
nor U7238 (N_7238,N_7080,N_7085);
nand U7239 (N_7239,N_7061,N_7007);
or U7240 (N_7240,N_7074,N_7114);
xor U7241 (N_7241,N_7109,N_7020);
nor U7242 (N_7242,N_7011,N_7111);
and U7243 (N_7243,N_7006,N_7025);
and U7244 (N_7244,N_7028,N_7085);
nand U7245 (N_7245,N_7069,N_7092);
xor U7246 (N_7246,N_7092,N_7101);
and U7247 (N_7247,N_7099,N_7059);
and U7248 (N_7248,N_7005,N_7121);
nor U7249 (N_7249,N_7008,N_7044);
and U7250 (N_7250,N_7239,N_7131);
or U7251 (N_7251,N_7225,N_7151);
nor U7252 (N_7252,N_7169,N_7193);
nor U7253 (N_7253,N_7187,N_7185);
or U7254 (N_7254,N_7170,N_7231);
and U7255 (N_7255,N_7223,N_7183);
nand U7256 (N_7256,N_7242,N_7135);
nor U7257 (N_7257,N_7129,N_7149);
xnor U7258 (N_7258,N_7217,N_7140);
and U7259 (N_7259,N_7199,N_7156);
nand U7260 (N_7260,N_7216,N_7164);
nor U7261 (N_7261,N_7235,N_7142);
nand U7262 (N_7262,N_7228,N_7227);
or U7263 (N_7263,N_7158,N_7200);
nor U7264 (N_7264,N_7148,N_7136);
or U7265 (N_7265,N_7236,N_7172);
and U7266 (N_7266,N_7245,N_7237);
and U7267 (N_7267,N_7204,N_7160);
nand U7268 (N_7268,N_7224,N_7229);
nor U7269 (N_7269,N_7146,N_7232);
nor U7270 (N_7270,N_7188,N_7210);
nand U7271 (N_7271,N_7144,N_7145);
nor U7272 (N_7272,N_7153,N_7189);
and U7273 (N_7273,N_7206,N_7141);
and U7274 (N_7274,N_7125,N_7152);
nand U7275 (N_7275,N_7196,N_7176);
nor U7276 (N_7276,N_7207,N_7127);
nand U7277 (N_7277,N_7157,N_7133);
nor U7278 (N_7278,N_7240,N_7226);
and U7279 (N_7279,N_7186,N_7179);
nor U7280 (N_7280,N_7191,N_7178);
nand U7281 (N_7281,N_7238,N_7246);
or U7282 (N_7282,N_7241,N_7173);
or U7283 (N_7283,N_7161,N_7213);
nor U7284 (N_7284,N_7150,N_7209);
or U7285 (N_7285,N_7132,N_7155);
xnor U7286 (N_7286,N_7190,N_7247);
xnor U7287 (N_7287,N_7138,N_7230);
xor U7288 (N_7288,N_7244,N_7215);
xnor U7289 (N_7289,N_7180,N_7197);
nand U7290 (N_7290,N_7182,N_7162);
xnor U7291 (N_7291,N_7208,N_7221);
nand U7292 (N_7292,N_7203,N_7184);
and U7293 (N_7293,N_7175,N_7181);
and U7294 (N_7294,N_7159,N_7166);
nor U7295 (N_7295,N_7205,N_7134);
and U7296 (N_7296,N_7165,N_7147);
nor U7297 (N_7297,N_7202,N_7163);
and U7298 (N_7298,N_7139,N_7154);
xnor U7299 (N_7299,N_7218,N_7192);
or U7300 (N_7300,N_7130,N_7222);
xor U7301 (N_7301,N_7234,N_7219);
xor U7302 (N_7302,N_7211,N_7171);
xnor U7303 (N_7303,N_7168,N_7220);
or U7304 (N_7304,N_7137,N_7201);
nand U7305 (N_7305,N_7174,N_7248);
or U7306 (N_7306,N_7249,N_7233);
or U7307 (N_7307,N_7212,N_7195);
nand U7308 (N_7308,N_7128,N_7198);
or U7309 (N_7309,N_7167,N_7177);
nand U7310 (N_7310,N_7194,N_7214);
and U7311 (N_7311,N_7143,N_7243);
or U7312 (N_7312,N_7126,N_7187);
nand U7313 (N_7313,N_7212,N_7204);
nor U7314 (N_7314,N_7188,N_7198);
nor U7315 (N_7315,N_7221,N_7128);
nor U7316 (N_7316,N_7137,N_7172);
and U7317 (N_7317,N_7242,N_7185);
or U7318 (N_7318,N_7244,N_7223);
or U7319 (N_7319,N_7137,N_7230);
xnor U7320 (N_7320,N_7231,N_7180);
and U7321 (N_7321,N_7156,N_7125);
or U7322 (N_7322,N_7191,N_7181);
and U7323 (N_7323,N_7175,N_7210);
nand U7324 (N_7324,N_7241,N_7188);
nand U7325 (N_7325,N_7231,N_7201);
and U7326 (N_7326,N_7180,N_7146);
and U7327 (N_7327,N_7211,N_7196);
and U7328 (N_7328,N_7201,N_7181);
nand U7329 (N_7329,N_7163,N_7140);
and U7330 (N_7330,N_7245,N_7182);
or U7331 (N_7331,N_7180,N_7176);
nor U7332 (N_7332,N_7198,N_7149);
xor U7333 (N_7333,N_7162,N_7185);
xor U7334 (N_7334,N_7135,N_7147);
and U7335 (N_7335,N_7213,N_7211);
and U7336 (N_7336,N_7143,N_7209);
and U7337 (N_7337,N_7160,N_7176);
nand U7338 (N_7338,N_7156,N_7173);
nand U7339 (N_7339,N_7138,N_7224);
nand U7340 (N_7340,N_7132,N_7140);
nand U7341 (N_7341,N_7180,N_7153);
nand U7342 (N_7342,N_7230,N_7240);
and U7343 (N_7343,N_7191,N_7225);
or U7344 (N_7344,N_7125,N_7207);
or U7345 (N_7345,N_7213,N_7183);
nor U7346 (N_7346,N_7192,N_7215);
nand U7347 (N_7347,N_7156,N_7179);
or U7348 (N_7348,N_7244,N_7159);
and U7349 (N_7349,N_7160,N_7227);
or U7350 (N_7350,N_7189,N_7172);
nor U7351 (N_7351,N_7204,N_7229);
nand U7352 (N_7352,N_7148,N_7229);
and U7353 (N_7353,N_7200,N_7146);
or U7354 (N_7354,N_7199,N_7160);
nand U7355 (N_7355,N_7232,N_7143);
nand U7356 (N_7356,N_7152,N_7222);
xnor U7357 (N_7357,N_7210,N_7228);
nor U7358 (N_7358,N_7164,N_7196);
and U7359 (N_7359,N_7156,N_7187);
nand U7360 (N_7360,N_7191,N_7188);
xnor U7361 (N_7361,N_7222,N_7214);
and U7362 (N_7362,N_7142,N_7162);
and U7363 (N_7363,N_7244,N_7209);
or U7364 (N_7364,N_7154,N_7216);
xor U7365 (N_7365,N_7215,N_7125);
or U7366 (N_7366,N_7134,N_7238);
nand U7367 (N_7367,N_7170,N_7241);
xnor U7368 (N_7368,N_7166,N_7147);
nor U7369 (N_7369,N_7232,N_7176);
and U7370 (N_7370,N_7162,N_7204);
and U7371 (N_7371,N_7194,N_7183);
xnor U7372 (N_7372,N_7211,N_7144);
and U7373 (N_7373,N_7157,N_7183);
xnor U7374 (N_7374,N_7173,N_7186);
nor U7375 (N_7375,N_7312,N_7355);
xnor U7376 (N_7376,N_7311,N_7303);
or U7377 (N_7377,N_7320,N_7300);
and U7378 (N_7378,N_7255,N_7275);
xnor U7379 (N_7379,N_7287,N_7285);
nand U7380 (N_7380,N_7309,N_7356);
nor U7381 (N_7381,N_7254,N_7273);
and U7382 (N_7382,N_7256,N_7374);
and U7383 (N_7383,N_7298,N_7340);
nand U7384 (N_7384,N_7253,N_7292);
and U7385 (N_7385,N_7357,N_7364);
nor U7386 (N_7386,N_7282,N_7269);
or U7387 (N_7387,N_7263,N_7302);
xor U7388 (N_7388,N_7349,N_7353);
nor U7389 (N_7389,N_7294,N_7286);
or U7390 (N_7390,N_7280,N_7332);
nor U7391 (N_7391,N_7278,N_7373);
nand U7392 (N_7392,N_7348,N_7328);
xor U7393 (N_7393,N_7371,N_7334);
nand U7394 (N_7394,N_7276,N_7317);
xor U7395 (N_7395,N_7274,N_7264);
or U7396 (N_7396,N_7283,N_7369);
nor U7397 (N_7397,N_7299,N_7365);
xor U7398 (N_7398,N_7338,N_7344);
nor U7399 (N_7399,N_7259,N_7277);
xnor U7400 (N_7400,N_7306,N_7296);
xor U7401 (N_7401,N_7367,N_7352);
nor U7402 (N_7402,N_7325,N_7323);
and U7403 (N_7403,N_7362,N_7262);
nor U7404 (N_7404,N_7326,N_7363);
nand U7405 (N_7405,N_7295,N_7370);
or U7406 (N_7406,N_7307,N_7272);
xor U7407 (N_7407,N_7347,N_7301);
xor U7408 (N_7408,N_7324,N_7341);
or U7409 (N_7409,N_7258,N_7316);
nor U7410 (N_7410,N_7315,N_7372);
nor U7411 (N_7411,N_7354,N_7322);
and U7412 (N_7412,N_7345,N_7358);
nor U7413 (N_7413,N_7251,N_7257);
and U7414 (N_7414,N_7271,N_7293);
nand U7415 (N_7415,N_7281,N_7368);
or U7416 (N_7416,N_7267,N_7318);
or U7417 (N_7417,N_7321,N_7360);
nand U7418 (N_7418,N_7310,N_7279);
or U7419 (N_7419,N_7337,N_7291);
or U7420 (N_7420,N_7304,N_7261);
or U7421 (N_7421,N_7314,N_7268);
nand U7422 (N_7422,N_7260,N_7361);
or U7423 (N_7423,N_7313,N_7342);
xor U7424 (N_7424,N_7319,N_7308);
nor U7425 (N_7425,N_7350,N_7366);
and U7426 (N_7426,N_7265,N_7329);
and U7427 (N_7427,N_7284,N_7333);
nand U7428 (N_7428,N_7331,N_7290);
or U7429 (N_7429,N_7359,N_7335);
nor U7430 (N_7430,N_7288,N_7250);
and U7431 (N_7431,N_7346,N_7266);
and U7432 (N_7432,N_7327,N_7351);
nand U7433 (N_7433,N_7289,N_7330);
nand U7434 (N_7434,N_7297,N_7343);
nor U7435 (N_7435,N_7305,N_7339);
nor U7436 (N_7436,N_7252,N_7270);
xnor U7437 (N_7437,N_7336,N_7300);
nor U7438 (N_7438,N_7370,N_7262);
and U7439 (N_7439,N_7358,N_7285);
xnor U7440 (N_7440,N_7284,N_7265);
or U7441 (N_7441,N_7295,N_7307);
and U7442 (N_7442,N_7353,N_7283);
or U7443 (N_7443,N_7365,N_7352);
or U7444 (N_7444,N_7286,N_7319);
nor U7445 (N_7445,N_7350,N_7250);
nand U7446 (N_7446,N_7326,N_7301);
or U7447 (N_7447,N_7309,N_7284);
nor U7448 (N_7448,N_7349,N_7373);
and U7449 (N_7449,N_7349,N_7277);
nand U7450 (N_7450,N_7301,N_7266);
nand U7451 (N_7451,N_7258,N_7335);
nor U7452 (N_7452,N_7360,N_7310);
nand U7453 (N_7453,N_7311,N_7349);
nor U7454 (N_7454,N_7309,N_7262);
and U7455 (N_7455,N_7370,N_7303);
and U7456 (N_7456,N_7252,N_7306);
nor U7457 (N_7457,N_7306,N_7360);
nor U7458 (N_7458,N_7329,N_7270);
and U7459 (N_7459,N_7325,N_7368);
nor U7460 (N_7460,N_7363,N_7332);
nor U7461 (N_7461,N_7251,N_7297);
nand U7462 (N_7462,N_7347,N_7320);
xor U7463 (N_7463,N_7267,N_7322);
or U7464 (N_7464,N_7351,N_7353);
and U7465 (N_7465,N_7372,N_7359);
nor U7466 (N_7466,N_7265,N_7318);
or U7467 (N_7467,N_7365,N_7265);
or U7468 (N_7468,N_7374,N_7313);
xnor U7469 (N_7469,N_7361,N_7261);
or U7470 (N_7470,N_7268,N_7373);
xor U7471 (N_7471,N_7359,N_7303);
and U7472 (N_7472,N_7306,N_7288);
nor U7473 (N_7473,N_7362,N_7280);
nand U7474 (N_7474,N_7371,N_7294);
or U7475 (N_7475,N_7352,N_7363);
and U7476 (N_7476,N_7263,N_7311);
nand U7477 (N_7477,N_7291,N_7345);
xnor U7478 (N_7478,N_7258,N_7322);
nor U7479 (N_7479,N_7374,N_7368);
xor U7480 (N_7480,N_7284,N_7370);
or U7481 (N_7481,N_7357,N_7371);
nand U7482 (N_7482,N_7352,N_7347);
or U7483 (N_7483,N_7281,N_7335);
and U7484 (N_7484,N_7355,N_7269);
nor U7485 (N_7485,N_7256,N_7343);
nand U7486 (N_7486,N_7333,N_7290);
and U7487 (N_7487,N_7326,N_7371);
nor U7488 (N_7488,N_7268,N_7324);
and U7489 (N_7489,N_7254,N_7343);
nand U7490 (N_7490,N_7257,N_7344);
or U7491 (N_7491,N_7329,N_7331);
nand U7492 (N_7492,N_7365,N_7362);
and U7493 (N_7493,N_7372,N_7329);
or U7494 (N_7494,N_7314,N_7252);
nor U7495 (N_7495,N_7369,N_7334);
or U7496 (N_7496,N_7266,N_7308);
and U7497 (N_7497,N_7267,N_7299);
nand U7498 (N_7498,N_7342,N_7345);
nor U7499 (N_7499,N_7270,N_7308);
nand U7500 (N_7500,N_7498,N_7464);
nor U7501 (N_7501,N_7421,N_7387);
nor U7502 (N_7502,N_7440,N_7423);
and U7503 (N_7503,N_7419,N_7436);
or U7504 (N_7504,N_7385,N_7470);
xor U7505 (N_7505,N_7394,N_7453);
nor U7506 (N_7506,N_7494,N_7396);
or U7507 (N_7507,N_7458,N_7401);
xor U7508 (N_7508,N_7376,N_7476);
nor U7509 (N_7509,N_7420,N_7456);
nand U7510 (N_7510,N_7441,N_7481);
xnor U7511 (N_7511,N_7479,N_7381);
nor U7512 (N_7512,N_7386,N_7474);
nand U7513 (N_7513,N_7461,N_7379);
xnor U7514 (N_7514,N_7391,N_7442);
nor U7515 (N_7515,N_7404,N_7432);
xnor U7516 (N_7516,N_7377,N_7499);
nand U7517 (N_7517,N_7465,N_7468);
or U7518 (N_7518,N_7443,N_7444);
nor U7519 (N_7519,N_7418,N_7478);
and U7520 (N_7520,N_7462,N_7435);
nand U7521 (N_7521,N_7490,N_7434);
xnor U7522 (N_7522,N_7407,N_7491);
or U7523 (N_7523,N_7492,N_7405);
xor U7524 (N_7524,N_7398,N_7378);
nand U7525 (N_7525,N_7452,N_7477);
or U7526 (N_7526,N_7451,N_7428);
xnor U7527 (N_7527,N_7411,N_7414);
nand U7528 (N_7528,N_7431,N_7466);
and U7529 (N_7529,N_7412,N_7493);
nand U7530 (N_7530,N_7449,N_7450);
nand U7531 (N_7531,N_7393,N_7399);
and U7532 (N_7532,N_7467,N_7427);
and U7533 (N_7533,N_7382,N_7406);
nor U7534 (N_7534,N_7390,N_7429);
nand U7535 (N_7535,N_7483,N_7383);
xnor U7536 (N_7536,N_7433,N_7489);
xor U7537 (N_7537,N_7475,N_7417);
or U7538 (N_7538,N_7375,N_7496);
or U7539 (N_7539,N_7430,N_7455);
and U7540 (N_7540,N_7488,N_7425);
and U7541 (N_7541,N_7472,N_7438);
or U7542 (N_7542,N_7392,N_7473);
xnor U7543 (N_7543,N_7437,N_7416);
nor U7544 (N_7544,N_7484,N_7426);
or U7545 (N_7545,N_7408,N_7469);
and U7546 (N_7546,N_7487,N_7454);
nand U7547 (N_7547,N_7497,N_7495);
nand U7548 (N_7548,N_7415,N_7413);
nor U7549 (N_7549,N_7388,N_7409);
or U7550 (N_7550,N_7400,N_7446);
or U7551 (N_7551,N_7389,N_7448);
or U7552 (N_7552,N_7485,N_7384);
nand U7553 (N_7553,N_7403,N_7457);
nand U7554 (N_7554,N_7482,N_7447);
nand U7555 (N_7555,N_7402,N_7395);
and U7556 (N_7556,N_7486,N_7397);
and U7557 (N_7557,N_7424,N_7460);
or U7558 (N_7558,N_7463,N_7480);
nor U7559 (N_7559,N_7471,N_7410);
and U7560 (N_7560,N_7422,N_7445);
nor U7561 (N_7561,N_7459,N_7380);
nand U7562 (N_7562,N_7439,N_7471);
xnor U7563 (N_7563,N_7447,N_7461);
nand U7564 (N_7564,N_7449,N_7379);
xor U7565 (N_7565,N_7428,N_7455);
nor U7566 (N_7566,N_7416,N_7497);
nand U7567 (N_7567,N_7452,N_7441);
nand U7568 (N_7568,N_7472,N_7424);
and U7569 (N_7569,N_7472,N_7464);
nand U7570 (N_7570,N_7414,N_7387);
or U7571 (N_7571,N_7388,N_7497);
and U7572 (N_7572,N_7469,N_7481);
nor U7573 (N_7573,N_7437,N_7390);
and U7574 (N_7574,N_7497,N_7375);
and U7575 (N_7575,N_7408,N_7467);
or U7576 (N_7576,N_7487,N_7394);
or U7577 (N_7577,N_7479,N_7387);
nand U7578 (N_7578,N_7420,N_7449);
and U7579 (N_7579,N_7435,N_7490);
nor U7580 (N_7580,N_7429,N_7420);
nor U7581 (N_7581,N_7437,N_7470);
nand U7582 (N_7582,N_7427,N_7482);
xnor U7583 (N_7583,N_7475,N_7493);
nor U7584 (N_7584,N_7416,N_7435);
or U7585 (N_7585,N_7451,N_7377);
nor U7586 (N_7586,N_7424,N_7454);
and U7587 (N_7587,N_7401,N_7378);
or U7588 (N_7588,N_7392,N_7444);
nor U7589 (N_7589,N_7484,N_7387);
and U7590 (N_7590,N_7442,N_7448);
nor U7591 (N_7591,N_7448,N_7429);
or U7592 (N_7592,N_7415,N_7385);
and U7593 (N_7593,N_7385,N_7399);
and U7594 (N_7594,N_7482,N_7466);
xor U7595 (N_7595,N_7456,N_7401);
and U7596 (N_7596,N_7412,N_7433);
nand U7597 (N_7597,N_7381,N_7481);
nor U7598 (N_7598,N_7432,N_7407);
and U7599 (N_7599,N_7382,N_7395);
and U7600 (N_7600,N_7439,N_7476);
and U7601 (N_7601,N_7465,N_7391);
nand U7602 (N_7602,N_7428,N_7376);
and U7603 (N_7603,N_7494,N_7406);
nand U7604 (N_7604,N_7433,N_7479);
nor U7605 (N_7605,N_7387,N_7437);
and U7606 (N_7606,N_7488,N_7445);
nor U7607 (N_7607,N_7445,N_7399);
nand U7608 (N_7608,N_7379,N_7382);
xnor U7609 (N_7609,N_7376,N_7496);
xnor U7610 (N_7610,N_7466,N_7375);
nor U7611 (N_7611,N_7471,N_7476);
nand U7612 (N_7612,N_7469,N_7447);
xnor U7613 (N_7613,N_7473,N_7486);
nand U7614 (N_7614,N_7414,N_7392);
or U7615 (N_7615,N_7428,N_7390);
nand U7616 (N_7616,N_7411,N_7452);
or U7617 (N_7617,N_7482,N_7393);
nor U7618 (N_7618,N_7493,N_7405);
nand U7619 (N_7619,N_7402,N_7401);
or U7620 (N_7620,N_7398,N_7428);
nor U7621 (N_7621,N_7400,N_7437);
xnor U7622 (N_7622,N_7390,N_7398);
nand U7623 (N_7623,N_7415,N_7477);
nand U7624 (N_7624,N_7448,N_7454);
or U7625 (N_7625,N_7509,N_7508);
xor U7626 (N_7626,N_7613,N_7528);
nor U7627 (N_7627,N_7507,N_7563);
xor U7628 (N_7628,N_7514,N_7558);
xor U7629 (N_7629,N_7607,N_7535);
nor U7630 (N_7630,N_7553,N_7540);
nand U7631 (N_7631,N_7516,N_7561);
nand U7632 (N_7632,N_7579,N_7590);
xnor U7633 (N_7633,N_7564,N_7538);
or U7634 (N_7634,N_7500,N_7578);
or U7635 (N_7635,N_7623,N_7622);
nand U7636 (N_7636,N_7596,N_7593);
xor U7637 (N_7637,N_7548,N_7527);
or U7638 (N_7638,N_7595,N_7525);
and U7639 (N_7639,N_7615,N_7611);
nand U7640 (N_7640,N_7599,N_7582);
nor U7641 (N_7641,N_7522,N_7619);
nand U7642 (N_7642,N_7505,N_7586);
and U7643 (N_7643,N_7600,N_7559);
nand U7644 (N_7644,N_7608,N_7542);
xnor U7645 (N_7645,N_7589,N_7618);
and U7646 (N_7646,N_7552,N_7620);
and U7647 (N_7647,N_7547,N_7512);
nand U7648 (N_7648,N_7501,N_7557);
and U7649 (N_7649,N_7592,N_7555);
xnor U7650 (N_7650,N_7565,N_7544);
nand U7651 (N_7651,N_7511,N_7549);
or U7652 (N_7652,N_7605,N_7574);
nand U7653 (N_7653,N_7606,N_7588);
nor U7654 (N_7654,N_7531,N_7576);
or U7655 (N_7655,N_7520,N_7510);
nor U7656 (N_7656,N_7621,N_7529);
xor U7657 (N_7657,N_7617,N_7585);
nor U7658 (N_7658,N_7541,N_7581);
nand U7659 (N_7659,N_7594,N_7568);
xor U7660 (N_7660,N_7572,N_7543);
and U7661 (N_7661,N_7598,N_7554);
or U7662 (N_7662,N_7515,N_7551);
or U7663 (N_7663,N_7519,N_7521);
nor U7664 (N_7664,N_7534,N_7597);
or U7665 (N_7665,N_7545,N_7567);
and U7666 (N_7666,N_7539,N_7612);
nand U7667 (N_7667,N_7506,N_7533);
nand U7668 (N_7668,N_7523,N_7569);
xnor U7669 (N_7669,N_7609,N_7546);
nand U7670 (N_7670,N_7614,N_7503);
or U7671 (N_7671,N_7616,N_7570);
and U7672 (N_7672,N_7560,N_7504);
or U7673 (N_7673,N_7537,N_7513);
xnor U7674 (N_7674,N_7573,N_7584);
xnor U7675 (N_7675,N_7610,N_7604);
nor U7676 (N_7676,N_7562,N_7526);
nor U7677 (N_7677,N_7575,N_7502);
xnor U7678 (N_7678,N_7580,N_7524);
nand U7679 (N_7679,N_7536,N_7591);
xor U7680 (N_7680,N_7603,N_7583);
nor U7681 (N_7681,N_7577,N_7601);
nand U7682 (N_7682,N_7602,N_7556);
and U7683 (N_7683,N_7566,N_7587);
nor U7684 (N_7684,N_7532,N_7530);
and U7685 (N_7685,N_7571,N_7518);
nor U7686 (N_7686,N_7517,N_7550);
nand U7687 (N_7687,N_7624,N_7534);
or U7688 (N_7688,N_7517,N_7569);
and U7689 (N_7689,N_7592,N_7558);
xor U7690 (N_7690,N_7515,N_7550);
xnor U7691 (N_7691,N_7621,N_7505);
xor U7692 (N_7692,N_7608,N_7519);
nor U7693 (N_7693,N_7579,N_7603);
and U7694 (N_7694,N_7518,N_7584);
nor U7695 (N_7695,N_7542,N_7541);
or U7696 (N_7696,N_7609,N_7575);
xnor U7697 (N_7697,N_7573,N_7559);
or U7698 (N_7698,N_7579,N_7567);
and U7699 (N_7699,N_7536,N_7568);
and U7700 (N_7700,N_7614,N_7608);
xor U7701 (N_7701,N_7520,N_7512);
nor U7702 (N_7702,N_7569,N_7586);
or U7703 (N_7703,N_7519,N_7574);
nand U7704 (N_7704,N_7607,N_7614);
and U7705 (N_7705,N_7610,N_7507);
and U7706 (N_7706,N_7624,N_7616);
and U7707 (N_7707,N_7552,N_7610);
xnor U7708 (N_7708,N_7571,N_7581);
or U7709 (N_7709,N_7522,N_7529);
nor U7710 (N_7710,N_7554,N_7596);
xnor U7711 (N_7711,N_7592,N_7501);
and U7712 (N_7712,N_7500,N_7551);
nand U7713 (N_7713,N_7606,N_7539);
nor U7714 (N_7714,N_7587,N_7597);
xnor U7715 (N_7715,N_7520,N_7529);
or U7716 (N_7716,N_7581,N_7618);
nand U7717 (N_7717,N_7519,N_7580);
xor U7718 (N_7718,N_7582,N_7539);
or U7719 (N_7719,N_7564,N_7622);
nor U7720 (N_7720,N_7581,N_7534);
nand U7721 (N_7721,N_7500,N_7537);
xor U7722 (N_7722,N_7560,N_7544);
nor U7723 (N_7723,N_7548,N_7589);
nor U7724 (N_7724,N_7553,N_7536);
xor U7725 (N_7725,N_7604,N_7611);
and U7726 (N_7726,N_7511,N_7608);
and U7727 (N_7727,N_7536,N_7619);
nand U7728 (N_7728,N_7547,N_7500);
and U7729 (N_7729,N_7561,N_7585);
and U7730 (N_7730,N_7614,N_7546);
xor U7731 (N_7731,N_7521,N_7623);
nor U7732 (N_7732,N_7566,N_7513);
xnor U7733 (N_7733,N_7549,N_7505);
or U7734 (N_7734,N_7514,N_7586);
nand U7735 (N_7735,N_7544,N_7502);
xnor U7736 (N_7736,N_7543,N_7545);
nand U7737 (N_7737,N_7546,N_7568);
nor U7738 (N_7738,N_7524,N_7601);
or U7739 (N_7739,N_7611,N_7574);
nand U7740 (N_7740,N_7593,N_7570);
xor U7741 (N_7741,N_7595,N_7593);
and U7742 (N_7742,N_7549,N_7542);
nor U7743 (N_7743,N_7508,N_7601);
and U7744 (N_7744,N_7596,N_7597);
nor U7745 (N_7745,N_7571,N_7569);
and U7746 (N_7746,N_7559,N_7533);
and U7747 (N_7747,N_7578,N_7591);
and U7748 (N_7748,N_7551,N_7581);
xnor U7749 (N_7749,N_7582,N_7579);
and U7750 (N_7750,N_7655,N_7678);
xor U7751 (N_7751,N_7746,N_7713);
or U7752 (N_7752,N_7705,N_7660);
nor U7753 (N_7753,N_7708,N_7654);
nand U7754 (N_7754,N_7729,N_7670);
and U7755 (N_7755,N_7679,N_7635);
xnor U7756 (N_7756,N_7683,N_7665);
nor U7757 (N_7757,N_7685,N_7711);
or U7758 (N_7758,N_7715,N_7658);
xor U7759 (N_7759,N_7677,N_7659);
or U7760 (N_7760,N_7687,N_7733);
nand U7761 (N_7761,N_7739,N_7731);
nand U7762 (N_7762,N_7641,N_7747);
and U7763 (N_7763,N_7627,N_7673);
xor U7764 (N_7764,N_7637,N_7682);
and U7765 (N_7765,N_7640,N_7642);
and U7766 (N_7766,N_7730,N_7676);
or U7767 (N_7767,N_7644,N_7662);
nor U7768 (N_7768,N_7681,N_7709);
or U7769 (N_7769,N_7671,N_7645);
and U7770 (N_7770,N_7699,N_7649);
nor U7771 (N_7771,N_7639,N_7720);
nor U7772 (N_7772,N_7738,N_7694);
xor U7773 (N_7773,N_7727,N_7634);
nand U7774 (N_7774,N_7629,N_7704);
xnor U7775 (N_7775,N_7668,N_7669);
xor U7776 (N_7776,N_7737,N_7672);
and U7777 (N_7777,N_7723,N_7698);
and U7778 (N_7778,N_7745,N_7651);
and U7779 (N_7779,N_7631,N_7716);
or U7780 (N_7780,N_7686,N_7736);
or U7781 (N_7781,N_7721,N_7718);
nor U7782 (N_7782,N_7706,N_7735);
xnor U7783 (N_7783,N_7633,N_7726);
or U7784 (N_7784,N_7701,N_7700);
nor U7785 (N_7785,N_7666,N_7722);
or U7786 (N_7786,N_7657,N_7697);
nor U7787 (N_7787,N_7710,N_7628);
nand U7788 (N_7788,N_7661,N_7734);
nand U7789 (N_7789,N_7725,N_7696);
and U7790 (N_7790,N_7732,N_7688);
and U7791 (N_7791,N_7689,N_7692);
and U7792 (N_7792,N_7653,N_7663);
nor U7793 (N_7793,N_7636,N_7744);
or U7794 (N_7794,N_7724,N_7648);
and U7795 (N_7795,N_7656,N_7728);
nor U7796 (N_7796,N_7695,N_7630);
and U7797 (N_7797,N_7664,N_7647);
nand U7798 (N_7798,N_7632,N_7652);
and U7799 (N_7799,N_7693,N_7625);
nand U7800 (N_7800,N_7749,N_7638);
or U7801 (N_7801,N_7684,N_7748);
nor U7802 (N_7802,N_7719,N_7626);
nor U7803 (N_7803,N_7702,N_7741);
or U7804 (N_7804,N_7740,N_7691);
xor U7805 (N_7805,N_7646,N_7707);
nand U7806 (N_7806,N_7643,N_7717);
nand U7807 (N_7807,N_7680,N_7650);
xnor U7808 (N_7808,N_7742,N_7667);
nand U7809 (N_7809,N_7703,N_7674);
xnor U7810 (N_7810,N_7714,N_7675);
nor U7811 (N_7811,N_7690,N_7712);
xor U7812 (N_7812,N_7743,N_7717);
and U7813 (N_7813,N_7689,N_7746);
and U7814 (N_7814,N_7631,N_7734);
nand U7815 (N_7815,N_7671,N_7664);
nand U7816 (N_7816,N_7654,N_7687);
nor U7817 (N_7817,N_7668,N_7700);
or U7818 (N_7818,N_7673,N_7695);
or U7819 (N_7819,N_7702,N_7665);
or U7820 (N_7820,N_7675,N_7722);
nand U7821 (N_7821,N_7628,N_7698);
nand U7822 (N_7822,N_7663,N_7709);
and U7823 (N_7823,N_7704,N_7627);
and U7824 (N_7824,N_7625,N_7679);
nor U7825 (N_7825,N_7663,N_7689);
nor U7826 (N_7826,N_7747,N_7632);
xnor U7827 (N_7827,N_7663,N_7725);
or U7828 (N_7828,N_7676,N_7719);
and U7829 (N_7829,N_7730,N_7655);
xor U7830 (N_7830,N_7671,N_7702);
nand U7831 (N_7831,N_7675,N_7662);
or U7832 (N_7832,N_7682,N_7722);
nor U7833 (N_7833,N_7732,N_7705);
nand U7834 (N_7834,N_7733,N_7714);
nand U7835 (N_7835,N_7674,N_7744);
and U7836 (N_7836,N_7741,N_7738);
nor U7837 (N_7837,N_7665,N_7629);
nand U7838 (N_7838,N_7656,N_7694);
and U7839 (N_7839,N_7725,N_7736);
xor U7840 (N_7840,N_7720,N_7644);
nand U7841 (N_7841,N_7632,N_7683);
nand U7842 (N_7842,N_7643,N_7662);
or U7843 (N_7843,N_7648,N_7706);
nand U7844 (N_7844,N_7672,N_7707);
and U7845 (N_7845,N_7734,N_7737);
nand U7846 (N_7846,N_7631,N_7681);
xor U7847 (N_7847,N_7678,N_7694);
nand U7848 (N_7848,N_7731,N_7728);
or U7849 (N_7849,N_7658,N_7632);
xnor U7850 (N_7850,N_7684,N_7672);
or U7851 (N_7851,N_7680,N_7664);
or U7852 (N_7852,N_7739,N_7633);
nor U7853 (N_7853,N_7679,N_7715);
and U7854 (N_7854,N_7637,N_7680);
and U7855 (N_7855,N_7742,N_7702);
nand U7856 (N_7856,N_7673,N_7736);
nor U7857 (N_7857,N_7708,N_7687);
and U7858 (N_7858,N_7723,N_7657);
xnor U7859 (N_7859,N_7730,N_7627);
xor U7860 (N_7860,N_7690,N_7668);
xnor U7861 (N_7861,N_7693,N_7731);
or U7862 (N_7862,N_7647,N_7680);
nand U7863 (N_7863,N_7640,N_7633);
or U7864 (N_7864,N_7636,N_7679);
and U7865 (N_7865,N_7638,N_7715);
xor U7866 (N_7866,N_7728,N_7736);
and U7867 (N_7867,N_7736,N_7715);
nand U7868 (N_7868,N_7711,N_7692);
nor U7869 (N_7869,N_7635,N_7669);
or U7870 (N_7870,N_7691,N_7742);
and U7871 (N_7871,N_7697,N_7648);
or U7872 (N_7872,N_7687,N_7704);
xnor U7873 (N_7873,N_7628,N_7638);
nand U7874 (N_7874,N_7744,N_7665);
nor U7875 (N_7875,N_7808,N_7849);
nand U7876 (N_7876,N_7858,N_7826);
and U7877 (N_7877,N_7837,N_7864);
nand U7878 (N_7878,N_7801,N_7870);
xor U7879 (N_7879,N_7798,N_7846);
nor U7880 (N_7880,N_7825,N_7852);
nand U7881 (N_7881,N_7788,N_7871);
nor U7882 (N_7882,N_7847,N_7772);
and U7883 (N_7883,N_7761,N_7765);
nand U7884 (N_7884,N_7799,N_7835);
nand U7885 (N_7885,N_7792,N_7797);
xnor U7886 (N_7886,N_7851,N_7755);
xor U7887 (N_7887,N_7818,N_7810);
nand U7888 (N_7888,N_7800,N_7831);
xor U7889 (N_7889,N_7840,N_7812);
xnor U7890 (N_7890,N_7865,N_7853);
or U7891 (N_7891,N_7859,N_7861);
xnor U7892 (N_7892,N_7796,N_7844);
and U7893 (N_7893,N_7839,N_7794);
or U7894 (N_7894,N_7752,N_7770);
or U7895 (N_7895,N_7814,N_7795);
nand U7896 (N_7896,N_7768,N_7819);
nor U7897 (N_7897,N_7764,N_7756);
xor U7898 (N_7898,N_7869,N_7760);
or U7899 (N_7899,N_7763,N_7766);
nand U7900 (N_7900,N_7780,N_7821);
or U7901 (N_7901,N_7813,N_7838);
xor U7902 (N_7902,N_7854,N_7784);
or U7903 (N_7903,N_7787,N_7811);
nor U7904 (N_7904,N_7750,N_7803);
nand U7905 (N_7905,N_7785,N_7751);
nor U7906 (N_7906,N_7805,N_7786);
or U7907 (N_7907,N_7867,N_7874);
nor U7908 (N_7908,N_7827,N_7868);
nor U7909 (N_7909,N_7775,N_7771);
nor U7910 (N_7910,N_7779,N_7832);
xnor U7911 (N_7911,N_7789,N_7767);
nor U7912 (N_7912,N_7866,N_7823);
nor U7913 (N_7913,N_7817,N_7862);
nand U7914 (N_7914,N_7807,N_7753);
xnor U7915 (N_7915,N_7873,N_7822);
xor U7916 (N_7916,N_7806,N_7816);
nor U7917 (N_7917,N_7863,N_7774);
xor U7918 (N_7918,N_7757,N_7843);
nand U7919 (N_7919,N_7769,N_7778);
or U7920 (N_7920,N_7824,N_7855);
or U7921 (N_7921,N_7872,N_7773);
nand U7922 (N_7922,N_7793,N_7828);
xor U7923 (N_7923,N_7783,N_7834);
xor U7924 (N_7924,N_7777,N_7860);
or U7925 (N_7925,N_7841,N_7848);
and U7926 (N_7926,N_7842,N_7836);
xor U7927 (N_7927,N_7758,N_7809);
xor U7928 (N_7928,N_7759,N_7833);
xnor U7929 (N_7929,N_7791,N_7850);
xnor U7930 (N_7930,N_7815,N_7776);
and U7931 (N_7931,N_7782,N_7856);
xor U7932 (N_7932,N_7820,N_7802);
xor U7933 (N_7933,N_7845,N_7754);
or U7934 (N_7934,N_7790,N_7762);
and U7935 (N_7935,N_7857,N_7830);
nand U7936 (N_7936,N_7781,N_7804);
and U7937 (N_7937,N_7829,N_7776);
nor U7938 (N_7938,N_7807,N_7795);
nand U7939 (N_7939,N_7846,N_7866);
nand U7940 (N_7940,N_7831,N_7855);
nor U7941 (N_7941,N_7791,N_7834);
or U7942 (N_7942,N_7788,N_7873);
and U7943 (N_7943,N_7775,N_7863);
nor U7944 (N_7944,N_7846,N_7860);
and U7945 (N_7945,N_7863,N_7773);
or U7946 (N_7946,N_7778,N_7857);
xor U7947 (N_7947,N_7762,N_7865);
xnor U7948 (N_7948,N_7843,N_7788);
or U7949 (N_7949,N_7816,N_7760);
nor U7950 (N_7950,N_7751,N_7831);
nand U7951 (N_7951,N_7808,N_7873);
nor U7952 (N_7952,N_7797,N_7782);
nor U7953 (N_7953,N_7813,N_7772);
or U7954 (N_7954,N_7765,N_7859);
nand U7955 (N_7955,N_7800,N_7763);
xnor U7956 (N_7956,N_7798,N_7801);
nand U7957 (N_7957,N_7800,N_7751);
and U7958 (N_7958,N_7754,N_7764);
nand U7959 (N_7959,N_7794,N_7780);
nand U7960 (N_7960,N_7838,N_7834);
or U7961 (N_7961,N_7820,N_7805);
nand U7962 (N_7962,N_7810,N_7842);
nand U7963 (N_7963,N_7827,N_7780);
xor U7964 (N_7964,N_7862,N_7871);
nand U7965 (N_7965,N_7870,N_7751);
nor U7966 (N_7966,N_7824,N_7866);
and U7967 (N_7967,N_7826,N_7832);
and U7968 (N_7968,N_7751,N_7779);
xnor U7969 (N_7969,N_7818,N_7837);
or U7970 (N_7970,N_7779,N_7814);
xnor U7971 (N_7971,N_7851,N_7761);
nor U7972 (N_7972,N_7871,N_7852);
and U7973 (N_7973,N_7794,N_7820);
or U7974 (N_7974,N_7758,N_7858);
or U7975 (N_7975,N_7768,N_7843);
and U7976 (N_7976,N_7754,N_7822);
nor U7977 (N_7977,N_7813,N_7827);
and U7978 (N_7978,N_7856,N_7750);
or U7979 (N_7979,N_7863,N_7829);
nand U7980 (N_7980,N_7824,N_7864);
and U7981 (N_7981,N_7833,N_7856);
xnor U7982 (N_7982,N_7868,N_7794);
or U7983 (N_7983,N_7766,N_7794);
nor U7984 (N_7984,N_7767,N_7845);
xor U7985 (N_7985,N_7770,N_7832);
nand U7986 (N_7986,N_7773,N_7811);
nor U7987 (N_7987,N_7820,N_7788);
nand U7988 (N_7988,N_7801,N_7750);
and U7989 (N_7989,N_7824,N_7764);
or U7990 (N_7990,N_7831,N_7872);
xor U7991 (N_7991,N_7787,N_7788);
xnor U7992 (N_7992,N_7810,N_7813);
xor U7993 (N_7993,N_7828,N_7865);
nor U7994 (N_7994,N_7801,N_7799);
nor U7995 (N_7995,N_7796,N_7790);
nand U7996 (N_7996,N_7821,N_7756);
xnor U7997 (N_7997,N_7805,N_7768);
xnor U7998 (N_7998,N_7793,N_7754);
nor U7999 (N_7999,N_7826,N_7777);
xnor U8000 (N_8000,N_7970,N_7991);
or U8001 (N_8001,N_7953,N_7976);
nand U8002 (N_8002,N_7906,N_7960);
or U8003 (N_8003,N_7936,N_7903);
nor U8004 (N_8004,N_7973,N_7956);
xnor U8005 (N_8005,N_7918,N_7877);
or U8006 (N_8006,N_7892,N_7886);
and U8007 (N_8007,N_7978,N_7919);
nand U8008 (N_8008,N_7997,N_7943);
nand U8009 (N_8009,N_7962,N_7964);
or U8010 (N_8010,N_7945,N_7900);
nor U8011 (N_8011,N_7916,N_7999);
and U8012 (N_8012,N_7954,N_7887);
or U8013 (N_8013,N_7898,N_7926);
and U8014 (N_8014,N_7947,N_7968);
nor U8015 (N_8015,N_7940,N_7975);
nand U8016 (N_8016,N_7984,N_7941);
nand U8017 (N_8017,N_7895,N_7883);
nand U8018 (N_8018,N_7986,N_7993);
xnor U8019 (N_8019,N_7980,N_7937);
nand U8020 (N_8020,N_7938,N_7929);
nor U8021 (N_8021,N_7952,N_7890);
nand U8022 (N_8022,N_7957,N_7989);
or U8023 (N_8023,N_7917,N_7927);
nand U8024 (N_8024,N_7889,N_7955);
nor U8025 (N_8025,N_7934,N_7963);
or U8026 (N_8026,N_7907,N_7987);
nor U8027 (N_8027,N_7914,N_7961);
and U8028 (N_8028,N_7995,N_7891);
nor U8029 (N_8029,N_7902,N_7884);
nand U8030 (N_8030,N_7879,N_7996);
nand U8031 (N_8031,N_7888,N_7972);
nand U8032 (N_8032,N_7958,N_7920);
or U8033 (N_8033,N_7933,N_7905);
xor U8034 (N_8034,N_7904,N_7913);
nor U8035 (N_8035,N_7959,N_7951);
xnor U8036 (N_8036,N_7910,N_7878);
nor U8037 (N_8037,N_7985,N_7935);
and U8038 (N_8038,N_7915,N_7876);
xnor U8039 (N_8039,N_7944,N_7983);
xor U8040 (N_8040,N_7924,N_7896);
or U8041 (N_8041,N_7946,N_7885);
or U8042 (N_8042,N_7930,N_7965);
nand U8043 (N_8043,N_7971,N_7948);
and U8044 (N_8044,N_7994,N_7909);
and U8045 (N_8045,N_7931,N_7998);
or U8046 (N_8046,N_7928,N_7967);
xnor U8047 (N_8047,N_7939,N_7881);
nand U8048 (N_8048,N_7974,N_7950);
nand U8049 (N_8049,N_7966,N_7880);
nor U8050 (N_8050,N_7875,N_7893);
or U8051 (N_8051,N_7901,N_7949);
xnor U8052 (N_8052,N_7897,N_7911);
xor U8053 (N_8053,N_7912,N_7981);
nor U8054 (N_8054,N_7942,N_7977);
nand U8055 (N_8055,N_7894,N_7882);
nor U8056 (N_8056,N_7979,N_7908);
nand U8057 (N_8057,N_7988,N_7992);
xor U8058 (N_8058,N_7932,N_7925);
or U8059 (N_8059,N_7921,N_7899);
and U8060 (N_8060,N_7922,N_7990);
and U8061 (N_8061,N_7969,N_7982);
xor U8062 (N_8062,N_7923,N_7907);
nand U8063 (N_8063,N_7958,N_7985);
or U8064 (N_8064,N_7926,N_7890);
nor U8065 (N_8065,N_7894,N_7925);
or U8066 (N_8066,N_7910,N_7934);
or U8067 (N_8067,N_7971,N_7970);
nor U8068 (N_8068,N_7985,N_7895);
or U8069 (N_8069,N_7911,N_7875);
or U8070 (N_8070,N_7968,N_7965);
nor U8071 (N_8071,N_7941,N_7959);
xor U8072 (N_8072,N_7952,N_7905);
xor U8073 (N_8073,N_7979,N_7980);
xnor U8074 (N_8074,N_7993,N_7915);
and U8075 (N_8075,N_7951,N_7917);
and U8076 (N_8076,N_7945,N_7926);
xnor U8077 (N_8077,N_7903,N_7998);
and U8078 (N_8078,N_7962,N_7957);
nand U8079 (N_8079,N_7998,N_7893);
nor U8080 (N_8080,N_7925,N_7992);
nand U8081 (N_8081,N_7947,N_7980);
or U8082 (N_8082,N_7945,N_7898);
nand U8083 (N_8083,N_7970,N_7884);
xor U8084 (N_8084,N_7939,N_7889);
nand U8085 (N_8085,N_7999,N_7982);
nor U8086 (N_8086,N_7952,N_7885);
xor U8087 (N_8087,N_7974,N_7886);
nor U8088 (N_8088,N_7922,N_7967);
nor U8089 (N_8089,N_7969,N_7994);
nand U8090 (N_8090,N_7986,N_7937);
and U8091 (N_8091,N_7941,N_7921);
and U8092 (N_8092,N_7996,N_7962);
xor U8093 (N_8093,N_7974,N_7920);
xnor U8094 (N_8094,N_7962,N_7991);
or U8095 (N_8095,N_7879,N_7892);
or U8096 (N_8096,N_7966,N_7958);
nand U8097 (N_8097,N_7963,N_7951);
nand U8098 (N_8098,N_7998,N_7987);
xor U8099 (N_8099,N_7971,N_7974);
or U8100 (N_8100,N_7992,N_7876);
nand U8101 (N_8101,N_7935,N_7952);
or U8102 (N_8102,N_7891,N_7938);
nand U8103 (N_8103,N_7947,N_7924);
nor U8104 (N_8104,N_7892,N_7909);
nor U8105 (N_8105,N_7931,N_7956);
nand U8106 (N_8106,N_7929,N_7957);
and U8107 (N_8107,N_7941,N_7914);
nor U8108 (N_8108,N_7992,N_7916);
nor U8109 (N_8109,N_7997,N_7884);
nand U8110 (N_8110,N_7945,N_7885);
nor U8111 (N_8111,N_7959,N_7990);
and U8112 (N_8112,N_7914,N_7926);
or U8113 (N_8113,N_7878,N_7875);
nand U8114 (N_8114,N_7907,N_7877);
and U8115 (N_8115,N_7888,N_7976);
nand U8116 (N_8116,N_7958,N_7899);
and U8117 (N_8117,N_7909,N_7880);
nand U8118 (N_8118,N_7894,N_7950);
nor U8119 (N_8119,N_7942,N_7983);
xnor U8120 (N_8120,N_7886,N_7920);
nor U8121 (N_8121,N_7991,N_7986);
nor U8122 (N_8122,N_7979,N_7882);
or U8123 (N_8123,N_7888,N_7921);
or U8124 (N_8124,N_7971,N_7985);
and U8125 (N_8125,N_8103,N_8090);
nand U8126 (N_8126,N_8119,N_8102);
xnor U8127 (N_8127,N_8000,N_8007);
or U8128 (N_8128,N_8124,N_8011);
and U8129 (N_8129,N_8113,N_8029);
or U8130 (N_8130,N_8104,N_8001);
xor U8131 (N_8131,N_8086,N_8053);
or U8132 (N_8132,N_8121,N_8031);
or U8133 (N_8133,N_8027,N_8005);
nor U8134 (N_8134,N_8016,N_8046);
or U8135 (N_8135,N_8115,N_8004);
nor U8136 (N_8136,N_8048,N_8019);
nor U8137 (N_8137,N_8110,N_8120);
nand U8138 (N_8138,N_8096,N_8038);
or U8139 (N_8139,N_8056,N_8050);
or U8140 (N_8140,N_8101,N_8018);
nor U8141 (N_8141,N_8085,N_8057);
xnor U8142 (N_8142,N_8002,N_8006);
and U8143 (N_8143,N_8095,N_8108);
and U8144 (N_8144,N_8064,N_8045);
or U8145 (N_8145,N_8030,N_8043);
and U8146 (N_8146,N_8062,N_8052);
and U8147 (N_8147,N_8015,N_8024);
or U8148 (N_8148,N_8073,N_8078);
xnor U8149 (N_8149,N_8058,N_8014);
and U8150 (N_8150,N_8072,N_8118);
nor U8151 (N_8151,N_8059,N_8068);
nor U8152 (N_8152,N_8079,N_8084);
or U8153 (N_8153,N_8063,N_8035);
and U8154 (N_8154,N_8039,N_8080);
nor U8155 (N_8155,N_8123,N_8069);
or U8156 (N_8156,N_8099,N_8100);
xor U8157 (N_8157,N_8026,N_8066);
xnor U8158 (N_8158,N_8122,N_8033);
or U8159 (N_8159,N_8034,N_8098);
or U8160 (N_8160,N_8105,N_8094);
nor U8161 (N_8161,N_8071,N_8044);
and U8162 (N_8162,N_8107,N_8061);
xor U8163 (N_8163,N_8021,N_8049);
xor U8164 (N_8164,N_8092,N_8028);
or U8165 (N_8165,N_8074,N_8093);
or U8166 (N_8166,N_8055,N_8091);
xnor U8167 (N_8167,N_8111,N_8017);
or U8168 (N_8168,N_8008,N_8012);
or U8169 (N_8169,N_8112,N_8054);
nor U8170 (N_8170,N_8060,N_8087);
and U8171 (N_8171,N_8020,N_8082);
xor U8172 (N_8172,N_8036,N_8117);
and U8173 (N_8173,N_8116,N_8106);
xor U8174 (N_8174,N_8047,N_8089);
and U8175 (N_8175,N_8083,N_8022);
or U8176 (N_8176,N_8081,N_8037);
and U8177 (N_8177,N_8076,N_8013);
nand U8178 (N_8178,N_8010,N_8067);
nor U8179 (N_8179,N_8041,N_8051);
and U8180 (N_8180,N_8032,N_8003);
nand U8181 (N_8181,N_8042,N_8088);
nor U8182 (N_8182,N_8114,N_8097);
and U8183 (N_8183,N_8023,N_8025);
and U8184 (N_8184,N_8009,N_8075);
and U8185 (N_8185,N_8077,N_8040);
or U8186 (N_8186,N_8109,N_8065);
or U8187 (N_8187,N_8070,N_8041);
and U8188 (N_8188,N_8101,N_8099);
and U8189 (N_8189,N_8097,N_8003);
or U8190 (N_8190,N_8043,N_8016);
nor U8191 (N_8191,N_8038,N_8037);
and U8192 (N_8192,N_8033,N_8049);
xor U8193 (N_8193,N_8084,N_8030);
nand U8194 (N_8194,N_8018,N_8117);
and U8195 (N_8195,N_8049,N_8027);
and U8196 (N_8196,N_8114,N_8053);
nand U8197 (N_8197,N_8083,N_8036);
or U8198 (N_8198,N_8001,N_8032);
nor U8199 (N_8199,N_8025,N_8072);
nand U8200 (N_8200,N_8070,N_8052);
nand U8201 (N_8201,N_8008,N_8024);
nand U8202 (N_8202,N_8077,N_8012);
xor U8203 (N_8203,N_8105,N_8066);
nor U8204 (N_8204,N_8093,N_8103);
xor U8205 (N_8205,N_8078,N_8082);
nand U8206 (N_8206,N_8080,N_8081);
nor U8207 (N_8207,N_8099,N_8052);
and U8208 (N_8208,N_8058,N_8056);
nor U8209 (N_8209,N_8058,N_8067);
or U8210 (N_8210,N_8013,N_8042);
or U8211 (N_8211,N_8012,N_8059);
nand U8212 (N_8212,N_8048,N_8072);
and U8213 (N_8213,N_8119,N_8028);
xnor U8214 (N_8214,N_8092,N_8041);
nand U8215 (N_8215,N_8027,N_8045);
and U8216 (N_8216,N_8011,N_8103);
and U8217 (N_8217,N_8074,N_8098);
or U8218 (N_8218,N_8119,N_8103);
or U8219 (N_8219,N_8074,N_8020);
nor U8220 (N_8220,N_8008,N_8111);
and U8221 (N_8221,N_8070,N_8026);
or U8222 (N_8222,N_8093,N_8078);
nand U8223 (N_8223,N_8110,N_8044);
or U8224 (N_8224,N_8026,N_8035);
nor U8225 (N_8225,N_8106,N_8072);
and U8226 (N_8226,N_8074,N_8038);
xor U8227 (N_8227,N_8022,N_8087);
nor U8228 (N_8228,N_8080,N_8002);
or U8229 (N_8229,N_8082,N_8091);
nand U8230 (N_8230,N_8031,N_8098);
xor U8231 (N_8231,N_8120,N_8013);
and U8232 (N_8232,N_8075,N_8083);
and U8233 (N_8233,N_8117,N_8039);
xnor U8234 (N_8234,N_8055,N_8107);
nor U8235 (N_8235,N_8049,N_8104);
or U8236 (N_8236,N_8000,N_8013);
xor U8237 (N_8237,N_8092,N_8089);
and U8238 (N_8238,N_8108,N_8105);
and U8239 (N_8239,N_8111,N_8102);
nand U8240 (N_8240,N_8111,N_8101);
xnor U8241 (N_8241,N_8063,N_8042);
nor U8242 (N_8242,N_8009,N_8104);
and U8243 (N_8243,N_8070,N_8099);
and U8244 (N_8244,N_8043,N_8015);
and U8245 (N_8245,N_8116,N_8062);
nor U8246 (N_8246,N_8071,N_8109);
xor U8247 (N_8247,N_8096,N_8020);
and U8248 (N_8248,N_8059,N_8072);
xnor U8249 (N_8249,N_8099,N_8009);
xor U8250 (N_8250,N_8150,N_8245);
and U8251 (N_8251,N_8142,N_8185);
nor U8252 (N_8252,N_8208,N_8194);
xnor U8253 (N_8253,N_8249,N_8146);
or U8254 (N_8254,N_8139,N_8247);
nand U8255 (N_8255,N_8205,N_8220);
and U8256 (N_8256,N_8243,N_8204);
or U8257 (N_8257,N_8212,N_8132);
nand U8258 (N_8258,N_8157,N_8173);
and U8259 (N_8259,N_8145,N_8129);
xnor U8260 (N_8260,N_8180,N_8154);
or U8261 (N_8261,N_8201,N_8228);
nand U8262 (N_8262,N_8156,N_8223);
and U8263 (N_8263,N_8147,N_8214);
nor U8264 (N_8264,N_8238,N_8234);
and U8265 (N_8265,N_8130,N_8237);
nand U8266 (N_8266,N_8176,N_8239);
xnor U8267 (N_8267,N_8169,N_8141);
nor U8268 (N_8268,N_8203,N_8213);
xnor U8269 (N_8269,N_8198,N_8232);
and U8270 (N_8270,N_8126,N_8192);
nand U8271 (N_8271,N_8226,N_8199);
and U8272 (N_8272,N_8229,N_8174);
nor U8273 (N_8273,N_8227,N_8196);
or U8274 (N_8274,N_8134,N_8159);
and U8275 (N_8275,N_8186,N_8200);
or U8276 (N_8276,N_8191,N_8144);
and U8277 (N_8277,N_8187,N_8155);
nor U8278 (N_8278,N_8182,N_8178);
nand U8279 (N_8279,N_8206,N_8236);
and U8280 (N_8280,N_8143,N_8184);
and U8281 (N_8281,N_8170,N_8193);
xnor U8282 (N_8282,N_8166,N_8222);
nor U8283 (N_8283,N_8165,N_8128);
nor U8284 (N_8284,N_8235,N_8195);
and U8285 (N_8285,N_8211,N_8153);
and U8286 (N_8286,N_8183,N_8127);
or U8287 (N_8287,N_8189,N_8190);
or U8288 (N_8288,N_8244,N_8188);
xnor U8289 (N_8289,N_8241,N_8240);
nand U8290 (N_8290,N_8172,N_8175);
xnor U8291 (N_8291,N_8224,N_8207);
or U8292 (N_8292,N_8160,N_8202);
xor U8293 (N_8293,N_8230,N_8221);
and U8294 (N_8294,N_8177,N_8181);
nand U8295 (N_8295,N_8168,N_8151);
and U8296 (N_8296,N_8162,N_8219);
or U8297 (N_8297,N_8246,N_8218);
nor U8298 (N_8298,N_8179,N_8136);
xor U8299 (N_8299,N_8210,N_8164);
nand U8300 (N_8300,N_8140,N_8233);
xor U8301 (N_8301,N_8248,N_8148);
and U8302 (N_8302,N_8197,N_8137);
or U8303 (N_8303,N_8217,N_8152);
and U8304 (N_8304,N_8131,N_8158);
nor U8305 (N_8305,N_8225,N_8242);
xor U8306 (N_8306,N_8149,N_8138);
nor U8307 (N_8307,N_8216,N_8125);
xor U8308 (N_8308,N_8163,N_8215);
xor U8309 (N_8309,N_8133,N_8135);
nor U8310 (N_8310,N_8161,N_8171);
and U8311 (N_8311,N_8231,N_8209);
nand U8312 (N_8312,N_8167,N_8238);
and U8313 (N_8313,N_8130,N_8240);
and U8314 (N_8314,N_8179,N_8201);
nor U8315 (N_8315,N_8149,N_8132);
or U8316 (N_8316,N_8245,N_8226);
or U8317 (N_8317,N_8169,N_8173);
or U8318 (N_8318,N_8217,N_8130);
and U8319 (N_8319,N_8226,N_8187);
nand U8320 (N_8320,N_8241,N_8220);
and U8321 (N_8321,N_8228,N_8136);
or U8322 (N_8322,N_8230,N_8175);
nor U8323 (N_8323,N_8237,N_8184);
xor U8324 (N_8324,N_8203,N_8125);
and U8325 (N_8325,N_8202,N_8224);
nand U8326 (N_8326,N_8230,N_8200);
nand U8327 (N_8327,N_8188,N_8143);
xor U8328 (N_8328,N_8239,N_8164);
nor U8329 (N_8329,N_8218,N_8153);
and U8330 (N_8330,N_8203,N_8222);
and U8331 (N_8331,N_8201,N_8211);
nand U8332 (N_8332,N_8248,N_8211);
nand U8333 (N_8333,N_8245,N_8222);
nand U8334 (N_8334,N_8166,N_8197);
xnor U8335 (N_8335,N_8202,N_8197);
or U8336 (N_8336,N_8179,N_8199);
nand U8337 (N_8337,N_8159,N_8132);
and U8338 (N_8338,N_8177,N_8147);
or U8339 (N_8339,N_8182,N_8220);
nand U8340 (N_8340,N_8159,N_8145);
xnor U8341 (N_8341,N_8134,N_8158);
nand U8342 (N_8342,N_8158,N_8205);
or U8343 (N_8343,N_8191,N_8229);
nand U8344 (N_8344,N_8185,N_8225);
nor U8345 (N_8345,N_8188,N_8132);
or U8346 (N_8346,N_8174,N_8162);
or U8347 (N_8347,N_8236,N_8164);
xor U8348 (N_8348,N_8139,N_8214);
and U8349 (N_8349,N_8212,N_8242);
and U8350 (N_8350,N_8233,N_8215);
or U8351 (N_8351,N_8221,N_8239);
xor U8352 (N_8352,N_8244,N_8249);
nand U8353 (N_8353,N_8186,N_8248);
or U8354 (N_8354,N_8139,N_8225);
and U8355 (N_8355,N_8240,N_8137);
and U8356 (N_8356,N_8203,N_8237);
nand U8357 (N_8357,N_8177,N_8234);
xnor U8358 (N_8358,N_8149,N_8207);
and U8359 (N_8359,N_8152,N_8149);
and U8360 (N_8360,N_8237,N_8195);
nor U8361 (N_8361,N_8157,N_8145);
and U8362 (N_8362,N_8132,N_8213);
and U8363 (N_8363,N_8238,N_8230);
xor U8364 (N_8364,N_8156,N_8202);
nor U8365 (N_8365,N_8150,N_8184);
nor U8366 (N_8366,N_8234,N_8214);
nand U8367 (N_8367,N_8174,N_8166);
or U8368 (N_8368,N_8242,N_8173);
nor U8369 (N_8369,N_8177,N_8169);
and U8370 (N_8370,N_8135,N_8180);
nand U8371 (N_8371,N_8201,N_8126);
or U8372 (N_8372,N_8179,N_8190);
nand U8373 (N_8373,N_8161,N_8141);
or U8374 (N_8374,N_8197,N_8236);
or U8375 (N_8375,N_8309,N_8288);
nand U8376 (N_8376,N_8266,N_8330);
nor U8377 (N_8377,N_8337,N_8310);
and U8378 (N_8378,N_8278,N_8374);
and U8379 (N_8379,N_8328,N_8301);
nand U8380 (N_8380,N_8324,N_8250);
and U8381 (N_8381,N_8360,N_8368);
and U8382 (N_8382,N_8280,N_8261);
or U8383 (N_8383,N_8274,N_8283);
nand U8384 (N_8384,N_8319,N_8355);
nor U8385 (N_8385,N_8289,N_8326);
nand U8386 (N_8386,N_8264,N_8253);
nand U8387 (N_8387,N_8372,N_8357);
or U8388 (N_8388,N_8300,N_8341);
nor U8389 (N_8389,N_8348,N_8263);
and U8390 (N_8390,N_8363,N_8316);
and U8391 (N_8391,N_8276,N_8292);
nand U8392 (N_8392,N_8268,N_8281);
and U8393 (N_8393,N_8270,N_8318);
nand U8394 (N_8394,N_8255,N_8259);
and U8395 (N_8395,N_8293,N_8313);
nand U8396 (N_8396,N_8359,N_8254);
or U8397 (N_8397,N_8345,N_8339);
and U8398 (N_8398,N_8371,N_8342);
or U8399 (N_8399,N_8267,N_8322);
xnor U8400 (N_8400,N_8251,N_8352);
nand U8401 (N_8401,N_8314,N_8304);
or U8402 (N_8402,N_8344,N_8290);
nor U8403 (N_8403,N_8347,N_8320);
nand U8404 (N_8404,N_8279,N_8362);
and U8405 (N_8405,N_8275,N_8265);
nand U8406 (N_8406,N_8295,N_8336);
and U8407 (N_8407,N_8284,N_8361);
nand U8408 (N_8408,N_8350,N_8269);
nand U8409 (N_8409,N_8356,N_8285);
nand U8410 (N_8410,N_8346,N_8365);
nor U8411 (N_8411,N_8306,N_8305);
nor U8412 (N_8412,N_8277,N_8303);
nor U8413 (N_8413,N_8286,N_8373);
and U8414 (N_8414,N_8351,N_8366);
and U8415 (N_8415,N_8291,N_8358);
nand U8416 (N_8416,N_8367,N_8369);
and U8417 (N_8417,N_8307,N_8312);
nor U8418 (N_8418,N_8332,N_8333);
xor U8419 (N_8419,N_8294,N_8335);
or U8420 (N_8420,N_8299,N_8297);
and U8421 (N_8421,N_8353,N_8354);
nand U8422 (N_8422,N_8331,N_8317);
xnor U8423 (N_8423,N_8272,N_8327);
nand U8424 (N_8424,N_8287,N_8329);
xnor U8425 (N_8425,N_8370,N_8340);
and U8426 (N_8426,N_8321,N_8349);
and U8427 (N_8427,N_8258,N_8260);
or U8428 (N_8428,N_8273,N_8252);
nor U8429 (N_8429,N_8343,N_8334);
xor U8430 (N_8430,N_8296,N_8298);
and U8431 (N_8431,N_8257,N_8256);
xor U8432 (N_8432,N_8311,N_8262);
and U8433 (N_8433,N_8315,N_8302);
nand U8434 (N_8434,N_8338,N_8323);
or U8435 (N_8435,N_8271,N_8282);
and U8436 (N_8436,N_8325,N_8308);
xnor U8437 (N_8437,N_8364,N_8272);
or U8438 (N_8438,N_8336,N_8310);
nand U8439 (N_8439,N_8267,N_8275);
nand U8440 (N_8440,N_8349,N_8326);
or U8441 (N_8441,N_8319,N_8362);
nor U8442 (N_8442,N_8279,N_8357);
and U8443 (N_8443,N_8354,N_8374);
nand U8444 (N_8444,N_8348,N_8284);
and U8445 (N_8445,N_8304,N_8251);
xor U8446 (N_8446,N_8349,N_8256);
xnor U8447 (N_8447,N_8318,N_8260);
and U8448 (N_8448,N_8310,N_8274);
nor U8449 (N_8449,N_8265,N_8308);
nand U8450 (N_8450,N_8373,N_8302);
or U8451 (N_8451,N_8308,N_8296);
and U8452 (N_8452,N_8371,N_8279);
nand U8453 (N_8453,N_8313,N_8308);
xor U8454 (N_8454,N_8343,N_8257);
xnor U8455 (N_8455,N_8324,N_8331);
xor U8456 (N_8456,N_8352,N_8349);
nand U8457 (N_8457,N_8339,N_8355);
xnor U8458 (N_8458,N_8253,N_8268);
nor U8459 (N_8459,N_8322,N_8271);
xnor U8460 (N_8460,N_8315,N_8255);
nand U8461 (N_8461,N_8304,N_8278);
nand U8462 (N_8462,N_8293,N_8364);
xnor U8463 (N_8463,N_8275,N_8320);
nor U8464 (N_8464,N_8275,N_8319);
nor U8465 (N_8465,N_8304,N_8257);
or U8466 (N_8466,N_8344,N_8356);
nor U8467 (N_8467,N_8308,N_8297);
nor U8468 (N_8468,N_8330,N_8303);
nor U8469 (N_8469,N_8262,N_8318);
nand U8470 (N_8470,N_8331,N_8349);
and U8471 (N_8471,N_8315,N_8312);
xnor U8472 (N_8472,N_8267,N_8318);
xor U8473 (N_8473,N_8279,N_8297);
and U8474 (N_8474,N_8364,N_8331);
or U8475 (N_8475,N_8349,N_8257);
and U8476 (N_8476,N_8259,N_8270);
xnor U8477 (N_8477,N_8365,N_8333);
nand U8478 (N_8478,N_8354,N_8258);
and U8479 (N_8479,N_8291,N_8251);
or U8480 (N_8480,N_8363,N_8269);
xor U8481 (N_8481,N_8255,N_8332);
or U8482 (N_8482,N_8270,N_8250);
or U8483 (N_8483,N_8308,N_8290);
nor U8484 (N_8484,N_8302,N_8329);
nand U8485 (N_8485,N_8264,N_8283);
and U8486 (N_8486,N_8253,N_8272);
and U8487 (N_8487,N_8341,N_8321);
xnor U8488 (N_8488,N_8257,N_8360);
nand U8489 (N_8489,N_8270,N_8258);
nand U8490 (N_8490,N_8358,N_8284);
nand U8491 (N_8491,N_8275,N_8353);
or U8492 (N_8492,N_8351,N_8337);
and U8493 (N_8493,N_8334,N_8299);
or U8494 (N_8494,N_8254,N_8356);
xnor U8495 (N_8495,N_8260,N_8351);
xnor U8496 (N_8496,N_8359,N_8336);
and U8497 (N_8497,N_8327,N_8300);
or U8498 (N_8498,N_8281,N_8310);
or U8499 (N_8499,N_8321,N_8294);
nand U8500 (N_8500,N_8428,N_8454);
xnor U8501 (N_8501,N_8495,N_8433);
xnor U8502 (N_8502,N_8473,N_8455);
xor U8503 (N_8503,N_8418,N_8393);
nor U8504 (N_8504,N_8416,N_8499);
nor U8505 (N_8505,N_8389,N_8436);
and U8506 (N_8506,N_8379,N_8440);
nor U8507 (N_8507,N_8470,N_8383);
or U8508 (N_8508,N_8480,N_8442);
nor U8509 (N_8509,N_8391,N_8491);
or U8510 (N_8510,N_8425,N_8384);
nand U8511 (N_8511,N_8435,N_8420);
xor U8512 (N_8512,N_8474,N_8401);
and U8513 (N_8513,N_8479,N_8465);
or U8514 (N_8514,N_8400,N_8478);
or U8515 (N_8515,N_8469,N_8388);
nand U8516 (N_8516,N_8487,N_8419);
nand U8517 (N_8517,N_8381,N_8430);
nor U8518 (N_8518,N_8498,N_8459);
nor U8519 (N_8519,N_8458,N_8407);
xnor U8520 (N_8520,N_8394,N_8448);
nor U8521 (N_8521,N_8444,N_8405);
xor U8522 (N_8522,N_8446,N_8457);
or U8523 (N_8523,N_8386,N_8408);
and U8524 (N_8524,N_8481,N_8493);
nand U8525 (N_8525,N_8378,N_8490);
or U8526 (N_8526,N_8464,N_8421);
and U8527 (N_8527,N_8392,N_8467);
nand U8528 (N_8528,N_8441,N_8427);
and U8529 (N_8529,N_8443,N_8417);
xnor U8530 (N_8530,N_8376,N_8486);
nand U8531 (N_8531,N_8380,N_8438);
or U8532 (N_8532,N_8468,N_8377);
and U8533 (N_8533,N_8496,N_8375);
and U8534 (N_8534,N_8456,N_8434);
and U8535 (N_8535,N_8385,N_8426);
xnor U8536 (N_8536,N_8382,N_8414);
or U8537 (N_8537,N_8453,N_8462);
nor U8538 (N_8538,N_8452,N_8409);
nor U8539 (N_8539,N_8399,N_8396);
or U8540 (N_8540,N_8411,N_8424);
nand U8541 (N_8541,N_8494,N_8492);
and U8542 (N_8542,N_8398,N_8484);
xor U8543 (N_8543,N_8403,N_8463);
nand U8544 (N_8544,N_8466,N_8497);
nor U8545 (N_8545,N_8475,N_8423);
xnor U8546 (N_8546,N_8429,N_8402);
nor U8547 (N_8547,N_8395,N_8445);
nor U8548 (N_8548,N_8476,N_8413);
nand U8549 (N_8549,N_8422,N_8449);
and U8550 (N_8550,N_8431,N_8483);
or U8551 (N_8551,N_8397,N_8477);
nand U8552 (N_8552,N_8415,N_8404);
or U8553 (N_8553,N_8485,N_8461);
xor U8554 (N_8554,N_8412,N_8482);
xor U8555 (N_8555,N_8460,N_8387);
xnor U8556 (N_8556,N_8471,N_8437);
and U8557 (N_8557,N_8472,N_8406);
or U8558 (N_8558,N_8488,N_8390);
xor U8559 (N_8559,N_8410,N_8432);
nand U8560 (N_8560,N_8447,N_8489);
nand U8561 (N_8561,N_8451,N_8450);
nand U8562 (N_8562,N_8439,N_8453);
xor U8563 (N_8563,N_8486,N_8396);
xnor U8564 (N_8564,N_8427,N_8478);
or U8565 (N_8565,N_8438,N_8436);
xor U8566 (N_8566,N_8423,N_8451);
and U8567 (N_8567,N_8396,N_8449);
nor U8568 (N_8568,N_8441,N_8434);
nor U8569 (N_8569,N_8401,N_8452);
and U8570 (N_8570,N_8453,N_8416);
nand U8571 (N_8571,N_8442,N_8383);
and U8572 (N_8572,N_8481,N_8476);
and U8573 (N_8573,N_8408,N_8464);
and U8574 (N_8574,N_8417,N_8467);
nor U8575 (N_8575,N_8434,N_8463);
or U8576 (N_8576,N_8379,N_8419);
or U8577 (N_8577,N_8440,N_8382);
xor U8578 (N_8578,N_8485,N_8497);
xor U8579 (N_8579,N_8419,N_8435);
and U8580 (N_8580,N_8470,N_8401);
nand U8581 (N_8581,N_8408,N_8431);
nor U8582 (N_8582,N_8407,N_8497);
nand U8583 (N_8583,N_8440,N_8409);
xor U8584 (N_8584,N_8386,N_8395);
nor U8585 (N_8585,N_8472,N_8411);
or U8586 (N_8586,N_8389,N_8420);
xor U8587 (N_8587,N_8404,N_8455);
xor U8588 (N_8588,N_8403,N_8451);
or U8589 (N_8589,N_8472,N_8385);
nand U8590 (N_8590,N_8431,N_8437);
nand U8591 (N_8591,N_8431,N_8423);
and U8592 (N_8592,N_8379,N_8475);
and U8593 (N_8593,N_8454,N_8471);
or U8594 (N_8594,N_8442,N_8396);
nor U8595 (N_8595,N_8495,N_8481);
xor U8596 (N_8596,N_8437,N_8440);
or U8597 (N_8597,N_8412,N_8392);
xor U8598 (N_8598,N_8447,N_8410);
or U8599 (N_8599,N_8450,N_8480);
xor U8600 (N_8600,N_8377,N_8491);
and U8601 (N_8601,N_8497,N_8384);
xnor U8602 (N_8602,N_8448,N_8395);
nand U8603 (N_8603,N_8450,N_8401);
nor U8604 (N_8604,N_8441,N_8398);
nand U8605 (N_8605,N_8390,N_8410);
nand U8606 (N_8606,N_8412,N_8375);
xnor U8607 (N_8607,N_8435,N_8434);
xor U8608 (N_8608,N_8426,N_8389);
xor U8609 (N_8609,N_8425,N_8467);
nand U8610 (N_8610,N_8398,N_8419);
nand U8611 (N_8611,N_8378,N_8405);
or U8612 (N_8612,N_8467,N_8470);
or U8613 (N_8613,N_8467,N_8463);
and U8614 (N_8614,N_8424,N_8377);
and U8615 (N_8615,N_8431,N_8418);
xnor U8616 (N_8616,N_8398,N_8438);
or U8617 (N_8617,N_8426,N_8392);
xor U8618 (N_8618,N_8376,N_8441);
and U8619 (N_8619,N_8445,N_8402);
xor U8620 (N_8620,N_8451,N_8441);
nand U8621 (N_8621,N_8495,N_8415);
and U8622 (N_8622,N_8456,N_8469);
nand U8623 (N_8623,N_8481,N_8416);
nor U8624 (N_8624,N_8478,N_8409);
xnor U8625 (N_8625,N_8556,N_8545);
xnor U8626 (N_8626,N_8618,N_8572);
nand U8627 (N_8627,N_8560,N_8519);
nand U8628 (N_8628,N_8528,N_8523);
and U8629 (N_8629,N_8579,N_8501);
xor U8630 (N_8630,N_8580,N_8571);
xnor U8631 (N_8631,N_8614,N_8553);
xor U8632 (N_8632,N_8540,N_8623);
xnor U8633 (N_8633,N_8596,N_8589);
and U8634 (N_8634,N_8535,N_8537);
or U8635 (N_8635,N_8550,N_8610);
or U8636 (N_8636,N_8597,N_8508);
xnor U8637 (N_8637,N_8506,N_8557);
and U8638 (N_8638,N_8539,N_8500);
xnor U8639 (N_8639,N_8530,N_8543);
or U8640 (N_8640,N_8600,N_8593);
and U8641 (N_8641,N_8541,N_8598);
nor U8642 (N_8642,N_8536,N_8559);
or U8643 (N_8643,N_8564,N_8522);
and U8644 (N_8644,N_8511,N_8554);
xnor U8645 (N_8645,N_8576,N_8574);
or U8646 (N_8646,N_8521,N_8585);
or U8647 (N_8647,N_8590,N_8599);
nand U8648 (N_8648,N_8586,N_8581);
or U8649 (N_8649,N_8578,N_8616);
and U8650 (N_8650,N_8575,N_8547);
and U8651 (N_8651,N_8617,N_8513);
nor U8652 (N_8652,N_8620,N_8619);
or U8653 (N_8653,N_8515,N_8551);
and U8654 (N_8654,N_8504,N_8605);
or U8655 (N_8655,N_8569,N_8505);
nor U8656 (N_8656,N_8549,N_8567);
nand U8657 (N_8657,N_8507,N_8516);
nor U8658 (N_8658,N_8583,N_8529);
nand U8659 (N_8659,N_8622,N_8573);
and U8660 (N_8660,N_8518,N_8595);
or U8661 (N_8661,N_8588,N_8555);
and U8662 (N_8662,N_8594,N_8612);
and U8663 (N_8663,N_8538,N_8608);
xor U8664 (N_8664,N_8558,N_8532);
and U8665 (N_8665,N_8542,N_8565);
nand U8666 (N_8666,N_8591,N_8624);
or U8667 (N_8667,N_8603,N_8602);
xor U8668 (N_8668,N_8517,N_8606);
nor U8669 (N_8669,N_8503,N_8604);
nand U8670 (N_8670,N_8531,N_8568);
nand U8671 (N_8671,N_8566,N_8607);
xor U8672 (N_8672,N_8527,N_8562);
and U8673 (N_8673,N_8544,N_8611);
or U8674 (N_8674,N_8548,N_8520);
and U8675 (N_8675,N_8524,N_8533);
nand U8676 (N_8676,N_8514,N_8552);
nor U8677 (N_8677,N_8502,N_8509);
nor U8678 (N_8678,N_8512,N_8534);
or U8679 (N_8679,N_8546,N_8592);
nand U8680 (N_8680,N_8584,N_8570);
nor U8681 (N_8681,N_8587,N_8615);
and U8682 (N_8682,N_8561,N_8601);
nand U8683 (N_8683,N_8621,N_8582);
nand U8684 (N_8684,N_8577,N_8526);
xor U8685 (N_8685,N_8563,N_8613);
nor U8686 (N_8686,N_8525,N_8510);
xor U8687 (N_8687,N_8609,N_8541);
xor U8688 (N_8688,N_8583,N_8570);
or U8689 (N_8689,N_8581,N_8561);
or U8690 (N_8690,N_8551,N_8574);
xor U8691 (N_8691,N_8606,N_8616);
nor U8692 (N_8692,N_8540,N_8573);
xor U8693 (N_8693,N_8603,N_8561);
or U8694 (N_8694,N_8566,N_8510);
nand U8695 (N_8695,N_8590,N_8546);
nor U8696 (N_8696,N_8501,N_8525);
xor U8697 (N_8697,N_8545,N_8521);
or U8698 (N_8698,N_8548,N_8621);
nand U8699 (N_8699,N_8612,N_8582);
xnor U8700 (N_8700,N_8552,N_8570);
nor U8701 (N_8701,N_8591,N_8598);
xnor U8702 (N_8702,N_8569,N_8555);
or U8703 (N_8703,N_8517,N_8504);
or U8704 (N_8704,N_8604,N_8507);
or U8705 (N_8705,N_8600,N_8616);
and U8706 (N_8706,N_8532,N_8572);
nor U8707 (N_8707,N_8507,N_8596);
nand U8708 (N_8708,N_8590,N_8501);
or U8709 (N_8709,N_8598,N_8536);
nand U8710 (N_8710,N_8541,N_8550);
and U8711 (N_8711,N_8551,N_8555);
xor U8712 (N_8712,N_8568,N_8600);
xor U8713 (N_8713,N_8529,N_8538);
or U8714 (N_8714,N_8584,N_8551);
nor U8715 (N_8715,N_8573,N_8530);
nor U8716 (N_8716,N_8576,N_8621);
and U8717 (N_8717,N_8618,N_8556);
xor U8718 (N_8718,N_8558,N_8588);
nand U8719 (N_8719,N_8550,N_8590);
xor U8720 (N_8720,N_8521,N_8592);
and U8721 (N_8721,N_8536,N_8620);
xor U8722 (N_8722,N_8502,N_8608);
nor U8723 (N_8723,N_8562,N_8572);
nor U8724 (N_8724,N_8538,N_8589);
and U8725 (N_8725,N_8540,N_8571);
nor U8726 (N_8726,N_8544,N_8543);
or U8727 (N_8727,N_8578,N_8567);
nor U8728 (N_8728,N_8503,N_8552);
and U8729 (N_8729,N_8602,N_8595);
and U8730 (N_8730,N_8525,N_8537);
and U8731 (N_8731,N_8519,N_8606);
and U8732 (N_8732,N_8521,N_8614);
and U8733 (N_8733,N_8536,N_8519);
or U8734 (N_8734,N_8535,N_8576);
or U8735 (N_8735,N_8566,N_8500);
nor U8736 (N_8736,N_8554,N_8517);
and U8737 (N_8737,N_8593,N_8607);
and U8738 (N_8738,N_8500,N_8542);
nand U8739 (N_8739,N_8553,N_8577);
nor U8740 (N_8740,N_8618,N_8623);
xor U8741 (N_8741,N_8513,N_8551);
nor U8742 (N_8742,N_8514,N_8585);
and U8743 (N_8743,N_8610,N_8587);
and U8744 (N_8744,N_8513,N_8527);
and U8745 (N_8745,N_8528,N_8576);
xnor U8746 (N_8746,N_8609,N_8580);
and U8747 (N_8747,N_8514,N_8607);
xnor U8748 (N_8748,N_8550,N_8509);
nand U8749 (N_8749,N_8552,N_8580);
xor U8750 (N_8750,N_8631,N_8721);
nand U8751 (N_8751,N_8724,N_8715);
nor U8752 (N_8752,N_8668,N_8705);
xor U8753 (N_8753,N_8704,N_8625);
and U8754 (N_8754,N_8744,N_8656);
nor U8755 (N_8755,N_8741,N_8711);
nor U8756 (N_8756,N_8740,N_8722);
xnor U8757 (N_8757,N_8676,N_8720);
or U8758 (N_8758,N_8727,N_8701);
or U8759 (N_8759,N_8695,N_8717);
and U8760 (N_8760,N_8641,N_8742);
or U8761 (N_8761,N_8645,N_8633);
nor U8762 (N_8762,N_8636,N_8630);
xor U8763 (N_8763,N_8643,N_8700);
nand U8764 (N_8764,N_8658,N_8670);
nand U8765 (N_8765,N_8659,N_8710);
nand U8766 (N_8766,N_8638,N_8708);
xnor U8767 (N_8767,N_8657,N_8689);
nand U8768 (N_8768,N_8714,N_8647);
xor U8769 (N_8769,N_8648,N_8665);
or U8770 (N_8770,N_8679,N_8719);
nand U8771 (N_8771,N_8640,N_8652);
or U8772 (N_8772,N_8716,N_8639);
nand U8773 (N_8773,N_8671,N_8677);
and U8774 (N_8774,N_8733,N_8726);
xor U8775 (N_8775,N_8650,N_8687);
and U8776 (N_8776,N_8725,N_8669);
and U8777 (N_8777,N_8694,N_8735);
xnor U8778 (N_8778,N_8723,N_8709);
nand U8779 (N_8779,N_8749,N_8731);
nor U8780 (N_8780,N_8651,N_8682);
xor U8781 (N_8781,N_8745,N_8626);
nor U8782 (N_8782,N_8748,N_8692);
or U8783 (N_8783,N_8703,N_8667);
xnor U8784 (N_8784,N_8663,N_8678);
and U8785 (N_8785,N_8644,N_8662);
nand U8786 (N_8786,N_8699,N_8718);
nor U8787 (N_8787,N_8693,N_8642);
xor U8788 (N_8788,N_8734,N_8673);
nand U8789 (N_8789,N_8681,N_8684);
nor U8790 (N_8790,N_8702,N_8696);
and U8791 (N_8791,N_8736,N_8634);
nand U8792 (N_8792,N_8738,N_8632);
and U8793 (N_8793,N_8646,N_8675);
xnor U8794 (N_8794,N_8664,N_8649);
xor U8795 (N_8795,N_8686,N_8747);
nor U8796 (N_8796,N_8674,N_8712);
xnor U8797 (N_8797,N_8629,N_8728);
or U8798 (N_8798,N_8661,N_8730);
or U8799 (N_8799,N_8729,N_8706);
nand U8800 (N_8800,N_8698,N_8628);
or U8801 (N_8801,N_8666,N_8697);
and U8802 (N_8802,N_8680,N_8732);
nor U8803 (N_8803,N_8683,N_8672);
xnor U8804 (N_8804,N_8660,N_8743);
and U8805 (N_8805,N_8713,N_8688);
and U8806 (N_8806,N_8690,N_8637);
xnor U8807 (N_8807,N_8635,N_8746);
and U8808 (N_8808,N_8627,N_8707);
xnor U8809 (N_8809,N_8737,N_8739);
xnor U8810 (N_8810,N_8685,N_8654);
nor U8811 (N_8811,N_8691,N_8655);
xor U8812 (N_8812,N_8653,N_8634);
xnor U8813 (N_8813,N_8657,N_8672);
nand U8814 (N_8814,N_8710,N_8636);
xor U8815 (N_8815,N_8687,N_8651);
nand U8816 (N_8816,N_8647,N_8641);
nor U8817 (N_8817,N_8741,N_8745);
or U8818 (N_8818,N_8701,N_8675);
and U8819 (N_8819,N_8660,N_8722);
nor U8820 (N_8820,N_8633,N_8626);
xnor U8821 (N_8821,N_8669,N_8740);
nand U8822 (N_8822,N_8721,N_8692);
and U8823 (N_8823,N_8633,N_8684);
nand U8824 (N_8824,N_8696,N_8664);
or U8825 (N_8825,N_8667,N_8677);
or U8826 (N_8826,N_8741,N_8685);
nand U8827 (N_8827,N_8660,N_8668);
nor U8828 (N_8828,N_8734,N_8706);
xor U8829 (N_8829,N_8662,N_8645);
or U8830 (N_8830,N_8680,N_8648);
nor U8831 (N_8831,N_8722,N_8643);
nor U8832 (N_8832,N_8638,N_8717);
nor U8833 (N_8833,N_8746,N_8664);
nand U8834 (N_8834,N_8673,N_8711);
nand U8835 (N_8835,N_8660,N_8747);
and U8836 (N_8836,N_8707,N_8659);
and U8837 (N_8837,N_8645,N_8715);
or U8838 (N_8838,N_8686,N_8657);
and U8839 (N_8839,N_8741,N_8719);
or U8840 (N_8840,N_8671,N_8645);
or U8841 (N_8841,N_8692,N_8651);
xor U8842 (N_8842,N_8724,N_8730);
nor U8843 (N_8843,N_8657,N_8713);
xnor U8844 (N_8844,N_8693,N_8663);
and U8845 (N_8845,N_8632,N_8663);
nor U8846 (N_8846,N_8678,N_8664);
nor U8847 (N_8847,N_8667,N_8627);
or U8848 (N_8848,N_8629,N_8681);
and U8849 (N_8849,N_8634,N_8638);
and U8850 (N_8850,N_8662,N_8748);
xnor U8851 (N_8851,N_8746,N_8738);
nor U8852 (N_8852,N_8672,N_8696);
nor U8853 (N_8853,N_8659,N_8655);
nand U8854 (N_8854,N_8732,N_8676);
and U8855 (N_8855,N_8629,N_8668);
nor U8856 (N_8856,N_8746,N_8628);
nand U8857 (N_8857,N_8665,N_8748);
xnor U8858 (N_8858,N_8664,N_8637);
or U8859 (N_8859,N_8743,N_8741);
xor U8860 (N_8860,N_8712,N_8633);
xor U8861 (N_8861,N_8707,N_8736);
nor U8862 (N_8862,N_8707,N_8671);
or U8863 (N_8863,N_8684,N_8678);
and U8864 (N_8864,N_8647,N_8693);
nand U8865 (N_8865,N_8724,N_8629);
or U8866 (N_8866,N_8728,N_8685);
nor U8867 (N_8867,N_8646,N_8727);
or U8868 (N_8868,N_8711,N_8667);
or U8869 (N_8869,N_8708,N_8712);
or U8870 (N_8870,N_8742,N_8635);
xnor U8871 (N_8871,N_8729,N_8629);
or U8872 (N_8872,N_8731,N_8745);
xnor U8873 (N_8873,N_8733,N_8654);
xor U8874 (N_8874,N_8731,N_8628);
or U8875 (N_8875,N_8833,N_8815);
nor U8876 (N_8876,N_8864,N_8769);
xnor U8877 (N_8877,N_8844,N_8836);
nor U8878 (N_8878,N_8859,N_8862);
xor U8879 (N_8879,N_8755,N_8814);
xor U8880 (N_8880,N_8783,N_8856);
nand U8881 (N_8881,N_8792,N_8820);
nor U8882 (N_8882,N_8763,N_8758);
nand U8883 (N_8883,N_8826,N_8781);
or U8884 (N_8884,N_8824,N_8766);
nor U8885 (N_8885,N_8762,N_8772);
or U8886 (N_8886,N_8838,N_8757);
xnor U8887 (N_8887,N_8827,N_8865);
and U8888 (N_8888,N_8837,N_8840);
or U8889 (N_8889,N_8795,N_8846);
or U8890 (N_8890,N_8855,N_8872);
or U8891 (N_8891,N_8848,N_8776);
and U8892 (N_8892,N_8871,N_8835);
and U8893 (N_8893,N_8851,N_8804);
nor U8894 (N_8894,N_8797,N_8828);
xor U8895 (N_8895,N_8812,N_8760);
xor U8896 (N_8896,N_8765,N_8782);
nor U8897 (N_8897,N_8800,N_8832);
and U8898 (N_8898,N_8759,N_8816);
or U8899 (N_8899,N_8813,N_8809);
nand U8900 (N_8900,N_8866,N_8869);
nand U8901 (N_8901,N_8790,N_8778);
nor U8902 (N_8902,N_8863,N_8791);
xor U8903 (N_8903,N_8806,N_8775);
and U8904 (N_8904,N_8874,N_8761);
and U8905 (N_8905,N_8798,N_8839);
xor U8906 (N_8906,N_8794,N_8787);
nor U8907 (N_8907,N_8857,N_8850);
nor U8908 (N_8908,N_8852,N_8785);
nand U8909 (N_8909,N_8829,N_8845);
or U8910 (N_8910,N_8831,N_8788);
nand U8911 (N_8911,N_8842,N_8751);
nor U8912 (N_8912,N_8823,N_8768);
nand U8913 (N_8913,N_8860,N_8771);
and U8914 (N_8914,N_8818,N_8841);
or U8915 (N_8915,N_8764,N_8817);
or U8916 (N_8916,N_8796,N_8822);
nand U8917 (N_8917,N_8861,N_8853);
xnor U8918 (N_8918,N_8805,N_8784);
or U8919 (N_8919,N_8801,N_8793);
xor U8920 (N_8920,N_8807,N_8867);
and U8921 (N_8921,N_8779,N_8750);
or U8922 (N_8922,N_8854,N_8858);
nand U8923 (N_8923,N_8780,N_8803);
or U8924 (N_8924,N_8808,N_8777);
xnor U8925 (N_8925,N_8786,N_8834);
or U8926 (N_8926,N_8756,N_8870);
nor U8927 (N_8927,N_8821,N_8847);
nor U8928 (N_8928,N_8819,N_8810);
and U8929 (N_8929,N_8811,N_8752);
or U8930 (N_8930,N_8873,N_8773);
or U8931 (N_8931,N_8789,N_8754);
xnor U8932 (N_8932,N_8825,N_8799);
and U8933 (N_8933,N_8770,N_8774);
nand U8934 (N_8934,N_8843,N_8767);
nand U8935 (N_8935,N_8753,N_8802);
xor U8936 (N_8936,N_8849,N_8868);
or U8937 (N_8937,N_8830,N_8858);
nor U8938 (N_8938,N_8857,N_8856);
xor U8939 (N_8939,N_8831,N_8783);
xor U8940 (N_8940,N_8838,N_8840);
nand U8941 (N_8941,N_8770,N_8871);
or U8942 (N_8942,N_8780,N_8841);
and U8943 (N_8943,N_8852,N_8805);
and U8944 (N_8944,N_8801,N_8769);
or U8945 (N_8945,N_8867,N_8780);
nand U8946 (N_8946,N_8871,N_8760);
and U8947 (N_8947,N_8771,N_8852);
nand U8948 (N_8948,N_8825,N_8769);
xnor U8949 (N_8949,N_8846,N_8858);
nand U8950 (N_8950,N_8836,N_8751);
nand U8951 (N_8951,N_8845,N_8779);
nand U8952 (N_8952,N_8806,N_8821);
and U8953 (N_8953,N_8801,N_8835);
and U8954 (N_8954,N_8860,N_8775);
or U8955 (N_8955,N_8835,N_8772);
nor U8956 (N_8956,N_8778,N_8817);
xor U8957 (N_8957,N_8802,N_8861);
nand U8958 (N_8958,N_8757,N_8794);
xor U8959 (N_8959,N_8798,N_8755);
nand U8960 (N_8960,N_8870,N_8805);
and U8961 (N_8961,N_8835,N_8800);
xnor U8962 (N_8962,N_8790,N_8795);
or U8963 (N_8963,N_8855,N_8823);
nor U8964 (N_8964,N_8817,N_8854);
or U8965 (N_8965,N_8867,N_8775);
nand U8966 (N_8966,N_8778,N_8874);
xnor U8967 (N_8967,N_8856,N_8806);
nor U8968 (N_8968,N_8750,N_8864);
nor U8969 (N_8969,N_8759,N_8847);
and U8970 (N_8970,N_8784,N_8782);
or U8971 (N_8971,N_8834,N_8849);
xor U8972 (N_8972,N_8776,N_8780);
or U8973 (N_8973,N_8807,N_8819);
and U8974 (N_8974,N_8815,N_8853);
and U8975 (N_8975,N_8814,N_8874);
and U8976 (N_8976,N_8778,N_8777);
or U8977 (N_8977,N_8856,N_8837);
nor U8978 (N_8978,N_8841,N_8839);
nand U8979 (N_8979,N_8758,N_8803);
nor U8980 (N_8980,N_8845,N_8818);
or U8981 (N_8981,N_8761,N_8838);
or U8982 (N_8982,N_8780,N_8840);
and U8983 (N_8983,N_8869,N_8857);
nor U8984 (N_8984,N_8772,N_8827);
and U8985 (N_8985,N_8827,N_8871);
and U8986 (N_8986,N_8761,N_8830);
or U8987 (N_8987,N_8825,N_8797);
nor U8988 (N_8988,N_8811,N_8830);
and U8989 (N_8989,N_8858,N_8827);
and U8990 (N_8990,N_8783,N_8829);
xnor U8991 (N_8991,N_8767,N_8834);
or U8992 (N_8992,N_8787,N_8830);
and U8993 (N_8993,N_8786,N_8845);
and U8994 (N_8994,N_8831,N_8841);
nand U8995 (N_8995,N_8802,N_8830);
xor U8996 (N_8996,N_8813,N_8841);
or U8997 (N_8997,N_8843,N_8793);
xnor U8998 (N_8998,N_8840,N_8760);
xor U8999 (N_8999,N_8863,N_8769);
or U9000 (N_9000,N_8884,N_8957);
xor U9001 (N_9001,N_8951,N_8988);
nor U9002 (N_9002,N_8992,N_8907);
nand U9003 (N_9003,N_8999,N_8952);
nor U9004 (N_9004,N_8985,N_8970);
and U9005 (N_9005,N_8955,N_8904);
xnor U9006 (N_9006,N_8891,N_8886);
nand U9007 (N_9007,N_8950,N_8944);
and U9008 (N_9008,N_8989,N_8905);
xor U9009 (N_9009,N_8991,N_8896);
xnor U9010 (N_9010,N_8908,N_8926);
and U9011 (N_9011,N_8946,N_8978);
and U9012 (N_9012,N_8986,N_8880);
and U9013 (N_9013,N_8960,N_8958);
nor U9014 (N_9014,N_8943,N_8897);
xor U9015 (N_9015,N_8939,N_8912);
nor U9016 (N_9016,N_8878,N_8979);
xnor U9017 (N_9017,N_8913,N_8882);
and U9018 (N_9018,N_8877,N_8935);
nand U9019 (N_9019,N_8929,N_8928);
xnor U9020 (N_9020,N_8881,N_8888);
nor U9021 (N_9021,N_8964,N_8915);
nand U9022 (N_9022,N_8909,N_8971);
or U9023 (N_9023,N_8981,N_8920);
nor U9024 (N_9024,N_8996,N_8901);
nand U9025 (N_9025,N_8953,N_8900);
nor U9026 (N_9026,N_8932,N_8956);
xnor U9027 (N_9027,N_8947,N_8889);
xor U9028 (N_9028,N_8919,N_8954);
nor U9029 (N_9029,N_8910,N_8994);
and U9030 (N_9030,N_8948,N_8937);
xor U9031 (N_9031,N_8895,N_8914);
nor U9032 (N_9032,N_8893,N_8906);
nand U9033 (N_9033,N_8990,N_8975);
nor U9034 (N_9034,N_8973,N_8961);
nor U9035 (N_9035,N_8918,N_8976);
nor U9036 (N_9036,N_8942,N_8892);
xor U9037 (N_9037,N_8945,N_8902);
or U9038 (N_9038,N_8894,N_8899);
and U9039 (N_9039,N_8917,N_8998);
nor U9040 (N_9040,N_8883,N_8966);
and U9041 (N_9041,N_8974,N_8982);
xnor U9042 (N_9042,N_8940,N_8969);
nand U9043 (N_9043,N_8938,N_8890);
nand U9044 (N_9044,N_8887,N_8987);
nor U9045 (N_9045,N_8925,N_8924);
or U9046 (N_9046,N_8927,N_8977);
nor U9047 (N_9047,N_8993,N_8941);
nor U9048 (N_9048,N_8963,N_8879);
xnor U9049 (N_9049,N_8922,N_8876);
or U9050 (N_9050,N_8875,N_8923);
xnor U9051 (N_9051,N_8934,N_8898);
xor U9052 (N_9052,N_8931,N_8968);
and U9053 (N_9053,N_8949,N_8959);
nand U9054 (N_9054,N_8936,N_8962);
nand U9055 (N_9055,N_8997,N_8921);
and U9056 (N_9056,N_8984,N_8995);
xor U9057 (N_9057,N_8980,N_8885);
and U9058 (N_9058,N_8933,N_8930);
and U9059 (N_9059,N_8972,N_8967);
or U9060 (N_9060,N_8903,N_8916);
xor U9061 (N_9061,N_8911,N_8965);
or U9062 (N_9062,N_8983,N_8885);
xor U9063 (N_9063,N_8974,N_8989);
nor U9064 (N_9064,N_8993,N_8890);
and U9065 (N_9065,N_8982,N_8882);
nor U9066 (N_9066,N_8916,N_8892);
xor U9067 (N_9067,N_8979,N_8903);
or U9068 (N_9068,N_8944,N_8909);
nor U9069 (N_9069,N_8900,N_8992);
or U9070 (N_9070,N_8907,N_8938);
or U9071 (N_9071,N_8998,N_8925);
and U9072 (N_9072,N_8970,N_8978);
and U9073 (N_9073,N_8970,N_8920);
xor U9074 (N_9074,N_8957,N_8973);
nand U9075 (N_9075,N_8894,N_8950);
and U9076 (N_9076,N_8938,N_8944);
nand U9077 (N_9077,N_8895,N_8989);
or U9078 (N_9078,N_8914,N_8908);
or U9079 (N_9079,N_8920,N_8875);
and U9080 (N_9080,N_8980,N_8975);
xor U9081 (N_9081,N_8967,N_8944);
and U9082 (N_9082,N_8994,N_8988);
or U9083 (N_9083,N_8899,N_8917);
and U9084 (N_9084,N_8880,N_8966);
or U9085 (N_9085,N_8959,N_8884);
and U9086 (N_9086,N_8906,N_8967);
and U9087 (N_9087,N_8985,N_8922);
xnor U9088 (N_9088,N_8986,N_8876);
and U9089 (N_9089,N_8933,N_8957);
xor U9090 (N_9090,N_8885,N_8981);
nand U9091 (N_9091,N_8989,N_8941);
nand U9092 (N_9092,N_8911,N_8923);
nand U9093 (N_9093,N_8906,N_8909);
xor U9094 (N_9094,N_8891,N_8961);
or U9095 (N_9095,N_8946,N_8921);
nor U9096 (N_9096,N_8902,N_8968);
xor U9097 (N_9097,N_8921,N_8905);
or U9098 (N_9098,N_8982,N_8907);
or U9099 (N_9099,N_8929,N_8911);
and U9100 (N_9100,N_8908,N_8918);
nand U9101 (N_9101,N_8951,N_8973);
xor U9102 (N_9102,N_8990,N_8877);
nand U9103 (N_9103,N_8910,N_8934);
nand U9104 (N_9104,N_8931,N_8927);
xnor U9105 (N_9105,N_8984,N_8972);
and U9106 (N_9106,N_8935,N_8951);
nor U9107 (N_9107,N_8886,N_8908);
nand U9108 (N_9108,N_8950,N_8994);
nor U9109 (N_9109,N_8962,N_8924);
or U9110 (N_9110,N_8888,N_8913);
or U9111 (N_9111,N_8900,N_8972);
xnor U9112 (N_9112,N_8993,N_8900);
or U9113 (N_9113,N_8981,N_8933);
nand U9114 (N_9114,N_8997,N_8951);
or U9115 (N_9115,N_8967,N_8879);
nand U9116 (N_9116,N_8926,N_8876);
and U9117 (N_9117,N_8998,N_8965);
nor U9118 (N_9118,N_8889,N_8953);
and U9119 (N_9119,N_8900,N_8901);
nor U9120 (N_9120,N_8967,N_8988);
and U9121 (N_9121,N_8978,N_8996);
nor U9122 (N_9122,N_8929,N_8948);
nor U9123 (N_9123,N_8910,N_8954);
nand U9124 (N_9124,N_8984,N_8960);
or U9125 (N_9125,N_9040,N_9021);
nor U9126 (N_9126,N_9063,N_9103);
and U9127 (N_9127,N_9037,N_9000);
xor U9128 (N_9128,N_9062,N_9032);
xor U9129 (N_9129,N_9115,N_9016);
nand U9130 (N_9130,N_9100,N_9017);
nor U9131 (N_9131,N_9117,N_9005);
nor U9132 (N_9132,N_9048,N_9084);
and U9133 (N_9133,N_9041,N_9098);
and U9134 (N_9134,N_9038,N_9124);
nor U9135 (N_9135,N_9045,N_9047);
nor U9136 (N_9136,N_9093,N_9061);
xnor U9137 (N_9137,N_9009,N_9057);
xnor U9138 (N_9138,N_9008,N_9027);
and U9139 (N_9139,N_9086,N_9119);
or U9140 (N_9140,N_9044,N_9050);
or U9141 (N_9141,N_9108,N_9074);
nand U9142 (N_9142,N_9043,N_9014);
xor U9143 (N_9143,N_9035,N_9122);
and U9144 (N_9144,N_9089,N_9055);
nor U9145 (N_9145,N_9070,N_9054);
nand U9146 (N_9146,N_9011,N_9007);
xor U9147 (N_9147,N_9082,N_9002);
and U9148 (N_9148,N_9022,N_9034);
nor U9149 (N_9149,N_9091,N_9097);
nor U9150 (N_9150,N_9026,N_9118);
or U9151 (N_9151,N_9042,N_9099);
or U9152 (N_9152,N_9107,N_9023);
nand U9153 (N_9153,N_9109,N_9024);
and U9154 (N_9154,N_9104,N_9094);
xnor U9155 (N_9155,N_9003,N_9033);
or U9156 (N_9156,N_9006,N_9036);
xnor U9157 (N_9157,N_9114,N_9105);
xnor U9158 (N_9158,N_9113,N_9073);
nor U9159 (N_9159,N_9081,N_9090);
or U9160 (N_9160,N_9092,N_9053);
xnor U9161 (N_9161,N_9101,N_9076);
xor U9162 (N_9162,N_9001,N_9088);
nand U9163 (N_9163,N_9039,N_9064);
xnor U9164 (N_9164,N_9067,N_9010);
xnor U9165 (N_9165,N_9075,N_9065);
nor U9166 (N_9166,N_9060,N_9110);
and U9167 (N_9167,N_9078,N_9020);
and U9168 (N_9168,N_9019,N_9112);
and U9169 (N_9169,N_9085,N_9087);
nand U9170 (N_9170,N_9051,N_9012);
and U9171 (N_9171,N_9072,N_9049);
nand U9172 (N_9172,N_9015,N_9079);
or U9173 (N_9173,N_9077,N_9068);
nor U9174 (N_9174,N_9059,N_9030);
nor U9175 (N_9175,N_9116,N_9004);
and U9176 (N_9176,N_9028,N_9120);
or U9177 (N_9177,N_9111,N_9018);
nand U9178 (N_9178,N_9121,N_9066);
or U9179 (N_9179,N_9106,N_9052);
nand U9180 (N_9180,N_9046,N_9029);
xor U9181 (N_9181,N_9056,N_9095);
nor U9182 (N_9182,N_9102,N_9083);
or U9183 (N_9183,N_9069,N_9031);
or U9184 (N_9184,N_9013,N_9071);
nor U9185 (N_9185,N_9025,N_9058);
xnor U9186 (N_9186,N_9096,N_9080);
or U9187 (N_9187,N_9123,N_9059);
and U9188 (N_9188,N_9076,N_9070);
xor U9189 (N_9189,N_9067,N_9096);
nand U9190 (N_9190,N_9000,N_9090);
and U9191 (N_9191,N_9054,N_9014);
xor U9192 (N_9192,N_9058,N_9071);
or U9193 (N_9193,N_9119,N_9043);
nand U9194 (N_9194,N_9062,N_9001);
nor U9195 (N_9195,N_9080,N_9071);
nand U9196 (N_9196,N_9044,N_9070);
and U9197 (N_9197,N_9087,N_9026);
nand U9198 (N_9198,N_9001,N_9109);
nand U9199 (N_9199,N_9070,N_9015);
and U9200 (N_9200,N_9012,N_9095);
and U9201 (N_9201,N_9019,N_9022);
nand U9202 (N_9202,N_9113,N_9104);
or U9203 (N_9203,N_9025,N_9087);
or U9204 (N_9204,N_9072,N_9024);
nor U9205 (N_9205,N_9123,N_9114);
and U9206 (N_9206,N_9018,N_9085);
or U9207 (N_9207,N_9087,N_9020);
xor U9208 (N_9208,N_9124,N_9087);
nor U9209 (N_9209,N_9023,N_9066);
or U9210 (N_9210,N_9117,N_9026);
nand U9211 (N_9211,N_9005,N_9088);
nand U9212 (N_9212,N_9096,N_9049);
nand U9213 (N_9213,N_9065,N_9050);
xor U9214 (N_9214,N_9040,N_9020);
xor U9215 (N_9215,N_9069,N_9067);
and U9216 (N_9216,N_9075,N_9104);
nand U9217 (N_9217,N_9015,N_9038);
or U9218 (N_9218,N_9040,N_9098);
and U9219 (N_9219,N_9103,N_9082);
nand U9220 (N_9220,N_9024,N_9094);
and U9221 (N_9221,N_9103,N_9010);
nand U9222 (N_9222,N_9088,N_9053);
nor U9223 (N_9223,N_9018,N_9080);
nor U9224 (N_9224,N_9038,N_9079);
or U9225 (N_9225,N_9025,N_9037);
and U9226 (N_9226,N_9029,N_9021);
nor U9227 (N_9227,N_9103,N_9083);
nor U9228 (N_9228,N_9059,N_9105);
xnor U9229 (N_9229,N_9009,N_9116);
nor U9230 (N_9230,N_9024,N_9018);
or U9231 (N_9231,N_9050,N_9043);
nor U9232 (N_9232,N_9081,N_9118);
and U9233 (N_9233,N_9029,N_9123);
and U9234 (N_9234,N_9070,N_9030);
nor U9235 (N_9235,N_9021,N_9112);
nor U9236 (N_9236,N_9007,N_9035);
or U9237 (N_9237,N_9061,N_9073);
or U9238 (N_9238,N_9038,N_9061);
nand U9239 (N_9239,N_9043,N_9031);
and U9240 (N_9240,N_9080,N_9059);
nor U9241 (N_9241,N_9070,N_9118);
xor U9242 (N_9242,N_9012,N_9116);
xnor U9243 (N_9243,N_9061,N_9111);
and U9244 (N_9244,N_9005,N_9015);
or U9245 (N_9245,N_9008,N_9025);
xor U9246 (N_9246,N_9027,N_9011);
xor U9247 (N_9247,N_9073,N_9081);
nand U9248 (N_9248,N_9045,N_9079);
xor U9249 (N_9249,N_9014,N_9083);
nand U9250 (N_9250,N_9219,N_9181);
nor U9251 (N_9251,N_9192,N_9220);
and U9252 (N_9252,N_9216,N_9193);
or U9253 (N_9253,N_9164,N_9187);
xnor U9254 (N_9254,N_9156,N_9130);
or U9255 (N_9255,N_9160,N_9234);
or U9256 (N_9256,N_9217,N_9168);
xor U9257 (N_9257,N_9236,N_9150);
xnor U9258 (N_9258,N_9157,N_9210);
nand U9259 (N_9259,N_9188,N_9245);
or U9260 (N_9260,N_9232,N_9136);
and U9261 (N_9261,N_9147,N_9227);
nand U9262 (N_9262,N_9151,N_9174);
and U9263 (N_9263,N_9247,N_9244);
and U9264 (N_9264,N_9185,N_9133);
and U9265 (N_9265,N_9145,N_9237);
xnor U9266 (N_9266,N_9129,N_9195);
or U9267 (N_9267,N_9177,N_9165);
nand U9268 (N_9268,N_9226,N_9198);
nand U9269 (N_9269,N_9146,N_9222);
xnor U9270 (N_9270,N_9186,N_9148);
or U9271 (N_9271,N_9200,N_9142);
nor U9272 (N_9272,N_9137,N_9138);
xor U9273 (N_9273,N_9240,N_9243);
nand U9274 (N_9274,N_9211,N_9125);
nand U9275 (N_9275,N_9149,N_9166);
or U9276 (N_9276,N_9159,N_9203);
nand U9277 (N_9277,N_9154,N_9158);
nand U9278 (N_9278,N_9246,N_9206);
or U9279 (N_9279,N_9249,N_9241);
xor U9280 (N_9280,N_9178,N_9205);
or U9281 (N_9281,N_9132,N_9171);
xor U9282 (N_9282,N_9152,N_9173);
nand U9283 (N_9283,N_9180,N_9127);
nand U9284 (N_9284,N_9134,N_9204);
or U9285 (N_9285,N_9162,N_9233);
nand U9286 (N_9286,N_9128,N_9170);
and U9287 (N_9287,N_9175,N_9163);
or U9288 (N_9288,N_9197,N_9229);
nand U9289 (N_9289,N_9135,N_9141);
nor U9290 (N_9290,N_9169,N_9196);
or U9291 (N_9291,N_9221,N_9207);
xor U9292 (N_9292,N_9126,N_9215);
or U9293 (N_9293,N_9223,N_9184);
or U9294 (N_9294,N_9248,N_9202);
and U9295 (N_9295,N_9161,N_9179);
nor U9296 (N_9296,N_9144,N_9201);
nor U9297 (N_9297,N_9213,N_9189);
nor U9298 (N_9298,N_9190,N_9191);
nor U9299 (N_9299,N_9224,N_9131);
and U9300 (N_9300,N_9155,N_9167);
or U9301 (N_9301,N_9194,N_9209);
and U9302 (N_9302,N_9238,N_9228);
nor U9303 (N_9303,N_9239,N_9176);
and U9304 (N_9304,N_9231,N_9183);
and U9305 (N_9305,N_9182,N_9208);
nor U9306 (N_9306,N_9212,N_9140);
nor U9307 (N_9307,N_9218,N_9230);
nor U9308 (N_9308,N_9153,N_9235);
nor U9309 (N_9309,N_9214,N_9242);
xnor U9310 (N_9310,N_9199,N_9225);
nand U9311 (N_9311,N_9139,N_9143);
xnor U9312 (N_9312,N_9172,N_9245);
xnor U9313 (N_9313,N_9178,N_9247);
nor U9314 (N_9314,N_9224,N_9214);
nor U9315 (N_9315,N_9135,N_9247);
xor U9316 (N_9316,N_9145,N_9238);
or U9317 (N_9317,N_9145,N_9155);
nand U9318 (N_9318,N_9191,N_9167);
nand U9319 (N_9319,N_9164,N_9150);
xnor U9320 (N_9320,N_9207,N_9247);
nand U9321 (N_9321,N_9204,N_9184);
or U9322 (N_9322,N_9154,N_9201);
nand U9323 (N_9323,N_9125,N_9206);
xor U9324 (N_9324,N_9196,N_9127);
nor U9325 (N_9325,N_9161,N_9216);
xnor U9326 (N_9326,N_9237,N_9225);
xnor U9327 (N_9327,N_9138,N_9139);
xnor U9328 (N_9328,N_9221,N_9187);
and U9329 (N_9329,N_9240,N_9209);
nand U9330 (N_9330,N_9225,N_9248);
or U9331 (N_9331,N_9163,N_9234);
or U9332 (N_9332,N_9208,N_9237);
or U9333 (N_9333,N_9233,N_9239);
or U9334 (N_9334,N_9186,N_9240);
nand U9335 (N_9335,N_9131,N_9178);
or U9336 (N_9336,N_9125,N_9236);
nor U9337 (N_9337,N_9166,N_9154);
xor U9338 (N_9338,N_9246,N_9230);
nand U9339 (N_9339,N_9183,N_9178);
nor U9340 (N_9340,N_9201,N_9165);
or U9341 (N_9341,N_9134,N_9156);
xor U9342 (N_9342,N_9138,N_9239);
and U9343 (N_9343,N_9145,N_9199);
nor U9344 (N_9344,N_9186,N_9163);
nor U9345 (N_9345,N_9246,N_9184);
nand U9346 (N_9346,N_9164,N_9241);
xnor U9347 (N_9347,N_9125,N_9201);
xor U9348 (N_9348,N_9190,N_9208);
and U9349 (N_9349,N_9230,N_9191);
or U9350 (N_9350,N_9197,N_9212);
or U9351 (N_9351,N_9176,N_9248);
nor U9352 (N_9352,N_9238,N_9136);
and U9353 (N_9353,N_9211,N_9132);
nor U9354 (N_9354,N_9215,N_9190);
nand U9355 (N_9355,N_9229,N_9181);
xnor U9356 (N_9356,N_9196,N_9192);
nand U9357 (N_9357,N_9208,N_9136);
xnor U9358 (N_9358,N_9134,N_9224);
or U9359 (N_9359,N_9136,N_9170);
nand U9360 (N_9360,N_9167,N_9215);
nor U9361 (N_9361,N_9185,N_9230);
and U9362 (N_9362,N_9210,N_9244);
nor U9363 (N_9363,N_9188,N_9159);
nand U9364 (N_9364,N_9132,N_9186);
and U9365 (N_9365,N_9198,N_9248);
xor U9366 (N_9366,N_9207,N_9196);
nand U9367 (N_9367,N_9140,N_9146);
nand U9368 (N_9368,N_9210,N_9164);
nand U9369 (N_9369,N_9151,N_9126);
or U9370 (N_9370,N_9126,N_9138);
xnor U9371 (N_9371,N_9217,N_9142);
or U9372 (N_9372,N_9155,N_9244);
and U9373 (N_9373,N_9227,N_9239);
nand U9374 (N_9374,N_9187,N_9141);
and U9375 (N_9375,N_9355,N_9268);
xnor U9376 (N_9376,N_9316,N_9318);
xnor U9377 (N_9377,N_9290,N_9307);
xnor U9378 (N_9378,N_9361,N_9280);
or U9379 (N_9379,N_9255,N_9374);
and U9380 (N_9380,N_9294,N_9363);
nor U9381 (N_9381,N_9257,N_9284);
xnor U9382 (N_9382,N_9253,N_9279);
xor U9383 (N_9383,N_9350,N_9304);
nor U9384 (N_9384,N_9315,N_9311);
nand U9385 (N_9385,N_9371,N_9260);
nand U9386 (N_9386,N_9299,N_9288);
or U9387 (N_9387,N_9306,N_9267);
xor U9388 (N_9388,N_9372,N_9254);
and U9389 (N_9389,N_9275,N_9333);
nor U9390 (N_9390,N_9259,N_9327);
nand U9391 (N_9391,N_9250,N_9302);
nand U9392 (N_9392,N_9310,N_9297);
nand U9393 (N_9393,N_9357,N_9330);
or U9394 (N_9394,N_9323,N_9359);
or U9395 (N_9395,N_9340,N_9272);
nor U9396 (N_9396,N_9348,N_9324);
and U9397 (N_9397,N_9341,N_9292);
nor U9398 (N_9398,N_9286,N_9370);
nand U9399 (N_9399,N_9252,N_9262);
and U9400 (N_9400,N_9256,N_9277);
nand U9401 (N_9401,N_9325,N_9271);
nand U9402 (N_9402,N_9308,N_9300);
nand U9403 (N_9403,N_9326,N_9356);
or U9404 (N_9404,N_9337,N_9344);
nand U9405 (N_9405,N_9328,N_9335);
and U9406 (N_9406,N_9332,N_9273);
xor U9407 (N_9407,N_9367,N_9261);
xnor U9408 (N_9408,N_9320,N_9338);
nor U9409 (N_9409,N_9276,N_9285);
or U9410 (N_9410,N_9281,N_9322);
xnor U9411 (N_9411,N_9289,N_9269);
and U9412 (N_9412,N_9369,N_9362);
or U9413 (N_9413,N_9274,N_9351);
or U9414 (N_9414,N_9305,N_9343);
or U9415 (N_9415,N_9321,N_9345);
nor U9416 (N_9416,N_9336,N_9301);
nand U9417 (N_9417,N_9296,N_9303);
nor U9418 (N_9418,N_9287,N_9331);
and U9419 (N_9419,N_9293,N_9282);
nor U9420 (N_9420,N_9373,N_9298);
and U9421 (N_9421,N_9295,N_9354);
or U9422 (N_9422,N_9329,N_9314);
nand U9423 (N_9423,N_9353,N_9365);
nand U9424 (N_9424,N_9352,N_9319);
or U9425 (N_9425,N_9266,N_9346);
and U9426 (N_9426,N_9334,N_9278);
or U9427 (N_9427,N_9317,N_9349);
xor U9428 (N_9428,N_9347,N_9339);
nor U9429 (N_9429,N_9364,N_9283);
nand U9430 (N_9430,N_9291,N_9264);
nor U9431 (N_9431,N_9309,N_9263);
and U9432 (N_9432,N_9270,N_9368);
nor U9433 (N_9433,N_9366,N_9358);
nor U9434 (N_9434,N_9313,N_9312);
or U9435 (N_9435,N_9251,N_9265);
nor U9436 (N_9436,N_9342,N_9360);
and U9437 (N_9437,N_9258,N_9277);
and U9438 (N_9438,N_9350,N_9310);
nand U9439 (N_9439,N_9350,N_9370);
and U9440 (N_9440,N_9346,N_9250);
xor U9441 (N_9441,N_9259,N_9331);
and U9442 (N_9442,N_9261,N_9302);
or U9443 (N_9443,N_9355,N_9287);
or U9444 (N_9444,N_9290,N_9316);
xor U9445 (N_9445,N_9322,N_9369);
and U9446 (N_9446,N_9373,N_9339);
and U9447 (N_9447,N_9332,N_9373);
nor U9448 (N_9448,N_9364,N_9281);
xnor U9449 (N_9449,N_9331,N_9260);
nand U9450 (N_9450,N_9275,N_9317);
nor U9451 (N_9451,N_9363,N_9310);
or U9452 (N_9452,N_9312,N_9338);
and U9453 (N_9453,N_9367,N_9267);
or U9454 (N_9454,N_9303,N_9334);
and U9455 (N_9455,N_9277,N_9288);
and U9456 (N_9456,N_9285,N_9261);
nand U9457 (N_9457,N_9302,N_9354);
nand U9458 (N_9458,N_9336,N_9344);
and U9459 (N_9459,N_9352,N_9338);
and U9460 (N_9460,N_9282,N_9332);
nor U9461 (N_9461,N_9361,N_9268);
nor U9462 (N_9462,N_9316,N_9257);
and U9463 (N_9463,N_9318,N_9261);
xnor U9464 (N_9464,N_9261,N_9284);
nand U9465 (N_9465,N_9348,N_9253);
xnor U9466 (N_9466,N_9370,N_9251);
nand U9467 (N_9467,N_9347,N_9351);
xnor U9468 (N_9468,N_9366,N_9313);
xnor U9469 (N_9469,N_9252,N_9345);
or U9470 (N_9470,N_9256,N_9273);
and U9471 (N_9471,N_9372,N_9266);
xor U9472 (N_9472,N_9369,N_9319);
and U9473 (N_9473,N_9344,N_9358);
and U9474 (N_9474,N_9277,N_9354);
xnor U9475 (N_9475,N_9362,N_9321);
nor U9476 (N_9476,N_9343,N_9292);
xnor U9477 (N_9477,N_9266,N_9369);
nand U9478 (N_9478,N_9349,N_9305);
xnor U9479 (N_9479,N_9355,N_9344);
nor U9480 (N_9480,N_9324,N_9300);
xor U9481 (N_9481,N_9318,N_9302);
and U9482 (N_9482,N_9362,N_9334);
xnor U9483 (N_9483,N_9348,N_9261);
nand U9484 (N_9484,N_9253,N_9290);
nor U9485 (N_9485,N_9306,N_9373);
or U9486 (N_9486,N_9324,N_9309);
nand U9487 (N_9487,N_9370,N_9358);
nand U9488 (N_9488,N_9261,N_9336);
and U9489 (N_9489,N_9314,N_9370);
nand U9490 (N_9490,N_9286,N_9368);
or U9491 (N_9491,N_9273,N_9303);
nand U9492 (N_9492,N_9277,N_9302);
nand U9493 (N_9493,N_9304,N_9347);
or U9494 (N_9494,N_9331,N_9364);
or U9495 (N_9495,N_9312,N_9276);
nor U9496 (N_9496,N_9357,N_9331);
nor U9497 (N_9497,N_9331,N_9322);
xor U9498 (N_9498,N_9296,N_9259);
and U9499 (N_9499,N_9348,N_9358);
nand U9500 (N_9500,N_9445,N_9497);
or U9501 (N_9501,N_9462,N_9381);
or U9502 (N_9502,N_9421,N_9392);
nand U9503 (N_9503,N_9436,N_9415);
nand U9504 (N_9504,N_9428,N_9480);
xor U9505 (N_9505,N_9396,N_9398);
xor U9506 (N_9506,N_9495,N_9444);
xnor U9507 (N_9507,N_9496,N_9401);
and U9508 (N_9508,N_9454,N_9399);
and U9509 (N_9509,N_9422,N_9426);
nor U9510 (N_9510,N_9489,N_9402);
xnor U9511 (N_9511,N_9490,N_9395);
nand U9512 (N_9512,N_9451,N_9457);
and U9513 (N_9513,N_9492,N_9471);
or U9514 (N_9514,N_9393,N_9382);
nor U9515 (N_9515,N_9408,N_9423);
and U9516 (N_9516,N_9377,N_9420);
or U9517 (N_9517,N_9453,N_9469);
or U9518 (N_9518,N_9390,N_9427);
nand U9519 (N_9519,N_9380,N_9447);
or U9520 (N_9520,N_9460,N_9413);
and U9521 (N_9521,N_9475,N_9476);
and U9522 (N_9522,N_9491,N_9403);
nor U9523 (N_9523,N_9433,N_9458);
nand U9524 (N_9524,N_9493,N_9431);
nand U9525 (N_9525,N_9483,N_9499);
nor U9526 (N_9526,N_9446,N_9441);
nor U9527 (N_9527,N_9459,N_9478);
nor U9528 (N_9528,N_9468,N_9411);
nor U9529 (N_9529,N_9467,N_9397);
nor U9530 (N_9530,N_9391,N_9388);
xor U9531 (N_9531,N_9494,N_9481);
and U9532 (N_9532,N_9455,N_9429);
nand U9533 (N_9533,N_9464,N_9410);
xor U9534 (N_9534,N_9498,N_9461);
xnor U9535 (N_9535,N_9409,N_9418);
and U9536 (N_9536,N_9473,N_9448);
nor U9537 (N_9537,N_9432,N_9407);
nand U9538 (N_9538,N_9470,N_9484);
xnor U9539 (N_9539,N_9442,N_9456);
and U9540 (N_9540,N_9387,N_9379);
or U9541 (N_9541,N_9463,N_9375);
and U9542 (N_9542,N_9383,N_9435);
and U9543 (N_9543,N_9440,N_9404);
nor U9544 (N_9544,N_9474,N_9376);
or U9545 (N_9545,N_9452,N_9472);
nor U9546 (N_9546,N_9419,N_9425);
and U9547 (N_9547,N_9389,N_9400);
and U9548 (N_9548,N_9405,N_9385);
or U9549 (N_9549,N_9479,N_9437);
nand U9550 (N_9550,N_9443,N_9394);
and U9551 (N_9551,N_9488,N_9414);
and U9552 (N_9552,N_9487,N_9417);
or U9553 (N_9553,N_9424,N_9450);
nor U9554 (N_9554,N_9386,N_9482);
nor U9555 (N_9555,N_9439,N_9449);
xor U9556 (N_9556,N_9485,N_9466);
and U9557 (N_9557,N_9378,N_9430);
xnor U9558 (N_9558,N_9416,N_9384);
nor U9559 (N_9559,N_9406,N_9465);
nand U9560 (N_9560,N_9486,N_9438);
nand U9561 (N_9561,N_9477,N_9434);
and U9562 (N_9562,N_9412,N_9397);
and U9563 (N_9563,N_9448,N_9406);
xor U9564 (N_9564,N_9460,N_9390);
and U9565 (N_9565,N_9482,N_9428);
or U9566 (N_9566,N_9494,N_9453);
nand U9567 (N_9567,N_9481,N_9403);
nor U9568 (N_9568,N_9475,N_9409);
or U9569 (N_9569,N_9476,N_9489);
xnor U9570 (N_9570,N_9449,N_9394);
nor U9571 (N_9571,N_9497,N_9478);
nand U9572 (N_9572,N_9419,N_9392);
or U9573 (N_9573,N_9472,N_9377);
or U9574 (N_9574,N_9386,N_9400);
nor U9575 (N_9575,N_9467,N_9463);
or U9576 (N_9576,N_9488,N_9481);
and U9577 (N_9577,N_9497,N_9385);
nor U9578 (N_9578,N_9379,N_9376);
xnor U9579 (N_9579,N_9382,N_9472);
and U9580 (N_9580,N_9401,N_9390);
nor U9581 (N_9581,N_9458,N_9472);
and U9582 (N_9582,N_9444,N_9456);
or U9583 (N_9583,N_9478,N_9415);
xor U9584 (N_9584,N_9419,N_9476);
or U9585 (N_9585,N_9499,N_9446);
or U9586 (N_9586,N_9487,N_9485);
nor U9587 (N_9587,N_9420,N_9411);
nand U9588 (N_9588,N_9496,N_9397);
nand U9589 (N_9589,N_9464,N_9419);
and U9590 (N_9590,N_9499,N_9403);
or U9591 (N_9591,N_9438,N_9472);
nand U9592 (N_9592,N_9457,N_9474);
nor U9593 (N_9593,N_9389,N_9397);
xnor U9594 (N_9594,N_9389,N_9385);
nand U9595 (N_9595,N_9496,N_9392);
nand U9596 (N_9596,N_9428,N_9388);
and U9597 (N_9597,N_9411,N_9497);
xnor U9598 (N_9598,N_9469,N_9376);
xnor U9599 (N_9599,N_9412,N_9468);
and U9600 (N_9600,N_9411,N_9427);
xor U9601 (N_9601,N_9410,N_9461);
nor U9602 (N_9602,N_9450,N_9485);
nor U9603 (N_9603,N_9420,N_9448);
xnor U9604 (N_9604,N_9487,N_9430);
and U9605 (N_9605,N_9375,N_9403);
or U9606 (N_9606,N_9440,N_9480);
xor U9607 (N_9607,N_9491,N_9482);
and U9608 (N_9608,N_9428,N_9483);
xnor U9609 (N_9609,N_9399,N_9464);
nor U9610 (N_9610,N_9423,N_9451);
and U9611 (N_9611,N_9400,N_9398);
xor U9612 (N_9612,N_9473,N_9431);
nor U9613 (N_9613,N_9435,N_9407);
or U9614 (N_9614,N_9494,N_9490);
or U9615 (N_9615,N_9453,N_9385);
or U9616 (N_9616,N_9474,N_9416);
xor U9617 (N_9617,N_9398,N_9393);
or U9618 (N_9618,N_9409,N_9441);
xor U9619 (N_9619,N_9381,N_9451);
nor U9620 (N_9620,N_9471,N_9438);
or U9621 (N_9621,N_9442,N_9446);
nand U9622 (N_9622,N_9499,N_9480);
nand U9623 (N_9623,N_9458,N_9395);
nor U9624 (N_9624,N_9380,N_9383);
or U9625 (N_9625,N_9500,N_9511);
or U9626 (N_9626,N_9604,N_9613);
nand U9627 (N_9627,N_9602,N_9546);
or U9628 (N_9628,N_9607,N_9502);
and U9629 (N_9629,N_9529,N_9547);
xnor U9630 (N_9630,N_9532,N_9519);
or U9631 (N_9631,N_9557,N_9622);
nand U9632 (N_9632,N_9563,N_9591);
nand U9633 (N_9633,N_9578,N_9612);
xnor U9634 (N_9634,N_9555,N_9538);
xnor U9635 (N_9635,N_9575,N_9520);
nor U9636 (N_9636,N_9553,N_9570);
nand U9637 (N_9637,N_9558,N_9611);
or U9638 (N_9638,N_9507,N_9624);
xnor U9639 (N_9639,N_9588,N_9550);
and U9640 (N_9640,N_9574,N_9534);
or U9641 (N_9641,N_9554,N_9504);
and U9642 (N_9642,N_9561,N_9527);
nand U9643 (N_9643,N_9597,N_9531);
or U9644 (N_9644,N_9526,N_9548);
nor U9645 (N_9645,N_9587,N_9608);
nor U9646 (N_9646,N_9543,N_9533);
and U9647 (N_9647,N_9586,N_9621);
nand U9648 (N_9648,N_9565,N_9521);
or U9649 (N_9649,N_9525,N_9559);
or U9650 (N_9650,N_9523,N_9589);
nand U9651 (N_9651,N_9584,N_9580);
nor U9652 (N_9652,N_9549,N_9616);
nand U9653 (N_9653,N_9556,N_9518);
nor U9654 (N_9654,N_9503,N_9596);
or U9655 (N_9655,N_9618,N_9540);
xor U9656 (N_9656,N_9517,N_9568);
nand U9657 (N_9657,N_9599,N_9620);
nand U9658 (N_9658,N_9590,N_9551);
nand U9659 (N_9659,N_9536,N_9542);
or U9660 (N_9660,N_9579,N_9583);
xor U9661 (N_9661,N_9585,N_9576);
and U9662 (N_9662,N_9567,N_9516);
nand U9663 (N_9663,N_9564,N_9506);
xnor U9664 (N_9664,N_9619,N_9566);
and U9665 (N_9665,N_9569,N_9512);
nor U9666 (N_9666,N_9539,N_9600);
nand U9667 (N_9667,N_9609,N_9508);
or U9668 (N_9668,N_9615,N_9617);
nor U9669 (N_9669,N_9514,N_9606);
or U9670 (N_9670,N_9535,N_9528);
or U9671 (N_9671,N_9515,N_9513);
xnor U9672 (N_9672,N_9501,N_9544);
and U9673 (N_9673,N_9560,N_9577);
nand U9674 (N_9674,N_9610,N_9530);
nor U9675 (N_9675,N_9605,N_9594);
nand U9676 (N_9676,N_9522,N_9545);
nor U9677 (N_9677,N_9509,N_9595);
or U9678 (N_9678,N_9541,N_9572);
and U9679 (N_9679,N_9601,N_9614);
nand U9680 (N_9680,N_9537,N_9603);
nand U9681 (N_9681,N_9581,N_9592);
nand U9682 (N_9682,N_9623,N_9582);
or U9683 (N_9683,N_9524,N_9562);
nand U9684 (N_9684,N_9571,N_9593);
nor U9685 (N_9685,N_9510,N_9505);
or U9686 (N_9686,N_9598,N_9552);
xor U9687 (N_9687,N_9573,N_9564);
nand U9688 (N_9688,N_9602,N_9551);
xor U9689 (N_9689,N_9574,N_9556);
nand U9690 (N_9690,N_9538,N_9585);
nand U9691 (N_9691,N_9536,N_9555);
and U9692 (N_9692,N_9535,N_9545);
or U9693 (N_9693,N_9551,N_9526);
xnor U9694 (N_9694,N_9619,N_9561);
and U9695 (N_9695,N_9538,N_9579);
nor U9696 (N_9696,N_9506,N_9550);
or U9697 (N_9697,N_9577,N_9589);
or U9698 (N_9698,N_9594,N_9577);
or U9699 (N_9699,N_9609,N_9591);
xor U9700 (N_9700,N_9562,N_9586);
nor U9701 (N_9701,N_9587,N_9546);
and U9702 (N_9702,N_9539,N_9552);
and U9703 (N_9703,N_9546,N_9599);
or U9704 (N_9704,N_9561,N_9577);
and U9705 (N_9705,N_9569,N_9530);
or U9706 (N_9706,N_9617,N_9533);
or U9707 (N_9707,N_9566,N_9528);
nand U9708 (N_9708,N_9543,N_9550);
nor U9709 (N_9709,N_9555,N_9534);
xnor U9710 (N_9710,N_9613,N_9558);
nand U9711 (N_9711,N_9518,N_9603);
xnor U9712 (N_9712,N_9535,N_9590);
xor U9713 (N_9713,N_9536,N_9623);
xor U9714 (N_9714,N_9545,N_9538);
nand U9715 (N_9715,N_9573,N_9609);
and U9716 (N_9716,N_9517,N_9582);
nand U9717 (N_9717,N_9579,N_9530);
and U9718 (N_9718,N_9571,N_9553);
xor U9719 (N_9719,N_9555,N_9575);
and U9720 (N_9720,N_9565,N_9537);
xor U9721 (N_9721,N_9617,N_9528);
and U9722 (N_9722,N_9549,N_9524);
nor U9723 (N_9723,N_9529,N_9563);
nand U9724 (N_9724,N_9614,N_9549);
or U9725 (N_9725,N_9558,N_9620);
xor U9726 (N_9726,N_9512,N_9592);
and U9727 (N_9727,N_9512,N_9555);
xnor U9728 (N_9728,N_9596,N_9533);
or U9729 (N_9729,N_9605,N_9617);
and U9730 (N_9730,N_9511,N_9554);
or U9731 (N_9731,N_9502,N_9610);
nor U9732 (N_9732,N_9531,N_9546);
xnor U9733 (N_9733,N_9548,N_9518);
nand U9734 (N_9734,N_9594,N_9549);
xor U9735 (N_9735,N_9611,N_9526);
nand U9736 (N_9736,N_9573,N_9611);
nor U9737 (N_9737,N_9523,N_9564);
nor U9738 (N_9738,N_9563,N_9611);
xnor U9739 (N_9739,N_9504,N_9609);
nand U9740 (N_9740,N_9512,N_9584);
and U9741 (N_9741,N_9599,N_9565);
nor U9742 (N_9742,N_9591,N_9570);
and U9743 (N_9743,N_9555,N_9598);
xor U9744 (N_9744,N_9503,N_9567);
nor U9745 (N_9745,N_9515,N_9530);
xor U9746 (N_9746,N_9615,N_9501);
xnor U9747 (N_9747,N_9532,N_9553);
xor U9748 (N_9748,N_9519,N_9603);
and U9749 (N_9749,N_9521,N_9604);
nor U9750 (N_9750,N_9659,N_9744);
nor U9751 (N_9751,N_9658,N_9674);
and U9752 (N_9752,N_9719,N_9687);
or U9753 (N_9753,N_9643,N_9640);
nand U9754 (N_9754,N_9668,N_9746);
nor U9755 (N_9755,N_9727,N_9696);
nor U9756 (N_9756,N_9691,N_9677);
nand U9757 (N_9757,N_9648,N_9655);
nor U9758 (N_9758,N_9637,N_9697);
nand U9759 (N_9759,N_9667,N_9704);
xor U9760 (N_9760,N_9701,N_9645);
nand U9761 (N_9761,N_9728,N_9625);
nor U9762 (N_9762,N_9663,N_9747);
or U9763 (N_9763,N_9725,N_9634);
or U9764 (N_9764,N_9694,N_9717);
nand U9765 (N_9765,N_9642,N_9683);
or U9766 (N_9766,N_9715,N_9630);
or U9767 (N_9767,N_9711,N_9678);
nor U9768 (N_9768,N_9628,N_9654);
nor U9769 (N_9769,N_9676,N_9735);
and U9770 (N_9770,N_9661,N_9722);
and U9771 (N_9771,N_9723,N_9749);
and U9772 (N_9772,N_9708,N_9656);
xnor U9773 (N_9773,N_9681,N_9660);
nand U9774 (N_9774,N_9695,N_9680);
nor U9775 (N_9775,N_9652,N_9703);
nand U9776 (N_9776,N_9626,N_9635);
nor U9777 (N_9777,N_9649,N_9627);
or U9778 (N_9778,N_9673,N_9650);
and U9779 (N_9779,N_9629,N_9631);
nor U9780 (N_9780,N_9718,N_9720);
nor U9781 (N_9781,N_9662,N_9716);
or U9782 (N_9782,N_9647,N_9726);
nand U9783 (N_9783,N_9707,N_9666);
nor U9784 (N_9784,N_9713,N_9679);
and U9785 (N_9785,N_9636,N_9734);
and U9786 (N_9786,N_9736,N_9669);
or U9787 (N_9787,N_9646,N_9633);
xor U9788 (N_9788,N_9644,N_9700);
and U9789 (N_9789,N_9732,N_9688);
or U9790 (N_9790,N_9748,N_9657);
or U9791 (N_9791,N_9664,N_9724);
nor U9792 (N_9792,N_9641,N_9682);
xor U9793 (N_9793,N_9743,N_9738);
and U9794 (N_9794,N_9686,N_9698);
nand U9795 (N_9795,N_9653,N_9737);
and U9796 (N_9796,N_9733,N_9731);
or U9797 (N_9797,N_9685,N_9702);
nor U9798 (N_9798,N_9742,N_9651);
and U9799 (N_9799,N_9670,N_9632);
and U9800 (N_9800,N_9714,N_9712);
xor U9801 (N_9801,N_9721,N_9665);
or U9802 (N_9802,N_9690,N_9699);
xor U9803 (N_9803,N_9672,N_9671);
nand U9804 (N_9804,N_9706,N_9739);
and U9805 (N_9805,N_9705,N_9638);
and U9806 (N_9806,N_9710,N_9675);
xor U9807 (N_9807,N_9692,N_9689);
xor U9808 (N_9808,N_9684,N_9741);
and U9809 (N_9809,N_9709,N_9639);
nand U9810 (N_9810,N_9740,N_9745);
nand U9811 (N_9811,N_9730,N_9729);
or U9812 (N_9812,N_9693,N_9718);
or U9813 (N_9813,N_9691,N_9728);
and U9814 (N_9814,N_9636,N_9647);
nor U9815 (N_9815,N_9722,N_9667);
and U9816 (N_9816,N_9639,N_9636);
nor U9817 (N_9817,N_9745,N_9739);
nor U9818 (N_9818,N_9660,N_9706);
xor U9819 (N_9819,N_9667,N_9730);
or U9820 (N_9820,N_9686,N_9730);
or U9821 (N_9821,N_9715,N_9666);
nand U9822 (N_9822,N_9707,N_9742);
and U9823 (N_9823,N_9705,N_9733);
xor U9824 (N_9824,N_9655,N_9713);
xnor U9825 (N_9825,N_9629,N_9658);
nand U9826 (N_9826,N_9728,N_9631);
or U9827 (N_9827,N_9718,N_9706);
and U9828 (N_9828,N_9652,N_9662);
nand U9829 (N_9829,N_9718,N_9660);
xnor U9830 (N_9830,N_9672,N_9686);
nand U9831 (N_9831,N_9689,N_9676);
nor U9832 (N_9832,N_9681,N_9706);
or U9833 (N_9833,N_9707,N_9710);
or U9834 (N_9834,N_9633,N_9719);
xnor U9835 (N_9835,N_9642,N_9732);
or U9836 (N_9836,N_9714,N_9667);
or U9837 (N_9837,N_9739,N_9730);
nor U9838 (N_9838,N_9737,N_9645);
nor U9839 (N_9839,N_9656,N_9637);
or U9840 (N_9840,N_9645,N_9666);
and U9841 (N_9841,N_9710,N_9656);
xor U9842 (N_9842,N_9670,N_9728);
nand U9843 (N_9843,N_9672,N_9703);
and U9844 (N_9844,N_9638,N_9702);
and U9845 (N_9845,N_9626,N_9715);
nand U9846 (N_9846,N_9731,N_9628);
nor U9847 (N_9847,N_9657,N_9734);
nand U9848 (N_9848,N_9625,N_9661);
and U9849 (N_9849,N_9699,N_9736);
and U9850 (N_9850,N_9669,N_9746);
xnor U9851 (N_9851,N_9706,N_9729);
nand U9852 (N_9852,N_9679,N_9636);
and U9853 (N_9853,N_9726,N_9677);
or U9854 (N_9854,N_9675,N_9692);
xnor U9855 (N_9855,N_9680,N_9658);
nor U9856 (N_9856,N_9747,N_9712);
and U9857 (N_9857,N_9738,N_9701);
or U9858 (N_9858,N_9702,N_9687);
and U9859 (N_9859,N_9703,N_9636);
and U9860 (N_9860,N_9635,N_9744);
and U9861 (N_9861,N_9732,N_9658);
nor U9862 (N_9862,N_9648,N_9682);
nand U9863 (N_9863,N_9713,N_9668);
nand U9864 (N_9864,N_9642,N_9694);
nor U9865 (N_9865,N_9636,N_9625);
xor U9866 (N_9866,N_9699,N_9692);
and U9867 (N_9867,N_9740,N_9708);
nand U9868 (N_9868,N_9678,N_9699);
and U9869 (N_9869,N_9672,N_9685);
and U9870 (N_9870,N_9633,N_9642);
nor U9871 (N_9871,N_9749,N_9633);
nor U9872 (N_9872,N_9689,N_9643);
xnor U9873 (N_9873,N_9690,N_9743);
xnor U9874 (N_9874,N_9700,N_9726);
xor U9875 (N_9875,N_9778,N_9869);
nor U9876 (N_9876,N_9800,N_9839);
nor U9877 (N_9877,N_9849,N_9847);
or U9878 (N_9878,N_9779,N_9809);
nand U9879 (N_9879,N_9850,N_9789);
nand U9880 (N_9880,N_9856,N_9807);
xnor U9881 (N_9881,N_9823,N_9765);
and U9882 (N_9882,N_9790,N_9803);
nand U9883 (N_9883,N_9845,N_9818);
or U9884 (N_9884,N_9859,N_9793);
nor U9885 (N_9885,N_9861,N_9771);
nor U9886 (N_9886,N_9851,N_9868);
nand U9887 (N_9887,N_9842,N_9768);
or U9888 (N_9888,N_9769,N_9794);
and U9889 (N_9889,N_9802,N_9792);
xnor U9890 (N_9890,N_9777,N_9812);
and U9891 (N_9891,N_9772,N_9864);
and U9892 (N_9892,N_9833,N_9784);
or U9893 (N_9893,N_9750,N_9820);
nand U9894 (N_9894,N_9834,N_9773);
and U9895 (N_9895,N_9835,N_9836);
xnor U9896 (N_9896,N_9806,N_9846);
nand U9897 (N_9897,N_9852,N_9811);
nand U9898 (N_9898,N_9873,N_9816);
nand U9899 (N_9899,N_9810,N_9813);
nor U9900 (N_9900,N_9756,N_9821);
and U9901 (N_9901,N_9841,N_9825);
xnor U9902 (N_9902,N_9840,N_9783);
and U9903 (N_9903,N_9843,N_9760);
or U9904 (N_9904,N_9801,N_9782);
and U9905 (N_9905,N_9791,N_9867);
nor U9906 (N_9906,N_9767,N_9826);
nor U9907 (N_9907,N_9755,N_9788);
or U9908 (N_9908,N_9831,N_9798);
nand U9909 (N_9909,N_9844,N_9838);
xor U9910 (N_9910,N_9837,N_9832);
nor U9911 (N_9911,N_9751,N_9795);
or U9912 (N_9912,N_9830,N_9866);
and U9913 (N_9913,N_9817,N_9787);
and U9914 (N_9914,N_9814,N_9785);
xor U9915 (N_9915,N_9815,N_9862);
and U9916 (N_9916,N_9829,N_9805);
or U9917 (N_9917,N_9797,N_9774);
nand U9918 (N_9918,N_9808,N_9824);
nand U9919 (N_9919,N_9799,N_9754);
or U9920 (N_9920,N_9871,N_9764);
nand U9921 (N_9921,N_9781,N_9858);
nor U9922 (N_9922,N_9855,N_9759);
nor U9923 (N_9923,N_9770,N_9762);
or U9924 (N_9924,N_9848,N_9872);
nor U9925 (N_9925,N_9757,N_9874);
or U9926 (N_9926,N_9780,N_9853);
xnor U9927 (N_9927,N_9865,N_9857);
nor U9928 (N_9928,N_9786,N_9863);
xnor U9929 (N_9929,N_9776,N_9763);
xnor U9930 (N_9930,N_9827,N_9753);
nor U9931 (N_9931,N_9804,N_9822);
nand U9932 (N_9932,N_9870,N_9761);
nor U9933 (N_9933,N_9752,N_9854);
xor U9934 (N_9934,N_9819,N_9775);
nand U9935 (N_9935,N_9766,N_9758);
xor U9936 (N_9936,N_9796,N_9860);
and U9937 (N_9937,N_9828,N_9820);
xor U9938 (N_9938,N_9816,N_9751);
xnor U9939 (N_9939,N_9848,N_9754);
nor U9940 (N_9940,N_9777,N_9786);
xnor U9941 (N_9941,N_9866,N_9859);
or U9942 (N_9942,N_9765,N_9768);
and U9943 (N_9943,N_9767,N_9865);
or U9944 (N_9944,N_9768,N_9816);
nor U9945 (N_9945,N_9804,N_9823);
and U9946 (N_9946,N_9871,N_9815);
xor U9947 (N_9947,N_9857,N_9830);
or U9948 (N_9948,N_9762,N_9852);
and U9949 (N_9949,N_9824,N_9855);
or U9950 (N_9950,N_9849,N_9804);
xnor U9951 (N_9951,N_9776,N_9864);
nand U9952 (N_9952,N_9855,N_9752);
or U9953 (N_9953,N_9809,N_9769);
nand U9954 (N_9954,N_9807,N_9752);
xnor U9955 (N_9955,N_9785,N_9777);
nor U9956 (N_9956,N_9802,N_9861);
xor U9957 (N_9957,N_9818,N_9831);
or U9958 (N_9958,N_9768,N_9802);
nand U9959 (N_9959,N_9873,N_9797);
nand U9960 (N_9960,N_9852,N_9797);
nand U9961 (N_9961,N_9822,N_9819);
nand U9962 (N_9962,N_9835,N_9851);
or U9963 (N_9963,N_9760,N_9820);
and U9964 (N_9964,N_9833,N_9780);
xor U9965 (N_9965,N_9856,N_9813);
xnor U9966 (N_9966,N_9769,N_9806);
nand U9967 (N_9967,N_9837,N_9838);
xnor U9968 (N_9968,N_9866,N_9831);
xor U9969 (N_9969,N_9823,N_9754);
xnor U9970 (N_9970,N_9819,N_9762);
nand U9971 (N_9971,N_9868,N_9859);
and U9972 (N_9972,N_9754,N_9750);
and U9973 (N_9973,N_9836,N_9863);
nor U9974 (N_9974,N_9769,N_9762);
or U9975 (N_9975,N_9757,N_9861);
or U9976 (N_9976,N_9757,N_9863);
nor U9977 (N_9977,N_9846,N_9817);
or U9978 (N_9978,N_9771,N_9836);
or U9979 (N_9979,N_9850,N_9762);
and U9980 (N_9980,N_9758,N_9774);
nor U9981 (N_9981,N_9834,N_9802);
and U9982 (N_9982,N_9776,N_9791);
or U9983 (N_9983,N_9811,N_9780);
and U9984 (N_9984,N_9835,N_9824);
xor U9985 (N_9985,N_9831,N_9770);
nor U9986 (N_9986,N_9851,N_9874);
xor U9987 (N_9987,N_9755,N_9825);
xor U9988 (N_9988,N_9815,N_9762);
nand U9989 (N_9989,N_9800,N_9836);
xor U9990 (N_9990,N_9801,N_9831);
xor U9991 (N_9991,N_9862,N_9816);
and U9992 (N_9992,N_9869,N_9802);
and U9993 (N_9993,N_9833,N_9851);
or U9994 (N_9994,N_9832,N_9865);
and U9995 (N_9995,N_9813,N_9818);
or U9996 (N_9996,N_9760,N_9765);
nor U9997 (N_9997,N_9760,N_9874);
xnor U9998 (N_9998,N_9756,N_9855);
and U9999 (N_9999,N_9787,N_9774);
xnor U10000 (N_10000,N_9931,N_9954);
nor U10001 (N_10001,N_9902,N_9979);
or U10002 (N_10002,N_9891,N_9896);
or U10003 (N_10003,N_9926,N_9962);
xnor U10004 (N_10004,N_9924,N_9980);
nor U10005 (N_10005,N_9916,N_9903);
nor U10006 (N_10006,N_9997,N_9978);
xor U10007 (N_10007,N_9950,N_9906);
and U10008 (N_10008,N_9967,N_9934);
or U10009 (N_10009,N_9933,N_9918);
nor U10010 (N_10010,N_9969,N_9942);
xnor U10011 (N_10011,N_9955,N_9911);
or U10012 (N_10012,N_9999,N_9889);
nand U10013 (N_10013,N_9876,N_9944);
and U10014 (N_10014,N_9881,N_9991);
and U10015 (N_10015,N_9935,N_9887);
and U10016 (N_10016,N_9905,N_9880);
and U10017 (N_10017,N_9912,N_9973);
or U10018 (N_10018,N_9992,N_9956);
and U10019 (N_10019,N_9976,N_9977);
nand U10020 (N_10020,N_9983,N_9927);
xnor U10021 (N_10021,N_9938,N_9958);
nor U10022 (N_10022,N_9882,N_9909);
nand U10023 (N_10023,N_9972,N_9930);
nor U10024 (N_10024,N_9932,N_9945);
and U10025 (N_10025,N_9937,N_9928);
xnor U10026 (N_10026,N_9960,N_9915);
xnor U10027 (N_10027,N_9975,N_9922);
xor U10028 (N_10028,N_9957,N_9949);
and U10029 (N_10029,N_9987,N_9895);
xnor U10030 (N_10030,N_9943,N_9948);
xor U10031 (N_10031,N_9974,N_9994);
nand U10032 (N_10032,N_9947,N_9951);
nor U10033 (N_10033,N_9885,N_9961);
or U10034 (N_10034,N_9995,N_9920);
xor U10035 (N_10035,N_9941,N_9883);
or U10036 (N_10036,N_9907,N_9996);
nand U10037 (N_10037,N_9879,N_9963);
xor U10038 (N_10038,N_9898,N_9959);
and U10039 (N_10039,N_9913,N_9910);
or U10040 (N_10040,N_9984,N_9993);
and U10041 (N_10041,N_9929,N_9964);
or U10042 (N_10042,N_9894,N_9990);
nor U10043 (N_10043,N_9982,N_9886);
xnor U10044 (N_10044,N_9875,N_9940);
or U10045 (N_10045,N_9893,N_9919);
nor U10046 (N_10046,N_9908,N_9914);
or U10047 (N_10047,N_9970,N_9900);
and U10048 (N_10048,N_9877,N_9888);
and U10049 (N_10049,N_9890,N_9936);
and U10050 (N_10050,N_9946,N_9925);
or U10051 (N_10051,N_9923,N_9985);
xor U10052 (N_10052,N_9897,N_9981);
and U10053 (N_10053,N_9884,N_9952);
or U10054 (N_10054,N_9971,N_9989);
xor U10055 (N_10055,N_9988,N_9917);
xor U10056 (N_10056,N_9892,N_9968);
xor U10057 (N_10057,N_9998,N_9953);
nand U10058 (N_10058,N_9899,N_9965);
nand U10059 (N_10059,N_9986,N_9904);
and U10060 (N_10060,N_9901,N_9966);
nor U10061 (N_10061,N_9939,N_9921);
xor U10062 (N_10062,N_9878,N_9992);
nand U10063 (N_10063,N_9892,N_9917);
or U10064 (N_10064,N_9971,N_9929);
nor U10065 (N_10065,N_9886,N_9964);
or U10066 (N_10066,N_9915,N_9930);
and U10067 (N_10067,N_9916,N_9906);
nand U10068 (N_10068,N_9996,N_9959);
and U10069 (N_10069,N_9989,N_9943);
xnor U10070 (N_10070,N_9897,N_9928);
nand U10071 (N_10071,N_9991,N_9950);
nor U10072 (N_10072,N_9942,N_9922);
xor U10073 (N_10073,N_9904,N_9921);
nand U10074 (N_10074,N_9997,N_9982);
nand U10075 (N_10075,N_9975,N_9934);
or U10076 (N_10076,N_9912,N_9949);
or U10077 (N_10077,N_9977,N_9988);
and U10078 (N_10078,N_9927,N_9949);
or U10079 (N_10079,N_9900,N_9984);
or U10080 (N_10080,N_9953,N_9900);
nand U10081 (N_10081,N_9992,N_9923);
nand U10082 (N_10082,N_9983,N_9878);
and U10083 (N_10083,N_9898,N_9937);
or U10084 (N_10084,N_9958,N_9939);
nand U10085 (N_10085,N_9948,N_9935);
xor U10086 (N_10086,N_9968,N_9998);
and U10087 (N_10087,N_9928,N_9998);
nand U10088 (N_10088,N_9949,N_9925);
nor U10089 (N_10089,N_9920,N_9906);
and U10090 (N_10090,N_9916,N_9929);
nor U10091 (N_10091,N_9909,N_9924);
or U10092 (N_10092,N_9969,N_9917);
nor U10093 (N_10093,N_9942,N_9879);
nor U10094 (N_10094,N_9901,N_9980);
or U10095 (N_10095,N_9987,N_9877);
nor U10096 (N_10096,N_9985,N_9974);
nand U10097 (N_10097,N_9992,N_9943);
nor U10098 (N_10098,N_9929,N_9943);
nand U10099 (N_10099,N_9996,N_9994);
nor U10100 (N_10100,N_9933,N_9926);
nand U10101 (N_10101,N_9876,N_9957);
xnor U10102 (N_10102,N_9954,N_9944);
or U10103 (N_10103,N_9989,N_9913);
nor U10104 (N_10104,N_9889,N_9922);
xor U10105 (N_10105,N_9992,N_9985);
nor U10106 (N_10106,N_9946,N_9928);
nor U10107 (N_10107,N_9918,N_9998);
and U10108 (N_10108,N_9952,N_9897);
nand U10109 (N_10109,N_9905,N_9910);
and U10110 (N_10110,N_9939,N_9879);
xnor U10111 (N_10111,N_9904,N_9930);
xor U10112 (N_10112,N_9933,N_9950);
nand U10113 (N_10113,N_9942,N_9900);
nor U10114 (N_10114,N_9893,N_9933);
nand U10115 (N_10115,N_9932,N_9993);
or U10116 (N_10116,N_9904,N_9911);
and U10117 (N_10117,N_9963,N_9997);
and U10118 (N_10118,N_9982,N_9961);
and U10119 (N_10119,N_9927,N_9918);
xnor U10120 (N_10120,N_9951,N_9964);
xnor U10121 (N_10121,N_9992,N_9959);
nand U10122 (N_10122,N_9891,N_9904);
xor U10123 (N_10123,N_9939,N_9894);
nand U10124 (N_10124,N_9981,N_9890);
nor U10125 (N_10125,N_10040,N_10083);
or U10126 (N_10126,N_10092,N_10084);
and U10127 (N_10127,N_10060,N_10070);
or U10128 (N_10128,N_10096,N_10042);
nor U10129 (N_10129,N_10036,N_10080);
nand U10130 (N_10130,N_10121,N_10056);
nand U10131 (N_10131,N_10038,N_10091);
nor U10132 (N_10132,N_10016,N_10035);
and U10133 (N_10133,N_10044,N_10032);
nor U10134 (N_10134,N_10100,N_10020);
or U10135 (N_10135,N_10079,N_10082);
nor U10136 (N_10136,N_10022,N_10025);
nand U10137 (N_10137,N_10002,N_10113);
or U10138 (N_10138,N_10021,N_10034);
nand U10139 (N_10139,N_10088,N_10041);
or U10140 (N_10140,N_10006,N_10061);
nand U10141 (N_10141,N_10017,N_10112);
nor U10142 (N_10142,N_10059,N_10069);
or U10143 (N_10143,N_10120,N_10124);
nand U10144 (N_10144,N_10028,N_10005);
nand U10145 (N_10145,N_10026,N_10118);
or U10146 (N_10146,N_10086,N_10107);
nand U10147 (N_10147,N_10076,N_10018);
and U10148 (N_10148,N_10010,N_10058);
and U10149 (N_10149,N_10001,N_10119);
or U10150 (N_10150,N_10098,N_10050);
and U10151 (N_10151,N_10049,N_10055);
nor U10152 (N_10152,N_10053,N_10000);
xor U10153 (N_10153,N_10093,N_10057);
nand U10154 (N_10154,N_10064,N_10008);
or U10155 (N_10155,N_10115,N_10014);
or U10156 (N_10156,N_10071,N_10110);
nand U10157 (N_10157,N_10030,N_10052);
nor U10158 (N_10158,N_10104,N_10012);
xor U10159 (N_10159,N_10033,N_10037);
xnor U10160 (N_10160,N_10085,N_10045);
xor U10161 (N_10161,N_10101,N_10072);
or U10162 (N_10162,N_10024,N_10013);
nand U10163 (N_10163,N_10095,N_10102);
or U10164 (N_10164,N_10090,N_10074);
nor U10165 (N_10165,N_10078,N_10027);
nand U10166 (N_10166,N_10073,N_10063);
nand U10167 (N_10167,N_10015,N_10051);
and U10168 (N_10168,N_10007,N_10117);
and U10169 (N_10169,N_10094,N_10106);
and U10170 (N_10170,N_10105,N_10048);
xnor U10171 (N_10171,N_10111,N_10068);
xnor U10172 (N_10172,N_10081,N_10023);
and U10173 (N_10173,N_10109,N_10062);
nor U10174 (N_10174,N_10054,N_10066);
nor U10175 (N_10175,N_10031,N_10047);
nor U10176 (N_10176,N_10019,N_10089);
and U10177 (N_10177,N_10067,N_10039);
or U10178 (N_10178,N_10108,N_10087);
nor U10179 (N_10179,N_10075,N_10116);
or U10180 (N_10180,N_10123,N_10114);
or U10181 (N_10181,N_10003,N_10099);
or U10182 (N_10182,N_10029,N_10011);
and U10183 (N_10183,N_10009,N_10077);
nor U10184 (N_10184,N_10097,N_10103);
or U10185 (N_10185,N_10122,N_10046);
nor U10186 (N_10186,N_10043,N_10004);
nor U10187 (N_10187,N_10065,N_10021);
or U10188 (N_10188,N_10037,N_10124);
nor U10189 (N_10189,N_10005,N_10118);
xnor U10190 (N_10190,N_10012,N_10024);
xor U10191 (N_10191,N_10026,N_10042);
and U10192 (N_10192,N_10042,N_10088);
nor U10193 (N_10193,N_10036,N_10005);
and U10194 (N_10194,N_10070,N_10062);
nand U10195 (N_10195,N_10047,N_10019);
xnor U10196 (N_10196,N_10030,N_10085);
xnor U10197 (N_10197,N_10018,N_10048);
nand U10198 (N_10198,N_10018,N_10115);
xor U10199 (N_10199,N_10014,N_10119);
xnor U10200 (N_10200,N_10029,N_10018);
xnor U10201 (N_10201,N_10120,N_10077);
nand U10202 (N_10202,N_10072,N_10112);
nor U10203 (N_10203,N_10013,N_10006);
nand U10204 (N_10204,N_10009,N_10037);
nor U10205 (N_10205,N_10032,N_10081);
or U10206 (N_10206,N_10009,N_10087);
nand U10207 (N_10207,N_10045,N_10044);
nor U10208 (N_10208,N_10069,N_10041);
nor U10209 (N_10209,N_10118,N_10059);
and U10210 (N_10210,N_10028,N_10000);
nand U10211 (N_10211,N_10068,N_10037);
and U10212 (N_10212,N_10096,N_10016);
nand U10213 (N_10213,N_10062,N_10106);
nor U10214 (N_10214,N_10103,N_10021);
or U10215 (N_10215,N_10059,N_10033);
nor U10216 (N_10216,N_10118,N_10047);
or U10217 (N_10217,N_10051,N_10104);
nand U10218 (N_10218,N_10115,N_10020);
nor U10219 (N_10219,N_10089,N_10091);
and U10220 (N_10220,N_10118,N_10074);
nor U10221 (N_10221,N_10043,N_10024);
or U10222 (N_10222,N_10106,N_10111);
xor U10223 (N_10223,N_10078,N_10040);
nor U10224 (N_10224,N_10116,N_10002);
nor U10225 (N_10225,N_10057,N_10109);
or U10226 (N_10226,N_10110,N_10056);
nor U10227 (N_10227,N_10078,N_10011);
nand U10228 (N_10228,N_10100,N_10073);
or U10229 (N_10229,N_10066,N_10015);
nand U10230 (N_10230,N_10022,N_10031);
or U10231 (N_10231,N_10051,N_10044);
xor U10232 (N_10232,N_10026,N_10115);
and U10233 (N_10233,N_10093,N_10120);
nor U10234 (N_10234,N_10069,N_10105);
nand U10235 (N_10235,N_10012,N_10089);
nor U10236 (N_10236,N_10059,N_10019);
nand U10237 (N_10237,N_10103,N_10082);
nor U10238 (N_10238,N_10030,N_10113);
or U10239 (N_10239,N_10124,N_10097);
nor U10240 (N_10240,N_10102,N_10032);
xnor U10241 (N_10241,N_10002,N_10044);
or U10242 (N_10242,N_10018,N_10007);
or U10243 (N_10243,N_10039,N_10012);
and U10244 (N_10244,N_10102,N_10034);
and U10245 (N_10245,N_10022,N_10095);
or U10246 (N_10246,N_10035,N_10115);
nor U10247 (N_10247,N_10082,N_10029);
or U10248 (N_10248,N_10069,N_10013);
or U10249 (N_10249,N_10095,N_10014);
nor U10250 (N_10250,N_10173,N_10180);
xnor U10251 (N_10251,N_10147,N_10139);
xnor U10252 (N_10252,N_10135,N_10216);
nor U10253 (N_10253,N_10241,N_10148);
xnor U10254 (N_10254,N_10245,N_10141);
and U10255 (N_10255,N_10214,N_10240);
nand U10256 (N_10256,N_10227,N_10158);
or U10257 (N_10257,N_10221,N_10249);
nor U10258 (N_10258,N_10143,N_10166);
xnor U10259 (N_10259,N_10235,N_10204);
or U10260 (N_10260,N_10194,N_10188);
nor U10261 (N_10261,N_10239,N_10223);
and U10262 (N_10262,N_10243,N_10185);
xor U10263 (N_10263,N_10154,N_10172);
or U10264 (N_10264,N_10137,N_10209);
nand U10265 (N_10265,N_10233,N_10232);
and U10266 (N_10266,N_10131,N_10190);
xnor U10267 (N_10267,N_10238,N_10201);
nor U10268 (N_10268,N_10242,N_10231);
xor U10269 (N_10269,N_10133,N_10163);
nand U10270 (N_10270,N_10217,N_10196);
or U10271 (N_10271,N_10181,N_10162);
nand U10272 (N_10272,N_10174,N_10213);
and U10273 (N_10273,N_10234,N_10220);
nor U10274 (N_10274,N_10145,N_10189);
xnor U10275 (N_10275,N_10205,N_10237);
or U10276 (N_10276,N_10192,N_10126);
nand U10277 (N_10277,N_10156,N_10164);
nand U10278 (N_10278,N_10210,N_10224);
nand U10279 (N_10279,N_10222,N_10215);
xor U10280 (N_10280,N_10130,N_10179);
or U10281 (N_10281,N_10208,N_10229);
nor U10282 (N_10282,N_10230,N_10197);
or U10283 (N_10283,N_10128,N_10127);
or U10284 (N_10284,N_10177,N_10155);
nand U10285 (N_10285,N_10142,N_10198);
nand U10286 (N_10286,N_10211,N_10152);
xnor U10287 (N_10287,N_10178,N_10183);
and U10288 (N_10288,N_10218,N_10169);
nand U10289 (N_10289,N_10132,N_10207);
nand U10290 (N_10290,N_10200,N_10193);
nand U10291 (N_10291,N_10182,N_10184);
and U10292 (N_10292,N_10244,N_10125);
and U10293 (N_10293,N_10160,N_10203);
or U10294 (N_10294,N_10136,N_10170);
xnor U10295 (N_10295,N_10134,N_10171);
nor U10296 (N_10296,N_10236,N_10161);
and U10297 (N_10297,N_10144,N_10168);
xnor U10298 (N_10298,N_10195,N_10138);
or U10299 (N_10299,N_10206,N_10165);
nand U10300 (N_10300,N_10226,N_10167);
or U10301 (N_10301,N_10176,N_10212);
nand U10302 (N_10302,N_10199,N_10159);
or U10303 (N_10303,N_10187,N_10153);
nand U10304 (N_10304,N_10149,N_10247);
nand U10305 (N_10305,N_10129,N_10248);
or U10306 (N_10306,N_10175,N_10228);
nand U10307 (N_10307,N_10202,N_10151);
nor U10308 (N_10308,N_10191,N_10146);
xnor U10309 (N_10309,N_10246,N_10157);
nand U10310 (N_10310,N_10140,N_10150);
nand U10311 (N_10311,N_10186,N_10225);
or U10312 (N_10312,N_10219,N_10190);
xnor U10313 (N_10313,N_10195,N_10241);
or U10314 (N_10314,N_10226,N_10228);
xor U10315 (N_10315,N_10222,N_10129);
or U10316 (N_10316,N_10214,N_10143);
xnor U10317 (N_10317,N_10160,N_10182);
or U10318 (N_10318,N_10155,N_10157);
or U10319 (N_10319,N_10177,N_10231);
and U10320 (N_10320,N_10129,N_10243);
and U10321 (N_10321,N_10227,N_10230);
or U10322 (N_10322,N_10206,N_10248);
nor U10323 (N_10323,N_10202,N_10163);
nor U10324 (N_10324,N_10129,N_10245);
and U10325 (N_10325,N_10240,N_10175);
nand U10326 (N_10326,N_10163,N_10232);
xor U10327 (N_10327,N_10194,N_10189);
nand U10328 (N_10328,N_10150,N_10237);
and U10329 (N_10329,N_10230,N_10175);
nand U10330 (N_10330,N_10155,N_10201);
xnor U10331 (N_10331,N_10202,N_10175);
xnor U10332 (N_10332,N_10141,N_10167);
and U10333 (N_10333,N_10127,N_10149);
or U10334 (N_10334,N_10187,N_10172);
nor U10335 (N_10335,N_10127,N_10202);
nor U10336 (N_10336,N_10190,N_10222);
nand U10337 (N_10337,N_10233,N_10222);
or U10338 (N_10338,N_10143,N_10148);
nor U10339 (N_10339,N_10171,N_10131);
nor U10340 (N_10340,N_10210,N_10204);
and U10341 (N_10341,N_10176,N_10172);
and U10342 (N_10342,N_10194,N_10148);
nand U10343 (N_10343,N_10126,N_10145);
xor U10344 (N_10344,N_10220,N_10216);
or U10345 (N_10345,N_10198,N_10216);
and U10346 (N_10346,N_10166,N_10154);
xnor U10347 (N_10347,N_10207,N_10223);
nand U10348 (N_10348,N_10175,N_10245);
nor U10349 (N_10349,N_10128,N_10160);
nor U10350 (N_10350,N_10192,N_10219);
nand U10351 (N_10351,N_10230,N_10143);
xor U10352 (N_10352,N_10203,N_10134);
xor U10353 (N_10353,N_10188,N_10176);
nor U10354 (N_10354,N_10241,N_10208);
and U10355 (N_10355,N_10221,N_10151);
nor U10356 (N_10356,N_10215,N_10146);
nor U10357 (N_10357,N_10238,N_10240);
xor U10358 (N_10358,N_10225,N_10218);
and U10359 (N_10359,N_10241,N_10128);
xor U10360 (N_10360,N_10247,N_10204);
and U10361 (N_10361,N_10137,N_10131);
xor U10362 (N_10362,N_10190,N_10194);
xnor U10363 (N_10363,N_10128,N_10171);
xnor U10364 (N_10364,N_10228,N_10171);
or U10365 (N_10365,N_10171,N_10199);
nor U10366 (N_10366,N_10206,N_10146);
nor U10367 (N_10367,N_10242,N_10180);
and U10368 (N_10368,N_10206,N_10179);
nand U10369 (N_10369,N_10143,N_10127);
nor U10370 (N_10370,N_10179,N_10211);
or U10371 (N_10371,N_10207,N_10198);
or U10372 (N_10372,N_10204,N_10201);
and U10373 (N_10373,N_10188,N_10127);
or U10374 (N_10374,N_10152,N_10172);
and U10375 (N_10375,N_10314,N_10263);
or U10376 (N_10376,N_10300,N_10364);
or U10377 (N_10377,N_10341,N_10354);
nand U10378 (N_10378,N_10260,N_10264);
nand U10379 (N_10379,N_10332,N_10326);
xnor U10380 (N_10380,N_10367,N_10339);
nand U10381 (N_10381,N_10271,N_10255);
nor U10382 (N_10382,N_10350,N_10338);
xnor U10383 (N_10383,N_10250,N_10374);
xnor U10384 (N_10384,N_10252,N_10340);
nor U10385 (N_10385,N_10315,N_10286);
or U10386 (N_10386,N_10336,N_10369);
nand U10387 (N_10387,N_10353,N_10360);
nand U10388 (N_10388,N_10371,N_10328);
or U10389 (N_10389,N_10358,N_10345);
or U10390 (N_10390,N_10362,N_10329);
nand U10391 (N_10391,N_10295,N_10261);
nor U10392 (N_10392,N_10357,N_10293);
or U10393 (N_10393,N_10279,N_10302);
or U10394 (N_10394,N_10283,N_10292);
nor U10395 (N_10395,N_10331,N_10299);
and U10396 (N_10396,N_10301,N_10370);
nand U10397 (N_10397,N_10285,N_10270);
and U10398 (N_10398,N_10257,N_10304);
and U10399 (N_10399,N_10344,N_10323);
xor U10400 (N_10400,N_10267,N_10346);
nand U10401 (N_10401,N_10309,N_10324);
or U10402 (N_10402,N_10278,N_10359);
or U10403 (N_10403,N_10281,N_10305);
nand U10404 (N_10404,N_10361,N_10320);
or U10405 (N_10405,N_10327,N_10254);
xor U10406 (N_10406,N_10363,N_10296);
or U10407 (N_10407,N_10337,N_10266);
xor U10408 (N_10408,N_10280,N_10335);
xor U10409 (N_10409,N_10258,N_10274);
nand U10410 (N_10410,N_10262,N_10298);
and U10411 (N_10411,N_10318,N_10275);
nand U10412 (N_10412,N_10330,N_10325);
nor U10413 (N_10413,N_10288,N_10321);
or U10414 (N_10414,N_10256,N_10308);
or U10415 (N_10415,N_10287,N_10273);
or U10416 (N_10416,N_10269,N_10277);
nand U10417 (N_10417,N_10322,N_10290);
and U10418 (N_10418,N_10303,N_10265);
nand U10419 (N_10419,N_10365,N_10333);
nand U10420 (N_10420,N_10373,N_10312);
nor U10421 (N_10421,N_10343,N_10282);
or U10422 (N_10422,N_10313,N_10276);
nor U10423 (N_10423,N_10356,N_10355);
nand U10424 (N_10424,N_10351,N_10366);
xnor U10425 (N_10425,N_10259,N_10294);
nor U10426 (N_10426,N_10307,N_10348);
nand U10427 (N_10427,N_10347,N_10284);
and U10428 (N_10428,N_10251,N_10253);
or U10429 (N_10429,N_10349,N_10297);
xnor U10430 (N_10430,N_10352,N_10289);
or U10431 (N_10431,N_10268,N_10306);
nand U10432 (N_10432,N_10310,N_10319);
or U10433 (N_10433,N_10334,N_10342);
or U10434 (N_10434,N_10317,N_10316);
nor U10435 (N_10435,N_10372,N_10368);
nor U10436 (N_10436,N_10272,N_10311);
or U10437 (N_10437,N_10291,N_10369);
nand U10438 (N_10438,N_10367,N_10321);
or U10439 (N_10439,N_10295,N_10314);
and U10440 (N_10440,N_10323,N_10267);
or U10441 (N_10441,N_10311,N_10295);
nand U10442 (N_10442,N_10354,N_10358);
nor U10443 (N_10443,N_10358,N_10261);
and U10444 (N_10444,N_10257,N_10368);
nand U10445 (N_10445,N_10260,N_10327);
xor U10446 (N_10446,N_10298,N_10277);
or U10447 (N_10447,N_10342,N_10268);
or U10448 (N_10448,N_10372,N_10260);
nand U10449 (N_10449,N_10331,N_10323);
nand U10450 (N_10450,N_10253,N_10318);
xor U10451 (N_10451,N_10332,N_10313);
and U10452 (N_10452,N_10311,N_10252);
or U10453 (N_10453,N_10274,N_10364);
and U10454 (N_10454,N_10332,N_10352);
or U10455 (N_10455,N_10255,N_10280);
nand U10456 (N_10456,N_10374,N_10260);
and U10457 (N_10457,N_10307,N_10365);
or U10458 (N_10458,N_10373,N_10256);
nor U10459 (N_10459,N_10304,N_10285);
nand U10460 (N_10460,N_10288,N_10374);
nand U10461 (N_10461,N_10316,N_10270);
or U10462 (N_10462,N_10252,N_10302);
nand U10463 (N_10463,N_10259,N_10257);
and U10464 (N_10464,N_10326,N_10374);
and U10465 (N_10465,N_10366,N_10364);
nand U10466 (N_10466,N_10342,N_10317);
and U10467 (N_10467,N_10327,N_10270);
or U10468 (N_10468,N_10300,N_10328);
nand U10469 (N_10469,N_10362,N_10259);
nand U10470 (N_10470,N_10328,N_10320);
xnor U10471 (N_10471,N_10257,N_10270);
xnor U10472 (N_10472,N_10263,N_10374);
or U10473 (N_10473,N_10340,N_10342);
and U10474 (N_10474,N_10264,N_10316);
xor U10475 (N_10475,N_10328,N_10297);
and U10476 (N_10476,N_10284,N_10372);
xor U10477 (N_10477,N_10274,N_10260);
and U10478 (N_10478,N_10366,N_10327);
xnor U10479 (N_10479,N_10317,N_10332);
xor U10480 (N_10480,N_10251,N_10272);
nor U10481 (N_10481,N_10297,N_10361);
xor U10482 (N_10482,N_10293,N_10373);
or U10483 (N_10483,N_10251,N_10277);
nand U10484 (N_10484,N_10363,N_10355);
xnor U10485 (N_10485,N_10338,N_10301);
or U10486 (N_10486,N_10257,N_10342);
nor U10487 (N_10487,N_10352,N_10312);
nor U10488 (N_10488,N_10320,N_10265);
nand U10489 (N_10489,N_10258,N_10317);
or U10490 (N_10490,N_10370,N_10283);
or U10491 (N_10491,N_10263,N_10287);
or U10492 (N_10492,N_10349,N_10270);
nand U10493 (N_10493,N_10348,N_10273);
and U10494 (N_10494,N_10354,N_10261);
nor U10495 (N_10495,N_10267,N_10334);
or U10496 (N_10496,N_10250,N_10315);
and U10497 (N_10497,N_10277,N_10309);
or U10498 (N_10498,N_10326,N_10368);
or U10499 (N_10499,N_10359,N_10306);
nand U10500 (N_10500,N_10493,N_10464);
or U10501 (N_10501,N_10391,N_10404);
nor U10502 (N_10502,N_10443,N_10417);
xnor U10503 (N_10503,N_10422,N_10480);
nand U10504 (N_10504,N_10385,N_10474);
nand U10505 (N_10505,N_10459,N_10497);
nand U10506 (N_10506,N_10454,N_10402);
and U10507 (N_10507,N_10495,N_10467);
nand U10508 (N_10508,N_10390,N_10438);
or U10509 (N_10509,N_10442,N_10416);
nand U10510 (N_10510,N_10396,N_10484);
nor U10511 (N_10511,N_10431,N_10476);
or U10512 (N_10512,N_10457,N_10434);
and U10513 (N_10513,N_10486,N_10469);
nand U10514 (N_10514,N_10489,N_10405);
nand U10515 (N_10515,N_10428,N_10392);
xor U10516 (N_10516,N_10458,N_10420);
nand U10517 (N_10517,N_10407,N_10432);
and U10518 (N_10518,N_10447,N_10379);
xor U10519 (N_10519,N_10389,N_10410);
nor U10520 (N_10520,N_10406,N_10452);
or U10521 (N_10521,N_10483,N_10475);
nor U10522 (N_10522,N_10424,N_10487);
or U10523 (N_10523,N_10426,N_10460);
xnor U10524 (N_10524,N_10393,N_10477);
or U10525 (N_10525,N_10440,N_10425);
xor U10526 (N_10526,N_10470,N_10384);
or U10527 (N_10527,N_10492,N_10398);
nand U10528 (N_10528,N_10387,N_10473);
or U10529 (N_10529,N_10419,N_10479);
nor U10530 (N_10530,N_10449,N_10439);
xor U10531 (N_10531,N_10435,N_10453);
nor U10532 (N_10532,N_10498,N_10378);
xor U10533 (N_10533,N_10490,N_10383);
xor U10534 (N_10534,N_10375,N_10418);
or U10535 (N_10535,N_10403,N_10494);
xor U10536 (N_10536,N_10394,N_10450);
nand U10537 (N_10537,N_10496,N_10478);
or U10538 (N_10538,N_10412,N_10433);
nand U10539 (N_10539,N_10485,N_10499);
and U10540 (N_10540,N_10421,N_10451);
and U10541 (N_10541,N_10488,N_10430);
xnor U10542 (N_10542,N_10414,N_10461);
nor U10543 (N_10543,N_10446,N_10411);
nand U10544 (N_10544,N_10399,N_10377);
and U10545 (N_10545,N_10444,N_10397);
nand U10546 (N_10546,N_10481,N_10400);
nor U10547 (N_10547,N_10466,N_10427);
and U10548 (N_10548,N_10382,N_10380);
xor U10549 (N_10549,N_10376,N_10441);
nand U10550 (N_10550,N_10462,N_10436);
nor U10551 (N_10551,N_10408,N_10471);
nand U10552 (N_10552,N_10437,N_10401);
nor U10553 (N_10553,N_10482,N_10465);
nor U10554 (N_10554,N_10448,N_10388);
xor U10555 (N_10555,N_10456,N_10381);
nor U10556 (N_10556,N_10472,N_10423);
xor U10557 (N_10557,N_10455,N_10468);
and U10558 (N_10558,N_10395,N_10415);
nand U10559 (N_10559,N_10445,N_10491);
nand U10560 (N_10560,N_10386,N_10413);
and U10561 (N_10561,N_10429,N_10409);
nor U10562 (N_10562,N_10463,N_10413);
and U10563 (N_10563,N_10447,N_10451);
nand U10564 (N_10564,N_10485,N_10433);
and U10565 (N_10565,N_10404,N_10460);
nand U10566 (N_10566,N_10444,N_10489);
nand U10567 (N_10567,N_10387,N_10446);
xnor U10568 (N_10568,N_10460,N_10390);
nor U10569 (N_10569,N_10405,N_10410);
nand U10570 (N_10570,N_10385,N_10499);
xnor U10571 (N_10571,N_10389,N_10377);
nor U10572 (N_10572,N_10464,N_10439);
xor U10573 (N_10573,N_10475,N_10385);
xnor U10574 (N_10574,N_10486,N_10388);
xor U10575 (N_10575,N_10406,N_10495);
or U10576 (N_10576,N_10428,N_10494);
nor U10577 (N_10577,N_10449,N_10436);
and U10578 (N_10578,N_10397,N_10440);
xor U10579 (N_10579,N_10424,N_10391);
nor U10580 (N_10580,N_10378,N_10464);
nand U10581 (N_10581,N_10418,N_10416);
nor U10582 (N_10582,N_10434,N_10381);
and U10583 (N_10583,N_10448,N_10384);
and U10584 (N_10584,N_10400,N_10430);
nand U10585 (N_10585,N_10396,N_10405);
nor U10586 (N_10586,N_10451,N_10453);
nor U10587 (N_10587,N_10402,N_10472);
xor U10588 (N_10588,N_10402,N_10468);
nand U10589 (N_10589,N_10450,N_10461);
nand U10590 (N_10590,N_10457,N_10378);
nand U10591 (N_10591,N_10423,N_10437);
nand U10592 (N_10592,N_10487,N_10467);
nand U10593 (N_10593,N_10404,N_10456);
or U10594 (N_10594,N_10475,N_10488);
nand U10595 (N_10595,N_10432,N_10408);
xnor U10596 (N_10596,N_10455,N_10453);
nand U10597 (N_10597,N_10498,N_10384);
and U10598 (N_10598,N_10409,N_10453);
or U10599 (N_10599,N_10491,N_10423);
and U10600 (N_10600,N_10390,N_10457);
and U10601 (N_10601,N_10453,N_10394);
or U10602 (N_10602,N_10393,N_10442);
and U10603 (N_10603,N_10376,N_10459);
nand U10604 (N_10604,N_10454,N_10395);
or U10605 (N_10605,N_10403,N_10448);
xnor U10606 (N_10606,N_10425,N_10412);
or U10607 (N_10607,N_10390,N_10477);
and U10608 (N_10608,N_10472,N_10395);
xnor U10609 (N_10609,N_10458,N_10478);
xor U10610 (N_10610,N_10448,N_10473);
or U10611 (N_10611,N_10495,N_10393);
xnor U10612 (N_10612,N_10437,N_10458);
xor U10613 (N_10613,N_10412,N_10447);
and U10614 (N_10614,N_10433,N_10479);
nand U10615 (N_10615,N_10494,N_10479);
or U10616 (N_10616,N_10474,N_10449);
nand U10617 (N_10617,N_10430,N_10468);
and U10618 (N_10618,N_10426,N_10471);
or U10619 (N_10619,N_10397,N_10384);
nor U10620 (N_10620,N_10401,N_10441);
and U10621 (N_10621,N_10494,N_10455);
nor U10622 (N_10622,N_10411,N_10434);
xor U10623 (N_10623,N_10436,N_10441);
and U10624 (N_10624,N_10448,N_10393);
nand U10625 (N_10625,N_10610,N_10560);
xnor U10626 (N_10626,N_10623,N_10596);
nand U10627 (N_10627,N_10508,N_10563);
and U10628 (N_10628,N_10602,N_10509);
or U10629 (N_10629,N_10561,N_10525);
nand U10630 (N_10630,N_10526,N_10583);
xor U10631 (N_10631,N_10512,N_10550);
nor U10632 (N_10632,N_10511,N_10555);
nand U10633 (N_10633,N_10578,N_10553);
xor U10634 (N_10634,N_10516,N_10503);
nand U10635 (N_10635,N_10570,N_10517);
and U10636 (N_10636,N_10539,N_10557);
nand U10637 (N_10637,N_10533,N_10510);
xnor U10638 (N_10638,N_10500,N_10567);
nand U10639 (N_10639,N_10600,N_10599);
or U10640 (N_10640,N_10554,N_10615);
xnor U10641 (N_10641,N_10513,N_10609);
and U10642 (N_10642,N_10579,N_10588);
nor U10643 (N_10643,N_10617,N_10594);
or U10644 (N_10644,N_10576,N_10520);
xnor U10645 (N_10645,N_10537,N_10522);
nand U10646 (N_10646,N_10584,N_10587);
xnor U10647 (N_10647,N_10548,N_10564);
xor U10648 (N_10648,N_10612,N_10603);
or U10649 (N_10649,N_10566,N_10532);
or U10650 (N_10650,N_10558,N_10574);
or U10651 (N_10651,N_10565,N_10589);
or U10652 (N_10652,N_10524,N_10595);
and U10653 (N_10653,N_10575,N_10620);
xnor U10654 (N_10654,N_10544,N_10569);
and U10655 (N_10655,N_10568,N_10530);
xor U10656 (N_10656,N_10573,N_10536);
nor U10657 (N_10657,N_10541,N_10556);
and U10658 (N_10658,N_10586,N_10506);
xor U10659 (N_10659,N_10505,N_10504);
nor U10660 (N_10660,N_10552,N_10580);
xor U10661 (N_10661,N_10519,N_10590);
and U10662 (N_10662,N_10604,N_10540);
nor U10663 (N_10663,N_10507,N_10622);
xnor U10664 (N_10664,N_10614,N_10597);
or U10665 (N_10665,N_10582,N_10585);
nand U10666 (N_10666,N_10502,N_10601);
xnor U10667 (N_10667,N_10514,N_10559);
xnor U10668 (N_10668,N_10535,N_10598);
nand U10669 (N_10669,N_10605,N_10593);
and U10670 (N_10670,N_10608,N_10542);
nand U10671 (N_10671,N_10591,N_10529);
and U10672 (N_10672,N_10523,N_10518);
and U10673 (N_10673,N_10624,N_10562);
or U10674 (N_10674,N_10581,N_10549);
or U10675 (N_10675,N_10592,N_10619);
nand U10676 (N_10676,N_10543,N_10528);
nor U10677 (N_10677,N_10545,N_10606);
or U10678 (N_10678,N_10571,N_10611);
nand U10679 (N_10679,N_10621,N_10613);
nor U10680 (N_10680,N_10527,N_10531);
nand U10681 (N_10681,N_10577,N_10534);
and U10682 (N_10682,N_10521,N_10616);
and U10683 (N_10683,N_10607,N_10538);
or U10684 (N_10684,N_10547,N_10618);
and U10685 (N_10685,N_10572,N_10546);
nand U10686 (N_10686,N_10515,N_10501);
nand U10687 (N_10687,N_10551,N_10504);
nor U10688 (N_10688,N_10587,N_10545);
or U10689 (N_10689,N_10617,N_10574);
nand U10690 (N_10690,N_10601,N_10550);
nand U10691 (N_10691,N_10530,N_10541);
nor U10692 (N_10692,N_10501,N_10555);
or U10693 (N_10693,N_10525,N_10564);
nand U10694 (N_10694,N_10544,N_10505);
nor U10695 (N_10695,N_10554,N_10558);
and U10696 (N_10696,N_10535,N_10532);
and U10697 (N_10697,N_10515,N_10509);
nand U10698 (N_10698,N_10518,N_10539);
nand U10699 (N_10699,N_10611,N_10516);
nor U10700 (N_10700,N_10522,N_10591);
or U10701 (N_10701,N_10621,N_10582);
nor U10702 (N_10702,N_10523,N_10566);
or U10703 (N_10703,N_10503,N_10533);
nand U10704 (N_10704,N_10558,N_10591);
nand U10705 (N_10705,N_10588,N_10587);
xnor U10706 (N_10706,N_10561,N_10616);
and U10707 (N_10707,N_10530,N_10521);
and U10708 (N_10708,N_10567,N_10524);
and U10709 (N_10709,N_10555,N_10559);
nor U10710 (N_10710,N_10529,N_10525);
and U10711 (N_10711,N_10514,N_10506);
nor U10712 (N_10712,N_10559,N_10566);
or U10713 (N_10713,N_10621,N_10508);
xor U10714 (N_10714,N_10575,N_10565);
nand U10715 (N_10715,N_10536,N_10599);
xnor U10716 (N_10716,N_10587,N_10532);
xor U10717 (N_10717,N_10593,N_10586);
or U10718 (N_10718,N_10581,N_10558);
or U10719 (N_10719,N_10610,N_10559);
or U10720 (N_10720,N_10535,N_10550);
or U10721 (N_10721,N_10606,N_10557);
or U10722 (N_10722,N_10549,N_10602);
or U10723 (N_10723,N_10530,N_10582);
or U10724 (N_10724,N_10543,N_10522);
nand U10725 (N_10725,N_10608,N_10516);
or U10726 (N_10726,N_10529,N_10575);
and U10727 (N_10727,N_10580,N_10585);
and U10728 (N_10728,N_10584,N_10596);
and U10729 (N_10729,N_10541,N_10584);
or U10730 (N_10730,N_10504,N_10576);
nor U10731 (N_10731,N_10529,N_10535);
xnor U10732 (N_10732,N_10560,N_10623);
or U10733 (N_10733,N_10536,N_10575);
nor U10734 (N_10734,N_10621,N_10521);
xor U10735 (N_10735,N_10606,N_10541);
nand U10736 (N_10736,N_10516,N_10600);
and U10737 (N_10737,N_10550,N_10537);
nand U10738 (N_10738,N_10595,N_10555);
nand U10739 (N_10739,N_10562,N_10507);
xnor U10740 (N_10740,N_10546,N_10524);
nand U10741 (N_10741,N_10591,N_10537);
nand U10742 (N_10742,N_10521,N_10509);
nand U10743 (N_10743,N_10544,N_10508);
nand U10744 (N_10744,N_10523,N_10525);
and U10745 (N_10745,N_10557,N_10578);
and U10746 (N_10746,N_10554,N_10533);
nor U10747 (N_10747,N_10501,N_10525);
nor U10748 (N_10748,N_10567,N_10504);
nand U10749 (N_10749,N_10604,N_10579);
nor U10750 (N_10750,N_10732,N_10669);
xnor U10751 (N_10751,N_10718,N_10641);
nor U10752 (N_10752,N_10722,N_10746);
nand U10753 (N_10753,N_10738,N_10630);
or U10754 (N_10754,N_10687,N_10657);
nand U10755 (N_10755,N_10675,N_10729);
or U10756 (N_10756,N_10717,N_10723);
nand U10757 (N_10757,N_10714,N_10685);
nor U10758 (N_10758,N_10631,N_10653);
xnor U10759 (N_10759,N_10670,N_10627);
and U10760 (N_10760,N_10740,N_10634);
and U10761 (N_10761,N_10743,N_10699);
nor U10762 (N_10762,N_10749,N_10643);
xnor U10763 (N_10763,N_10705,N_10642);
nand U10764 (N_10764,N_10688,N_10659);
nand U10765 (N_10765,N_10737,N_10721);
xnor U10766 (N_10766,N_10745,N_10635);
xnor U10767 (N_10767,N_10628,N_10692);
and U10768 (N_10768,N_10695,N_10734);
nand U10769 (N_10769,N_10702,N_10678);
xor U10770 (N_10770,N_10681,N_10629);
xnor U10771 (N_10771,N_10638,N_10704);
xor U10772 (N_10772,N_10713,N_10671);
or U10773 (N_10773,N_10694,N_10683);
nor U10774 (N_10774,N_10667,N_10654);
and U10775 (N_10775,N_10662,N_10645);
or U10776 (N_10776,N_10733,N_10655);
nand U10777 (N_10777,N_10739,N_10710);
nor U10778 (N_10778,N_10700,N_10697);
or U10779 (N_10779,N_10680,N_10625);
xor U10780 (N_10780,N_10663,N_10696);
xor U10781 (N_10781,N_10682,N_10731);
nand U10782 (N_10782,N_10646,N_10665);
nand U10783 (N_10783,N_10715,N_10652);
nor U10784 (N_10784,N_10689,N_10686);
and U10785 (N_10785,N_10649,N_10742);
or U10786 (N_10786,N_10719,N_10632);
nor U10787 (N_10787,N_10650,N_10724);
xor U10788 (N_10788,N_10708,N_10673);
or U10789 (N_10789,N_10661,N_10691);
xor U10790 (N_10790,N_10648,N_10636);
nand U10791 (N_10791,N_10706,N_10651);
xor U10792 (N_10792,N_10698,N_10660);
or U10793 (N_10793,N_10677,N_10703);
nand U10794 (N_10794,N_10720,N_10716);
and U10795 (N_10795,N_10728,N_10640);
and U10796 (N_10796,N_10672,N_10747);
or U10797 (N_10797,N_10709,N_10727);
xor U10798 (N_10798,N_10712,N_10730);
xor U10799 (N_10799,N_10626,N_10725);
nor U10800 (N_10800,N_10644,N_10637);
or U10801 (N_10801,N_10748,N_10684);
xnor U10802 (N_10802,N_10701,N_10741);
nor U10803 (N_10803,N_10726,N_10633);
and U10804 (N_10804,N_10707,N_10668);
nand U10805 (N_10805,N_10656,N_10676);
nand U10806 (N_10806,N_10679,N_10711);
nand U10807 (N_10807,N_10674,N_10647);
nor U10808 (N_10808,N_10664,N_10735);
nand U10809 (N_10809,N_10690,N_10693);
and U10810 (N_10810,N_10736,N_10658);
or U10811 (N_10811,N_10666,N_10744);
xor U10812 (N_10812,N_10639,N_10747);
and U10813 (N_10813,N_10724,N_10705);
xnor U10814 (N_10814,N_10626,N_10683);
nor U10815 (N_10815,N_10731,N_10707);
nand U10816 (N_10816,N_10659,N_10744);
nor U10817 (N_10817,N_10726,N_10690);
nand U10818 (N_10818,N_10746,N_10714);
and U10819 (N_10819,N_10654,N_10740);
or U10820 (N_10820,N_10724,N_10743);
xor U10821 (N_10821,N_10675,N_10663);
or U10822 (N_10822,N_10713,N_10748);
nand U10823 (N_10823,N_10709,N_10631);
and U10824 (N_10824,N_10684,N_10724);
nand U10825 (N_10825,N_10662,N_10739);
xnor U10826 (N_10826,N_10679,N_10714);
or U10827 (N_10827,N_10728,N_10704);
nand U10828 (N_10828,N_10741,N_10634);
and U10829 (N_10829,N_10702,N_10642);
nor U10830 (N_10830,N_10644,N_10693);
nor U10831 (N_10831,N_10695,N_10689);
and U10832 (N_10832,N_10746,N_10692);
xor U10833 (N_10833,N_10654,N_10707);
nor U10834 (N_10834,N_10689,N_10728);
or U10835 (N_10835,N_10718,N_10646);
xnor U10836 (N_10836,N_10626,N_10733);
xor U10837 (N_10837,N_10737,N_10722);
or U10838 (N_10838,N_10738,N_10676);
xnor U10839 (N_10839,N_10700,N_10651);
nand U10840 (N_10840,N_10747,N_10677);
xor U10841 (N_10841,N_10722,N_10632);
nand U10842 (N_10842,N_10729,N_10657);
nand U10843 (N_10843,N_10698,N_10711);
nand U10844 (N_10844,N_10626,N_10654);
xnor U10845 (N_10845,N_10743,N_10632);
nor U10846 (N_10846,N_10673,N_10677);
nand U10847 (N_10847,N_10633,N_10657);
xnor U10848 (N_10848,N_10671,N_10695);
nor U10849 (N_10849,N_10694,N_10646);
and U10850 (N_10850,N_10643,N_10625);
and U10851 (N_10851,N_10665,N_10714);
or U10852 (N_10852,N_10722,N_10721);
or U10853 (N_10853,N_10704,N_10745);
nor U10854 (N_10854,N_10708,N_10691);
nor U10855 (N_10855,N_10683,N_10646);
or U10856 (N_10856,N_10725,N_10682);
or U10857 (N_10857,N_10690,N_10698);
xor U10858 (N_10858,N_10666,N_10702);
xor U10859 (N_10859,N_10701,N_10710);
nor U10860 (N_10860,N_10684,N_10730);
xor U10861 (N_10861,N_10681,N_10703);
nor U10862 (N_10862,N_10668,N_10719);
nor U10863 (N_10863,N_10703,N_10628);
nand U10864 (N_10864,N_10708,N_10715);
xnor U10865 (N_10865,N_10642,N_10703);
or U10866 (N_10866,N_10696,N_10637);
and U10867 (N_10867,N_10640,N_10628);
and U10868 (N_10868,N_10728,N_10698);
nand U10869 (N_10869,N_10689,N_10680);
or U10870 (N_10870,N_10660,N_10638);
xnor U10871 (N_10871,N_10704,N_10631);
and U10872 (N_10872,N_10711,N_10651);
and U10873 (N_10873,N_10746,N_10716);
or U10874 (N_10874,N_10737,N_10704);
or U10875 (N_10875,N_10791,N_10844);
or U10876 (N_10876,N_10807,N_10826);
and U10877 (N_10877,N_10871,N_10783);
nand U10878 (N_10878,N_10780,N_10828);
or U10879 (N_10879,N_10757,N_10766);
nor U10880 (N_10880,N_10767,N_10794);
nor U10881 (N_10881,N_10778,N_10869);
and U10882 (N_10882,N_10792,N_10761);
or U10883 (N_10883,N_10795,N_10831);
or U10884 (N_10884,N_10867,N_10755);
xnor U10885 (N_10885,N_10835,N_10864);
nand U10886 (N_10886,N_10827,N_10808);
or U10887 (N_10887,N_10858,N_10769);
nand U10888 (N_10888,N_10809,N_10830);
and U10889 (N_10889,N_10756,N_10845);
xnor U10890 (N_10890,N_10825,N_10852);
xor U10891 (N_10891,N_10870,N_10764);
or U10892 (N_10892,N_10861,N_10829);
and U10893 (N_10893,N_10823,N_10788);
nor U10894 (N_10894,N_10874,N_10855);
xor U10895 (N_10895,N_10799,N_10853);
nor U10896 (N_10896,N_10873,N_10754);
nand U10897 (N_10897,N_10866,N_10805);
nand U10898 (N_10898,N_10860,N_10787);
and U10899 (N_10899,N_10840,N_10782);
or U10900 (N_10900,N_10772,N_10859);
and U10901 (N_10901,N_10850,N_10802);
and U10902 (N_10902,N_10848,N_10773);
and U10903 (N_10903,N_10762,N_10753);
xor U10904 (N_10904,N_10774,N_10810);
or U10905 (N_10905,N_10834,N_10775);
xor U10906 (N_10906,N_10833,N_10847);
and U10907 (N_10907,N_10843,N_10770);
xnor U10908 (N_10908,N_10818,N_10846);
or U10909 (N_10909,N_10832,N_10765);
or U10910 (N_10910,N_10781,N_10816);
nand U10911 (N_10911,N_10813,N_10763);
nor U10912 (N_10912,N_10814,N_10842);
xor U10913 (N_10913,N_10856,N_10758);
nand U10914 (N_10914,N_10820,N_10872);
and U10915 (N_10915,N_10798,N_10821);
nor U10916 (N_10916,N_10849,N_10812);
nor U10917 (N_10917,N_10790,N_10854);
nand U10918 (N_10918,N_10785,N_10751);
xnor U10919 (N_10919,N_10759,N_10803);
or U10920 (N_10920,N_10804,N_10811);
or U10921 (N_10921,N_10796,N_10865);
and U10922 (N_10922,N_10771,N_10760);
and U10923 (N_10923,N_10824,N_10837);
nand U10924 (N_10924,N_10779,N_10793);
xnor U10925 (N_10925,N_10863,N_10750);
nand U10926 (N_10926,N_10836,N_10801);
xnor U10927 (N_10927,N_10822,N_10776);
nor U10928 (N_10928,N_10857,N_10868);
and U10929 (N_10929,N_10817,N_10806);
nor U10930 (N_10930,N_10851,N_10784);
nand U10931 (N_10931,N_10841,N_10768);
nand U10932 (N_10932,N_10815,N_10752);
and U10933 (N_10933,N_10838,N_10862);
and U10934 (N_10934,N_10797,N_10839);
and U10935 (N_10935,N_10786,N_10819);
and U10936 (N_10936,N_10777,N_10789);
and U10937 (N_10937,N_10800,N_10779);
nand U10938 (N_10938,N_10753,N_10798);
nand U10939 (N_10939,N_10804,N_10796);
and U10940 (N_10940,N_10814,N_10788);
or U10941 (N_10941,N_10781,N_10768);
nor U10942 (N_10942,N_10812,N_10753);
or U10943 (N_10943,N_10784,N_10832);
nand U10944 (N_10944,N_10871,N_10807);
or U10945 (N_10945,N_10773,N_10787);
xor U10946 (N_10946,N_10808,N_10810);
or U10947 (N_10947,N_10805,N_10868);
xnor U10948 (N_10948,N_10778,N_10834);
nor U10949 (N_10949,N_10821,N_10804);
nand U10950 (N_10950,N_10834,N_10793);
nand U10951 (N_10951,N_10785,N_10807);
nand U10952 (N_10952,N_10779,N_10811);
and U10953 (N_10953,N_10825,N_10771);
or U10954 (N_10954,N_10782,N_10791);
nor U10955 (N_10955,N_10865,N_10772);
nand U10956 (N_10956,N_10821,N_10842);
and U10957 (N_10957,N_10874,N_10854);
or U10958 (N_10958,N_10863,N_10844);
and U10959 (N_10959,N_10845,N_10821);
xor U10960 (N_10960,N_10840,N_10809);
xor U10961 (N_10961,N_10777,N_10830);
nand U10962 (N_10962,N_10846,N_10835);
nor U10963 (N_10963,N_10803,N_10843);
and U10964 (N_10964,N_10752,N_10763);
nor U10965 (N_10965,N_10823,N_10872);
or U10966 (N_10966,N_10838,N_10800);
nor U10967 (N_10967,N_10762,N_10827);
xnor U10968 (N_10968,N_10830,N_10769);
and U10969 (N_10969,N_10842,N_10832);
xor U10970 (N_10970,N_10855,N_10815);
and U10971 (N_10971,N_10798,N_10808);
xnor U10972 (N_10972,N_10813,N_10846);
or U10973 (N_10973,N_10782,N_10752);
nor U10974 (N_10974,N_10828,N_10816);
and U10975 (N_10975,N_10830,N_10780);
nor U10976 (N_10976,N_10805,N_10763);
nand U10977 (N_10977,N_10817,N_10848);
nor U10978 (N_10978,N_10812,N_10869);
nand U10979 (N_10979,N_10798,N_10835);
or U10980 (N_10980,N_10837,N_10803);
or U10981 (N_10981,N_10757,N_10767);
or U10982 (N_10982,N_10854,N_10813);
nor U10983 (N_10983,N_10863,N_10852);
nor U10984 (N_10984,N_10832,N_10864);
and U10985 (N_10985,N_10872,N_10819);
xor U10986 (N_10986,N_10834,N_10871);
and U10987 (N_10987,N_10793,N_10837);
or U10988 (N_10988,N_10863,N_10781);
nor U10989 (N_10989,N_10794,N_10798);
nand U10990 (N_10990,N_10821,N_10766);
nand U10991 (N_10991,N_10847,N_10812);
or U10992 (N_10992,N_10838,N_10819);
nor U10993 (N_10993,N_10754,N_10833);
and U10994 (N_10994,N_10787,N_10866);
or U10995 (N_10995,N_10771,N_10781);
xor U10996 (N_10996,N_10860,N_10759);
nor U10997 (N_10997,N_10853,N_10862);
nor U10998 (N_10998,N_10830,N_10820);
nor U10999 (N_10999,N_10771,N_10759);
nor U11000 (N_11000,N_10955,N_10876);
and U11001 (N_11001,N_10934,N_10921);
nand U11002 (N_11002,N_10912,N_10940);
and U11003 (N_11003,N_10987,N_10936);
nor U11004 (N_11004,N_10883,N_10910);
xor U11005 (N_11005,N_10959,N_10970);
xnor U11006 (N_11006,N_10995,N_10957);
xor U11007 (N_11007,N_10996,N_10889);
or U11008 (N_11008,N_10964,N_10941);
xor U11009 (N_11009,N_10911,N_10960);
nand U11010 (N_11010,N_10985,N_10965);
xor U11011 (N_11011,N_10926,N_10950);
nand U11012 (N_11012,N_10875,N_10978);
or U11013 (N_11013,N_10902,N_10947);
and U11014 (N_11014,N_10887,N_10915);
or U11015 (N_11015,N_10924,N_10945);
xnor U11016 (N_11016,N_10882,N_10937);
nor U11017 (N_11017,N_10962,N_10949);
xnor U11018 (N_11018,N_10899,N_10886);
and U11019 (N_11019,N_10977,N_10929);
nor U11020 (N_11020,N_10956,N_10923);
nand U11021 (N_11021,N_10999,N_10958);
nand U11022 (N_11022,N_10991,N_10907);
xnor U11023 (N_11023,N_10988,N_10908);
nor U11024 (N_11024,N_10881,N_10946);
nand U11025 (N_11025,N_10884,N_10896);
nor U11026 (N_11026,N_10888,N_10925);
or U11027 (N_11027,N_10933,N_10984);
or U11028 (N_11028,N_10990,N_10976);
and U11029 (N_11029,N_10890,N_10952);
xor U11030 (N_11030,N_10944,N_10967);
or U11031 (N_11031,N_10993,N_10916);
nand U11032 (N_11032,N_10894,N_10909);
xor U11033 (N_11033,N_10939,N_10906);
or U11034 (N_11034,N_10974,N_10892);
nor U11035 (N_11035,N_10966,N_10877);
nor U11036 (N_11036,N_10903,N_10953);
nor U11037 (N_11037,N_10922,N_10969);
or U11038 (N_11038,N_10880,N_10973);
nand U11039 (N_11039,N_10900,N_10963);
or U11040 (N_11040,N_10986,N_10917);
nand U11041 (N_11041,N_10983,N_10975);
and U11042 (N_11042,N_10972,N_10885);
nand U11043 (N_11043,N_10931,N_10997);
nor U11044 (N_11044,N_10914,N_10954);
and U11045 (N_11045,N_10992,N_10920);
nand U11046 (N_11046,N_10895,N_10981);
nand U11047 (N_11047,N_10893,N_10971);
or U11048 (N_11048,N_10968,N_10979);
xnor U11049 (N_11049,N_10994,N_10989);
or U11050 (N_11050,N_10879,N_10898);
xnor U11051 (N_11051,N_10982,N_10998);
nor U11052 (N_11052,N_10901,N_10943);
nor U11053 (N_11053,N_10951,N_10948);
xnor U11054 (N_11054,N_10961,N_10878);
xor U11055 (N_11055,N_10980,N_10935);
and U11056 (N_11056,N_10932,N_10905);
nand U11057 (N_11057,N_10919,N_10927);
and U11058 (N_11058,N_10897,N_10913);
or U11059 (N_11059,N_10904,N_10938);
nor U11060 (N_11060,N_10891,N_10918);
nand U11061 (N_11061,N_10930,N_10942);
xor U11062 (N_11062,N_10928,N_10932);
and U11063 (N_11063,N_10954,N_10898);
nand U11064 (N_11064,N_10946,N_10903);
nand U11065 (N_11065,N_10999,N_10930);
and U11066 (N_11066,N_10936,N_10934);
or U11067 (N_11067,N_10984,N_10884);
nand U11068 (N_11068,N_10946,N_10886);
nand U11069 (N_11069,N_10970,N_10891);
nand U11070 (N_11070,N_10966,N_10916);
nand U11071 (N_11071,N_10878,N_10900);
and U11072 (N_11072,N_10942,N_10953);
xnor U11073 (N_11073,N_10990,N_10983);
xnor U11074 (N_11074,N_10995,N_10941);
and U11075 (N_11075,N_10980,N_10982);
nor U11076 (N_11076,N_10906,N_10966);
xnor U11077 (N_11077,N_10881,N_10931);
and U11078 (N_11078,N_10956,N_10888);
nand U11079 (N_11079,N_10971,N_10977);
nor U11080 (N_11080,N_10914,N_10876);
nand U11081 (N_11081,N_10975,N_10889);
nand U11082 (N_11082,N_10968,N_10906);
nor U11083 (N_11083,N_10891,N_10906);
and U11084 (N_11084,N_10896,N_10882);
nand U11085 (N_11085,N_10954,N_10890);
and U11086 (N_11086,N_10933,N_10996);
nor U11087 (N_11087,N_10888,N_10959);
nor U11088 (N_11088,N_10876,N_10946);
xnor U11089 (N_11089,N_10967,N_10958);
xnor U11090 (N_11090,N_10945,N_10951);
xnor U11091 (N_11091,N_10982,N_10913);
or U11092 (N_11092,N_10926,N_10958);
nand U11093 (N_11093,N_10911,N_10963);
nor U11094 (N_11094,N_10961,N_10993);
nand U11095 (N_11095,N_10911,N_10880);
nor U11096 (N_11096,N_10960,N_10971);
or U11097 (N_11097,N_10978,N_10974);
nor U11098 (N_11098,N_10964,N_10929);
nand U11099 (N_11099,N_10961,N_10915);
nor U11100 (N_11100,N_10958,N_10941);
and U11101 (N_11101,N_10883,N_10980);
xor U11102 (N_11102,N_10966,N_10881);
nand U11103 (N_11103,N_10985,N_10876);
xnor U11104 (N_11104,N_10986,N_10962);
nand U11105 (N_11105,N_10892,N_10913);
and U11106 (N_11106,N_10917,N_10941);
xor U11107 (N_11107,N_10945,N_10888);
nand U11108 (N_11108,N_10961,N_10952);
nor U11109 (N_11109,N_10983,N_10993);
nand U11110 (N_11110,N_10960,N_10961);
xnor U11111 (N_11111,N_10923,N_10894);
xnor U11112 (N_11112,N_10989,N_10928);
or U11113 (N_11113,N_10923,N_10888);
or U11114 (N_11114,N_10930,N_10899);
and U11115 (N_11115,N_10994,N_10979);
and U11116 (N_11116,N_10999,N_10952);
xnor U11117 (N_11117,N_10888,N_10891);
nor U11118 (N_11118,N_10878,N_10953);
nor U11119 (N_11119,N_10946,N_10983);
and U11120 (N_11120,N_10978,N_10959);
or U11121 (N_11121,N_10939,N_10934);
nand U11122 (N_11122,N_10967,N_10906);
nor U11123 (N_11123,N_10947,N_10900);
nor U11124 (N_11124,N_10884,N_10938);
and U11125 (N_11125,N_11020,N_11109);
xor U11126 (N_11126,N_11074,N_11013);
and U11127 (N_11127,N_11025,N_11064);
and U11128 (N_11128,N_11040,N_11017);
xor U11129 (N_11129,N_11090,N_11079);
or U11130 (N_11130,N_11031,N_11097);
nor U11131 (N_11131,N_11016,N_11118);
and U11132 (N_11132,N_11052,N_11026);
or U11133 (N_11133,N_11093,N_11063);
nor U11134 (N_11134,N_11046,N_11080);
xnor U11135 (N_11135,N_11022,N_11023);
and U11136 (N_11136,N_11009,N_11120);
nand U11137 (N_11137,N_11030,N_11027);
nor U11138 (N_11138,N_11028,N_11113);
nand U11139 (N_11139,N_11123,N_11011);
xor U11140 (N_11140,N_11024,N_11049);
and U11141 (N_11141,N_11057,N_11065);
and U11142 (N_11142,N_11042,N_11048);
xor U11143 (N_11143,N_11116,N_11095);
and U11144 (N_11144,N_11088,N_11117);
nor U11145 (N_11145,N_11000,N_11102);
nor U11146 (N_11146,N_11043,N_11121);
nor U11147 (N_11147,N_11050,N_11099);
nand U11148 (N_11148,N_11094,N_11003);
or U11149 (N_11149,N_11119,N_11053);
and U11150 (N_11150,N_11107,N_11037);
or U11151 (N_11151,N_11014,N_11012);
xnor U11152 (N_11152,N_11045,N_11007);
nand U11153 (N_11153,N_11056,N_11115);
nand U11154 (N_11154,N_11008,N_11066);
nand U11155 (N_11155,N_11082,N_11104);
nand U11156 (N_11156,N_11069,N_11114);
nor U11157 (N_11157,N_11038,N_11015);
and U11158 (N_11158,N_11071,N_11033);
nand U11159 (N_11159,N_11077,N_11036);
nor U11160 (N_11160,N_11112,N_11061);
or U11161 (N_11161,N_11047,N_11096);
nand U11162 (N_11162,N_11086,N_11006);
and U11163 (N_11163,N_11092,N_11068);
nand U11164 (N_11164,N_11041,N_11083);
nor U11165 (N_11165,N_11089,N_11058);
nor U11166 (N_11166,N_11039,N_11076);
nor U11167 (N_11167,N_11098,N_11073);
or U11168 (N_11168,N_11070,N_11067);
or U11169 (N_11169,N_11111,N_11062);
or U11170 (N_11170,N_11124,N_11010);
or U11171 (N_11171,N_11075,N_11029);
xor U11172 (N_11172,N_11019,N_11085);
or U11173 (N_11173,N_11005,N_11004);
or U11174 (N_11174,N_11032,N_11091);
or U11175 (N_11175,N_11072,N_11101);
nand U11176 (N_11176,N_11059,N_11002);
or U11177 (N_11177,N_11087,N_11021);
nand U11178 (N_11178,N_11100,N_11105);
or U11179 (N_11179,N_11122,N_11044);
and U11180 (N_11180,N_11035,N_11110);
nor U11181 (N_11181,N_11060,N_11078);
xnor U11182 (N_11182,N_11034,N_11106);
or U11183 (N_11183,N_11108,N_11001);
nor U11184 (N_11184,N_11084,N_11055);
and U11185 (N_11185,N_11081,N_11018);
nand U11186 (N_11186,N_11054,N_11103);
nand U11187 (N_11187,N_11051,N_11121);
and U11188 (N_11188,N_11112,N_11004);
nor U11189 (N_11189,N_11120,N_11124);
nor U11190 (N_11190,N_11092,N_11040);
nand U11191 (N_11191,N_11024,N_11000);
or U11192 (N_11192,N_11120,N_11017);
and U11193 (N_11193,N_11095,N_11103);
xor U11194 (N_11194,N_11030,N_11012);
nor U11195 (N_11195,N_11003,N_11064);
nand U11196 (N_11196,N_11087,N_11035);
and U11197 (N_11197,N_11077,N_11000);
and U11198 (N_11198,N_11086,N_11046);
xor U11199 (N_11199,N_11078,N_11071);
nand U11200 (N_11200,N_11024,N_11112);
nand U11201 (N_11201,N_11014,N_11045);
nand U11202 (N_11202,N_11067,N_11043);
nand U11203 (N_11203,N_11063,N_11038);
nor U11204 (N_11204,N_11123,N_11059);
nand U11205 (N_11205,N_11058,N_11122);
or U11206 (N_11206,N_11049,N_11068);
and U11207 (N_11207,N_11120,N_11107);
nor U11208 (N_11208,N_11011,N_11083);
or U11209 (N_11209,N_11069,N_11031);
nand U11210 (N_11210,N_11020,N_11001);
nand U11211 (N_11211,N_11076,N_11056);
or U11212 (N_11212,N_11049,N_11022);
or U11213 (N_11213,N_11074,N_11043);
nor U11214 (N_11214,N_11090,N_11068);
and U11215 (N_11215,N_11069,N_11090);
nand U11216 (N_11216,N_11031,N_11024);
and U11217 (N_11217,N_11109,N_11124);
nand U11218 (N_11218,N_11036,N_11001);
and U11219 (N_11219,N_11073,N_11042);
xnor U11220 (N_11220,N_11023,N_11076);
and U11221 (N_11221,N_11029,N_11107);
nand U11222 (N_11222,N_11021,N_11012);
and U11223 (N_11223,N_11096,N_11054);
or U11224 (N_11224,N_11038,N_11092);
nor U11225 (N_11225,N_11098,N_11024);
or U11226 (N_11226,N_11025,N_11081);
nand U11227 (N_11227,N_11040,N_11117);
nor U11228 (N_11228,N_11097,N_11011);
xor U11229 (N_11229,N_11081,N_11036);
nor U11230 (N_11230,N_11120,N_11092);
nand U11231 (N_11231,N_11057,N_11095);
nor U11232 (N_11232,N_11044,N_11120);
nor U11233 (N_11233,N_11097,N_11065);
nor U11234 (N_11234,N_11017,N_11098);
or U11235 (N_11235,N_11067,N_11044);
or U11236 (N_11236,N_11105,N_11058);
and U11237 (N_11237,N_11042,N_11023);
and U11238 (N_11238,N_11114,N_11112);
and U11239 (N_11239,N_11039,N_11089);
xor U11240 (N_11240,N_11027,N_11123);
xnor U11241 (N_11241,N_11074,N_11037);
xnor U11242 (N_11242,N_11062,N_11044);
or U11243 (N_11243,N_11008,N_11022);
or U11244 (N_11244,N_11068,N_11010);
nor U11245 (N_11245,N_11005,N_11085);
or U11246 (N_11246,N_11091,N_11100);
nor U11247 (N_11247,N_11002,N_11083);
nor U11248 (N_11248,N_11124,N_11104);
or U11249 (N_11249,N_11091,N_11045);
nor U11250 (N_11250,N_11140,N_11166);
xor U11251 (N_11251,N_11144,N_11164);
nand U11252 (N_11252,N_11243,N_11229);
xor U11253 (N_11253,N_11141,N_11177);
nand U11254 (N_11254,N_11242,N_11218);
and U11255 (N_11255,N_11220,N_11215);
or U11256 (N_11256,N_11226,N_11214);
nand U11257 (N_11257,N_11222,N_11155);
or U11258 (N_11258,N_11247,N_11148);
xnor U11259 (N_11259,N_11162,N_11188);
nor U11260 (N_11260,N_11216,N_11134);
xnor U11261 (N_11261,N_11232,N_11126);
xnor U11262 (N_11262,N_11190,N_11183);
nor U11263 (N_11263,N_11241,N_11153);
nand U11264 (N_11264,N_11187,N_11131);
nor U11265 (N_11265,N_11202,N_11201);
and U11266 (N_11266,N_11150,N_11180);
nor U11267 (N_11267,N_11221,N_11132);
and U11268 (N_11268,N_11173,N_11240);
nand U11269 (N_11269,N_11195,N_11125);
nand U11270 (N_11270,N_11175,N_11204);
xor U11271 (N_11271,N_11233,N_11239);
xnor U11272 (N_11272,N_11182,N_11217);
nor U11273 (N_11273,N_11196,N_11244);
xor U11274 (N_11274,N_11205,N_11209);
or U11275 (N_11275,N_11186,N_11228);
xnor U11276 (N_11276,N_11169,N_11178);
nor U11277 (N_11277,N_11245,N_11230);
and U11278 (N_11278,N_11189,N_11197);
xnor U11279 (N_11279,N_11158,N_11168);
nor U11280 (N_11280,N_11185,N_11200);
xor U11281 (N_11281,N_11129,N_11149);
xor U11282 (N_11282,N_11194,N_11238);
nor U11283 (N_11283,N_11223,N_11213);
or U11284 (N_11284,N_11234,N_11151);
xor U11285 (N_11285,N_11237,N_11210);
nor U11286 (N_11286,N_11224,N_11193);
xnor U11287 (N_11287,N_11248,N_11137);
nand U11288 (N_11288,N_11143,N_11211);
xnor U11289 (N_11289,N_11225,N_11179);
xnor U11290 (N_11290,N_11147,N_11246);
nand U11291 (N_11291,N_11249,N_11163);
or U11292 (N_11292,N_11174,N_11172);
nor U11293 (N_11293,N_11231,N_11127);
nand U11294 (N_11294,N_11154,N_11138);
nand U11295 (N_11295,N_11171,N_11184);
xnor U11296 (N_11296,N_11145,N_11136);
nand U11297 (N_11297,N_11192,N_11156);
and U11298 (N_11298,N_11176,N_11128);
nand U11299 (N_11299,N_11135,N_11207);
or U11300 (N_11300,N_11236,N_11142);
nand U11301 (N_11301,N_11152,N_11206);
and U11302 (N_11302,N_11160,N_11203);
nor U11303 (N_11303,N_11139,N_11199);
and U11304 (N_11304,N_11159,N_11167);
and U11305 (N_11305,N_11165,N_11208);
nand U11306 (N_11306,N_11133,N_11146);
xnor U11307 (N_11307,N_11170,N_11161);
xnor U11308 (N_11308,N_11157,N_11191);
or U11309 (N_11309,N_11181,N_11235);
nand U11310 (N_11310,N_11212,N_11219);
xor U11311 (N_11311,N_11227,N_11198);
xor U11312 (N_11312,N_11130,N_11138);
and U11313 (N_11313,N_11151,N_11220);
xnor U11314 (N_11314,N_11234,N_11192);
nor U11315 (N_11315,N_11126,N_11159);
nand U11316 (N_11316,N_11187,N_11237);
xor U11317 (N_11317,N_11231,N_11156);
nor U11318 (N_11318,N_11226,N_11171);
nand U11319 (N_11319,N_11195,N_11183);
nand U11320 (N_11320,N_11155,N_11227);
or U11321 (N_11321,N_11186,N_11235);
or U11322 (N_11322,N_11203,N_11175);
nand U11323 (N_11323,N_11246,N_11159);
xnor U11324 (N_11324,N_11197,N_11157);
nor U11325 (N_11325,N_11199,N_11141);
xor U11326 (N_11326,N_11217,N_11179);
nand U11327 (N_11327,N_11242,N_11208);
or U11328 (N_11328,N_11170,N_11197);
nand U11329 (N_11329,N_11134,N_11211);
and U11330 (N_11330,N_11160,N_11241);
nand U11331 (N_11331,N_11159,N_11161);
nor U11332 (N_11332,N_11163,N_11177);
nor U11333 (N_11333,N_11183,N_11187);
nor U11334 (N_11334,N_11196,N_11213);
xnor U11335 (N_11335,N_11154,N_11242);
xor U11336 (N_11336,N_11132,N_11193);
nand U11337 (N_11337,N_11209,N_11165);
xor U11338 (N_11338,N_11125,N_11244);
nor U11339 (N_11339,N_11228,N_11235);
or U11340 (N_11340,N_11236,N_11249);
nor U11341 (N_11341,N_11176,N_11164);
and U11342 (N_11342,N_11202,N_11189);
nor U11343 (N_11343,N_11173,N_11216);
nand U11344 (N_11344,N_11142,N_11152);
nand U11345 (N_11345,N_11233,N_11142);
and U11346 (N_11346,N_11158,N_11247);
nor U11347 (N_11347,N_11212,N_11171);
nor U11348 (N_11348,N_11238,N_11188);
and U11349 (N_11349,N_11126,N_11154);
nor U11350 (N_11350,N_11235,N_11133);
and U11351 (N_11351,N_11184,N_11177);
and U11352 (N_11352,N_11166,N_11240);
nand U11353 (N_11353,N_11137,N_11224);
and U11354 (N_11354,N_11135,N_11245);
xnor U11355 (N_11355,N_11218,N_11131);
and U11356 (N_11356,N_11192,N_11195);
or U11357 (N_11357,N_11167,N_11237);
xor U11358 (N_11358,N_11145,N_11174);
or U11359 (N_11359,N_11241,N_11168);
or U11360 (N_11360,N_11239,N_11212);
or U11361 (N_11361,N_11228,N_11193);
nand U11362 (N_11362,N_11235,N_11172);
and U11363 (N_11363,N_11133,N_11200);
nor U11364 (N_11364,N_11192,N_11243);
nand U11365 (N_11365,N_11239,N_11231);
nand U11366 (N_11366,N_11200,N_11177);
nor U11367 (N_11367,N_11207,N_11225);
and U11368 (N_11368,N_11188,N_11200);
xnor U11369 (N_11369,N_11143,N_11163);
or U11370 (N_11370,N_11217,N_11128);
nand U11371 (N_11371,N_11199,N_11164);
nand U11372 (N_11372,N_11229,N_11225);
nor U11373 (N_11373,N_11196,N_11136);
nand U11374 (N_11374,N_11203,N_11170);
or U11375 (N_11375,N_11288,N_11320);
or U11376 (N_11376,N_11305,N_11309);
nand U11377 (N_11377,N_11364,N_11265);
and U11378 (N_11378,N_11303,N_11337);
xnor U11379 (N_11379,N_11319,N_11297);
nand U11380 (N_11380,N_11322,N_11366);
nor U11381 (N_11381,N_11277,N_11349);
nand U11382 (N_11382,N_11283,N_11291);
or U11383 (N_11383,N_11374,N_11368);
or U11384 (N_11384,N_11345,N_11369);
or U11385 (N_11385,N_11346,N_11355);
xnor U11386 (N_11386,N_11284,N_11257);
or U11387 (N_11387,N_11372,N_11348);
and U11388 (N_11388,N_11271,N_11285);
or U11389 (N_11389,N_11344,N_11365);
nand U11390 (N_11390,N_11316,N_11286);
and U11391 (N_11391,N_11292,N_11282);
or U11392 (N_11392,N_11312,N_11264);
or U11393 (N_11393,N_11301,N_11325);
nand U11394 (N_11394,N_11278,N_11304);
nand U11395 (N_11395,N_11335,N_11317);
and U11396 (N_11396,N_11332,N_11266);
nor U11397 (N_11397,N_11333,N_11347);
nor U11398 (N_11398,N_11358,N_11315);
xor U11399 (N_11399,N_11294,N_11270);
and U11400 (N_11400,N_11362,N_11261);
or U11401 (N_11401,N_11253,N_11295);
xor U11402 (N_11402,N_11326,N_11371);
and U11403 (N_11403,N_11354,N_11339);
and U11404 (N_11404,N_11328,N_11268);
or U11405 (N_11405,N_11280,N_11334);
nand U11406 (N_11406,N_11308,N_11272);
nor U11407 (N_11407,N_11323,N_11298);
and U11408 (N_11408,N_11356,N_11363);
nor U11409 (N_11409,N_11299,N_11342);
or U11410 (N_11410,N_11330,N_11256);
xor U11411 (N_11411,N_11359,N_11350);
xnor U11412 (N_11412,N_11273,N_11293);
xor U11413 (N_11413,N_11289,N_11343);
or U11414 (N_11414,N_11275,N_11267);
and U11415 (N_11415,N_11357,N_11311);
xnor U11416 (N_11416,N_11338,N_11281);
and U11417 (N_11417,N_11353,N_11321);
nor U11418 (N_11418,N_11314,N_11262);
nand U11419 (N_11419,N_11331,N_11263);
and U11420 (N_11420,N_11300,N_11290);
or U11421 (N_11421,N_11279,N_11370);
and U11422 (N_11422,N_11250,N_11361);
nand U11423 (N_11423,N_11276,N_11313);
nor U11424 (N_11424,N_11306,N_11254);
or U11425 (N_11425,N_11324,N_11341);
or U11426 (N_11426,N_11274,N_11269);
xnor U11427 (N_11427,N_11258,N_11259);
and U11428 (N_11428,N_11340,N_11336);
and U11429 (N_11429,N_11373,N_11367);
or U11430 (N_11430,N_11307,N_11296);
xor U11431 (N_11431,N_11327,N_11329);
or U11432 (N_11432,N_11252,N_11287);
or U11433 (N_11433,N_11260,N_11352);
xnor U11434 (N_11434,N_11251,N_11310);
and U11435 (N_11435,N_11302,N_11318);
xor U11436 (N_11436,N_11255,N_11360);
nand U11437 (N_11437,N_11351,N_11353);
and U11438 (N_11438,N_11331,N_11352);
and U11439 (N_11439,N_11310,N_11361);
or U11440 (N_11440,N_11336,N_11306);
and U11441 (N_11441,N_11288,N_11279);
nor U11442 (N_11442,N_11341,N_11280);
xor U11443 (N_11443,N_11317,N_11372);
or U11444 (N_11444,N_11307,N_11255);
and U11445 (N_11445,N_11335,N_11312);
or U11446 (N_11446,N_11343,N_11252);
or U11447 (N_11447,N_11361,N_11355);
nor U11448 (N_11448,N_11297,N_11309);
or U11449 (N_11449,N_11335,N_11328);
and U11450 (N_11450,N_11367,N_11294);
xnor U11451 (N_11451,N_11346,N_11282);
and U11452 (N_11452,N_11372,N_11327);
and U11453 (N_11453,N_11373,N_11268);
or U11454 (N_11454,N_11272,N_11295);
or U11455 (N_11455,N_11335,N_11351);
nand U11456 (N_11456,N_11326,N_11277);
or U11457 (N_11457,N_11369,N_11269);
or U11458 (N_11458,N_11304,N_11269);
and U11459 (N_11459,N_11332,N_11302);
nor U11460 (N_11460,N_11271,N_11260);
nand U11461 (N_11461,N_11266,N_11283);
and U11462 (N_11462,N_11304,N_11279);
or U11463 (N_11463,N_11369,N_11364);
or U11464 (N_11464,N_11326,N_11253);
and U11465 (N_11465,N_11295,N_11349);
nand U11466 (N_11466,N_11297,N_11259);
nand U11467 (N_11467,N_11296,N_11284);
xnor U11468 (N_11468,N_11365,N_11337);
nor U11469 (N_11469,N_11345,N_11367);
xor U11470 (N_11470,N_11364,N_11359);
and U11471 (N_11471,N_11326,N_11346);
nand U11472 (N_11472,N_11365,N_11259);
xnor U11473 (N_11473,N_11310,N_11294);
nor U11474 (N_11474,N_11290,N_11337);
or U11475 (N_11475,N_11373,N_11281);
or U11476 (N_11476,N_11347,N_11372);
xnor U11477 (N_11477,N_11299,N_11349);
and U11478 (N_11478,N_11329,N_11320);
nor U11479 (N_11479,N_11300,N_11373);
or U11480 (N_11480,N_11293,N_11370);
or U11481 (N_11481,N_11338,N_11336);
and U11482 (N_11482,N_11272,N_11343);
and U11483 (N_11483,N_11308,N_11343);
or U11484 (N_11484,N_11268,N_11251);
xor U11485 (N_11485,N_11350,N_11340);
and U11486 (N_11486,N_11299,N_11358);
or U11487 (N_11487,N_11263,N_11306);
nor U11488 (N_11488,N_11287,N_11302);
or U11489 (N_11489,N_11282,N_11340);
or U11490 (N_11490,N_11324,N_11270);
and U11491 (N_11491,N_11303,N_11271);
nor U11492 (N_11492,N_11344,N_11260);
xnor U11493 (N_11493,N_11312,N_11305);
and U11494 (N_11494,N_11275,N_11367);
nand U11495 (N_11495,N_11302,N_11356);
nor U11496 (N_11496,N_11363,N_11264);
nor U11497 (N_11497,N_11265,N_11287);
and U11498 (N_11498,N_11328,N_11254);
xnor U11499 (N_11499,N_11297,N_11367);
or U11500 (N_11500,N_11465,N_11472);
and U11501 (N_11501,N_11461,N_11409);
nor U11502 (N_11502,N_11483,N_11473);
nand U11503 (N_11503,N_11450,N_11419);
xor U11504 (N_11504,N_11444,N_11448);
or U11505 (N_11505,N_11453,N_11435);
xor U11506 (N_11506,N_11449,N_11454);
nor U11507 (N_11507,N_11396,N_11385);
and U11508 (N_11508,N_11482,N_11430);
or U11509 (N_11509,N_11407,N_11457);
xor U11510 (N_11510,N_11437,N_11443);
nor U11511 (N_11511,N_11375,N_11428);
and U11512 (N_11512,N_11476,N_11411);
xor U11513 (N_11513,N_11418,N_11378);
nand U11514 (N_11514,N_11460,N_11478);
or U11515 (N_11515,N_11466,N_11467);
and U11516 (N_11516,N_11434,N_11459);
xnor U11517 (N_11517,N_11455,N_11391);
and U11518 (N_11518,N_11384,N_11489);
or U11519 (N_11519,N_11484,N_11416);
or U11520 (N_11520,N_11410,N_11399);
or U11521 (N_11521,N_11492,N_11441);
xor U11522 (N_11522,N_11417,N_11487);
nor U11523 (N_11523,N_11442,N_11490);
xor U11524 (N_11524,N_11382,N_11446);
xnor U11525 (N_11525,N_11408,N_11451);
nand U11526 (N_11526,N_11422,N_11377);
nand U11527 (N_11527,N_11423,N_11494);
and U11528 (N_11528,N_11447,N_11479);
or U11529 (N_11529,N_11421,N_11499);
or U11530 (N_11530,N_11398,N_11493);
and U11531 (N_11531,N_11456,N_11471);
nand U11532 (N_11532,N_11406,N_11431);
and U11533 (N_11533,N_11429,N_11438);
or U11534 (N_11534,N_11386,N_11393);
nand U11535 (N_11535,N_11425,N_11464);
nand U11536 (N_11536,N_11432,N_11394);
nand U11537 (N_11537,N_11498,N_11427);
nor U11538 (N_11538,N_11496,N_11475);
nor U11539 (N_11539,N_11470,N_11424);
nor U11540 (N_11540,N_11420,N_11445);
nand U11541 (N_11541,N_11388,N_11403);
nor U11542 (N_11542,N_11488,N_11426);
or U11543 (N_11543,N_11477,N_11486);
nor U11544 (N_11544,N_11390,N_11469);
xor U11545 (N_11545,N_11401,N_11405);
xnor U11546 (N_11546,N_11452,N_11497);
or U11547 (N_11547,N_11491,N_11415);
or U11548 (N_11548,N_11402,N_11440);
xnor U11549 (N_11549,N_11474,N_11413);
nand U11550 (N_11550,N_11404,N_11414);
or U11551 (N_11551,N_11392,N_11481);
xnor U11552 (N_11552,N_11412,N_11439);
nand U11553 (N_11553,N_11379,N_11380);
or U11554 (N_11554,N_11480,N_11376);
xnor U11555 (N_11555,N_11436,N_11395);
and U11556 (N_11556,N_11458,N_11383);
or U11557 (N_11557,N_11381,N_11389);
and U11558 (N_11558,N_11468,N_11397);
xnor U11559 (N_11559,N_11462,N_11485);
xor U11560 (N_11560,N_11387,N_11463);
xor U11561 (N_11561,N_11495,N_11433);
xnor U11562 (N_11562,N_11400,N_11380);
nand U11563 (N_11563,N_11465,N_11406);
and U11564 (N_11564,N_11430,N_11432);
or U11565 (N_11565,N_11409,N_11403);
nand U11566 (N_11566,N_11451,N_11438);
nor U11567 (N_11567,N_11467,N_11462);
nand U11568 (N_11568,N_11486,N_11393);
nand U11569 (N_11569,N_11409,N_11450);
or U11570 (N_11570,N_11414,N_11377);
xnor U11571 (N_11571,N_11438,N_11494);
or U11572 (N_11572,N_11388,N_11420);
xnor U11573 (N_11573,N_11413,N_11496);
xor U11574 (N_11574,N_11413,N_11461);
nor U11575 (N_11575,N_11495,N_11442);
or U11576 (N_11576,N_11429,N_11432);
and U11577 (N_11577,N_11440,N_11463);
nand U11578 (N_11578,N_11397,N_11434);
nand U11579 (N_11579,N_11428,N_11495);
or U11580 (N_11580,N_11444,N_11456);
or U11581 (N_11581,N_11481,N_11427);
and U11582 (N_11582,N_11400,N_11376);
nor U11583 (N_11583,N_11409,N_11415);
nand U11584 (N_11584,N_11442,N_11478);
and U11585 (N_11585,N_11497,N_11438);
xor U11586 (N_11586,N_11394,N_11436);
or U11587 (N_11587,N_11415,N_11380);
nand U11588 (N_11588,N_11447,N_11483);
nand U11589 (N_11589,N_11417,N_11474);
nor U11590 (N_11590,N_11430,N_11453);
nand U11591 (N_11591,N_11461,N_11381);
or U11592 (N_11592,N_11387,N_11461);
and U11593 (N_11593,N_11474,N_11486);
xor U11594 (N_11594,N_11407,N_11415);
nand U11595 (N_11595,N_11377,N_11490);
nor U11596 (N_11596,N_11418,N_11466);
nand U11597 (N_11597,N_11471,N_11467);
xnor U11598 (N_11598,N_11415,N_11452);
and U11599 (N_11599,N_11465,N_11474);
nand U11600 (N_11600,N_11493,N_11421);
nand U11601 (N_11601,N_11463,N_11446);
xor U11602 (N_11602,N_11390,N_11418);
xor U11603 (N_11603,N_11448,N_11456);
or U11604 (N_11604,N_11428,N_11388);
and U11605 (N_11605,N_11386,N_11420);
nor U11606 (N_11606,N_11397,N_11459);
nor U11607 (N_11607,N_11452,N_11413);
and U11608 (N_11608,N_11472,N_11461);
nand U11609 (N_11609,N_11487,N_11460);
xor U11610 (N_11610,N_11461,N_11424);
or U11611 (N_11611,N_11384,N_11493);
nor U11612 (N_11612,N_11499,N_11494);
and U11613 (N_11613,N_11474,N_11378);
and U11614 (N_11614,N_11448,N_11492);
and U11615 (N_11615,N_11382,N_11424);
or U11616 (N_11616,N_11376,N_11415);
or U11617 (N_11617,N_11426,N_11487);
xnor U11618 (N_11618,N_11470,N_11395);
xnor U11619 (N_11619,N_11459,N_11385);
or U11620 (N_11620,N_11457,N_11375);
xor U11621 (N_11621,N_11444,N_11474);
nand U11622 (N_11622,N_11393,N_11382);
and U11623 (N_11623,N_11472,N_11400);
xor U11624 (N_11624,N_11490,N_11462);
nor U11625 (N_11625,N_11510,N_11519);
xnor U11626 (N_11626,N_11541,N_11526);
or U11627 (N_11627,N_11528,N_11571);
or U11628 (N_11628,N_11582,N_11624);
xor U11629 (N_11629,N_11524,N_11566);
nor U11630 (N_11630,N_11618,N_11532);
nand U11631 (N_11631,N_11548,N_11513);
nor U11632 (N_11632,N_11504,N_11577);
and U11633 (N_11633,N_11515,N_11575);
xor U11634 (N_11634,N_11549,N_11563);
nand U11635 (N_11635,N_11505,N_11500);
and U11636 (N_11636,N_11611,N_11544);
and U11637 (N_11637,N_11557,N_11605);
nor U11638 (N_11638,N_11543,N_11597);
nor U11639 (N_11639,N_11570,N_11572);
xor U11640 (N_11640,N_11554,N_11591);
and U11641 (N_11641,N_11607,N_11603);
nor U11642 (N_11642,N_11531,N_11521);
xor U11643 (N_11643,N_11514,N_11621);
or U11644 (N_11644,N_11583,N_11527);
and U11645 (N_11645,N_11609,N_11517);
xor U11646 (N_11646,N_11562,N_11596);
or U11647 (N_11647,N_11550,N_11534);
and U11648 (N_11648,N_11602,N_11536);
nor U11649 (N_11649,N_11601,N_11599);
nor U11650 (N_11650,N_11606,N_11567);
nor U11651 (N_11651,N_11545,N_11556);
nand U11652 (N_11652,N_11580,N_11559);
nand U11653 (N_11653,N_11579,N_11574);
xor U11654 (N_11654,N_11530,N_11622);
nand U11655 (N_11655,N_11551,N_11581);
xor U11656 (N_11656,N_11509,N_11612);
and U11657 (N_11657,N_11589,N_11565);
nor U11658 (N_11658,N_11615,N_11529);
nand U11659 (N_11659,N_11560,N_11573);
nor U11660 (N_11660,N_11569,N_11542);
nand U11661 (N_11661,N_11588,N_11507);
and U11662 (N_11662,N_11568,N_11539);
xnor U11663 (N_11663,N_11546,N_11604);
nand U11664 (N_11664,N_11564,N_11614);
nor U11665 (N_11665,N_11585,N_11584);
nor U11666 (N_11666,N_11561,N_11533);
or U11667 (N_11667,N_11506,N_11520);
xor U11668 (N_11668,N_11553,N_11501);
nand U11669 (N_11669,N_11518,N_11587);
nand U11670 (N_11670,N_11525,N_11616);
xor U11671 (N_11671,N_11600,N_11512);
and U11672 (N_11672,N_11590,N_11578);
or U11673 (N_11673,N_11508,N_11523);
and U11674 (N_11674,N_11537,N_11592);
or U11675 (N_11675,N_11552,N_11516);
nor U11676 (N_11676,N_11598,N_11535);
xnor U11677 (N_11677,N_11522,N_11595);
and U11678 (N_11678,N_11576,N_11547);
xor U11679 (N_11679,N_11623,N_11503);
nand U11680 (N_11680,N_11617,N_11610);
xor U11681 (N_11681,N_11619,N_11538);
xnor U11682 (N_11682,N_11594,N_11502);
nand U11683 (N_11683,N_11555,N_11593);
nor U11684 (N_11684,N_11511,N_11540);
nor U11685 (N_11685,N_11558,N_11620);
nand U11686 (N_11686,N_11613,N_11608);
nor U11687 (N_11687,N_11586,N_11515);
nor U11688 (N_11688,N_11552,N_11601);
nand U11689 (N_11689,N_11549,N_11584);
xor U11690 (N_11690,N_11616,N_11622);
nor U11691 (N_11691,N_11560,N_11606);
nand U11692 (N_11692,N_11593,N_11549);
xnor U11693 (N_11693,N_11514,N_11574);
nand U11694 (N_11694,N_11552,N_11589);
and U11695 (N_11695,N_11543,N_11569);
or U11696 (N_11696,N_11514,N_11617);
and U11697 (N_11697,N_11616,N_11577);
or U11698 (N_11698,N_11608,N_11583);
and U11699 (N_11699,N_11572,N_11607);
and U11700 (N_11700,N_11577,N_11558);
nor U11701 (N_11701,N_11518,N_11584);
nor U11702 (N_11702,N_11537,N_11607);
or U11703 (N_11703,N_11543,N_11619);
xor U11704 (N_11704,N_11535,N_11522);
or U11705 (N_11705,N_11507,N_11597);
xor U11706 (N_11706,N_11604,N_11540);
xor U11707 (N_11707,N_11613,N_11521);
xor U11708 (N_11708,N_11545,N_11517);
xor U11709 (N_11709,N_11597,N_11574);
xnor U11710 (N_11710,N_11552,N_11570);
or U11711 (N_11711,N_11526,N_11624);
nor U11712 (N_11712,N_11621,N_11556);
or U11713 (N_11713,N_11580,N_11618);
or U11714 (N_11714,N_11550,N_11599);
xor U11715 (N_11715,N_11571,N_11620);
xnor U11716 (N_11716,N_11557,N_11507);
and U11717 (N_11717,N_11576,N_11603);
or U11718 (N_11718,N_11601,N_11512);
nor U11719 (N_11719,N_11612,N_11581);
xnor U11720 (N_11720,N_11514,N_11619);
xor U11721 (N_11721,N_11553,N_11526);
nor U11722 (N_11722,N_11585,N_11601);
nor U11723 (N_11723,N_11556,N_11584);
nand U11724 (N_11724,N_11501,N_11558);
or U11725 (N_11725,N_11541,N_11564);
or U11726 (N_11726,N_11585,N_11550);
and U11727 (N_11727,N_11590,N_11558);
nor U11728 (N_11728,N_11621,N_11589);
or U11729 (N_11729,N_11602,N_11622);
nand U11730 (N_11730,N_11515,N_11525);
and U11731 (N_11731,N_11592,N_11568);
or U11732 (N_11732,N_11616,N_11624);
nor U11733 (N_11733,N_11515,N_11528);
nand U11734 (N_11734,N_11606,N_11516);
and U11735 (N_11735,N_11533,N_11502);
and U11736 (N_11736,N_11607,N_11602);
xor U11737 (N_11737,N_11575,N_11501);
and U11738 (N_11738,N_11518,N_11545);
nor U11739 (N_11739,N_11507,N_11553);
or U11740 (N_11740,N_11555,N_11520);
or U11741 (N_11741,N_11510,N_11531);
nand U11742 (N_11742,N_11578,N_11601);
nor U11743 (N_11743,N_11515,N_11518);
or U11744 (N_11744,N_11600,N_11585);
or U11745 (N_11745,N_11553,N_11568);
and U11746 (N_11746,N_11506,N_11581);
nor U11747 (N_11747,N_11586,N_11502);
xor U11748 (N_11748,N_11549,N_11524);
nor U11749 (N_11749,N_11555,N_11609);
xor U11750 (N_11750,N_11700,N_11708);
nor U11751 (N_11751,N_11686,N_11645);
nor U11752 (N_11752,N_11681,N_11637);
nor U11753 (N_11753,N_11650,N_11732);
or U11754 (N_11754,N_11662,N_11736);
or U11755 (N_11755,N_11719,N_11715);
nand U11756 (N_11756,N_11655,N_11740);
nor U11757 (N_11757,N_11647,N_11717);
or U11758 (N_11758,N_11685,N_11633);
and U11759 (N_11759,N_11729,N_11742);
or U11760 (N_11760,N_11730,N_11677);
xor U11761 (N_11761,N_11628,N_11682);
nor U11762 (N_11762,N_11627,N_11687);
nor U11763 (N_11763,N_11716,N_11698);
or U11764 (N_11764,N_11705,N_11709);
nand U11765 (N_11765,N_11739,N_11651);
or U11766 (N_11766,N_11733,N_11672);
nor U11767 (N_11767,N_11718,N_11741);
and U11768 (N_11768,N_11663,N_11666);
nor U11769 (N_11769,N_11659,N_11643);
nor U11770 (N_11770,N_11638,N_11690);
and U11771 (N_11771,N_11722,N_11669);
or U11772 (N_11772,N_11629,N_11703);
nor U11773 (N_11773,N_11713,N_11695);
xor U11774 (N_11774,N_11679,N_11726);
and U11775 (N_11775,N_11671,N_11704);
nor U11776 (N_11776,N_11711,N_11693);
and U11777 (N_11777,N_11689,N_11684);
nand U11778 (N_11778,N_11696,N_11664);
or U11779 (N_11779,N_11652,N_11721);
nor U11780 (N_11780,N_11714,N_11646);
nor U11781 (N_11781,N_11680,N_11660);
nand U11782 (N_11782,N_11727,N_11744);
nand U11783 (N_11783,N_11735,N_11699);
nor U11784 (N_11784,N_11737,N_11747);
nand U11785 (N_11785,N_11707,N_11697);
and U11786 (N_11786,N_11745,N_11632);
xor U11787 (N_11787,N_11683,N_11720);
or U11788 (N_11788,N_11728,N_11670);
or U11789 (N_11789,N_11654,N_11641);
and U11790 (N_11790,N_11657,N_11626);
and U11791 (N_11791,N_11706,N_11631);
or U11792 (N_11792,N_11702,N_11743);
xnor U11793 (N_11793,N_11636,N_11749);
nor U11794 (N_11794,N_11653,N_11691);
or U11795 (N_11795,N_11658,N_11692);
nor U11796 (N_11796,N_11639,N_11640);
nor U11797 (N_11797,N_11649,N_11675);
nor U11798 (N_11798,N_11642,N_11644);
or U11799 (N_11799,N_11738,N_11688);
or U11800 (N_11800,N_11723,N_11731);
or U11801 (N_11801,N_11712,N_11676);
nand U11802 (N_11802,N_11630,N_11661);
xnor U11803 (N_11803,N_11625,N_11674);
or U11804 (N_11804,N_11725,N_11667);
xnor U11805 (N_11805,N_11635,N_11724);
xor U11806 (N_11806,N_11656,N_11648);
and U11807 (N_11807,N_11634,N_11734);
or U11808 (N_11808,N_11665,N_11710);
or U11809 (N_11809,N_11694,N_11701);
and U11810 (N_11810,N_11746,N_11668);
nand U11811 (N_11811,N_11748,N_11673);
nand U11812 (N_11812,N_11678,N_11712);
and U11813 (N_11813,N_11706,N_11647);
xor U11814 (N_11814,N_11731,N_11698);
and U11815 (N_11815,N_11667,N_11698);
nor U11816 (N_11816,N_11703,N_11687);
and U11817 (N_11817,N_11701,N_11699);
or U11818 (N_11818,N_11712,N_11640);
and U11819 (N_11819,N_11742,N_11628);
nand U11820 (N_11820,N_11650,N_11638);
nor U11821 (N_11821,N_11644,N_11726);
nor U11822 (N_11822,N_11694,N_11663);
and U11823 (N_11823,N_11739,N_11700);
xor U11824 (N_11824,N_11724,N_11742);
xnor U11825 (N_11825,N_11740,N_11719);
nand U11826 (N_11826,N_11677,N_11724);
or U11827 (N_11827,N_11684,N_11749);
and U11828 (N_11828,N_11740,N_11634);
nor U11829 (N_11829,N_11655,N_11679);
nor U11830 (N_11830,N_11633,N_11702);
and U11831 (N_11831,N_11711,N_11747);
or U11832 (N_11832,N_11724,N_11646);
nor U11833 (N_11833,N_11685,N_11638);
or U11834 (N_11834,N_11683,N_11677);
nand U11835 (N_11835,N_11736,N_11710);
xnor U11836 (N_11836,N_11718,N_11735);
or U11837 (N_11837,N_11717,N_11688);
and U11838 (N_11838,N_11711,N_11632);
nor U11839 (N_11839,N_11695,N_11640);
and U11840 (N_11840,N_11660,N_11675);
or U11841 (N_11841,N_11731,N_11722);
nor U11842 (N_11842,N_11722,N_11702);
nor U11843 (N_11843,N_11650,N_11689);
xnor U11844 (N_11844,N_11745,N_11700);
xor U11845 (N_11845,N_11653,N_11745);
xnor U11846 (N_11846,N_11714,N_11749);
nor U11847 (N_11847,N_11692,N_11739);
nor U11848 (N_11848,N_11709,N_11651);
nor U11849 (N_11849,N_11660,N_11677);
or U11850 (N_11850,N_11726,N_11687);
or U11851 (N_11851,N_11742,N_11671);
nor U11852 (N_11852,N_11632,N_11685);
nand U11853 (N_11853,N_11692,N_11736);
or U11854 (N_11854,N_11746,N_11674);
nor U11855 (N_11855,N_11713,N_11659);
and U11856 (N_11856,N_11746,N_11730);
or U11857 (N_11857,N_11640,N_11645);
or U11858 (N_11858,N_11625,N_11700);
and U11859 (N_11859,N_11722,N_11641);
xnor U11860 (N_11860,N_11735,N_11722);
and U11861 (N_11861,N_11701,N_11665);
nand U11862 (N_11862,N_11693,N_11740);
nand U11863 (N_11863,N_11666,N_11702);
nor U11864 (N_11864,N_11686,N_11718);
nor U11865 (N_11865,N_11704,N_11689);
nand U11866 (N_11866,N_11694,N_11724);
nor U11867 (N_11867,N_11709,N_11676);
and U11868 (N_11868,N_11726,N_11695);
nor U11869 (N_11869,N_11655,N_11696);
xnor U11870 (N_11870,N_11720,N_11658);
nand U11871 (N_11871,N_11629,N_11685);
nor U11872 (N_11872,N_11738,N_11631);
or U11873 (N_11873,N_11737,N_11652);
xnor U11874 (N_11874,N_11663,N_11658);
or U11875 (N_11875,N_11770,N_11849);
and U11876 (N_11876,N_11766,N_11862);
xor U11877 (N_11877,N_11807,N_11780);
and U11878 (N_11878,N_11762,N_11859);
xor U11879 (N_11879,N_11855,N_11751);
nor U11880 (N_11880,N_11767,N_11827);
nand U11881 (N_11881,N_11847,N_11823);
and U11882 (N_11882,N_11860,N_11870);
nand U11883 (N_11883,N_11818,N_11834);
or U11884 (N_11884,N_11777,N_11810);
nor U11885 (N_11885,N_11843,N_11757);
nand U11886 (N_11886,N_11836,N_11785);
or U11887 (N_11887,N_11853,N_11801);
nand U11888 (N_11888,N_11789,N_11851);
and U11889 (N_11889,N_11848,N_11799);
xnor U11890 (N_11890,N_11750,N_11873);
nand U11891 (N_11891,N_11779,N_11782);
and U11892 (N_11892,N_11763,N_11798);
and U11893 (N_11893,N_11771,N_11866);
and U11894 (N_11894,N_11815,N_11755);
nand U11895 (N_11895,N_11761,N_11788);
nor U11896 (N_11896,N_11800,N_11772);
and U11897 (N_11897,N_11787,N_11756);
nor U11898 (N_11898,N_11809,N_11857);
or U11899 (N_11899,N_11841,N_11858);
and U11900 (N_11900,N_11820,N_11812);
nor U11901 (N_11901,N_11765,N_11861);
or U11902 (N_11902,N_11792,N_11869);
nor U11903 (N_11903,N_11794,N_11838);
nand U11904 (N_11904,N_11835,N_11839);
and U11905 (N_11905,N_11790,N_11783);
nand U11906 (N_11906,N_11846,N_11774);
xnor U11907 (N_11907,N_11753,N_11797);
xor U11908 (N_11908,N_11872,N_11865);
nand U11909 (N_11909,N_11840,N_11842);
and U11910 (N_11910,N_11795,N_11850);
and U11911 (N_11911,N_11864,N_11829);
nor U11912 (N_11912,N_11806,N_11821);
or U11913 (N_11913,N_11811,N_11773);
or U11914 (N_11914,N_11808,N_11805);
and U11915 (N_11915,N_11837,N_11804);
and U11916 (N_11916,N_11819,N_11775);
xor U11917 (N_11917,N_11764,N_11874);
and U11918 (N_11918,N_11814,N_11754);
nand U11919 (N_11919,N_11752,N_11871);
xnor U11920 (N_11920,N_11803,N_11867);
or U11921 (N_11921,N_11816,N_11852);
and U11922 (N_11922,N_11786,N_11758);
nand U11923 (N_11923,N_11828,N_11796);
or U11924 (N_11924,N_11832,N_11813);
nand U11925 (N_11925,N_11854,N_11802);
nand U11926 (N_11926,N_11822,N_11791);
and U11927 (N_11927,N_11776,N_11824);
xor U11928 (N_11928,N_11759,N_11784);
nor U11929 (N_11929,N_11778,N_11826);
nor U11930 (N_11930,N_11781,N_11817);
nor U11931 (N_11931,N_11825,N_11856);
nor U11932 (N_11932,N_11793,N_11863);
nor U11933 (N_11933,N_11833,N_11831);
nand U11934 (N_11934,N_11769,N_11844);
or U11935 (N_11935,N_11845,N_11868);
and U11936 (N_11936,N_11760,N_11768);
nand U11937 (N_11937,N_11830,N_11757);
nor U11938 (N_11938,N_11858,N_11793);
xnor U11939 (N_11939,N_11859,N_11823);
and U11940 (N_11940,N_11844,N_11792);
or U11941 (N_11941,N_11802,N_11817);
nand U11942 (N_11942,N_11830,N_11766);
nand U11943 (N_11943,N_11849,N_11806);
and U11944 (N_11944,N_11834,N_11825);
and U11945 (N_11945,N_11872,N_11765);
or U11946 (N_11946,N_11830,N_11869);
xor U11947 (N_11947,N_11839,N_11769);
xnor U11948 (N_11948,N_11784,N_11863);
nor U11949 (N_11949,N_11788,N_11852);
and U11950 (N_11950,N_11783,N_11768);
nor U11951 (N_11951,N_11786,N_11790);
xnor U11952 (N_11952,N_11754,N_11774);
and U11953 (N_11953,N_11754,N_11869);
nand U11954 (N_11954,N_11812,N_11769);
nand U11955 (N_11955,N_11855,N_11849);
nand U11956 (N_11956,N_11822,N_11874);
nand U11957 (N_11957,N_11854,N_11805);
or U11958 (N_11958,N_11762,N_11802);
xnor U11959 (N_11959,N_11790,N_11835);
or U11960 (N_11960,N_11873,N_11755);
nor U11961 (N_11961,N_11756,N_11760);
nand U11962 (N_11962,N_11792,N_11813);
or U11963 (N_11963,N_11846,N_11779);
and U11964 (N_11964,N_11853,N_11768);
nand U11965 (N_11965,N_11828,N_11795);
or U11966 (N_11966,N_11821,N_11834);
or U11967 (N_11967,N_11844,N_11800);
nor U11968 (N_11968,N_11799,N_11852);
nand U11969 (N_11969,N_11785,N_11803);
xor U11970 (N_11970,N_11784,N_11860);
nand U11971 (N_11971,N_11856,N_11827);
nand U11972 (N_11972,N_11812,N_11843);
nand U11973 (N_11973,N_11799,N_11779);
xor U11974 (N_11974,N_11871,N_11809);
and U11975 (N_11975,N_11859,N_11842);
nand U11976 (N_11976,N_11787,N_11754);
or U11977 (N_11977,N_11788,N_11858);
and U11978 (N_11978,N_11758,N_11828);
nand U11979 (N_11979,N_11841,N_11859);
and U11980 (N_11980,N_11847,N_11765);
and U11981 (N_11981,N_11860,N_11850);
nand U11982 (N_11982,N_11789,N_11825);
and U11983 (N_11983,N_11808,N_11803);
and U11984 (N_11984,N_11845,N_11838);
nor U11985 (N_11985,N_11809,N_11842);
nor U11986 (N_11986,N_11821,N_11822);
or U11987 (N_11987,N_11847,N_11784);
nor U11988 (N_11988,N_11786,N_11860);
or U11989 (N_11989,N_11799,N_11844);
xnor U11990 (N_11990,N_11768,N_11823);
xnor U11991 (N_11991,N_11845,N_11862);
nor U11992 (N_11992,N_11772,N_11774);
xnor U11993 (N_11993,N_11766,N_11794);
nand U11994 (N_11994,N_11777,N_11833);
or U11995 (N_11995,N_11837,N_11868);
xor U11996 (N_11996,N_11757,N_11767);
and U11997 (N_11997,N_11789,N_11837);
and U11998 (N_11998,N_11836,N_11864);
xor U11999 (N_11999,N_11829,N_11806);
or U12000 (N_12000,N_11992,N_11940);
and U12001 (N_12001,N_11955,N_11917);
or U12002 (N_12002,N_11904,N_11979);
xor U12003 (N_12003,N_11893,N_11889);
and U12004 (N_12004,N_11910,N_11951);
xnor U12005 (N_12005,N_11954,N_11916);
xor U12006 (N_12006,N_11999,N_11898);
and U12007 (N_12007,N_11943,N_11989);
xor U12008 (N_12008,N_11931,N_11947);
nor U12009 (N_12009,N_11982,N_11965);
xor U12010 (N_12010,N_11974,N_11990);
nand U12011 (N_12011,N_11949,N_11977);
or U12012 (N_12012,N_11913,N_11983);
and U12013 (N_12013,N_11972,N_11875);
xor U12014 (N_12014,N_11883,N_11905);
nand U12015 (N_12015,N_11919,N_11876);
and U12016 (N_12016,N_11878,N_11900);
and U12017 (N_12017,N_11909,N_11994);
or U12018 (N_12018,N_11918,N_11894);
or U12019 (N_12019,N_11920,N_11890);
xnor U12020 (N_12020,N_11968,N_11901);
xnor U12021 (N_12021,N_11886,N_11888);
nor U12022 (N_12022,N_11932,N_11899);
and U12023 (N_12023,N_11958,N_11877);
nor U12024 (N_12024,N_11988,N_11880);
nor U12025 (N_12025,N_11936,N_11906);
nor U12026 (N_12026,N_11976,N_11928);
nand U12027 (N_12027,N_11925,N_11892);
and U12028 (N_12028,N_11957,N_11963);
and U12029 (N_12029,N_11978,N_11945);
nand U12030 (N_12030,N_11911,N_11950);
or U12031 (N_12031,N_11922,N_11896);
xnor U12032 (N_12032,N_11929,N_11907);
nand U12033 (N_12033,N_11998,N_11996);
nor U12034 (N_12034,N_11985,N_11882);
or U12035 (N_12035,N_11964,N_11956);
nor U12036 (N_12036,N_11946,N_11897);
xor U12037 (N_12037,N_11912,N_11961);
and U12038 (N_12038,N_11891,N_11970);
or U12039 (N_12039,N_11923,N_11881);
or U12040 (N_12040,N_11942,N_11980);
nor U12041 (N_12041,N_11987,N_11941);
and U12042 (N_12042,N_11937,N_11973);
or U12043 (N_12043,N_11966,N_11884);
nand U12044 (N_12044,N_11991,N_11935);
xnor U12045 (N_12045,N_11938,N_11887);
nand U12046 (N_12046,N_11952,N_11914);
nor U12047 (N_12047,N_11986,N_11993);
and U12048 (N_12048,N_11926,N_11967);
nor U12049 (N_12049,N_11948,N_11981);
xor U12050 (N_12050,N_11924,N_11930);
or U12051 (N_12051,N_11984,N_11939);
and U12052 (N_12052,N_11879,N_11885);
and U12053 (N_12053,N_11934,N_11962);
xor U12054 (N_12054,N_11921,N_11944);
nand U12055 (N_12055,N_11903,N_11960);
xnor U12056 (N_12056,N_11915,N_11902);
nand U12057 (N_12057,N_11927,N_11971);
xor U12058 (N_12058,N_11908,N_11997);
or U12059 (N_12059,N_11959,N_11969);
or U12060 (N_12060,N_11895,N_11933);
or U12061 (N_12061,N_11953,N_11975);
or U12062 (N_12062,N_11995,N_11946);
nand U12063 (N_12063,N_11933,N_11959);
xor U12064 (N_12064,N_11998,N_11902);
and U12065 (N_12065,N_11989,N_11983);
nor U12066 (N_12066,N_11995,N_11951);
and U12067 (N_12067,N_11949,N_11906);
nand U12068 (N_12068,N_11902,N_11997);
xor U12069 (N_12069,N_11949,N_11896);
xor U12070 (N_12070,N_11922,N_11883);
nor U12071 (N_12071,N_11971,N_11953);
nor U12072 (N_12072,N_11916,N_11880);
xnor U12073 (N_12073,N_11966,N_11982);
nor U12074 (N_12074,N_11877,N_11988);
or U12075 (N_12075,N_11962,N_11991);
and U12076 (N_12076,N_11898,N_11896);
and U12077 (N_12077,N_11993,N_11965);
and U12078 (N_12078,N_11966,N_11906);
nand U12079 (N_12079,N_11927,N_11921);
xnor U12080 (N_12080,N_11958,N_11961);
xnor U12081 (N_12081,N_11963,N_11967);
nand U12082 (N_12082,N_11948,N_11934);
nand U12083 (N_12083,N_11963,N_11960);
and U12084 (N_12084,N_11998,N_11995);
xor U12085 (N_12085,N_11994,N_11954);
or U12086 (N_12086,N_11942,N_11957);
nand U12087 (N_12087,N_11927,N_11966);
nand U12088 (N_12088,N_11932,N_11882);
and U12089 (N_12089,N_11902,N_11913);
xnor U12090 (N_12090,N_11910,N_11928);
xnor U12091 (N_12091,N_11979,N_11877);
nand U12092 (N_12092,N_11977,N_11895);
or U12093 (N_12093,N_11998,N_11876);
nand U12094 (N_12094,N_11928,N_11980);
nor U12095 (N_12095,N_11944,N_11908);
or U12096 (N_12096,N_11988,N_11909);
xor U12097 (N_12097,N_11950,N_11942);
nor U12098 (N_12098,N_11922,N_11908);
nand U12099 (N_12099,N_11892,N_11975);
nand U12100 (N_12100,N_11900,N_11944);
xor U12101 (N_12101,N_11927,N_11928);
and U12102 (N_12102,N_11954,N_11997);
or U12103 (N_12103,N_11957,N_11965);
xor U12104 (N_12104,N_11997,N_11996);
nand U12105 (N_12105,N_11977,N_11953);
or U12106 (N_12106,N_11927,N_11948);
and U12107 (N_12107,N_11980,N_11882);
nor U12108 (N_12108,N_11881,N_11936);
nor U12109 (N_12109,N_11898,N_11919);
or U12110 (N_12110,N_11920,N_11984);
nand U12111 (N_12111,N_11913,N_11973);
nor U12112 (N_12112,N_11889,N_11952);
nand U12113 (N_12113,N_11878,N_11950);
nand U12114 (N_12114,N_11945,N_11900);
or U12115 (N_12115,N_11978,N_11982);
and U12116 (N_12116,N_11897,N_11943);
nand U12117 (N_12117,N_11952,N_11922);
xnor U12118 (N_12118,N_11923,N_11974);
nand U12119 (N_12119,N_11907,N_11885);
nor U12120 (N_12120,N_11932,N_11964);
xor U12121 (N_12121,N_11919,N_11943);
nor U12122 (N_12122,N_11940,N_11981);
xor U12123 (N_12123,N_11999,N_11948);
nand U12124 (N_12124,N_11897,N_11992);
or U12125 (N_12125,N_12029,N_12001);
nor U12126 (N_12126,N_12074,N_12114);
and U12127 (N_12127,N_12084,N_12046);
nand U12128 (N_12128,N_12061,N_12078);
or U12129 (N_12129,N_12119,N_12092);
or U12130 (N_12130,N_12097,N_12003);
xor U12131 (N_12131,N_12017,N_12016);
xor U12132 (N_12132,N_12025,N_12073);
and U12133 (N_12133,N_12056,N_12039);
and U12134 (N_12134,N_12015,N_12008);
nor U12135 (N_12135,N_12040,N_12101);
or U12136 (N_12136,N_12090,N_12072);
and U12137 (N_12137,N_12045,N_12051);
and U12138 (N_12138,N_12018,N_12005);
and U12139 (N_12139,N_12027,N_12105);
xor U12140 (N_12140,N_12067,N_12120);
or U12141 (N_12141,N_12075,N_12026);
or U12142 (N_12142,N_12108,N_12011);
xor U12143 (N_12143,N_12116,N_12009);
nand U12144 (N_12144,N_12000,N_12110);
nor U12145 (N_12145,N_12047,N_12021);
xor U12146 (N_12146,N_12107,N_12080);
xnor U12147 (N_12147,N_12041,N_12062);
nor U12148 (N_12148,N_12004,N_12054);
and U12149 (N_12149,N_12082,N_12006);
and U12150 (N_12150,N_12057,N_12094);
nor U12151 (N_12151,N_12081,N_12099);
xnor U12152 (N_12152,N_12030,N_12065);
or U12153 (N_12153,N_12024,N_12034);
nor U12154 (N_12154,N_12118,N_12020);
nand U12155 (N_12155,N_12010,N_12071);
or U12156 (N_12156,N_12044,N_12070);
nand U12157 (N_12157,N_12106,N_12088);
nand U12158 (N_12158,N_12083,N_12066);
nor U12159 (N_12159,N_12022,N_12069);
and U12160 (N_12160,N_12013,N_12122);
and U12161 (N_12161,N_12037,N_12113);
and U12162 (N_12162,N_12058,N_12085);
xor U12163 (N_12163,N_12063,N_12035);
nand U12164 (N_12164,N_12033,N_12077);
nor U12165 (N_12165,N_12098,N_12096);
or U12166 (N_12166,N_12007,N_12059);
nor U12167 (N_12167,N_12031,N_12002);
nor U12168 (N_12168,N_12111,N_12050);
and U12169 (N_12169,N_12032,N_12093);
and U12170 (N_12170,N_12053,N_12112);
or U12171 (N_12171,N_12079,N_12068);
xor U12172 (N_12172,N_12087,N_12049);
or U12173 (N_12173,N_12028,N_12042);
xnor U12174 (N_12174,N_12052,N_12102);
nand U12175 (N_12175,N_12121,N_12036);
and U12176 (N_12176,N_12100,N_12043);
xor U12177 (N_12177,N_12115,N_12038);
or U12178 (N_12178,N_12012,N_12095);
and U12179 (N_12179,N_12104,N_12014);
or U12180 (N_12180,N_12109,N_12023);
or U12181 (N_12181,N_12124,N_12086);
nand U12182 (N_12182,N_12123,N_12117);
nand U12183 (N_12183,N_12019,N_12089);
nand U12184 (N_12184,N_12091,N_12103);
and U12185 (N_12185,N_12048,N_12076);
xnor U12186 (N_12186,N_12055,N_12064);
nand U12187 (N_12187,N_12060,N_12057);
and U12188 (N_12188,N_12017,N_12035);
or U12189 (N_12189,N_12034,N_12066);
and U12190 (N_12190,N_12055,N_12121);
nor U12191 (N_12191,N_12060,N_12020);
or U12192 (N_12192,N_12026,N_12095);
and U12193 (N_12193,N_12123,N_12029);
or U12194 (N_12194,N_12104,N_12025);
nor U12195 (N_12195,N_12031,N_12000);
nand U12196 (N_12196,N_12000,N_12074);
or U12197 (N_12197,N_12086,N_12003);
xor U12198 (N_12198,N_12007,N_12042);
and U12199 (N_12199,N_12087,N_12007);
and U12200 (N_12200,N_12024,N_12108);
and U12201 (N_12201,N_12108,N_12123);
nand U12202 (N_12202,N_12063,N_12028);
xnor U12203 (N_12203,N_12031,N_12071);
and U12204 (N_12204,N_12054,N_12029);
nor U12205 (N_12205,N_12047,N_12082);
nor U12206 (N_12206,N_12027,N_12078);
and U12207 (N_12207,N_12005,N_12087);
or U12208 (N_12208,N_12059,N_12056);
or U12209 (N_12209,N_12030,N_12021);
xor U12210 (N_12210,N_12111,N_12092);
nand U12211 (N_12211,N_12033,N_12056);
xnor U12212 (N_12212,N_12076,N_12047);
and U12213 (N_12213,N_12027,N_12065);
nor U12214 (N_12214,N_12059,N_12092);
nand U12215 (N_12215,N_12108,N_12060);
or U12216 (N_12216,N_12103,N_12039);
or U12217 (N_12217,N_12117,N_12075);
xor U12218 (N_12218,N_12092,N_12080);
or U12219 (N_12219,N_12035,N_12030);
xnor U12220 (N_12220,N_12121,N_12001);
or U12221 (N_12221,N_12056,N_12058);
and U12222 (N_12222,N_12060,N_12030);
and U12223 (N_12223,N_12010,N_12068);
nand U12224 (N_12224,N_12025,N_12054);
nor U12225 (N_12225,N_12023,N_12095);
nor U12226 (N_12226,N_12118,N_12044);
xnor U12227 (N_12227,N_12091,N_12019);
nor U12228 (N_12228,N_12056,N_12050);
and U12229 (N_12229,N_12085,N_12026);
nor U12230 (N_12230,N_12016,N_12042);
or U12231 (N_12231,N_12076,N_12078);
nor U12232 (N_12232,N_12003,N_12002);
xor U12233 (N_12233,N_12069,N_12078);
nor U12234 (N_12234,N_12123,N_12092);
or U12235 (N_12235,N_12006,N_12005);
or U12236 (N_12236,N_12117,N_12021);
nand U12237 (N_12237,N_12022,N_12103);
xor U12238 (N_12238,N_12035,N_12049);
xor U12239 (N_12239,N_12040,N_12089);
and U12240 (N_12240,N_12065,N_12105);
and U12241 (N_12241,N_12049,N_12072);
xor U12242 (N_12242,N_12017,N_12034);
or U12243 (N_12243,N_12100,N_12003);
nand U12244 (N_12244,N_12000,N_12070);
xnor U12245 (N_12245,N_12042,N_12047);
xnor U12246 (N_12246,N_12002,N_12105);
and U12247 (N_12247,N_12005,N_12110);
or U12248 (N_12248,N_12084,N_12092);
xor U12249 (N_12249,N_12035,N_12022);
and U12250 (N_12250,N_12170,N_12162);
nand U12251 (N_12251,N_12190,N_12214);
xnor U12252 (N_12252,N_12146,N_12210);
or U12253 (N_12253,N_12127,N_12248);
nor U12254 (N_12254,N_12174,N_12237);
xor U12255 (N_12255,N_12159,N_12219);
or U12256 (N_12256,N_12187,N_12129);
or U12257 (N_12257,N_12220,N_12239);
xnor U12258 (N_12258,N_12201,N_12236);
nor U12259 (N_12259,N_12185,N_12224);
and U12260 (N_12260,N_12143,N_12157);
nand U12261 (N_12261,N_12246,N_12227);
nor U12262 (N_12262,N_12206,N_12141);
and U12263 (N_12263,N_12166,N_12148);
nand U12264 (N_12264,N_12208,N_12238);
nand U12265 (N_12265,N_12173,N_12182);
or U12266 (N_12266,N_12126,N_12144);
xor U12267 (N_12267,N_12192,N_12131);
or U12268 (N_12268,N_12197,N_12149);
or U12269 (N_12269,N_12194,N_12135);
nand U12270 (N_12270,N_12142,N_12198);
or U12271 (N_12271,N_12223,N_12235);
and U12272 (N_12272,N_12152,N_12177);
and U12273 (N_12273,N_12195,N_12139);
and U12274 (N_12274,N_12172,N_12178);
xnor U12275 (N_12275,N_12154,N_12186);
xor U12276 (N_12276,N_12233,N_12232);
xor U12277 (N_12277,N_12245,N_12169);
and U12278 (N_12278,N_12132,N_12140);
and U12279 (N_12279,N_12189,N_12156);
xor U12280 (N_12280,N_12130,N_12171);
xor U12281 (N_12281,N_12193,N_12145);
and U12282 (N_12282,N_12138,N_12215);
or U12283 (N_12283,N_12168,N_12134);
xnor U12284 (N_12284,N_12242,N_12241);
or U12285 (N_12285,N_12228,N_12153);
and U12286 (N_12286,N_12133,N_12243);
nor U12287 (N_12287,N_12217,N_12125);
or U12288 (N_12288,N_12229,N_12222);
nor U12289 (N_12289,N_12183,N_12164);
nor U12290 (N_12290,N_12163,N_12176);
nor U12291 (N_12291,N_12200,N_12188);
nor U12292 (N_12292,N_12211,N_12207);
or U12293 (N_12293,N_12137,N_12158);
nor U12294 (N_12294,N_12181,N_12226);
nand U12295 (N_12295,N_12204,N_12244);
xnor U12296 (N_12296,N_12205,N_12199);
or U12297 (N_12297,N_12209,N_12128);
and U12298 (N_12298,N_12203,N_12213);
and U12299 (N_12299,N_12184,N_12225);
nor U12300 (N_12300,N_12216,N_12212);
and U12301 (N_12301,N_12191,N_12165);
and U12302 (N_12302,N_12150,N_12136);
and U12303 (N_12303,N_12247,N_12151);
nor U12304 (N_12304,N_12175,N_12167);
nor U12305 (N_12305,N_12249,N_12160);
xnor U12306 (N_12306,N_12231,N_12234);
or U12307 (N_12307,N_12218,N_12230);
and U12308 (N_12308,N_12147,N_12240);
and U12309 (N_12309,N_12179,N_12221);
xnor U12310 (N_12310,N_12196,N_12155);
nor U12311 (N_12311,N_12161,N_12180);
xnor U12312 (N_12312,N_12202,N_12184);
xor U12313 (N_12313,N_12226,N_12192);
or U12314 (N_12314,N_12228,N_12125);
and U12315 (N_12315,N_12125,N_12133);
xor U12316 (N_12316,N_12174,N_12204);
nand U12317 (N_12317,N_12213,N_12193);
nor U12318 (N_12318,N_12184,N_12170);
xor U12319 (N_12319,N_12225,N_12191);
xnor U12320 (N_12320,N_12172,N_12199);
nor U12321 (N_12321,N_12213,N_12175);
nand U12322 (N_12322,N_12220,N_12211);
and U12323 (N_12323,N_12198,N_12222);
or U12324 (N_12324,N_12150,N_12197);
nor U12325 (N_12325,N_12247,N_12180);
xor U12326 (N_12326,N_12216,N_12204);
nand U12327 (N_12327,N_12193,N_12159);
nand U12328 (N_12328,N_12175,N_12201);
and U12329 (N_12329,N_12246,N_12232);
nor U12330 (N_12330,N_12197,N_12233);
or U12331 (N_12331,N_12239,N_12173);
and U12332 (N_12332,N_12203,N_12177);
nor U12333 (N_12333,N_12204,N_12229);
nor U12334 (N_12334,N_12200,N_12192);
and U12335 (N_12335,N_12176,N_12212);
and U12336 (N_12336,N_12226,N_12187);
nor U12337 (N_12337,N_12193,N_12227);
and U12338 (N_12338,N_12197,N_12136);
nand U12339 (N_12339,N_12207,N_12188);
or U12340 (N_12340,N_12194,N_12196);
nor U12341 (N_12341,N_12138,N_12248);
nor U12342 (N_12342,N_12188,N_12131);
and U12343 (N_12343,N_12237,N_12155);
or U12344 (N_12344,N_12148,N_12245);
nor U12345 (N_12345,N_12229,N_12166);
and U12346 (N_12346,N_12242,N_12199);
nand U12347 (N_12347,N_12156,N_12214);
nor U12348 (N_12348,N_12247,N_12217);
or U12349 (N_12349,N_12138,N_12218);
or U12350 (N_12350,N_12171,N_12246);
xnor U12351 (N_12351,N_12131,N_12128);
xor U12352 (N_12352,N_12226,N_12184);
nor U12353 (N_12353,N_12233,N_12142);
nor U12354 (N_12354,N_12230,N_12206);
or U12355 (N_12355,N_12202,N_12197);
or U12356 (N_12356,N_12177,N_12157);
nand U12357 (N_12357,N_12168,N_12184);
xnor U12358 (N_12358,N_12152,N_12138);
and U12359 (N_12359,N_12175,N_12165);
or U12360 (N_12360,N_12243,N_12126);
and U12361 (N_12361,N_12156,N_12237);
and U12362 (N_12362,N_12194,N_12147);
nor U12363 (N_12363,N_12126,N_12146);
nor U12364 (N_12364,N_12154,N_12143);
nor U12365 (N_12365,N_12164,N_12241);
nor U12366 (N_12366,N_12226,N_12194);
nand U12367 (N_12367,N_12155,N_12178);
xor U12368 (N_12368,N_12173,N_12199);
or U12369 (N_12369,N_12212,N_12222);
or U12370 (N_12370,N_12170,N_12150);
xnor U12371 (N_12371,N_12216,N_12137);
or U12372 (N_12372,N_12126,N_12130);
or U12373 (N_12373,N_12170,N_12148);
nor U12374 (N_12374,N_12152,N_12239);
xor U12375 (N_12375,N_12305,N_12276);
nand U12376 (N_12376,N_12313,N_12366);
and U12377 (N_12377,N_12250,N_12288);
nor U12378 (N_12378,N_12298,N_12311);
nor U12379 (N_12379,N_12279,N_12343);
and U12380 (N_12380,N_12331,N_12261);
nand U12381 (N_12381,N_12360,N_12334);
and U12382 (N_12382,N_12340,N_12365);
and U12383 (N_12383,N_12287,N_12253);
and U12384 (N_12384,N_12310,N_12282);
nor U12385 (N_12385,N_12319,N_12280);
xor U12386 (N_12386,N_12351,N_12352);
nor U12387 (N_12387,N_12344,N_12339);
nor U12388 (N_12388,N_12369,N_12306);
nor U12389 (N_12389,N_12347,N_12284);
nand U12390 (N_12390,N_12266,N_12314);
nor U12391 (N_12391,N_12309,N_12254);
nand U12392 (N_12392,N_12286,N_12257);
xor U12393 (N_12393,N_12350,N_12324);
xnor U12394 (N_12394,N_12322,N_12269);
and U12395 (N_12395,N_12353,N_12291);
nand U12396 (N_12396,N_12283,N_12275);
and U12397 (N_12397,N_12321,N_12373);
xor U12398 (N_12398,N_12255,N_12308);
and U12399 (N_12399,N_12290,N_12312);
nor U12400 (N_12400,N_12357,N_12317);
xnor U12401 (N_12401,N_12271,N_12333);
or U12402 (N_12402,N_12364,N_12278);
and U12403 (N_12403,N_12328,N_12337);
and U12404 (N_12404,N_12281,N_12295);
xnor U12405 (N_12405,N_12267,N_12318);
xor U12406 (N_12406,N_12263,N_12374);
nor U12407 (N_12407,N_12265,N_12341);
xnor U12408 (N_12408,N_12358,N_12260);
and U12409 (N_12409,N_12277,N_12329);
nor U12410 (N_12410,N_12330,N_12348);
and U12411 (N_12411,N_12345,N_12355);
nor U12412 (N_12412,N_12259,N_12300);
xnor U12413 (N_12413,N_12307,N_12264);
nor U12414 (N_12414,N_12285,N_12299);
nor U12415 (N_12415,N_12293,N_12258);
xnor U12416 (N_12416,N_12272,N_12297);
nand U12417 (N_12417,N_12371,N_12372);
xnor U12418 (N_12418,N_12289,N_12303);
and U12419 (N_12419,N_12294,N_12320);
and U12420 (N_12420,N_12323,N_12354);
and U12421 (N_12421,N_12302,N_12251);
nor U12422 (N_12422,N_12359,N_12367);
xor U12423 (N_12423,N_12262,N_12292);
and U12424 (N_12424,N_12368,N_12346);
nand U12425 (N_12425,N_12332,N_12335);
and U12426 (N_12426,N_12342,N_12296);
and U12427 (N_12427,N_12304,N_12326);
nor U12428 (N_12428,N_12316,N_12270);
or U12429 (N_12429,N_12252,N_12361);
nor U12430 (N_12430,N_12336,N_12370);
xnor U12431 (N_12431,N_12268,N_12301);
and U12432 (N_12432,N_12327,N_12356);
nor U12433 (N_12433,N_12273,N_12362);
nor U12434 (N_12434,N_12349,N_12256);
nor U12435 (N_12435,N_12274,N_12325);
nand U12436 (N_12436,N_12363,N_12315);
or U12437 (N_12437,N_12338,N_12281);
or U12438 (N_12438,N_12261,N_12255);
or U12439 (N_12439,N_12368,N_12369);
nand U12440 (N_12440,N_12260,N_12301);
and U12441 (N_12441,N_12319,N_12342);
nand U12442 (N_12442,N_12335,N_12360);
xor U12443 (N_12443,N_12267,N_12336);
nor U12444 (N_12444,N_12365,N_12321);
nand U12445 (N_12445,N_12284,N_12279);
or U12446 (N_12446,N_12337,N_12343);
and U12447 (N_12447,N_12258,N_12275);
nor U12448 (N_12448,N_12367,N_12323);
nand U12449 (N_12449,N_12364,N_12253);
xor U12450 (N_12450,N_12333,N_12334);
xor U12451 (N_12451,N_12316,N_12339);
nand U12452 (N_12452,N_12285,N_12365);
nand U12453 (N_12453,N_12309,N_12322);
nand U12454 (N_12454,N_12285,N_12280);
or U12455 (N_12455,N_12331,N_12338);
nand U12456 (N_12456,N_12259,N_12270);
xnor U12457 (N_12457,N_12256,N_12260);
and U12458 (N_12458,N_12282,N_12300);
xor U12459 (N_12459,N_12273,N_12292);
and U12460 (N_12460,N_12357,N_12312);
or U12461 (N_12461,N_12373,N_12356);
nor U12462 (N_12462,N_12309,N_12330);
nand U12463 (N_12463,N_12290,N_12314);
and U12464 (N_12464,N_12294,N_12290);
xnor U12465 (N_12465,N_12264,N_12319);
nor U12466 (N_12466,N_12321,N_12334);
xor U12467 (N_12467,N_12342,N_12282);
nand U12468 (N_12468,N_12263,N_12268);
and U12469 (N_12469,N_12264,N_12337);
or U12470 (N_12470,N_12302,N_12271);
nand U12471 (N_12471,N_12251,N_12267);
and U12472 (N_12472,N_12314,N_12278);
xor U12473 (N_12473,N_12348,N_12288);
nor U12474 (N_12474,N_12277,N_12350);
or U12475 (N_12475,N_12290,N_12252);
or U12476 (N_12476,N_12252,N_12272);
or U12477 (N_12477,N_12311,N_12328);
xor U12478 (N_12478,N_12292,N_12316);
xnor U12479 (N_12479,N_12299,N_12254);
xor U12480 (N_12480,N_12275,N_12254);
and U12481 (N_12481,N_12351,N_12301);
or U12482 (N_12482,N_12290,N_12289);
or U12483 (N_12483,N_12286,N_12370);
and U12484 (N_12484,N_12263,N_12300);
xor U12485 (N_12485,N_12311,N_12340);
nor U12486 (N_12486,N_12329,N_12335);
nor U12487 (N_12487,N_12252,N_12344);
xnor U12488 (N_12488,N_12326,N_12364);
xnor U12489 (N_12489,N_12368,N_12268);
xnor U12490 (N_12490,N_12356,N_12265);
xor U12491 (N_12491,N_12295,N_12307);
or U12492 (N_12492,N_12360,N_12343);
xor U12493 (N_12493,N_12259,N_12299);
or U12494 (N_12494,N_12326,N_12316);
nand U12495 (N_12495,N_12294,N_12373);
or U12496 (N_12496,N_12295,N_12372);
nor U12497 (N_12497,N_12260,N_12278);
or U12498 (N_12498,N_12338,N_12265);
nand U12499 (N_12499,N_12257,N_12260);
nand U12500 (N_12500,N_12447,N_12410);
xor U12501 (N_12501,N_12430,N_12412);
xor U12502 (N_12502,N_12448,N_12418);
or U12503 (N_12503,N_12454,N_12428);
nor U12504 (N_12504,N_12484,N_12432);
xor U12505 (N_12505,N_12473,N_12439);
and U12506 (N_12506,N_12396,N_12438);
or U12507 (N_12507,N_12393,N_12476);
or U12508 (N_12508,N_12463,N_12490);
and U12509 (N_12509,N_12485,N_12383);
and U12510 (N_12510,N_12386,N_12458);
and U12511 (N_12511,N_12422,N_12480);
nor U12512 (N_12512,N_12378,N_12414);
or U12513 (N_12513,N_12379,N_12468);
xnor U12514 (N_12514,N_12382,N_12376);
nor U12515 (N_12515,N_12459,N_12391);
xor U12516 (N_12516,N_12472,N_12498);
nand U12517 (N_12517,N_12471,N_12395);
or U12518 (N_12518,N_12429,N_12478);
and U12519 (N_12519,N_12402,N_12403);
and U12520 (N_12520,N_12392,N_12408);
nand U12521 (N_12521,N_12488,N_12474);
nand U12522 (N_12522,N_12457,N_12416);
or U12523 (N_12523,N_12375,N_12420);
xnor U12524 (N_12524,N_12495,N_12437);
xnor U12525 (N_12525,N_12445,N_12435);
nor U12526 (N_12526,N_12387,N_12426);
xor U12527 (N_12527,N_12441,N_12423);
xor U12528 (N_12528,N_12405,N_12398);
nand U12529 (N_12529,N_12464,N_12433);
nand U12530 (N_12530,N_12483,N_12467);
or U12531 (N_12531,N_12466,N_12446);
or U12532 (N_12532,N_12440,N_12499);
or U12533 (N_12533,N_12479,N_12452);
nand U12534 (N_12534,N_12453,N_12406);
or U12535 (N_12535,N_12431,N_12489);
nor U12536 (N_12536,N_12424,N_12427);
or U12537 (N_12537,N_12462,N_12425);
nor U12538 (N_12538,N_12384,N_12497);
and U12539 (N_12539,N_12401,N_12477);
nand U12540 (N_12540,N_12450,N_12496);
or U12541 (N_12541,N_12409,N_12492);
or U12542 (N_12542,N_12436,N_12443);
nand U12543 (N_12543,N_12461,N_12460);
nand U12544 (N_12544,N_12482,N_12469);
or U12545 (N_12545,N_12442,N_12465);
xnor U12546 (N_12546,N_12470,N_12417);
nand U12547 (N_12547,N_12397,N_12377);
or U12548 (N_12548,N_12444,N_12455);
xor U12549 (N_12549,N_12421,N_12413);
xor U12550 (N_12550,N_12381,N_12388);
nor U12551 (N_12551,N_12451,N_12487);
and U12552 (N_12552,N_12411,N_12380);
or U12553 (N_12553,N_12456,N_12399);
and U12554 (N_12554,N_12400,N_12494);
nor U12555 (N_12555,N_12407,N_12434);
or U12556 (N_12556,N_12449,N_12475);
or U12557 (N_12557,N_12389,N_12481);
xor U12558 (N_12558,N_12404,N_12390);
nand U12559 (N_12559,N_12493,N_12415);
xnor U12560 (N_12560,N_12419,N_12491);
xnor U12561 (N_12561,N_12486,N_12385);
nor U12562 (N_12562,N_12394,N_12478);
nor U12563 (N_12563,N_12446,N_12395);
nand U12564 (N_12564,N_12447,N_12469);
and U12565 (N_12565,N_12433,N_12481);
nor U12566 (N_12566,N_12457,N_12449);
and U12567 (N_12567,N_12442,N_12496);
nor U12568 (N_12568,N_12396,N_12408);
xor U12569 (N_12569,N_12415,N_12385);
xor U12570 (N_12570,N_12394,N_12439);
xnor U12571 (N_12571,N_12404,N_12463);
nand U12572 (N_12572,N_12486,N_12490);
nand U12573 (N_12573,N_12418,N_12460);
nand U12574 (N_12574,N_12448,N_12410);
xor U12575 (N_12575,N_12423,N_12394);
nor U12576 (N_12576,N_12483,N_12459);
xnor U12577 (N_12577,N_12473,N_12454);
or U12578 (N_12578,N_12461,N_12458);
nand U12579 (N_12579,N_12476,N_12493);
nor U12580 (N_12580,N_12478,N_12413);
xor U12581 (N_12581,N_12458,N_12411);
xor U12582 (N_12582,N_12443,N_12398);
and U12583 (N_12583,N_12455,N_12463);
or U12584 (N_12584,N_12493,N_12392);
nor U12585 (N_12585,N_12424,N_12436);
xnor U12586 (N_12586,N_12473,N_12470);
nand U12587 (N_12587,N_12426,N_12381);
and U12588 (N_12588,N_12407,N_12450);
and U12589 (N_12589,N_12418,N_12496);
and U12590 (N_12590,N_12496,N_12396);
and U12591 (N_12591,N_12416,N_12410);
and U12592 (N_12592,N_12419,N_12437);
nor U12593 (N_12593,N_12468,N_12395);
and U12594 (N_12594,N_12391,N_12414);
nand U12595 (N_12595,N_12464,N_12434);
and U12596 (N_12596,N_12443,N_12429);
or U12597 (N_12597,N_12438,N_12430);
and U12598 (N_12598,N_12481,N_12482);
or U12599 (N_12599,N_12458,N_12415);
nor U12600 (N_12600,N_12483,N_12463);
xor U12601 (N_12601,N_12383,N_12394);
and U12602 (N_12602,N_12441,N_12389);
or U12603 (N_12603,N_12480,N_12451);
nand U12604 (N_12604,N_12428,N_12423);
nand U12605 (N_12605,N_12457,N_12479);
nor U12606 (N_12606,N_12435,N_12441);
xor U12607 (N_12607,N_12490,N_12394);
and U12608 (N_12608,N_12443,N_12392);
nor U12609 (N_12609,N_12401,N_12437);
xnor U12610 (N_12610,N_12447,N_12401);
nand U12611 (N_12611,N_12417,N_12492);
xnor U12612 (N_12612,N_12479,N_12404);
xor U12613 (N_12613,N_12432,N_12443);
or U12614 (N_12614,N_12444,N_12394);
and U12615 (N_12615,N_12418,N_12489);
xor U12616 (N_12616,N_12377,N_12444);
nand U12617 (N_12617,N_12477,N_12379);
or U12618 (N_12618,N_12443,N_12394);
xor U12619 (N_12619,N_12474,N_12489);
nor U12620 (N_12620,N_12499,N_12405);
nor U12621 (N_12621,N_12447,N_12419);
and U12622 (N_12622,N_12418,N_12422);
nor U12623 (N_12623,N_12464,N_12426);
nor U12624 (N_12624,N_12443,N_12471);
and U12625 (N_12625,N_12593,N_12609);
nand U12626 (N_12626,N_12574,N_12567);
nor U12627 (N_12627,N_12605,N_12542);
and U12628 (N_12628,N_12581,N_12559);
nor U12629 (N_12629,N_12508,N_12513);
nand U12630 (N_12630,N_12604,N_12509);
xnor U12631 (N_12631,N_12622,N_12552);
nand U12632 (N_12632,N_12511,N_12590);
nand U12633 (N_12633,N_12502,N_12585);
and U12634 (N_12634,N_12596,N_12527);
and U12635 (N_12635,N_12594,N_12578);
nand U12636 (N_12636,N_12565,N_12560);
nor U12637 (N_12637,N_12541,N_12617);
and U12638 (N_12638,N_12548,N_12606);
and U12639 (N_12639,N_12603,N_12523);
or U12640 (N_12640,N_12558,N_12612);
or U12641 (N_12641,N_12517,N_12607);
xnor U12642 (N_12642,N_12529,N_12564);
nor U12643 (N_12643,N_12544,N_12610);
or U12644 (N_12644,N_12507,N_12501);
nor U12645 (N_12645,N_12537,N_12549);
xnor U12646 (N_12646,N_12561,N_12533);
and U12647 (N_12647,N_12528,N_12599);
nand U12648 (N_12648,N_12583,N_12600);
nor U12649 (N_12649,N_12525,N_12614);
xnor U12650 (N_12650,N_12536,N_12582);
and U12651 (N_12651,N_12589,N_12597);
and U12652 (N_12652,N_12505,N_12521);
and U12653 (N_12653,N_12503,N_12515);
nand U12654 (N_12654,N_12551,N_12563);
or U12655 (N_12655,N_12504,N_12598);
or U12656 (N_12656,N_12516,N_12601);
nand U12657 (N_12657,N_12530,N_12579);
and U12658 (N_12658,N_12514,N_12569);
xnor U12659 (N_12659,N_12512,N_12571);
nand U12660 (N_12660,N_12587,N_12539);
and U12661 (N_12661,N_12608,N_12538);
and U12662 (N_12662,N_12577,N_12510);
xor U12663 (N_12663,N_12506,N_12613);
or U12664 (N_12664,N_12588,N_12531);
or U12665 (N_12665,N_12621,N_12500);
xnor U12666 (N_12666,N_12592,N_12572);
xnor U12667 (N_12667,N_12553,N_12618);
and U12668 (N_12668,N_12620,N_12543);
nor U12669 (N_12669,N_12557,N_12573);
xor U12670 (N_12670,N_12535,N_12550);
and U12671 (N_12671,N_12580,N_12562);
or U12672 (N_12672,N_12570,N_12545);
xor U12673 (N_12673,N_12595,N_12611);
nor U12674 (N_12674,N_12584,N_12555);
and U12675 (N_12675,N_12524,N_12616);
xor U12676 (N_12676,N_12519,N_12566);
nand U12677 (N_12677,N_12540,N_12619);
nor U12678 (N_12678,N_12586,N_12575);
or U12679 (N_12679,N_12554,N_12522);
and U12680 (N_12680,N_12623,N_12546);
nand U12681 (N_12681,N_12624,N_12547);
and U12682 (N_12682,N_12526,N_12568);
nand U12683 (N_12683,N_12556,N_12532);
nand U12684 (N_12684,N_12534,N_12518);
and U12685 (N_12685,N_12615,N_12576);
xnor U12686 (N_12686,N_12591,N_12520);
and U12687 (N_12687,N_12602,N_12606);
nand U12688 (N_12688,N_12542,N_12561);
xnor U12689 (N_12689,N_12613,N_12532);
and U12690 (N_12690,N_12516,N_12590);
xor U12691 (N_12691,N_12528,N_12504);
nor U12692 (N_12692,N_12577,N_12505);
xnor U12693 (N_12693,N_12596,N_12616);
or U12694 (N_12694,N_12554,N_12569);
xor U12695 (N_12695,N_12507,N_12562);
xor U12696 (N_12696,N_12536,N_12624);
or U12697 (N_12697,N_12522,N_12619);
nand U12698 (N_12698,N_12598,N_12550);
nand U12699 (N_12699,N_12501,N_12539);
or U12700 (N_12700,N_12547,N_12621);
nand U12701 (N_12701,N_12519,N_12583);
xnor U12702 (N_12702,N_12568,N_12519);
or U12703 (N_12703,N_12542,N_12614);
nor U12704 (N_12704,N_12549,N_12587);
nor U12705 (N_12705,N_12527,N_12520);
and U12706 (N_12706,N_12518,N_12557);
nor U12707 (N_12707,N_12604,N_12612);
and U12708 (N_12708,N_12559,N_12549);
nor U12709 (N_12709,N_12590,N_12533);
nor U12710 (N_12710,N_12522,N_12556);
xnor U12711 (N_12711,N_12553,N_12595);
or U12712 (N_12712,N_12506,N_12602);
xor U12713 (N_12713,N_12541,N_12538);
xnor U12714 (N_12714,N_12507,N_12540);
nand U12715 (N_12715,N_12622,N_12536);
or U12716 (N_12716,N_12601,N_12604);
nor U12717 (N_12717,N_12599,N_12566);
nand U12718 (N_12718,N_12503,N_12567);
or U12719 (N_12719,N_12583,N_12534);
nor U12720 (N_12720,N_12507,N_12531);
xor U12721 (N_12721,N_12579,N_12613);
nor U12722 (N_12722,N_12594,N_12611);
nand U12723 (N_12723,N_12598,N_12558);
xnor U12724 (N_12724,N_12519,N_12523);
nand U12725 (N_12725,N_12572,N_12589);
and U12726 (N_12726,N_12603,N_12560);
xor U12727 (N_12727,N_12608,N_12549);
xnor U12728 (N_12728,N_12503,N_12574);
or U12729 (N_12729,N_12524,N_12559);
or U12730 (N_12730,N_12527,N_12592);
xor U12731 (N_12731,N_12504,N_12547);
xnor U12732 (N_12732,N_12590,N_12588);
nand U12733 (N_12733,N_12500,N_12617);
and U12734 (N_12734,N_12605,N_12611);
xnor U12735 (N_12735,N_12534,N_12598);
nor U12736 (N_12736,N_12588,N_12571);
or U12737 (N_12737,N_12555,N_12624);
nor U12738 (N_12738,N_12548,N_12509);
or U12739 (N_12739,N_12543,N_12539);
or U12740 (N_12740,N_12565,N_12527);
nor U12741 (N_12741,N_12550,N_12595);
xnor U12742 (N_12742,N_12558,N_12501);
or U12743 (N_12743,N_12606,N_12560);
or U12744 (N_12744,N_12559,N_12598);
xnor U12745 (N_12745,N_12513,N_12515);
xor U12746 (N_12746,N_12608,N_12529);
nand U12747 (N_12747,N_12575,N_12587);
nand U12748 (N_12748,N_12556,N_12577);
nand U12749 (N_12749,N_12614,N_12555);
xor U12750 (N_12750,N_12734,N_12736);
and U12751 (N_12751,N_12724,N_12689);
nand U12752 (N_12752,N_12728,N_12729);
and U12753 (N_12753,N_12672,N_12662);
or U12754 (N_12754,N_12705,N_12687);
or U12755 (N_12755,N_12680,N_12716);
and U12756 (N_12756,N_12715,N_12733);
nor U12757 (N_12757,N_12629,N_12703);
or U12758 (N_12758,N_12747,N_12684);
xnor U12759 (N_12759,N_12735,N_12657);
nand U12760 (N_12760,N_12661,N_12732);
or U12761 (N_12761,N_12633,N_12706);
nor U12762 (N_12762,N_12685,N_12659);
and U12763 (N_12763,N_12656,N_12737);
nand U12764 (N_12764,N_12713,N_12683);
or U12765 (N_12765,N_12696,N_12697);
nor U12766 (N_12766,N_12677,N_12653);
xnor U12767 (N_12767,N_12693,N_12692);
or U12768 (N_12768,N_12695,N_12627);
nand U12769 (N_12769,N_12675,N_12634);
nor U12770 (N_12770,N_12682,N_12690);
and U12771 (N_12771,N_12708,N_12730);
or U12772 (N_12772,N_12666,N_12643);
and U12773 (N_12773,N_12649,N_12671);
xnor U12774 (N_12774,N_12707,N_12714);
and U12775 (N_12775,N_12731,N_12678);
nor U12776 (N_12776,N_12668,N_12748);
nand U12777 (N_12777,N_12632,N_12630);
and U12778 (N_12778,N_12717,N_12628);
xnor U12779 (N_12779,N_12647,N_12741);
and U12780 (N_12780,N_12694,N_12646);
or U12781 (N_12781,N_12669,N_12652);
nand U12782 (N_12782,N_12740,N_12704);
xnor U12783 (N_12783,N_12650,N_12654);
and U12784 (N_12784,N_12644,N_12641);
nand U12785 (N_12785,N_12681,N_12636);
or U12786 (N_12786,N_12699,N_12660);
nand U12787 (N_12787,N_12665,N_12749);
nand U12788 (N_12788,N_12742,N_12664);
and U12789 (N_12789,N_12637,N_12727);
and U12790 (N_12790,N_12743,N_12723);
nand U12791 (N_12791,N_12702,N_12710);
nand U12792 (N_12792,N_12726,N_12712);
or U12793 (N_12793,N_12635,N_12711);
nor U12794 (N_12794,N_12739,N_12686);
and U12795 (N_12795,N_12709,N_12746);
nand U12796 (N_12796,N_12691,N_12700);
nor U12797 (N_12797,N_12722,N_12667);
nand U12798 (N_12798,N_12721,N_12701);
or U12799 (N_12799,N_12719,N_12655);
or U12800 (N_12800,N_12679,N_12745);
nand U12801 (N_12801,N_12663,N_12648);
or U12802 (N_12802,N_12698,N_12625);
or U12803 (N_12803,N_12626,N_12744);
nand U12804 (N_12804,N_12658,N_12688);
xnor U12805 (N_12805,N_12640,N_12720);
nor U12806 (N_12806,N_12725,N_12676);
nand U12807 (N_12807,N_12638,N_12718);
xnor U12808 (N_12808,N_12639,N_12673);
nand U12809 (N_12809,N_12674,N_12631);
xor U12810 (N_12810,N_12642,N_12645);
and U12811 (N_12811,N_12670,N_12651);
nand U12812 (N_12812,N_12738,N_12646);
xor U12813 (N_12813,N_12640,N_12748);
xor U12814 (N_12814,N_12745,N_12663);
nor U12815 (N_12815,N_12742,N_12703);
xnor U12816 (N_12816,N_12627,N_12663);
or U12817 (N_12817,N_12695,N_12733);
nand U12818 (N_12818,N_12649,N_12740);
or U12819 (N_12819,N_12649,N_12673);
and U12820 (N_12820,N_12677,N_12701);
nor U12821 (N_12821,N_12658,N_12717);
nor U12822 (N_12822,N_12686,N_12725);
nand U12823 (N_12823,N_12673,N_12725);
or U12824 (N_12824,N_12721,N_12667);
nor U12825 (N_12825,N_12741,N_12712);
and U12826 (N_12826,N_12714,N_12671);
xnor U12827 (N_12827,N_12745,N_12630);
nand U12828 (N_12828,N_12701,N_12685);
and U12829 (N_12829,N_12658,N_12715);
or U12830 (N_12830,N_12648,N_12717);
nor U12831 (N_12831,N_12680,N_12630);
xnor U12832 (N_12832,N_12677,N_12652);
nor U12833 (N_12833,N_12711,N_12668);
and U12834 (N_12834,N_12725,N_12695);
or U12835 (N_12835,N_12692,N_12641);
nand U12836 (N_12836,N_12733,N_12673);
xor U12837 (N_12837,N_12730,N_12686);
nand U12838 (N_12838,N_12746,N_12686);
xnor U12839 (N_12839,N_12667,N_12707);
nand U12840 (N_12840,N_12712,N_12661);
and U12841 (N_12841,N_12684,N_12730);
nor U12842 (N_12842,N_12672,N_12728);
nor U12843 (N_12843,N_12720,N_12694);
nor U12844 (N_12844,N_12667,N_12626);
xnor U12845 (N_12845,N_12679,N_12732);
nor U12846 (N_12846,N_12673,N_12729);
nand U12847 (N_12847,N_12695,N_12683);
nand U12848 (N_12848,N_12696,N_12674);
and U12849 (N_12849,N_12720,N_12716);
and U12850 (N_12850,N_12638,N_12653);
nand U12851 (N_12851,N_12653,N_12676);
or U12852 (N_12852,N_12694,N_12740);
nor U12853 (N_12853,N_12626,N_12695);
nor U12854 (N_12854,N_12660,N_12698);
xor U12855 (N_12855,N_12688,N_12645);
nand U12856 (N_12856,N_12684,N_12661);
and U12857 (N_12857,N_12714,N_12650);
nand U12858 (N_12858,N_12698,N_12735);
xor U12859 (N_12859,N_12671,N_12730);
or U12860 (N_12860,N_12729,N_12627);
or U12861 (N_12861,N_12680,N_12652);
or U12862 (N_12862,N_12670,N_12701);
nor U12863 (N_12863,N_12680,N_12725);
xnor U12864 (N_12864,N_12625,N_12711);
nor U12865 (N_12865,N_12719,N_12727);
nor U12866 (N_12866,N_12701,N_12659);
nor U12867 (N_12867,N_12738,N_12718);
and U12868 (N_12868,N_12748,N_12636);
nor U12869 (N_12869,N_12627,N_12740);
nor U12870 (N_12870,N_12723,N_12744);
xnor U12871 (N_12871,N_12662,N_12684);
and U12872 (N_12872,N_12718,N_12654);
nor U12873 (N_12873,N_12669,N_12707);
nor U12874 (N_12874,N_12720,N_12691);
nor U12875 (N_12875,N_12772,N_12804);
xor U12876 (N_12876,N_12849,N_12788);
and U12877 (N_12877,N_12858,N_12817);
or U12878 (N_12878,N_12783,N_12866);
or U12879 (N_12879,N_12800,N_12865);
nor U12880 (N_12880,N_12765,N_12854);
xor U12881 (N_12881,N_12845,N_12853);
nor U12882 (N_12882,N_12777,N_12795);
nand U12883 (N_12883,N_12776,N_12870);
nor U12884 (N_12884,N_12869,N_12806);
or U12885 (N_12885,N_12770,N_12771);
nor U12886 (N_12886,N_12864,N_12852);
and U12887 (N_12887,N_12827,N_12822);
xnor U12888 (N_12888,N_12818,N_12820);
nand U12889 (N_12889,N_12829,N_12833);
or U12890 (N_12890,N_12764,N_12802);
xnor U12891 (N_12891,N_12782,N_12803);
nor U12892 (N_12892,N_12757,N_12848);
xnor U12893 (N_12893,N_12775,N_12767);
and U12894 (N_12894,N_12758,N_12756);
and U12895 (N_12895,N_12808,N_12796);
and U12896 (N_12896,N_12840,N_12786);
nor U12897 (N_12897,N_12787,N_12768);
nor U12898 (N_12898,N_12752,N_12760);
xor U12899 (N_12899,N_12762,N_12813);
nand U12900 (N_12900,N_12792,N_12780);
or U12901 (N_12901,N_12801,N_12798);
nand U12902 (N_12902,N_12789,N_12834);
xnor U12903 (N_12903,N_12794,N_12831);
nor U12904 (N_12904,N_12812,N_12807);
xor U12905 (N_12905,N_12826,N_12846);
nor U12906 (N_12906,N_12781,N_12830);
or U12907 (N_12907,N_12868,N_12797);
and U12908 (N_12908,N_12815,N_12816);
xnor U12909 (N_12909,N_12860,N_12809);
nor U12910 (N_12910,N_12751,N_12824);
xnor U12911 (N_12911,N_12773,N_12839);
xnor U12912 (N_12912,N_12754,N_12874);
xnor U12913 (N_12913,N_12763,N_12872);
or U12914 (N_12914,N_12810,N_12766);
or U12915 (N_12915,N_12842,N_12837);
nor U12916 (N_12916,N_12863,N_12873);
nor U12917 (N_12917,N_12841,N_12814);
xnor U12918 (N_12918,N_12753,N_12750);
nor U12919 (N_12919,N_12805,N_12862);
and U12920 (N_12920,N_12851,N_12867);
nor U12921 (N_12921,N_12850,N_12779);
nor U12922 (N_12922,N_12784,N_12769);
xnor U12923 (N_12923,N_12755,N_12857);
and U12924 (N_12924,N_12856,N_12871);
nor U12925 (N_12925,N_12832,N_12861);
xnor U12926 (N_12926,N_12759,N_12843);
and U12927 (N_12927,N_12828,N_12859);
nor U12928 (N_12928,N_12821,N_12823);
or U12929 (N_12929,N_12844,N_12790);
nor U12930 (N_12930,N_12836,N_12835);
and U12931 (N_12931,N_12774,N_12838);
or U12932 (N_12932,N_12799,N_12847);
nand U12933 (N_12933,N_12855,N_12793);
xor U12934 (N_12934,N_12791,N_12785);
and U12935 (N_12935,N_12819,N_12761);
nor U12936 (N_12936,N_12811,N_12778);
or U12937 (N_12937,N_12825,N_12801);
and U12938 (N_12938,N_12773,N_12813);
nor U12939 (N_12939,N_12816,N_12866);
nand U12940 (N_12940,N_12868,N_12840);
xor U12941 (N_12941,N_12758,N_12769);
xnor U12942 (N_12942,N_12857,N_12816);
or U12943 (N_12943,N_12798,N_12800);
and U12944 (N_12944,N_12791,N_12810);
nor U12945 (N_12945,N_12783,N_12789);
nor U12946 (N_12946,N_12845,N_12824);
nand U12947 (N_12947,N_12790,N_12865);
xor U12948 (N_12948,N_12764,N_12808);
nand U12949 (N_12949,N_12773,N_12769);
nand U12950 (N_12950,N_12765,N_12860);
xor U12951 (N_12951,N_12861,N_12803);
nor U12952 (N_12952,N_12797,N_12829);
and U12953 (N_12953,N_12773,N_12823);
and U12954 (N_12954,N_12842,N_12858);
nand U12955 (N_12955,N_12814,N_12840);
or U12956 (N_12956,N_12788,N_12818);
and U12957 (N_12957,N_12832,N_12797);
xor U12958 (N_12958,N_12871,N_12817);
or U12959 (N_12959,N_12782,N_12827);
xnor U12960 (N_12960,N_12767,N_12799);
nor U12961 (N_12961,N_12858,N_12762);
or U12962 (N_12962,N_12871,N_12836);
nor U12963 (N_12963,N_12837,N_12839);
or U12964 (N_12964,N_12827,N_12856);
or U12965 (N_12965,N_12872,N_12779);
or U12966 (N_12966,N_12808,N_12771);
xor U12967 (N_12967,N_12861,N_12840);
xor U12968 (N_12968,N_12835,N_12764);
xor U12969 (N_12969,N_12766,N_12840);
xnor U12970 (N_12970,N_12769,N_12803);
and U12971 (N_12971,N_12785,N_12834);
or U12972 (N_12972,N_12810,N_12780);
nor U12973 (N_12973,N_12801,N_12827);
nor U12974 (N_12974,N_12791,N_12861);
nor U12975 (N_12975,N_12755,N_12817);
and U12976 (N_12976,N_12874,N_12857);
xnor U12977 (N_12977,N_12850,N_12782);
nor U12978 (N_12978,N_12831,N_12865);
and U12979 (N_12979,N_12854,N_12818);
xnor U12980 (N_12980,N_12862,N_12768);
xor U12981 (N_12981,N_12752,N_12825);
nand U12982 (N_12982,N_12833,N_12843);
nand U12983 (N_12983,N_12780,N_12837);
or U12984 (N_12984,N_12855,N_12803);
nor U12985 (N_12985,N_12794,N_12795);
or U12986 (N_12986,N_12802,N_12864);
or U12987 (N_12987,N_12822,N_12776);
and U12988 (N_12988,N_12872,N_12825);
nand U12989 (N_12989,N_12797,N_12809);
xnor U12990 (N_12990,N_12869,N_12778);
nand U12991 (N_12991,N_12809,N_12785);
nand U12992 (N_12992,N_12874,N_12838);
xor U12993 (N_12993,N_12810,N_12812);
nor U12994 (N_12994,N_12867,N_12753);
or U12995 (N_12995,N_12822,N_12809);
and U12996 (N_12996,N_12834,N_12782);
or U12997 (N_12997,N_12847,N_12873);
and U12998 (N_12998,N_12836,N_12850);
nor U12999 (N_12999,N_12812,N_12860);
nor U13000 (N_13000,N_12948,N_12884);
and U13001 (N_13001,N_12999,N_12984);
and U13002 (N_13002,N_12977,N_12877);
xnor U13003 (N_13003,N_12940,N_12972);
xnor U13004 (N_13004,N_12934,N_12979);
nand U13005 (N_13005,N_12880,N_12971);
nand U13006 (N_13006,N_12896,N_12911);
or U13007 (N_13007,N_12997,N_12891);
or U13008 (N_13008,N_12969,N_12919);
nand U13009 (N_13009,N_12962,N_12909);
nand U13010 (N_13010,N_12956,N_12889);
nor U13011 (N_13011,N_12927,N_12907);
or U13012 (N_13012,N_12921,N_12903);
and U13013 (N_13013,N_12916,N_12967);
or U13014 (N_13014,N_12937,N_12964);
xnor U13015 (N_13015,N_12996,N_12938);
and U13016 (N_13016,N_12876,N_12883);
nand U13017 (N_13017,N_12914,N_12913);
or U13018 (N_13018,N_12924,N_12894);
xnor U13019 (N_13019,N_12970,N_12881);
nor U13020 (N_13020,N_12885,N_12987);
nand U13021 (N_13021,N_12928,N_12974);
nor U13022 (N_13022,N_12993,N_12922);
xor U13023 (N_13023,N_12912,N_12918);
or U13024 (N_13024,N_12910,N_12930);
nor U13025 (N_13025,N_12958,N_12886);
xnor U13026 (N_13026,N_12933,N_12989);
nand U13027 (N_13027,N_12892,N_12920);
nand U13028 (N_13028,N_12900,N_12925);
nor U13029 (N_13029,N_12961,N_12953);
and U13030 (N_13030,N_12973,N_12943);
nand U13031 (N_13031,N_12990,N_12992);
xor U13032 (N_13032,N_12917,N_12942);
nand U13033 (N_13033,N_12965,N_12890);
nor U13034 (N_13034,N_12939,N_12986);
and U13035 (N_13035,N_12879,N_12976);
nand U13036 (N_13036,N_12905,N_12949);
nor U13037 (N_13037,N_12915,N_12945);
nor U13038 (N_13038,N_12955,N_12929);
or U13039 (N_13039,N_12982,N_12931);
and U13040 (N_13040,N_12946,N_12935);
nor U13041 (N_13041,N_12926,N_12954);
nor U13042 (N_13042,N_12947,N_12959);
or U13043 (N_13043,N_12998,N_12980);
nand U13044 (N_13044,N_12897,N_12963);
or U13045 (N_13045,N_12951,N_12991);
nand U13046 (N_13046,N_12878,N_12944);
and U13047 (N_13047,N_12904,N_12975);
xnor U13048 (N_13048,N_12985,N_12950);
nor U13049 (N_13049,N_12952,N_12901);
nor U13050 (N_13050,N_12899,N_12902);
and U13051 (N_13051,N_12906,N_12966);
or U13052 (N_13052,N_12875,N_12968);
nand U13053 (N_13053,N_12908,N_12898);
nor U13054 (N_13054,N_12895,N_12932);
xor U13055 (N_13055,N_12941,N_12995);
xnor U13056 (N_13056,N_12983,N_12893);
xor U13057 (N_13057,N_12887,N_12994);
or U13058 (N_13058,N_12888,N_12957);
or U13059 (N_13059,N_12936,N_12978);
or U13060 (N_13060,N_12960,N_12882);
or U13061 (N_13061,N_12988,N_12923);
or U13062 (N_13062,N_12981,N_12994);
xnor U13063 (N_13063,N_12984,N_12954);
nor U13064 (N_13064,N_12981,N_12889);
nor U13065 (N_13065,N_12882,N_12964);
and U13066 (N_13066,N_12880,N_12994);
xnor U13067 (N_13067,N_12903,N_12993);
and U13068 (N_13068,N_12908,N_12930);
nor U13069 (N_13069,N_12972,N_12992);
and U13070 (N_13070,N_12992,N_12947);
nand U13071 (N_13071,N_12898,N_12907);
nand U13072 (N_13072,N_12961,N_12999);
nand U13073 (N_13073,N_12917,N_12936);
nor U13074 (N_13074,N_12997,N_12881);
nor U13075 (N_13075,N_12970,N_12973);
and U13076 (N_13076,N_12985,N_12997);
or U13077 (N_13077,N_12916,N_12931);
xnor U13078 (N_13078,N_12948,N_12921);
or U13079 (N_13079,N_12926,N_12955);
xor U13080 (N_13080,N_12886,N_12960);
xor U13081 (N_13081,N_12971,N_12948);
or U13082 (N_13082,N_12971,N_12964);
and U13083 (N_13083,N_12966,N_12967);
nand U13084 (N_13084,N_12894,N_12965);
xnor U13085 (N_13085,N_12963,N_12910);
or U13086 (N_13086,N_12976,N_12959);
nand U13087 (N_13087,N_12916,N_12883);
and U13088 (N_13088,N_12894,N_12888);
xor U13089 (N_13089,N_12877,N_12962);
nand U13090 (N_13090,N_12962,N_12886);
or U13091 (N_13091,N_12942,N_12916);
nand U13092 (N_13092,N_12959,N_12966);
or U13093 (N_13093,N_12906,N_12936);
nand U13094 (N_13094,N_12991,N_12972);
xnor U13095 (N_13095,N_12969,N_12912);
nand U13096 (N_13096,N_12977,N_12886);
nor U13097 (N_13097,N_12877,N_12964);
xnor U13098 (N_13098,N_12892,N_12958);
xor U13099 (N_13099,N_12932,N_12995);
nor U13100 (N_13100,N_12888,N_12919);
and U13101 (N_13101,N_12881,N_12940);
or U13102 (N_13102,N_12966,N_12983);
xnor U13103 (N_13103,N_12963,N_12916);
or U13104 (N_13104,N_12956,N_12989);
nand U13105 (N_13105,N_12979,N_12886);
xnor U13106 (N_13106,N_12898,N_12901);
and U13107 (N_13107,N_12999,N_12957);
nor U13108 (N_13108,N_12942,N_12937);
nand U13109 (N_13109,N_12884,N_12920);
xor U13110 (N_13110,N_12956,N_12966);
nand U13111 (N_13111,N_12882,N_12899);
xor U13112 (N_13112,N_12960,N_12949);
xor U13113 (N_13113,N_12903,N_12988);
or U13114 (N_13114,N_12879,N_12973);
xnor U13115 (N_13115,N_12986,N_12926);
or U13116 (N_13116,N_12950,N_12930);
nand U13117 (N_13117,N_12993,N_12927);
nand U13118 (N_13118,N_12978,N_12966);
nand U13119 (N_13119,N_12993,N_12959);
xor U13120 (N_13120,N_12993,N_12995);
nor U13121 (N_13121,N_12999,N_12978);
xor U13122 (N_13122,N_12884,N_12984);
xnor U13123 (N_13123,N_12901,N_12959);
nand U13124 (N_13124,N_12884,N_12915);
or U13125 (N_13125,N_13035,N_13047);
and U13126 (N_13126,N_13083,N_13032);
nor U13127 (N_13127,N_13050,N_13055);
and U13128 (N_13128,N_13098,N_13054);
nand U13129 (N_13129,N_13096,N_13076);
xor U13130 (N_13130,N_13124,N_13013);
nor U13131 (N_13131,N_13010,N_13068);
nand U13132 (N_13132,N_13116,N_13052);
or U13133 (N_13133,N_13058,N_13106);
or U13134 (N_13134,N_13060,N_13049);
and U13135 (N_13135,N_13005,N_13003);
nor U13136 (N_13136,N_13123,N_13079);
nand U13137 (N_13137,N_13048,N_13030);
nand U13138 (N_13138,N_13109,N_13080);
and U13139 (N_13139,N_13007,N_13034);
nand U13140 (N_13140,N_13000,N_13008);
nor U13141 (N_13141,N_13094,N_13115);
nor U13142 (N_13142,N_13018,N_13072);
nor U13143 (N_13143,N_13037,N_13011);
nor U13144 (N_13144,N_13103,N_13053);
or U13145 (N_13145,N_13099,N_13121);
nand U13146 (N_13146,N_13042,N_13108);
xor U13147 (N_13147,N_13046,N_13090);
nand U13148 (N_13148,N_13095,N_13002);
and U13149 (N_13149,N_13012,N_13105);
and U13150 (N_13150,N_13069,N_13081);
xor U13151 (N_13151,N_13022,N_13017);
or U13152 (N_13152,N_13014,N_13088);
and U13153 (N_13153,N_13016,N_13062);
nand U13154 (N_13154,N_13006,N_13025);
or U13155 (N_13155,N_13019,N_13070);
or U13156 (N_13156,N_13015,N_13036);
xnor U13157 (N_13157,N_13112,N_13033);
and U13158 (N_13158,N_13078,N_13114);
nand U13159 (N_13159,N_13093,N_13028);
nor U13160 (N_13160,N_13041,N_13085);
and U13161 (N_13161,N_13092,N_13084);
or U13162 (N_13162,N_13021,N_13104);
and U13163 (N_13163,N_13059,N_13029);
xnor U13164 (N_13164,N_13040,N_13110);
nand U13165 (N_13165,N_13120,N_13009);
xnor U13166 (N_13166,N_13087,N_13119);
nand U13167 (N_13167,N_13097,N_13107);
or U13168 (N_13168,N_13073,N_13113);
xnor U13169 (N_13169,N_13086,N_13122);
or U13170 (N_13170,N_13024,N_13039);
nor U13171 (N_13171,N_13027,N_13082);
nand U13172 (N_13172,N_13067,N_13089);
xnor U13173 (N_13173,N_13066,N_13074);
and U13174 (N_13174,N_13004,N_13111);
and U13175 (N_13175,N_13101,N_13044);
nand U13176 (N_13176,N_13038,N_13075);
nor U13177 (N_13177,N_13057,N_13061);
nor U13178 (N_13178,N_13031,N_13001);
xnor U13179 (N_13179,N_13091,N_13118);
nand U13180 (N_13180,N_13020,N_13117);
or U13181 (N_13181,N_13100,N_13056);
xor U13182 (N_13182,N_13063,N_13023);
or U13183 (N_13183,N_13064,N_13026);
xnor U13184 (N_13184,N_13043,N_13102);
or U13185 (N_13185,N_13077,N_13051);
xnor U13186 (N_13186,N_13071,N_13045);
nand U13187 (N_13187,N_13065,N_13041);
xor U13188 (N_13188,N_13096,N_13099);
and U13189 (N_13189,N_13044,N_13072);
xor U13190 (N_13190,N_13096,N_13017);
or U13191 (N_13191,N_13119,N_13113);
xnor U13192 (N_13192,N_13074,N_13033);
and U13193 (N_13193,N_13064,N_13023);
xnor U13194 (N_13194,N_13063,N_13115);
and U13195 (N_13195,N_13029,N_13114);
xnor U13196 (N_13196,N_13028,N_13079);
nor U13197 (N_13197,N_13013,N_13091);
and U13198 (N_13198,N_13039,N_13032);
or U13199 (N_13199,N_13045,N_13102);
and U13200 (N_13200,N_13091,N_13109);
nor U13201 (N_13201,N_13024,N_13090);
nor U13202 (N_13202,N_13123,N_13067);
nor U13203 (N_13203,N_13041,N_13077);
nand U13204 (N_13204,N_13095,N_13010);
or U13205 (N_13205,N_13016,N_13093);
nand U13206 (N_13206,N_13047,N_13037);
and U13207 (N_13207,N_13071,N_13060);
or U13208 (N_13208,N_13077,N_13048);
nor U13209 (N_13209,N_13098,N_13084);
nor U13210 (N_13210,N_13005,N_13061);
nand U13211 (N_13211,N_13112,N_13019);
xnor U13212 (N_13212,N_13100,N_13028);
nand U13213 (N_13213,N_13009,N_13092);
nor U13214 (N_13214,N_13055,N_13037);
and U13215 (N_13215,N_13108,N_13058);
nand U13216 (N_13216,N_13033,N_13078);
and U13217 (N_13217,N_13029,N_13100);
or U13218 (N_13218,N_13098,N_13108);
and U13219 (N_13219,N_13107,N_13022);
and U13220 (N_13220,N_13102,N_13063);
nor U13221 (N_13221,N_13051,N_13074);
xor U13222 (N_13222,N_13020,N_13039);
nor U13223 (N_13223,N_13078,N_13064);
nand U13224 (N_13224,N_13079,N_13001);
and U13225 (N_13225,N_13081,N_13079);
nor U13226 (N_13226,N_13124,N_13104);
and U13227 (N_13227,N_13050,N_13003);
nor U13228 (N_13228,N_13107,N_13085);
nor U13229 (N_13229,N_13020,N_13075);
nor U13230 (N_13230,N_13123,N_13055);
or U13231 (N_13231,N_13075,N_13025);
nand U13232 (N_13232,N_13042,N_13121);
and U13233 (N_13233,N_13009,N_13101);
or U13234 (N_13234,N_13000,N_13078);
nand U13235 (N_13235,N_13054,N_13074);
and U13236 (N_13236,N_13050,N_13092);
and U13237 (N_13237,N_13061,N_13122);
and U13238 (N_13238,N_13112,N_13011);
xnor U13239 (N_13239,N_13033,N_13079);
or U13240 (N_13240,N_13006,N_13091);
or U13241 (N_13241,N_13001,N_13093);
xor U13242 (N_13242,N_13077,N_13018);
or U13243 (N_13243,N_13009,N_13121);
nor U13244 (N_13244,N_13084,N_13121);
nand U13245 (N_13245,N_13080,N_13121);
nand U13246 (N_13246,N_13100,N_13006);
or U13247 (N_13247,N_13028,N_13095);
and U13248 (N_13248,N_13034,N_13113);
or U13249 (N_13249,N_13095,N_13096);
nand U13250 (N_13250,N_13227,N_13198);
xnor U13251 (N_13251,N_13223,N_13245);
xor U13252 (N_13252,N_13215,N_13141);
and U13253 (N_13253,N_13193,N_13160);
xor U13254 (N_13254,N_13219,N_13211);
and U13255 (N_13255,N_13186,N_13133);
and U13256 (N_13256,N_13226,N_13145);
and U13257 (N_13257,N_13221,N_13137);
or U13258 (N_13258,N_13248,N_13178);
and U13259 (N_13259,N_13243,N_13242);
nand U13260 (N_13260,N_13154,N_13138);
nor U13261 (N_13261,N_13241,N_13161);
xor U13262 (N_13262,N_13187,N_13142);
xor U13263 (N_13263,N_13130,N_13188);
nor U13264 (N_13264,N_13170,N_13239);
and U13265 (N_13265,N_13225,N_13201);
nand U13266 (N_13266,N_13234,N_13204);
nor U13267 (N_13267,N_13126,N_13228);
and U13268 (N_13268,N_13217,N_13155);
or U13269 (N_13269,N_13191,N_13205);
xor U13270 (N_13270,N_13182,N_13180);
or U13271 (N_13271,N_13199,N_13168);
nand U13272 (N_13272,N_13238,N_13203);
nand U13273 (N_13273,N_13236,N_13165);
nand U13274 (N_13274,N_13131,N_13202);
and U13275 (N_13275,N_13212,N_13240);
nor U13276 (N_13276,N_13148,N_13136);
or U13277 (N_13277,N_13172,N_13218);
nand U13278 (N_13278,N_13197,N_13195);
nand U13279 (N_13279,N_13153,N_13229);
or U13280 (N_13280,N_13149,N_13214);
nand U13281 (N_13281,N_13237,N_13175);
nand U13282 (N_13282,N_13179,N_13176);
nor U13283 (N_13283,N_13139,N_13190);
xor U13284 (N_13284,N_13220,N_13213);
xor U13285 (N_13285,N_13183,N_13135);
nor U13286 (N_13286,N_13207,N_13127);
xor U13287 (N_13287,N_13162,N_13128);
or U13288 (N_13288,N_13209,N_13158);
xnor U13289 (N_13289,N_13184,N_13224);
xnor U13290 (N_13290,N_13156,N_13167);
and U13291 (N_13291,N_13164,N_13166);
and U13292 (N_13292,N_13134,N_13129);
and U13293 (N_13293,N_13146,N_13125);
and U13294 (N_13294,N_13152,N_13157);
or U13295 (N_13295,N_13140,N_13150);
or U13296 (N_13296,N_13246,N_13159);
and U13297 (N_13297,N_13169,N_13231);
nand U13298 (N_13298,N_13174,N_13208);
nand U13299 (N_13299,N_13244,N_13192);
or U13300 (N_13300,N_13143,N_13206);
xnor U13301 (N_13301,N_13185,N_13144);
or U13302 (N_13302,N_13222,N_13147);
or U13303 (N_13303,N_13173,N_13189);
nand U13304 (N_13304,N_13200,N_13177);
or U13305 (N_13305,N_13230,N_13249);
xor U13306 (N_13306,N_13232,N_13194);
xor U13307 (N_13307,N_13163,N_13216);
nand U13308 (N_13308,N_13132,N_13196);
nand U13309 (N_13309,N_13235,N_13151);
nand U13310 (N_13310,N_13171,N_13233);
nor U13311 (N_13311,N_13210,N_13181);
or U13312 (N_13312,N_13247,N_13195);
and U13313 (N_13313,N_13169,N_13156);
or U13314 (N_13314,N_13184,N_13223);
and U13315 (N_13315,N_13142,N_13220);
nor U13316 (N_13316,N_13245,N_13201);
xor U13317 (N_13317,N_13204,N_13181);
and U13318 (N_13318,N_13204,N_13158);
nor U13319 (N_13319,N_13191,N_13217);
or U13320 (N_13320,N_13147,N_13198);
or U13321 (N_13321,N_13221,N_13225);
nor U13322 (N_13322,N_13213,N_13229);
nor U13323 (N_13323,N_13198,N_13156);
nand U13324 (N_13324,N_13226,N_13151);
or U13325 (N_13325,N_13238,N_13192);
nand U13326 (N_13326,N_13184,N_13227);
and U13327 (N_13327,N_13206,N_13230);
nor U13328 (N_13328,N_13158,N_13201);
or U13329 (N_13329,N_13229,N_13224);
nor U13330 (N_13330,N_13148,N_13181);
nor U13331 (N_13331,N_13175,N_13208);
nand U13332 (N_13332,N_13206,N_13165);
nor U13333 (N_13333,N_13184,N_13218);
or U13334 (N_13334,N_13128,N_13211);
nor U13335 (N_13335,N_13126,N_13170);
nor U13336 (N_13336,N_13152,N_13153);
nor U13337 (N_13337,N_13174,N_13155);
and U13338 (N_13338,N_13218,N_13129);
xnor U13339 (N_13339,N_13127,N_13219);
xnor U13340 (N_13340,N_13236,N_13183);
nand U13341 (N_13341,N_13228,N_13185);
or U13342 (N_13342,N_13143,N_13243);
and U13343 (N_13343,N_13196,N_13186);
and U13344 (N_13344,N_13126,N_13194);
xnor U13345 (N_13345,N_13134,N_13170);
xnor U13346 (N_13346,N_13185,N_13199);
or U13347 (N_13347,N_13239,N_13199);
or U13348 (N_13348,N_13182,N_13166);
and U13349 (N_13349,N_13214,N_13186);
nand U13350 (N_13350,N_13155,N_13238);
nand U13351 (N_13351,N_13137,N_13153);
xor U13352 (N_13352,N_13132,N_13229);
and U13353 (N_13353,N_13204,N_13186);
and U13354 (N_13354,N_13205,N_13167);
and U13355 (N_13355,N_13212,N_13207);
xnor U13356 (N_13356,N_13222,N_13232);
nand U13357 (N_13357,N_13167,N_13199);
or U13358 (N_13358,N_13178,N_13236);
xor U13359 (N_13359,N_13168,N_13212);
xnor U13360 (N_13360,N_13197,N_13149);
nor U13361 (N_13361,N_13210,N_13128);
nand U13362 (N_13362,N_13162,N_13127);
nand U13363 (N_13363,N_13178,N_13153);
nor U13364 (N_13364,N_13206,N_13238);
nand U13365 (N_13365,N_13126,N_13219);
nor U13366 (N_13366,N_13202,N_13156);
and U13367 (N_13367,N_13242,N_13127);
and U13368 (N_13368,N_13231,N_13126);
or U13369 (N_13369,N_13211,N_13192);
or U13370 (N_13370,N_13153,N_13166);
nand U13371 (N_13371,N_13242,N_13154);
or U13372 (N_13372,N_13206,N_13210);
nor U13373 (N_13373,N_13127,N_13229);
or U13374 (N_13374,N_13199,N_13234);
xnor U13375 (N_13375,N_13356,N_13311);
or U13376 (N_13376,N_13358,N_13339);
xnor U13377 (N_13377,N_13346,N_13261);
nor U13378 (N_13378,N_13326,N_13351);
and U13379 (N_13379,N_13255,N_13372);
nand U13380 (N_13380,N_13312,N_13287);
xor U13381 (N_13381,N_13363,N_13341);
nor U13382 (N_13382,N_13270,N_13253);
nand U13383 (N_13383,N_13268,N_13316);
or U13384 (N_13384,N_13303,N_13335);
nor U13385 (N_13385,N_13337,N_13264);
nor U13386 (N_13386,N_13265,N_13362);
xnor U13387 (N_13387,N_13294,N_13347);
or U13388 (N_13388,N_13350,N_13252);
nand U13389 (N_13389,N_13323,N_13327);
or U13390 (N_13390,N_13359,N_13319);
nor U13391 (N_13391,N_13353,N_13330);
and U13392 (N_13392,N_13277,N_13259);
or U13393 (N_13393,N_13299,N_13297);
and U13394 (N_13394,N_13331,N_13352);
nor U13395 (N_13395,N_13364,N_13269);
xor U13396 (N_13396,N_13320,N_13355);
nor U13397 (N_13397,N_13317,N_13283);
nor U13398 (N_13398,N_13266,N_13344);
and U13399 (N_13399,N_13334,N_13325);
nor U13400 (N_13400,N_13286,N_13354);
nor U13401 (N_13401,N_13298,N_13285);
nor U13402 (N_13402,N_13342,N_13302);
or U13403 (N_13403,N_13371,N_13257);
or U13404 (N_13404,N_13365,N_13292);
and U13405 (N_13405,N_13310,N_13276);
xor U13406 (N_13406,N_13289,N_13338);
nand U13407 (N_13407,N_13306,N_13258);
nand U13408 (N_13408,N_13263,N_13280);
and U13409 (N_13409,N_13281,N_13274);
nor U13410 (N_13410,N_13332,N_13251);
nor U13411 (N_13411,N_13307,N_13357);
nor U13412 (N_13412,N_13315,N_13328);
and U13413 (N_13413,N_13288,N_13300);
nand U13414 (N_13414,N_13275,N_13305);
nor U13415 (N_13415,N_13296,N_13278);
xor U13416 (N_13416,N_13295,N_13260);
xor U13417 (N_13417,N_13343,N_13308);
xor U13418 (N_13418,N_13322,N_13267);
and U13419 (N_13419,N_13290,N_13368);
nor U13420 (N_13420,N_13272,N_13348);
nor U13421 (N_13421,N_13271,N_13324);
or U13422 (N_13422,N_13340,N_13250);
xor U13423 (N_13423,N_13279,N_13321);
nand U13424 (N_13424,N_13313,N_13370);
and U13425 (N_13425,N_13336,N_13273);
xnor U13426 (N_13426,N_13329,N_13291);
nor U13427 (N_13427,N_13304,N_13284);
nand U13428 (N_13428,N_13333,N_13361);
xnor U13429 (N_13429,N_13366,N_13318);
nand U13430 (N_13430,N_13369,N_13301);
nor U13431 (N_13431,N_13314,N_13254);
nand U13432 (N_13432,N_13345,N_13256);
nor U13433 (N_13433,N_13360,N_13282);
or U13434 (N_13434,N_13293,N_13309);
nor U13435 (N_13435,N_13374,N_13367);
xnor U13436 (N_13436,N_13373,N_13349);
xor U13437 (N_13437,N_13262,N_13359);
or U13438 (N_13438,N_13373,N_13320);
nor U13439 (N_13439,N_13307,N_13356);
xor U13440 (N_13440,N_13357,N_13308);
nand U13441 (N_13441,N_13315,N_13357);
nor U13442 (N_13442,N_13329,N_13264);
nand U13443 (N_13443,N_13305,N_13366);
and U13444 (N_13444,N_13272,N_13309);
and U13445 (N_13445,N_13294,N_13349);
or U13446 (N_13446,N_13311,N_13352);
nor U13447 (N_13447,N_13289,N_13307);
and U13448 (N_13448,N_13372,N_13323);
and U13449 (N_13449,N_13333,N_13253);
xor U13450 (N_13450,N_13296,N_13304);
nor U13451 (N_13451,N_13261,N_13359);
xor U13452 (N_13452,N_13288,N_13319);
and U13453 (N_13453,N_13333,N_13312);
and U13454 (N_13454,N_13368,N_13284);
nor U13455 (N_13455,N_13355,N_13333);
nand U13456 (N_13456,N_13328,N_13277);
nand U13457 (N_13457,N_13333,N_13258);
nor U13458 (N_13458,N_13288,N_13316);
or U13459 (N_13459,N_13256,N_13297);
and U13460 (N_13460,N_13341,N_13343);
or U13461 (N_13461,N_13355,N_13265);
xnor U13462 (N_13462,N_13335,N_13251);
nand U13463 (N_13463,N_13324,N_13265);
nor U13464 (N_13464,N_13354,N_13360);
or U13465 (N_13465,N_13262,N_13259);
xnor U13466 (N_13466,N_13289,N_13254);
nand U13467 (N_13467,N_13268,N_13370);
and U13468 (N_13468,N_13347,N_13335);
nor U13469 (N_13469,N_13277,N_13312);
nor U13470 (N_13470,N_13283,N_13266);
nand U13471 (N_13471,N_13353,N_13348);
and U13472 (N_13472,N_13308,N_13365);
or U13473 (N_13473,N_13291,N_13353);
and U13474 (N_13474,N_13366,N_13283);
nor U13475 (N_13475,N_13367,N_13298);
and U13476 (N_13476,N_13356,N_13308);
nor U13477 (N_13477,N_13253,N_13338);
and U13478 (N_13478,N_13346,N_13300);
xor U13479 (N_13479,N_13282,N_13272);
or U13480 (N_13480,N_13312,N_13344);
nor U13481 (N_13481,N_13310,N_13320);
nand U13482 (N_13482,N_13280,N_13347);
and U13483 (N_13483,N_13301,N_13347);
and U13484 (N_13484,N_13362,N_13261);
nor U13485 (N_13485,N_13298,N_13316);
xor U13486 (N_13486,N_13343,N_13317);
nor U13487 (N_13487,N_13366,N_13347);
and U13488 (N_13488,N_13305,N_13259);
or U13489 (N_13489,N_13297,N_13257);
xnor U13490 (N_13490,N_13255,N_13346);
nand U13491 (N_13491,N_13285,N_13356);
nand U13492 (N_13492,N_13299,N_13274);
nor U13493 (N_13493,N_13323,N_13284);
and U13494 (N_13494,N_13278,N_13314);
nand U13495 (N_13495,N_13353,N_13299);
nand U13496 (N_13496,N_13334,N_13276);
and U13497 (N_13497,N_13357,N_13294);
xor U13498 (N_13498,N_13360,N_13253);
and U13499 (N_13499,N_13262,N_13307);
nand U13500 (N_13500,N_13413,N_13392);
or U13501 (N_13501,N_13437,N_13452);
and U13502 (N_13502,N_13435,N_13398);
nor U13503 (N_13503,N_13471,N_13430);
nand U13504 (N_13504,N_13462,N_13376);
xnor U13505 (N_13505,N_13414,N_13388);
nor U13506 (N_13506,N_13459,N_13434);
nor U13507 (N_13507,N_13383,N_13492);
and U13508 (N_13508,N_13410,N_13389);
xor U13509 (N_13509,N_13404,N_13440);
nor U13510 (N_13510,N_13451,N_13443);
nand U13511 (N_13511,N_13401,N_13381);
nand U13512 (N_13512,N_13424,N_13411);
xnor U13513 (N_13513,N_13466,N_13453);
and U13514 (N_13514,N_13409,N_13419);
nand U13515 (N_13515,N_13490,N_13436);
and U13516 (N_13516,N_13426,N_13432);
or U13517 (N_13517,N_13438,N_13461);
xor U13518 (N_13518,N_13416,N_13463);
nand U13519 (N_13519,N_13470,N_13449);
nand U13520 (N_13520,N_13429,N_13395);
nand U13521 (N_13521,N_13464,N_13380);
or U13522 (N_13522,N_13390,N_13397);
xor U13523 (N_13523,N_13495,N_13442);
nand U13524 (N_13524,N_13387,N_13486);
or U13525 (N_13525,N_13445,N_13427);
xor U13526 (N_13526,N_13483,N_13420);
nand U13527 (N_13527,N_13407,N_13402);
nand U13528 (N_13528,N_13405,N_13487);
nor U13529 (N_13529,N_13473,N_13396);
and U13530 (N_13530,N_13481,N_13493);
or U13531 (N_13531,N_13446,N_13384);
nor U13532 (N_13532,N_13391,N_13458);
nor U13533 (N_13533,N_13467,N_13423);
xnor U13534 (N_13534,N_13491,N_13468);
and U13535 (N_13535,N_13499,N_13476);
or U13536 (N_13536,N_13386,N_13417);
and U13537 (N_13537,N_13441,N_13496);
or U13538 (N_13538,N_13484,N_13379);
and U13539 (N_13539,N_13480,N_13469);
xor U13540 (N_13540,N_13465,N_13393);
xor U13541 (N_13541,N_13428,N_13497);
or U13542 (N_13542,N_13450,N_13394);
or U13543 (N_13543,N_13412,N_13457);
or U13544 (N_13544,N_13474,N_13375);
and U13545 (N_13545,N_13482,N_13455);
xor U13546 (N_13546,N_13415,N_13399);
nand U13547 (N_13547,N_13378,N_13439);
nand U13548 (N_13548,N_13422,N_13475);
or U13549 (N_13549,N_13385,N_13377);
nor U13550 (N_13550,N_13485,N_13406);
nor U13551 (N_13551,N_13421,N_13403);
and U13552 (N_13552,N_13448,N_13456);
nor U13553 (N_13553,N_13488,N_13447);
nand U13554 (N_13554,N_13477,N_13382);
or U13555 (N_13555,N_13433,N_13454);
nand U13556 (N_13556,N_13408,N_13444);
nor U13557 (N_13557,N_13494,N_13479);
xor U13558 (N_13558,N_13418,N_13472);
or U13559 (N_13559,N_13431,N_13425);
nor U13560 (N_13560,N_13478,N_13498);
or U13561 (N_13561,N_13460,N_13400);
nand U13562 (N_13562,N_13489,N_13403);
nor U13563 (N_13563,N_13432,N_13386);
or U13564 (N_13564,N_13496,N_13404);
xor U13565 (N_13565,N_13425,N_13428);
or U13566 (N_13566,N_13426,N_13462);
xor U13567 (N_13567,N_13493,N_13477);
nor U13568 (N_13568,N_13393,N_13444);
xnor U13569 (N_13569,N_13418,N_13459);
nand U13570 (N_13570,N_13484,N_13474);
or U13571 (N_13571,N_13412,N_13481);
nand U13572 (N_13572,N_13473,N_13379);
and U13573 (N_13573,N_13466,N_13376);
nor U13574 (N_13574,N_13411,N_13488);
and U13575 (N_13575,N_13481,N_13384);
xor U13576 (N_13576,N_13460,N_13382);
and U13577 (N_13577,N_13429,N_13488);
and U13578 (N_13578,N_13416,N_13415);
xnor U13579 (N_13579,N_13444,N_13463);
nor U13580 (N_13580,N_13413,N_13488);
or U13581 (N_13581,N_13387,N_13400);
xnor U13582 (N_13582,N_13382,N_13398);
nor U13583 (N_13583,N_13497,N_13446);
or U13584 (N_13584,N_13401,N_13407);
nand U13585 (N_13585,N_13430,N_13425);
nand U13586 (N_13586,N_13468,N_13399);
nor U13587 (N_13587,N_13425,N_13382);
nor U13588 (N_13588,N_13437,N_13384);
nand U13589 (N_13589,N_13379,N_13385);
nor U13590 (N_13590,N_13455,N_13471);
nor U13591 (N_13591,N_13469,N_13385);
xor U13592 (N_13592,N_13476,N_13378);
xnor U13593 (N_13593,N_13421,N_13417);
and U13594 (N_13594,N_13422,N_13483);
or U13595 (N_13595,N_13442,N_13445);
or U13596 (N_13596,N_13457,N_13467);
xnor U13597 (N_13597,N_13424,N_13489);
xor U13598 (N_13598,N_13420,N_13484);
nand U13599 (N_13599,N_13483,N_13456);
nand U13600 (N_13600,N_13456,N_13485);
and U13601 (N_13601,N_13376,N_13485);
xnor U13602 (N_13602,N_13469,N_13432);
xnor U13603 (N_13603,N_13384,N_13417);
or U13604 (N_13604,N_13447,N_13467);
or U13605 (N_13605,N_13395,N_13393);
nand U13606 (N_13606,N_13375,N_13389);
nor U13607 (N_13607,N_13410,N_13432);
nand U13608 (N_13608,N_13446,N_13375);
nand U13609 (N_13609,N_13399,N_13441);
nand U13610 (N_13610,N_13429,N_13490);
xor U13611 (N_13611,N_13436,N_13456);
xor U13612 (N_13612,N_13390,N_13493);
xor U13613 (N_13613,N_13460,N_13386);
nor U13614 (N_13614,N_13479,N_13405);
or U13615 (N_13615,N_13452,N_13471);
xor U13616 (N_13616,N_13393,N_13380);
xor U13617 (N_13617,N_13440,N_13473);
and U13618 (N_13618,N_13407,N_13494);
and U13619 (N_13619,N_13440,N_13407);
and U13620 (N_13620,N_13397,N_13460);
or U13621 (N_13621,N_13380,N_13383);
nor U13622 (N_13622,N_13378,N_13446);
xor U13623 (N_13623,N_13497,N_13438);
xnor U13624 (N_13624,N_13388,N_13484);
nor U13625 (N_13625,N_13595,N_13532);
nor U13626 (N_13626,N_13517,N_13516);
xor U13627 (N_13627,N_13530,N_13520);
xnor U13628 (N_13628,N_13577,N_13536);
nand U13629 (N_13629,N_13620,N_13579);
xor U13630 (N_13630,N_13539,N_13552);
xnor U13631 (N_13631,N_13515,N_13564);
nand U13632 (N_13632,N_13575,N_13518);
nor U13633 (N_13633,N_13533,N_13583);
nand U13634 (N_13634,N_13510,N_13611);
nor U13635 (N_13635,N_13580,N_13567);
and U13636 (N_13636,N_13589,N_13555);
xnor U13637 (N_13637,N_13599,N_13556);
xnor U13638 (N_13638,N_13565,N_13561);
nand U13639 (N_13639,N_13519,N_13607);
and U13640 (N_13640,N_13571,N_13598);
xor U13641 (N_13641,N_13616,N_13551);
nand U13642 (N_13642,N_13542,N_13506);
nand U13643 (N_13643,N_13509,N_13608);
and U13644 (N_13644,N_13544,N_13553);
or U13645 (N_13645,N_13524,N_13572);
nand U13646 (N_13646,N_13568,N_13507);
or U13647 (N_13647,N_13514,N_13581);
xor U13648 (N_13648,N_13601,N_13610);
or U13649 (N_13649,N_13606,N_13508);
and U13650 (N_13650,N_13502,N_13574);
nand U13651 (N_13651,N_13623,N_13535);
nand U13652 (N_13652,N_13554,N_13604);
and U13653 (N_13653,N_13602,N_13569);
nor U13654 (N_13654,N_13600,N_13513);
nand U13655 (N_13655,N_13566,N_13558);
or U13656 (N_13656,N_13585,N_13547);
or U13657 (N_13657,N_13541,N_13503);
or U13658 (N_13658,N_13527,N_13545);
or U13659 (N_13659,N_13563,N_13578);
nand U13660 (N_13660,N_13549,N_13605);
or U13661 (N_13661,N_13531,N_13543);
and U13662 (N_13662,N_13612,N_13624);
or U13663 (N_13663,N_13609,N_13614);
nand U13664 (N_13664,N_13560,N_13621);
xnor U13665 (N_13665,N_13592,N_13573);
nor U13666 (N_13666,N_13500,N_13504);
or U13667 (N_13667,N_13590,N_13562);
nor U13668 (N_13668,N_13529,N_13617);
or U13669 (N_13669,N_13523,N_13587);
nor U13670 (N_13670,N_13512,N_13522);
nor U13671 (N_13671,N_13538,N_13588);
xor U13672 (N_13672,N_13586,N_13570);
xnor U13673 (N_13673,N_13534,N_13505);
xor U13674 (N_13674,N_13559,N_13584);
nor U13675 (N_13675,N_13501,N_13594);
xnor U13676 (N_13676,N_13526,N_13525);
xor U13677 (N_13677,N_13591,N_13528);
xnor U13678 (N_13678,N_13540,N_13603);
or U13679 (N_13679,N_13619,N_13511);
nand U13680 (N_13680,N_13593,N_13557);
and U13681 (N_13681,N_13613,N_13550);
or U13682 (N_13682,N_13596,N_13521);
nor U13683 (N_13683,N_13576,N_13546);
xnor U13684 (N_13684,N_13615,N_13548);
and U13685 (N_13685,N_13537,N_13582);
xnor U13686 (N_13686,N_13622,N_13618);
nor U13687 (N_13687,N_13597,N_13513);
nand U13688 (N_13688,N_13569,N_13504);
nor U13689 (N_13689,N_13516,N_13535);
or U13690 (N_13690,N_13518,N_13527);
and U13691 (N_13691,N_13570,N_13534);
nor U13692 (N_13692,N_13587,N_13571);
and U13693 (N_13693,N_13522,N_13549);
or U13694 (N_13694,N_13537,N_13504);
or U13695 (N_13695,N_13515,N_13523);
and U13696 (N_13696,N_13516,N_13593);
or U13697 (N_13697,N_13590,N_13576);
nand U13698 (N_13698,N_13608,N_13539);
nor U13699 (N_13699,N_13581,N_13563);
or U13700 (N_13700,N_13582,N_13610);
or U13701 (N_13701,N_13520,N_13549);
nor U13702 (N_13702,N_13603,N_13520);
nor U13703 (N_13703,N_13572,N_13598);
or U13704 (N_13704,N_13622,N_13543);
and U13705 (N_13705,N_13578,N_13591);
and U13706 (N_13706,N_13566,N_13601);
and U13707 (N_13707,N_13624,N_13555);
nor U13708 (N_13708,N_13622,N_13623);
nor U13709 (N_13709,N_13502,N_13608);
or U13710 (N_13710,N_13613,N_13581);
xnor U13711 (N_13711,N_13507,N_13596);
nand U13712 (N_13712,N_13575,N_13574);
nor U13713 (N_13713,N_13534,N_13546);
and U13714 (N_13714,N_13512,N_13596);
xnor U13715 (N_13715,N_13563,N_13521);
nor U13716 (N_13716,N_13599,N_13545);
xor U13717 (N_13717,N_13591,N_13575);
nand U13718 (N_13718,N_13623,N_13553);
nor U13719 (N_13719,N_13611,N_13575);
nor U13720 (N_13720,N_13588,N_13602);
or U13721 (N_13721,N_13618,N_13565);
and U13722 (N_13722,N_13509,N_13531);
nor U13723 (N_13723,N_13578,N_13618);
or U13724 (N_13724,N_13541,N_13552);
nor U13725 (N_13725,N_13609,N_13563);
nor U13726 (N_13726,N_13608,N_13505);
xor U13727 (N_13727,N_13595,N_13552);
nand U13728 (N_13728,N_13502,N_13571);
xnor U13729 (N_13729,N_13571,N_13552);
nor U13730 (N_13730,N_13574,N_13554);
xor U13731 (N_13731,N_13502,N_13550);
xnor U13732 (N_13732,N_13535,N_13504);
nor U13733 (N_13733,N_13556,N_13563);
or U13734 (N_13734,N_13527,N_13596);
nor U13735 (N_13735,N_13614,N_13591);
nor U13736 (N_13736,N_13596,N_13550);
and U13737 (N_13737,N_13501,N_13583);
nor U13738 (N_13738,N_13568,N_13595);
nand U13739 (N_13739,N_13594,N_13613);
xnor U13740 (N_13740,N_13553,N_13594);
and U13741 (N_13741,N_13576,N_13595);
and U13742 (N_13742,N_13612,N_13568);
nand U13743 (N_13743,N_13502,N_13617);
or U13744 (N_13744,N_13585,N_13603);
and U13745 (N_13745,N_13586,N_13515);
xnor U13746 (N_13746,N_13536,N_13513);
or U13747 (N_13747,N_13537,N_13602);
xnor U13748 (N_13748,N_13536,N_13501);
or U13749 (N_13749,N_13507,N_13567);
and U13750 (N_13750,N_13687,N_13700);
xnor U13751 (N_13751,N_13630,N_13627);
or U13752 (N_13752,N_13738,N_13660);
xor U13753 (N_13753,N_13680,N_13723);
and U13754 (N_13754,N_13737,N_13646);
xnor U13755 (N_13755,N_13747,N_13672);
xnor U13756 (N_13756,N_13724,N_13742);
nor U13757 (N_13757,N_13749,N_13695);
nand U13758 (N_13758,N_13639,N_13744);
and U13759 (N_13759,N_13642,N_13625);
or U13760 (N_13760,N_13740,N_13676);
xor U13761 (N_13761,N_13734,N_13631);
nand U13762 (N_13762,N_13716,N_13665);
nand U13763 (N_13763,N_13645,N_13638);
nor U13764 (N_13764,N_13629,N_13654);
nand U13765 (N_13765,N_13713,N_13636);
nor U13766 (N_13766,N_13691,N_13682);
nand U13767 (N_13767,N_13667,N_13641);
or U13768 (N_13768,N_13733,N_13649);
and U13769 (N_13769,N_13739,N_13628);
and U13770 (N_13770,N_13640,N_13675);
xor U13771 (N_13771,N_13717,N_13666);
or U13772 (N_13772,N_13719,N_13729);
and U13773 (N_13773,N_13726,N_13648);
or U13774 (N_13774,N_13702,N_13690);
or U13775 (N_13775,N_13634,N_13709);
xor U13776 (N_13776,N_13678,N_13721);
nor U13777 (N_13777,N_13712,N_13741);
nand U13778 (N_13778,N_13635,N_13657);
xnor U13779 (N_13779,N_13650,N_13699);
and U13780 (N_13780,N_13688,N_13673);
nand U13781 (N_13781,N_13732,N_13663);
nand U13782 (N_13782,N_13668,N_13633);
and U13783 (N_13783,N_13664,N_13743);
and U13784 (N_13784,N_13707,N_13693);
xor U13785 (N_13785,N_13658,N_13661);
or U13786 (N_13786,N_13725,N_13647);
and U13787 (N_13787,N_13683,N_13643);
nor U13788 (N_13788,N_13670,N_13727);
or U13789 (N_13789,N_13656,N_13731);
nor U13790 (N_13790,N_13706,N_13708);
and U13791 (N_13791,N_13689,N_13748);
and U13792 (N_13792,N_13644,N_13718);
or U13793 (N_13793,N_13626,N_13653);
and U13794 (N_13794,N_13685,N_13637);
and U13795 (N_13795,N_13681,N_13704);
nand U13796 (N_13796,N_13651,N_13715);
nor U13797 (N_13797,N_13655,N_13659);
nor U13798 (N_13798,N_13694,N_13703);
xor U13799 (N_13799,N_13710,N_13720);
nor U13800 (N_13800,N_13686,N_13714);
xor U13801 (N_13801,N_13698,N_13679);
nand U13802 (N_13802,N_13728,N_13696);
nand U13803 (N_13803,N_13652,N_13662);
or U13804 (N_13804,N_13669,N_13632);
xnor U13805 (N_13805,N_13722,N_13730);
nand U13806 (N_13806,N_13671,N_13674);
nand U13807 (N_13807,N_13684,N_13692);
and U13808 (N_13808,N_13735,N_13677);
xnor U13809 (N_13809,N_13701,N_13705);
or U13810 (N_13810,N_13745,N_13711);
xnor U13811 (N_13811,N_13736,N_13697);
or U13812 (N_13812,N_13746,N_13656);
and U13813 (N_13813,N_13638,N_13643);
nand U13814 (N_13814,N_13732,N_13699);
nand U13815 (N_13815,N_13742,N_13749);
nor U13816 (N_13816,N_13715,N_13692);
and U13817 (N_13817,N_13664,N_13694);
nor U13818 (N_13818,N_13629,N_13725);
nor U13819 (N_13819,N_13718,N_13626);
or U13820 (N_13820,N_13639,N_13659);
nor U13821 (N_13821,N_13659,N_13652);
and U13822 (N_13822,N_13631,N_13644);
or U13823 (N_13823,N_13697,N_13671);
and U13824 (N_13824,N_13740,N_13730);
xor U13825 (N_13825,N_13710,N_13655);
and U13826 (N_13826,N_13674,N_13731);
and U13827 (N_13827,N_13670,N_13669);
xnor U13828 (N_13828,N_13674,N_13703);
xnor U13829 (N_13829,N_13675,N_13714);
nor U13830 (N_13830,N_13630,N_13736);
and U13831 (N_13831,N_13725,N_13745);
nor U13832 (N_13832,N_13697,N_13651);
or U13833 (N_13833,N_13724,N_13709);
and U13834 (N_13834,N_13672,N_13697);
nand U13835 (N_13835,N_13747,N_13704);
and U13836 (N_13836,N_13648,N_13732);
nand U13837 (N_13837,N_13746,N_13658);
or U13838 (N_13838,N_13627,N_13628);
or U13839 (N_13839,N_13669,N_13672);
xnor U13840 (N_13840,N_13649,N_13661);
nor U13841 (N_13841,N_13711,N_13738);
nand U13842 (N_13842,N_13653,N_13748);
xor U13843 (N_13843,N_13665,N_13668);
nor U13844 (N_13844,N_13728,N_13700);
nand U13845 (N_13845,N_13631,N_13635);
and U13846 (N_13846,N_13689,N_13678);
nor U13847 (N_13847,N_13665,N_13640);
nor U13848 (N_13848,N_13691,N_13731);
or U13849 (N_13849,N_13739,N_13652);
or U13850 (N_13850,N_13701,N_13723);
or U13851 (N_13851,N_13637,N_13675);
nor U13852 (N_13852,N_13704,N_13723);
and U13853 (N_13853,N_13745,N_13706);
and U13854 (N_13854,N_13690,N_13664);
or U13855 (N_13855,N_13668,N_13694);
nor U13856 (N_13856,N_13710,N_13628);
nand U13857 (N_13857,N_13705,N_13661);
nand U13858 (N_13858,N_13669,N_13724);
xor U13859 (N_13859,N_13651,N_13637);
or U13860 (N_13860,N_13703,N_13700);
xor U13861 (N_13861,N_13649,N_13628);
nand U13862 (N_13862,N_13680,N_13686);
xnor U13863 (N_13863,N_13664,N_13654);
and U13864 (N_13864,N_13646,N_13665);
or U13865 (N_13865,N_13635,N_13666);
nor U13866 (N_13866,N_13682,N_13643);
or U13867 (N_13867,N_13674,N_13649);
xor U13868 (N_13868,N_13666,N_13745);
and U13869 (N_13869,N_13672,N_13740);
nor U13870 (N_13870,N_13670,N_13658);
nor U13871 (N_13871,N_13708,N_13732);
nand U13872 (N_13872,N_13713,N_13672);
or U13873 (N_13873,N_13681,N_13669);
or U13874 (N_13874,N_13749,N_13713);
nor U13875 (N_13875,N_13782,N_13872);
and U13876 (N_13876,N_13806,N_13772);
nand U13877 (N_13877,N_13862,N_13774);
xor U13878 (N_13878,N_13771,N_13834);
xnor U13879 (N_13879,N_13765,N_13792);
nand U13880 (N_13880,N_13819,N_13830);
nand U13881 (N_13881,N_13785,N_13768);
or U13882 (N_13882,N_13803,N_13776);
or U13883 (N_13883,N_13754,N_13863);
xnor U13884 (N_13884,N_13851,N_13760);
nand U13885 (N_13885,N_13859,N_13786);
or U13886 (N_13886,N_13815,N_13758);
nand U13887 (N_13887,N_13751,N_13807);
nor U13888 (N_13888,N_13844,N_13867);
or U13889 (N_13889,N_13823,N_13854);
nand U13890 (N_13890,N_13865,N_13802);
nand U13891 (N_13891,N_13769,N_13864);
or U13892 (N_13892,N_13812,N_13857);
xor U13893 (N_13893,N_13753,N_13842);
xnor U13894 (N_13894,N_13779,N_13836);
nor U13895 (N_13895,N_13831,N_13797);
and U13896 (N_13896,N_13853,N_13759);
xor U13897 (N_13897,N_13874,N_13809);
nand U13898 (N_13898,N_13808,N_13794);
or U13899 (N_13899,N_13852,N_13840);
xor U13900 (N_13900,N_13843,N_13773);
nand U13901 (N_13901,N_13817,N_13798);
nor U13902 (N_13902,N_13833,N_13821);
xnor U13903 (N_13903,N_13757,N_13849);
nand U13904 (N_13904,N_13832,N_13778);
nor U13905 (N_13905,N_13861,N_13869);
nand U13906 (N_13906,N_13847,N_13777);
xor U13907 (N_13907,N_13795,N_13837);
xnor U13908 (N_13908,N_13766,N_13791);
xnor U13909 (N_13909,N_13820,N_13784);
nor U13910 (N_13910,N_13755,N_13846);
xnor U13911 (N_13911,N_13767,N_13873);
xnor U13912 (N_13912,N_13860,N_13845);
nand U13913 (N_13913,N_13848,N_13870);
xnor U13914 (N_13914,N_13855,N_13871);
or U13915 (N_13915,N_13826,N_13829);
xor U13916 (N_13916,N_13762,N_13801);
and U13917 (N_13917,N_13796,N_13813);
nand U13918 (N_13918,N_13788,N_13841);
and U13919 (N_13919,N_13800,N_13763);
or U13920 (N_13920,N_13824,N_13816);
nand U13921 (N_13921,N_13799,N_13814);
and U13922 (N_13922,N_13827,N_13856);
nor U13923 (N_13923,N_13858,N_13750);
or U13924 (N_13924,N_13839,N_13761);
nor U13925 (N_13925,N_13805,N_13764);
or U13926 (N_13926,N_13838,N_13793);
nor U13927 (N_13927,N_13783,N_13850);
and U13928 (N_13928,N_13811,N_13789);
xor U13929 (N_13929,N_13752,N_13868);
nand U13930 (N_13930,N_13790,N_13775);
xor U13931 (N_13931,N_13756,N_13828);
or U13932 (N_13932,N_13825,N_13804);
or U13933 (N_13933,N_13818,N_13787);
or U13934 (N_13934,N_13822,N_13866);
xor U13935 (N_13935,N_13835,N_13810);
nand U13936 (N_13936,N_13770,N_13780);
nor U13937 (N_13937,N_13781,N_13843);
and U13938 (N_13938,N_13851,N_13828);
nand U13939 (N_13939,N_13823,N_13812);
nor U13940 (N_13940,N_13788,N_13798);
or U13941 (N_13941,N_13787,N_13758);
or U13942 (N_13942,N_13874,N_13787);
and U13943 (N_13943,N_13861,N_13758);
xnor U13944 (N_13944,N_13840,N_13757);
and U13945 (N_13945,N_13787,N_13782);
and U13946 (N_13946,N_13817,N_13815);
or U13947 (N_13947,N_13797,N_13809);
nor U13948 (N_13948,N_13781,N_13833);
xnor U13949 (N_13949,N_13796,N_13755);
and U13950 (N_13950,N_13801,N_13846);
or U13951 (N_13951,N_13796,N_13848);
xnor U13952 (N_13952,N_13780,N_13787);
nor U13953 (N_13953,N_13841,N_13792);
nand U13954 (N_13954,N_13834,N_13786);
or U13955 (N_13955,N_13789,N_13855);
xnor U13956 (N_13956,N_13752,N_13823);
xnor U13957 (N_13957,N_13859,N_13857);
or U13958 (N_13958,N_13854,N_13852);
or U13959 (N_13959,N_13764,N_13788);
nor U13960 (N_13960,N_13791,N_13845);
or U13961 (N_13961,N_13758,N_13828);
xnor U13962 (N_13962,N_13849,N_13824);
nand U13963 (N_13963,N_13859,N_13766);
nand U13964 (N_13964,N_13781,N_13776);
nor U13965 (N_13965,N_13853,N_13865);
nand U13966 (N_13966,N_13831,N_13833);
and U13967 (N_13967,N_13757,N_13869);
or U13968 (N_13968,N_13823,N_13852);
nor U13969 (N_13969,N_13796,N_13787);
xor U13970 (N_13970,N_13766,N_13788);
and U13971 (N_13971,N_13872,N_13804);
nor U13972 (N_13972,N_13811,N_13871);
and U13973 (N_13973,N_13853,N_13796);
nor U13974 (N_13974,N_13840,N_13779);
nand U13975 (N_13975,N_13778,N_13809);
nor U13976 (N_13976,N_13772,N_13757);
or U13977 (N_13977,N_13851,N_13792);
or U13978 (N_13978,N_13776,N_13840);
or U13979 (N_13979,N_13829,N_13774);
nand U13980 (N_13980,N_13786,N_13794);
nor U13981 (N_13981,N_13815,N_13775);
xnor U13982 (N_13982,N_13799,N_13819);
or U13983 (N_13983,N_13868,N_13813);
xnor U13984 (N_13984,N_13830,N_13846);
nand U13985 (N_13985,N_13826,N_13783);
nand U13986 (N_13986,N_13753,N_13826);
or U13987 (N_13987,N_13848,N_13813);
xor U13988 (N_13988,N_13816,N_13858);
nor U13989 (N_13989,N_13805,N_13822);
nor U13990 (N_13990,N_13791,N_13768);
xor U13991 (N_13991,N_13753,N_13839);
xnor U13992 (N_13992,N_13841,N_13765);
nor U13993 (N_13993,N_13783,N_13750);
xor U13994 (N_13994,N_13798,N_13855);
xor U13995 (N_13995,N_13781,N_13841);
nand U13996 (N_13996,N_13862,N_13835);
or U13997 (N_13997,N_13791,N_13819);
and U13998 (N_13998,N_13870,N_13770);
xor U13999 (N_13999,N_13794,N_13807);
nor U14000 (N_14000,N_13993,N_13992);
and U14001 (N_14001,N_13917,N_13981);
nor U14002 (N_14002,N_13902,N_13911);
nor U14003 (N_14003,N_13878,N_13875);
xor U14004 (N_14004,N_13975,N_13988);
xor U14005 (N_14005,N_13966,N_13926);
nor U14006 (N_14006,N_13890,N_13983);
nand U14007 (N_14007,N_13901,N_13951);
nand U14008 (N_14008,N_13877,N_13896);
nand U14009 (N_14009,N_13893,N_13997);
xor U14010 (N_14010,N_13887,N_13944);
nor U14011 (N_14011,N_13996,N_13880);
nor U14012 (N_14012,N_13967,N_13977);
nand U14013 (N_14013,N_13956,N_13888);
and U14014 (N_14014,N_13908,N_13943);
and U14015 (N_14015,N_13980,N_13925);
nor U14016 (N_14016,N_13936,N_13960);
and U14017 (N_14017,N_13898,N_13892);
or U14018 (N_14018,N_13891,N_13919);
and U14019 (N_14019,N_13924,N_13986);
nor U14020 (N_14020,N_13939,N_13881);
nor U14021 (N_14021,N_13922,N_13894);
and U14022 (N_14022,N_13928,N_13954);
nor U14023 (N_14023,N_13950,N_13914);
nand U14024 (N_14024,N_13978,N_13923);
nor U14025 (N_14025,N_13903,N_13952);
nand U14026 (N_14026,N_13948,N_13945);
and U14027 (N_14027,N_13906,N_13886);
nor U14028 (N_14028,N_13985,N_13913);
nand U14029 (N_14029,N_13968,N_13969);
or U14030 (N_14030,N_13920,N_13889);
and U14031 (N_14031,N_13971,N_13912);
and U14032 (N_14032,N_13904,N_13937);
xnor U14033 (N_14033,N_13909,N_13883);
xor U14034 (N_14034,N_13905,N_13982);
nand U14035 (N_14035,N_13938,N_13907);
nand U14036 (N_14036,N_13984,N_13910);
or U14037 (N_14037,N_13929,N_13882);
or U14038 (N_14038,N_13972,N_13973);
nand U14039 (N_14039,N_13958,N_13884);
nor U14040 (N_14040,N_13940,N_13930);
or U14041 (N_14041,N_13942,N_13963);
or U14042 (N_14042,N_13932,N_13897);
nand U14043 (N_14043,N_13987,N_13931);
and U14044 (N_14044,N_13949,N_13899);
nand U14045 (N_14045,N_13970,N_13876);
xnor U14046 (N_14046,N_13916,N_13991);
nand U14047 (N_14047,N_13915,N_13941);
xor U14048 (N_14048,N_13961,N_13974);
nand U14049 (N_14049,N_13918,N_13979);
or U14050 (N_14050,N_13999,N_13895);
nand U14051 (N_14051,N_13927,N_13933);
nand U14052 (N_14052,N_13976,N_13879);
xor U14053 (N_14053,N_13900,N_13955);
and U14054 (N_14054,N_13994,N_13998);
and U14055 (N_14055,N_13990,N_13953);
or U14056 (N_14056,N_13965,N_13934);
and U14057 (N_14057,N_13957,N_13946);
or U14058 (N_14058,N_13959,N_13921);
or U14059 (N_14059,N_13962,N_13964);
or U14060 (N_14060,N_13995,N_13885);
and U14061 (N_14061,N_13947,N_13935);
xnor U14062 (N_14062,N_13989,N_13936);
xnor U14063 (N_14063,N_13876,N_13938);
and U14064 (N_14064,N_13924,N_13907);
nand U14065 (N_14065,N_13938,N_13951);
and U14066 (N_14066,N_13921,N_13926);
or U14067 (N_14067,N_13943,N_13975);
and U14068 (N_14068,N_13940,N_13879);
and U14069 (N_14069,N_13946,N_13915);
nand U14070 (N_14070,N_13920,N_13919);
nor U14071 (N_14071,N_13993,N_13996);
or U14072 (N_14072,N_13911,N_13901);
xnor U14073 (N_14073,N_13927,N_13959);
nor U14074 (N_14074,N_13972,N_13962);
and U14075 (N_14075,N_13906,N_13900);
nor U14076 (N_14076,N_13910,N_13999);
xnor U14077 (N_14077,N_13892,N_13972);
and U14078 (N_14078,N_13917,N_13907);
nor U14079 (N_14079,N_13952,N_13961);
nor U14080 (N_14080,N_13916,N_13971);
and U14081 (N_14081,N_13877,N_13961);
nor U14082 (N_14082,N_13962,N_13921);
and U14083 (N_14083,N_13879,N_13918);
nand U14084 (N_14084,N_13922,N_13959);
xor U14085 (N_14085,N_13927,N_13890);
and U14086 (N_14086,N_13967,N_13892);
nor U14087 (N_14087,N_13888,N_13995);
nor U14088 (N_14088,N_13940,N_13935);
or U14089 (N_14089,N_13886,N_13961);
or U14090 (N_14090,N_13877,N_13936);
or U14091 (N_14091,N_13970,N_13875);
and U14092 (N_14092,N_13931,N_13958);
or U14093 (N_14093,N_13948,N_13974);
and U14094 (N_14094,N_13923,N_13960);
or U14095 (N_14095,N_13974,N_13954);
xnor U14096 (N_14096,N_13876,N_13889);
or U14097 (N_14097,N_13905,N_13940);
nor U14098 (N_14098,N_13940,N_13972);
or U14099 (N_14099,N_13951,N_13982);
or U14100 (N_14100,N_13934,N_13877);
nor U14101 (N_14101,N_13909,N_13884);
xnor U14102 (N_14102,N_13901,N_13956);
and U14103 (N_14103,N_13988,N_13947);
xor U14104 (N_14104,N_13903,N_13899);
or U14105 (N_14105,N_13949,N_13979);
or U14106 (N_14106,N_13888,N_13920);
nand U14107 (N_14107,N_13960,N_13898);
or U14108 (N_14108,N_13929,N_13877);
or U14109 (N_14109,N_13975,N_13942);
and U14110 (N_14110,N_13904,N_13988);
nor U14111 (N_14111,N_13923,N_13974);
nor U14112 (N_14112,N_13918,N_13898);
nor U14113 (N_14113,N_13977,N_13988);
and U14114 (N_14114,N_13984,N_13917);
or U14115 (N_14115,N_13926,N_13918);
or U14116 (N_14116,N_13968,N_13882);
xnor U14117 (N_14117,N_13956,N_13927);
nor U14118 (N_14118,N_13975,N_13926);
or U14119 (N_14119,N_13929,N_13905);
nor U14120 (N_14120,N_13894,N_13885);
and U14121 (N_14121,N_13969,N_13974);
xnor U14122 (N_14122,N_13965,N_13897);
xnor U14123 (N_14123,N_13975,N_13913);
nor U14124 (N_14124,N_13982,N_13901);
nor U14125 (N_14125,N_14106,N_14088);
xnor U14126 (N_14126,N_14066,N_14037);
and U14127 (N_14127,N_14003,N_14072);
nand U14128 (N_14128,N_14043,N_14027);
or U14129 (N_14129,N_14019,N_14060);
xnor U14130 (N_14130,N_14046,N_14095);
xnor U14131 (N_14131,N_14102,N_14036);
xnor U14132 (N_14132,N_14111,N_14109);
xor U14133 (N_14133,N_14086,N_14098);
and U14134 (N_14134,N_14040,N_14114);
nor U14135 (N_14135,N_14052,N_14068);
xnor U14136 (N_14136,N_14108,N_14117);
nor U14137 (N_14137,N_14084,N_14023);
and U14138 (N_14138,N_14124,N_14085);
xnor U14139 (N_14139,N_14089,N_14034);
nand U14140 (N_14140,N_14122,N_14024);
nand U14141 (N_14141,N_14081,N_14025);
nor U14142 (N_14142,N_14011,N_14042);
and U14143 (N_14143,N_14035,N_14105);
nor U14144 (N_14144,N_14009,N_14041);
nand U14145 (N_14145,N_14064,N_14116);
and U14146 (N_14146,N_14073,N_14031);
or U14147 (N_14147,N_14000,N_14075);
and U14148 (N_14148,N_14110,N_14100);
nor U14149 (N_14149,N_14014,N_14058);
and U14150 (N_14150,N_14113,N_14006);
xnor U14151 (N_14151,N_14022,N_14033);
or U14152 (N_14152,N_14069,N_14047);
and U14153 (N_14153,N_14028,N_14056);
nor U14154 (N_14154,N_14120,N_14017);
nor U14155 (N_14155,N_14063,N_14032);
or U14156 (N_14156,N_14071,N_14078);
nand U14157 (N_14157,N_14079,N_14112);
nor U14158 (N_14158,N_14039,N_14065);
or U14159 (N_14159,N_14004,N_14044);
nor U14160 (N_14160,N_14107,N_14092);
nor U14161 (N_14161,N_14093,N_14061);
nor U14162 (N_14162,N_14118,N_14050);
nor U14163 (N_14163,N_14097,N_14059);
nand U14164 (N_14164,N_14103,N_14076);
nand U14165 (N_14165,N_14094,N_14074);
and U14166 (N_14166,N_14021,N_14018);
nor U14167 (N_14167,N_14099,N_14082);
and U14168 (N_14168,N_14070,N_14077);
xor U14169 (N_14169,N_14045,N_14001);
xnor U14170 (N_14170,N_14055,N_14062);
nor U14171 (N_14171,N_14013,N_14090);
or U14172 (N_14172,N_14051,N_14067);
xor U14173 (N_14173,N_14030,N_14007);
nand U14174 (N_14174,N_14104,N_14115);
nand U14175 (N_14175,N_14080,N_14012);
xor U14176 (N_14176,N_14010,N_14101);
and U14177 (N_14177,N_14015,N_14096);
nor U14178 (N_14178,N_14016,N_14049);
nor U14179 (N_14179,N_14053,N_14020);
nor U14180 (N_14180,N_14002,N_14123);
nand U14181 (N_14181,N_14057,N_14029);
xor U14182 (N_14182,N_14008,N_14087);
or U14183 (N_14183,N_14054,N_14119);
nand U14184 (N_14184,N_14005,N_14083);
nand U14185 (N_14185,N_14038,N_14026);
xnor U14186 (N_14186,N_14121,N_14048);
nand U14187 (N_14187,N_14091,N_14070);
nand U14188 (N_14188,N_14034,N_14009);
or U14189 (N_14189,N_14023,N_14054);
and U14190 (N_14190,N_14033,N_14113);
and U14191 (N_14191,N_14095,N_14042);
or U14192 (N_14192,N_14044,N_14033);
xor U14193 (N_14193,N_14089,N_14108);
xor U14194 (N_14194,N_14081,N_14066);
xnor U14195 (N_14195,N_14082,N_14002);
or U14196 (N_14196,N_14014,N_14027);
and U14197 (N_14197,N_14025,N_14000);
and U14198 (N_14198,N_14053,N_14042);
nor U14199 (N_14199,N_14065,N_14054);
and U14200 (N_14200,N_14096,N_14040);
xnor U14201 (N_14201,N_14060,N_14063);
xnor U14202 (N_14202,N_14099,N_14124);
or U14203 (N_14203,N_14082,N_14064);
xor U14204 (N_14204,N_14116,N_14016);
or U14205 (N_14205,N_14091,N_14079);
or U14206 (N_14206,N_14012,N_14098);
nand U14207 (N_14207,N_14023,N_14049);
nand U14208 (N_14208,N_14082,N_14026);
and U14209 (N_14209,N_14108,N_14019);
and U14210 (N_14210,N_14078,N_14059);
nand U14211 (N_14211,N_14071,N_14039);
nand U14212 (N_14212,N_14012,N_14014);
and U14213 (N_14213,N_14036,N_14065);
xor U14214 (N_14214,N_14012,N_14034);
or U14215 (N_14215,N_14091,N_14064);
and U14216 (N_14216,N_14121,N_14085);
nand U14217 (N_14217,N_14036,N_14080);
xor U14218 (N_14218,N_14100,N_14060);
nor U14219 (N_14219,N_14078,N_14097);
or U14220 (N_14220,N_14121,N_14007);
xor U14221 (N_14221,N_14083,N_14099);
and U14222 (N_14222,N_14054,N_14063);
and U14223 (N_14223,N_14011,N_14068);
or U14224 (N_14224,N_14022,N_14090);
nor U14225 (N_14225,N_14106,N_14014);
and U14226 (N_14226,N_14100,N_14084);
and U14227 (N_14227,N_14073,N_14100);
nor U14228 (N_14228,N_14013,N_14106);
xnor U14229 (N_14229,N_14052,N_14094);
nand U14230 (N_14230,N_14013,N_14043);
nor U14231 (N_14231,N_14041,N_14091);
nand U14232 (N_14232,N_14066,N_14053);
xor U14233 (N_14233,N_14005,N_14062);
nor U14234 (N_14234,N_14009,N_14003);
nand U14235 (N_14235,N_14124,N_14119);
nor U14236 (N_14236,N_14040,N_14074);
xor U14237 (N_14237,N_14082,N_14077);
or U14238 (N_14238,N_14019,N_14037);
nand U14239 (N_14239,N_14090,N_14066);
and U14240 (N_14240,N_14037,N_14111);
nor U14241 (N_14241,N_14058,N_14022);
or U14242 (N_14242,N_14117,N_14101);
and U14243 (N_14243,N_14035,N_14058);
xnor U14244 (N_14244,N_14124,N_14047);
and U14245 (N_14245,N_14061,N_14070);
or U14246 (N_14246,N_14097,N_14114);
nor U14247 (N_14247,N_14070,N_14022);
nand U14248 (N_14248,N_14077,N_14030);
nand U14249 (N_14249,N_14094,N_14077);
and U14250 (N_14250,N_14162,N_14217);
or U14251 (N_14251,N_14163,N_14233);
and U14252 (N_14252,N_14213,N_14142);
or U14253 (N_14253,N_14204,N_14199);
nand U14254 (N_14254,N_14237,N_14160);
and U14255 (N_14255,N_14170,N_14208);
or U14256 (N_14256,N_14143,N_14182);
or U14257 (N_14257,N_14235,N_14169);
nand U14258 (N_14258,N_14206,N_14165);
xor U14259 (N_14259,N_14212,N_14228);
xnor U14260 (N_14260,N_14152,N_14161);
or U14261 (N_14261,N_14234,N_14148);
and U14262 (N_14262,N_14242,N_14133);
xnor U14263 (N_14263,N_14175,N_14154);
xor U14264 (N_14264,N_14164,N_14211);
xnor U14265 (N_14265,N_14177,N_14136);
nand U14266 (N_14266,N_14202,N_14224);
nor U14267 (N_14267,N_14210,N_14195);
or U14268 (N_14268,N_14125,N_14178);
or U14269 (N_14269,N_14155,N_14138);
nor U14270 (N_14270,N_14127,N_14205);
nand U14271 (N_14271,N_14185,N_14215);
xnor U14272 (N_14272,N_14229,N_14227);
nand U14273 (N_14273,N_14158,N_14201);
nor U14274 (N_14274,N_14189,N_14172);
nand U14275 (N_14275,N_14140,N_14244);
or U14276 (N_14276,N_14187,N_14128);
and U14277 (N_14277,N_14139,N_14248);
nand U14278 (N_14278,N_14145,N_14222);
and U14279 (N_14279,N_14219,N_14176);
and U14280 (N_14280,N_14239,N_14173);
or U14281 (N_14281,N_14184,N_14153);
nor U14282 (N_14282,N_14156,N_14192);
xor U14283 (N_14283,N_14240,N_14246);
and U14284 (N_14284,N_14194,N_14198);
nand U14285 (N_14285,N_14238,N_14207);
and U14286 (N_14286,N_14157,N_14183);
and U14287 (N_14287,N_14221,N_14134);
xnor U14288 (N_14288,N_14146,N_14193);
or U14289 (N_14289,N_14191,N_14166);
nor U14290 (N_14290,N_14159,N_14231);
xnor U14291 (N_14291,N_14174,N_14179);
xnor U14292 (N_14292,N_14147,N_14132);
nor U14293 (N_14293,N_14190,N_14214);
or U14294 (N_14294,N_14232,N_14225);
nor U14295 (N_14295,N_14186,N_14188);
and U14296 (N_14296,N_14196,N_14137);
or U14297 (N_14297,N_14247,N_14131);
or U14298 (N_14298,N_14135,N_14168);
nor U14299 (N_14299,N_14200,N_14141);
nor U14300 (N_14300,N_14236,N_14151);
xnor U14301 (N_14301,N_14167,N_14150);
or U14302 (N_14302,N_14216,N_14180);
nor U14303 (N_14303,N_14209,N_14181);
or U14304 (N_14304,N_14149,N_14241);
nand U14305 (N_14305,N_14197,N_14203);
nor U14306 (N_14306,N_14230,N_14245);
and U14307 (N_14307,N_14223,N_14171);
and U14308 (N_14308,N_14218,N_14130);
xor U14309 (N_14309,N_14249,N_14220);
nand U14310 (N_14310,N_14126,N_14129);
nor U14311 (N_14311,N_14226,N_14144);
nor U14312 (N_14312,N_14243,N_14136);
or U14313 (N_14313,N_14128,N_14205);
or U14314 (N_14314,N_14241,N_14214);
nor U14315 (N_14315,N_14185,N_14167);
xnor U14316 (N_14316,N_14226,N_14156);
nand U14317 (N_14317,N_14184,N_14227);
xor U14318 (N_14318,N_14187,N_14245);
or U14319 (N_14319,N_14133,N_14136);
nor U14320 (N_14320,N_14165,N_14190);
xnor U14321 (N_14321,N_14242,N_14196);
or U14322 (N_14322,N_14195,N_14130);
and U14323 (N_14323,N_14204,N_14139);
xnor U14324 (N_14324,N_14208,N_14131);
nand U14325 (N_14325,N_14237,N_14233);
or U14326 (N_14326,N_14226,N_14242);
xnor U14327 (N_14327,N_14130,N_14166);
nand U14328 (N_14328,N_14170,N_14245);
nor U14329 (N_14329,N_14233,N_14126);
nand U14330 (N_14330,N_14129,N_14162);
nand U14331 (N_14331,N_14188,N_14168);
and U14332 (N_14332,N_14179,N_14164);
and U14333 (N_14333,N_14223,N_14129);
nand U14334 (N_14334,N_14203,N_14234);
xor U14335 (N_14335,N_14230,N_14201);
and U14336 (N_14336,N_14151,N_14176);
nand U14337 (N_14337,N_14197,N_14141);
and U14338 (N_14338,N_14230,N_14154);
xnor U14339 (N_14339,N_14187,N_14194);
nand U14340 (N_14340,N_14212,N_14223);
xor U14341 (N_14341,N_14197,N_14214);
xor U14342 (N_14342,N_14217,N_14226);
or U14343 (N_14343,N_14208,N_14211);
or U14344 (N_14344,N_14190,N_14232);
and U14345 (N_14345,N_14164,N_14153);
and U14346 (N_14346,N_14167,N_14135);
nor U14347 (N_14347,N_14126,N_14241);
nor U14348 (N_14348,N_14144,N_14146);
or U14349 (N_14349,N_14228,N_14179);
or U14350 (N_14350,N_14235,N_14248);
nand U14351 (N_14351,N_14246,N_14135);
and U14352 (N_14352,N_14196,N_14232);
and U14353 (N_14353,N_14221,N_14166);
xnor U14354 (N_14354,N_14194,N_14163);
nor U14355 (N_14355,N_14229,N_14211);
nand U14356 (N_14356,N_14198,N_14213);
xnor U14357 (N_14357,N_14165,N_14138);
nand U14358 (N_14358,N_14178,N_14181);
or U14359 (N_14359,N_14129,N_14198);
xor U14360 (N_14360,N_14164,N_14224);
nor U14361 (N_14361,N_14186,N_14237);
nand U14362 (N_14362,N_14152,N_14135);
nand U14363 (N_14363,N_14138,N_14193);
or U14364 (N_14364,N_14235,N_14158);
and U14365 (N_14365,N_14225,N_14167);
or U14366 (N_14366,N_14243,N_14152);
or U14367 (N_14367,N_14206,N_14139);
nor U14368 (N_14368,N_14215,N_14171);
and U14369 (N_14369,N_14221,N_14206);
or U14370 (N_14370,N_14213,N_14135);
xnor U14371 (N_14371,N_14226,N_14193);
nand U14372 (N_14372,N_14232,N_14145);
and U14373 (N_14373,N_14136,N_14209);
and U14374 (N_14374,N_14220,N_14201);
and U14375 (N_14375,N_14310,N_14361);
nand U14376 (N_14376,N_14366,N_14253);
and U14377 (N_14377,N_14345,N_14303);
nand U14378 (N_14378,N_14250,N_14285);
and U14379 (N_14379,N_14371,N_14286);
nor U14380 (N_14380,N_14355,N_14270);
nand U14381 (N_14381,N_14298,N_14331);
nor U14382 (N_14382,N_14322,N_14284);
xor U14383 (N_14383,N_14280,N_14306);
xnor U14384 (N_14384,N_14316,N_14269);
xnor U14385 (N_14385,N_14254,N_14255);
xnor U14386 (N_14386,N_14292,N_14334);
and U14387 (N_14387,N_14335,N_14300);
and U14388 (N_14388,N_14328,N_14343);
nand U14389 (N_14389,N_14260,N_14323);
and U14390 (N_14390,N_14266,N_14327);
and U14391 (N_14391,N_14281,N_14311);
xnor U14392 (N_14392,N_14329,N_14352);
and U14393 (N_14393,N_14305,N_14271);
or U14394 (N_14394,N_14337,N_14349);
xor U14395 (N_14395,N_14297,N_14291);
and U14396 (N_14396,N_14293,N_14353);
xnor U14397 (N_14397,N_14350,N_14273);
nor U14398 (N_14398,N_14276,N_14338);
nand U14399 (N_14399,N_14346,N_14364);
xnor U14400 (N_14400,N_14301,N_14360);
and U14401 (N_14401,N_14369,N_14272);
nor U14402 (N_14402,N_14330,N_14308);
and U14403 (N_14403,N_14319,N_14288);
nor U14404 (N_14404,N_14264,N_14356);
xnor U14405 (N_14405,N_14372,N_14374);
nor U14406 (N_14406,N_14370,N_14252);
nand U14407 (N_14407,N_14274,N_14296);
xnor U14408 (N_14408,N_14351,N_14283);
and U14409 (N_14409,N_14348,N_14268);
or U14410 (N_14410,N_14290,N_14367);
and U14411 (N_14411,N_14363,N_14258);
nor U14412 (N_14412,N_14262,N_14318);
and U14413 (N_14413,N_14321,N_14315);
and U14414 (N_14414,N_14314,N_14261);
xnor U14415 (N_14415,N_14295,N_14362);
nand U14416 (N_14416,N_14302,N_14275);
xor U14417 (N_14417,N_14251,N_14373);
or U14418 (N_14418,N_14307,N_14333);
xnor U14419 (N_14419,N_14336,N_14289);
xnor U14420 (N_14420,N_14309,N_14278);
nand U14421 (N_14421,N_14265,N_14359);
and U14422 (N_14422,N_14357,N_14257);
xor U14423 (N_14423,N_14332,N_14368);
nor U14424 (N_14424,N_14326,N_14324);
or U14425 (N_14425,N_14299,N_14277);
nor U14426 (N_14426,N_14325,N_14339);
nor U14427 (N_14427,N_14342,N_14358);
and U14428 (N_14428,N_14256,N_14347);
nand U14429 (N_14429,N_14312,N_14304);
nor U14430 (N_14430,N_14354,N_14279);
or U14431 (N_14431,N_14259,N_14320);
and U14432 (N_14432,N_14287,N_14344);
xnor U14433 (N_14433,N_14263,N_14267);
nor U14434 (N_14434,N_14282,N_14365);
nor U14435 (N_14435,N_14341,N_14313);
nor U14436 (N_14436,N_14340,N_14317);
xnor U14437 (N_14437,N_14294,N_14348);
nand U14438 (N_14438,N_14258,N_14361);
and U14439 (N_14439,N_14296,N_14340);
and U14440 (N_14440,N_14324,N_14348);
nand U14441 (N_14441,N_14266,N_14338);
nor U14442 (N_14442,N_14277,N_14303);
or U14443 (N_14443,N_14291,N_14303);
nor U14444 (N_14444,N_14295,N_14367);
or U14445 (N_14445,N_14277,N_14373);
xor U14446 (N_14446,N_14296,N_14363);
and U14447 (N_14447,N_14271,N_14303);
nand U14448 (N_14448,N_14371,N_14279);
nor U14449 (N_14449,N_14302,N_14361);
xor U14450 (N_14450,N_14339,N_14271);
and U14451 (N_14451,N_14307,N_14327);
xor U14452 (N_14452,N_14270,N_14279);
or U14453 (N_14453,N_14300,N_14314);
nor U14454 (N_14454,N_14321,N_14363);
nand U14455 (N_14455,N_14309,N_14348);
nand U14456 (N_14456,N_14273,N_14268);
xor U14457 (N_14457,N_14374,N_14296);
nand U14458 (N_14458,N_14306,N_14318);
xnor U14459 (N_14459,N_14315,N_14296);
nor U14460 (N_14460,N_14267,N_14348);
xor U14461 (N_14461,N_14335,N_14366);
xnor U14462 (N_14462,N_14367,N_14278);
nand U14463 (N_14463,N_14314,N_14359);
or U14464 (N_14464,N_14349,N_14322);
and U14465 (N_14465,N_14285,N_14357);
xor U14466 (N_14466,N_14304,N_14369);
xnor U14467 (N_14467,N_14312,N_14357);
xnor U14468 (N_14468,N_14263,N_14303);
nor U14469 (N_14469,N_14302,N_14265);
xor U14470 (N_14470,N_14343,N_14268);
nor U14471 (N_14471,N_14326,N_14269);
or U14472 (N_14472,N_14358,N_14260);
nand U14473 (N_14473,N_14312,N_14303);
or U14474 (N_14474,N_14254,N_14340);
xnor U14475 (N_14475,N_14287,N_14369);
and U14476 (N_14476,N_14297,N_14327);
and U14477 (N_14477,N_14285,N_14362);
and U14478 (N_14478,N_14297,N_14360);
or U14479 (N_14479,N_14367,N_14315);
nand U14480 (N_14480,N_14357,N_14279);
nand U14481 (N_14481,N_14263,N_14259);
nor U14482 (N_14482,N_14371,N_14253);
nand U14483 (N_14483,N_14280,N_14366);
nand U14484 (N_14484,N_14335,N_14352);
or U14485 (N_14485,N_14312,N_14279);
nand U14486 (N_14486,N_14333,N_14320);
and U14487 (N_14487,N_14339,N_14278);
and U14488 (N_14488,N_14270,N_14325);
nand U14489 (N_14489,N_14355,N_14357);
xor U14490 (N_14490,N_14321,N_14371);
and U14491 (N_14491,N_14361,N_14344);
nand U14492 (N_14492,N_14257,N_14266);
and U14493 (N_14493,N_14333,N_14362);
xor U14494 (N_14494,N_14274,N_14261);
and U14495 (N_14495,N_14274,N_14255);
xor U14496 (N_14496,N_14310,N_14343);
nor U14497 (N_14497,N_14328,N_14331);
or U14498 (N_14498,N_14330,N_14316);
and U14499 (N_14499,N_14355,N_14363);
nor U14500 (N_14500,N_14398,N_14414);
nor U14501 (N_14501,N_14421,N_14494);
nor U14502 (N_14502,N_14420,N_14472);
nand U14503 (N_14503,N_14385,N_14445);
and U14504 (N_14504,N_14430,N_14479);
nor U14505 (N_14505,N_14489,N_14426);
nand U14506 (N_14506,N_14419,N_14463);
and U14507 (N_14507,N_14418,N_14381);
and U14508 (N_14508,N_14412,N_14496);
and U14509 (N_14509,N_14406,N_14485);
xor U14510 (N_14510,N_14393,N_14492);
or U14511 (N_14511,N_14391,N_14447);
xnor U14512 (N_14512,N_14399,N_14411);
or U14513 (N_14513,N_14495,N_14466);
nor U14514 (N_14514,N_14481,N_14439);
and U14515 (N_14515,N_14467,N_14490);
and U14516 (N_14516,N_14386,N_14474);
nor U14517 (N_14517,N_14395,N_14498);
nor U14518 (N_14518,N_14440,N_14422);
or U14519 (N_14519,N_14459,N_14401);
and U14520 (N_14520,N_14499,N_14497);
nor U14521 (N_14521,N_14377,N_14450);
or U14522 (N_14522,N_14407,N_14375);
nand U14523 (N_14523,N_14392,N_14464);
nor U14524 (N_14524,N_14473,N_14390);
nand U14525 (N_14525,N_14409,N_14442);
or U14526 (N_14526,N_14451,N_14404);
nand U14527 (N_14527,N_14475,N_14470);
nor U14528 (N_14528,N_14413,N_14455);
nor U14529 (N_14529,N_14482,N_14376);
nand U14530 (N_14530,N_14471,N_14437);
xnor U14531 (N_14531,N_14394,N_14428);
xor U14532 (N_14532,N_14405,N_14378);
nor U14533 (N_14533,N_14478,N_14432);
and U14534 (N_14534,N_14462,N_14434);
xor U14535 (N_14535,N_14410,N_14427);
or U14536 (N_14536,N_14446,N_14436);
and U14537 (N_14537,N_14469,N_14480);
xnor U14538 (N_14538,N_14382,N_14441);
nand U14539 (N_14539,N_14443,N_14477);
nand U14540 (N_14540,N_14408,N_14415);
nand U14541 (N_14541,N_14433,N_14487);
xor U14542 (N_14542,N_14454,N_14380);
and U14543 (N_14543,N_14402,N_14461);
nor U14544 (N_14544,N_14429,N_14488);
nand U14545 (N_14545,N_14396,N_14493);
or U14546 (N_14546,N_14400,N_14465);
or U14547 (N_14547,N_14423,N_14384);
and U14548 (N_14548,N_14460,N_14424);
xnor U14549 (N_14549,N_14458,N_14476);
nand U14550 (N_14550,N_14456,N_14416);
nand U14551 (N_14551,N_14448,N_14444);
and U14552 (N_14552,N_14484,N_14468);
and U14553 (N_14553,N_14452,N_14486);
or U14554 (N_14554,N_14438,N_14403);
nor U14555 (N_14555,N_14379,N_14457);
and U14556 (N_14556,N_14383,N_14417);
nand U14557 (N_14557,N_14388,N_14449);
nor U14558 (N_14558,N_14389,N_14491);
nand U14559 (N_14559,N_14483,N_14453);
or U14560 (N_14560,N_14431,N_14397);
nand U14561 (N_14561,N_14435,N_14425);
nand U14562 (N_14562,N_14387,N_14495);
xor U14563 (N_14563,N_14390,N_14447);
and U14564 (N_14564,N_14421,N_14450);
and U14565 (N_14565,N_14400,N_14408);
and U14566 (N_14566,N_14451,N_14420);
nor U14567 (N_14567,N_14419,N_14492);
and U14568 (N_14568,N_14434,N_14454);
xor U14569 (N_14569,N_14488,N_14483);
xor U14570 (N_14570,N_14378,N_14393);
nor U14571 (N_14571,N_14480,N_14434);
or U14572 (N_14572,N_14420,N_14381);
or U14573 (N_14573,N_14467,N_14404);
xor U14574 (N_14574,N_14385,N_14379);
or U14575 (N_14575,N_14426,N_14376);
xor U14576 (N_14576,N_14418,N_14445);
nand U14577 (N_14577,N_14459,N_14387);
xnor U14578 (N_14578,N_14401,N_14405);
and U14579 (N_14579,N_14381,N_14470);
nor U14580 (N_14580,N_14489,N_14467);
nor U14581 (N_14581,N_14408,N_14484);
or U14582 (N_14582,N_14496,N_14435);
xor U14583 (N_14583,N_14423,N_14485);
nand U14584 (N_14584,N_14418,N_14428);
nand U14585 (N_14585,N_14454,N_14413);
xor U14586 (N_14586,N_14395,N_14457);
nor U14587 (N_14587,N_14400,N_14432);
or U14588 (N_14588,N_14393,N_14422);
nor U14589 (N_14589,N_14417,N_14479);
and U14590 (N_14590,N_14398,N_14465);
nand U14591 (N_14591,N_14420,N_14498);
nor U14592 (N_14592,N_14464,N_14405);
nor U14593 (N_14593,N_14472,N_14494);
or U14594 (N_14594,N_14401,N_14470);
and U14595 (N_14595,N_14457,N_14491);
xnor U14596 (N_14596,N_14387,N_14409);
xor U14597 (N_14597,N_14414,N_14434);
or U14598 (N_14598,N_14380,N_14427);
xnor U14599 (N_14599,N_14379,N_14383);
xnor U14600 (N_14600,N_14496,N_14491);
or U14601 (N_14601,N_14396,N_14390);
or U14602 (N_14602,N_14375,N_14480);
or U14603 (N_14603,N_14466,N_14426);
xor U14604 (N_14604,N_14485,N_14457);
xnor U14605 (N_14605,N_14404,N_14469);
and U14606 (N_14606,N_14403,N_14375);
xor U14607 (N_14607,N_14492,N_14391);
and U14608 (N_14608,N_14446,N_14459);
xor U14609 (N_14609,N_14467,N_14408);
nor U14610 (N_14610,N_14399,N_14435);
xor U14611 (N_14611,N_14404,N_14491);
xnor U14612 (N_14612,N_14491,N_14420);
xor U14613 (N_14613,N_14425,N_14416);
nand U14614 (N_14614,N_14376,N_14392);
nand U14615 (N_14615,N_14494,N_14392);
or U14616 (N_14616,N_14415,N_14401);
nor U14617 (N_14617,N_14428,N_14407);
nor U14618 (N_14618,N_14400,N_14427);
nor U14619 (N_14619,N_14445,N_14379);
nor U14620 (N_14620,N_14455,N_14421);
nor U14621 (N_14621,N_14388,N_14390);
nand U14622 (N_14622,N_14388,N_14440);
or U14623 (N_14623,N_14454,N_14495);
or U14624 (N_14624,N_14377,N_14393);
or U14625 (N_14625,N_14516,N_14559);
and U14626 (N_14626,N_14517,N_14565);
nor U14627 (N_14627,N_14608,N_14612);
xor U14628 (N_14628,N_14503,N_14539);
and U14629 (N_14629,N_14561,N_14550);
nor U14630 (N_14630,N_14577,N_14569);
or U14631 (N_14631,N_14578,N_14515);
nor U14632 (N_14632,N_14568,N_14560);
nor U14633 (N_14633,N_14573,N_14620);
and U14634 (N_14634,N_14596,N_14558);
and U14635 (N_14635,N_14556,N_14501);
nor U14636 (N_14636,N_14521,N_14604);
xor U14637 (N_14637,N_14532,N_14609);
nand U14638 (N_14638,N_14555,N_14504);
nand U14639 (N_14639,N_14616,N_14520);
nand U14640 (N_14640,N_14571,N_14621);
nand U14641 (N_14641,N_14584,N_14524);
or U14642 (N_14642,N_14614,N_14528);
and U14643 (N_14643,N_14522,N_14570);
and U14644 (N_14644,N_14598,N_14576);
xor U14645 (N_14645,N_14589,N_14533);
nand U14646 (N_14646,N_14563,N_14567);
xor U14647 (N_14647,N_14557,N_14518);
and U14648 (N_14648,N_14549,N_14613);
nand U14649 (N_14649,N_14583,N_14574);
nor U14650 (N_14650,N_14538,N_14602);
xnor U14651 (N_14651,N_14509,N_14500);
and U14652 (N_14652,N_14552,N_14605);
nand U14653 (N_14653,N_14548,N_14588);
and U14654 (N_14654,N_14553,N_14601);
and U14655 (N_14655,N_14600,N_14511);
nand U14656 (N_14656,N_14530,N_14527);
nand U14657 (N_14657,N_14606,N_14512);
and U14658 (N_14658,N_14531,N_14513);
xnor U14659 (N_14659,N_14547,N_14542);
or U14660 (N_14660,N_14525,N_14590);
nor U14661 (N_14661,N_14541,N_14610);
nand U14662 (N_14662,N_14566,N_14523);
and U14663 (N_14663,N_14505,N_14595);
or U14664 (N_14664,N_14599,N_14607);
or U14665 (N_14665,N_14535,N_14617);
nor U14666 (N_14666,N_14510,N_14585);
nor U14667 (N_14667,N_14575,N_14546);
nand U14668 (N_14668,N_14580,N_14507);
nand U14669 (N_14669,N_14623,N_14579);
and U14670 (N_14670,N_14587,N_14562);
xnor U14671 (N_14671,N_14611,N_14537);
and U14672 (N_14672,N_14545,N_14591);
nand U14673 (N_14673,N_14615,N_14514);
and U14674 (N_14674,N_14506,N_14624);
nor U14675 (N_14675,N_14581,N_14582);
and U14676 (N_14676,N_14618,N_14519);
nor U14677 (N_14677,N_14536,N_14502);
and U14678 (N_14678,N_14593,N_14554);
or U14679 (N_14679,N_14544,N_14540);
nand U14680 (N_14680,N_14594,N_14508);
or U14681 (N_14681,N_14534,N_14526);
or U14682 (N_14682,N_14551,N_14586);
nor U14683 (N_14683,N_14619,N_14592);
nand U14684 (N_14684,N_14564,N_14572);
nor U14685 (N_14685,N_14603,N_14597);
xor U14686 (N_14686,N_14622,N_14529);
and U14687 (N_14687,N_14543,N_14615);
or U14688 (N_14688,N_14574,N_14538);
nand U14689 (N_14689,N_14500,N_14590);
nor U14690 (N_14690,N_14510,N_14561);
nor U14691 (N_14691,N_14514,N_14585);
and U14692 (N_14692,N_14603,N_14571);
nor U14693 (N_14693,N_14616,N_14589);
and U14694 (N_14694,N_14618,N_14522);
xnor U14695 (N_14695,N_14584,N_14599);
and U14696 (N_14696,N_14585,N_14624);
and U14697 (N_14697,N_14513,N_14525);
nand U14698 (N_14698,N_14550,N_14590);
nor U14699 (N_14699,N_14623,N_14514);
and U14700 (N_14700,N_14535,N_14573);
nor U14701 (N_14701,N_14588,N_14590);
xnor U14702 (N_14702,N_14532,N_14551);
or U14703 (N_14703,N_14582,N_14536);
nor U14704 (N_14704,N_14612,N_14526);
nor U14705 (N_14705,N_14590,N_14506);
or U14706 (N_14706,N_14561,N_14622);
and U14707 (N_14707,N_14516,N_14591);
nand U14708 (N_14708,N_14528,N_14514);
nor U14709 (N_14709,N_14590,N_14577);
nor U14710 (N_14710,N_14536,N_14623);
nor U14711 (N_14711,N_14595,N_14549);
xnor U14712 (N_14712,N_14509,N_14610);
nand U14713 (N_14713,N_14544,N_14606);
and U14714 (N_14714,N_14604,N_14532);
or U14715 (N_14715,N_14515,N_14588);
nor U14716 (N_14716,N_14609,N_14522);
xor U14717 (N_14717,N_14532,N_14531);
nand U14718 (N_14718,N_14528,N_14529);
or U14719 (N_14719,N_14558,N_14623);
or U14720 (N_14720,N_14597,N_14592);
nand U14721 (N_14721,N_14618,N_14617);
xnor U14722 (N_14722,N_14514,N_14532);
or U14723 (N_14723,N_14543,N_14514);
nand U14724 (N_14724,N_14591,N_14550);
nor U14725 (N_14725,N_14609,N_14619);
xor U14726 (N_14726,N_14583,N_14571);
nand U14727 (N_14727,N_14561,N_14506);
nor U14728 (N_14728,N_14505,N_14597);
nand U14729 (N_14729,N_14620,N_14568);
xnor U14730 (N_14730,N_14585,N_14543);
or U14731 (N_14731,N_14615,N_14613);
nand U14732 (N_14732,N_14597,N_14535);
or U14733 (N_14733,N_14592,N_14502);
xnor U14734 (N_14734,N_14545,N_14558);
nor U14735 (N_14735,N_14621,N_14545);
or U14736 (N_14736,N_14551,N_14621);
nor U14737 (N_14737,N_14505,N_14527);
nor U14738 (N_14738,N_14567,N_14606);
xor U14739 (N_14739,N_14579,N_14609);
or U14740 (N_14740,N_14545,N_14575);
or U14741 (N_14741,N_14614,N_14600);
xnor U14742 (N_14742,N_14509,N_14512);
nor U14743 (N_14743,N_14500,N_14600);
nand U14744 (N_14744,N_14571,N_14584);
and U14745 (N_14745,N_14595,N_14616);
and U14746 (N_14746,N_14580,N_14512);
or U14747 (N_14747,N_14624,N_14526);
xor U14748 (N_14748,N_14621,N_14538);
xor U14749 (N_14749,N_14500,N_14617);
nor U14750 (N_14750,N_14747,N_14663);
or U14751 (N_14751,N_14717,N_14665);
nor U14752 (N_14752,N_14642,N_14728);
nand U14753 (N_14753,N_14742,N_14690);
and U14754 (N_14754,N_14704,N_14645);
xor U14755 (N_14755,N_14748,N_14653);
xor U14756 (N_14756,N_14701,N_14672);
or U14757 (N_14757,N_14629,N_14686);
nor U14758 (N_14758,N_14678,N_14698);
and U14759 (N_14759,N_14721,N_14711);
or U14760 (N_14760,N_14627,N_14716);
nor U14761 (N_14761,N_14709,N_14705);
or U14762 (N_14762,N_14730,N_14676);
nand U14763 (N_14763,N_14710,N_14659);
xor U14764 (N_14764,N_14666,N_14682);
or U14765 (N_14765,N_14700,N_14719);
nand U14766 (N_14766,N_14648,N_14674);
nor U14767 (N_14767,N_14675,N_14688);
and U14768 (N_14768,N_14691,N_14743);
xnor U14769 (N_14769,N_14727,N_14737);
xor U14770 (N_14770,N_14685,N_14637);
or U14771 (N_14771,N_14706,N_14702);
and U14772 (N_14772,N_14712,N_14630);
nand U14773 (N_14773,N_14739,N_14673);
xor U14774 (N_14774,N_14655,N_14651);
and U14775 (N_14775,N_14646,N_14632);
nor U14776 (N_14776,N_14699,N_14631);
nand U14777 (N_14777,N_14635,N_14692);
nor U14778 (N_14778,N_14724,N_14720);
nand U14779 (N_14779,N_14677,N_14654);
xor U14780 (N_14780,N_14734,N_14625);
nor U14781 (N_14781,N_14650,N_14643);
or U14782 (N_14782,N_14644,N_14715);
nand U14783 (N_14783,N_14729,N_14733);
nor U14784 (N_14784,N_14664,N_14722);
and U14785 (N_14785,N_14696,N_14639);
nor U14786 (N_14786,N_14660,N_14723);
or U14787 (N_14787,N_14670,N_14687);
and U14788 (N_14788,N_14647,N_14640);
xor U14789 (N_14789,N_14735,N_14638);
or U14790 (N_14790,N_14740,N_14626);
or U14791 (N_14791,N_14746,N_14671);
nand U14792 (N_14792,N_14628,N_14732);
or U14793 (N_14793,N_14636,N_14658);
xnor U14794 (N_14794,N_14683,N_14694);
or U14795 (N_14795,N_14652,N_14725);
and U14796 (N_14796,N_14669,N_14741);
and U14797 (N_14797,N_14703,N_14649);
nor U14798 (N_14798,N_14641,N_14714);
nand U14799 (N_14799,N_14738,N_14634);
and U14800 (N_14800,N_14693,N_14726);
nand U14801 (N_14801,N_14689,N_14684);
xor U14802 (N_14802,N_14662,N_14745);
and U14803 (N_14803,N_14718,N_14656);
nand U14804 (N_14804,N_14749,N_14679);
nand U14805 (N_14805,N_14713,N_14667);
xor U14806 (N_14806,N_14633,N_14657);
or U14807 (N_14807,N_14707,N_14697);
xor U14808 (N_14808,N_14708,N_14681);
xnor U14809 (N_14809,N_14668,N_14736);
xor U14810 (N_14810,N_14680,N_14744);
nor U14811 (N_14811,N_14695,N_14731);
nand U14812 (N_14812,N_14661,N_14650);
or U14813 (N_14813,N_14742,N_14669);
nor U14814 (N_14814,N_14747,N_14635);
and U14815 (N_14815,N_14634,N_14644);
nor U14816 (N_14816,N_14738,N_14648);
xor U14817 (N_14817,N_14649,N_14715);
and U14818 (N_14818,N_14739,N_14642);
xor U14819 (N_14819,N_14625,N_14708);
xnor U14820 (N_14820,N_14671,N_14719);
or U14821 (N_14821,N_14632,N_14682);
nand U14822 (N_14822,N_14640,N_14625);
nand U14823 (N_14823,N_14696,N_14642);
nand U14824 (N_14824,N_14702,N_14672);
nor U14825 (N_14825,N_14728,N_14718);
and U14826 (N_14826,N_14748,N_14693);
or U14827 (N_14827,N_14713,N_14741);
or U14828 (N_14828,N_14644,N_14665);
nand U14829 (N_14829,N_14657,N_14654);
or U14830 (N_14830,N_14627,N_14719);
or U14831 (N_14831,N_14748,N_14674);
nand U14832 (N_14832,N_14664,N_14628);
and U14833 (N_14833,N_14627,N_14713);
or U14834 (N_14834,N_14635,N_14652);
nand U14835 (N_14835,N_14697,N_14667);
or U14836 (N_14836,N_14656,N_14674);
or U14837 (N_14837,N_14702,N_14734);
nand U14838 (N_14838,N_14642,N_14746);
or U14839 (N_14839,N_14712,N_14629);
nand U14840 (N_14840,N_14669,N_14688);
nor U14841 (N_14841,N_14685,N_14684);
nor U14842 (N_14842,N_14677,N_14706);
nor U14843 (N_14843,N_14659,N_14664);
nand U14844 (N_14844,N_14687,N_14664);
xnor U14845 (N_14845,N_14641,N_14741);
and U14846 (N_14846,N_14650,N_14631);
xnor U14847 (N_14847,N_14695,N_14662);
xor U14848 (N_14848,N_14644,N_14737);
and U14849 (N_14849,N_14723,N_14625);
or U14850 (N_14850,N_14682,N_14669);
nor U14851 (N_14851,N_14741,N_14727);
nor U14852 (N_14852,N_14697,N_14677);
nor U14853 (N_14853,N_14648,N_14707);
nor U14854 (N_14854,N_14633,N_14655);
xor U14855 (N_14855,N_14674,N_14743);
xor U14856 (N_14856,N_14697,N_14647);
xor U14857 (N_14857,N_14731,N_14656);
nor U14858 (N_14858,N_14638,N_14627);
nor U14859 (N_14859,N_14701,N_14719);
nand U14860 (N_14860,N_14685,N_14749);
or U14861 (N_14861,N_14739,N_14684);
and U14862 (N_14862,N_14729,N_14652);
nor U14863 (N_14863,N_14682,N_14626);
and U14864 (N_14864,N_14734,N_14689);
and U14865 (N_14865,N_14671,N_14729);
nor U14866 (N_14866,N_14675,N_14632);
xnor U14867 (N_14867,N_14695,N_14677);
xor U14868 (N_14868,N_14666,N_14689);
nor U14869 (N_14869,N_14666,N_14630);
and U14870 (N_14870,N_14721,N_14641);
nor U14871 (N_14871,N_14741,N_14635);
or U14872 (N_14872,N_14628,N_14631);
and U14873 (N_14873,N_14636,N_14641);
nand U14874 (N_14874,N_14663,N_14670);
xor U14875 (N_14875,N_14873,N_14806);
nor U14876 (N_14876,N_14781,N_14761);
or U14877 (N_14877,N_14790,N_14858);
xnor U14878 (N_14878,N_14778,N_14773);
xnor U14879 (N_14879,N_14839,N_14819);
xnor U14880 (N_14880,N_14789,N_14857);
nor U14881 (N_14881,N_14853,N_14808);
and U14882 (N_14882,N_14829,N_14838);
xnor U14883 (N_14883,N_14792,N_14787);
nor U14884 (N_14884,N_14834,N_14764);
nand U14885 (N_14885,N_14804,N_14822);
and U14886 (N_14886,N_14774,N_14862);
or U14887 (N_14887,N_14813,N_14828);
nor U14888 (N_14888,N_14840,N_14771);
or U14889 (N_14889,N_14831,N_14807);
or U14890 (N_14890,N_14805,N_14768);
nor U14891 (N_14891,N_14785,N_14802);
nand U14892 (N_14892,N_14752,N_14765);
and U14893 (N_14893,N_14824,N_14796);
or U14894 (N_14894,N_14830,N_14863);
xnor U14895 (N_14895,N_14793,N_14815);
or U14896 (N_14896,N_14810,N_14860);
xnor U14897 (N_14897,N_14842,N_14850);
or U14898 (N_14898,N_14855,N_14820);
or U14899 (N_14899,N_14835,N_14788);
xnor U14900 (N_14900,N_14870,N_14868);
and U14901 (N_14901,N_14811,N_14803);
nand U14902 (N_14902,N_14758,N_14864);
and U14903 (N_14903,N_14756,N_14812);
nand U14904 (N_14904,N_14776,N_14872);
or U14905 (N_14905,N_14800,N_14851);
nor U14906 (N_14906,N_14801,N_14780);
nor U14907 (N_14907,N_14825,N_14844);
and U14908 (N_14908,N_14823,N_14854);
and U14909 (N_14909,N_14799,N_14762);
nand U14910 (N_14910,N_14757,N_14843);
nand U14911 (N_14911,N_14755,N_14861);
or U14912 (N_14912,N_14777,N_14772);
nand U14913 (N_14913,N_14809,N_14874);
nor U14914 (N_14914,N_14763,N_14841);
xnor U14915 (N_14915,N_14852,N_14786);
or U14916 (N_14916,N_14782,N_14856);
nand U14917 (N_14917,N_14848,N_14816);
nand U14918 (N_14918,N_14817,N_14759);
nand U14919 (N_14919,N_14770,N_14871);
xor U14920 (N_14920,N_14836,N_14798);
nand U14921 (N_14921,N_14795,N_14775);
or U14922 (N_14922,N_14769,N_14754);
xnor U14923 (N_14923,N_14784,N_14869);
nand U14924 (N_14924,N_14753,N_14750);
or U14925 (N_14925,N_14767,N_14814);
nor U14926 (N_14926,N_14783,N_14833);
nand U14927 (N_14927,N_14865,N_14818);
xnor U14928 (N_14928,N_14766,N_14751);
xor U14929 (N_14929,N_14791,N_14866);
nand U14930 (N_14930,N_14827,N_14832);
and U14931 (N_14931,N_14847,N_14779);
xnor U14932 (N_14932,N_14837,N_14845);
xnor U14933 (N_14933,N_14846,N_14760);
nor U14934 (N_14934,N_14867,N_14859);
nor U14935 (N_14935,N_14849,N_14821);
nor U14936 (N_14936,N_14794,N_14797);
and U14937 (N_14937,N_14826,N_14813);
nand U14938 (N_14938,N_14800,N_14808);
and U14939 (N_14939,N_14829,N_14855);
and U14940 (N_14940,N_14780,N_14779);
or U14941 (N_14941,N_14843,N_14803);
xor U14942 (N_14942,N_14864,N_14854);
xor U14943 (N_14943,N_14819,N_14786);
and U14944 (N_14944,N_14841,N_14872);
or U14945 (N_14945,N_14764,N_14781);
or U14946 (N_14946,N_14785,N_14825);
or U14947 (N_14947,N_14835,N_14828);
or U14948 (N_14948,N_14867,N_14841);
and U14949 (N_14949,N_14811,N_14849);
nand U14950 (N_14950,N_14862,N_14758);
nor U14951 (N_14951,N_14834,N_14825);
nand U14952 (N_14952,N_14859,N_14836);
xor U14953 (N_14953,N_14807,N_14791);
xor U14954 (N_14954,N_14808,N_14772);
nor U14955 (N_14955,N_14809,N_14841);
or U14956 (N_14956,N_14826,N_14808);
xnor U14957 (N_14957,N_14779,N_14870);
nor U14958 (N_14958,N_14765,N_14841);
nor U14959 (N_14959,N_14855,N_14755);
and U14960 (N_14960,N_14865,N_14751);
nand U14961 (N_14961,N_14778,N_14762);
nand U14962 (N_14962,N_14793,N_14832);
nand U14963 (N_14963,N_14803,N_14853);
or U14964 (N_14964,N_14841,N_14787);
nor U14965 (N_14965,N_14799,N_14848);
xor U14966 (N_14966,N_14792,N_14833);
nand U14967 (N_14967,N_14842,N_14859);
xor U14968 (N_14968,N_14751,N_14789);
or U14969 (N_14969,N_14773,N_14844);
nand U14970 (N_14970,N_14789,N_14800);
nor U14971 (N_14971,N_14756,N_14750);
xor U14972 (N_14972,N_14811,N_14752);
nor U14973 (N_14973,N_14807,N_14862);
or U14974 (N_14974,N_14840,N_14859);
xor U14975 (N_14975,N_14782,N_14822);
nor U14976 (N_14976,N_14801,N_14841);
nand U14977 (N_14977,N_14756,N_14774);
nand U14978 (N_14978,N_14816,N_14756);
or U14979 (N_14979,N_14842,N_14829);
nor U14980 (N_14980,N_14824,N_14851);
nor U14981 (N_14981,N_14822,N_14868);
nor U14982 (N_14982,N_14783,N_14771);
or U14983 (N_14983,N_14779,N_14831);
or U14984 (N_14984,N_14816,N_14872);
nor U14985 (N_14985,N_14752,N_14841);
xor U14986 (N_14986,N_14801,N_14819);
nand U14987 (N_14987,N_14752,N_14756);
nor U14988 (N_14988,N_14848,N_14755);
xnor U14989 (N_14989,N_14836,N_14797);
nor U14990 (N_14990,N_14871,N_14788);
and U14991 (N_14991,N_14758,N_14823);
nor U14992 (N_14992,N_14849,N_14874);
nor U14993 (N_14993,N_14856,N_14821);
or U14994 (N_14994,N_14753,N_14863);
nor U14995 (N_14995,N_14764,N_14840);
and U14996 (N_14996,N_14754,N_14849);
and U14997 (N_14997,N_14762,N_14812);
nand U14998 (N_14998,N_14759,N_14756);
xnor U14999 (N_14999,N_14755,N_14813);
or UO_0 (O_0,N_14924,N_14878);
or UO_1 (O_1,N_14949,N_14976);
and UO_2 (O_2,N_14894,N_14967);
or UO_3 (O_3,N_14985,N_14981);
nand UO_4 (O_4,N_14897,N_14944);
nor UO_5 (O_5,N_14912,N_14956);
nor UO_6 (O_6,N_14896,N_14902);
and UO_7 (O_7,N_14990,N_14950);
nand UO_8 (O_8,N_14887,N_14995);
nand UO_9 (O_9,N_14997,N_14921);
xnor UO_10 (O_10,N_14890,N_14983);
or UO_11 (O_11,N_14938,N_14946);
and UO_12 (O_12,N_14885,N_14920);
xnor UO_13 (O_13,N_14988,N_14982);
nor UO_14 (O_14,N_14906,N_14891);
or UO_15 (O_15,N_14909,N_14880);
nand UO_16 (O_16,N_14927,N_14966);
xor UO_17 (O_17,N_14994,N_14971);
or UO_18 (O_18,N_14952,N_14913);
nand UO_19 (O_19,N_14934,N_14953);
xor UO_20 (O_20,N_14964,N_14963);
nor UO_21 (O_21,N_14892,N_14879);
nor UO_22 (O_22,N_14926,N_14875);
xor UO_23 (O_23,N_14889,N_14992);
xor UO_24 (O_24,N_14961,N_14914);
nand UO_25 (O_25,N_14908,N_14960);
and UO_26 (O_26,N_14905,N_14939);
xor UO_27 (O_27,N_14987,N_14947);
nor UO_28 (O_28,N_14991,N_14907);
xor UO_29 (O_29,N_14959,N_14957);
nand UO_30 (O_30,N_14942,N_14936);
nand UO_31 (O_31,N_14911,N_14888);
xnor UO_32 (O_32,N_14900,N_14999);
and UO_33 (O_33,N_14901,N_14965);
nand UO_34 (O_34,N_14923,N_14979);
nor UO_35 (O_35,N_14932,N_14882);
and UO_36 (O_36,N_14883,N_14916);
nand UO_37 (O_37,N_14929,N_14922);
nor UO_38 (O_38,N_14931,N_14954);
nand UO_39 (O_39,N_14917,N_14975);
xnor UO_40 (O_40,N_14903,N_14893);
and UO_41 (O_41,N_14970,N_14881);
and UO_42 (O_42,N_14940,N_14996);
nor UO_43 (O_43,N_14877,N_14969);
and UO_44 (O_44,N_14943,N_14904);
nor UO_45 (O_45,N_14977,N_14986);
or UO_46 (O_46,N_14918,N_14973);
xor UO_47 (O_47,N_14958,N_14895);
nand UO_48 (O_48,N_14993,N_14968);
nor UO_49 (O_49,N_14962,N_14935);
xor UO_50 (O_50,N_14886,N_14948);
nand UO_51 (O_51,N_14980,N_14915);
and UO_52 (O_52,N_14925,N_14984);
nor UO_53 (O_53,N_14876,N_14972);
or UO_54 (O_54,N_14884,N_14937);
and UO_55 (O_55,N_14998,N_14989);
or UO_56 (O_56,N_14941,N_14955);
or UO_57 (O_57,N_14974,N_14898);
and UO_58 (O_58,N_14910,N_14928);
nor UO_59 (O_59,N_14945,N_14951);
nor UO_60 (O_60,N_14919,N_14933);
nand UO_61 (O_61,N_14930,N_14978);
and UO_62 (O_62,N_14899,N_14974);
nor UO_63 (O_63,N_14950,N_14996);
and UO_64 (O_64,N_14963,N_14983);
and UO_65 (O_65,N_14966,N_14877);
xor UO_66 (O_66,N_14878,N_14989);
xor UO_67 (O_67,N_14896,N_14928);
nor UO_68 (O_68,N_14914,N_14958);
nand UO_69 (O_69,N_14913,N_14924);
xnor UO_70 (O_70,N_14883,N_14989);
and UO_71 (O_71,N_14892,N_14900);
and UO_72 (O_72,N_14988,N_14929);
and UO_73 (O_73,N_14987,N_14919);
and UO_74 (O_74,N_14875,N_14954);
nor UO_75 (O_75,N_14955,N_14907);
nor UO_76 (O_76,N_14978,N_14903);
nor UO_77 (O_77,N_14979,N_14929);
nor UO_78 (O_78,N_14948,N_14969);
xnor UO_79 (O_79,N_14953,N_14924);
nand UO_80 (O_80,N_14879,N_14888);
and UO_81 (O_81,N_14963,N_14878);
and UO_82 (O_82,N_14922,N_14967);
and UO_83 (O_83,N_14968,N_14890);
or UO_84 (O_84,N_14964,N_14902);
xor UO_85 (O_85,N_14983,N_14977);
nor UO_86 (O_86,N_14936,N_14956);
nor UO_87 (O_87,N_14930,N_14886);
nand UO_88 (O_88,N_14908,N_14966);
or UO_89 (O_89,N_14982,N_14910);
nor UO_90 (O_90,N_14878,N_14919);
nand UO_91 (O_91,N_14936,N_14945);
xor UO_92 (O_92,N_14976,N_14968);
xnor UO_93 (O_93,N_14956,N_14891);
nor UO_94 (O_94,N_14931,N_14972);
nor UO_95 (O_95,N_14936,N_14901);
or UO_96 (O_96,N_14912,N_14882);
and UO_97 (O_97,N_14940,N_14968);
xnor UO_98 (O_98,N_14875,N_14994);
nand UO_99 (O_99,N_14982,N_14991);
xor UO_100 (O_100,N_14945,N_14934);
nand UO_101 (O_101,N_14920,N_14941);
nor UO_102 (O_102,N_14918,N_14907);
nand UO_103 (O_103,N_14945,N_14994);
nor UO_104 (O_104,N_14933,N_14989);
and UO_105 (O_105,N_14888,N_14984);
nand UO_106 (O_106,N_14928,N_14989);
and UO_107 (O_107,N_14876,N_14980);
nand UO_108 (O_108,N_14994,N_14955);
nor UO_109 (O_109,N_14976,N_14892);
and UO_110 (O_110,N_14907,N_14909);
and UO_111 (O_111,N_14988,N_14963);
or UO_112 (O_112,N_14885,N_14974);
and UO_113 (O_113,N_14962,N_14987);
nand UO_114 (O_114,N_14966,N_14926);
xnor UO_115 (O_115,N_14931,N_14978);
and UO_116 (O_116,N_14928,N_14958);
and UO_117 (O_117,N_14884,N_14965);
nor UO_118 (O_118,N_14946,N_14904);
nand UO_119 (O_119,N_14997,N_14941);
nand UO_120 (O_120,N_14937,N_14998);
nor UO_121 (O_121,N_14915,N_14911);
nand UO_122 (O_122,N_14948,N_14917);
nand UO_123 (O_123,N_14919,N_14979);
and UO_124 (O_124,N_14962,N_14882);
nand UO_125 (O_125,N_14906,N_14911);
xor UO_126 (O_126,N_14922,N_14964);
nor UO_127 (O_127,N_14922,N_14876);
or UO_128 (O_128,N_14895,N_14985);
nand UO_129 (O_129,N_14917,N_14953);
xnor UO_130 (O_130,N_14924,N_14934);
nand UO_131 (O_131,N_14944,N_14991);
and UO_132 (O_132,N_14994,N_14932);
nand UO_133 (O_133,N_14983,N_14978);
or UO_134 (O_134,N_14997,N_14984);
and UO_135 (O_135,N_14914,N_14966);
xnor UO_136 (O_136,N_14884,N_14953);
or UO_137 (O_137,N_14999,N_14913);
xor UO_138 (O_138,N_14981,N_14926);
xnor UO_139 (O_139,N_14904,N_14921);
nor UO_140 (O_140,N_14928,N_14996);
xnor UO_141 (O_141,N_14925,N_14955);
xnor UO_142 (O_142,N_14901,N_14968);
or UO_143 (O_143,N_14954,N_14967);
or UO_144 (O_144,N_14904,N_14995);
or UO_145 (O_145,N_14980,N_14957);
or UO_146 (O_146,N_14998,N_14881);
nand UO_147 (O_147,N_14952,N_14978);
nor UO_148 (O_148,N_14879,N_14886);
nand UO_149 (O_149,N_14876,N_14924);
nor UO_150 (O_150,N_14996,N_14906);
or UO_151 (O_151,N_14879,N_14977);
and UO_152 (O_152,N_14959,N_14981);
and UO_153 (O_153,N_14882,N_14897);
xor UO_154 (O_154,N_14959,N_14953);
nand UO_155 (O_155,N_14954,N_14941);
xor UO_156 (O_156,N_14893,N_14888);
nand UO_157 (O_157,N_14990,N_14885);
or UO_158 (O_158,N_14902,N_14943);
or UO_159 (O_159,N_14911,N_14962);
xor UO_160 (O_160,N_14962,N_14942);
nor UO_161 (O_161,N_14906,N_14887);
nand UO_162 (O_162,N_14916,N_14885);
nand UO_163 (O_163,N_14993,N_14888);
nand UO_164 (O_164,N_14923,N_14976);
nand UO_165 (O_165,N_14945,N_14876);
and UO_166 (O_166,N_14948,N_14964);
or UO_167 (O_167,N_14996,N_14989);
nand UO_168 (O_168,N_14884,N_14928);
or UO_169 (O_169,N_14882,N_14884);
and UO_170 (O_170,N_14932,N_14977);
and UO_171 (O_171,N_14913,N_14970);
nor UO_172 (O_172,N_14947,N_14972);
and UO_173 (O_173,N_14902,N_14962);
xor UO_174 (O_174,N_14886,N_14893);
and UO_175 (O_175,N_14986,N_14955);
xnor UO_176 (O_176,N_14958,N_14952);
nand UO_177 (O_177,N_14957,N_14981);
nand UO_178 (O_178,N_14991,N_14961);
nor UO_179 (O_179,N_14950,N_14974);
xor UO_180 (O_180,N_14993,N_14916);
xor UO_181 (O_181,N_14978,N_14883);
nand UO_182 (O_182,N_14930,N_14952);
nand UO_183 (O_183,N_14913,N_14875);
nand UO_184 (O_184,N_14905,N_14986);
nand UO_185 (O_185,N_14987,N_14932);
nand UO_186 (O_186,N_14908,N_14927);
nand UO_187 (O_187,N_14935,N_14937);
nand UO_188 (O_188,N_14906,N_14875);
xnor UO_189 (O_189,N_14996,N_14975);
nor UO_190 (O_190,N_14964,N_14952);
nor UO_191 (O_191,N_14910,N_14915);
nand UO_192 (O_192,N_14971,N_14950);
xnor UO_193 (O_193,N_14950,N_14949);
nor UO_194 (O_194,N_14952,N_14877);
or UO_195 (O_195,N_14895,N_14991);
and UO_196 (O_196,N_14976,N_14882);
nand UO_197 (O_197,N_14948,N_14996);
nor UO_198 (O_198,N_14942,N_14944);
or UO_199 (O_199,N_14912,N_14934);
or UO_200 (O_200,N_14916,N_14879);
or UO_201 (O_201,N_14879,N_14952);
nand UO_202 (O_202,N_14882,N_14935);
nor UO_203 (O_203,N_14978,N_14979);
and UO_204 (O_204,N_14920,N_14971);
or UO_205 (O_205,N_14955,N_14895);
or UO_206 (O_206,N_14941,N_14913);
nand UO_207 (O_207,N_14888,N_14896);
nor UO_208 (O_208,N_14910,N_14957);
and UO_209 (O_209,N_14934,N_14908);
or UO_210 (O_210,N_14950,N_14970);
nor UO_211 (O_211,N_14888,N_14995);
and UO_212 (O_212,N_14986,N_14961);
or UO_213 (O_213,N_14900,N_14982);
or UO_214 (O_214,N_14904,N_14932);
and UO_215 (O_215,N_14998,N_14976);
nand UO_216 (O_216,N_14986,N_14953);
nand UO_217 (O_217,N_14946,N_14894);
xnor UO_218 (O_218,N_14933,N_14937);
or UO_219 (O_219,N_14882,N_14989);
or UO_220 (O_220,N_14954,N_14983);
nand UO_221 (O_221,N_14967,N_14943);
or UO_222 (O_222,N_14917,N_14928);
nor UO_223 (O_223,N_14918,N_14978);
or UO_224 (O_224,N_14992,N_14911);
or UO_225 (O_225,N_14877,N_14991);
xnor UO_226 (O_226,N_14897,N_14986);
nand UO_227 (O_227,N_14981,N_14966);
or UO_228 (O_228,N_14948,N_14985);
and UO_229 (O_229,N_14917,N_14964);
or UO_230 (O_230,N_14916,N_14910);
nand UO_231 (O_231,N_14880,N_14976);
nand UO_232 (O_232,N_14915,N_14993);
and UO_233 (O_233,N_14951,N_14954);
nor UO_234 (O_234,N_14967,N_14879);
and UO_235 (O_235,N_14875,N_14894);
xnor UO_236 (O_236,N_14939,N_14967);
xnor UO_237 (O_237,N_14934,N_14899);
nand UO_238 (O_238,N_14920,N_14909);
or UO_239 (O_239,N_14899,N_14925);
and UO_240 (O_240,N_14991,N_14981);
or UO_241 (O_241,N_14994,N_14978);
nor UO_242 (O_242,N_14922,N_14939);
nand UO_243 (O_243,N_14875,N_14949);
nor UO_244 (O_244,N_14912,N_14947);
xnor UO_245 (O_245,N_14951,N_14960);
and UO_246 (O_246,N_14915,N_14955);
or UO_247 (O_247,N_14901,N_14894);
nand UO_248 (O_248,N_14993,N_14987);
and UO_249 (O_249,N_14928,N_14993);
or UO_250 (O_250,N_14878,N_14911);
xnor UO_251 (O_251,N_14936,N_14964);
nand UO_252 (O_252,N_14918,N_14931);
nand UO_253 (O_253,N_14897,N_14966);
nor UO_254 (O_254,N_14969,N_14903);
or UO_255 (O_255,N_14960,N_14922);
nand UO_256 (O_256,N_14973,N_14934);
nor UO_257 (O_257,N_14887,N_14923);
nand UO_258 (O_258,N_14884,N_14911);
and UO_259 (O_259,N_14905,N_14895);
nand UO_260 (O_260,N_14984,N_14958);
nand UO_261 (O_261,N_14919,N_14876);
or UO_262 (O_262,N_14945,N_14886);
and UO_263 (O_263,N_14929,N_14952);
nor UO_264 (O_264,N_14984,N_14884);
nor UO_265 (O_265,N_14879,N_14889);
nor UO_266 (O_266,N_14907,N_14899);
nand UO_267 (O_267,N_14884,N_14894);
or UO_268 (O_268,N_14995,N_14881);
nand UO_269 (O_269,N_14983,N_14903);
nand UO_270 (O_270,N_14877,N_14901);
or UO_271 (O_271,N_14982,N_14909);
nand UO_272 (O_272,N_14939,N_14999);
nor UO_273 (O_273,N_14876,N_14957);
nor UO_274 (O_274,N_14912,N_14935);
or UO_275 (O_275,N_14925,N_14904);
and UO_276 (O_276,N_14894,N_14959);
and UO_277 (O_277,N_14934,N_14896);
nor UO_278 (O_278,N_14960,N_14943);
xnor UO_279 (O_279,N_14948,N_14951);
nor UO_280 (O_280,N_14935,N_14969);
or UO_281 (O_281,N_14880,N_14883);
nor UO_282 (O_282,N_14910,N_14966);
nor UO_283 (O_283,N_14963,N_14894);
nor UO_284 (O_284,N_14960,N_14975);
nor UO_285 (O_285,N_14937,N_14951);
or UO_286 (O_286,N_14878,N_14875);
and UO_287 (O_287,N_14881,N_14953);
xor UO_288 (O_288,N_14936,N_14882);
and UO_289 (O_289,N_14931,N_14957);
and UO_290 (O_290,N_14940,N_14974);
or UO_291 (O_291,N_14983,N_14966);
xor UO_292 (O_292,N_14970,N_14984);
nor UO_293 (O_293,N_14934,N_14959);
nand UO_294 (O_294,N_14955,N_14918);
nand UO_295 (O_295,N_14904,N_14891);
xnor UO_296 (O_296,N_14970,N_14910);
nor UO_297 (O_297,N_14998,N_14944);
nor UO_298 (O_298,N_14963,N_14979);
or UO_299 (O_299,N_14880,N_14950);
nor UO_300 (O_300,N_14977,N_14995);
and UO_301 (O_301,N_14880,N_14894);
and UO_302 (O_302,N_14922,N_14892);
xor UO_303 (O_303,N_14915,N_14995);
or UO_304 (O_304,N_14945,N_14924);
xor UO_305 (O_305,N_14975,N_14966);
or UO_306 (O_306,N_14904,N_14958);
and UO_307 (O_307,N_14897,N_14968);
and UO_308 (O_308,N_14950,N_14998);
and UO_309 (O_309,N_14884,N_14940);
nor UO_310 (O_310,N_14924,N_14941);
and UO_311 (O_311,N_14973,N_14949);
nor UO_312 (O_312,N_14922,N_14887);
nor UO_313 (O_313,N_14991,N_14972);
nand UO_314 (O_314,N_14930,N_14908);
nand UO_315 (O_315,N_14920,N_14887);
and UO_316 (O_316,N_14929,N_14942);
xnor UO_317 (O_317,N_14957,N_14964);
nand UO_318 (O_318,N_14988,N_14907);
nand UO_319 (O_319,N_14993,N_14879);
and UO_320 (O_320,N_14918,N_14912);
xor UO_321 (O_321,N_14884,N_14966);
nor UO_322 (O_322,N_14889,N_14977);
nor UO_323 (O_323,N_14983,N_14972);
xnor UO_324 (O_324,N_14941,N_14978);
nand UO_325 (O_325,N_14930,N_14936);
and UO_326 (O_326,N_14998,N_14947);
or UO_327 (O_327,N_14982,N_14878);
xnor UO_328 (O_328,N_14918,N_14975);
xor UO_329 (O_329,N_14966,N_14976);
nor UO_330 (O_330,N_14940,N_14890);
xnor UO_331 (O_331,N_14990,N_14936);
or UO_332 (O_332,N_14883,N_14887);
nand UO_333 (O_333,N_14931,N_14952);
xor UO_334 (O_334,N_14932,N_14988);
or UO_335 (O_335,N_14998,N_14964);
nor UO_336 (O_336,N_14920,N_14921);
and UO_337 (O_337,N_14936,N_14983);
xnor UO_338 (O_338,N_14980,N_14914);
nor UO_339 (O_339,N_14991,N_14899);
and UO_340 (O_340,N_14884,N_14880);
or UO_341 (O_341,N_14941,N_14974);
or UO_342 (O_342,N_14893,N_14991);
nor UO_343 (O_343,N_14967,N_14908);
nor UO_344 (O_344,N_14985,N_14983);
or UO_345 (O_345,N_14968,N_14921);
or UO_346 (O_346,N_14957,N_14984);
or UO_347 (O_347,N_14964,N_14999);
nor UO_348 (O_348,N_14983,N_14941);
or UO_349 (O_349,N_14974,N_14880);
xor UO_350 (O_350,N_14972,N_14927);
nor UO_351 (O_351,N_14898,N_14968);
nor UO_352 (O_352,N_14879,N_14883);
or UO_353 (O_353,N_14948,N_14999);
nand UO_354 (O_354,N_14969,N_14952);
nor UO_355 (O_355,N_14885,N_14948);
xnor UO_356 (O_356,N_14962,N_14885);
nand UO_357 (O_357,N_14946,N_14932);
or UO_358 (O_358,N_14981,N_14922);
and UO_359 (O_359,N_14891,N_14999);
and UO_360 (O_360,N_14985,N_14893);
or UO_361 (O_361,N_14889,N_14979);
or UO_362 (O_362,N_14998,N_14877);
nand UO_363 (O_363,N_14969,N_14896);
nor UO_364 (O_364,N_14904,N_14991);
xnor UO_365 (O_365,N_14955,N_14929);
and UO_366 (O_366,N_14970,N_14995);
nor UO_367 (O_367,N_14975,N_14900);
xnor UO_368 (O_368,N_14884,N_14908);
xnor UO_369 (O_369,N_14887,N_14987);
and UO_370 (O_370,N_14898,N_14877);
and UO_371 (O_371,N_14980,N_14898);
nor UO_372 (O_372,N_14931,N_14913);
or UO_373 (O_373,N_14943,N_14977);
and UO_374 (O_374,N_14990,N_14942);
nand UO_375 (O_375,N_14983,N_14914);
xor UO_376 (O_376,N_14966,N_14934);
or UO_377 (O_377,N_14976,N_14969);
nor UO_378 (O_378,N_14998,N_14915);
nor UO_379 (O_379,N_14878,N_14962);
nor UO_380 (O_380,N_14915,N_14938);
and UO_381 (O_381,N_14987,N_14959);
xor UO_382 (O_382,N_14955,N_14891);
or UO_383 (O_383,N_14884,N_14981);
nor UO_384 (O_384,N_14985,N_14877);
xnor UO_385 (O_385,N_14915,N_14987);
and UO_386 (O_386,N_14953,N_14907);
nand UO_387 (O_387,N_14935,N_14925);
nor UO_388 (O_388,N_14989,N_14966);
and UO_389 (O_389,N_14933,N_14918);
or UO_390 (O_390,N_14937,N_14939);
and UO_391 (O_391,N_14971,N_14960);
nor UO_392 (O_392,N_14988,N_14945);
nand UO_393 (O_393,N_14982,N_14978);
nand UO_394 (O_394,N_14933,N_14958);
xnor UO_395 (O_395,N_14980,N_14952);
or UO_396 (O_396,N_14894,N_14900);
or UO_397 (O_397,N_14988,N_14880);
nand UO_398 (O_398,N_14938,N_14943);
or UO_399 (O_399,N_14993,N_14974);
xnor UO_400 (O_400,N_14875,N_14987);
nand UO_401 (O_401,N_14965,N_14937);
or UO_402 (O_402,N_14889,N_14893);
or UO_403 (O_403,N_14933,N_14882);
nand UO_404 (O_404,N_14940,N_14984);
nand UO_405 (O_405,N_14968,N_14924);
and UO_406 (O_406,N_14945,N_14948);
and UO_407 (O_407,N_14931,N_14966);
nand UO_408 (O_408,N_14959,N_14944);
or UO_409 (O_409,N_14982,N_14901);
nor UO_410 (O_410,N_14901,N_14930);
or UO_411 (O_411,N_14878,N_14994);
xor UO_412 (O_412,N_14973,N_14901);
nor UO_413 (O_413,N_14968,N_14965);
and UO_414 (O_414,N_14884,N_14944);
or UO_415 (O_415,N_14979,N_14909);
or UO_416 (O_416,N_14952,N_14893);
and UO_417 (O_417,N_14948,N_14938);
xor UO_418 (O_418,N_14896,N_14900);
nand UO_419 (O_419,N_14946,N_14926);
or UO_420 (O_420,N_14932,N_14934);
nor UO_421 (O_421,N_14980,N_14953);
xor UO_422 (O_422,N_14990,N_14991);
nor UO_423 (O_423,N_14922,N_14928);
xnor UO_424 (O_424,N_14951,N_14941);
xnor UO_425 (O_425,N_14947,N_14917);
or UO_426 (O_426,N_14889,N_14927);
nor UO_427 (O_427,N_14953,N_14960);
nand UO_428 (O_428,N_14998,N_14891);
and UO_429 (O_429,N_14975,N_14958);
and UO_430 (O_430,N_14907,N_14977);
nand UO_431 (O_431,N_14955,N_14983);
nand UO_432 (O_432,N_14977,N_14880);
nand UO_433 (O_433,N_14972,N_14966);
nor UO_434 (O_434,N_14902,N_14993);
and UO_435 (O_435,N_14911,N_14986);
or UO_436 (O_436,N_14934,N_14905);
and UO_437 (O_437,N_14975,N_14970);
and UO_438 (O_438,N_14892,N_14953);
or UO_439 (O_439,N_14909,N_14883);
xnor UO_440 (O_440,N_14898,N_14881);
xor UO_441 (O_441,N_14908,N_14952);
and UO_442 (O_442,N_14936,N_14925);
or UO_443 (O_443,N_14899,N_14982);
nand UO_444 (O_444,N_14989,N_14995);
or UO_445 (O_445,N_14888,N_14954);
or UO_446 (O_446,N_14878,N_14971);
or UO_447 (O_447,N_14952,N_14943);
nand UO_448 (O_448,N_14921,N_14885);
xor UO_449 (O_449,N_14885,N_14971);
and UO_450 (O_450,N_14992,N_14985);
xor UO_451 (O_451,N_14961,N_14895);
nor UO_452 (O_452,N_14926,N_14942);
nor UO_453 (O_453,N_14905,N_14968);
and UO_454 (O_454,N_14932,N_14966);
nor UO_455 (O_455,N_14954,N_14982);
and UO_456 (O_456,N_14935,N_14940);
nand UO_457 (O_457,N_14883,N_14977);
nand UO_458 (O_458,N_14997,N_14881);
and UO_459 (O_459,N_14938,N_14910);
and UO_460 (O_460,N_14938,N_14967);
nor UO_461 (O_461,N_14934,N_14944);
xnor UO_462 (O_462,N_14994,N_14898);
and UO_463 (O_463,N_14985,N_14962);
nand UO_464 (O_464,N_14909,N_14956);
or UO_465 (O_465,N_14882,N_14885);
or UO_466 (O_466,N_14875,N_14961);
and UO_467 (O_467,N_14876,N_14878);
xnor UO_468 (O_468,N_14946,N_14959);
and UO_469 (O_469,N_14906,N_14984);
nor UO_470 (O_470,N_14956,N_14901);
or UO_471 (O_471,N_14910,N_14964);
and UO_472 (O_472,N_14912,N_14973);
and UO_473 (O_473,N_14956,N_14995);
and UO_474 (O_474,N_14888,N_14991);
xnor UO_475 (O_475,N_14941,N_14952);
or UO_476 (O_476,N_14897,N_14952);
or UO_477 (O_477,N_14964,N_14930);
nand UO_478 (O_478,N_14961,N_14997);
nand UO_479 (O_479,N_14939,N_14876);
nor UO_480 (O_480,N_14954,N_14944);
or UO_481 (O_481,N_14904,N_14964);
nor UO_482 (O_482,N_14959,N_14954);
and UO_483 (O_483,N_14986,N_14928);
and UO_484 (O_484,N_14973,N_14889);
or UO_485 (O_485,N_14911,N_14889);
nor UO_486 (O_486,N_14903,N_14875);
or UO_487 (O_487,N_14917,N_14999);
or UO_488 (O_488,N_14952,N_14900);
nand UO_489 (O_489,N_14971,N_14987);
or UO_490 (O_490,N_14998,N_14967);
nand UO_491 (O_491,N_14975,N_14941);
and UO_492 (O_492,N_14915,N_14949);
nor UO_493 (O_493,N_14892,N_14934);
and UO_494 (O_494,N_14937,N_14888);
nand UO_495 (O_495,N_14915,N_14895);
xor UO_496 (O_496,N_14970,N_14949);
xnor UO_497 (O_497,N_14928,N_14974);
and UO_498 (O_498,N_14961,N_14940);
nand UO_499 (O_499,N_14904,N_14915);
nand UO_500 (O_500,N_14975,N_14937);
or UO_501 (O_501,N_14964,N_14925);
and UO_502 (O_502,N_14896,N_14948);
xor UO_503 (O_503,N_14978,N_14996);
and UO_504 (O_504,N_14994,N_14912);
nand UO_505 (O_505,N_14975,N_14984);
and UO_506 (O_506,N_14946,N_14916);
and UO_507 (O_507,N_14965,N_14977);
xor UO_508 (O_508,N_14891,N_14896);
xor UO_509 (O_509,N_14969,N_14898);
and UO_510 (O_510,N_14946,N_14988);
xnor UO_511 (O_511,N_14909,N_14911);
nand UO_512 (O_512,N_14893,N_14945);
or UO_513 (O_513,N_14897,N_14995);
xnor UO_514 (O_514,N_14971,N_14948);
xnor UO_515 (O_515,N_14991,N_14916);
xnor UO_516 (O_516,N_14981,N_14956);
nor UO_517 (O_517,N_14878,N_14987);
and UO_518 (O_518,N_14999,N_14993);
nand UO_519 (O_519,N_14893,N_14881);
nand UO_520 (O_520,N_14976,N_14965);
nor UO_521 (O_521,N_14882,N_14991);
nor UO_522 (O_522,N_14909,N_14950);
and UO_523 (O_523,N_14927,N_14893);
and UO_524 (O_524,N_14975,N_14992);
or UO_525 (O_525,N_14969,N_14906);
and UO_526 (O_526,N_14988,N_14927);
or UO_527 (O_527,N_14913,N_14929);
nand UO_528 (O_528,N_14984,N_14894);
and UO_529 (O_529,N_14875,N_14955);
nand UO_530 (O_530,N_14986,N_14919);
xnor UO_531 (O_531,N_14999,N_14894);
xnor UO_532 (O_532,N_14976,N_14930);
or UO_533 (O_533,N_14876,N_14956);
xnor UO_534 (O_534,N_14882,N_14914);
and UO_535 (O_535,N_14967,N_14976);
nand UO_536 (O_536,N_14949,N_14927);
nand UO_537 (O_537,N_14999,N_14881);
nand UO_538 (O_538,N_14986,N_14888);
nand UO_539 (O_539,N_14876,N_14997);
or UO_540 (O_540,N_14884,N_14901);
nand UO_541 (O_541,N_14940,N_14917);
nor UO_542 (O_542,N_14934,N_14911);
xnor UO_543 (O_543,N_14917,N_14899);
nor UO_544 (O_544,N_14973,N_14928);
or UO_545 (O_545,N_14905,N_14882);
nand UO_546 (O_546,N_14920,N_14932);
nand UO_547 (O_547,N_14878,N_14927);
or UO_548 (O_548,N_14935,N_14971);
nand UO_549 (O_549,N_14935,N_14876);
nand UO_550 (O_550,N_14992,N_14954);
nand UO_551 (O_551,N_14969,N_14929);
nand UO_552 (O_552,N_14947,N_14962);
xnor UO_553 (O_553,N_14909,N_14914);
xnor UO_554 (O_554,N_14978,N_14887);
nor UO_555 (O_555,N_14923,N_14946);
and UO_556 (O_556,N_14958,N_14949);
nor UO_557 (O_557,N_14989,N_14960);
and UO_558 (O_558,N_14939,N_14972);
nand UO_559 (O_559,N_14990,N_14986);
and UO_560 (O_560,N_14904,N_14997);
nand UO_561 (O_561,N_14935,N_14909);
xor UO_562 (O_562,N_14975,N_14936);
nor UO_563 (O_563,N_14934,N_14884);
xnor UO_564 (O_564,N_14891,N_14878);
nand UO_565 (O_565,N_14925,N_14937);
nor UO_566 (O_566,N_14906,N_14881);
or UO_567 (O_567,N_14962,N_14936);
xor UO_568 (O_568,N_14920,N_14991);
nor UO_569 (O_569,N_14901,N_14893);
or UO_570 (O_570,N_14944,N_14890);
and UO_571 (O_571,N_14952,N_14971);
nand UO_572 (O_572,N_14913,N_14998);
nor UO_573 (O_573,N_14880,N_14968);
xnor UO_574 (O_574,N_14977,N_14952);
or UO_575 (O_575,N_14978,N_14998);
nor UO_576 (O_576,N_14923,N_14886);
nand UO_577 (O_577,N_14938,N_14977);
nor UO_578 (O_578,N_14897,N_14931);
and UO_579 (O_579,N_14905,N_14994);
xnor UO_580 (O_580,N_14942,N_14920);
or UO_581 (O_581,N_14894,N_14925);
nor UO_582 (O_582,N_14950,N_14904);
and UO_583 (O_583,N_14995,N_14918);
or UO_584 (O_584,N_14913,N_14976);
and UO_585 (O_585,N_14952,N_14998);
or UO_586 (O_586,N_14947,N_14958);
and UO_587 (O_587,N_14885,N_14909);
or UO_588 (O_588,N_14934,N_14971);
and UO_589 (O_589,N_14901,N_14911);
or UO_590 (O_590,N_14899,N_14884);
or UO_591 (O_591,N_14905,N_14894);
nand UO_592 (O_592,N_14941,N_14968);
nor UO_593 (O_593,N_14940,N_14948);
or UO_594 (O_594,N_14992,N_14881);
or UO_595 (O_595,N_14946,N_14939);
xor UO_596 (O_596,N_14981,N_14933);
nand UO_597 (O_597,N_14901,N_14994);
or UO_598 (O_598,N_14921,N_14887);
nor UO_599 (O_599,N_14986,N_14958);
xor UO_600 (O_600,N_14925,N_14942);
nor UO_601 (O_601,N_14925,N_14944);
and UO_602 (O_602,N_14985,N_14968);
nand UO_603 (O_603,N_14954,N_14937);
xor UO_604 (O_604,N_14932,N_14984);
nand UO_605 (O_605,N_14994,N_14910);
or UO_606 (O_606,N_14953,N_14891);
nor UO_607 (O_607,N_14950,N_14916);
and UO_608 (O_608,N_14900,N_14984);
nor UO_609 (O_609,N_14883,N_14900);
xor UO_610 (O_610,N_14923,N_14897);
or UO_611 (O_611,N_14875,N_14892);
and UO_612 (O_612,N_14979,N_14936);
xor UO_613 (O_613,N_14952,N_14935);
nor UO_614 (O_614,N_14885,N_14891);
or UO_615 (O_615,N_14879,N_14998);
or UO_616 (O_616,N_14910,N_14948);
or UO_617 (O_617,N_14995,N_14901);
nand UO_618 (O_618,N_14977,N_14980);
nand UO_619 (O_619,N_14968,N_14923);
nand UO_620 (O_620,N_14957,N_14937);
or UO_621 (O_621,N_14946,N_14956);
nor UO_622 (O_622,N_14980,N_14970);
xnor UO_623 (O_623,N_14941,N_14936);
and UO_624 (O_624,N_14875,N_14888);
nor UO_625 (O_625,N_14954,N_14915);
and UO_626 (O_626,N_14920,N_14876);
and UO_627 (O_627,N_14884,N_14887);
and UO_628 (O_628,N_14887,N_14892);
nand UO_629 (O_629,N_14911,N_14954);
and UO_630 (O_630,N_14970,N_14974);
and UO_631 (O_631,N_14913,N_14940);
nor UO_632 (O_632,N_14972,N_14906);
and UO_633 (O_633,N_14990,N_14880);
or UO_634 (O_634,N_14892,N_14995);
nand UO_635 (O_635,N_14932,N_14978);
xnor UO_636 (O_636,N_14971,N_14993);
xnor UO_637 (O_637,N_14970,N_14978);
nand UO_638 (O_638,N_14903,N_14921);
nor UO_639 (O_639,N_14994,N_14986);
and UO_640 (O_640,N_14968,N_14918);
or UO_641 (O_641,N_14973,N_14941);
nand UO_642 (O_642,N_14895,N_14937);
xor UO_643 (O_643,N_14983,N_14952);
nor UO_644 (O_644,N_14902,N_14970);
and UO_645 (O_645,N_14946,N_14907);
nor UO_646 (O_646,N_14917,N_14982);
nor UO_647 (O_647,N_14988,N_14900);
or UO_648 (O_648,N_14974,N_14989);
xnor UO_649 (O_649,N_14903,N_14922);
nor UO_650 (O_650,N_14878,N_14992);
nand UO_651 (O_651,N_14945,N_14882);
or UO_652 (O_652,N_14997,N_14918);
or UO_653 (O_653,N_14970,N_14899);
nand UO_654 (O_654,N_14958,N_14890);
and UO_655 (O_655,N_14973,N_14974);
nand UO_656 (O_656,N_14990,N_14931);
or UO_657 (O_657,N_14932,N_14921);
nor UO_658 (O_658,N_14984,N_14953);
or UO_659 (O_659,N_14901,N_14919);
nor UO_660 (O_660,N_14895,N_14909);
and UO_661 (O_661,N_14901,N_14888);
xnor UO_662 (O_662,N_14971,N_14905);
nor UO_663 (O_663,N_14950,N_14922);
nand UO_664 (O_664,N_14976,N_14934);
and UO_665 (O_665,N_14961,N_14901);
or UO_666 (O_666,N_14933,N_14925);
and UO_667 (O_667,N_14920,N_14951);
and UO_668 (O_668,N_14963,N_14928);
or UO_669 (O_669,N_14957,N_14881);
and UO_670 (O_670,N_14943,N_14976);
nand UO_671 (O_671,N_14917,N_14894);
xnor UO_672 (O_672,N_14947,N_14935);
nand UO_673 (O_673,N_14989,N_14939);
and UO_674 (O_674,N_14966,N_14990);
nor UO_675 (O_675,N_14881,N_14894);
nor UO_676 (O_676,N_14905,N_14898);
nand UO_677 (O_677,N_14890,N_14923);
or UO_678 (O_678,N_14887,N_14901);
nand UO_679 (O_679,N_14885,N_14881);
or UO_680 (O_680,N_14900,N_14915);
nand UO_681 (O_681,N_14993,N_14930);
nor UO_682 (O_682,N_14901,N_14926);
nor UO_683 (O_683,N_14939,N_14893);
or UO_684 (O_684,N_14997,N_14990);
nand UO_685 (O_685,N_14966,N_14984);
xor UO_686 (O_686,N_14975,N_14907);
and UO_687 (O_687,N_14883,N_14971);
or UO_688 (O_688,N_14889,N_14942);
or UO_689 (O_689,N_14965,N_14898);
nor UO_690 (O_690,N_14929,N_14920);
xor UO_691 (O_691,N_14881,N_14972);
and UO_692 (O_692,N_14951,N_14955);
nor UO_693 (O_693,N_14971,N_14989);
and UO_694 (O_694,N_14885,N_14877);
and UO_695 (O_695,N_14997,N_14934);
nor UO_696 (O_696,N_14937,N_14940);
xor UO_697 (O_697,N_14984,N_14939);
nand UO_698 (O_698,N_14880,N_14992);
or UO_699 (O_699,N_14957,N_14918);
xor UO_700 (O_700,N_14879,N_14981);
nand UO_701 (O_701,N_14897,N_14891);
and UO_702 (O_702,N_14941,N_14958);
or UO_703 (O_703,N_14960,N_14958);
xor UO_704 (O_704,N_14883,N_14966);
nand UO_705 (O_705,N_14915,N_14982);
or UO_706 (O_706,N_14986,N_14964);
or UO_707 (O_707,N_14967,N_14884);
nor UO_708 (O_708,N_14904,N_14957);
and UO_709 (O_709,N_14915,N_14892);
nand UO_710 (O_710,N_14900,N_14973);
and UO_711 (O_711,N_14945,N_14922);
xor UO_712 (O_712,N_14920,N_14956);
nor UO_713 (O_713,N_14979,N_14949);
and UO_714 (O_714,N_14923,N_14917);
nor UO_715 (O_715,N_14907,N_14931);
nand UO_716 (O_716,N_14951,N_14935);
and UO_717 (O_717,N_14916,N_14973);
and UO_718 (O_718,N_14989,N_14951);
nand UO_719 (O_719,N_14929,N_14957);
nand UO_720 (O_720,N_14971,N_14946);
nor UO_721 (O_721,N_14987,N_14990);
nand UO_722 (O_722,N_14906,N_14940);
and UO_723 (O_723,N_14948,N_14977);
xnor UO_724 (O_724,N_14960,N_14959);
nand UO_725 (O_725,N_14945,N_14979);
nor UO_726 (O_726,N_14926,N_14899);
xor UO_727 (O_727,N_14905,N_14944);
nor UO_728 (O_728,N_14908,N_14916);
or UO_729 (O_729,N_14943,N_14992);
or UO_730 (O_730,N_14890,N_14951);
or UO_731 (O_731,N_14944,N_14985);
nor UO_732 (O_732,N_14986,N_14920);
nand UO_733 (O_733,N_14966,N_14986);
nand UO_734 (O_734,N_14916,N_14982);
nand UO_735 (O_735,N_14887,N_14936);
and UO_736 (O_736,N_14965,N_14926);
and UO_737 (O_737,N_14903,N_14987);
xnor UO_738 (O_738,N_14901,N_14947);
xor UO_739 (O_739,N_14915,N_14974);
nor UO_740 (O_740,N_14950,N_14910);
nand UO_741 (O_741,N_14958,N_14916);
or UO_742 (O_742,N_14900,N_14991);
nor UO_743 (O_743,N_14962,N_14932);
xor UO_744 (O_744,N_14996,N_14965);
and UO_745 (O_745,N_14986,N_14881);
or UO_746 (O_746,N_14900,N_14891);
or UO_747 (O_747,N_14936,N_14875);
nor UO_748 (O_748,N_14972,N_14961);
nand UO_749 (O_749,N_14976,N_14914);
and UO_750 (O_750,N_14992,N_14979);
or UO_751 (O_751,N_14888,N_14967);
nand UO_752 (O_752,N_14929,N_14900);
xor UO_753 (O_753,N_14907,N_14905);
xor UO_754 (O_754,N_14934,N_14900);
and UO_755 (O_755,N_14938,N_14893);
or UO_756 (O_756,N_14987,N_14944);
or UO_757 (O_757,N_14991,N_14875);
nand UO_758 (O_758,N_14982,N_14895);
xnor UO_759 (O_759,N_14984,N_14903);
xnor UO_760 (O_760,N_14908,N_14928);
nor UO_761 (O_761,N_14979,N_14985);
or UO_762 (O_762,N_14890,N_14994);
xnor UO_763 (O_763,N_14975,N_14964);
nand UO_764 (O_764,N_14949,N_14888);
nor UO_765 (O_765,N_14890,N_14876);
or UO_766 (O_766,N_14988,N_14993);
nor UO_767 (O_767,N_14905,N_14964);
nand UO_768 (O_768,N_14929,N_14917);
nor UO_769 (O_769,N_14917,N_14902);
nor UO_770 (O_770,N_14920,N_14926);
or UO_771 (O_771,N_14955,N_14878);
or UO_772 (O_772,N_14898,N_14986);
nand UO_773 (O_773,N_14949,N_14887);
nand UO_774 (O_774,N_14950,N_14993);
nor UO_775 (O_775,N_14898,N_14989);
nand UO_776 (O_776,N_14879,N_14910);
nand UO_777 (O_777,N_14999,N_14957);
and UO_778 (O_778,N_14916,N_14875);
or UO_779 (O_779,N_14901,N_14932);
nand UO_780 (O_780,N_14883,N_14892);
xnor UO_781 (O_781,N_14975,N_14912);
nor UO_782 (O_782,N_14928,N_14912);
or UO_783 (O_783,N_14879,N_14887);
or UO_784 (O_784,N_14918,N_14921);
nand UO_785 (O_785,N_14929,N_14949);
or UO_786 (O_786,N_14980,N_14991);
and UO_787 (O_787,N_14918,N_14917);
or UO_788 (O_788,N_14887,N_14990);
or UO_789 (O_789,N_14897,N_14908);
or UO_790 (O_790,N_14987,N_14986);
or UO_791 (O_791,N_14977,N_14926);
nor UO_792 (O_792,N_14923,N_14982);
or UO_793 (O_793,N_14977,N_14920);
and UO_794 (O_794,N_14881,N_14900);
xnor UO_795 (O_795,N_14891,N_14884);
nor UO_796 (O_796,N_14897,N_14886);
and UO_797 (O_797,N_14965,N_14961);
or UO_798 (O_798,N_14972,N_14903);
and UO_799 (O_799,N_14953,N_14893);
nor UO_800 (O_800,N_14890,N_14939);
or UO_801 (O_801,N_14955,N_14950);
or UO_802 (O_802,N_14920,N_14967);
nor UO_803 (O_803,N_14882,N_14880);
or UO_804 (O_804,N_14962,N_14923);
nor UO_805 (O_805,N_14954,N_14994);
nor UO_806 (O_806,N_14959,N_14927);
xor UO_807 (O_807,N_14985,N_14959);
and UO_808 (O_808,N_14881,N_14926);
xor UO_809 (O_809,N_14900,N_14913);
xnor UO_810 (O_810,N_14991,N_14977);
nor UO_811 (O_811,N_14877,N_14987);
xor UO_812 (O_812,N_14998,N_14999);
nor UO_813 (O_813,N_14952,N_14904);
nand UO_814 (O_814,N_14962,N_14954);
or UO_815 (O_815,N_14934,N_14964);
or UO_816 (O_816,N_14965,N_14957);
xnor UO_817 (O_817,N_14878,N_14896);
or UO_818 (O_818,N_14908,N_14925);
nor UO_819 (O_819,N_14880,N_14926);
and UO_820 (O_820,N_14943,N_14944);
nand UO_821 (O_821,N_14933,N_14947);
nand UO_822 (O_822,N_14976,N_14932);
nand UO_823 (O_823,N_14925,N_14987);
nor UO_824 (O_824,N_14926,N_14882);
and UO_825 (O_825,N_14924,N_14937);
xnor UO_826 (O_826,N_14913,N_14968);
xor UO_827 (O_827,N_14897,N_14965);
nor UO_828 (O_828,N_14976,N_14985);
nand UO_829 (O_829,N_14940,N_14923);
nand UO_830 (O_830,N_14930,N_14971);
xor UO_831 (O_831,N_14934,N_14889);
or UO_832 (O_832,N_14995,N_14896);
nor UO_833 (O_833,N_14908,N_14986);
nand UO_834 (O_834,N_14905,N_14927);
nor UO_835 (O_835,N_14962,N_14993);
nand UO_836 (O_836,N_14992,N_14974);
xor UO_837 (O_837,N_14896,N_14997);
and UO_838 (O_838,N_14959,N_14943);
xor UO_839 (O_839,N_14943,N_14966);
nand UO_840 (O_840,N_14897,N_14956);
and UO_841 (O_841,N_14882,N_14995);
or UO_842 (O_842,N_14886,N_14983);
nor UO_843 (O_843,N_14916,N_14972);
xnor UO_844 (O_844,N_14907,N_14996);
or UO_845 (O_845,N_14970,N_14903);
nor UO_846 (O_846,N_14999,N_14988);
nand UO_847 (O_847,N_14900,N_14906);
or UO_848 (O_848,N_14975,N_14908);
xor UO_849 (O_849,N_14880,N_14896);
xor UO_850 (O_850,N_14889,N_14888);
and UO_851 (O_851,N_14908,N_14977);
nand UO_852 (O_852,N_14990,N_14930);
nand UO_853 (O_853,N_14926,N_14936);
xnor UO_854 (O_854,N_14990,N_14884);
xnor UO_855 (O_855,N_14917,N_14980);
xnor UO_856 (O_856,N_14893,N_14954);
nand UO_857 (O_857,N_14886,N_14951);
nand UO_858 (O_858,N_14967,N_14877);
and UO_859 (O_859,N_14990,N_14954);
nor UO_860 (O_860,N_14960,N_14969);
or UO_861 (O_861,N_14930,N_14955);
xor UO_862 (O_862,N_14921,N_14884);
xnor UO_863 (O_863,N_14956,N_14964);
or UO_864 (O_864,N_14883,N_14917);
xnor UO_865 (O_865,N_14875,N_14993);
nand UO_866 (O_866,N_14998,N_14946);
and UO_867 (O_867,N_14960,N_14957);
and UO_868 (O_868,N_14975,N_14962);
nand UO_869 (O_869,N_14891,N_14905);
or UO_870 (O_870,N_14991,N_14996);
xnor UO_871 (O_871,N_14999,N_14953);
or UO_872 (O_872,N_14962,N_14982);
nand UO_873 (O_873,N_14918,N_14983);
nand UO_874 (O_874,N_14993,N_14941);
or UO_875 (O_875,N_14878,N_14941);
and UO_876 (O_876,N_14918,N_14969);
nor UO_877 (O_877,N_14928,N_14941);
nand UO_878 (O_878,N_14938,N_14996);
nor UO_879 (O_879,N_14946,N_14943);
and UO_880 (O_880,N_14887,N_14937);
xor UO_881 (O_881,N_14898,N_14998);
or UO_882 (O_882,N_14980,N_14959);
xnor UO_883 (O_883,N_14928,N_14997);
or UO_884 (O_884,N_14888,N_14912);
nand UO_885 (O_885,N_14932,N_14877);
or UO_886 (O_886,N_14963,N_14962);
xor UO_887 (O_887,N_14887,N_14964);
and UO_888 (O_888,N_14937,N_14938);
or UO_889 (O_889,N_14900,N_14950);
nor UO_890 (O_890,N_14955,N_14906);
nand UO_891 (O_891,N_14915,N_14906);
nand UO_892 (O_892,N_14944,N_14963);
and UO_893 (O_893,N_14984,N_14913);
nor UO_894 (O_894,N_14878,N_14937);
or UO_895 (O_895,N_14994,N_14998);
xor UO_896 (O_896,N_14949,N_14991);
xor UO_897 (O_897,N_14928,N_14878);
and UO_898 (O_898,N_14883,N_14924);
nor UO_899 (O_899,N_14935,N_14930);
xnor UO_900 (O_900,N_14896,N_14960);
or UO_901 (O_901,N_14917,N_14954);
and UO_902 (O_902,N_14958,N_14935);
nor UO_903 (O_903,N_14942,N_14902);
and UO_904 (O_904,N_14900,N_14922);
or UO_905 (O_905,N_14915,N_14989);
xnor UO_906 (O_906,N_14914,N_14895);
xor UO_907 (O_907,N_14880,N_14906);
xor UO_908 (O_908,N_14989,N_14908);
and UO_909 (O_909,N_14955,N_14998);
xor UO_910 (O_910,N_14953,N_14945);
xor UO_911 (O_911,N_14932,N_14922);
or UO_912 (O_912,N_14977,N_14940);
nor UO_913 (O_913,N_14919,N_14905);
nor UO_914 (O_914,N_14917,N_14886);
and UO_915 (O_915,N_14983,N_14953);
and UO_916 (O_916,N_14908,N_14972);
xor UO_917 (O_917,N_14909,N_14962);
xnor UO_918 (O_918,N_14925,N_14959);
or UO_919 (O_919,N_14917,N_14912);
xor UO_920 (O_920,N_14919,N_14892);
or UO_921 (O_921,N_14991,N_14956);
nor UO_922 (O_922,N_14927,N_14882);
nor UO_923 (O_923,N_14984,N_14936);
or UO_924 (O_924,N_14962,N_14901);
or UO_925 (O_925,N_14948,N_14939);
nand UO_926 (O_926,N_14981,N_14930);
nand UO_927 (O_927,N_14909,N_14966);
xor UO_928 (O_928,N_14943,N_14968);
and UO_929 (O_929,N_14918,N_14942);
xor UO_930 (O_930,N_14980,N_14993);
or UO_931 (O_931,N_14920,N_14985);
xnor UO_932 (O_932,N_14941,N_14985);
nor UO_933 (O_933,N_14897,N_14973);
and UO_934 (O_934,N_14878,N_14965);
or UO_935 (O_935,N_14885,N_14915);
or UO_936 (O_936,N_14972,N_14880);
or UO_937 (O_937,N_14883,N_14931);
nand UO_938 (O_938,N_14977,N_14928);
or UO_939 (O_939,N_14881,N_14887);
or UO_940 (O_940,N_14997,N_14900);
xnor UO_941 (O_941,N_14881,N_14932);
xor UO_942 (O_942,N_14941,N_14879);
xnor UO_943 (O_943,N_14887,N_14968);
or UO_944 (O_944,N_14924,N_14969);
nand UO_945 (O_945,N_14951,N_14979);
xnor UO_946 (O_946,N_14979,N_14984);
and UO_947 (O_947,N_14989,N_14893);
xor UO_948 (O_948,N_14936,N_14910);
or UO_949 (O_949,N_14982,N_14965);
or UO_950 (O_950,N_14984,N_14990);
nor UO_951 (O_951,N_14994,N_14968);
xor UO_952 (O_952,N_14890,N_14904);
nand UO_953 (O_953,N_14901,N_14987);
and UO_954 (O_954,N_14959,N_14890);
or UO_955 (O_955,N_14916,N_14920);
nand UO_956 (O_956,N_14906,N_14962);
nand UO_957 (O_957,N_14917,N_14897);
xor UO_958 (O_958,N_14954,N_14881);
nor UO_959 (O_959,N_14916,N_14933);
and UO_960 (O_960,N_14926,N_14932);
xnor UO_961 (O_961,N_14984,N_14995);
nor UO_962 (O_962,N_14908,N_14878);
or UO_963 (O_963,N_14965,N_14880);
or UO_964 (O_964,N_14878,N_14888);
and UO_965 (O_965,N_14893,N_14937);
nand UO_966 (O_966,N_14924,N_14919);
nor UO_967 (O_967,N_14942,N_14949);
nand UO_968 (O_968,N_14948,N_14967);
nand UO_969 (O_969,N_14995,N_14898);
nand UO_970 (O_970,N_14975,N_14952);
and UO_971 (O_971,N_14959,N_14884);
or UO_972 (O_972,N_14876,N_14911);
nor UO_973 (O_973,N_14969,N_14965);
and UO_974 (O_974,N_14888,N_14940);
nand UO_975 (O_975,N_14926,N_14904);
and UO_976 (O_976,N_14889,N_14928);
and UO_977 (O_977,N_14969,N_14958);
nand UO_978 (O_978,N_14955,N_14935);
nand UO_979 (O_979,N_14921,N_14925);
or UO_980 (O_980,N_14902,N_14958);
or UO_981 (O_981,N_14940,N_14912);
and UO_982 (O_982,N_14917,N_14890);
nand UO_983 (O_983,N_14936,N_14913);
nor UO_984 (O_984,N_14909,N_14904);
nor UO_985 (O_985,N_14980,N_14956);
xor UO_986 (O_986,N_14967,N_14975);
xor UO_987 (O_987,N_14996,N_14962);
nand UO_988 (O_988,N_14912,N_14920);
nor UO_989 (O_989,N_14982,N_14944);
xnor UO_990 (O_990,N_14971,N_14978);
or UO_991 (O_991,N_14993,N_14935);
xor UO_992 (O_992,N_14964,N_14908);
nand UO_993 (O_993,N_14912,N_14971);
xnor UO_994 (O_994,N_14899,N_14956);
or UO_995 (O_995,N_14975,N_14894);
or UO_996 (O_996,N_14949,N_14981);
and UO_997 (O_997,N_14974,N_14926);
nand UO_998 (O_998,N_14937,N_14891);
or UO_999 (O_999,N_14975,N_14878);
and UO_1000 (O_1000,N_14947,N_14940);
nand UO_1001 (O_1001,N_14911,N_14925);
or UO_1002 (O_1002,N_14916,N_14956);
nor UO_1003 (O_1003,N_14986,N_14975);
xor UO_1004 (O_1004,N_14989,N_14929);
or UO_1005 (O_1005,N_14943,N_14909);
nand UO_1006 (O_1006,N_14919,N_14967);
nor UO_1007 (O_1007,N_14903,N_14958);
xor UO_1008 (O_1008,N_14990,N_14922);
or UO_1009 (O_1009,N_14950,N_14959);
nand UO_1010 (O_1010,N_14927,N_14901);
xor UO_1011 (O_1011,N_14980,N_14998);
nand UO_1012 (O_1012,N_14959,N_14897);
or UO_1013 (O_1013,N_14921,N_14935);
or UO_1014 (O_1014,N_14998,N_14914);
nand UO_1015 (O_1015,N_14913,N_14897);
xor UO_1016 (O_1016,N_14881,N_14964);
and UO_1017 (O_1017,N_14927,N_14912);
or UO_1018 (O_1018,N_14992,N_14926);
nor UO_1019 (O_1019,N_14946,N_14921);
xnor UO_1020 (O_1020,N_14893,N_14924);
or UO_1021 (O_1021,N_14924,N_14925);
nor UO_1022 (O_1022,N_14967,N_14983);
nor UO_1023 (O_1023,N_14943,N_14999);
and UO_1024 (O_1024,N_14953,N_14985);
nand UO_1025 (O_1025,N_14953,N_14939);
or UO_1026 (O_1026,N_14955,N_14997);
xnor UO_1027 (O_1027,N_14888,N_14989);
and UO_1028 (O_1028,N_14946,N_14878);
nor UO_1029 (O_1029,N_14910,N_14930);
nor UO_1030 (O_1030,N_14916,N_14892);
and UO_1031 (O_1031,N_14942,N_14888);
xnor UO_1032 (O_1032,N_14887,N_14939);
and UO_1033 (O_1033,N_14978,N_14995);
nor UO_1034 (O_1034,N_14911,N_14922);
xor UO_1035 (O_1035,N_14963,N_14966);
or UO_1036 (O_1036,N_14977,N_14963);
nand UO_1037 (O_1037,N_14931,N_14950);
nor UO_1038 (O_1038,N_14996,N_14969);
nor UO_1039 (O_1039,N_14916,N_14961);
or UO_1040 (O_1040,N_14892,N_14912);
nor UO_1041 (O_1041,N_14994,N_14951);
nand UO_1042 (O_1042,N_14986,N_14900);
xnor UO_1043 (O_1043,N_14937,N_14900);
nor UO_1044 (O_1044,N_14875,N_14884);
nor UO_1045 (O_1045,N_14892,N_14990);
xor UO_1046 (O_1046,N_14924,N_14996);
nor UO_1047 (O_1047,N_14936,N_14890);
or UO_1048 (O_1048,N_14886,N_14969);
and UO_1049 (O_1049,N_14935,N_14973);
nor UO_1050 (O_1050,N_14931,N_14949);
xnor UO_1051 (O_1051,N_14898,N_14963);
and UO_1052 (O_1052,N_14989,N_14991);
nand UO_1053 (O_1053,N_14933,N_14976);
and UO_1054 (O_1054,N_14994,N_14993);
nand UO_1055 (O_1055,N_14893,N_14950);
xnor UO_1056 (O_1056,N_14942,N_14882);
xnor UO_1057 (O_1057,N_14962,N_14999);
or UO_1058 (O_1058,N_14994,N_14965);
nand UO_1059 (O_1059,N_14944,N_14914);
nor UO_1060 (O_1060,N_14923,N_14879);
or UO_1061 (O_1061,N_14918,N_14941);
nor UO_1062 (O_1062,N_14895,N_14925);
or UO_1063 (O_1063,N_14883,N_14985);
nor UO_1064 (O_1064,N_14968,N_14974);
or UO_1065 (O_1065,N_14885,N_14924);
and UO_1066 (O_1066,N_14919,N_14992);
nand UO_1067 (O_1067,N_14959,N_14993);
nor UO_1068 (O_1068,N_14914,N_14965);
or UO_1069 (O_1069,N_14983,N_14875);
nor UO_1070 (O_1070,N_14994,N_14907);
nand UO_1071 (O_1071,N_14879,N_14930);
nor UO_1072 (O_1072,N_14919,N_14926);
and UO_1073 (O_1073,N_14988,N_14914);
xnor UO_1074 (O_1074,N_14877,N_14935);
xor UO_1075 (O_1075,N_14973,N_14875);
nand UO_1076 (O_1076,N_14962,N_14907);
and UO_1077 (O_1077,N_14955,N_14988);
nor UO_1078 (O_1078,N_14989,N_14968);
nor UO_1079 (O_1079,N_14994,N_14942);
nand UO_1080 (O_1080,N_14947,N_14999);
nand UO_1081 (O_1081,N_14926,N_14945);
or UO_1082 (O_1082,N_14879,N_14912);
and UO_1083 (O_1083,N_14977,N_14881);
or UO_1084 (O_1084,N_14987,N_14955);
and UO_1085 (O_1085,N_14978,N_14972);
and UO_1086 (O_1086,N_14979,N_14888);
xor UO_1087 (O_1087,N_14891,N_14970);
xor UO_1088 (O_1088,N_14890,N_14975);
xnor UO_1089 (O_1089,N_14926,N_14985);
or UO_1090 (O_1090,N_14929,N_14884);
nand UO_1091 (O_1091,N_14957,N_14920);
xor UO_1092 (O_1092,N_14978,N_14902);
xnor UO_1093 (O_1093,N_14942,N_14934);
xor UO_1094 (O_1094,N_14956,N_14953);
and UO_1095 (O_1095,N_14973,N_14936);
nand UO_1096 (O_1096,N_14954,N_14939);
nand UO_1097 (O_1097,N_14955,N_14999);
xnor UO_1098 (O_1098,N_14922,N_14889);
and UO_1099 (O_1099,N_14922,N_14979);
and UO_1100 (O_1100,N_14944,N_14876);
nand UO_1101 (O_1101,N_14925,N_14891);
xnor UO_1102 (O_1102,N_14915,N_14902);
xor UO_1103 (O_1103,N_14996,N_14944);
and UO_1104 (O_1104,N_14977,N_14925);
xor UO_1105 (O_1105,N_14905,N_14876);
or UO_1106 (O_1106,N_14993,N_14899);
xor UO_1107 (O_1107,N_14930,N_14926);
and UO_1108 (O_1108,N_14934,N_14957);
nor UO_1109 (O_1109,N_14904,N_14917);
nand UO_1110 (O_1110,N_14997,N_14945);
or UO_1111 (O_1111,N_14956,N_14974);
nor UO_1112 (O_1112,N_14960,N_14963);
nor UO_1113 (O_1113,N_14886,N_14915);
or UO_1114 (O_1114,N_14979,N_14969);
nor UO_1115 (O_1115,N_14972,N_14932);
or UO_1116 (O_1116,N_14881,N_14903);
and UO_1117 (O_1117,N_14894,N_14921);
or UO_1118 (O_1118,N_14916,N_14925);
and UO_1119 (O_1119,N_14963,N_14933);
nor UO_1120 (O_1120,N_14970,N_14979);
and UO_1121 (O_1121,N_14977,N_14924);
nor UO_1122 (O_1122,N_14919,N_14953);
nand UO_1123 (O_1123,N_14884,N_14877);
xor UO_1124 (O_1124,N_14994,N_14880);
xnor UO_1125 (O_1125,N_14947,N_14945);
nor UO_1126 (O_1126,N_14884,N_14939);
nor UO_1127 (O_1127,N_14948,N_14905);
xor UO_1128 (O_1128,N_14919,N_14886);
or UO_1129 (O_1129,N_14969,N_14881);
and UO_1130 (O_1130,N_14961,N_14933);
nor UO_1131 (O_1131,N_14896,N_14890);
nand UO_1132 (O_1132,N_14956,N_14992);
or UO_1133 (O_1133,N_14895,N_14924);
or UO_1134 (O_1134,N_14998,N_14959);
xnor UO_1135 (O_1135,N_14950,N_14889);
nor UO_1136 (O_1136,N_14996,N_14937);
or UO_1137 (O_1137,N_14963,N_14895);
or UO_1138 (O_1138,N_14986,N_14932);
xor UO_1139 (O_1139,N_14904,N_14882);
nor UO_1140 (O_1140,N_14886,N_14972);
or UO_1141 (O_1141,N_14934,N_14974);
xnor UO_1142 (O_1142,N_14969,N_14988);
xnor UO_1143 (O_1143,N_14889,N_14877);
nand UO_1144 (O_1144,N_14931,N_14977);
xnor UO_1145 (O_1145,N_14900,N_14876);
nor UO_1146 (O_1146,N_14934,N_14933);
and UO_1147 (O_1147,N_14904,N_14919);
xnor UO_1148 (O_1148,N_14937,N_14918);
nand UO_1149 (O_1149,N_14892,N_14918);
nand UO_1150 (O_1150,N_14947,N_14949);
or UO_1151 (O_1151,N_14924,N_14891);
nand UO_1152 (O_1152,N_14974,N_14929);
nor UO_1153 (O_1153,N_14971,N_14951);
and UO_1154 (O_1154,N_14900,N_14901);
nand UO_1155 (O_1155,N_14897,N_14958);
or UO_1156 (O_1156,N_14959,N_14918);
nor UO_1157 (O_1157,N_14912,N_14979);
nor UO_1158 (O_1158,N_14987,N_14978);
nand UO_1159 (O_1159,N_14962,N_14881);
and UO_1160 (O_1160,N_14961,N_14959);
or UO_1161 (O_1161,N_14943,N_14963);
or UO_1162 (O_1162,N_14947,N_14913);
nand UO_1163 (O_1163,N_14975,N_14882);
xnor UO_1164 (O_1164,N_14897,N_14900);
nor UO_1165 (O_1165,N_14935,N_14903);
and UO_1166 (O_1166,N_14909,N_14997);
and UO_1167 (O_1167,N_14886,N_14901);
or UO_1168 (O_1168,N_14988,N_14956);
nor UO_1169 (O_1169,N_14992,N_14983);
and UO_1170 (O_1170,N_14887,N_14924);
and UO_1171 (O_1171,N_14990,N_14995);
nand UO_1172 (O_1172,N_14974,N_14882);
nand UO_1173 (O_1173,N_14955,N_14909);
nor UO_1174 (O_1174,N_14901,N_14891);
nor UO_1175 (O_1175,N_14930,N_14884);
nor UO_1176 (O_1176,N_14898,N_14888);
nor UO_1177 (O_1177,N_14931,N_14989);
or UO_1178 (O_1178,N_14923,N_14924);
and UO_1179 (O_1179,N_14893,N_14962);
or UO_1180 (O_1180,N_14884,N_14980);
nand UO_1181 (O_1181,N_14888,N_14971);
nand UO_1182 (O_1182,N_14911,N_14980);
xnor UO_1183 (O_1183,N_14929,N_14999);
and UO_1184 (O_1184,N_14974,N_14958);
xor UO_1185 (O_1185,N_14963,N_14956);
xor UO_1186 (O_1186,N_14951,N_14880);
and UO_1187 (O_1187,N_14981,N_14920);
or UO_1188 (O_1188,N_14945,N_14961);
xor UO_1189 (O_1189,N_14927,N_14877);
nand UO_1190 (O_1190,N_14904,N_14896);
or UO_1191 (O_1191,N_14933,N_14879);
nand UO_1192 (O_1192,N_14900,N_14886);
nand UO_1193 (O_1193,N_14957,N_14995);
and UO_1194 (O_1194,N_14882,N_14958);
or UO_1195 (O_1195,N_14903,N_14959);
nor UO_1196 (O_1196,N_14972,N_14992);
and UO_1197 (O_1197,N_14983,N_14927);
nor UO_1198 (O_1198,N_14961,N_14950);
and UO_1199 (O_1199,N_14929,N_14937);
xnor UO_1200 (O_1200,N_14986,N_14991);
xnor UO_1201 (O_1201,N_14879,N_14909);
and UO_1202 (O_1202,N_14936,N_14954);
xnor UO_1203 (O_1203,N_14990,N_14940);
or UO_1204 (O_1204,N_14935,N_14995);
nand UO_1205 (O_1205,N_14953,N_14936);
and UO_1206 (O_1206,N_14954,N_14882);
xor UO_1207 (O_1207,N_14996,N_14893);
nand UO_1208 (O_1208,N_14978,N_14950);
or UO_1209 (O_1209,N_14948,N_14990);
xor UO_1210 (O_1210,N_14898,N_14979);
and UO_1211 (O_1211,N_14961,N_14992);
or UO_1212 (O_1212,N_14918,N_14913);
nor UO_1213 (O_1213,N_14923,N_14955);
xnor UO_1214 (O_1214,N_14907,N_14928);
nor UO_1215 (O_1215,N_14877,N_14984);
nor UO_1216 (O_1216,N_14948,N_14920);
nor UO_1217 (O_1217,N_14925,N_14913);
xnor UO_1218 (O_1218,N_14985,N_14898);
and UO_1219 (O_1219,N_14965,N_14974);
or UO_1220 (O_1220,N_14931,N_14891);
xor UO_1221 (O_1221,N_14992,N_14933);
or UO_1222 (O_1222,N_14941,N_14931);
and UO_1223 (O_1223,N_14953,N_14949);
or UO_1224 (O_1224,N_14986,N_14886);
or UO_1225 (O_1225,N_14936,N_14916);
nor UO_1226 (O_1226,N_14897,N_14894);
xnor UO_1227 (O_1227,N_14913,N_14986);
or UO_1228 (O_1228,N_14969,N_14934);
or UO_1229 (O_1229,N_14950,N_14895);
nor UO_1230 (O_1230,N_14922,N_14925);
or UO_1231 (O_1231,N_14887,N_14916);
nor UO_1232 (O_1232,N_14890,N_14922);
nand UO_1233 (O_1233,N_14925,N_14991);
or UO_1234 (O_1234,N_14899,N_14937);
and UO_1235 (O_1235,N_14966,N_14944);
nor UO_1236 (O_1236,N_14952,N_14945);
nand UO_1237 (O_1237,N_14981,N_14992);
xnor UO_1238 (O_1238,N_14961,N_14880);
xnor UO_1239 (O_1239,N_14994,N_14977);
nor UO_1240 (O_1240,N_14955,N_14970);
nand UO_1241 (O_1241,N_14941,N_14946);
or UO_1242 (O_1242,N_14899,N_14915);
or UO_1243 (O_1243,N_14908,N_14905);
or UO_1244 (O_1244,N_14999,N_14884);
or UO_1245 (O_1245,N_14905,N_14953);
xnor UO_1246 (O_1246,N_14919,N_14983);
nor UO_1247 (O_1247,N_14893,N_14926);
or UO_1248 (O_1248,N_14954,N_14988);
nor UO_1249 (O_1249,N_14988,N_14944);
xor UO_1250 (O_1250,N_14914,N_14923);
or UO_1251 (O_1251,N_14966,N_14896);
and UO_1252 (O_1252,N_14942,N_14912);
or UO_1253 (O_1253,N_14978,N_14981);
xor UO_1254 (O_1254,N_14946,N_14901);
or UO_1255 (O_1255,N_14875,N_14970);
nor UO_1256 (O_1256,N_14938,N_14958);
xor UO_1257 (O_1257,N_14909,N_14902);
or UO_1258 (O_1258,N_14900,N_14931);
xnor UO_1259 (O_1259,N_14979,N_14892);
nor UO_1260 (O_1260,N_14921,N_14933);
or UO_1261 (O_1261,N_14966,N_14997);
nor UO_1262 (O_1262,N_14890,N_14998);
xnor UO_1263 (O_1263,N_14877,N_14875);
xnor UO_1264 (O_1264,N_14951,N_14943);
and UO_1265 (O_1265,N_14894,N_14893);
or UO_1266 (O_1266,N_14972,N_14929);
or UO_1267 (O_1267,N_14921,N_14900);
nor UO_1268 (O_1268,N_14988,N_14942);
xor UO_1269 (O_1269,N_14985,N_14888);
and UO_1270 (O_1270,N_14997,N_14969);
and UO_1271 (O_1271,N_14950,N_14883);
or UO_1272 (O_1272,N_14980,N_14960);
nand UO_1273 (O_1273,N_14997,N_14998);
nand UO_1274 (O_1274,N_14919,N_14920);
nor UO_1275 (O_1275,N_14929,N_14991);
nor UO_1276 (O_1276,N_14903,N_14937);
or UO_1277 (O_1277,N_14990,N_14935);
or UO_1278 (O_1278,N_14928,N_14995);
xor UO_1279 (O_1279,N_14926,N_14941);
nor UO_1280 (O_1280,N_14989,N_14930);
nand UO_1281 (O_1281,N_14876,N_14913);
nand UO_1282 (O_1282,N_14931,N_14924);
nor UO_1283 (O_1283,N_14965,N_14924);
and UO_1284 (O_1284,N_14948,N_14994);
nand UO_1285 (O_1285,N_14992,N_14886);
or UO_1286 (O_1286,N_14905,N_14957);
and UO_1287 (O_1287,N_14910,N_14947);
and UO_1288 (O_1288,N_14997,N_14948);
nor UO_1289 (O_1289,N_14905,N_14892);
or UO_1290 (O_1290,N_14985,N_14996);
nor UO_1291 (O_1291,N_14916,N_14945);
or UO_1292 (O_1292,N_14948,N_14925);
xor UO_1293 (O_1293,N_14896,N_14955);
or UO_1294 (O_1294,N_14920,N_14886);
nor UO_1295 (O_1295,N_14943,N_14911);
and UO_1296 (O_1296,N_14945,N_14923);
xnor UO_1297 (O_1297,N_14988,N_14901);
and UO_1298 (O_1298,N_14877,N_14973);
and UO_1299 (O_1299,N_14914,N_14950);
nand UO_1300 (O_1300,N_14963,N_14892);
nor UO_1301 (O_1301,N_14939,N_14906);
nand UO_1302 (O_1302,N_14976,N_14875);
and UO_1303 (O_1303,N_14917,N_14916);
and UO_1304 (O_1304,N_14993,N_14966);
xnor UO_1305 (O_1305,N_14971,N_14936);
nand UO_1306 (O_1306,N_14953,N_14914);
or UO_1307 (O_1307,N_14908,N_14957);
or UO_1308 (O_1308,N_14902,N_14893);
xor UO_1309 (O_1309,N_14956,N_14929);
and UO_1310 (O_1310,N_14973,N_14970);
or UO_1311 (O_1311,N_14984,N_14978);
xnor UO_1312 (O_1312,N_14939,N_14898);
nand UO_1313 (O_1313,N_14902,N_14928);
xor UO_1314 (O_1314,N_14915,N_14943);
xor UO_1315 (O_1315,N_14944,N_14919);
and UO_1316 (O_1316,N_14924,N_14880);
xnor UO_1317 (O_1317,N_14944,N_14912);
nand UO_1318 (O_1318,N_14937,N_14898);
xor UO_1319 (O_1319,N_14903,N_14905);
and UO_1320 (O_1320,N_14928,N_14966);
or UO_1321 (O_1321,N_14881,N_14909);
and UO_1322 (O_1322,N_14931,N_14947);
and UO_1323 (O_1323,N_14964,N_14969);
nand UO_1324 (O_1324,N_14899,N_14945);
nor UO_1325 (O_1325,N_14995,N_14950);
nor UO_1326 (O_1326,N_14972,N_14988);
xor UO_1327 (O_1327,N_14975,N_14935);
nand UO_1328 (O_1328,N_14967,N_14903);
nand UO_1329 (O_1329,N_14963,N_14990);
nor UO_1330 (O_1330,N_14929,N_14919);
xor UO_1331 (O_1331,N_14903,N_14940);
nor UO_1332 (O_1332,N_14905,N_14881);
and UO_1333 (O_1333,N_14887,N_14914);
or UO_1334 (O_1334,N_14970,N_14928);
and UO_1335 (O_1335,N_14997,N_14943);
xor UO_1336 (O_1336,N_14888,N_14900);
or UO_1337 (O_1337,N_14945,N_14995);
or UO_1338 (O_1338,N_14936,N_14902);
or UO_1339 (O_1339,N_14933,N_14955);
xor UO_1340 (O_1340,N_14903,N_14917);
and UO_1341 (O_1341,N_14992,N_14887);
or UO_1342 (O_1342,N_14916,N_14898);
and UO_1343 (O_1343,N_14968,N_14946);
nand UO_1344 (O_1344,N_14956,N_14962);
and UO_1345 (O_1345,N_14965,N_14998);
and UO_1346 (O_1346,N_14952,N_14990);
or UO_1347 (O_1347,N_14954,N_14908);
nand UO_1348 (O_1348,N_14903,N_14949);
nor UO_1349 (O_1349,N_14940,N_14982);
xor UO_1350 (O_1350,N_14914,N_14993);
or UO_1351 (O_1351,N_14907,N_14912);
or UO_1352 (O_1352,N_14958,N_14966);
xor UO_1353 (O_1353,N_14974,N_14912);
xnor UO_1354 (O_1354,N_14883,N_14910);
xor UO_1355 (O_1355,N_14990,N_14933);
and UO_1356 (O_1356,N_14965,N_14894);
nand UO_1357 (O_1357,N_14987,N_14892);
or UO_1358 (O_1358,N_14963,N_14921);
and UO_1359 (O_1359,N_14934,N_14987);
xnor UO_1360 (O_1360,N_14997,N_14968);
and UO_1361 (O_1361,N_14943,N_14964);
and UO_1362 (O_1362,N_14988,N_14931);
and UO_1363 (O_1363,N_14999,N_14987);
and UO_1364 (O_1364,N_14950,N_14976);
and UO_1365 (O_1365,N_14886,N_14909);
xnor UO_1366 (O_1366,N_14930,N_14940);
xor UO_1367 (O_1367,N_14974,N_14981);
xnor UO_1368 (O_1368,N_14915,N_14994);
or UO_1369 (O_1369,N_14974,N_14978);
and UO_1370 (O_1370,N_14884,N_14932);
xor UO_1371 (O_1371,N_14988,N_14913);
or UO_1372 (O_1372,N_14912,N_14941);
nand UO_1373 (O_1373,N_14998,N_14966);
nand UO_1374 (O_1374,N_14983,N_14885);
and UO_1375 (O_1375,N_14977,N_14927);
and UO_1376 (O_1376,N_14950,N_14917);
or UO_1377 (O_1377,N_14957,N_14976);
xor UO_1378 (O_1378,N_14918,N_14903);
nor UO_1379 (O_1379,N_14934,N_14904);
nand UO_1380 (O_1380,N_14917,N_14994);
xnor UO_1381 (O_1381,N_14899,N_14946);
and UO_1382 (O_1382,N_14979,N_14907);
nand UO_1383 (O_1383,N_14921,N_14924);
or UO_1384 (O_1384,N_14957,N_14886);
or UO_1385 (O_1385,N_14884,N_14914);
xnor UO_1386 (O_1386,N_14929,N_14901);
xor UO_1387 (O_1387,N_14905,N_14923);
xor UO_1388 (O_1388,N_14883,N_14876);
or UO_1389 (O_1389,N_14920,N_14894);
and UO_1390 (O_1390,N_14959,N_14887);
or UO_1391 (O_1391,N_14942,N_14943);
nand UO_1392 (O_1392,N_14908,N_14956);
nor UO_1393 (O_1393,N_14893,N_14980);
or UO_1394 (O_1394,N_14996,N_14897);
xor UO_1395 (O_1395,N_14984,N_14967);
nor UO_1396 (O_1396,N_14958,N_14917);
or UO_1397 (O_1397,N_14966,N_14970);
nand UO_1398 (O_1398,N_14987,N_14970);
xnor UO_1399 (O_1399,N_14909,N_14995);
and UO_1400 (O_1400,N_14950,N_14968);
and UO_1401 (O_1401,N_14897,N_14890);
nor UO_1402 (O_1402,N_14980,N_14899);
xnor UO_1403 (O_1403,N_14920,N_14976);
nand UO_1404 (O_1404,N_14960,N_14956);
and UO_1405 (O_1405,N_14904,N_14969);
xnor UO_1406 (O_1406,N_14999,N_14974);
nor UO_1407 (O_1407,N_14877,N_14970);
xor UO_1408 (O_1408,N_14995,N_14994);
nand UO_1409 (O_1409,N_14920,N_14960);
and UO_1410 (O_1410,N_14890,N_14971);
and UO_1411 (O_1411,N_14912,N_14961);
xnor UO_1412 (O_1412,N_14971,N_14983);
nand UO_1413 (O_1413,N_14917,N_14882);
nor UO_1414 (O_1414,N_14901,N_14990);
nor UO_1415 (O_1415,N_14989,N_14918);
and UO_1416 (O_1416,N_14952,N_14911);
nand UO_1417 (O_1417,N_14973,N_14904);
nand UO_1418 (O_1418,N_14880,N_14897);
xnor UO_1419 (O_1419,N_14973,N_14920);
xnor UO_1420 (O_1420,N_14880,N_14947);
and UO_1421 (O_1421,N_14892,N_14927);
nor UO_1422 (O_1422,N_14927,N_14951);
nand UO_1423 (O_1423,N_14915,N_14962);
xnor UO_1424 (O_1424,N_14955,N_14947);
nand UO_1425 (O_1425,N_14926,N_14900);
or UO_1426 (O_1426,N_14911,N_14879);
or UO_1427 (O_1427,N_14941,N_14945);
and UO_1428 (O_1428,N_14878,N_14995);
or UO_1429 (O_1429,N_14944,N_14964);
or UO_1430 (O_1430,N_14963,N_14938);
or UO_1431 (O_1431,N_14991,N_14947);
nand UO_1432 (O_1432,N_14947,N_14973);
nand UO_1433 (O_1433,N_14974,N_14895);
nor UO_1434 (O_1434,N_14926,N_14891);
nand UO_1435 (O_1435,N_14899,N_14936);
nor UO_1436 (O_1436,N_14948,N_14882);
nand UO_1437 (O_1437,N_14972,N_14997);
or UO_1438 (O_1438,N_14895,N_14892);
xnor UO_1439 (O_1439,N_14983,N_14951);
xor UO_1440 (O_1440,N_14919,N_14881);
xor UO_1441 (O_1441,N_14894,N_14908);
or UO_1442 (O_1442,N_14935,N_14978);
xor UO_1443 (O_1443,N_14924,N_14992);
and UO_1444 (O_1444,N_14989,N_14903);
nor UO_1445 (O_1445,N_14935,N_14934);
nor UO_1446 (O_1446,N_14915,N_14999);
or UO_1447 (O_1447,N_14951,N_14911);
xnor UO_1448 (O_1448,N_14906,N_14950);
and UO_1449 (O_1449,N_14945,N_14887);
and UO_1450 (O_1450,N_14965,N_14946);
xnor UO_1451 (O_1451,N_14946,N_14937);
and UO_1452 (O_1452,N_14943,N_14880);
and UO_1453 (O_1453,N_14933,N_14993);
nand UO_1454 (O_1454,N_14943,N_14897);
and UO_1455 (O_1455,N_14922,N_14989);
and UO_1456 (O_1456,N_14948,N_14884);
and UO_1457 (O_1457,N_14891,N_14986);
xnor UO_1458 (O_1458,N_14949,N_14912);
nand UO_1459 (O_1459,N_14936,N_14896);
xnor UO_1460 (O_1460,N_14961,N_14996);
and UO_1461 (O_1461,N_14973,N_14960);
or UO_1462 (O_1462,N_14959,N_14914);
or UO_1463 (O_1463,N_14941,N_14981);
xor UO_1464 (O_1464,N_14995,N_14939);
nor UO_1465 (O_1465,N_14973,N_14965);
nand UO_1466 (O_1466,N_14959,N_14921);
or UO_1467 (O_1467,N_14924,N_14936);
nor UO_1468 (O_1468,N_14941,N_14980);
or UO_1469 (O_1469,N_14933,N_14984);
xnor UO_1470 (O_1470,N_14908,N_14968);
or UO_1471 (O_1471,N_14895,N_14953);
nand UO_1472 (O_1472,N_14885,N_14933);
or UO_1473 (O_1473,N_14899,N_14923);
xor UO_1474 (O_1474,N_14959,N_14964);
nor UO_1475 (O_1475,N_14897,N_14889);
xor UO_1476 (O_1476,N_14923,N_14916);
or UO_1477 (O_1477,N_14956,N_14919);
or UO_1478 (O_1478,N_14983,N_14893);
nand UO_1479 (O_1479,N_14975,N_14956);
nor UO_1480 (O_1480,N_14887,N_14989);
and UO_1481 (O_1481,N_14932,N_14898);
and UO_1482 (O_1482,N_14974,N_14991);
and UO_1483 (O_1483,N_14911,N_14985);
or UO_1484 (O_1484,N_14961,N_14900);
or UO_1485 (O_1485,N_14947,N_14967);
nand UO_1486 (O_1486,N_14992,N_14936);
or UO_1487 (O_1487,N_14972,N_14887);
nand UO_1488 (O_1488,N_14979,N_14981);
xnor UO_1489 (O_1489,N_14935,N_14898);
nor UO_1490 (O_1490,N_14898,N_14970);
or UO_1491 (O_1491,N_14887,N_14985);
and UO_1492 (O_1492,N_14888,N_14987);
and UO_1493 (O_1493,N_14888,N_14952);
nand UO_1494 (O_1494,N_14892,N_14978);
or UO_1495 (O_1495,N_14978,N_14969);
nor UO_1496 (O_1496,N_14947,N_14969);
or UO_1497 (O_1497,N_14970,N_14953);
and UO_1498 (O_1498,N_14946,N_14960);
xnor UO_1499 (O_1499,N_14911,N_14959);
or UO_1500 (O_1500,N_14931,N_14962);
and UO_1501 (O_1501,N_14904,N_14927);
nand UO_1502 (O_1502,N_14957,N_14919);
and UO_1503 (O_1503,N_14998,N_14931);
nand UO_1504 (O_1504,N_14953,N_14964);
nand UO_1505 (O_1505,N_14987,N_14998);
xor UO_1506 (O_1506,N_14878,N_14968);
or UO_1507 (O_1507,N_14991,N_14890);
nor UO_1508 (O_1508,N_14940,N_14989);
nand UO_1509 (O_1509,N_14899,N_14898);
nand UO_1510 (O_1510,N_14878,N_14930);
and UO_1511 (O_1511,N_14906,N_14924);
and UO_1512 (O_1512,N_14978,N_14890);
nand UO_1513 (O_1513,N_14888,N_14969);
nor UO_1514 (O_1514,N_14898,N_14891);
nor UO_1515 (O_1515,N_14895,N_14908);
xor UO_1516 (O_1516,N_14963,N_14999);
xnor UO_1517 (O_1517,N_14927,N_14895);
xor UO_1518 (O_1518,N_14982,N_14893);
or UO_1519 (O_1519,N_14917,N_14931);
nor UO_1520 (O_1520,N_14964,N_14927);
nor UO_1521 (O_1521,N_14964,N_14995);
nor UO_1522 (O_1522,N_14999,N_14966);
xnor UO_1523 (O_1523,N_14907,N_14893);
nor UO_1524 (O_1524,N_14891,N_14921);
xor UO_1525 (O_1525,N_14981,N_14953);
and UO_1526 (O_1526,N_14902,N_14918);
and UO_1527 (O_1527,N_14926,N_14878);
nand UO_1528 (O_1528,N_14986,N_14914);
nor UO_1529 (O_1529,N_14929,N_14906);
xor UO_1530 (O_1530,N_14880,N_14917);
and UO_1531 (O_1531,N_14963,N_14987);
xnor UO_1532 (O_1532,N_14892,N_14952);
or UO_1533 (O_1533,N_14915,N_14997);
or UO_1534 (O_1534,N_14982,N_14898);
nor UO_1535 (O_1535,N_14939,N_14997);
and UO_1536 (O_1536,N_14881,N_14942);
nor UO_1537 (O_1537,N_14967,N_14907);
and UO_1538 (O_1538,N_14990,N_14897);
xnor UO_1539 (O_1539,N_14889,N_14985);
and UO_1540 (O_1540,N_14965,N_14930);
or UO_1541 (O_1541,N_14997,N_14922);
and UO_1542 (O_1542,N_14969,N_14955);
nor UO_1543 (O_1543,N_14976,N_14996);
xor UO_1544 (O_1544,N_14892,N_14897);
xor UO_1545 (O_1545,N_14924,N_14932);
nand UO_1546 (O_1546,N_14917,N_14978);
nor UO_1547 (O_1547,N_14983,N_14892);
xor UO_1548 (O_1548,N_14979,N_14991);
or UO_1549 (O_1549,N_14918,N_14894);
nor UO_1550 (O_1550,N_14912,N_14926);
xor UO_1551 (O_1551,N_14943,N_14893);
xor UO_1552 (O_1552,N_14998,N_14922);
or UO_1553 (O_1553,N_14898,N_14908);
nor UO_1554 (O_1554,N_14977,N_14972);
or UO_1555 (O_1555,N_14976,N_14908);
xnor UO_1556 (O_1556,N_14927,N_14986);
nor UO_1557 (O_1557,N_14898,N_14910);
xnor UO_1558 (O_1558,N_14927,N_14945);
xor UO_1559 (O_1559,N_14961,N_14988);
and UO_1560 (O_1560,N_14994,N_14997);
nand UO_1561 (O_1561,N_14911,N_14913);
and UO_1562 (O_1562,N_14951,N_14995);
xor UO_1563 (O_1563,N_14951,N_14970);
or UO_1564 (O_1564,N_14895,N_14884);
or UO_1565 (O_1565,N_14956,N_14993);
nor UO_1566 (O_1566,N_14879,N_14997);
xor UO_1567 (O_1567,N_14949,N_14987);
and UO_1568 (O_1568,N_14883,N_14903);
xor UO_1569 (O_1569,N_14955,N_14965);
xor UO_1570 (O_1570,N_14934,N_14999);
nand UO_1571 (O_1571,N_14879,N_14999);
xnor UO_1572 (O_1572,N_14894,N_14909);
or UO_1573 (O_1573,N_14918,N_14976);
and UO_1574 (O_1574,N_14953,N_14923);
nor UO_1575 (O_1575,N_14979,N_14934);
xor UO_1576 (O_1576,N_14935,N_14980);
nand UO_1577 (O_1577,N_14923,N_14948);
nor UO_1578 (O_1578,N_14933,N_14968);
nand UO_1579 (O_1579,N_14896,N_14907);
and UO_1580 (O_1580,N_14958,N_14998);
nor UO_1581 (O_1581,N_14990,N_14996);
xor UO_1582 (O_1582,N_14924,N_14981);
or UO_1583 (O_1583,N_14899,N_14979);
nor UO_1584 (O_1584,N_14997,N_14954);
xnor UO_1585 (O_1585,N_14964,N_14945);
nand UO_1586 (O_1586,N_14894,N_14981);
nor UO_1587 (O_1587,N_14922,N_14976);
xor UO_1588 (O_1588,N_14990,N_14958);
nand UO_1589 (O_1589,N_14907,N_14984);
and UO_1590 (O_1590,N_14906,N_14889);
xnor UO_1591 (O_1591,N_14898,N_14972);
nor UO_1592 (O_1592,N_14885,N_14954);
nor UO_1593 (O_1593,N_14916,N_14924);
nor UO_1594 (O_1594,N_14887,N_14955);
nor UO_1595 (O_1595,N_14935,N_14885);
and UO_1596 (O_1596,N_14956,N_14969);
or UO_1597 (O_1597,N_14916,N_14921);
nand UO_1598 (O_1598,N_14885,N_14940);
nor UO_1599 (O_1599,N_14892,N_14929);
xor UO_1600 (O_1600,N_14968,N_14998);
xnor UO_1601 (O_1601,N_14988,N_14909);
nor UO_1602 (O_1602,N_14976,N_14899);
xnor UO_1603 (O_1603,N_14922,N_14924);
nor UO_1604 (O_1604,N_14927,N_14941);
nand UO_1605 (O_1605,N_14938,N_14947);
and UO_1606 (O_1606,N_14983,N_14895);
or UO_1607 (O_1607,N_14906,N_14968);
and UO_1608 (O_1608,N_14897,N_14919);
and UO_1609 (O_1609,N_14977,N_14984);
nand UO_1610 (O_1610,N_14993,N_14898);
or UO_1611 (O_1611,N_14965,N_14922);
xnor UO_1612 (O_1612,N_14985,N_14878);
nor UO_1613 (O_1613,N_14955,N_14904);
or UO_1614 (O_1614,N_14897,N_14920);
or UO_1615 (O_1615,N_14937,N_14973);
nand UO_1616 (O_1616,N_14875,N_14890);
and UO_1617 (O_1617,N_14948,N_14979);
and UO_1618 (O_1618,N_14972,N_14875);
nor UO_1619 (O_1619,N_14898,N_14973);
or UO_1620 (O_1620,N_14970,N_14945);
and UO_1621 (O_1621,N_14982,N_14924);
or UO_1622 (O_1622,N_14907,N_14894);
or UO_1623 (O_1623,N_14975,N_14893);
or UO_1624 (O_1624,N_14987,N_14921);
or UO_1625 (O_1625,N_14893,N_14920);
nor UO_1626 (O_1626,N_14959,N_14904);
xnor UO_1627 (O_1627,N_14910,N_14939);
and UO_1628 (O_1628,N_14912,N_14991);
and UO_1629 (O_1629,N_14926,N_14970);
and UO_1630 (O_1630,N_14901,N_14935);
xnor UO_1631 (O_1631,N_14993,N_14920);
nor UO_1632 (O_1632,N_14957,N_14891);
nand UO_1633 (O_1633,N_14999,N_14887);
nor UO_1634 (O_1634,N_14947,N_14926);
nand UO_1635 (O_1635,N_14962,N_14976);
xnor UO_1636 (O_1636,N_14941,N_14896);
and UO_1637 (O_1637,N_14938,N_14987);
nand UO_1638 (O_1638,N_14936,N_14974);
nand UO_1639 (O_1639,N_14973,N_14899);
and UO_1640 (O_1640,N_14994,N_14981);
or UO_1641 (O_1641,N_14916,N_14886);
and UO_1642 (O_1642,N_14992,N_14877);
nand UO_1643 (O_1643,N_14951,N_14940);
and UO_1644 (O_1644,N_14916,N_14957);
and UO_1645 (O_1645,N_14894,N_14916);
xor UO_1646 (O_1646,N_14968,N_14896);
and UO_1647 (O_1647,N_14963,N_14970);
nand UO_1648 (O_1648,N_14963,N_14936);
xor UO_1649 (O_1649,N_14957,N_14988);
xnor UO_1650 (O_1650,N_14971,N_14967);
nor UO_1651 (O_1651,N_14954,N_14950);
or UO_1652 (O_1652,N_14973,N_14923);
or UO_1653 (O_1653,N_14993,N_14948);
xnor UO_1654 (O_1654,N_14934,N_14897);
nand UO_1655 (O_1655,N_14897,N_14957);
and UO_1656 (O_1656,N_14929,N_14902);
and UO_1657 (O_1657,N_14949,N_14939);
xnor UO_1658 (O_1658,N_14877,N_14921);
or UO_1659 (O_1659,N_14893,N_14919);
and UO_1660 (O_1660,N_14998,N_14882);
xnor UO_1661 (O_1661,N_14954,N_14894);
and UO_1662 (O_1662,N_14882,N_14983);
and UO_1663 (O_1663,N_14899,N_14995);
and UO_1664 (O_1664,N_14965,N_14932);
xor UO_1665 (O_1665,N_14941,N_14908);
xor UO_1666 (O_1666,N_14929,N_14997);
nand UO_1667 (O_1667,N_14882,N_14889);
and UO_1668 (O_1668,N_14957,N_14938);
nor UO_1669 (O_1669,N_14980,N_14894);
and UO_1670 (O_1670,N_14898,N_14941);
nand UO_1671 (O_1671,N_14889,N_14891);
xor UO_1672 (O_1672,N_14995,N_14914);
and UO_1673 (O_1673,N_14992,N_14897);
nor UO_1674 (O_1674,N_14877,N_14948);
nand UO_1675 (O_1675,N_14907,N_14888);
and UO_1676 (O_1676,N_14877,N_14983);
and UO_1677 (O_1677,N_14920,N_14889);
xnor UO_1678 (O_1678,N_14887,N_14994);
and UO_1679 (O_1679,N_14919,N_14887);
and UO_1680 (O_1680,N_14928,N_14914);
nand UO_1681 (O_1681,N_14975,N_14928);
xnor UO_1682 (O_1682,N_14964,N_14903);
and UO_1683 (O_1683,N_14921,N_14886);
xnor UO_1684 (O_1684,N_14954,N_14925);
xnor UO_1685 (O_1685,N_14891,N_14933);
and UO_1686 (O_1686,N_14908,N_14938);
nor UO_1687 (O_1687,N_14984,N_14994);
nor UO_1688 (O_1688,N_14999,N_14945);
nand UO_1689 (O_1689,N_14903,N_14994);
or UO_1690 (O_1690,N_14913,N_14964);
xnor UO_1691 (O_1691,N_14922,N_14949);
nor UO_1692 (O_1692,N_14934,N_14948);
nand UO_1693 (O_1693,N_14901,N_14914);
nor UO_1694 (O_1694,N_14882,N_14952);
nor UO_1695 (O_1695,N_14983,N_14940);
and UO_1696 (O_1696,N_14901,N_14922);
and UO_1697 (O_1697,N_14885,N_14887);
nand UO_1698 (O_1698,N_14883,N_14953);
and UO_1699 (O_1699,N_14926,N_14923);
nor UO_1700 (O_1700,N_14977,N_14914);
nor UO_1701 (O_1701,N_14953,N_14876);
nand UO_1702 (O_1702,N_14951,N_14996);
xnor UO_1703 (O_1703,N_14970,N_14907);
xnor UO_1704 (O_1704,N_14924,N_14958);
nand UO_1705 (O_1705,N_14977,N_14891);
and UO_1706 (O_1706,N_14906,N_14920);
or UO_1707 (O_1707,N_14960,N_14934);
nand UO_1708 (O_1708,N_14977,N_14954);
or UO_1709 (O_1709,N_14887,N_14932);
or UO_1710 (O_1710,N_14940,N_14975);
and UO_1711 (O_1711,N_14882,N_14972);
xnor UO_1712 (O_1712,N_14960,N_14970);
nor UO_1713 (O_1713,N_14993,N_14949);
nand UO_1714 (O_1714,N_14971,N_14985);
or UO_1715 (O_1715,N_14982,N_14881);
nand UO_1716 (O_1716,N_14978,N_14968);
or UO_1717 (O_1717,N_14992,N_14959);
xnor UO_1718 (O_1718,N_14990,N_14928);
nand UO_1719 (O_1719,N_14928,N_14944);
or UO_1720 (O_1720,N_14930,N_14907);
nor UO_1721 (O_1721,N_14878,N_14993);
nand UO_1722 (O_1722,N_14986,N_14963);
nor UO_1723 (O_1723,N_14933,N_14951);
nor UO_1724 (O_1724,N_14928,N_14976);
xnor UO_1725 (O_1725,N_14959,N_14963);
and UO_1726 (O_1726,N_14987,N_14940);
or UO_1727 (O_1727,N_14971,N_14962);
nand UO_1728 (O_1728,N_14885,N_14941);
xor UO_1729 (O_1729,N_14948,N_14959);
nand UO_1730 (O_1730,N_14966,N_14888);
or UO_1731 (O_1731,N_14972,N_14951);
or UO_1732 (O_1732,N_14925,N_14906);
and UO_1733 (O_1733,N_14919,N_14949);
xnor UO_1734 (O_1734,N_14906,N_14877);
xnor UO_1735 (O_1735,N_14932,N_14907);
nor UO_1736 (O_1736,N_14881,N_14966);
or UO_1737 (O_1737,N_14947,N_14996);
xnor UO_1738 (O_1738,N_14960,N_14911);
or UO_1739 (O_1739,N_14954,N_14922);
nand UO_1740 (O_1740,N_14912,N_14989);
nand UO_1741 (O_1741,N_14941,N_14894);
or UO_1742 (O_1742,N_14971,N_14884);
xor UO_1743 (O_1743,N_14957,N_14973);
nor UO_1744 (O_1744,N_14875,N_14922);
nor UO_1745 (O_1745,N_14932,N_14979);
xnor UO_1746 (O_1746,N_14890,N_14921);
nor UO_1747 (O_1747,N_14925,N_14900);
nor UO_1748 (O_1748,N_14961,N_14904);
nand UO_1749 (O_1749,N_14904,N_14885);
or UO_1750 (O_1750,N_14962,N_14900);
nor UO_1751 (O_1751,N_14955,N_14967);
nand UO_1752 (O_1752,N_14899,N_14950);
and UO_1753 (O_1753,N_14980,N_14963);
and UO_1754 (O_1754,N_14976,N_14973);
and UO_1755 (O_1755,N_14949,N_14975);
or UO_1756 (O_1756,N_14881,N_14884);
and UO_1757 (O_1757,N_14966,N_14917);
or UO_1758 (O_1758,N_14968,N_14942);
or UO_1759 (O_1759,N_14880,N_14905);
and UO_1760 (O_1760,N_14914,N_14892);
nor UO_1761 (O_1761,N_14893,N_14898);
or UO_1762 (O_1762,N_14967,N_14880);
or UO_1763 (O_1763,N_14966,N_14948);
or UO_1764 (O_1764,N_14932,N_14990);
nor UO_1765 (O_1765,N_14897,N_14899);
nor UO_1766 (O_1766,N_14964,N_14891);
xor UO_1767 (O_1767,N_14891,N_14984);
or UO_1768 (O_1768,N_14946,N_14892);
or UO_1769 (O_1769,N_14894,N_14887);
nand UO_1770 (O_1770,N_14933,N_14915);
nor UO_1771 (O_1771,N_14898,N_14931);
and UO_1772 (O_1772,N_14918,N_14949);
xnor UO_1773 (O_1773,N_14940,N_14965);
or UO_1774 (O_1774,N_14922,N_14898);
and UO_1775 (O_1775,N_14886,N_14954);
and UO_1776 (O_1776,N_14923,N_14911);
nand UO_1777 (O_1777,N_14985,N_14957);
xor UO_1778 (O_1778,N_14975,N_14905);
nand UO_1779 (O_1779,N_14916,N_14988);
or UO_1780 (O_1780,N_14918,N_14998);
xor UO_1781 (O_1781,N_14886,N_14931);
xnor UO_1782 (O_1782,N_14882,N_14901);
and UO_1783 (O_1783,N_14930,N_14957);
xnor UO_1784 (O_1784,N_14992,N_14918);
nor UO_1785 (O_1785,N_14876,N_14943);
or UO_1786 (O_1786,N_14993,N_14927);
nor UO_1787 (O_1787,N_14962,N_14894);
xnor UO_1788 (O_1788,N_14977,N_14997);
and UO_1789 (O_1789,N_14992,N_14938);
nor UO_1790 (O_1790,N_14974,N_14975);
nand UO_1791 (O_1791,N_14995,N_14987);
nor UO_1792 (O_1792,N_14911,N_14908);
or UO_1793 (O_1793,N_14979,N_14904);
and UO_1794 (O_1794,N_14978,N_14997);
nor UO_1795 (O_1795,N_14991,N_14960);
nand UO_1796 (O_1796,N_14935,N_14910);
xnor UO_1797 (O_1797,N_14891,N_14943);
nand UO_1798 (O_1798,N_14980,N_14947);
xnor UO_1799 (O_1799,N_14877,N_14928);
and UO_1800 (O_1800,N_14989,N_14964);
xor UO_1801 (O_1801,N_14888,N_14963);
nor UO_1802 (O_1802,N_14926,N_14991);
or UO_1803 (O_1803,N_14958,N_14965);
nand UO_1804 (O_1804,N_14921,N_14953);
xor UO_1805 (O_1805,N_14960,N_14974);
or UO_1806 (O_1806,N_14913,N_14877);
xor UO_1807 (O_1807,N_14977,N_14998);
or UO_1808 (O_1808,N_14980,N_14891);
nand UO_1809 (O_1809,N_14960,N_14899);
and UO_1810 (O_1810,N_14911,N_14885);
xor UO_1811 (O_1811,N_14953,N_14938);
and UO_1812 (O_1812,N_14931,N_14974);
and UO_1813 (O_1813,N_14934,N_14950);
or UO_1814 (O_1814,N_14978,N_14915);
nor UO_1815 (O_1815,N_14903,N_14945);
nand UO_1816 (O_1816,N_14977,N_14973);
nand UO_1817 (O_1817,N_14943,N_14973);
nor UO_1818 (O_1818,N_14881,N_14914);
xnor UO_1819 (O_1819,N_14875,N_14990);
xor UO_1820 (O_1820,N_14937,N_14989);
and UO_1821 (O_1821,N_14899,N_14895);
nand UO_1822 (O_1822,N_14971,N_14899);
or UO_1823 (O_1823,N_14905,N_14890);
nand UO_1824 (O_1824,N_14997,N_14903);
nand UO_1825 (O_1825,N_14932,N_14886);
xnor UO_1826 (O_1826,N_14937,N_14892);
nor UO_1827 (O_1827,N_14928,N_14950);
or UO_1828 (O_1828,N_14891,N_14922);
nand UO_1829 (O_1829,N_14952,N_14994);
nor UO_1830 (O_1830,N_14931,N_14979);
nor UO_1831 (O_1831,N_14911,N_14881);
xnor UO_1832 (O_1832,N_14984,N_14919);
xnor UO_1833 (O_1833,N_14960,N_14893);
and UO_1834 (O_1834,N_14878,N_14990);
or UO_1835 (O_1835,N_14936,N_14934);
nand UO_1836 (O_1836,N_14964,N_14924);
xor UO_1837 (O_1837,N_14943,N_14912);
or UO_1838 (O_1838,N_14930,N_14958);
nand UO_1839 (O_1839,N_14909,N_14967);
xor UO_1840 (O_1840,N_14919,N_14974);
or UO_1841 (O_1841,N_14906,N_14930);
and UO_1842 (O_1842,N_14951,N_14964);
and UO_1843 (O_1843,N_14933,N_14883);
and UO_1844 (O_1844,N_14948,N_14946);
nand UO_1845 (O_1845,N_14928,N_14948);
nor UO_1846 (O_1846,N_14909,N_14975);
and UO_1847 (O_1847,N_14943,N_14883);
nor UO_1848 (O_1848,N_14886,N_14999);
or UO_1849 (O_1849,N_14953,N_14935);
or UO_1850 (O_1850,N_14976,N_14988);
and UO_1851 (O_1851,N_14891,N_14907);
or UO_1852 (O_1852,N_14918,N_14887);
or UO_1853 (O_1853,N_14944,N_14948);
nand UO_1854 (O_1854,N_14913,N_14896);
or UO_1855 (O_1855,N_14959,N_14875);
nor UO_1856 (O_1856,N_14914,N_14924);
xor UO_1857 (O_1857,N_14993,N_14997);
nor UO_1858 (O_1858,N_14909,N_14945);
or UO_1859 (O_1859,N_14932,N_14968);
or UO_1860 (O_1860,N_14975,N_14933);
or UO_1861 (O_1861,N_14925,N_14876);
nand UO_1862 (O_1862,N_14939,N_14914);
nor UO_1863 (O_1863,N_14886,N_14942);
xnor UO_1864 (O_1864,N_14896,N_14956);
nor UO_1865 (O_1865,N_14927,N_14979);
or UO_1866 (O_1866,N_14891,N_14892);
nor UO_1867 (O_1867,N_14885,N_14875);
nor UO_1868 (O_1868,N_14932,N_14969);
nand UO_1869 (O_1869,N_14969,N_14876);
nand UO_1870 (O_1870,N_14966,N_14961);
and UO_1871 (O_1871,N_14913,N_14942);
xnor UO_1872 (O_1872,N_14989,N_14984);
nor UO_1873 (O_1873,N_14910,N_14876);
and UO_1874 (O_1874,N_14997,N_14911);
and UO_1875 (O_1875,N_14875,N_14938);
nand UO_1876 (O_1876,N_14975,N_14927);
xnor UO_1877 (O_1877,N_14997,N_14914);
or UO_1878 (O_1878,N_14963,N_14900);
nor UO_1879 (O_1879,N_14923,N_14889);
xor UO_1880 (O_1880,N_14953,N_14971);
nand UO_1881 (O_1881,N_14925,N_14969);
xnor UO_1882 (O_1882,N_14938,N_14980);
or UO_1883 (O_1883,N_14980,N_14948);
xnor UO_1884 (O_1884,N_14909,N_14952);
nor UO_1885 (O_1885,N_14985,N_14875);
nand UO_1886 (O_1886,N_14911,N_14948);
xor UO_1887 (O_1887,N_14921,N_14896);
or UO_1888 (O_1888,N_14951,N_14913);
or UO_1889 (O_1889,N_14991,N_14967);
or UO_1890 (O_1890,N_14943,N_14925);
nor UO_1891 (O_1891,N_14920,N_14936);
nor UO_1892 (O_1892,N_14998,N_14981);
and UO_1893 (O_1893,N_14999,N_14986);
nand UO_1894 (O_1894,N_14962,N_14916);
nor UO_1895 (O_1895,N_14902,N_14887);
xnor UO_1896 (O_1896,N_14914,N_14954);
nor UO_1897 (O_1897,N_14969,N_14889);
xor UO_1898 (O_1898,N_14988,N_14984);
xnor UO_1899 (O_1899,N_14952,N_14991);
nor UO_1900 (O_1900,N_14900,N_14998);
nor UO_1901 (O_1901,N_14906,N_14948);
or UO_1902 (O_1902,N_14944,N_14965);
or UO_1903 (O_1903,N_14875,N_14960);
nor UO_1904 (O_1904,N_14995,N_14999);
or UO_1905 (O_1905,N_14950,N_14937);
or UO_1906 (O_1906,N_14962,N_14904);
or UO_1907 (O_1907,N_14920,N_14961);
or UO_1908 (O_1908,N_14906,N_14957);
and UO_1909 (O_1909,N_14958,N_14907);
xnor UO_1910 (O_1910,N_14939,N_14938);
xnor UO_1911 (O_1911,N_14948,N_14953);
nor UO_1912 (O_1912,N_14941,N_14907);
nor UO_1913 (O_1913,N_14990,N_14968);
or UO_1914 (O_1914,N_14968,N_14912);
xor UO_1915 (O_1915,N_14878,N_14909);
or UO_1916 (O_1916,N_14995,N_14953);
and UO_1917 (O_1917,N_14957,N_14903);
nor UO_1918 (O_1918,N_14956,N_14933);
or UO_1919 (O_1919,N_14976,N_14953);
xor UO_1920 (O_1920,N_14995,N_14933);
nand UO_1921 (O_1921,N_14944,N_14920);
nor UO_1922 (O_1922,N_14957,N_14884);
nand UO_1923 (O_1923,N_14955,N_14972);
xor UO_1924 (O_1924,N_14875,N_14989);
nor UO_1925 (O_1925,N_14928,N_14949);
and UO_1926 (O_1926,N_14927,N_14971);
and UO_1927 (O_1927,N_14955,N_14942);
or UO_1928 (O_1928,N_14888,N_14973);
and UO_1929 (O_1929,N_14898,N_14903);
or UO_1930 (O_1930,N_14947,N_14974);
xor UO_1931 (O_1931,N_14970,N_14972);
and UO_1932 (O_1932,N_14931,N_14991);
nand UO_1933 (O_1933,N_14914,N_14938);
nor UO_1934 (O_1934,N_14990,N_14926);
xnor UO_1935 (O_1935,N_14890,N_14885);
xor UO_1936 (O_1936,N_14957,N_14875);
and UO_1937 (O_1937,N_14925,N_14892);
nor UO_1938 (O_1938,N_14904,N_14975);
or UO_1939 (O_1939,N_14920,N_14979);
or UO_1940 (O_1940,N_14999,N_14895);
xor UO_1941 (O_1941,N_14911,N_14926);
xor UO_1942 (O_1942,N_14970,N_14916);
xor UO_1943 (O_1943,N_14920,N_14982);
and UO_1944 (O_1944,N_14963,N_14915);
nand UO_1945 (O_1945,N_14969,N_14961);
and UO_1946 (O_1946,N_14913,N_14930);
or UO_1947 (O_1947,N_14999,N_14946);
nand UO_1948 (O_1948,N_14960,N_14982);
nor UO_1949 (O_1949,N_14967,N_14957);
and UO_1950 (O_1950,N_14971,N_14941);
nand UO_1951 (O_1951,N_14979,N_14887);
xnor UO_1952 (O_1952,N_14893,N_14914);
or UO_1953 (O_1953,N_14996,N_14953);
nor UO_1954 (O_1954,N_14904,N_14907);
xnor UO_1955 (O_1955,N_14957,N_14970);
or UO_1956 (O_1956,N_14931,N_14910);
or UO_1957 (O_1957,N_14930,N_14933);
nor UO_1958 (O_1958,N_14992,N_14895);
nand UO_1959 (O_1959,N_14907,N_14924);
nand UO_1960 (O_1960,N_14937,N_14943);
xnor UO_1961 (O_1961,N_14974,N_14930);
and UO_1962 (O_1962,N_14972,N_14996);
or UO_1963 (O_1963,N_14984,N_14898);
and UO_1964 (O_1964,N_14908,N_14883);
nand UO_1965 (O_1965,N_14908,N_14984);
nand UO_1966 (O_1966,N_14922,N_14893);
nor UO_1967 (O_1967,N_14974,N_14906);
nor UO_1968 (O_1968,N_14973,N_14962);
nor UO_1969 (O_1969,N_14948,N_14955);
or UO_1970 (O_1970,N_14904,N_14963);
nand UO_1971 (O_1971,N_14930,N_14903);
nand UO_1972 (O_1972,N_14966,N_14920);
xnor UO_1973 (O_1973,N_14982,N_14903);
xor UO_1974 (O_1974,N_14992,N_14935);
nor UO_1975 (O_1975,N_14931,N_14951);
and UO_1976 (O_1976,N_14883,N_14970);
nor UO_1977 (O_1977,N_14903,N_14928);
xor UO_1978 (O_1978,N_14917,N_14977);
or UO_1979 (O_1979,N_14949,N_14938);
nand UO_1980 (O_1980,N_14904,N_14901);
or UO_1981 (O_1981,N_14995,N_14980);
xnor UO_1982 (O_1982,N_14915,N_14928);
or UO_1983 (O_1983,N_14935,N_14927);
nor UO_1984 (O_1984,N_14980,N_14961);
and UO_1985 (O_1985,N_14909,N_14891);
xnor UO_1986 (O_1986,N_14927,N_14939);
or UO_1987 (O_1987,N_14975,N_14945);
xnor UO_1988 (O_1988,N_14930,N_14914);
nor UO_1989 (O_1989,N_14912,N_14925);
or UO_1990 (O_1990,N_14888,N_14970);
nor UO_1991 (O_1991,N_14926,N_14894);
nor UO_1992 (O_1992,N_14912,N_14950);
or UO_1993 (O_1993,N_14907,N_14917);
or UO_1994 (O_1994,N_14971,N_14988);
nor UO_1995 (O_1995,N_14934,N_14907);
xor UO_1996 (O_1996,N_14932,N_14953);
and UO_1997 (O_1997,N_14941,N_14944);
nand UO_1998 (O_1998,N_14944,N_14896);
and UO_1999 (O_1999,N_14881,N_14904);
endmodule