module basic_500_3000_500_50_levels_2xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_222,In_438);
nor U1 (N_1,In_147,In_345);
nor U2 (N_2,In_121,In_252);
and U3 (N_3,In_436,In_298);
nand U4 (N_4,In_233,In_212);
or U5 (N_5,In_17,In_208);
nand U6 (N_6,In_346,In_154);
xor U7 (N_7,In_482,In_397);
and U8 (N_8,In_465,In_267);
or U9 (N_9,In_162,In_423);
or U10 (N_10,In_83,In_125);
nor U11 (N_11,In_30,In_200);
and U12 (N_12,In_170,In_98);
and U13 (N_13,In_94,In_152);
and U14 (N_14,In_248,In_112);
xor U15 (N_15,In_54,In_488);
or U16 (N_16,In_241,In_366);
nand U17 (N_17,In_149,In_450);
nand U18 (N_18,In_281,In_424);
and U19 (N_19,In_19,In_431);
and U20 (N_20,In_9,In_275);
xor U21 (N_21,In_335,In_484);
nand U22 (N_22,In_184,In_257);
and U23 (N_23,In_317,In_109);
or U24 (N_24,In_140,In_115);
nor U25 (N_25,In_59,In_62);
nand U26 (N_26,In_455,In_81);
xnor U27 (N_27,In_35,In_290);
nor U28 (N_28,In_453,In_235);
nand U29 (N_29,In_202,In_4);
nor U30 (N_30,In_467,In_437);
nor U31 (N_31,In_21,In_119);
or U32 (N_32,In_60,In_64);
nor U33 (N_33,In_318,In_31);
nor U34 (N_34,In_263,In_176);
nand U35 (N_35,In_230,In_478);
nor U36 (N_36,In_144,In_320);
or U37 (N_37,In_280,In_404);
and U38 (N_38,In_487,In_11);
xnor U39 (N_39,In_292,In_414);
or U40 (N_40,In_143,In_429);
or U41 (N_41,In_495,In_169);
nand U42 (N_42,In_206,In_16);
nand U43 (N_43,In_387,In_293);
or U44 (N_44,In_354,In_457);
nand U45 (N_45,In_174,In_40);
xor U46 (N_46,In_390,In_371);
nor U47 (N_47,In_385,In_89);
or U48 (N_48,In_444,In_71);
or U49 (N_49,In_256,In_175);
or U50 (N_50,In_418,In_203);
nor U51 (N_51,In_427,In_462);
nor U52 (N_52,In_39,In_114);
or U53 (N_53,In_38,In_379);
nor U54 (N_54,In_351,In_168);
nor U55 (N_55,In_128,In_376);
nand U56 (N_56,In_461,In_349);
or U57 (N_57,In_157,In_215);
nor U58 (N_58,In_85,In_6);
and U59 (N_59,In_459,In_130);
nand U60 (N_60,In_244,In_245);
nor U61 (N_61,In_44,In_250);
xor U62 (N_62,In_211,In_166);
or U63 (N_63,In_363,In_118);
nand U64 (N_64,In_246,In_116);
and U65 (N_65,In_402,In_75);
nor U66 (N_66,In_122,In_391);
nor U67 (N_67,In_434,In_481);
nor U68 (N_68,In_111,In_13);
or U69 (N_69,In_260,N_0);
nand U70 (N_70,In_213,N_46);
nand U71 (N_71,In_441,In_494);
or U72 (N_72,In_289,In_229);
or U73 (N_73,N_43,N_9);
or U74 (N_74,In_56,In_113);
or U75 (N_75,In_8,In_433);
nand U76 (N_76,In_324,In_53);
nand U77 (N_77,In_463,In_350);
nor U78 (N_78,N_16,In_399);
nor U79 (N_79,N_59,In_356);
or U80 (N_80,In_348,In_172);
nand U81 (N_81,In_492,In_377);
nor U82 (N_82,In_406,In_447);
and U83 (N_83,In_384,In_160);
nor U84 (N_84,N_54,In_491);
nand U85 (N_85,In_332,In_150);
nand U86 (N_86,In_67,N_39);
or U87 (N_87,N_52,In_196);
and U88 (N_88,In_221,In_254);
nand U89 (N_89,In_37,In_417);
or U90 (N_90,In_278,In_55);
nor U91 (N_91,In_7,N_40);
nand U92 (N_92,In_271,In_133);
or U93 (N_93,In_104,In_338);
or U94 (N_94,In_291,In_234);
and U95 (N_95,In_117,In_473);
nor U96 (N_96,In_333,In_2);
nor U97 (N_97,In_32,In_153);
nand U98 (N_98,In_120,N_36);
xor U99 (N_99,In_177,In_41);
or U100 (N_100,In_309,In_102);
nor U101 (N_101,In_329,In_312);
nor U102 (N_102,In_23,In_425);
nand U103 (N_103,In_151,N_33);
nand U104 (N_104,In_28,In_321);
nor U105 (N_105,In_158,N_11);
and U106 (N_106,N_20,In_330);
nand U107 (N_107,N_26,In_472);
nor U108 (N_108,In_378,In_15);
nor U109 (N_109,In_58,In_322);
nor U110 (N_110,In_411,In_82);
nor U111 (N_111,In_258,In_276);
xnor U112 (N_112,In_136,In_355);
nor U113 (N_113,In_381,In_451);
nor U114 (N_114,In_323,In_311);
nand U115 (N_115,N_42,In_307);
or U116 (N_116,In_180,In_446);
or U117 (N_117,In_22,In_14);
nand U118 (N_118,In_480,In_420);
nor U119 (N_119,In_223,In_192);
nand U120 (N_120,N_24,N_15);
nor U121 (N_121,In_301,In_123);
and U122 (N_122,In_382,N_92);
and U123 (N_123,N_95,In_101);
nand U124 (N_124,In_242,N_99);
or U125 (N_125,In_489,In_392);
and U126 (N_126,N_115,In_443);
or U127 (N_127,In_1,In_238);
nor U128 (N_128,In_45,In_224);
and U129 (N_129,N_97,N_63);
nand U130 (N_130,In_181,In_262);
and U131 (N_131,In_264,In_156);
nand U132 (N_132,N_1,In_103);
nor U133 (N_133,In_398,In_148);
nor U134 (N_134,In_20,In_146);
or U135 (N_135,In_226,In_27);
or U136 (N_136,In_90,In_91);
nor U137 (N_137,N_41,N_58);
nand U138 (N_138,In_78,In_72);
or U139 (N_139,N_34,In_303);
or U140 (N_140,In_395,In_445);
nor U141 (N_141,In_442,N_98);
and U142 (N_142,In_225,In_483);
nor U143 (N_143,In_449,In_84);
nor U144 (N_144,In_372,In_97);
or U145 (N_145,In_132,In_24);
nor U146 (N_146,In_173,In_138);
nor U147 (N_147,In_409,In_400);
or U148 (N_148,In_485,In_458);
and U149 (N_149,N_69,N_14);
nand U150 (N_150,N_65,N_112);
nand U151 (N_151,In_369,In_195);
nor U152 (N_152,N_76,In_219);
nor U153 (N_153,N_103,In_426);
nor U154 (N_154,In_314,N_109);
xnor U155 (N_155,In_99,In_407);
nor U156 (N_156,In_209,In_336);
nand U157 (N_157,In_210,In_474);
and U158 (N_158,In_190,In_393);
and U159 (N_159,In_137,In_493);
and U160 (N_160,N_116,In_295);
nor U161 (N_161,In_204,In_183);
or U162 (N_162,In_305,N_7);
and U163 (N_163,In_316,In_340);
nor U164 (N_164,N_2,In_499);
and U165 (N_165,In_86,In_268);
and U166 (N_166,In_178,In_415);
and U167 (N_167,In_334,N_93);
nor U168 (N_168,In_77,In_161);
and U169 (N_169,N_110,In_331);
nand U170 (N_170,N_104,N_77);
nor U171 (N_171,N_72,In_454);
and U172 (N_172,In_105,N_81);
nand U173 (N_173,In_251,N_4);
nand U174 (N_174,In_341,In_42);
nand U175 (N_175,In_185,N_38);
and U176 (N_176,In_401,In_93);
and U177 (N_177,In_73,In_139);
nor U178 (N_178,In_218,In_421);
and U179 (N_179,In_142,In_496);
or U180 (N_180,N_29,In_106);
or U181 (N_181,In_359,N_133);
nand U182 (N_182,N_83,N_27);
nor U183 (N_183,In_70,N_144);
or U184 (N_184,N_66,In_205);
nand U185 (N_185,N_96,N_113);
nor U186 (N_186,In_279,In_422);
or U187 (N_187,N_161,In_327);
or U188 (N_188,N_114,In_273);
and U189 (N_189,In_88,In_325);
and U190 (N_190,In_300,N_145);
or U191 (N_191,In_48,In_237);
and U192 (N_192,In_383,In_339);
nand U193 (N_193,In_274,N_19);
nand U194 (N_194,In_107,N_118);
nor U195 (N_195,In_46,In_374);
or U196 (N_196,N_130,In_337);
and U197 (N_197,In_470,In_272);
nand U198 (N_198,N_84,N_175);
nor U199 (N_199,N_122,N_160);
nand U200 (N_200,In_34,N_50);
or U201 (N_201,In_412,N_171);
nor U202 (N_202,In_286,N_79);
nand U203 (N_203,In_214,N_28);
xor U204 (N_204,N_154,In_50);
nand U205 (N_205,In_33,N_151);
nor U206 (N_206,In_182,In_498);
and U207 (N_207,In_108,N_176);
nor U208 (N_208,N_148,In_231);
nand U209 (N_209,N_5,N_30);
and U210 (N_210,N_155,N_90);
and U211 (N_211,In_308,N_117);
or U212 (N_212,N_6,N_60);
nor U213 (N_213,In_468,In_131);
nor U214 (N_214,N_80,In_179);
nand U215 (N_215,In_164,N_106);
and U216 (N_216,In_353,In_306);
or U217 (N_217,In_207,In_460);
nand U218 (N_218,N_147,In_29);
and U219 (N_219,N_153,N_53);
nand U220 (N_220,N_73,In_287);
nand U221 (N_221,In_456,In_247);
or U222 (N_222,In_373,In_66);
nor U223 (N_223,N_25,In_466);
nor U224 (N_224,N_45,In_253);
and U225 (N_225,In_430,In_171);
or U226 (N_226,N_13,N_68);
xnor U227 (N_227,In_471,In_198);
or U228 (N_228,In_47,N_71);
nor U229 (N_229,N_86,In_201);
nor U230 (N_230,N_88,In_328);
or U231 (N_231,In_186,In_394);
and U232 (N_232,In_490,N_164);
or U233 (N_233,In_259,In_266);
and U234 (N_234,N_49,In_360);
nand U235 (N_235,In_52,In_448);
and U236 (N_236,N_55,In_367);
and U237 (N_237,N_124,In_63);
nor U238 (N_238,N_174,N_18);
nor U239 (N_239,N_17,N_74);
or U240 (N_240,In_134,In_477);
or U241 (N_241,N_162,N_220);
nor U242 (N_242,N_163,N_172);
xor U243 (N_243,In_165,N_180);
nor U244 (N_244,N_173,N_152);
nor U245 (N_245,N_166,N_100);
nand U246 (N_246,In_76,In_313);
xnor U247 (N_247,In_326,N_120);
or U248 (N_248,In_232,N_181);
and U249 (N_249,N_212,In_310);
nor U250 (N_250,N_199,N_121);
nor U251 (N_251,In_261,In_194);
nand U252 (N_252,N_47,In_159);
nand U253 (N_253,In_364,N_134);
nor U254 (N_254,In_475,In_380);
and U255 (N_255,In_155,N_137);
or U256 (N_256,In_435,In_297);
xor U257 (N_257,In_216,In_243);
nor U258 (N_258,In_296,N_101);
and U259 (N_259,In_368,In_74);
nor U260 (N_260,N_139,N_111);
nand U261 (N_261,In_342,N_123);
and U262 (N_262,In_69,In_189);
or U263 (N_263,N_158,N_203);
xor U264 (N_264,In_249,In_188);
and U265 (N_265,N_8,N_128);
and U266 (N_266,N_156,N_142);
or U267 (N_267,N_56,N_184);
and U268 (N_268,In_5,N_75);
nand U269 (N_269,In_288,N_215);
nand U270 (N_270,In_358,N_192);
nand U271 (N_271,In_439,In_95);
or U272 (N_272,N_165,N_188);
or U273 (N_273,In_476,N_22);
or U274 (N_274,N_61,In_452);
or U275 (N_275,N_170,N_223);
or U276 (N_276,In_92,N_205);
or U277 (N_277,In_270,N_189);
nand U278 (N_278,In_197,In_26);
or U279 (N_279,In_343,N_194);
or U280 (N_280,N_229,N_127);
and U281 (N_281,N_102,N_21);
nor U282 (N_282,In_255,N_233);
and U283 (N_283,N_169,N_235);
and U284 (N_284,N_230,N_231);
nand U285 (N_285,In_65,N_178);
nand U286 (N_286,N_211,In_277);
nand U287 (N_287,In_187,N_177);
nor U288 (N_288,N_91,In_486);
and U289 (N_289,N_143,N_204);
or U290 (N_290,In_3,In_294);
nand U291 (N_291,In_283,N_32);
nor U292 (N_292,N_195,N_227);
nor U293 (N_293,In_413,In_61);
nand U294 (N_294,In_469,N_214);
nor U295 (N_295,In_10,N_135);
nor U296 (N_296,N_236,In_135);
nand U297 (N_297,N_208,N_224);
nand U298 (N_298,N_217,N_222);
nor U299 (N_299,N_57,In_428);
nand U300 (N_300,In_124,In_167);
nor U301 (N_301,In_362,N_48);
nand U302 (N_302,In_80,N_105);
and U303 (N_303,N_271,N_89);
or U304 (N_304,In_304,In_193);
nand U305 (N_305,N_209,N_244);
nor U306 (N_306,In_141,N_168);
or U307 (N_307,N_213,N_256);
or U308 (N_308,N_182,N_284);
or U309 (N_309,N_258,N_70);
nand U310 (N_310,In_375,N_248);
or U311 (N_311,In_36,In_217);
and U312 (N_312,N_239,In_269);
nor U313 (N_313,In_396,N_296);
or U314 (N_314,In_68,N_249);
or U315 (N_315,N_275,N_290);
xnor U316 (N_316,N_291,In_361);
and U317 (N_317,N_285,In_299);
and U318 (N_318,N_264,In_12);
nand U319 (N_319,N_108,In_302);
or U320 (N_320,N_260,In_126);
nand U321 (N_321,In_479,N_234);
nand U322 (N_322,N_263,In_419);
nor U323 (N_323,N_140,In_100);
nand U324 (N_324,In_18,N_62);
or U325 (N_325,N_270,In_87);
nand U326 (N_326,N_150,N_255);
nand U327 (N_327,N_250,N_119);
nor U328 (N_328,N_23,N_136);
nand U329 (N_329,In_79,N_219);
nand U330 (N_330,In_410,In_228);
and U331 (N_331,N_85,N_293);
nor U332 (N_332,N_240,N_228);
nor U333 (N_333,In_51,N_294);
nor U334 (N_334,N_51,N_297);
nor U335 (N_335,N_226,N_78);
or U336 (N_336,N_201,N_276);
or U337 (N_337,N_67,In_389);
xnor U338 (N_338,N_274,In_464);
nor U339 (N_339,In_416,N_246);
nor U340 (N_340,N_267,N_196);
and U341 (N_341,In_403,N_149);
and U342 (N_342,N_159,In_25);
or U343 (N_343,N_247,N_131);
nor U344 (N_344,In_319,N_207);
nand U345 (N_345,N_31,In_497);
or U346 (N_346,N_254,N_286);
xnor U347 (N_347,N_125,N_252);
and U348 (N_348,N_253,N_281);
or U349 (N_349,N_266,N_232);
nor U350 (N_350,N_243,N_257);
nor U351 (N_351,N_241,N_280);
nand U352 (N_352,N_126,N_185);
nand U353 (N_353,In_265,N_197);
or U354 (N_354,N_265,N_269);
or U355 (N_355,In_315,In_220);
nand U356 (N_356,In_285,N_190);
and U357 (N_357,N_183,In_432);
or U358 (N_358,N_10,In_405);
and U359 (N_359,N_295,N_157);
nand U360 (N_360,N_306,N_341);
or U361 (N_361,N_318,N_262);
nor U362 (N_362,N_332,N_268);
nor U363 (N_363,N_309,N_329);
nor U364 (N_364,In_43,N_87);
and U365 (N_365,N_216,N_310);
or U366 (N_366,N_301,In_110);
or U367 (N_367,N_358,In_284);
or U368 (N_368,N_251,N_64);
and U369 (N_369,N_356,N_304);
nor U370 (N_370,N_289,N_359);
nor U371 (N_371,N_357,In_145);
and U372 (N_372,N_287,N_12);
nor U373 (N_373,In_0,N_333);
or U374 (N_374,In_388,N_334);
nor U375 (N_375,N_307,N_340);
or U376 (N_376,N_336,N_354);
nor U377 (N_377,In_347,N_300);
nand U378 (N_378,N_138,N_179);
or U379 (N_379,In_344,In_49);
and U380 (N_380,N_338,N_339);
and U381 (N_381,In_440,N_346);
nor U382 (N_382,N_344,N_351);
and U383 (N_383,N_242,In_127);
nand U384 (N_384,In_365,N_319);
or U385 (N_385,N_191,N_210);
nor U386 (N_386,N_349,N_311);
and U387 (N_387,N_331,In_240);
nand U388 (N_388,N_305,N_343);
nand U389 (N_389,N_321,In_57);
nor U390 (N_390,N_322,N_299);
nor U391 (N_391,N_328,N_308);
xnor U392 (N_392,In_227,In_239);
and U393 (N_393,N_193,N_107);
and U394 (N_394,N_94,N_261);
and U395 (N_395,N_272,N_279);
and U396 (N_396,N_326,In_386);
or U397 (N_397,In_357,N_292);
or U398 (N_398,N_187,N_303);
nor U399 (N_399,N_316,N_167);
nand U400 (N_400,N_348,N_206);
and U401 (N_401,N_202,N_259);
or U402 (N_402,N_129,N_317);
or U403 (N_403,In_129,N_320);
or U404 (N_404,N_225,N_282);
nand U405 (N_405,N_221,N_245);
or U406 (N_406,N_323,N_342);
and U407 (N_407,N_352,N_298);
nor U408 (N_408,In_191,In_163);
nand U409 (N_409,N_345,N_302);
nand U410 (N_410,N_198,N_325);
and U411 (N_411,In_236,In_370);
or U412 (N_412,N_283,N_312);
nor U413 (N_413,N_146,N_278);
or U414 (N_414,N_3,In_199);
nor U415 (N_415,N_238,N_353);
nor U416 (N_416,N_315,N_337);
and U417 (N_417,In_352,N_141);
and U418 (N_418,N_44,N_327);
and U419 (N_419,N_186,N_335);
nand U420 (N_420,N_414,N_402);
nor U421 (N_421,N_393,N_132);
nor U422 (N_422,N_368,N_394);
or U423 (N_423,N_365,N_389);
nor U424 (N_424,N_380,N_406);
nand U425 (N_425,N_399,N_237);
nor U426 (N_426,N_350,N_387);
and U427 (N_427,N_417,N_377);
or U428 (N_428,N_381,N_415);
or U429 (N_429,In_408,N_403);
and U430 (N_430,N_363,N_374);
nand U431 (N_431,N_371,N_386);
nand U432 (N_432,N_378,N_412);
and U433 (N_433,N_364,N_273);
or U434 (N_434,N_362,N_218);
or U435 (N_435,N_375,N_418);
nand U436 (N_436,N_411,N_416);
and U437 (N_437,N_395,N_409);
xnor U438 (N_438,N_383,N_324);
and U439 (N_439,N_288,N_382);
nor U440 (N_440,N_392,N_366);
or U441 (N_441,N_369,N_372);
nor U442 (N_442,In_282,N_388);
nand U443 (N_443,N_397,N_410);
or U444 (N_444,N_370,N_367);
nor U445 (N_445,N_35,N_407);
nand U446 (N_446,N_37,In_96);
nor U447 (N_447,N_401,N_82);
nor U448 (N_448,N_313,N_413);
nand U449 (N_449,N_355,N_314);
nand U450 (N_450,N_400,N_277);
and U451 (N_451,N_373,N_384);
nand U452 (N_452,N_360,N_347);
nor U453 (N_453,N_200,N_408);
or U454 (N_454,N_405,N_398);
nand U455 (N_455,N_361,N_385);
nor U456 (N_456,N_419,N_390);
or U457 (N_457,N_379,N_396);
or U458 (N_458,N_391,N_330);
nor U459 (N_459,N_376,N_404);
or U460 (N_460,N_365,N_415);
nand U461 (N_461,N_412,N_403);
xor U462 (N_462,N_82,N_389);
and U463 (N_463,N_388,N_365);
or U464 (N_464,N_385,N_408);
nor U465 (N_465,N_390,N_411);
and U466 (N_466,N_347,N_361);
and U467 (N_467,N_366,N_324);
or U468 (N_468,N_371,N_35);
or U469 (N_469,N_273,N_390);
nand U470 (N_470,N_411,N_413);
nor U471 (N_471,N_408,N_37);
nand U472 (N_472,N_391,N_35);
nand U473 (N_473,N_82,N_273);
nor U474 (N_474,N_384,N_200);
nand U475 (N_475,N_404,N_200);
and U476 (N_476,In_96,N_386);
nor U477 (N_477,N_400,N_35);
nand U478 (N_478,N_406,N_379);
nand U479 (N_479,N_393,N_414);
and U480 (N_480,N_429,N_426);
and U481 (N_481,N_428,N_441);
xor U482 (N_482,N_430,N_465);
and U483 (N_483,N_434,N_467);
and U484 (N_484,N_421,N_433);
and U485 (N_485,N_446,N_439);
nand U486 (N_486,N_438,N_425);
nand U487 (N_487,N_455,N_463);
and U488 (N_488,N_459,N_452);
and U489 (N_489,N_473,N_450);
nor U490 (N_490,N_431,N_474);
nand U491 (N_491,N_478,N_466);
nor U492 (N_492,N_443,N_432);
and U493 (N_493,N_424,N_462);
or U494 (N_494,N_427,N_472);
nand U495 (N_495,N_454,N_470);
or U496 (N_496,N_471,N_420);
nand U497 (N_497,N_449,N_460);
or U498 (N_498,N_475,N_423);
or U499 (N_499,N_447,N_440);
nand U500 (N_500,N_457,N_469);
nand U501 (N_501,N_453,N_422);
nand U502 (N_502,N_442,N_461);
nand U503 (N_503,N_451,N_437);
nand U504 (N_504,N_468,N_444);
and U505 (N_505,N_476,N_445);
nor U506 (N_506,N_458,N_477);
and U507 (N_507,N_435,N_448);
and U508 (N_508,N_464,N_436);
nor U509 (N_509,N_479,N_456);
and U510 (N_510,N_437,N_460);
and U511 (N_511,N_469,N_466);
nand U512 (N_512,N_449,N_452);
nor U513 (N_513,N_459,N_451);
or U514 (N_514,N_475,N_449);
and U515 (N_515,N_440,N_444);
nand U516 (N_516,N_429,N_448);
and U517 (N_517,N_435,N_468);
and U518 (N_518,N_429,N_463);
or U519 (N_519,N_449,N_463);
or U520 (N_520,N_459,N_470);
nand U521 (N_521,N_449,N_439);
nand U522 (N_522,N_473,N_471);
or U523 (N_523,N_465,N_437);
or U524 (N_524,N_452,N_467);
nand U525 (N_525,N_435,N_440);
and U526 (N_526,N_436,N_432);
xor U527 (N_527,N_473,N_474);
and U528 (N_528,N_462,N_459);
and U529 (N_529,N_475,N_448);
and U530 (N_530,N_460,N_427);
nor U531 (N_531,N_450,N_448);
or U532 (N_532,N_467,N_420);
or U533 (N_533,N_446,N_461);
or U534 (N_534,N_437,N_426);
and U535 (N_535,N_436,N_460);
xor U536 (N_536,N_474,N_444);
nor U537 (N_537,N_427,N_428);
nand U538 (N_538,N_438,N_458);
nor U539 (N_539,N_459,N_475);
nor U540 (N_540,N_510,N_482);
and U541 (N_541,N_514,N_502);
nor U542 (N_542,N_492,N_524);
or U543 (N_543,N_501,N_516);
nand U544 (N_544,N_533,N_512);
and U545 (N_545,N_522,N_538);
nor U546 (N_546,N_519,N_525);
nand U547 (N_547,N_534,N_489);
nor U548 (N_548,N_520,N_517);
nand U549 (N_549,N_513,N_523);
nand U550 (N_550,N_506,N_503);
or U551 (N_551,N_521,N_488);
or U552 (N_552,N_498,N_485);
nor U553 (N_553,N_481,N_531);
nor U554 (N_554,N_515,N_486);
or U555 (N_555,N_497,N_536);
nand U556 (N_556,N_537,N_480);
and U557 (N_557,N_490,N_532);
and U558 (N_558,N_518,N_528);
and U559 (N_559,N_527,N_491);
xor U560 (N_560,N_499,N_535);
nand U561 (N_561,N_511,N_487);
nand U562 (N_562,N_494,N_500);
nor U563 (N_563,N_504,N_508);
and U564 (N_564,N_483,N_526);
nand U565 (N_565,N_530,N_495);
and U566 (N_566,N_539,N_509);
or U567 (N_567,N_507,N_529);
nor U568 (N_568,N_484,N_496);
nor U569 (N_569,N_493,N_505);
nor U570 (N_570,N_504,N_512);
or U571 (N_571,N_507,N_516);
nand U572 (N_572,N_526,N_494);
nand U573 (N_573,N_508,N_505);
or U574 (N_574,N_481,N_537);
nand U575 (N_575,N_510,N_530);
or U576 (N_576,N_503,N_489);
nor U577 (N_577,N_539,N_530);
and U578 (N_578,N_511,N_523);
nor U579 (N_579,N_511,N_519);
nor U580 (N_580,N_523,N_488);
and U581 (N_581,N_529,N_503);
and U582 (N_582,N_481,N_530);
nor U583 (N_583,N_481,N_492);
and U584 (N_584,N_532,N_487);
or U585 (N_585,N_483,N_493);
nand U586 (N_586,N_539,N_493);
or U587 (N_587,N_525,N_520);
nor U588 (N_588,N_530,N_491);
or U589 (N_589,N_508,N_531);
and U590 (N_590,N_517,N_532);
nor U591 (N_591,N_488,N_525);
and U592 (N_592,N_510,N_522);
nand U593 (N_593,N_535,N_517);
nor U594 (N_594,N_505,N_511);
or U595 (N_595,N_500,N_483);
or U596 (N_596,N_485,N_496);
or U597 (N_597,N_480,N_499);
xor U598 (N_598,N_525,N_517);
nor U599 (N_599,N_528,N_525);
nor U600 (N_600,N_580,N_587);
nand U601 (N_601,N_588,N_558);
nor U602 (N_602,N_555,N_573);
and U603 (N_603,N_597,N_563);
and U604 (N_604,N_557,N_541);
and U605 (N_605,N_585,N_546);
and U606 (N_606,N_540,N_543);
nand U607 (N_607,N_582,N_599);
and U608 (N_608,N_544,N_575);
or U609 (N_609,N_559,N_561);
or U610 (N_610,N_545,N_566);
or U611 (N_611,N_598,N_581);
nand U612 (N_612,N_562,N_567);
and U613 (N_613,N_590,N_589);
nor U614 (N_614,N_548,N_552);
nand U615 (N_615,N_560,N_551);
nand U616 (N_616,N_593,N_568);
nand U617 (N_617,N_595,N_596);
or U618 (N_618,N_594,N_564);
nand U619 (N_619,N_550,N_578);
nand U620 (N_620,N_572,N_574);
nand U621 (N_621,N_592,N_553);
nand U622 (N_622,N_579,N_569);
and U623 (N_623,N_577,N_549);
and U624 (N_624,N_547,N_570);
nand U625 (N_625,N_542,N_571);
xnor U626 (N_626,N_576,N_583);
nor U627 (N_627,N_554,N_586);
nor U628 (N_628,N_556,N_565);
or U629 (N_629,N_591,N_584);
and U630 (N_630,N_589,N_578);
and U631 (N_631,N_589,N_574);
and U632 (N_632,N_570,N_557);
nor U633 (N_633,N_585,N_573);
nor U634 (N_634,N_593,N_596);
nand U635 (N_635,N_546,N_555);
nand U636 (N_636,N_569,N_553);
nand U637 (N_637,N_594,N_595);
or U638 (N_638,N_582,N_566);
nor U639 (N_639,N_595,N_566);
and U640 (N_640,N_590,N_562);
nor U641 (N_641,N_563,N_592);
xnor U642 (N_642,N_563,N_572);
nand U643 (N_643,N_559,N_585);
nor U644 (N_644,N_556,N_566);
nand U645 (N_645,N_549,N_547);
nor U646 (N_646,N_599,N_591);
and U647 (N_647,N_591,N_594);
and U648 (N_648,N_551,N_559);
or U649 (N_649,N_568,N_557);
nor U650 (N_650,N_568,N_540);
and U651 (N_651,N_575,N_592);
or U652 (N_652,N_566,N_542);
nand U653 (N_653,N_550,N_543);
and U654 (N_654,N_552,N_568);
nor U655 (N_655,N_590,N_594);
or U656 (N_656,N_577,N_556);
and U657 (N_657,N_544,N_595);
nor U658 (N_658,N_545,N_587);
and U659 (N_659,N_568,N_571);
or U660 (N_660,N_621,N_602);
or U661 (N_661,N_608,N_601);
xnor U662 (N_662,N_625,N_606);
xnor U663 (N_663,N_639,N_644);
and U664 (N_664,N_642,N_658);
xnor U665 (N_665,N_646,N_652);
nor U666 (N_666,N_649,N_628);
and U667 (N_667,N_631,N_650);
and U668 (N_668,N_630,N_635);
nand U669 (N_669,N_615,N_604);
or U670 (N_670,N_612,N_610);
and U671 (N_671,N_647,N_623);
and U672 (N_672,N_651,N_654);
and U673 (N_673,N_643,N_619);
or U674 (N_674,N_636,N_622);
or U675 (N_675,N_616,N_618);
nand U676 (N_676,N_629,N_603);
nand U677 (N_677,N_638,N_645);
nor U678 (N_678,N_659,N_600);
or U679 (N_679,N_627,N_637);
nor U680 (N_680,N_633,N_634);
nor U681 (N_681,N_611,N_620);
nor U682 (N_682,N_648,N_640);
and U683 (N_683,N_613,N_614);
nor U684 (N_684,N_632,N_641);
xnor U685 (N_685,N_657,N_605);
or U686 (N_686,N_653,N_607);
nor U687 (N_687,N_656,N_617);
nand U688 (N_688,N_609,N_624);
and U689 (N_689,N_626,N_655);
nor U690 (N_690,N_625,N_643);
nor U691 (N_691,N_606,N_622);
nor U692 (N_692,N_608,N_635);
nor U693 (N_693,N_635,N_637);
nor U694 (N_694,N_640,N_618);
or U695 (N_695,N_600,N_612);
and U696 (N_696,N_657,N_648);
xnor U697 (N_697,N_649,N_611);
or U698 (N_698,N_647,N_610);
nand U699 (N_699,N_613,N_649);
nor U700 (N_700,N_652,N_604);
nor U701 (N_701,N_654,N_647);
and U702 (N_702,N_654,N_606);
xor U703 (N_703,N_643,N_637);
and U704 (N_704,N_610,N_613);
and U705 (N_705,N_628,N_624);
and U706 (N_706,N_625,N_631);
or U707 (N_707,N_607,N_625);
xnor U708 (N_708,N_656,N_622);
nor U709 (N_709,N_649,N_641);
and U710 (N_710,N_600,N_626);
and U711 (N_711,N_604,N_609);
nor U712 (N_712,N_614,N_611);
and U713 (N_713,N_617,N_600);
nor U714 (N_714,N_643,N_636);
nor U715 (N_715,N_604,N_626);
nand U716 (N_716,N_604,N_605);
nand U717 (N_717,N_617,N_657);
nand U718 (N_718,N_651,N_604);
nand U719 (N_719,N_634,N_639);
nand U720 (N_720,N_679,N_680);
nand U721 (N_721,N_697,N_666);
nand U722 (N_722,N_714,N_671);
and U723 (N_723,N_688,N_672);
nand U724 (N_724,N_673,N_707);
or U725 (N_725,N_681,N_670);
nand U726 (N_726,N_718,N_694);
nor U727 (N_727,N_665,N_660);
and U728 (N_728,N_683,N_690);
nor U729 (N_729,N_662,N_715);
and U730 (N_730,N_696,N_709);
and U731 (N_731,N_684,N_675);
or U732 (N_732,N_695,N_668);
or U733 (N_733,N_692,N_678);
or U734 (N_734,N_699,N_708);
nor U735 (N_735,N_677,N_703);
nor U736 (N_736,N_711,N_682);
or U737 (N_737,N_663,N_704);
nor U738 (N_738,N_719,N_710);
xnor U739 (N_739,N_686,N_693);
nor U740 (N_740,N_705,N_664);
nor U741 (N_741,N_706,N_691);
and U742 (N_742,N_713,N_716);
and U743 (N_743,N_689,N_698);
nor U744 (N_744,N_717,N_701);
and U745 (N_745,N_667,N_687);
and U746 (N_746,N_674,N_712);
and U747 (N_747,N_676,N_700);
nand U748 (N_748,N_669,N_685);
xnor U749 (N_749,N_661,N_702);
and U750 (N_750,N_667,N_675);
nand U751 (N_751,N_662,N_690);
nor U752 (N_752,N_685,N_708);
or U753 (N_753,N_690,N_672);
or U754 (N_754,N_711,N_718);
nand U755 (N_755,N_714,N_672);
nand U756 (N_756,N_698,N_678);
nand U757 (N_757,N_708,N_677);
nand U758 (N_758,N_703,N_687);
nand U759 (N_759,N_666,N_699);
nand U760 (N_760,N_704,N_703);
xor U761 (N_761,N_707,N_665);
nand U762 (N_762,N_661,N_685);
or U763 (N_763,N_708,N_707);
nor U764 (N_764,N_678,N_675);
and U765 (N_765,N_701,N_676);
xor U766 (N_766,N_705,N_710);
and U767 (N_767,N_677,N_717);
nand U768 (N_768,N_688,N_698);
nand U769 (N_769,N_678,N_668);
nand U770 (N_770,N_671,N_663);
or U771 (N_771,N_682,N_661);
nand U772 (N_772,N_716,N_698);
nor U773 (N_773,N_695,N_690);
nor U774 (N_774,N_682,N_687);
or U775 (N_775,N_677,N_676);
xnor U776 (N_776,N_716,N_679);
and U777 (N_777,N_681,N_704);
nor U778 (N_778,N_692,N_718);
or U779 (N_779,N_664,N_706);
or U780 (N_780,N_769,N_743);
xor U781 (N_781,N_756,N_752);
nand U782 (N_782,N_744,N_727);
nor U783 (N_783,N_724,N_768);
nand U784 (N_784,N_770,N_757);
nand U785 (N_785,N_758,N_746);
or U786 (N_786,N_736,N_740);
xor U787 (N_787,N_738,N_729);
nor U788 (N_788,N_763,N_749);
nor U789 (N_789,N_778,N_753);
nor U790 (N_790,N_750,N_774);
nand U791 (N_791,N_734,N_742);
nor U792 (N_792,N_720,N_755);
or U793 (N_793,N_751,N_762);
or U794 (N_794,N_721,N_772);
nand U795 (N_795,N_765,N_733);
or U796 (N_796,N_730,N_726);
and U797 (N_797,N_732,N_779);
and U798 (N_798,N_767,N_722);
or U799 (N_799,N_741,N_748);
xnor U800 (N_800,N_728,N_723);
and U801 (N_801,N_754,N_775);
nand U802 (N_802,N_760,N_735);
and U803 (N_803,N_745,N_739);
nor U804 (N_804,N_725,N_773);
or U805 (N_805,N_737,N_759);
and U806 (N_806,N_747,N_771);
nor U807 (N_807,N_776,N_764);
nand U808 (N_808,N_766,N_731);
xnor U809 (N_809,N_761,N_777);
and U810 (N_810,N_766,N_758);
or U811 (N_811,N_733,N_731);
nor U812 (N_812,N_725,N_760);
nor U813 (N_813,N_729,N_741);
or U814 (N_814,N_728,N_760);
and U815 (N_815,N_728,N_742);
and U816 (N_816,N_771,N_749);
and U817 (N_817,N_745,N_772);
and U818 (N_818,N_766,N_762);
or U819 (N_819,N_770,N_742);
nor U820 (N_820,N_721,N_737);
nor U821 (N_821,N_749,N_742);
nor U822 (N_822,N_734,N_761);
or U823 (N_823,N_741,N_769);
and U824 (N_824,N_725,N_738);
nor U825 (N_825,N_775,N_779);
nor U826 (N_826,N_726,N_747);
nand U827 (N_827,N_756,N_753);
and U828 (N_828,N_753,N_738);
or U829 (N_829,N_754,N_739);
or U830 (N_830,N_736,N_778);
and U831 (N_831,N_733,N_750);
and U832 (N_832,N_749,N_730);
nor U833 (N_833,N_735,N_767);
or U834 (N_834,N_720,N_739);
nor U835 (N_835,N_759,N_760);
or U836 (N_836,N_761,N_751);
or U837 (N_837,N_778,N_767);
nand U838 (N_838,N_741,N_751);
nand U839 (N_839,N_726,N_728);
nand U840 (N_840,N_783,N_832);
nand U841 (N_841,N_797,N_792);
nand U842 (N_842,N_799,N_814);
nor U843 (N_843,N_817,N_823);
and U844 (N_844,N_806,N_786);
nand U845 (N_845,N_834,N_830);
and U846 (N_846,N_801,N_811);
nor U847 (N_847,N_795,N_827);
nor U848 (N_848,N_816,N_829);
and U849 (N_849,N_788,N_784);
nand U850 (N_850,N_805,N_826);
and U851 (N_851,N_813,N_822);
nand U852 (N_852,N_803,N_836);
nand U853 (N_853,N_807,N_782);
and U854 (N_854,N_820,N_835);
or U855 (N_855,N_787,N_791);
or U856 (N_856,N_812,N_810);
nand U857 (N_857,N_838,N_796);
nand U858 (N_858,N_825,N_780);
nor U859 (N_859,N_831,N_819);
nor U860 (N_860,N_818,N_833);
nand U861 (N_861,N_809,N_821);
nor U862 (N_862,N_781,N_839);
nand U863 (N_863,N_824,N_790);
and U864 (N_864,N_802,N_794);
nor U865 (N_865,N_800,N_828);
nand U866 (N_866,N_808,N_789);
and U867 (N_867,N_785,N_815);
and U868 (N_868,N_804,N_837);
and U869 (N_869,N_798,N_793);
nand U870 (N_870,N_793,N_805);
and U871 (N_871,N_833,N_839);
nor U872 (N_872,N_813,N_797);
nand U873 (N_873,N_824,N_795);
or U874 (N_874,N_809,N_839);
nand U875 (N_875,N_794,N_816);
nand U876 (N_876,N_823,N_818);
nand U877 (N_877,N_785,N_806);
nor U878 (N_878,N_799,N_816);
or U879 (N_879,N_799,N_802);
and U880 (N_880,N_809,N_820);
nor U881 (N_881,N_798,N_831);
or U882 (N_882,N_822,N_805);
nor U883 (N_883,N_828,N_802);
or U884 (N_884,N_816,N_795);
nand U885 (N_885,N_812,N_833);
or U886 (N_886,N_797,N_833);
or U887 (N_887,N_794,N_786);
nand U888 (N_888,N_809,N_819);
nand U889 (N_889,N_795,N_784);
nand U890 (N_890,N_828,N_830);
nor U891 (N_891,N_821,N_784);
nand U892 (N_892,N_787,N_824);
and U893 (N_893,N_839,N_794);
or U894 (N_894,N_819,N_838);
nand U895 (N_895,N_815,N_806);
nor U896 (N_896,N_821,N_833);
nor U897 (N_897,N_792,N_818);
xor U898 (N_898,N_809,N_828);
nand U899 (N_899,N_803,N_829);
nand U900 (N_900,N_872,N_852);
or U901 (N_901,N_848,N_873);
nor U902 (N_902,N_875,N_841);
nand U903 (N_903,N_879,N_874);
and U904 (N_904,N_858,N_888);
or U905 (N_905,N_886,N_876);
nor U906 (N_906,N_894,N_869);
and U907 (N_907,N_882,N_860);
or U908 (N_908,N_880,N_863);
nand U909 (N_909,N_878,N_857);
or U910 (N_910,N_889,N_847);
nor U911 (N_911,N_866,N_849);
or U912 (N_912,N_898,N_868);
and U913 (N_913,N_897,N_853);
and U914 (N_914,N_883,N_864);
and U915 (N_915,N_884,N_843);
nor U916 (N_916,N_896,N_893);
and U917 (N_917,N_877,N_851);
or U918 (N_918,N_870,N_850);
and U919 (N_919,N_891,N_861);
or U920 (N_920,N_842,N_867);
nand U921 (N_921,N_890,N_856);
nand U922 (N_922,N_859,N_899);
or U923 (N_923,N_885,N_855);
nor U924 (N_924,N_854,N_895);
or U925 (N_925,N_845,N_881);
xnor U926 (N_926,N_887,N_844);
and U927 (N_927,N_865,N_892);
nand U928 (N_928,N_862,N_871);
xnor U929 (N_929,N_840,N_846);
nor U930 (N_930,N_891,N_890);
and U931 (N_931,N_896,N_867);
or U932 (N_932,N_865,N_863);
and U933 (N_933,N_890,N_877);
or U934 (N_934,N_897,N_883);
nor U935 (N_935,N_874,N_847);
or U936 (N_936,N_843,N_849);
and U937 (N_937,N_854,N_859);
and U938 (N_938,N_844,N_877);
nand U939 (N_939,N_862,N_844);
nor U940 (N_940,N_845,N_878);
or U941 (N_941,N_852,N_861);
nor U942 (N_942,N_873,N_899);
and U943 (N_943,N_840,N_889);
and U944 (N_944,N_876,N_878);
and U945 (N_945,N_892,N_884);
or U946 (N_946,N_858,N_881);
or U947 (N_947,N_863,N_854);
and U948 (N_948,N_883,N_850);
nand U949 (N_949,N_857,N_863);
and U950 (N_950,N_873,N_867);
and U951 (N_951,N_873,N_857);
nand U952 (N_952,N_845,N_849);
nor U953 (N_953,N_852,N_844);
nand U954 (N_954,N_882,N_867);
or U955 (N_955,N_868,N_846);
and U956 (N_956,N_850,N_876);
xor U957 (N_957,N_869,N_866);
nand U958 (N_958,N_857,N_860);
and U959 (N_959,N_898,N_855);
nand U960 (N_960,N_905,N_903);
nor U961 (N_961,N_929,N_914);
and U962 (N_962,N_944,N_939);
or U963 (N_963,N_911,N_928);
and U964 (N_964,N_935,N_910);
or U965 (N_965,N_933,N_925);
nand U966 (N_966,N_924,N_920);
nor U967 (N_967,N_936,N_950);
nor U968 (N_968,N_908,N_947);
nor U969 (N_969,N_918,N_948);
or U970 (N_970,N_930,N_907);
or U971 (N_971,N_912,N_915);
xnor U972 (N_972,N_904,N_949);
and U973 (N_973,N_931,N_957);
and U974 (N_974,N_916,N_959);
or U975 (N_975,N_937,N_906);
nor U976 (N_976,N_951,N_923);
nand U977 (N_977,N_954,N_900);
and U978 (N_978,N_926,N_934);
nor U979 (N_979,N_901,N_919);
xor U980 (N_980,N_938,N_958);
nand U981 (N_981,N_955,N_922);
nand U982 (N_982,N_913,N_956);
or U983 (N_983,N_941,N_909);
and U984 (N_984,N_940,N_945);
or U985 (N_985,N_953,N_927);
nor U986 (N_986,N_917,N_902);
or U987 (N_987,N_952,N_932);
or U988 (N_988,N_946,N_942);
nor U989 (N_989,N_943,N_921);
or U990 (N_990,N_902,N_943);
or U991 (N_991,N_912,N_940);
nand U992 (N_992,N_923,N_952);
and U993 (N_993,N_900,N_946);
or U994 (N_994,N_923,N_959);
or U995 (N_995,N_902,N_923);
and U996 (N_996,N_953,N_908);
and U997 (N_997,N_950,N_949);
nand U998 (N_998,N_912,N_904);
and U999 (N_999,N_946,N_918);
and U1000 (N_1000,N_924,N_945);
and U1001 (N_1001,N_945,N_902);
nor U1002 (N_1002,N_949,N_942);
or U1003 (N_1003,N_945,N_925);
or U1004 (N_1004,N_949,N_955);
nand U1005 (N_1005,N_936,N_930);
nand U1006 (N_1006,N_924,N_946);
or U1007 (N_1007,N_918,N_916);
or U1008 (N_1008,N_918,N_915);
or U1009 (N_1009,N_906,N_942);
or U1010 (N_1010,N_910,N_938);
or U1011 (N_1011,N_900,N_937);
or U1012 (N_1012,N_919,N_957);
and U1013 (N_1013,N_919,N_940);
or U1014 (N_1014,N_934,N_920);
nand U1015 (N_1015,N_901,N_937);
nor U1016 (N_1016,N_957,N_922);
or U1017 (N_1017,N_928,N_923);
or U1018 (N_1018,N_957,N_926);
or U1019 (N_1019,N_953,N_943);
nand U1020 (N_1020,N_981,N_1009);
nand U1021 (N_1021,N_994,N_1012);
nor U1022 (N_1022,N_980,N_965);
nand U1023 (N_1023,N_1001,N_999);
or U1024 (N_1024,N_986,N_982);
nor U1025 (N_1025,N_990,N_1013);
and U1026 (N_1026,N_985,N_991);
nor U1027 (N_1027,N_993,N_977);
and U1028 (N_1028,N_997,N_984);
nand U1029 (N_1029,N_1019,N_960);
or U1030 (N_1030,N_988,N_1002);
and U1031 (N_1031,N_1008,N_972);
nand U1032 (N_1032,N_1005,N_976);
nor U1033 (N_1033,N_966,N_969);
nand U1034 (N_1034,N_989,N_1000);
or U1035 (N_1035,N_1010,N_961);
nand U1036 (N_1036,N_963,N_978);
and U1037 (N_1037,N_987,N_995);
or U1038 (N_1038,N_992,N_983);
nor U1039 (N_1039,N_962,N_1014);
or U1040 (N_1040,N_964,N_1018);
nor U1041 (N_1041,N_1007,N_968);
nand U1042 (N_1042,N_975,N_1003);
nand U1043 (N_1043,N_1017,N_1011);
or U1044 (N_1044,N_1004,N_971);
or U1045 (N_1045,N_1006,N_973);
nand U1046 (N_1046,N_998,N_974);
nand U1047 (N_1047,N_979,N_1015);
or U1048 (N_1048,N_970,N_967);
and U1049 (N_1049,N_1016,N_996);
or U1050 (N_1050,N_966,N_988);
nor U1051 (N_1051,N_980,N_968);
nor U1052 (N_1052,N_965,N_1001);
or U1053 (N_1053,N_962,N_1009);
and U1054 (N_1054,N_1016,N_1000);
nor U1055 (N_1055,N_976,N_979);
nor U1056 (N_1056,N_962,N_986);
nor U1057 (N_1057,N_965,N_1003);
or U1058 (N_1058,N_969,N_1006);
nand U1059 (N_1059,N_994,N_973);
nand U1060 (N_1060,N_993,N_983);
or U1061 (N_1061,N_976,N_996);
nand U1062 (N_1062,N_1000,N_1009);
nand U1063 (N_1063,N_989,N_998);
nor U1064 (N_1064,N_1005,N_974);
or U1065 (N_1065,N_1004,N_1011);
nor U1066 (N_1066,N_980,N_1013);
or U1067 (N_1067,N_1019,N_1012);
or U1068 (N_1068,N_1011,N_967);
or U1069 (N_1069,N_995,N_971);
nand U1070 (N_1070,N_978,N_977);
or U1071 (N_1071,N_960,N_966);
or U1072 (N_1072,N_1010,N_1012);
nor U1073 (N_1073,N_970,N_989);
nor U1074 (N_1074,N_996,N_1003);
and U1075 (N_1075,N_969,N_964);
or U1076 (N_1076,N_997,N_1007);
nor U1077 (N_1077,N_968,N_1003);
or U1078 (N_1078,N_972,N_990);
nor U1079 (N_1079,N_963,N_970);
and U1080 (N_1080,N_1077,N_1046);
nor U1081 (N_1081,N_1065,N_1020);
xor U1082 (N_1082,N_1068,N_1052);
nor U1083 (N_1083,N_1022,N_1072);
nand U1084 (N_1084,N_1028,N_1054);
and U1085 (N_1085,N_1033,N_1056);
nor U1086 (N_1086,N_1053,N_1074);
and U1087 (N_1087,N_1025,N_1048);
or U1088 (N_1088,N_1038,N_1039);
xor U1089 (N_1089,N_1061,N_1023);
nor U1090 (N_1090,N_1035,N_1030);
and U1091 (N_1091,N_1079,N_1041);
nand U1092 (N_1092,N_1026,N_1027);
nor U1093 (N_1093,N_1059,N_1051);
and U1094 (N_1094,N_1024,N_1067);
xnor U1095 (N_1095,N_1032,N_1078);
nand U1096 (N_1096,N_1073,N_1036);
xnor U1097 (N_1097,N_1045,N_1040);
nor U1098 (N_1098,N_1063,N_1031);
or U1099 (N_1099,N_1049,N_1057);
and U1100 (N_1100,N_1037,N_1034);
and U1101 (N_1101,N_1043,N_1044);
and U1102 (N_1102,N_1060,N_1070);
nand U1103 (N_1103,N_1066,N_1055);
and U1104 (N_1104,N_1076,N_1064);
or U1105 (N_1105,N_1058,N_1021);
and U1106 (N_1106,N_1069,N_1075);
or U1107 (N_1107,N_1042,N_1050);
and U1108 (N_1108,N_1029,N_1047);
nand U1109 (N_1109,N_1062,N_1071);
nor U1110 (N_1110,N_1054,N_1069);
or U1111 (N_1111,N_1069,N_1021);
or U1112 (N_1112,N_1063,N_1076);
and U1113 (N_1113,N_1044,N_1067);
or U1114 (N_1114,N_1062,N_1024);
nor U1115 (N_1115,N_1047,N_1041);
or U1116 (N_1116,N_1061,N_1027);
or U1117 (N_1117,N_1064,N_1028);
nand U1118 (N_1118,N_1059,N_1061);
and U1119 (N_1119,N_1034,N_1046);
or U1120 (N_1120,N_1035,N_1074);
nor U1121 (N_1121,N_1030,N_1071);
or U1122 (N_1122,N_1022,N_1038);
nor U1123 (N_1123,N_1024,N_1074);
or U1124 (N_1124,N_1052,N_1043);
nand U1125 (N_1125,N_1069,N_1079);
and U1126 (N_1126,N_1061,N_1071);
or U1127 (N_1127,N_1062,N_1026);
or U1128 (N_1128,N_1026,N_1073);
nand U1129 (N_1129,N_1033,N_1075);
or U1130 (N_1130,N_1069,N_1033);
or U1131 (N_1131,N_1057,N_1079);
nor U1132 (N_1132,N_1033,N_1040);
nor U1133 (N_1133,N_1078,N_1067);
nor U1134 (N_1134,N_1066,N_1078);
and U1135 (N_1135,N_1020,N_1076);
nand U1136 (N_1136,N_1078,N_1033);
xnor U1137 (N_1137,N_1023,N_1066);
nand U1138 (N_1138,N_1063,N_1020);
or U1139 (N_1139,N_1076,N_1046);
nand U1140 (N_1140,N_1128,N_1096);
and U1141 (N_1141,N_1109,N_1114);
nor U1142 (N_1142,N_1101,N_1130);
nor U1143 (N_1143,N_1117,N_1083);
or U1144 (N_1144,N_1087,N_1107);
or U1145 (N_1145,N_1106,N_1137);
nor U1146 (N_1146,N_1103,N_1102);
nand U1147 (N_1147,N_1092,N_1124);
nand U1148 (N_1148,N_1131,N_1081);
nor U1149 (N_1149,N_1120,N_1085);
or U1150 (N_1150,N_1119,N_1091);
nand U1151 (N_1151,N_1121,N_1104);
nand U1152 (N_1152,N_1111,N_1113);
and U1153 (N_1153,N_1116,N_1097);
or U1154 (N_1154,N_1088,N_1133);
and U1155 (N_1155,N_1129,N_1086);
or U1156 (N_1156,N_1108,N_1084);
or U1157 (N_1157,N_1110,N_1093);
nand U1158 (N_1158,N_1115,N_1098);
nor U1159 (N_1159,N_1094,N_1100);
and U1160 (N_1160,N_1122,N_1112);
and U1161 (N_1161,N_1080,N_1132);
xnor U1162 (N_1162,N_1099,N_1089);
or U1163 (N_1163,N_1127,N_1090);
nor U1164 (N_1164,N_1082,N_1105);
or U1165 (N_1165,N_1126,N_1138);
nand U1166 (N_1166,N_1136,N_1095);
xnor U1167 (N_1167,N_1134,N_1118);
and U1168 (N_1168,N_1125,N_1135);
nand U1169 (N_1169,N_1139,N_1123);
or U1170 (N_1170,N_1114,N_1093);
nor U1171 (N_1171,N_1081,N_1121);
nand U1172 (N_1172,N_1099,N_1110);
xor U1173 (N_1173,N_1121,N_1084);
and U1174 (N_1174,N_1107,N_1099);
nand U1175 (N_1175,N_1089,N_1081);
or U1176 (N_1176,N_1101,N_1134);
or U1177 (N_1177,N_1107,N_1115);
and U1178 (N_1178,N_1111,N_1105);
or U1179 (N_1179,N_1086,N_1106);
nand U1180 (N_1180,N_1138,N_1120);
nand U1181 (N_1181,N_1124,N_1080);
nand U1182 (N_1182,N_1117,N_1098);
nand U1183 (N_1183,N_1136,N_1121);
nor U1184 (N_1184,N_1124,N_1097);
nand U1185 (N_1185,N_1116,N_1114);
and U1186 (N_1186,N_1102,N_1082);
nand U1187 (N_1187,N_1103,N_1105);
nand U1188 (N_1188,N_1090,N_1138);
and U1189 (N_1189,N_1127,N_1125);
or U1190 (N_1190,N_1119,N_1123);
and U1191 (N_1191,N_1137,N_1096);
nand U1192 (N_1192,N_1086,N_1108);
or U1193 (N_1193,N_1088,N_1134);
and U1194 (N_1194,N_1133,N_1103);
nor U1195 (N_1195,N_1102,N_1134);
or U1196 (N_1196,N_1110,N_1088);
and U1197 (N_1197,N_1109,N_1121);
nor U1198 (N_1198,N_1085,N_1122);
and U1199 (N_1199,N_1125,N_1086);
xnor U1200 (N_1200,N_1172,N_1148);
nand U1201 (N_1201,N_1198,N_1187);
nor U1202 (N_1202,N_1159,N_1168);
or U1203 (N_1203,N_1170,N_1150);
and U1204 (N_1204,N_1186,N_1183);
or U1205 (N_1205,N_1179,N_1140);
or U1206 (N_1206,N_1195,N_1165);
nand U1207 (N_1207,N_1151,N_1152);
nand U1208 (N_1208,N_1142,N_1192);
nand U1209 (N_1209,N_1155,N_1191);
nor U1210 (N_1210,N_1177,N_1145);
nand U1211 (N_1211,N_1161,N_1182);
xnor U1212 (N_1212,N_1189,N_1181);
nand U1213 (N_1213,N_1146,N_1174);
or U1214 (N_1214,N_1164,N_1178);
and U1215 (N_1215,N_1169,N_1163);
nand U1216 (N_1216,N_1194,N_1156);
and U1217 (N_1217,N_1173,N_1193);
and U1218 (N_1218,N_1171,N_1176);
or U1219 (N_1219,N_1153,N_1141);
nand U1220 (N_1220,N_1154,N_1166);
xnor U1221 (N_1221,N_1147,N_1157);
nand U1222 (N_1222,N_1180,N_1199);
and U1223 (N_1223,N_1144,N_1196);
nor U1224 (N_1224,N_1162,N_1158);
nor U1225 (N_1225,N_1167,N_1197);
nor U1226 (N_1226,N_1149,N_1185);
nor U1227 (N_1227,N_1175,N_1184);
and U1228 (N_1228,N_1143,N_1188);
or U1229 (N_1229,N_1190,N_1160);
and U1230 (N_1230,N_1185,N_1159);
nand U1231 (N_1231,N_1148,N_1162);
nand U1232 (N_1232,N_1189,N_1141);
nand U1233 (N_1233,N_1174,N_1198);
and U1234 (N_1234,N_1153,N_1161);
nand U1235 (N_1235,N_1184,N_1170);
and U1236 (N_1236,N_1151,N_1167);
and U1237 (N_1237,N_1166,N_1142);
or U1238 (N_1238,N_1150,N_1185);
nor U1239 (N_1239,N_1194,N_1182);
or U1240 (N_1240,N_1183,N_1198);
nand U1241 (N_1241,N_1197,N_1159);
or U1242 (N_1242,N_1178,N_1190);
nand U1243 (N_1243,N_1180,N_1183);
and U1244 (N_1244,N_1140,N_1176);
nand U1245 (N_1245,N_1169,N_1159);
xor U1246 (N_1246,N_1143,N_1182);
nor U1247 (N_1247,N_1186,N_1163);
or U1248 (N_1248,N_1151,N_1169);
or U1249 (N_1249,N_1176,N_1159);
nand U1250 (N_1250,N_1170,N_1185);
xor U1251 (N_1251,N_1188,N_1149);
or U1252 (N_1252,N_1170,N_1141);
nand U1253 (N_1253,N_1174,N_1183);
nand U1254 (N_1254,N_1141,N_1199);
and U1255 (N_1255,N_1168,N_1173);
and U1256 (N_1256,N_1181,N_1187);
and U1257 (N_1257,N_1142,N_1178);
and U1258 (N_1258,N_1189,N_1169);
or U1259 (N_1259,N_1176,N_1153);
or U1260 (N_1260,N_1230,N_1201);
nor U1261 (N_1261,N_1258,N_1212);
and U1262 (N_1262,N_1203,N_1207);
nor U1263 (N_1263,N_1236,N_1259);
nand U1264 (N_1264,N_1217,N_1220);
nor U1265 (N_1265,N_1243,N_1246);
nor U1266 (N_1266,N_1218,N_1224);
nand U1267 (N_1267,N_1245,N_1238);
or U1268 (N_1268,N_1233,N_1209);
nor U1269 (N_1269,N_1222,N_1249);
or U1270 (N_1270,N_1204,N_1241);
nor U1271 (N_1271,N_1208,N_1255);
nor U1272 (N_1272,N_1239,N_1205);
and U1273 (N_1273,N_1248,N_1211);
nor U1274 (N_1274,N_1219,N_1251);
nand U1275 (N_1275,N_1227,N_1225);
nand U1276 (N_1276,N_1223,N_1253);
or U1277 (N_1277,N_1206,N_1250);
nand U1278 (N_1278,N_1226,N_1231);
and U1279 (N_1279,N_1234,N_1242);
nand U1280 (N_1280,N_1244,N_1257);
nor U1281 (N_1281,N_1247,N_1215);
or U1282 (N_1282,N_1221,N_1232);
nor U1283 (N_1283,N_1254,N_1200);
and U1284 (N_1284,N_1229,N_1214);
and U1285 (N_1285,N_1237,N_1240);
nand U1286 (N_1286,N_1235,N_1202);
xnor U1287 (N_1287,N_1213,N_1210);
and U1288 (N_1288,N_1228,N_1216);
or U1289 (N_1289,N_1252,N_1256);
or U1290 (N_1290,N_1226,N_1203);
and U1291 (N_1291,N_1226,N_1235);
or U1292 (N_1292,N_1244,N_1255);
or U1293 (N_1293,N_1202,N_1211);
and U1294 (N_1294,N_1227,N_1244);
or U1295 (N_1295,N_1229,N_1216);
nor U1296 (N_1296,N_1208,N_1203);
or U1297 (N_1297,N_1257,N_1200);
or U1298 (N_1298,N_1213,N_1256);
and U1299 (N_1299,N_1257,N_1232);
and U1300 (N_1300,N_1230,N_1248);
or U1301 (N_1301,N_1202,N_1255);
and U1302 (N_1302,N_1206,N_1229);
and U1303 (N_1303,N_1245,N_1248);
and U1304 (N_1304,N_1222,N_1217);
nor U1305 (N_1305,N_1203,N_1251);
nand U1306 (N_1306,N_1258,N_1216);
nor U1307 (N_1307,N_1228,N_1246);
nor U1308 (N_1308,N_1210,N_1212);
nand U1309 (N_1309,N_1237,N_1228);
or U1310 (N_1310,N_1258,N_1245);
nand U1311 (N_1311,N_1237,N_1242);
nor U1312 (N_1312,N_1243,N_1203);
and U1313 (N_1313,N_1253,N_1236);
nand U1314 (N_1314,N_1203,N_1238);
nand U1315 (N_1315,N_1238,N_1216);
or U1316 (N_1316,N_1234,N_1212);
nand U1317 (N_1317,N_1242,N_1210);
and U1318 (N_1318,N_1222,N_1250);
nand U1319 (N_1319,N_1206,N_1254);
nor U1320 (N_1320,N_1270,N_1310);
nor U1321 (N_1321,N_1309,N_1266);
nor U1322 (N_1322,N_1276,N_1278);
nor U1323 (N_1323,N_1287,N_1274);
or U1324 (N_1324,N_1281,N_1279);
or U1325 (N_1325,N_1265,N_1282);
or U1326 (N_1326,N_1316,N_1303);
nand U1327 (N_1327,N_1271,N_1298);
or U1328 (N_1328,N_1285,N_1299);
nor U1329 (N_1329,N_1305,N_1277);
nand U1330 (N_1330,N_1313,N_1283);
and U1331 (N_1331,N_1302,N_1262);
nor U1332 (N_1332,N_1267,N_1263);
nand U1333 (N_1333,N_1289,N_1264);
nor U1334 (N_1334,N_1296,N_1288);
or U1335 (N_1335,N_1273,N_1272);
or U1336 (N_1336,N_1314,N_1300);
nor U1337 (N_1337,N_1268,N_1312);
nor U1338 (N_1338,N_1297,N_1306);
nor U1339 (N_1339,N_1293,N_1290);
and U1340 (N_1340,N_1318,N_1294);
nor U1341 (N_1341,N_1319,N_1307);
xnor U1342 (N_1342,N_1286,N_1260);
and U1343 (N_1343,N_1304,N_1275);
and U1344 (N_1344,N_1301,N_1308);
and U1345 (N_1345,N_1291,N_1280);
nand U1346 (N_1346,N_1295,N_1261);
nand U1347 (N_1347,N_1269,N_1284);
nand U1348 (N_1348,N_1292,N_1315);
nand U1349 (N_1349,N_1311,N_1317);
or U1350 (N_1350,N_1263,N_1296);
nor U1351 (N_1351,N_1263,N_1304);
and U1352 (N_1352,N_1303,N_1271);
or U1353 (N_1353,N_1282,N_1272);
nor U1354 (N_1354,N_1264,N_1300);
or U1355 (N_1355,N_1273,N_1285);
nor U1356 (N_1356,N_1281,N_1317);
and U1357 (N_1357,N_1265,N_1261);
or U1358 (N_1358,N_1302,N_1279);
nand U1359 (N_1359,N_1299,N_1309);
nand U1360 (N_1360,N_1298,N_1275);
xnor U1361 (N_1361,N_1268,N_1317);
nand U1362 (N_1362,N_1277,N_1313);
or U1363 (N_1363,N_1289,N_1311);
nor U1364 (N_1364,N_1270,N_1282);
and U1365 (N_1365,N_1313,N_1267);
nand U1366 (N_1366,N_1297,N_1313);
nand U1367 (N_1367,N_1289,N_1310);
nand U1368 (N_1368,N_1293,N_1277);
and U1369 (N_1369,N_1271,N_1314);
and U1370 (N_1370,N_1297,N_1276);
nand U1371 (N_1371,N_1264,N_1306);
and U1372 (N_1372,N_1300,N_1292);
nor U1373 (N_1373,N_1284,N_1317);
and U1374 (N_1374,N_1263,N_1270);
or U1375 (N_1375,N_1268,N_1263);
or U1376 (N_1376,N_1261,N_1270);
or U1377 (N_1377,N_1306,N_1312);
nor U1378 (N_1378,N_1261,N_1264);
and U1379 (N_1379,N_1288,N_1291);
nor U1380 (N_1380,N_1341,N_1377);
nor U1381 (N_1381,N_1354,N_1359);
and U1382 (N_1382,N_1362,N_1333);
nand U1383 (N_1383,N_1339,N_1324);
nor U1384 (N_1384,N_1357,N_1371);
nor U1385 (N_1385,N_1358,N_1326);
or U1386 (N_1386,N_1334,N_1355);
nor U1387 (N_1387,N_1348,N_1369);
or U1388 (N_1388,N_1370,N_1321);
nor U1389 (N_1389,N_1378,N_1323);
and U1390 (N_1390,N_1379,N_1350);
or U1391 (N_1391,N_1353,N_1366);
and U1392 (N_1392,N_1360,N_1336);
and U1393 (N_1393,N_1340,N_1364);
or U1394 (N_1394,N_1356,N_1349);
xnor U1395 (N_1395,N_1347,N_1375);
or U1396 (N_1396,N_1376,N_1367);
or U1397 (N_1397,N_1363,N_1346);
and U1398 (N_1398,N_1372,N_1332);
nand U1399 (N_1399,N_1322,N_1328);
nor U1400 (N_1400,N_1351,N_1344);
and U1401 (N_1401,N_1330,N_1368);
or U1402 (N_1402,N_1374,N_1320);
and U1403 (N_1403,N_1373,N_1337);
nand U1404 (N_1404,N_1345,N_1331);
xor U1405 (N_1405,N_1342,N_1361);
nor U1406 (N_1406,N_1338,N_1352);
nand U1407 (N_1407,N_1329,N_1335);
nand U1408 (N_1408,N_1365,N_1343);
or U1409 (N_1409,N_1327,N_1325);
nor U1410 (N_1410,N_1371,N_1339);
nor U1411 (N_1411,N_1337,N_1351);
or U1412 (N_1412,N_1344,N_1378);
nor U1413 (N_1413,N_1330,N_1334);
nand U1414 (N_1414,N_1377,N_1370);
nand U1415 (N_1415,N_1364,N_1375);
nand U1416 (N_1416,N_1343,N_1370);
nand U1417 (N_1417,N_1344,N_1367);
nor U1418 (N_1418,N_1373,N_1376);
or U1419 (N_1419,N_1330,N_1346);
xor U1420 (N_1420,N_1360,N_1359);
nand U1421 (N_1421,N_1320,N_1349);
or U1422 (N_1422,N_1352,N_1323);
nor U1423 (N_1423,N_1320,N_1330);
and U1424 (N_1424,N_1348,N_1370);
and U1425 (N_1425,N_1329,N_1366);
nor U1426 (N_1426,N_1327,N_1365);
and U1427 (N_1427,N_1369,N_1362);
or U1428 (N_1428,N_1362,N_1346);
or U1429 (N_1429,N_1375,N_1341);
or U1430 (N_1430,N_1358,N_1324);
nand U1431 (N_1431,N_1366,N_1350);
or U1432 (N_1432,N_1322,N_1365);
or U1433 (N_1433,N_1346,N_1373);
nor U1434 (N_1434,N_1374,N_1340);
or U1435 (N_1435,N_1367,N_1355);
nand U1436 (N_1436,N_1358,N_1334);
or U1437 (N_1437,N_1320,N_1350);
nor U1438 (N_1438,N_1359,N_1372);
or U1439 (N_1439,N_1362,N_1352);
or U1440 (N_1440,N_1394,N_1424);
and U1441 (N_1441,N_1411,N_1420);
nand U1442 (N_1442,N_1383,N_1431);
nand U1443 (N_1443,N_1400,N_1432);
nor U1444 (N_1444,N_1412,N_1435);
and U1445 (N_1445,N_1415,N_1428);
nand U1446 (N_1446,N_1398,N_1439);
xnor U1447 (N_1447,N_1392,N_1436);
nor U1448 (N_1448,N_1417,N_1429);
and U1449 (N_1449,N_1393,N_1416);
or U1450 (N_1450,N_1410,N_1401);
nor U1451 (N_1451,N_1382,N_1399);
nand U1452 (N_1452,N_1387,N_1381);
or U1453 (N_1453,N_1437,N_1395);
nor U1454 (N_1454,N_1385,N_1407);
nand U1455 (N_1455,N_1404,N_1426);
xor U1456 (N_1456,N_1388,N_1430);
or U1457 (N_1457,N_1409,N_1419);
nor U1458 (N_1458,N_1438,N_1423);
or U1459 (N_1459,N_1402,N_1413);
nor U1460 (N_1460,N_1389,N_1434);
and U1461 (N_1461,N_1406,N_1425);
or U1462 (N_1462,N_1427,N_1396);
and U1463 (N_1463,N_1397,N_1418);
and U1464 (N_1464,N_1391,N_1380);
nand U1465 (N_1465,N_1384,N_1421);
nand U1466 (N_1466,N_1408,N_1433);
nor U1467 (N_1467,N_1414,N_1422);
nor U1468 (N_1468,N_1386,N_1403);
and U1469 (N_1469,N_1390,N_1405);
and U1470 (N_1470,N_1383,N_1416);
nor U1471 (N_1471,N_1428,N_1420);
nand U1472 (N_1472,N_1411,N_1433);
nand U1473 (N_1473,N_1435,N_1396);
nand U1474 (N_1474,N_1434,N_1384);
or U1475 (N_1475,N_1406,N_1416);
and U1476 (N_1476,N_1417,N_1410);
nor U1477 (N_1477,N_1403,N_1410);
nand U1478 (N_1478,N_1408,N_1380);
or U1479 (N_1479,N_1437,N_1438);
and U1480 (N_1480,N_1395,N_1392);
nor U1481 (N_1481,N_1427,N_1428);
nand U1482 (N_1482,N_1404,N_1388);
nor U1483 (N_1483,N_1389,N_1397);
nand U1484 (N_1484,N_1391,N_1388);
and U1485 (N_1485,N_1411,N_1405);
or U1486 (N_1486,N_1392,N_1434);
or U1487 (N_1487,N_1395,N_1407);
or U1488 (N_1488,N_1382,N_1400);
nand U1489 (N_1489,N_1387,N_1410);
or U1490 (N_1490,N_1400,N_1392);
nand U1491 (N_1491,N_1394,N_1430);
nor U1492 (N_1492,N_1438,N_1386);
nor U1493 (N_1493,N_1382,N_1390);
or U1494 (N_1494,N_1380,N_1406);
and U1495 (N_1495,N_1387,N_1394);
nor U1496 (N_1496,N_1412,N_1411);
nand U1497 (N_1497,N_1432,N_1388);
or U1498 (N_1498,N_1405,N_1427);
nand U1499 (N_1499,N_1415,N_1413);
and U1500 (N_1500,N_1459,N_1447);
and U1501 (N_1501,N_1465,N_1491);
and U1502 (N_1502,N_1446,N_1450);
nand U1503 (N_1503,N_1480,N_1473);
or U1504 (N_1504,N_1474,N_1444);
nand U1505 (N_1505,N_1443,N_1485);
and U1506 (N_1506,N_1497,N_1471);
or U1507 (N_1507,N_1453,N_1489);
or U1508 (N_1508,N_1448,N_1445);
or U1509 (N_1509,N_1498,N_1470);
nor U1510 (N_1510,N_1496,N_1455);
or U1511 (N_1511,N_1463,N_1440);
nor U1512 (N_1512,N_1449,N_1486);
or U1513 (N_1513,N_1468,N_1457);
nor U1514 (N_1514,N_1475,N_1456);
nor U1515 (N_1515,N_1482,N_1487);
nor U1516 (N_1516,N_1483,N_1462);
and U1517 (N_1517,N_1484,N_1454);
or U1518 (N_1518,N_1452,N_1464);
nor U1519 (N_1519,N_1490,N_1495);
nor U1520 (N_1520,N_1467,N_1493);
xnor U1521 (N_1521,N_1494,N_1460);
or U1522 (N_1522,N_1499,N_1441);
or U1523 (N_1523,N_1461,N_1492);
nand U1524 (N_1524,N_1478,N_1479);
or U1525 (N_1525,N_1476,N_1472);
or U1526 (N_1526,N_1488,N_1481);
nand U1527 (N_1527,N_1477,N_1469);
nor U1528 (N_1528,N_1458,N_1466);
and U1529 (N_1529,N_1442,N_1451);
xnor U1530 (N_1530,N_1442,N_1471);
nand U1531 (N_1531,N_1446,N_1489);
or U1532 (N_1532,N_1493,N_1485);
or U1533 (N_1533,N_1465,N_1463);
and U1534 (N_1534,N_1491,N_1479);
nand U1535 (N_1535,N_1478,N_1447);
nand U1536 (N_1536,N_1493,N_1480);
and U1537 (N_1537,N_1476,N_1496);
nor U1538 (N_1538,N_1486,N_1492);
or U1539 (N_1539,N_1470,N_1487);
and U1540 (N_1540,N_1484,N_1452);
nor U1541 (N_1541,N_1444,N_1442);
or U1542 (N_1542,N_1444,N_1440);
or U1543 (N_1543,N_1442,N_1450);
or U1544 (N_1544,N_1462,N_1476);
or U1545 (N_1545,N_1484,N_1488);
and U1546 (N_1546,N_1453,N_1497);
nor U1547 (N_1547,N_1480,N_1492);
nand U1548 (N_1548,N_1442,N_1486);
and U1549 (N_1549,N_1494,N_1489);
and U1550 (N_1550,N_1458,N_1452);
and U1551 (N_1551,N_1475,N_1491);
nand U1552 (N_1552,N_1491,N_1449);
nand U1553 (N_1553,N_1481,N_1494);
nor U1554 (N_1554,N_1474,N_1459);
nor U1555 (N_1555,N_1481,N_1485);
and U1556 (N_1556,N_1471,N_1495);
nor U1557 (N_1557,N_1463,N_1479);
nand U1558 (N_1558,N_1499,N_1473);
nand U1559 (N_1559,N_1458,N_1442);
nor U1560 (N_1560,N_1533,N_1535);
and U1561 (N_1561,N_1545,N_1538);
or U1562 (N_1562,N_1518,N_1507);
or U1563 (N_1563,N_1546,N_1536);
nand U1564 (N_1564,N_1532,N_1511);
nand U1565 (N_1565,N_1557,N_1549);
nor U1566 (N_1566,N_1504,N_1520);
nor U1567 (N_1567,N_1502,N_1550);
and U1568 (N_1568,N_1558,N_1509);
nor U1569 (N_1569,N_1528,N_1534);
nand U1570 (N_1570,N_1503,N_1543);
nand U1571 (N_1571,N_1510,N_1512);
nand U1572 (N_1572,N_1553,N_1526);
and U1573 (N_1573,N_1519,N_1552);
nor U1574 (N_1574,N_1506,N_1539);
nand U1575 (N_1575,N_1554,N_1500);
and U1576 (N_1576,N_1505,N_1525);
nand U1577 (N_1577,N_1541,N_1537);
nor U1578 (N_1578,N_1555,N_1508);
nor U1579 (N_1579,N_1531,N_1540);
nor U1580 (N_1580,N_1524,N_1551);
or U1581 (N_1581,N_1530,N_1515);
or U1582 (N_1582,N_1544,N_1522);
or U1583 (N_1583,N_1527,N_1513);
and U1584 (N_1584,N_1547,N_1529);
and U1585 (N_1585,N_1521,N_1548);
and U1586 (N_1586,N_1514,N_1516);
and U1587 (N_1587,N_1517,N_1523);
or U1588 (N_1588,N_1559,N_1556);
nor U1589 (N_1589,N_1542,N_1501);
or U1590 (N_1590,N_1533,N_1504);
and U1591 (N_1591,N_1533,N_1544);
nor U1592 (N_1592,N_1554,N_1544);
nor U1593 (N_1593,N_1516,N_1517);
nand U1594 (N_1594,N_1542,N_1511);
and U1595 (N_1595,N_1538,N_1501);
nand U1596 (N_1596,N_1501,N_1547);
nor U1597 (N_1597,N_1541,N_1502);
nor U1598 (N_1598,N_1502,N_1523);
nor U1599 (N_1599,N_1550,N_1545);
or U1600 (N_1600,N_1534,N_1520);
or U1601 (N_1601,N_1521,N_1523);
and U1602 (N_1602,N_1547,N_1500);
or U1603 (N_1603,N_1527,N_1536);
nor U1604 (N_1604,N_1555,N_1509);
nand U1605 (N_1605,N_1505,N_1508);
nor U1606 (N_1606,N_1557,N_1538);
and U1607 (N_1607,N_1547,N_1506);
and U1608 (N_1608,N_1525,N_1508);
nand U1609 (N_1609,N_1521,N_1527);
xor U1610 (N_1610,N_1503,N_1504);
or U1611 (N_1611,N_1502,N_1507);
and U1612 (N_1612,N_1521,N_1505);
or U1613 (N_1613,N_1534,N_1509);
nand U1614 (N_1614,N_1541,N_1526);
nand U1615 (N_1615,N_1509,N_1551);
and U1616 (N_1616,N_1538,N_1552);
and U1617 (N_1617,N_1558,N_1501);
nand U1618 (N_1618,N_1518,N_1556);
or U1619 (N_1619,N_1505,N_1507);
nand U1620 (N_1620,N_1564,N_1611);
or U1621 (N_1621,N_1596,N_1587);
nor U1622 (N_1622,N_1589,N_1616);
nor U1623 (N_1623,N_1588,N_1570);
and U1624 (N_1624,N_1583,N_1579);
and U1625 (N_1625,N_1561,N_1591);
and U1626 (N_1626,N_1614,N_1573);
nand U1627 (N_1627,N_1574,N_1562);
nand U1628 (N_1628,N_1590,N_1592);
and U1629 (N_1629,N_1563,N_1577);
and U1630 (N_1630,N_1607,N_1604);
nand U1631 (N_1631,N_1602,N_1615);
and U1632 (N_1632,N_1560,N_1618);
nor U1633 (N_1633,N_1609,N_1608);
or U1634 (N_1634,N_1600,N_1568);
xor U1635 (N_1635,N_1581,N_1593);
and U1636 (N_1636,N_1603,N_1601);
or U1637 (N_1637,N_1572,N_1565);
and U1638 (N_1638,N_1571,N_1595);
nor U1639 (N_1639,N_1586,N_1599);
nor U1640 (N_1640,N_1594,N_1597);
nand U1641 (N_1641,N_1567,N_1569);
and U1642 (N_1642,N_1606,N_1605);
nor U1643 (N_1643,N_1613,N_1582);
or U1644 (N_1644,N_1584,N_1610);
or U1645 (N_1645,N_1580,N_1566);
and U1646 (N_1646,N_1585,N_1598);
or U1647 (N_1647,N_1578,N_1612);
nor U1648 (N_1648,N_1619,N_1575);
nand U1649 (N_1649,N_1576,N_1617);
or U1650 (N_1650,N_1572,N_1614);
or U1651 (N_1651,N_1603,N_1591);
nor U1652 (N_1652,N_1613,N_1564);
or U1653 (N_1653,N_1571,N_1565);
nor U1654 (N_1654,N_1593,N_1608);
nor U1655 (N_1655,N_1607,N_1561);
and U1656 (N_1656,N_1575,N_1564);
and U1657 (N_1657,N_1583,N_1582);
nand U1658 (N_1658,N_1560,N_1566);
nor U1659 (N_1659,N_1562,N_1617);
nor U1660 (N_1660,N_1604,N_1588);
nand U1661 (N_1661,N_1570,N_1600);
nand U1662 (N_1662,N_1565,N_1575);
nor U1663 (N_1663,N_1581,N_1567);
nand U1664 (N_1664,N_1562,N_1585);
or U1665 (N_1665,N_1618,N_1601);
and U1666 (N_1666,N_1586,N_1577);
nand U1667 (N_1667,N_1590,N_1574);
or U1668 (N_1668,N_1596,N_1608);
nor U1669 (N_1669,N_1597,N_1582);
and U1670 (N_1670,N_1614,N_1580);
nand U1671 (N_1671,N_1619,N_1563);
nor U1672 (N_1672,N_1581,N_1562);
and U1673 (N_1673,N_1589,N_1598);
nor U1674 (N_1674,N_1575,N_1560);
and U1675 (N_1675,N_1609,N_1591);
and U1676 (N_1676,N_1595,N_1563);
nor U1677 (N_1677,N_1570,N_1607);
nor U1678 (N_1678,N_1574,N_1594);
nor U1679 (N_1679,N_1619,N_1589);
nor U1680 (N_1680,N_1621,N_1676);
and U1681 (N_1681,N_1646,N_1642);
nor U1682 (N_1682,N_1653,N_1647);
nor U1683 (N_1683,N_1672,N_1641);
or U1684 (N_1684,N_1645,N_1678);
nor U1685 (N_1685,N_1664,N_1666);
or U1686 (N_1686,N_1656,N_1628);
or U1687 (N_1687,N_1669,N_1667);
or U1688 (N_1688,N_1662,N_1626);
nor U1689 (N_1689,N_1630,N_1632);
nor U1690 (N_1690,N_1650,N_1637);
nand U1691 (N_1691,N_1640,N_1655);
and U1692 (N_1692,N_1643,N_1638);
nand U1693 (N_1693,N_1674,N_1624);
and U1694 (N_1694,N_1623,N_1654);
and U1695 (N_1695,N_1673,N_1663);
nand U1696 (N_1696,N_1644,N_1651);
or U1697 (N_1697,N_1649,N_1629);
or U1698 (N_1698,N_1679,N_1657);
or U1699 (N_1699,N_1635,N_1633);
nor U1700 (N_1700,N_1660,N_1639);
nand U1701 (N_1701,N_1670,N_1625);
nand U1702 (N_1702,N_1668,N_1636);
nand U1703 (N_1703,N_1620,N_1622);
nand U1704 (N_1704,N_1627,N_1634);
and U1705 (N_1705,N_1631,N_1677);
nand U1706 (N_1706,N_1658,N_1665);
or U1707 (N_1707,N_1652,N_1659);
or U1708 (N_1708,N_1671,N_1661);
nor U1709 (N_1709,N_1648,N_1675);
or U1710 (N_1710,N_1641,N_1633);
or U1711 (N_1711,N_1678,N_1669);
or U1712 (N_1712,N_1676,N_1647);
nand U1713 (N_1713,N_1665,N_1643);
and U1714 (N_1714,N_1622,N_1624);
or U1715 (N_1715,N_1670,N_1676);
nand U1716 (N_1716,N_1672,N_1677);
and U1717 (N_1717,N_1627,N_1623);
or U1718 (N_1718,N_1679,N_1673);
or U1719 (N_1719,N_1669,N_1646);
xor U1720 (N_1720,N_1659,N_1667);
xnor U1721 (N_1721,N_1669,N_1626);
or U1722 (N_1722,N_1661,N_1633);
xor U1723 (N_1723,N_1663,N_1630);
or U1724 (N_1724,N_1673,N_1654);
or U1725 (N_1725,N_1677,N_1666);
or U1726 (N_1726,N_1653,N_1635);
or U1727 (N_1727,N_1643,N_1631);
or U1728 (N_1728,N_1636,N_1673);
and U1729 (N_1729,N_1649,N_1670);
nand U1730 (N_1730,N_1639,N_1648);
xnor U1731 (N_1731,N_1653,N_1641);
or U1732 (N_1732,N_1664,N_1675);
and U1733 (N_1733,N_1620,N_1624);
nor U1734 (N_1734,N_1638,N_1644);
or U1735 (N_1735,N_1626,N_1634);
nand U1736 (N_1736,N_1666,N_1652);
or U1737 (N_1737,N_1648,N_1673);
and U1738 (N_1738,N_1661,N_1643);
or U1739 (N_1739,N_1630,N_1626);
or U1740 (N_1740,N_1703,N_1734);
xnor U1741 (N_1741,N_1683,N_1701);
and U1742 (N_1742,N_1716,N_1736);
or U1743 (N_1743,N_1682,N_1697);
and U1744 (N_1744,N_1691,N_1728);
nand U1745 (N_1745,N_1706,N_1702);
nand U1746 (N_1746,N_1727,N_1729);
nor U1747 (N_1747,N_1709,N_1695);
or U1748 (N_1748,N_1684,N_1721);
or U1749 (N_1749,N_1719,N_1693);
nor U1750 (N_1750,N_1688,N_1720);
nor U1751 (N_1751,N_1685,N_1717);
nand U1752 (N_1752,N_1733,N_1699);
or U1753 (N_1753,N_1714,N_1686);
and U1754 (N_1754,N_1726,N_1698);
nor U1755 (N_1755,N_1724,N_1687);
or U1756 (N_1756,N_1704,N_1680);
or U1757 (N_1757,N_1737,N_1681);
and U1758 (N_1758,N_1713,N_1692);
and U1759 (N_1759,N_1708,N_1725);
nand U1760 (N_1760,N_1707,N_1696);
nand U1761 (N_1761,N_1722,N_1705);
or U1762 (N_1762,N_1690,N_1700);
xor U1763 (N_1763,N_1718,N_1732);
and U1764 (N_1764,N_1689,N_1730);
nor U1765 (N_1765,N_1712,N_1738);
nand U1766 (N_1766,N_1739,N_1710);
nand U1767 (N_1767,N_1694,N_1711);
nor U1768 (N_1768,N_1723,N_1715);
nor U1769 (N_1769,N_1731,N_1735);
nor U1770 (N_1770,N_1688,N_1717);
or U1771 (N_1771,N_1704,N_1718);
xor U1772 (N_1772,N_1715,N_1688);
nand U1773 (N_1773,N_1681,N_1705);
nor U1774 (N_1774,N_1739,N_1689);
or U1775 (N_1775,N_1714,N_1688);
nor U1776 (N_1776,N_1704,N_1685);
and U1777 (N_1777,N_1737,N_1716);
and U1778 (N_1778,N_1699,N_1739);
nor U1779 (N_1779,N_1721,N_1720);
or U1780 (N_1780,N_1716,N_1686);
and U1781 (N_1781,N_1737,N_1703);
nand U1782 (N_1782,N_1735,N_1707);
and U1783 (N_1783,N_1723,N_1712);
nor U1784 (N_1784,N_1725,N_1688);
nor U1785 (N_1785,N_1680,N_1706);
and U1786 (N_1786,N_1723,N_1695);
nor U1787 (N_1787,N_1688,N_1686);
nor U1788 (N_1788,N_1687,N_1727);
or U1789 (N_1789,N_1695,N_1685);
or U1790 (N_1790,N_1729,N_1711);
nor U1791 (N_1791,N_1683,N_1732);
nor U1792 (N_1792,N_1706,N_1722);
or U1793 (N_1793,N_1685,N_1693);
and U1794 (N_1794,N_1725,N_1735);
nor U1795 (N_1795,N_1685,N_1729);
or U1796 (N_1796,N_1728,N_1686);
or U1797 (N_1797,N_1714,N_1732);
or U1798 (N_1798,N_1716,N_1705);
and U1799 (N_1799,N_1739,N_1707);
and U1800 (N_1800,N_1755,N_1774);
or U1801 (N_1801,N_1747,N_1753);
or U1802 (N_1802,N_1743,N_1761);
xor U1803 (N_1803,N_1799,N_1760);
and U1804 (N_1804,N_1784,N_1778);
or U1805 (N_1805,N_1756,N_1757);
nor U1806 (N_1806,N_1793,N_1762);
or U1807 (N_1807,N_1790,N_1789);
nor U1808 (N_1808,N_1770,N_1740);
nand U1809 (N_1809,N_1779,N_1748);
and U1810 (N_1810,N_1785,N_1752);
nor U1811 (N_1811,N_1768,N_1754);
and U1812 (N_1812,N_1741,N_1777);
or U1813 (N_1813,N_1750,N_1765);
nand U1814 (N_1814,N_1749,N_1783);
or U1815 (N_1815,N_1742,N_1782);
nor U1816 (N_1816,N_1795,N_1764);
nand U1817 (N_1817,N_1773,N_1767);
and U1818 (N_1818,N_1781,N_1744);
nand U1819 (N_1819,N_1745,N_1792);
and U1820 (N_1820,N_1772,N_1776);
nand U1821 (N_1821,N_1775,N_1796);
nand U1822 (N_1822,N_1763,N_1751);
nor U1823 (N_1823,N_1766,N_1798);
nand U1824 (N_1824,N_1791,N_1746);
nand U1825 (N_1825,N_1794,N_1787);
xnor U1826 (N_1826,N_1788,N_1769);
xnor U1827 (N_1827,N_1758,N_1797);
or U1828 (N_1828,N_1780,N_1786);
and U1829 (N_1829,N_1759,N_1771);
or U1830 (N_1830,N_1769,N_1741);
nor U1831 (N_1831,N_1755,N_1760);
nor U1832 (N_1832,N_1782,N_1788);
nand U1833 (N_1833,N_1753,N_1778);
and U1834 (N_1834,N_1753,N_1784);
nor U1835 (N_1835,N_1775,N_1759);
nand U1836 (N_1836,N_1796,N_1794);
nand U1837 (N_1837,N_1758,N_1756);
nand U1838 (N_1838,N_1773,N_1764);
nor U1839 (N_1839,N_1752,N_1740);
and U1840 (N_1840,N_1753,N_1791);
nor U1841 (N_1841,N_1776,N_1771);
nor U1842 (N_1842,N_1787,N_1759);
or U1843 (N_1843,N_1768,N_1755);
or U1844 (N_1844,N_1752,N_1773);
or U1845 (N_1845,N_1781,N_1796);
or U1846 (N_1846,N_1748,N_1796);
nor U1847 (N_1847,N_1757,N_1796);
nand U1848 (N_1848,N_1774,N_1746);
nand U1849 (N_1849,N_1757,N_1760);
nor U1850 (N_1850,N_1777,N_1755);
nor U1851 (N_1851,N_1748,N_1771);
nand U1852 (N_1852,N_1798,N_1786);
and U1853 (N_1853,N_1784,N_1771);
nor U1854 (N_1854,N_1790,N_1745);
xnor U1855 (N_1855,N_1787,N_1774);
nor U1856 (N_1856,N_1777,N_1764);
nor U1857 (N_1857,N_1753,N_1745);
nand U1858 (N_1858,N_1787,N_1769);
nor U1859 (N_1859,N_1782,N_1756);
nor U1860 (N_1860,N_1819,N_1801);
or U1861 (N_1861,N_1843,N_1825);
xnor U1862 (N_1862,N_1855,N_1836);
and U1863 (N_1863,N_1847,N_1858);
and U1864 (N_1864,N_1829,N_1802);
nand U1865 (N_1865,N_1850,N_1822);
nand U1866 (N_1866,N_1828,N_1811);
nand U1867 (N_1867,N_1837,N_1817);
and U1868 (N_1868,N_1851,N_1834);
or U1869 (N_1869,N_1835,N_1852);
or U1870 (N_1870,N_1857,N_1823);
and U1871 (N_1871,N_1821,N_1814);
or U1872 (N_1872,N_1842,N_1804);
and U1873 (N_1873,N_1846,N_1854);
nand U1874 (N_1874,N_1813,N_1853);
or U1875 (N_1875,N_1830,N_1856);
or U1876 (N_1876,N_1810,N_1820);
or U1877 (N_1877,N_1859,N_1845);
nand U1878 (N_1878,N_1806,N_1849);
or U1879 (N_1879,N_1839,N_1815);
nor U1880 (N_1880,N_1827,N_1844);
nor U1881 (N_1881,N_1826,N_1840);
nor U1882 (N_1882,N_1812,N_1805);
or U1883 (N_1883,N_1807,N_1831);
nor U1884 (N_1884,N_1800,N_1841);
or U1885 (N_1885,N_1816,N_1824);
nor U1886 (N_1886,N_1803,N_1838);
nor U1887 (N_1887,N_1832,N_1848);
and U1888 (N_1888,N_1818,N_1808);
nor U1889 (N_1889,N_1809,N_1833);
nand U1890 (N_1890,N_1818,N_1830);
or U1891 (N_1891,N_1826,N_1801);
and U1892 (N_1892,N_1856,N_1840);
nand U1893 (N_1893,N_1835,N_1843);
nor U1894 (N_1894,N_1829,N_1844);
or U1895 (N_1895,N_1827,N_1840);
nand U1896 (N_1896,N_1825,N_1810);
nand U1897 (N_1897,N_1810,N_1819);
and U1898 (N_1898,N_1831,N_1822);
or U1899 (N_1899,N_1822,N_1829);
nor U1900 (N_1900,N_1845,N_1851);
and U1901 (N_1901,N_1809,N_1815);
nand U1902 (N_1902,N_1803,N_1852);
nand U1903 (N_1903,N_1816,N_1804);
or U1904 (N_1904,N_1841,N_1842);
and U1905 (N_1905,N_1800,N_1814);
and U1906 (N_1906,N_1842,N_1829);
or U1907 (N_1907,N_1820,N_1806);
or U1908 (N_1908,N_1822,N_1809);
nor U1909 (N_1909,N_1804,N_1855);
nand U1910 (N_1910,N_1856,N_1841);
nor U1911 (N_1911,N_1802,N_1833);
and U1912 (N_1912,N_1849,N_1811);
or U1913 (N_1913,N_1815,N_1855);
and U1914 (N_1914,N_1814,N_1846);
nand U1915 (N_1915,N_1819,N_1845);
and U1916 (N_1916,N_1827,N_1857);
nor U1917 (N_1917,N_1850,N_1801);
and U1918 (N_1918,N_1839,N_1858);
nand U1919 (N_1919,N_1859,N_1825);
nor U1920 (N_1920,N_1889,N_1861);
nand U1921 (N_1921,N_1894,N_1875);
and U1922 (N_1922,N_1892,N_1880);
nand U1923 (N_1923,N_1905,N_1907);
and U1924 (N_1924,N_1915,N_1873);
or U1925 (N_1925,N_1887,N_1908);
and U1926 (N_1926,N_1884,N_1866);
and U1927 (N_1927,N_1895,N_1865);
nand U1928 (N_1928,N_1913,N_1896);
nor U1929 (N_1929,N_1898,N_1882);
or U1930 (N_1930,N_1891,N_1899);
and U1931 (N_1931,N_1919,N_1888);
nor U1932 (N_1932,N_1863,N_1874);
or U1933 (N_1933,N_1869,N_1914);
nor U1934 (N_1934,N_1909,N_1878);
nand U1935 (N_1935,N_1877,N_1872);
nand U1936 (N_1936,N_1904,N_1912);
nand U1937 (N_1937,N_1864,N_1906);
and U1938 (N_1938,N_1870,N_1886);
or U1939 (N_1939,N_1910,N_1871);
and U1940 (N_1940,N_1916,N_1911);
or U1941 (N_1941,N_1867,N_1902);
and U1942 (N_1942,N_1868,N_1893);
and U1943 (N_1943,N_1917,N_1876);
or U1944 (N_1944,N_1890,N_1918);
and U1945 (N_1945,N_1900,N_1879);
or U1946 (N_1946,N_1903,N_1901);
or U1947 (N_1947,N_1862,N_1897);
nor U1948 (N_1948,N_1881,N_1883);
nand U1949 (N_1949,N_1885,N_1860);
nor U1950 (N_1950,N_1862,N_1888);
or U1951 (N_1951,N_1915,N_1867);
and U1952 (N_1952,N_1861,N_1909);
nor U1953 (N_1953,N_1877,N_1906);
nor U1954 (N_1954,N_1869,N_1888);
and U1955 (N_1955,N_1901,N_1861);
or U1956 (N_1956,N_1915,N_1902);
xor U1957 (N_1957,N_1889,N_1906);
and U1958 (N_1958,N_1917,N_1880);
and U1959 (N_1959,N_1876,N_1903);
nor U1960 (N_1960,N_1871,N_1915);
and U1961 (N_1961,N_1867,N_1907);
and U1962 (N_1962,N_1866,N_1881);
nand U1963 (N_1963,N_1892,N_1867);
or U1964 (N_1964,N_1898,N_1902);
and U1965 (N_1965,N_1881,N_1860);
nor U1966 (N_1966,N_1885,N_1884);
nor U1967 (N_1967,N_1883,N_1889);
nand U1968 (N_1968,N_1918,N_1883);
nand U1969 (N_1969,N_1864,N_1901);
and U1970 (N_1970,N_1883,N_1873);
nor U1971 (N_1971,N_1864,N_1918);
nand U1972 (N_1972,N_1887,N_1897);
or U1973 (N_1973,N_1868,N_1885);
nand U1974 (N_1974,N_1863,N_1866);
nand U1975 (N_1975,N_1870,N_1891);
nor U1976 (N_1976,N_1897,N_1902);
nor U1977 (N_1977,N_1918,N_1908);
nor U1978 (N_1978,N_1871,N_1877);
and U1979 (N_1979,N_1901,N_1874);
nand U1980 (N_1980,N_1940,N_1924);
nor U1981 (N_1981,N_1952,N_1921);
or U1982 (N_1982,N_1935,N_1922);
nand U1983 (N_1983,N_1943,N_1964);
nand U1984 (N_1984,N_1933,N_1955);
nor U1985 (N_1985,N_1967,N_1936);
nand U1986 (N_1986,N_1966,N_1975);
nor U1987 (N_1987,N_1971,N_1972);
nor U1988 (N_1988,N_1979,N_1944);
nand U1989 (N_1989,N_1978,N_1925);
and U1990 (N_1990,N_1958,N_1934);
nor U1991 (N_1991,N_1928,N_1923);
or U1992 (N_1992,N_1954,N_1950);
nor U1993 (N_1993,N_1942,N_1956);
and U1994 (N_1994,N_1931,N_1977);
and U1995 (N_1995,N_1937,N_1945);
and U1996 (N_1996,N_1974,N_1951);
and U1997 (N_1997,N_1949,N_1947);
or U1998 (N_1998,N_1962,N_1920);
nor U1999 (N_1999,N_1929,N_1941);
nand U2000 (N_2000,N_1938,N_1953);
and U2001 (N_2001,N_1976,N_1959);
nor U2002 (N_2002,N_1957,N_1968);
or U2003 (N_2003,N_1961,N_1927);
nand U2004 (N_2004,N_1973,N_1946);
nand U2005 (N_2005,N_1963,N_1960);
and U2006 (N_2006,N_1930,N_1970);
or U2007 (N_2007,N_1965,N_1948);
nand U2008 (N_2008,N_1932,N_1969);
nor U2009 (N_2009,N_1926,N_1939);
nand U2010 (N_2010,N_1964,N_1969);
and U2011 (N_2011,N_1971,N_1920);
and U2012 (N_2012,N_1935,N_1967);
nor U2013 (N_2013,N_1958,N_1931);
nor U2014 (N_2014,N_1963,N_1945);
nand U2015 (N_2015,N_1923,N_1933);
and U2016 (N_2016,N_1935,N_1948);
nor U2017 (N_2017,N_1921,N_1944);
and U2018 (N_2018,N_1966,N_1953);
nor U2019 (N_2019,N_1977,N_1963);
nor U2020 (N_2020,N_1929,N_1970);
nand U2021 (N_2021,N_1959,N_1975);
nand U2022 (N_2022,N_1956,N_1968);
and U2023 (N_2023,N_1948,N_1975);
nor U2024 (N_2024,N_1946,N_1949);
nor U2025 (N_2025,N_1924,N_1945);
or U2026 (N_2026,N_1979,N_1971);
nand U2027 (N_2027,N_1926,N_1930);
nor U2028 (N_2028,N_1978,N_1922);
nor U2029 (N_2029,N_1922,N_1924);
or U2030 (N_2030,N_1954,N_1930);
and U2031 (N_2031,N_1957,N_1948);
and U2032 (N_2032,N_1969,N_1931);
and U2033 (N_2033,N_1928,N_1978);
or U2034 (N_2034,N_1933,N_1945);
nand U2035 (N_2035,N_1963,N_1937);
and U2036 (N_2036,N_1933,N_1924);
nor U2037 (N_2037,N_1930,N_1967);
nand U2038 (N_2038,N_1957,N_1939);
nand U2039 (N_2039,N_1977,N_1935);
or U2040 (N_2040,N_2011,N_1983);
xor U2041 (N_2041,N_1999,N_1997);
nor U2042 (N_2042,N_2017,N_2006);
or U2043 (N_2043,N_2005,N_2010);
nand U2044 (N_2044,N_2007,N_2009);
or U2045 (N_2045,N_2028,N_2020);
nor U2046 (N_2046,N_2036,N_1992);
or U2047 (N_2047,N_2031,N_1990);
or U2048 (N_2048,N_2029,N_2024);
nor U2049 (N_2049,N_2019,N_2033);
nand U2050 (N_2050,N_2000,N_2030);
nand U2051 (N_2051,N_1986,N_2012);
or U2052 (N_2052,N_2008,N_2003);
and U2053 (N_2053,N_1987,N_2026);
and U2054 (N_2054,N_2034,N_2032);
xnor U2055 (N_2055,N_2001,N_1991);
nand U2056 (N_2056,N_1988,N_2039);
nand U2057 (N_2057,N_1980,N_2023);
or U2058 (N_2058,N_1993,N_1985);
and U2059 (N_2059,N_2016,N_1981);
nor U2060 (N_2060,N_2035,N_2015);
or U2061 (N_2061,N_1982,N_2022);
or U2062 (N_2062,N_2002,N_2037);
or U2063 (N_2063,N_2013,N_2004);
or U2064 (N_2064,N_1995,N_1984);
and U2065 (N_2065,N_2021,N_2025);
nand U2066 (N_2066,N_2014,N_2018);
nand U2067 (N_2067,N_1996,N_2027);
nand U2068 (N_2068,N_2038,N_1998);
nand U2069 (N_2069,N_1989,N_1994);
and U2070 (N_2070,N_1998,N_2004);
and U2071 (N_2071,N_2022,N_2031);
and U2072 (N_2072,N_2021,N_2037);
or U2073 (N_2073,N_1991,N_2021);
or U2074 (N_2074,N_2015,N_1988);
and U2075 (N_2075,N_2038,N_1985);
or U2076 (N_2076,N_2036,N_2026);
nand U2077 (N_2077,N_2026,N_1980);
or U2078 (N_2078,N_2012,N_2039);
or U2079 (N_2079,N_2007,N_2022);
nor U2080 (N_2080,N_1999,N_2006);
nand U2081 (N_2081,N_1980,N_2013);
nor U2082 (N_2082,N_2015,N_2022);
and U2083 (N_2083,N_2031,N_1994);
nand U2084 (N_2084,N_1988,N_2034);
and U2085 (N_2085,N_1993,N_2029);
nor U2086 (N_2086,N_2012,N_2019);
and U2087 (N_2087,N_1990,N_2021);
nor U2088 (N_2088,N_1985,N_2001);
xnor U2089 (N_2089,N_2032,N_2033);
and U2090 (N_2090,N_2011,N_2007);
nand U2091 (N_2091,N_2007,N_1980);
nand U2092 (N_2092,N_1996,N_1994);
nor U2093 (N_2093,N_2001,N_2004);
nand U2094 (N_2094,N_1987,N_1998);
and U2095 (N_2095,N_1994,N_2013);
and U2096 (N_2096,N_2001,N_2006);
and U2097 (N_2097,N_2028,N_2026);
and U2098 (N_2098,N_2038,N_2036);
nor U2099 (N_2099,N_2002,N_2017);
and U2100 (N_2100,N_2084,N_2090);
or U2101 (N_2101,N_2086,N_2057);
nor U2102 (N_2102,N_2070,N_2048);
and U2103 (N_2103,N_2062,N_2046);
or U2104 (N_2104,N_2042,N_2093);
and U2105 (N_2105,N_2098,N_2050);
and U2106 (N_2106,N_2068,N_2079);
and U2107 (N_2107,N_2091,N_2044);
nand U2108 (N_2108,N_2097,N_2071);
and U2109 (N_2109,N_2052,N_2040);
and U2110 (N_2110,N_2082,N_2095);
or U2111 (N_2111,N_2054,N_2077);
nand U2112 (N_2112,N_2063,N_2094);
and U2113 (N_2113,N_2053,N_2092);
nor U2114 (N_2114,N_2059,N_2069);
or U2115 (N_2115,N_2087,N_2061);
or U2116 (N_2116,N_2088,N_2043);
or U2117 (N_2117,N_2072,N_2083);
nor U2118 (N_2118,N_2075,N_2073);
nor U2119 (N_2119,N_2080,N_2099);
nand U2120 (N_2120,N_2056,N_2060);
nor U2121 (N_2121,N_2065,N_2064);
nor U2122 (N_2122,N_2078,N_2076);
nor U2123 (N_2123,N_2074,N_2051);
and U2124 (N_2124,N_2067,N_2089);
or U2125 (N_2125,N_2049,N_2055);
or U2126 (N_2126,N_2081,N_2058);
or U2127 (N_2127,N_2041,N_2045);
and U2128 (N_2128,N_2085,N_2066);
or U2129 (N_2129,N_2047,N_2096);
and U2130 (N_2130,N_2070,N_2045);
nand U2131 (N_2131,N_2055,N_2067);
and U2132 (N_2132,N_2080,N_2095);
xnor U2133 (N_2133,N_2081,N_2078);
or U2134 (N_2134,N_2058,N_2071);
nor U2135 (N_2135,N_2046,N_2090);
nor U2136 (N_2136,N_2088,N_2042);
or U2137 (N_2137,N_2069,N_2045);
and U2138 (N_2138,N_2096,N_2070);
or U2139 (N_2139,N_2068,N_2094);
xor U2140 (N_2140,N_2073,N_2043);
nor U2141 (N_2141,N_2074,N_2084);
xor U2142 (N_2142,N_2099,N_2045);
nor U2143 (N_2143,N_2075,N_2045);
nor U2144 (N_2144,N_2074,N_2079);
or U2145 (N_2145,N_2092,N_2069);
or U2146 (N_2146,N_2077,N_2059);
and U2147 (N_2147,N_2076,N_2093);
and U2148 (N_2148,N_2059,N_2066);
and U2149 (N_2149,N_2056,N_2075);
or U2150 (N_2150,N_2087,N_2065);
and U2151 (N_2151,N_2072,N_2040);
xnor U2152 (N_2152,N_2041,N_2043);
xnor U2153 (N_2153,N_2067,N_2062);
nand U2154 (N_2154,N_2079,N_2093);
nand U2155 (N_2155,N_2041,N_2072);
nor U2156 (N_2156,N_2071,N_2065);
or U2157 (N_2157,N_2099,N_2073);
nor U2158 (N_2158,N_2097,N_2047);
nor U2159 (N_2159,N_2086,N_2044);
nor U2160 (N_2160,N_2133,N_2144);
nor U2161 (N_2161,N_2146,N_2151);
or U2162 (N_2162,N_2105,N_2153);
and U2163 (N_2163,N_2139,N_2113);
nor U2164 (N_2164,N_2134,N_2138);
or U2165 (N_2165,N_2100,N_2159);
or U2166 (N_2166,N_2130,N_2136);
nor U2167 (N_2167,N_2127,N_2121);
nor U2168 (N_2168,N_2118,N_2123);
or U2169 (N_2169,N_2106,N_2116);
and U2170 (N_2170,N_2117,N_2128);
nand U2171 (N_2171,N_2152,N_2135);
and U2172 (N_2172,N_2110,N_2141);
or U2173 (N_2173,N_2112,N_2119);
nand U2174 (N_2174,N_2115,N_2108);
or U2175 (N_2175,N_2114,N_2129);
and U2176 (N_2176,N_2132,N_2157);
or U2177 (N_2177,N_2148,N_2154);
nor U2178 (N_2178,N_2156,N_2158);
or U2179 (N_2179,N_2102,N_2147);
nor U2180 (N_2180,N_2143,N_2111);
or U2181 (N_2181,N_2104,N_2142);
nor U2182 (N_2182,N_2124,N_2150);
or U2183 (N_2183,N_2103,N_2126);
nor U2184 (N_2184,N_2145,N_2137);
and U2185 (N_2185,N_2101,N_2122);
nor U2186 (N_2186,N_2120,N_2125);
and U2187 (N_2187,N_2109,N_2107);
nor U2188 (N_2188,N_2149,N_2131);
xnor U2189 (N_2189,N_2140,N_2155);
nand U2190 (N_2190,N_2103,N_2107);
nand U2191 (N_2191,N_2126,N_2146);
nor U2192 (N_2192,N_2121,N_2135);
and U2193 (N_2193,N_2134,N_2123);
nand U2194 (N_2194,N_2148,N_2125);
or U2195 (N_2195,N_2121,N_2136);
xnor U2196 (N_2196,N_2126,N_2139);
nor U2197 (N_2197,N_2104,N_2101);
nor U2198 (N_2198,N_2147,N_2132);
nand U2199 (N_2199,N_2151,N_2106);
nand U2200 (N_2200,N_2151,N_2134);
and U2201 (N_2201,N_2114,N_2143);
or U2202 (N_2202,N_2134,N_2102);
nand U2203 (N_2203,N_2136,N_2126);
and U2204 (N_2204,N_2119,N_2148);
or U2205 (N_2205,N_2136,N_2141);
and U2206 (N_2206,N_2137,N_2121);
xor U2207 (N_2207,N_2140,N_2141);
xor U2208 (N_2208,N_2115,N_2149);
nand U2209 (N_2209,N_2152,N_2106);
and U2210 (N_2210,N_2151,N_2132);
nand U2211 (N_2211,N_2127,N_2124);
nor U2212 (N_2212,N_2159,N_2138);
nand U2213 (N_2213,N_2110,N_2114);
or U2214 (N_2214,N_2119,N_2101);
or U2215 (N_2215,N_2157,N_2134);
or U2216 (N_2216,N_2137,N_2116);
or U2217 (N_2217,N_2136,N_2125);
and U2218 (N_2218,N_2134,N_2133);
nand U2219 (N_2219,N_2156,N_2119);
and U2220 (N_2220,N_2172,N_2184);
or U2221 (N_2221,N_2163,N_2175);
and U2222 (N_2222,N_2208,N_2201);
nor U2223 (N_2223,N_2178,N_2194);
and U2224 (N_2224,N_2162,N_2204);
or U2225 (N_2225,N_2215,N_2193);
or U2226 (N_2226,N_2190,N_2214);
nor U2227 (N_2227,N_2164,N_2197);
and U2228 (N_2228,N_2181,N_2199);
nor U2229 (N_2229,N_2174,N_2182);
or U2230 (N_2230,N_2173,N_2196);
nor U2231 (N_2231,N_2216,N_2189);
or U2232 (N_2232,N_2192,N_2212);
and U2233 (N_2233,N_2177,N_2179);
and U2234 (N_2234,N_2191,N_2202);
nor U2235 (N_2235,N_2183,N_2167);
nor U2236 (N_2236,N_2219,N_2170);
and U2237 (N_2237,N_2217,N_2188);
nand U2238 (N_2238,N_2166,N_2198);
and U2239 (N_2239,N_2165,N_2160);
xnor U2240 (N_2240,N_2213,N_2168);
nor U2241 (N_2241,N_2206,N_2211);
or U2242 (N_2242,N_2185,N_2207);
nor U2243 (N_2243,N_2203,N_2171);
nand U2244 (N_2244,N_2195,N_2209);
and U2245 (N_2245,N_2186,N_2180);
and U2246 (N_2246,N_2205,N_2169);
or U2247 (N_2247,N_2161,N_2187);
and U2248 (N_2248,N_2176,N_2210);
nand U2249 (N_2249,N_2200,N_2218);
and U2250 (N_2250,N_2213,N_2210);
and U2251 (N_2251,N_2215,N_2205);
and U2252 (N_2252,N_2194,N_2204);
and U2253 (N_2253,N_2179,N_2192);
nand U2254 (N_2254,N_2178,N_2176);
nor U2255 (N_2255,N_2218,N_2188);
and U2256 (N_2256,N_2188,N_2161);
and U2257 (N_2257,N_2174,N_2192);
and U2258 (N_2258,N_2212,N_2174);
and U2259 (N_2259,N_2218,N_2210);
nor U2260 (N_2260,N_2188,N_2213);
or U2261 (N_2261,N_2167,N_2201);
nor U2262 (N_2262,N_2202,N_2196);
or U2263 (N_2263,N_2181,N_2215);
and U2264 (N_2264,N_2193,N_2182);
or U2265 (N_2265,N_2182,N_2192);
and U2266 (N_2266,N_2218,N_2174);
nor U2267 (N_2267,N_2197,N_2172);
nor U2268 (N_2268,N_2206,N_2185);
xnor U2269 (N_2269,N_2211,N_2162);
or U2270 (N_2270,N_2177,N_2187);
nand U2271 (N_2271,N_2161,N_2183);
nand U2272 (N_2272,N_2218,N_2184);
nor U2273 (N_2273,N_2217,N_2176);
nand U2274 (N_2274,N_2166,N_2171);
or U2275 (N_2275,N_2201,N_2213);
nor U2276 (N_2276,N_2186,N_2161);
or U2277 (N_2277,N_2205,N_2176);
and U2278 (N_2278,N_2181,N_2217);
nor U2279 (N_2279,N_2215,N_2174);
and U2280 (N_2280,N_2247,N_2250);
and U2281 (N_2281,N_2221,N_2244);
nor U2282 (N_2282,N_2245,N_2269);
nor U2283 (N_2283,N_2236,N_2252);
nand U2284 (N_2284,N_2253,N_2265);
nor U2285 (N_2285,N_2274,N_2273);
or U2286 (N_2286,N_2224,N_2268);
nor U2287 (N_2287,N_2223,N_2238);
nand U2288 (N_2288,N_2260,N_2271);
nor U2289 (N_2289,N_2258,N_2241);
nor U2290 (N_2290,N_2266,N_2228);
nor U2291 (N_2291,N_2225,N_2233);
nand U2292 (N_2292,N_2270,N_2279);
or U2293 (N_2293,N_2259,N_2226);
and U2294 (N_2294,N_2255,N_2276);
nor U2295 (N_2295,N_2264,N_2277);
or U2296 (N_2296,N_2262,N_2248);
nand U2297 (N_2297,N_2240,N_2275);
or U2298 (N_2298,N_2222,N_2235);
nor U2299 (N_2299,N_2239,N_2254);
or U2300 (N_2300,N_2227,N_2232);
nor U2301 (N_2301,N_2256,N_2242);
or U2302 (N_2302,N_2267,N_2272);
nand U2303 (N_2303,N_2261,N_2237);
nor U2304 (N_2304,N_2243,N_2246);
nand U2305 (N_2305,N_2229,N_2231);
or U2306 (N_2306,N_2257,N_2278);
nand U2307 (N_2307,N_2251,N_2220);
and U2308 (N_2308,N_2230,N_2249);
and U2309 (N_2309,N_2263,N_2234);
and U2310 (N_2310,N_2220,N_2246);
nand U2311 (N_2311,N_2262,N_2259);
and U2312 (N_2312,N_2269,N_2277);
and U2313 (N_2313,N_2274,N_2227);
or U2314 (N_2314,N_2267,N_2259);
nand U2315 (N_2315,N_2220,N_2279);
and U2316 (N_2316,N_2250,N_2234);
or U2317 (N_2317,N_2279,N_2246);
nand U2318 (N_2318,N_2272,N_2220);
or U2319 (N_2319,N_2250,N_2256);
nor U2320 (N_2320,N_2245,N_2264);
and U2321 (N_2321,N_2266,N_2229);
nor U2322 (N_2322,N_2239,N_2234);
nand U2323 (N_2323,N_2230,N_2220);
nor U2324 (N_2324,N_2253,N_2261);
and U2325 (N_2325,N_2244,N_2279);
or U2326 (N_2326,N_2253,N_2220);
or U2327 (N_2327,N_2245,N_2250);
or U2328 (N_2328,N_2263,N_2271);
nor U2329 (N_2329,N_2246,N_2221);
nand U2330 (N_2330,N_2258,N_2231);
or U2331 (N_2331,N_2230,N_2245);
or U2332 (N_2332,N_2246,N_2258);
nor U2333 (N_2333,N_2249,N_2246);
nor U2334 (N_2334,N_2264,N_2224);
and U2335 (N_2335,N_2274,N_2272);
nor U2336 (N_2336,N_2235,N_2249);
nand U2337 (N_2337,N_2251,N_2226);
nor U2338 (N_2338,N_2254,N_2268);
or U2339 (N_2339,N_2224,N_2220);
nor U2340 (N_2340,N_2292,N_2283);
nor U2341 (N_2341,N_2321,N_2324);
nor U2342 (N_2342,N_2290,N_2334);
nand U2343 (N_2343,N_2286,N_2301);
or U2344 (N_2344,N_2287,N_2282);
nor U2345 (N_2345,N_2300,N_2288);
and U2346 (N_2346,N_2338,N_2323);
nand U2347 (N_2347,N_2336,N_2305);
and U2348 (N_2348,N_2337,N_2308);
nor U2349 (N_2349,N_2326,N_2296);
or U2350 (N_2350,N_2328,N_2293);
or U2351 (N_2351,N_2318,N_2291);
or U2352 (N_2352,N_2317,N_2325);
or U2353 (N_2353,N_2322,N_2284);
nor U2354 (N_2354,N_2299,N_2297);
nand U2355 (N_2355,N_2302,N_2294);
and U2356 (N_2356,N_2289,N_2309);
nor U2357 (N_2357,N_2319,N_2330);
and U2358 (N_2358,N_2320,N_2313);
nor U2359 (N_2359,N_2331,N_2307);
nor U2360 (N_2360,N_2281,N_2306);
nand U2361 (N_2361,N_2315,N_2304);
or U2362 (N_2362,N_2335,N_2312);
and U2363 (N_2363,N_2332,N_2327);
or U2364 (N_2364,N_2333,N_2280);
nand U2365 (N_2365,N_2285,N_2311);
or U2366 (N_2366,N_2298,N_2295);
nand U2367 (N_2367,N_2329,N_2310);
xor U2368 (N_2368,N_2303,N_2314);
nor U2369 (N_2369,N_2339,N_2316);
nor U2370 (N_2370,N_2336,N_2283);
and U2371 (N_2371,N_2301,N_2285);
and U2372 (N_2372,N_2282,N_2311);
nor U2373 (N_2373,N_2298,N_2292);
and U2374 (N_2374,N_2308,N_2327);
nand U2375 (N_2375,N_2291,N_2334);
nor U2376 (N_2376,N_2336,N_2299);
or U2377 (N_2377,N_2285,N_2297);
and U2378 (N_2378,N_2332,N_2313);
nand U2379 (N_2379,N_2288,N_2298);
nor U2380 (N_2380,N_2336,N_2317);
nand U2381 (N_2381,N_2323,N_2298);
or U2382 (N_2382,N_2327,N_2319);
nand U2383 (N_2383,N_2326,N_2299);
nand U2384 (N_2384,N_2280,N_2320);
or U2385 (N_2385,N_2338,N_2293);
and U2386 (N_2386,N_2282,N_2293);
or U2387 (N_2387,N_2332,N_2284);
nor U2388 (N_2388,N_2297,N_2332);
nor U2389 (N_2389,N_2303,N_2291);
nand U2390 (N_2390,N_2338,N_2321);
nand U2391 (N_2391,N_2312,N_2289);
and U2392 (N_2392,N_2283,N_2301);
or U2393 (N_2393,N_2335,N_2282);
nor U2394 (N_2394,N_2332,N_2316);
or U2395 (N_2395,N_2297,N_2316);
nand U2396 (N_2396,N_2315,N_2326);
and U2397 (N_2397,N_2320,N_2304);
nor U2398 (N_2398,N_2328,N_2332);
or U2399 (N_2399,N_2289,N_2294);
nand U2400 (N_2400,N_2360,N_2347);
and U2401 (N_2401,N_2385,N_2383);
nand U2402 (N_2402,N_2378,N_2389);
nor U2403 (N_2403,N_2364,N_2371);
or U2404 (N_2404,N_2367,N_2393);
nand U2405 (N_2405,N_2386,N_2399);
or U2406 (N_2406,N_2398,N_2397);
nand U2407 (N_2407,N_2354,N_2340);
nor U2408 (N_2408,N_2372,N_2350);
nand U2409 (N_2409,N_2362,N_2343);
or U2410 (N_2410,N_2377,N_2363);
nor U2411 (N_2411,N_2352,N_2342);
nor U2412 (N_2412,N_2341,N_2387);
nand U2413 (N_2413,N_2382,N_2388);
and U2414 (N_2414,N_2353,N_2368);
or U2415 (N_2415,N_2370,N_2379);
or U2416 (N_2416,N_2355,N_2348);
nor U2417 (N_2417,N_2380,N_2366);
nor U2418 (N_2418,N_2365,N_2395);
or U2419 (N_2419,N_2394,N_2381);
nor U2420 (N_2420,N_2361,N_2359);
and U2421 (N_2421,N_2376,N_2373);
nand U2422 (N_2422,N_2396,N_2356);
or U2423 (N_2423,N_2384,N_2391);
or U2424 (N_2424,N_2392,N_2358);
nor U2425 (N_2425,N_2357,N_2390);
nor U2426 (N_2426,N_2349,N_2375);
and U2427 (N_2427,N_2346,N_2344);
and U2428 (N_2428,N_2374,N_2345);
or U2429 (N_2429,N_2351,N_2369);
nor U2430 (N_2430,N_2357,N_2362);
and U2431 (N_2431,N_2356,N_2366);
or U2432 (N_2432,N_2389,N_2341);
or U2433 (N_2433,N_2373,N_2389);
nor U2434 (N_2434,N_2358,N_2364);
and U2435 (N_2435,N_2340,N_2356);
nand U2436 (N_2436,N_2383,N_2369);
nand U2437 (N_2437,N_2384,N_2370);
or U2438 (N_2438,N_2392,N_2394);
and U2439 (N_2439,N_2343,N_2387);
nor U2440 (N_2440,N_2359,N_2392);
and U2441 (N_2441,N_2365,N_2347);
or U2442 (N_2442,N_2370,N_2385);
nor U2443 (N_2443,N_2383,N_2368);
xor U2444 (N_2444,N_2365,N_2370);
nand U2445 (N_2445,N_2363,N_2399);
nor U2446 (N_2446,N_2396,N_2378);
nand U2447 (N_2447,N_2363,N_2369);
and U2448 (N_2448,N_2363,N_2371);
nor U2449 (N_2449,N_2362,N_2356);
nor U2450 (N_2450,N_2378,N_2379);
or U2451 (N_2451,N_2387,N_2360);
nor U2452 (N_2452,N_2366,N_2376);
or U2453 (N_2453,N_2395,N_2360);
nand U2454 (N_2454,N_2380,N_2393);
or U2455 (N_2455,N_2382,N_2380);
and U2456 (N_2456,N_2382,N_2356);
or U2457 (N_2457,N_2360,N_2370);
nor U2458 (N_2458,N_2357,N_2346);
nor U2459 (N_2459,N_2369,N_2387);
or U2460 (N_2460,N_2436,N_2401);
nand U2461 (N_2461,N_2438,N_2406);
and U2462 (N_2462,N_2452,N_2433);
nand U2463 (N_2463,N_2430,N_2448);
and U2464 (N_2464,N_2421,N_2420);
nand U2465 (N_2465,N_2423,N_2447);
or U2466 (N_2466,N_2437,N_2409);
and U2467 (N_2467,N_2427,N_2455);
and U2468 (N_2468,N_2419,N_2414);
nand U2469 (N_2469,N_2454,N_2458);
nor U2470 (N_2470,N_2413,N_2429);
and U2471 (N_2471,N_2416,N_2435);
nor U2472 (N_2472,N_2442,N_2418);
and U2473 (N_2473,N_2411,N_2431);
nor U2474 (N_2474,N_2417,N_2441);
xor U2475 (N_2475,N_2426,N_2456);
or U2476 (N_2476,N_2434,N_2453);
and U2477 (N_2477,N_2439,N_2443);
nand U2478 (N_2478,N_2405,N_2459);
or U2479 (N_2479,N_2408,N_2407);
or U2480 (N_2480,N_2404,N_2422);
nand U2481 (N_2481,N_2432,N_2400);
nor U2482 (N_2482,N_2450,N_2428);
nand U2483 (N_2483,N_2410,N_2451);
nand U2484 (N_2484,N_2415,N_2425);
or U2485 (N_2485,N_2446,N_2412);
and U2486 (N_2486,N_2445,N_2444);
nor U2487 (N_2487,N_2457,N_2402);
nand U2488 (N_2488,N_2449,N_2403);
nor U2489 (N_2489,N_2440,N_2424);
and U2490 (N_2490,N_2425,N_2447);
nor U2491 (N_2491,N_2436,N_2408);
nand U2492 (N_2492,N_2451,N_2401);
or U2493 (N_2493,N_2450,N_2425);
and U2494 (N_2494,N_2432,N_2412);
and U2495 (N_2495,N_2429,N_2418);
or U2496 (N_2496,N_2412,N_2444);
nor U2497 (N_2497,N_2455,N_2412);
nor U2498 (N_2498,N_2428,N_2439);
and U2499 (N_2499,N_2455,N_2429);
nand U2500 (N_2500,N_2416,N_2446);
or U2501 (N_2501,N_2404,N_2456);
nand U2502 (N_2502,N_2443,N_2418);
and U2503 (N_2503,N_2411,N_2426);
nand U2504 (N_2504,N_2428,N_2458);
and U2505 (N_2505,N_2445,N_2450);
nand U2506 (N_2506,N_2421,N_2450);
nand U2507 (N_2507,N_2457,N_2423);
nand U2508 (N_2508,N_2436,N_2432);
and U2509 (N_2509,N_2418,N_2445);
nor U2510 (N_2510,N_2418,N_2420);
or U2511 (N_2511,N_2415,N_2431);
nor U2512 (N_2512,N_2457,N_2411);
or U2513 (N_2513,N_2407,N_2414);
and U2514 (N_2514,N_2434,N_2411);
nor U2515 (N_2515,N_2420,N_2410);
nor U2516 (N_2516,N_2414,N_2444);
nand U2517 (N_2517,N_2421,N_2422);
nand U2518 (N_2518,N_2406,N_2403);
nand U2519 (N_2519,N_2406,N_2408);
xor U2520 (N_2520,N_2517,N_2487);
and U2521 (N_2521,N_2475,N_2518);
nor U2522 (N_2522,N_2503,N_2462);
nor U2523 (N_2523,N_2498,N_2477);
or U2524 (N_2524,N_2497,N_2469);
nor U2525 (N_2525,N_2511,N_2467);
or U2526 (N_2526,N_2484,N_2508);
or U2527 (N_2527,N_2505,N_2483);
and U2528 (N_2528,N_2500,N_2479);
nor U2529 (N_2529,N_2465,N_2512);
nand U2530 (N_2530,N_2496,N_2472);
or U2531 (N_2531,N_2489,N_2506);
or U2532 (N_2532,N_2481,N_2485);
and U2533 (N_2533,N_2499,N_2492);
nand U2534 (N_2534,N_2510,N_2507);
and U2535 (N_2535,N_2471,N_2468);
nor U2536 (N_2536,N_2491,N_2474);
and U2537 (N_2537,N_2470,N_2478);
and U2538 (N_2538,N_2460,N_2488);
or U2539 (N_2539,N_2486,N_2495);
nand U2540 (N_2540,N_2501,N_2504);
nor U2541 (N_2541,N_2493,N_2494);
nor U2542 (N_2542,N_2473,N_2480);
and U2543 (N_2543,N_2516,N_2513);
and U2544 (N_2544,N_2476,N_2515);
or U2545 (N_2545,N_2463,N_2514);
or U2546 (N_2546,N_2490,N_2482);
nor U2547 (N_2547,N_2466,N_2519);
or U2548 (N_2548,N_2464,N_2502);
nand U2549 (N_2549,N_2461,N_2509);
nor U2550 (N_2550,N_2489,N_2497);
or U2551 (N_2551,N_2501,N_2486);
nand U2552 (N_2552,N_2494,N_2474);
and U2553 (N_2553,N_2461,N_2463);
and U2554 (N_2554,N_2464,N_2461);
xor U2555 (N_2555,N_2500,N_2461);
nand U2556 (N_2556,N_2496,N_2518);
or U2557 (N_2557,N_2487,N_2488);
nand U2558 (N_2558,N_2509,N_2465);
nor U2559 (N_2559,N_2488,N_2508);
nand U2560 (N_2560,N_2497,N_2467);
nand U2561 (N_2561,N_2478,N_2493);
and U2562 (N_2562,N_2467,N_2474);
nor U2563 (N_2563,N_2512,N_2506);
and U2564 (N_2564,N_2500,N_2510);
and U2565 (N_2565,N_2502,N_2496);
nor U2566 (N_2566,N_2469,N_2491);
and U2567 (N_2567,N_2466,N_2500);
nor U2568 (N_2568,N_2500,N_2512);
and U2569 (N_2569,N_2518,N_2485);
or U2570 (N_2570,N_2480,N_2488);
nor U2571 (N_2571,N_2488,N_2510);
or U2572 (N_2572,N_2462,N_2490);
or U2573 (N_2573,N_2499,N_2467);
nand U2574 (N_2574,N_2511,N_2514);
or U2575 (N_2575,N_2475,N_2461);
nand U2576 (N_2576,N_2497,N_2460);
and U2577 (N_2577,N_2497,N_2506);
nor U2578 (N_2578,N_2491,N_2481);
nand U2579 (N_2579,N_2514,N_2492);
or U2580 (N_2580,N_2572,N_2533);
nor U2581 (N_2581,N_2544,N_2555);
nor U2582 (N_2582,N_2570,N_2547);
or U2583 (N_2583,N_2545,N_2569);
nor U2584 (N_2584,N_2556,N_2577);
xor U2585 (N_2585,N_2534,N_2575);
or U2586 (N_2586,N_2562,N_2537);
or U2587 (N_2587,N_2531,N_2530);
nand U2588 (N_2588,N_2558,N_2520);
nand U2589 (N_2589,N_2538,N_2535);
or U2590 (N_2590,N_2554,N_2543);
or U2591 (N_2591,N_2529,N_2527);
nand U2592 (N_2592,N_2561,N_2523);
nor U2593 (N_2593,N_2563,N_2576);
nor U2594 (N_2594,N_2548,N_2566);
nor U2595 (N_2595,N_2542,N_2578);
and U2596 (N_2596,N_2564,N_2568);
and U2597 (N_2597,N_2553,N_2571);
nand U2598 (N_2598,N_2525,N_2551);
nand U2599 (N_2599,N_2573,N_2557);
and U2600 (N_2600,N_2579,N_2567);
or U2601 (N_2601,N_2574,N_2539);
nand U2602 (N_2602,N_2536,N_2549);
nor U2603 (N_2603,N_2552,N_2532);
nor U2604 (N_2604,N_2526,N_2541);
and U2605 (N_2605,N_2546,N_2560);
nand U2606 (N_2606,N_2550,N_2522);
or U2607 (N_2607,N_2521,N_2565);
and U2608 (N_2608,N_2540,N_2528);
or U2609 (N_2609,N_2524,N_2559);
nand U2610 (N_2610,N_2561,N_2534);
and U2611 (N_2611,N_2573,N_2534);
nand U2612 (N_2612,N_2551,N_2534);
or U2613 (N_2613,N_2520,N_2571);
nor U2614 (N_2614,N_2547,N_2521);
nand U2615 (N_2615,N_2540,N_2541);
and U2616 (N_2616,N_2561,N_2555);
or U2617 (N_2617,N_2525,N_2556);
nand U2618 (N_2618,N_2552,N_2554);
nand U2619 (N_2619,N_2529,N_2558);
nand U2620 (N_2620,N_2521,N_2555);
nand U2621 (N_2621,N_2545,N_2579);
xor U2622 (N_2622,N_2575,N_2541);
nand U2623 (N_2623,N_2550,N_2538);
nor U2624 (N_2624,N_2546,N_2548);
nor U2625 (N_2625,N_2557,N_2578);
nand U2626 (N_2626,N_2558,N_2566);
and U2627 (N_2627,N_2538,N_2522);
nor U2628 (N_2628,N_2569,N_2562);
nand U2629 (N_2629,N_2567,N_2572);
xnor U2630 (N_2630,N_2555,N_2569);
and U2631 (N_2631,N_2563,N_2557);
nand U2632 (N_2632,N_2556,N_2575);
and U2633 (N_2633,N_2546,N_2574);
and U2634 (N_2634,N_2562,N_2531);
nor U2635 (N_2635,N_2544,N_2533);
and U2636 (N_2636,N_2541,N_2548);
and U2637 (N_2637,N_2574,N_2536);
nand U2638 (N_2638,N_2528,N_2568);
and U2639 (N_2639,N_2532,N_2554);
nand U2640 (N_2640,N_2605,N_2615);
nor U2641 (N_2641,N_2597,N_2634);
nor U2642 (N_2642,N_2600,N_2580);
nand U2643 (N_2643,N_2619,N_2636);
or U2644 (N_2644,N_2626,N_2593);
or U2645 (N_2645,N_2627,N_2628);
nand U2646 (N_2646,N_2630,N_2604);
or U2647 (N_2647,N_2603,N_2638);
or U2648 (N_2648,N_2620,N_2583);
nand U2649 (N_2649,N_2629,N_2595);
nor U2650 (N_2650,N_2581,N_2588);
nand U2651 (N_2651,N_2598,N_2606);
nor U2652 (N_2652,N_2635,N_2594);
nand U2653 (N_2653,N_2612,N_2609);
or U2654 (N_2654,N_2616,N_2632);
nand U2655 (N_2655,N_2624,N_2599);
and U2656 (N_2656,N_2622,N_2585);
nor U2657 (N_2657,N_2607,N_2623);
and U2658 (N_2658,N_2592,N_2611);
and U2659 (N_2659,N_2617,N_2590);
nor U2660 (N_2660,N_2621,N_2582);
xor U2661 (N_2661,N_2591,N_2596);
and U2662 (N_2662,N_2584,N_2586);
nand U2663 (N_2663,N_2601,N_2614);
nor U2664 (N_2664,N_2610,N_2631);
nand U2665 (N_2665,N_2587,N_2637);
nor U2666 (N_2666,N_2589,N_2625);
or U2667 (N_2667,N_2602,N_2613);
or U2668 (N_2668,N_2633,N_2639);
and U2669 (N_2669,N_2608,N_2618);
nor U2670 (N_2670,N_2632,N_2592);
nor U2671 (N_2671,N_2626,N_2592);
xnor U2672 (N_2672,N_2635,N_2582);
nor U2673 (N_2673,N_2607,N_2589);
and U2674 (N_2674,N_2592,N_2610);
nor U2675 (N_2675,N_2633,N_2605);
nor U2676 (N_2676,N_2638,N_2592);
nand U2677 (N_2677,N_2602,N_2587);
and U2678 (N_2678,N_2614,N_2586);
and U2679 (N_2679,N_2626,N_2632);
nor U2680 (N_2680,N_2606,N_2592);
nor U2681 (N_2681,N_2585,N_2633);
nor U2682 (N_2682,N_2634,N_2584);
nand U2683 (N_2683,N_2597,N_2613);
or U2684 (N_2684,N_2629,N_2623);
nand U2685 (N_2685,N_2630,N_2590);
nand U2686 (N_2686,N_2636,N_2614);
nand U2687 (N_2687,N_2631,N_2634);
or U2688 (N_2688,N_2605,N_2586);
and U2689 (N_2689,N_2586,N_2630);
nand U2690 (N_2690,N_2623,N_2580);
nand U2691 (N_2691,N_2622,N_2589);
and U2692 (N_2692,N_2636,N_2615);
xor U2693 (N_2693,N_2627,N_2630);
nor U2694 (N_2694,N_2632,N_2607);
nand U2695 (N_2695,N_2621,N_2622);
or U2696 (N_2696,N_2617,N_2639);
or U2697 (N_2697,N_2602,N_2607);
nand U2698 (N_2698,N_2620,N_2592);
nor U2699 (N_2699,N_2590,N_2616);
and U2700 (N_2700,N_2657,N_2665);
or U2701 (N_2701,N_2642,N_2643);
and U2702 (N_2702,N_2645,N_2663);
or U2703 (N_2703,N_2678,N_2644);
and U2704 (N_2704,N_2694,N_2697);
or U2705 (N_2705,N_2660,N_2688);
nor U2706 (N_2706,N_2653,N_2681);
and U2707 (N_2707,N_2683,N_2649);
and U2708 (N_2708,N_2671,N_2661);
and U2709 (N_2709,N_2680,N_2658);
and U2710 (N_2710,N_2652,N_2648);
nand U2711 (N_2711,N_2667,N_2654);
xnor U2712 (N_2712,N_2672,N_2679);
or U2713 (N_2713,N_2695,N_2677);
or U2714 (N_2714,N_2662,N_2673);
or U2715 (N_2715,N_2696,N_2698);
and U2716 (N_2716,N_2685,N_2666);
and U2717 (N_2717,N_2651,N_2676);
or U2718 (N_2718,N_2670,N_2690);
nand U2719 (N_2719,N_2641,N_2656);
nand U2720 (N_2720,N_2693,N_2686);
nand U2721 (N_2721,N_2689,N_2664);
nand U2722 (N_2722,N_2650,N_2640);
xor U2723 (N_2723,N_2699,N_2675);
nor U2724 (N_2724,N_2668,N_2692);
nand U2725 (N_2725,N_2659,N_2687);
or U2726 (N_2726,N_2647,N_2646);
nand U2727 (N_2727,N_2669,N_2674);
nand U2728 (N_2728,N_2691,N_2684);
or U2729 (N_2729,N_2682,N_2655);
and U2730 (N_2730,N_2643,N_2681);
nor U2731 (N_2731,N_2691,N_2688);
and U2732 (N_2732,N_2658,N_2687);
and U2733 (N_2733,N_2687,N_2696);
and U2734 (N_2734,N_2689,N_2651);
or U2735 (N_2735,N_2653,N_2669);
nor U2736 (N_2736,N_2672,N_2683);
or U2737 (N_2737,N_2681,N_2668);
nor U2738 (N_2738,N_2689,N_2643);
nand U2739 (N_2739,N_2668,N_2697);
and U2740 (N_2740,N_2671,N_2676);
nor U2741 (N_2741,N_2644,N_2692);
and U2742 (N_2742,N_2644,N_2654);
nor U2743 (N_2743,N_2668,N_2686);
nor U2744 (N_2744,N_2660,N_2681);
or U2745 (N_2745,N_2670,N_2686);
and U2746 (N_2746,N_2676,N_2679);
nor U2747 (N_2747,N_2664,N_2668);
and U2748 (N_2748,N_2654,N_2663);
and U2749 (N_2749,N_2657,N_2695);
and U2750 (N_2750,N_2665,N_2666);
and U2751 (N_2751,N_2665,N_2689);
nor U2752 (N_2752,N_2668,N_2688);
and U2753 (N_2753,N_2661,N_2665);
and U2754 (N_2754,N_2661,N_2693);
and U2755 (N_2755,N_2690,N_2656);
or U2756 (N_2756,N_2643,N_2680);
and U2757 (N_2757,N_2655,N_2693);
and U2758 (N_2758,N_2692,N_2699);
or U2759 (N_2759,N_2642,N_2679);
nor U2760 (N_2760,N_2738,N_2704);
nor U2761 (N_2761,N_2718,N_2700);
and U2762 (N_2762,N_2729,N_2746);
and U2763 (N_2763,N_2701,N_2748);
and U2764 (N_2764,N_2706,N_2745);
nor U2765 (N_2765,N_2740,N_2717);
or U2766 (N_2766,N_2741,N_2758);
or U2767 (N_2767,N_2742,N_2719);
and U2768 (N_2768,N_2713,N_2733);
nor U2769 (N_2769,N_2727,N_2725);
nand U2770 (N_2770,N_2723,N_2722);
and U2771 (N_2771,N_2721,N_2759);
or U2772 (N_2772,N_2737,N_2724);
and U2773 (N_2773,N_2711,N_2712);
or U2774 (N_2774,N_2732,N_2730);
and U2775 (N_2775,N_2747,N_2710);
or U2776 (N_2776,N_2750,N_2754);
nand U2777 (N_2777,N_2702,N_2720);
xor U2778 (N_2778,N_2715,N_2749);
or U2779 (N_2779,N_2707,N_2752);
nand U2780 (N_2780,N_2751,N_2735);
and U2781 (N_2781,N_2716,N_2756);
nand U2782 (N_2782,N_2709,N_2708);
or U2783 (N_2783,N_2755,N_2726);
or U2784 (N_2784,N_2753,N_2734);
nand U2785 (N_2785,N_2757,N_2705);
or U2786 (N_2786,N_2744,N_2743);
or U2787 (N_2787,N_2728,N_2714);
and U2788 (N_2788,N_2736,N_2731);
nand U2789 (N_2789,N_2703,N_2739);
and U2790 (N_2790,N_2759,N_2747);
nor U2791 (N_2791,N_2730,N_2706);
or U2792 (N_2792,N_2748,N_2728);
or U2793 (N_2793,N_2726,N_2746);
or U2794 (N_2794,N_2707,N_2745);
and U2795 (N_2795,N_2743,N_2729);
nand U2796 (N_2796,N_2710,N_2707);
and U2797 (N_2797,N_2706,N_2754);
nand U2798 (N_2798,N_2754,N_2743);
or U2799 (N_2799,N_2751,N_2748);
nor U2800 (N_2800,N_2724,N_2741);
or U2801 (N_2801,N_2751,N_2754);
and U2802 (N_2802,N_2759,N_2723);
nor U2803 (N_2803,N_2758,N_2713);
and U2804 (N_2804,N_2759,N_2751);
or U2805 (N_2805,N_2747,N_2703);
nor U2806 (N_2806,N_2722,N_2710);
and U2807 (N_2807,N_2747,N_2756);
nand U2808 (N_2808,N_2707,N_2738);
and U2809 (N_2809,N_2721,N_2716);
nor U2810 (N_2810,N_2705,N_2736);
and U2811 (N_2811,N_2737,N_2708);
and U2812 (N_2812,N_2703,N_2700);
nor U2813 (N_2813,N_2728,N_2758);
nand U2814 (N_2814,N_2714,N_2751);
or U2815 (N_2815,N_2713,N_2711);
and U2816 (N_2816,N_2716,N_2745);
nor U2817 (N_2817,N_2743,N_2739);
nor U2818 (N_2818,N_2732,N_2750);
xnor U2819 (N_2819,N_2714,N_2729);
nand U2820 (N_2820,N_2788,N_2809);
and U2821 (N_2821,N_2764,N_2813);
or U2822 (N_2822,N_2789,N_2811);
or U2823 (N_2823,N_2778,N_2795);
or U2824 (N_2824,N_2782,N_2793);
and U2825 (N_2825,N_2763,N_2803);
nor U2826 (N_2826,N_2779,N_2799);
nand U2827 (N_2827,N_2765,N_2781);
nor U2828 (N_2828,N_2819,N_2770);
or U2829 (N_2829,N_2807,N_2776);
or U2830 (N_2830,N_2797,N_2780);
or U2831 (N_2831,N_2818,N_2766);
and U2832 (N_2832,N_2810,N_2798);
nor U2833 (N_2833,N_2773,N_2787);
nor U2834 (N_2834,N_2815,N_2804);
nand U2835 (N_2835,N_2768,N_2805);
nor U2836 (N_2836,N_2777,N_2784);
nor U2837 (N_2837,N_2808,N_2801);
nand U2838 (N_2838,N_2800,N_2760);
and U2839 (N_2839,N_2812,N_2771);
or U2840 (N_2840,N_2761,N_2796);
nor U2841 (N_2841,N_2775,N_2785);
or U2842 (N_2842,N_2786,N_2792);
nand U2843 (N_2843,N_2816,N_2767);
nand U2844 (N_2844,N_2806,N_2772);
nor U2845 (N_2845,N_2790,N_2817);
nand U2846 (N_2846,N_2783,N_2769);
and U2847 (N_2847,N_2791,N_2762);
nand U2848 (N_2848,N_2802,N_2794);
nor U2849 (N_2849,N_2774,N_2814);
nand U2850 (N_2850,N_2768,N_2761);
and U2851 (N_2851,N_2791,N_2778);
and U2852 (N_2852,N_2764,N_2761);
nor U2853 (N_2853,N_2777,N_2776);
and U2854 (N_2854,N_2804,N_2791);
nand U2855 (N_2855,N_2791,N_2783);
or U2856 (N_2856,N_2768,N_2787);
xnor U2857 (N_2857,N_2814,N_2782);
or U2858 (N_2858,N_2771,N_2776);
nand U2859 (N_2859,N_2771,N_2783);
nor U2860 (N_2860,N_2770,N_2784);
nand U2861 (N_2861,N_2797,N_2798);
nor U2862 (N_2862,N_2810,N_2801);
nand U2863 (N_2863,N_2790,N_2803);
or U2864 (N_2864,N_2811,N_2799);
nor U2865 (N_2865,N_2765,N_2782);
nor U2866 (N_2866,N_2808,N_2803);
nand U2867 (N_2867,N_2806,N_2768);
and U2868 (N_2868,N_2767,N_2804);
or U2869 (N_2869,N_2794,N_2813);
or U2870 (N_2870,N_2794,N_2782);
nor U2871 (N_2871,N_2761,N_2770);
xor U2872 (N_2872,N_2791,N_2802);
nor U2873 (N_2873,N_2766,N_2772);
and U2874 (N_2874,N_2787,N_2789);
nor U2875 (N_2875,N_2788,N_2771);
nand U2876 (N_2876,N_2812,N_2789);
nor U2877 (N_2877,N_2793,N_2817);
xnor U2878 (N_2878,N_2808,N_2800);
nand U2879 (N_2879,N_2813,N_2795);
and U2880 (N_2880,N_2875,N_2830);
nor U2881 (N_2881,N_2849,N_2874);
nor U2882 (N_2882,N_2857,N_2862);
or U2883 (N_2883,N_2867,N_2828);
or U2884 (N_2884,N_2823,N_2853);
nand U2885 (N_2885,N_2842,N_2822);
nor U2886 (N_2886,N_2858,N_2824);
nor U2887 (N_2887,N_2868,N_2865);
nand U2888 (N_2888,N_2860,N_2847);
nor U2889 (N_2889,N_2854,N_2852);
nand U2890 (N_2890,N_2846,N_2851);
nand U2891 (N_2891,N_2826,N_2859);
nand U2892 (N_2892,N_2873,N_2864);
nor U2893 (N_2893,N_2877,N_2821);
nor U2894 (N_2894,N_2856,N_2871);
and U2895 (N_2895,N_2840,N_2835);
nor U2896 (N_2896,N_2827,N_2869);
nand U2897 (N_2897,N_2837,N_2855);
nand U2898 (N_2898,N_2845,N_2825);
or U2899 (N_2899,N_2844,N_2850);
nand U2900 (N_2900,N_2829,N_2872);
nand U2901 (N_2901,N_2870,N_2841);
nor U2902 (N_2902,N_2836,N_2838);
nand U2903 (N_2903,N_2831,N_2863);
nand U2904 (N_2904,N_2876,N_2820);
and U2905 (N_2905,N_2839,N_2848);
and U2906 (N_2906,N_2879,N_2833);
or U2907 (N_2907,N_2832,N_2866);
nand U2908 (N_2908,N_2843,N_2861);
and U2909 (N_2909,N_2834,N_2878);
nor U2910 (N_2910,N_2856,N_2863);
nor U2911 (N_2911,N_2845,N_2851);
or U2912 (N_2912,N_2856,N_2875);
nand U2913 (N_2913,N_2867,N_2830);
nor U2914 (N_2914,N_2820,N_2826);
and U2915 (N_2915,N_2869,N_2839);
or U2916 (N_2916,N_2835,N_2822);
or U2917 (N_2917,N_2848,N_2856);
nor U2918 (N_2918,N_2879,N_2874);
nand U2919 (N_2919,N_2833,N_2851);
nor U2920 (N_2920,N_2870,N_2848);
or U2921 (N_2921,N_2856,N_2829);
and U2922 (N_2922,N_2842,N_2825);
nand U2923 (N_2923,N_2852,N_2872);
nor U2924 (N_2924,N_2830,N_2825);
and U2925 (N_2925,N_2835,N_2827);
nand U2926 (N_2926,N_2875,N_2854);
nor U2927 (N_2927,N_2859,N_2838);
and U2928 (N_2928,N_2856,N_2835);
nor U2929 (N_2929,N_2867,N_2853);
or U2930 (N_2930,N_2849,N_2853);
or U2931 (N_2931,N_2847,N_2858);
nor U2932 (N_2932,N_2837,N_2844);
nand U2933 (N_2933,N_2857,N_2841);
nor U2934 (N_2934,N_2825,N_2876);
nor U2935 (N_2935,N_2823,N_2824);
and U2936 (N_2936,N_2877,N_2824);
or U2937 (N_2937,N_2821,N_2835);
or U2938 (N_2938,N_2869,N_2860);
nor U2939 (N_2939,N_2856,N_2851);
nor U2940 (N_2940,N_2887,N_2910);
nand U2941 (N_2941,N_2902,N_2907);
or U2942 (N_2942,N_2933,N_2886);
and U2943 (N_2943,N_2921,N_2911);
nor U2944 (N_2944,N_2930,N_2881);
nand U2945 (N_2945,N_2913,N_2920);
nor U2946 (N_2946,N_2939,N_2885);
nand U2947 (N_2947,N_2912,N_2891);
nor U2948 (N_2948,N_2928,N_2882);
and U2949 (N_2949,N_2927,N_2905);
and U2950 (N_2950,N_2892,N_2925);
or U2951 (N_2951,N_2918,N_2903);
or U2952 (N_2952,N_2896,N_2916);
or U2953 (N_2953,N_2924,N_2897);
nand U2954 (N_2954,N_2900,N_2936);
nand U2955 (N_2955,N_2934,N_2922);
or U2956 (N_2956,N_2938,N_2931);
and U2957 (N_2957,N_2909,N_2880);
or U2958 (N_2958,N_2889,N_2890);
and U2959 (N_2959,N_2895,N_2884);
or U2960 (N_2960,N_2898,N_2906);
nor U2961 (N_2961,N_2914,N_2904);
or U2962 (N_2962,N_2917,N_2901);
nor U2963 (N_2963,N_2888,N_2899);
xor U2964 (N_2964,N_2883,N_2908);
nand U2965 (N_2965,N_2937,N_2926);
nor U2966 (N_2966,N_2894,N_2929);
nor U2967 (N_2967,N_2932,N_2893);
nand U2968 (N_2968,N_2915,N_2923);
or U2969 (N_2969,N_2919,N_2935);
nand U2970 (N_2970,N_2915,N_2932);
nand U2971 (N_2971,N_2897,N_2889);
or U2972 (N_2972,N_2898,N_2932);
nor U2973 (N_2973,N_2912,N_2918);
or U2974 (N_2974,N_2934,N_2901);
nor U2975 (N_2975,N_2892,N_2880);
or U2976 (N_2976,N_2890,N_2909);
or U2977 (N_2977,N_2895,N_2883);
and U2978 (N_2978,N_2929,N_2928);
and U2979 (N_2979,N_2919,N_2896);
or U2980 (N_2980,N_2907,N_2900);
or U2981 (N_2981,N_2908,N_2891);
or U2982 (N_2982,N_2909,N_2881);
or U2983 (N_2983,N_2925,N_2904);
and U2984 (N_2984,N_2915,N_2899);
and U2985 (N_2985,N_2905,N_2901);
or U2986 (N_2986,N_2911,N_2885);
nand U2987 (N_2987,N_2905,N_2883);
and U2988 (N_2988,N_2907,N_2930);
nor U2989 (N_2989,N_2927,N_2929);
nand U2990 (N_2990,N_2907,N_2880);
and U2991 (N_2991,N_2888,N_2904);
or U2992 (N_2992,N_2895,N_2918);
nor U2993 (N_2993,N_2912,N_2911);
and U2994 (N_2994,N_2931,N_2898);
nor U2995 (N_2995,N_2883,N_2899);
and U2996 (N_2996,N_2911,N_2910);
and U2997 (N_2997,N_2916,N_2924);
nand U2998 (N_2998,N_2926,N_2912);
nand U2999 (N_2999,N_2888,N_2930);
or UO_0 (O_0,N_2995,N_2996);
and UO_1 (O_1,N_2954,N_2985);
and UO_2 (O_2,N_2951,N_2940);
or UO_3 (O_3,N_2957,N_2947);
and UO_4 (O_4,N_2946,N_2973);
nand UO_5 (O_5,N_2977,N_2961);
and UO_6 (O_6,N_2964,N_2943);
nor UO_7 (O_7,N_2994,N_2990);
nor UO_8 (O_8,N_2992,N_2980);
nand UO_9 (O_9,N_2959,N_2942);
nor UO_10 (O_10,N_2955,N_2952);
or UO_11 (O_11,N_2971,N_2944);
nand UO_12 (O_12,N_2989,N_2993);
or UO_13 (O_13,N_2982,N_2974);
nor UO_14 (O_14,N_2970,N_2963);
nor UO_15 (O_15,N_2962,N_2965);
nand UO_16 (O_16,N_2953,N_2967);
or UO_17 (O_17,N_2972,N_2986);
or UO_18 (O_18,N_2956,N_2968);
or UO_19 (O_19,N_2987,N_2978);
or UO_20 (O_20,N_2969,N_2966);
or UO_21 (O_21,N_2960,N_2975);
or UO_22 (O_22,N_2958,N_2991);
nand UO_23 (O_23,N_2979,N_2941);
or UO_24 (O_24,N_2997,N_2984);
nor UO_25 (O_25,N_2948,N_2999);
and UO_26 (O_26,N_2981,N_2949);
nor UO_27 (O_27,N_2976,N_2945);
nor UO_28 (O_28,N_2998,N_2983);
and UO_29 (O_29,N_2988,N_2950);
and UO_30 (O_30,N_2981,N_2950);
nand UO_31 (O_31,N_2961,N_2956);
nand UO_32 (O_32,N_2962,N_2990);
or UO_33 (O_33,N_2958,N_2951);
and UO_34 (O_34,N_2949,N_2966);
or UO_35 (O_35,N_2978,N_2945);
nand UO_36 (O_36,N_2977,N_2990);
nand UO_37 (O_37,N_2958,N_2956);
nor UO_38 (O_38,N_2971,N_2960);
or UO_39 (O_39,N_2978,N_2999);
or UO_40 (O_40,N_2944,N_2973);
or UO_41 (O_41,N_2992,N_2940);
nand UO_42 (O_42,N_2946,N_2996);
and UO_43 (O_43,N_2987,N_2942);
and UO_44 (O_44,N_2979,N_2969);
and UO_45 (O_45,N_2990,N_2981);
or UO_46 (O_46,N_2964,N_2952);
nor UO_47 (O_47,N_2955,N_2999);
or UO_48 (O_48,N_2949,N_2959);
or UO_49 (O_49,N_2973,N_2977);
and UO_50 (O_50,N_2943,N_2947);
and UO_51 (O_51,N_2956,N_2979);
or UO_52 (O_52,N_2968,N_2976);
and UO_53 (O_53,N_2980,N_2981);
and UO_54 (O_54,N_2944,N_2978);
nand UO_55 (O_55,N_2964,N_2953);
nor UO_56 (O_56,N_2980,N_2974);
nor UO_57 (O_57,N_2981,N_2996);
or UO_58 (O_58,N_2991,N_2981);
nand UO_59 (O_59,N_2956,N_2996);
or UO_60 (O_60,N_2950,N_2989);
nand UO_61 (O_61,N_2991,N_2943);
nand UO_62 (O_62,N_2954,N_2978);
nand UO_63 (O_63,N_2996,N_2976);
and UO_64 (O_64,N_2953,N_2975);
nand UO_65 (O_65,N_2960,N_2993);
or UO_66 (O_66,N_2997,N_2959);
nand UO_67 (O_67,N_2958,N_2973);
or UO_68 (O_68,N_2984,N_2975);
or UO_69 (O_69,N_2957,N_2982);
or UO_70 (O_70,N_2955,N_2975);
and UO_71 (O_71,N_2946,N_2998);
nand UO_72 (O_72,N_2970,N_2968);
nor UO_73 (O_73,N_2983,N_2972);
and UO_74 (O_74,N_2983,N_2976);
nor UO_75 (O_75,N_2940,N_2998);
nand UO_76 (O_76,N_2997,N_2967);
and UO_77 (O_77,N_2983,N_2940);
nor UO_78 (O_78,N_2959,N_2965);
and UO_79 (O_79,N_2949,N_2943);
and UO_80 (O_80,N_2962,N_2991);
nand UO_81 (O_81,N_2940,N_2997);
or UO_82 (O_82,N_2976,N_2985);
nand UO_83 (O_83,N_2976,N_2987);
and UO_84 (O_84,N_2948,N_2996);
nand UO_85 (O_85,N_2998,N_2994);
nand UO_86 (O_86,N_2977,N_2985);
or UO_87 (O_87,N_2945,N_2997);
nand UO_88 (O_88,N_2993,N_2962);
nor UO_89 (O_89,N_2943,N_2950);
nor UO_90 (O_90,N_2944,N_2992);
nor UO_91 (O_91,N_2987,N_2996);
nand UO_92 (O_92,N_2959,N_2976);
nor UO_93 (O_93,N_2980,N_2979);
and UO_94 (O_94,N_2944,N_2946);
and UO_95 (O_95,N_2974,N_2978);
nor UO_96 (O_96,N_2940,N_2944);
and UO_97 (O_97,N_2945,N_2946);
xnor UO_98 (O_98,N_2990,N_2970);
and UO_99 (O_99,N_2966,N_2956);
nor UO_100 (O_100,N_2946,N_2986);
nor UO_101 (O_101,N_2976,N_2989);
or UO_102 (O_102,N_2972,N_2950);
or UO_103 (O_103,N_2966,N_2974);
and UO_104 (O_104,N_2949,N_2951);
or UO_105 (O_105,N_2988,N_2987);
nand UO_106 (O_106,N_2995,N_2946);
or UO_107 (O_107,N_2958,N_2960);
and UO_108 (O_108,N_2955,N_2949);
nand UO_109 (O_109,N_2997,N_2981);
and UO_110 (O_110,N_2983,N_2962);
or UO_111 (O_111,N_2965,N_2971);
or UO_112 (O_112,N_2956,N_2991);
and UO_113 (O_113,N_2972,N_2965);
nor UO_114 (O_114,N_2958,N_2940);
nor UO_115 (O_115,N_2961,N_2992);
or UO_116 (O_116,N_2959,N_2963);
nor UO_117 (O_117,N_2945,N_2944);
nor UO_118 (O_118,N_2994,N_2972);
and UO_119 (O_119,N_2949,N_2999);
nand UO_120 (O_120,N_2986,N_2992);
nor UO_121 (O_121,N_2999,N_2962);
and UO_122 (O_122,N_2998,N_2970);
nor UO_123 (O_123,N_2992,N_2978);
or UO_124 (O_124,N_2955,N_2941);
nor UO_125 (O_125,N_2995,N_2990);
nor UO_126 (O_126,N_2967,N_2974);
or UO_127 (O_127,N_2996,N_2969);
nor UO_128 (O_128,N_2966,N_2988);
and UO_129 (O_129,N_2981,N_2958);
nand UO_130 (O_130,N_2979,N_2994);
and UO_131 (O_131,N_2985,N_2988);
nor UO_132 (O_132,N_2959,N_2983);
nor UO_133 (O_133,N_2960,N_2988);
nand UO_134 (O_134,N_2953,N_2987);
and UO_135 (O_135,N_2993,N_2971);
nand UO_136 (O_136,N_2985,N_2992);
and UO_137 (O_137,N_2965,N_2967);
nand UO_138 (O_138,N_2954,N_2997);
or UO_139 (O_139,N_2963,N_2943);
or UO_140 (O_140,N_2945,N_2967);
or UO_141 (O_141,N_2969,N_2970);
nor UO_142 (O_142,N_2940,N_2977);
nand UO_143 (O_143,N_2960,N_2944);
and UO_144 (O_144,N_2996,N_2991);
or UO_145 (O_145,N_2968,N_2965);
nor UO_146 (O_146,N_2957,N_2992);
nor UO_147 (O_147,N_2966,N_2976);
and UO_148 (O_148,N_2999,N_2947);
nor UO_149 (O_149,N_2962,N_2966);
nand UO_150 (O_150,N_2980,N_2970);
or UO_151 (O_151,N_2940,N_2948);
or UO_152 (O_152,N_2943,N_2956);
nor UO_153 (O_153,N_2992,N_2952);
and UO_154 (O_154,N_2991,N_2959);
nor UO_155 (O_155,N_2947,N_2996);
or UO_156 (O_156,N_2997,N_2998);
nand UO_157 (O_157,N_2980,N_2942);
nand UO_158 (O_158,N_2959,N_2960);
nand UO_159 (O_159,N_2965,N_2954);
and UO_160 (O_160,N_2949,N_2968);
and UO_161 (O_161,N_2991,N_2997);
or UO_162 (O_162,N_2948,N_2990);
nor UO_163 (O_163,N_2993,N_2959);
xnor UO_164 (O_164,N_2985,N_2973);
nand UO_165 (O_165,N_2973,N_2945);
nand UO_166 (O_166,N_2989,N_2971);
and UO_167 (O_167,N_2999,N_2986);
nand UO_168 (O_168,N_2985,N_2990);
and UO_169 (O_169,N_2991,N_2978);
and UO_170 (O_170,N_2943,N_2967);
nand UO_171 (O_171,N_2940,N_2954);
nor UO_172 (O_172,N_2959,N_2990);
nor UO_173 (O_173,N_2941,N_2971);
nand UO_174 (O_174,N_2958,N_2968);
or UO_175 (O_175,N_2945,N_2941);
nor UO_176 (O_176,N_2987,N_2964);
nand UO_177 (O_177,N_2992,N_2959);
and UO_178 (O_178,N_2958,N_2998);
nor UO_179 (O_179,N_2984,N_2961);
nor UO_180 (O_180,N_2970,N_2987);
or UO_181 (O_181,N_2977,N_2947);
or UO_182 (O_182,N_2948,N_2944);
or UO_183 (O_183,N_2997,N_2970);
and UO_184 (O_184,N_2966,N_2991);
and UO_185 (O_185,N_2968,N_2962);
and UO_186 (O_186,N_2963,N_2953);
nor UO_187 (O_187,N_2997,N_2955);
nor UO_188 (O_188,N_2948,N_2986);
and UO_189 (O_189,N_2949,N_2947);
nand UO_190 (O_190,N_2972,N_2948);
nor UO_191 (O_191,N_2971,N_2940);
or UO_192 (O_192,N_2995,N_2940);
and UO_193 (O_193,N_2978,N_2968);
or UO_194 (O_194,N_2982,N_2964);
and UO_195 (O_195,N_2946,N_2979);
and UO_196 (O_196,N_2993,N_2944);
or UO_197 (O_197,N_2984,N_2958);
and UO_198 (O_198,N_2958,N_2950);
and UO_199 (O_199,N_2988,N_2956);
and UO_200 (O_200,N_2959,N_2958);
nor UO_201 (O_201,N_2962,N_2977);
or UO_202 (O_202,N_2966,N_2982);
xor UO_203 (O_203,N_2948,N_2954);
nand UO_204 (O_204,N_2945,N_2966);
and UO_205 (O_205,N_2986,N_2990);
nor UO_206 (O_206,N_2956,N_2959);
and UO_207 (O_207,N_2982,N_2955);
nor UO_208 (O_208,N_2991,N_2951);
or UO_209 (O_209,N_2971,N_2942);
or UO_210 (O_210,N_2995,N_2988);
and UO_211 (O_211,N_2959,N_2978);
nor UO_212 (O_212,N_2951,N_2995);
or UO_213 (O_213,N_2975,N_2980);
and UO_214 (O_214,N_2999,N_2983);
or UO_215 (O_215,N_2956,N_2951);
or UO_216 (O_216,N_2940,N_2987);
and UO_217 (O_217,N_2940,N_2972);
or UO_218 (O_218,N_2963,N_2942);
nand UO_219 (O_219,N_2966,N_2973);
nor UO_220 (O_220,N_2991,N_2961);
nor UO_221 (O_221,N_2982,N_2962);
xnor UO_222 (O_222,N_2943,N_2998);
or UO_223 (O_223,N_2972,N_2951);
or UO_224 (O_224,N_2956,N_2977);
nand UO_225 (O_225,N_2981,N_2979);
or UO_226 (O_226,N_2986,N_2973);
xor UO_227 (O_227,N_2976,N_2981);
xor UO_228 (O_228,N_2991,N_2948);
nor UO_229 (O_229,N_2941,N_2967);
nand UO_230 (O_230,N_2971,N_2948);
and UO_231 (O_231,N_2967,N_2950);
nand UO_232 (O_232,N_2989,N_2974);
or UO_233 (O_233,N_2999,N_2957);
or UO_234 (O_234,N_2990,N_2946);
and UO_235 (O_235,N_2965,N_2966);
nor UO_236 (O_236,N_2984,N_2944);
nor UO_237 (O_237,N_2952,N_2974);
nand UO_238 (O_238,N_2995,N_2998);
nand UO_239 (O_239,N_2951,N_2988);
and UO_240 (O_240,N_2951,N_2959);
and UO_241 (O_241,N_2955,N_2984);
or UO_242 (O_242,N_2956,N_2989);
nor UO_243 (O_243,N_2942,N_2978);
nor UO_244 (O_244,N_2998,N_2964);
nor UO_245 (O_245,N_2977,N_2954);
and UO_246 (O_246,N_2977,N_2959);
xor UO_247 (O_247,N_2995,N_2959);
or UO_248 (O_248,N_2966,N_2986);
nand UO_249 (O_249,N_2985,N_2967);
xor UO_250 (O_250,N_2999,N_2995);
and UO_251 (O_251,N_2975,N_2976);
nor UO_252 (O_252,N_2961,N_2976);
and UO_253 (O_253,N_2980,N_2991);
nand UO_254 (O_254,N_2956,N_2980);
nor UO_255 (O_255,N_2989,N_2980);
and UO_256 (O_256,N_2998,N_2979);
and UO_257 (O_257,N_2988,N_2963);
and UO_258 (O_258,N_2964,N_2946);
or UO_259 (O_259,N_2980,N_2972);
nor UO_260 (O_260,N_2988,N_2989);
nand UO_261 (O_261,N_2972,N_2988);
nand UO_262 (O_262,N_2963,N_2978);
nand UO_263 (O_263,N_2988,N_2971);
xor UO_264 (O_264,N_2958,N_2975);
xor UO_265 (O_265,N_2971,N_2963);
nand UO_266 (O_266,N_2975,N_2947);
xor UO_267 (O_267,N_2970,N_2983);
nand UO_268 (O_268,N_2954,N_2951);
nand UO_269 (O_269,N_2974,N_2992);
nand UO_270 (O_270,N_2988,N_2953);
or UO_271 (O_271,N_2953,N_2949);
nor UO_272 (O_272,N_2949,N_2952);
or UO_273 (O_273,N_2952,N_2975);
and UO_274 (O_274,N_2941,N_2948);
nand UO_275 (O_275,N_2940,N_2989);
nand UO_276 (O_276,N_2999,N_2979);
nor UO_277 (O_277,N_2961,N_2946);
and UO_278 (O_278,N_2975,N_2956);
nor UO_279 (O_279,N_2945,N_2979);
nand UO_280 (O_280,N_2945,N_2988);
or UO_281 (O_281,N_2944,N_2953);
nor UO_282 (O_282,N_2941,N_2963);
xor UO_283 (O_283,N_2981,N_2993);
and UO_284 (O_284,N_2953,N_2976);
and UO_285 (O_285,N_2943,N_2976);
or UO_286 (O_286,N_2982,N_2985);
nand UO_287 (O_287,N_2959,N_2973);
or UO_288 (O_288,N_2968,N_2940);
and UO_289 (O_289,N_2968,N_2971);
or UO_290 (O_290,N_2993,N_2966);
nor UO_291 (O_291,N_2979,N_2984);
nor UO_292 (O_292,N_2992,N_2973);
and UO_293 (O_293,N_2947,N_2986);
nor UO_294 (O_294,N_2999,N_2972);
and UO_295 (O_295,N_2992,N_2994);
nor UO_296 (O_296,N_2954,N_2941);
nor UO_297 (O_297,N_2968,N_2954);
or UO_298 (O_298,N_2966,N_2971);
or UO_299 (O_299,N_2999,N_2991);
nor UO_300 (O_300,N_2946,N_2974);
and UO_301 (O_301,N_2941,N_2977);
nor UO_302 (O_302,N_2960,N_2984);
or UO_303 (O_303,N_2945,N_2954);
nor UO_304 (O_304,N_2961,N_2998);
nor UO_305 (O_305,N_2991,N_2963);
and UO_306 (O_306,N_2954,N_2970);
nor UO_307 (O_307,N_2978,N_2986);
and UO_308 (O_308,N_2988,N_2978);
or UO_309 (O_309,N_2951,N_2950);
or UO_310 (O_310,N_2980,N_2944);
nor UO_311 (O_311,N_2943,N_2972);
xnor UO_312 (O_312,N_2958,N_2946);
nand UO_313 (O_313,N_2994,N_2986);
nand UO_314 (O_314,N_2999,N_2966);
or UO_315 (O_315,N_2995,N_2983);
nand UO_316 (O_316,N_2997,N_2960);
or UO_317 (O_317,N_2961,N_2979);
nand UO_318 (O_318,N_2991,N_2975);
and UO_319 (O_319,N_2949,N_2972);
and UO_320 (O_320,N_2951,N_2998);
nand UO_321 (O_321,N_2969,N_2992);
nand UO_322 (O_322,N_2979,N_2940);
and UO_323 (O_323,N_2992,N_2951);
or UO_324 (O_324,N_2998,N_2992);
nand UO_325 (O_325,N_2992,N_2971);
nor UO_326 (O_326,N_2943,N_2992);
nor UO_327 (O_327,N_2994,N_2942);
nor UO_328 (O_328,N_2957,N_2963);
nor UO_329 (O_329,N_2961,N_2957);
nor UO_330 (O_330,N_2943,N_2995);
nand UO_331 (O_331,N_2961,N_2985);
or UO_332 (O_332,N_2994,N_2977);
xor UO_333 (O_333,N_2989,N_2949);
nand UO_334 (O_334,N_2977,N_2983);
and UO_335 (O_335,N_2976,N_2991);
nor UO_336 (O_336,N_2968,N_2975);
and UO_337 (O_337,N_2991,N_2971);
or UO_338 (O_338,N_2956,N_2973);
or UO_339 (O_339,N_2965,N_2996);
and UO_340 (O_340,N_2940,N_2946);
or UO_341 (O_341,N_2978,N_2980);
nand UO_342 (O_342,N_2982,N_2983);
nor UO_343 (O_343,N_2977,N_2945);
nor UO_344 (O_344,N_2964,N_2992);
or UO_345 (O_345,N_2987,N_2951);
nor UO_346 (O_346,N_2947,N_2945);
nand UO_347 (O_347,N_2941,N_2975);
and UO_348 (O_348,N_2965,N_2980);
or UO_349 (O_349,N_2971,N_2964);
and UO_350 (O_350,N_2991,N_2986);
nor UO_351 (O_351,N_2958,N_2983);
or UO_352 (O_352,N_2950,N_2991);
and UO_353 (O_353,N_2988,N_2973);
and UO_354 (O_354,N_2958,N_2989);
nand UO_355 (O_355,N_2942,N_2976);
or UO_356 (O_356,N_2969,N_2960);
and UO_357 (O_357,N_2967,N_2952);
xor UO_358 (O_358,N_2993,N_2969);
and UO_359 (O_359,N_2944,N_2954);
and UO_360 (O_360,N_2970,N_2947);
and UO_361 (O_361,N_2947,N_2941);
nand UO_362 (O_362,N_2961,N_2974);
and UO_363 (O_363,N_2943,N_2987);
and UO_364 (O_364,N_2951,N_2977);
or UO_365 (O_365,N_2943,N_2944);
or UO_366 (O_366,N_2940,N_2996);
or UO_367 (O_367,N_2986,N_2993);
nand UO_368 (O_368,N_2988,N_2957);
nor UO_369 (O_369,N_2985,N_2949);
nand UO_370 (O_370,N_2988,N_2970);
nor UO_371 (O_371,N_2990,N_2999);
and UO_372 (O_372,N_2984,N_2989);
nor UO_373 (O_373,N_2998,N_2953);
nor UO_374 (O_374,N_2992,N_2995);
or UO_375 (O_375,N_2959,N_2964);
or UO_376 (O_376,N_2947,N_2995);
nand UO_377 (O_377,N_2949,N_2962);
and UO_378 (O_378,N_2980,N_2976);
or UO_379 (O_379,N_2991,N_2972);
and UO_380 (O_380,N_2999,N_2956);
nor UO_381 (O_381,N_2940,N_2973);
and UO_382 (O_382,N_2943,N_2996);
and UO_383 (O_383,N_2985,N_2997);
nor UO_384 (O_384,N_2948,N_2980);
and UO_385 (O_385,N_2953,N_2961);
nand UO_386 (O_386,N_2952,N_2942);
nor UO_387 (O_387,N_2969,N_2995);
nand UO_388 (O_388,N_2950,N_2954);
nor UO_389 (O_389,N_2986,N_2954);
nor UO_390 (O_390,N_2940,N_2969);
and UO_391 (O_391,N_2963,N_2977);
nand UO_392 (O_392,N_2953,N_2969);
nand UO_393 (O_393,N_2982,N_2984);
nor UO_394 (O_394,N_2971,N_2945);
or UO_395 (O_395,N_2953,N_2955);
nor UO_396 (O_396,N_2959,N_2996);
nand UO_397 (O_397,N_2977,N_2997);
nand UO_398 (O_398,N_2988,N_2961);
or UO_399 (O_399,N_2965,N_2994);
and UO_400 (O_400,N_2952,N_2986);
nor UO_401 (O_401,N_2971,N_2954);
and UO_402 (O_402,N_2941,N_2989);
and UO_403 (O_403,N_2989,N_2947);
nor UO_404 (O_404,N_2998,N_2950);
xor UO_405 (O_405,N_2943,N_2985);
nand UO_406 (O_406,N_2976,N_2995);
nor UO_407 (O_407,N_2981,N_2989);
or UO_408 (O_408,N_2993,N_2949);
nor UO_409 (O_409,N_2994,N_2953);
nor UO_410 (O_410,N_2967,N_2966);
and UO_411 (O_411,N_2996,N_2951);
or UO_412 (O_412,N_2961,N_2959);
and UO_413 (O_413,N_2983,N_2997);
nor UO_414 (O_414,N_2949,N_2976);
nor UO_415 (O_415,N_2967,N_2980);
or UO_416 (O_416,N_2995,N_2942);
nor UO_417 (O_417,N_2966,N_2992);
nor UO_418 (O_418,N_2947,N_2954);
or UO_419 (O_419,N_2949,N_2958);
or UO_420 (O_420,N_2947,N_2955);
nand UO_421 (O_421,N_2947,N_2967);
nor UO_422 (O_422,N_2962,N_2981);
nand UO_423 (O_423,N_2975,N_2967);
nor UO_424 (O_424,N_2980,N_2946);
nor UO_425 (O_425,N_2982,N_2943);
or UO_426 (O_426,N_2980,N_2971);
nor UO_427 (O_427,N_2953,N_2979);
nand UO_428 (O_428,N_2972,N_2962);
or UO_429 (O_429,N_2996,N_2950);
or UO_430 (O_430,N_2946,N_2969);
and UO_431 (O_431,N_2996,N_2984);
nor UO_432 (O_432,N_2995,N_2944);
nand UO_433 (O_433,N_2977,N_2986);
nand UO_434 (O_434,N_2984,N_2986);
nand UO_435 (O_435,N_2993,N_2980);
nor UO_436 (O_436,N_2984,N_2977);
and UO_437 (O_437,N_2975,N_2966);
nand UO_438 (O_438,N_2949,N_2990);
or UO_439 (O_439,N_2975,N_2946);
nor UO_440 (O_440,N_2948,N_2958);
nand UO_441 (O_441,N_2995,N_2977);
nor UO_442 (O_442,N_2990,N_2997);
nand UO_443 (O_443,N_2964,N_2966);
and UO_444 (O_444,N_2991,N_2946);
and UO_445 (O_445,N_2999,N_2973);
nor UO_446 (O_446,N_2989,N_2968);
and UO_447 (O_447,N_2941,N_2996);
nand UO_448 (O_448,N_2990,N_2992);
and UO_449 (O_449,N_2948,N_2945);
or UO_450 (O_450,N_2985,N_2979);
nand UO_451 (O_451,N_2944,N_2958);
and UO_452 (O_452,N_2972,N_2996);
nand UO_453 (O_453,N_2981,N_2965);
xnor UO_454 (O_454,N_2997,N_2947);
nor UO_455 (O_455,N_2965,N_2982);
nor UO_456 (O_456,N_2978,N_2961);
or UO_457 (O_457,N_2969,N_2973);
nor UO_458 (O_458,N_2952,N_2984);
nand UO_459 (O_459,N_2946,N_2963);
nor UO_460 (O_460,N_2978,N_2984);
nand UO_461 (O_461,N_2942,N_2958);
or UO_462 (O_462,N_2979,N_2962);
or UO_463 (O_463,N_2979,N_2992);
xor UO_464 (O_464,N_2942,N_2949);
nand UO_465 (O_465,N_2943,N_2977);
and UO_466 (O_466,N_2983,N_2952);
nor UO_467 (O_467,N_2971,N_2956);
nor UO_468 (O_468,N_2980,N_2986);
nand UO_469 (O_469,N_2978,N_2996);
or UO_470 (O_470,N_2947,N_2985);
or UO_471 (O_471,N_2984,N_2940);
nand UO_472 (O_472,N_2982,N_2975);
or UO_473 (O_473,N_2948,N_2994);
and UO_474 (O_474,N_2989,N_2975);
and UO_475 (O_475,N_2970,N_2949);
nand UO_476 (O_476,N_2985,N_2983);
nand UO_477 (O_477,N_2972,N_2942);
or UO_478 (O_478,N_2981,N_2985);
nor UO_479 (O_479,N_2960,N_2981);
nor UO_480 (O_480,N_2994,N_2973);
nor UO_481 (O_481,N_2971,N_2979);
and UO_482 (O_482,N_2940,N_2981);
xnor UO_483 (O_483,N_2974,N_2996);
nor UO_484 (O_484,N_2989,N_2966);
nor UO_485 (O_485,N_2990,N_2945);
nor UO_486 (O_486,N_2985,N_2987);
nand UO_487 (O_487,N_2958,N_2964);
nor UO_488 (O_488,N_2965,N_2974);
nor UO_489 (O_489,N_2994,N_2957);
or UO_490 (O_490,N_2977,N_2970);
nor UO_491 (O_491,N_2970,N_2944);
nand UO_492 (O_492,N_2997,N_2989);
and UO_493 (O_493,N_2954,N_2949);
nor UO_494 (O_494,N_2942,N_2999);
nand UO_495 (O_495,N_2953,N_2983);
nor UO_496 (O_496,N_2960,N_2994);
nand UO_497 (O_497,N_2952,N_2972);
and UO_498 (O_498,N_2989,N_2995);
or UO_499 (O_499,N_2998,N_2956);
endmodule