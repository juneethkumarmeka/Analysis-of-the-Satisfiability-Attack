module basic_500_3000_500_15_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_102,In_100);
or U1 (N_1,In_467,In_349);
and U2 (N_2,In_436,In_141);
nor U3 (N_3,In_125,In_220);
nor U4 (N_4,In_275,In_137);
nor U5 (N_5,In_7,In_442);
or U6 (N_6,In_21,In_138);
nand U7 (N_7,In_147,In_129);
nand U8 (N_8,In_395,In_152);
nand U9 (N_9,In_0,In_381);
nand U10 (N_10,In_469,In_203);
or U11 (N_11,In_418,In_95);
or U12 (N_12,In_456,In_330);
nor U13 (N_13,In_72,In_475);
or U14 (N_14,In_334,In_422);
nor U15 (N_15,In_339,In_325);
and U16 (N_16,In_459,In_350);
xor U17 (N_17,In_342,In_87);
nor U18 (N_18,In_289,In_435);
and U19 (N_19,In_460,In_341);
nand U20 (N_20,In_321,In_242);
xor U21 (N_21,In_133,In_382);
and U22 (N_22,In_298,In_450);
and U23 (N_23,In_486,In_54);
or U24 (N_24,In_304,In_157);
nand U25 (N_25,In_358,In_481);
or U26 (N_26,In_470,In_445);
nor U27 (N_27,In_66,In_288);
nor U28 (N_28,In_114,In_367);
and U29 (N_29,In_361,In_338);
and U30 (N_30,In_463,In_256);
or U31 (N_31,In_85,In_491);
nand U32 (N_32,In_294,In_162);
xor U33 (N_33,In_441,In_187);
xor U34 (N_34,In_226,In_354);
nor U35 (N_35,In_42,In_202);
nand U36 (N_36,In_167,In_8);
nor U37 (N_37,In_483,In_245);
and U38 (N_38,In_472,In_179);
nand U39 (N_39,In_130,In_253);
xnor U40 (N_40,In_91,In_333);
nand U41 (N_41,In_433,In_163);
nand U42 (N_42,In_28,In_158);
and U43 (N_43,In_399,In_112);
or U44 (N_44,In_105,In_420);
or U45 (N_45,In_410,In_171);
xnor U46 (N_46,In_413,In_353);
or U47 (N_47,In_232,In_207);
nor U48 (N_48,In_113,In_303);
nand U49 (N_49,In_89,In_444);
nand U50 (N_50,In_53,In_364);
and U51 (N_51,In_192,In_336);
or U52 (N_52,In_498,In_430);
nand U53 (N_53,In_379,In_396);
xnor U54 (N_54,In_58,In_238);
nand U55 (N_55,In_33,In_205);
or U56 (N_56,In_188,In_165);
nor U57 (N_57,In_313,In_380);
and U58 (N_58,In_284,In_328);
or U59 (N_59,In_327,In_219);
and U60 (N_60,In_305,In_216);
nand U61 (N_61,In_355,In_371);
nor U62 (N_62,In_293,In_168);
nand U63 (N_63,In_123,In_79);
or U64 (N_64,In_34,In_406);
or U65 (N_65,In_269,In_57);
or U66 (N_66,In_356,In_485);
and U67 (N_67,In_128,In_496);
nor U68 (N_68,In_309,In_368);
or U69 (N_69,In_393,In_191);
xnor U70 (N_70,In_223,In_94);
nand U71 (N_71,In_407,In_97);
xnor U72 (N_72,In_440,In_365);
nor U73 (N_73,In_416,In_77);
and U74 (N_74,In_434,In_24);
nor U75 (N_75,In_65,In_131);
nor U76 (N_76,In_111,In_47);
xnor U77 (N_77,In_46,In_98);
or U78 (N_78,In_262,In_474);
nor U79 (N_79,In_362,In_489);
xnor U80 (N_80,In_84,In_344);
xnor U81 (N_81,In_447,In_493);
nor U82 (N_82,In_295,In_3);
xor U83 (N_83,In_118,In_1);
or U84 (N_84,In_88,In_259);
nor U85 (N_85,In_117,In_190);
nand U86 (N_86,In_124,In_5);
or U87 (N_87,In_211,In_348);
and U88 (N_88,In_161,In_222);
xor U89 (N_89,In_408,In_227);
xor U90 (N_90,In_306,In_308);
or U91 (N_91,In_80,In_402);
and U92 (N_92,In_268,In_264);
or U93 (N_93,In_400,In_409);
nor U94 (N_94,In_311,In_215);
or U95 (N_95,In_153,In_283);
and U96 (N_96,In_213,In_499);
nor U97 (N_97,In_43,In_329);
xnor U98 (N_98,In_140,In_487);
nor U99 (N_99,In_18,In_240);
nand U100 (N_100,In_482,In_70);
xor U101 (N_101,In_476,In_189);
and U102 (N_102,In_297,In_390);
xnor U103 (N_103,In_360,In_438);
nand U104 (N_104,In_225,In_170);
xor U105 (N_105,In_398,In_174);
or U106 (N_106,In_116,In_107);
xnor U107 (N_107,In_462,In_307);
xor U108 (N_108,In_431,In_250);
or U109 (N_109,In_40,In_51);
and U110 (N_110,In_251,In_108);
and U111 (N_111,In_455,In_119);
nor U112 (N_112,In_217,In_263);
and U113 (N_113,In_201,In_452);
nor U114 (N_114,In_258,In_479);
nor U115 (N_115,In_428,In_224);
or U116 (N_116,In_101,In_468);
xor U117 (N_117,In_247,In_443);
nor U118 (N_118,In_279,In_50);
and U119 (N_119,In_175,In_302);
nand U120 (N_120,In_415,In_372);
nor U121 (N_121,In_246,In_121);
nor U122 (N_122,In_331,In_271);
nor U123 (N_123,In_86,In_347);
nor U124 (N_124,In_241,In_414);
xor U125 (N_125,In_480,In_404);
nor U126 (N_126,In_494,In_44);
nand U127 (N_127,In_437,In_388);
or U128 (N_128,In_159,In_52);
or U129 (N_129,In_451,In_461);
nor U130 (N_130,In_373,In_290);
nor U131 (N_131,In_149,In_243);
nand U132 (N_132,In_204,In_239);
and U133 (N_133,In_104,In_343);
xor U134 (N_134,In_25,In_424);
nand U135 (N_135,In_139,In_335);
nand U136 (N_136,In_249,In_230);
xor U137 (N_137,In_26,In_6);
and U138 (N_138,In_401,In_370);
xor U139 (N_139,In_495,In_48);
and U140 (N_140,In_120,In_312);
or U141 (N_141,In_425,In_292);
and U142 (N_142,In_314,In_352);
nand U143 (N_143,In_69,In_369);
and U144 (N_144,In_62,In_439);
nor U145 (N_145,In_169,In_197);
and U146 (N_146,In_71,In_200);
nor U147 (N_147,In_75,In_142);
and U148 (N_148,In_454,In_233);
and U149 (N_149,In_173,In_31);
and U150 (N_150,In_260,In_229);
nand U151 (N_151,In_15,In_81);
and U152 (N_152,In_411,In_180);
and U153 (N_153,In_377,In_340);
and U154 (N_154,In_417,In_389);
nor U155 (N_155,In_196,In_134);
xor U156 (N_156,In_27,In_2);
nor U157 (N_157,In_11,In_255);
nor U158 (N_158,In_148,In_317);
nand U159 (N_159,In_273,In_392);
or U160 (N_160,In_199,In_41);
or U161 (N_161,In_301,In_237);
nand U162 (N_162,In_277,In_266);
nor U163 (N_163,In_310,In_144);
and U164 (N_164,In_135,In_16);
and U165 (N_165,In_109,In_429);
nand U166 (N_166,In_9,In_166);
and U167 (N_167,In_235,In_29);
and U168 (N_168,In_272,In_160);
or U169 (N_169,In_198,In_56);
nor U170 (N_170,In_453,In_82);
and U171 (N_171,In_126,In_244);
and U172 (N_172,In_385,In_68);
and U173 (N_173,In_218,In_276);
nand U174 (N_174,In_146,In_186);
and U175 (N_175,In_90,In_99);
nand U176 (N_176,In_359,In_67);
xnor U177 (N_177,In_92,In_194);
or U178 (N_178,In_384,In_181);
xor U179 (N_179,In_136,In_35);
nor U180 (N_180,In_150,In_281);
xor U181 (N_181,In_326,In_208);
or U182 (N_182,In_19,In_346);
and U183 (N_183,In_465,In_300);
and U184 (N_184,In_466,In_457);
nor U185 (N_185,In_387,In_405);
or U186 (N_186,In_60,In_285);
xnor U187 (N_187,In_497,In_156);
xor U188 (N_188,In_257,In_363);
nand U189 (N_189,In_478,In_151);
xor U190 (N_190,In_164,In_177);
or U191 (N_191,In_299,In_261);
nand U192 (N_192,In_426,In_74);
and U193 (N_193,In_378,In_63);
nand U194 (N_194,In_403,In_446);
nand U195 (N_195,In_397,In_287);
nor U196 (N_196,In_10,In_316);
nor U197 (N_197,In_83,In_22);
xor U198 (N_198,In_391,In_449);
or U199 (N_199,In_351,In_145);
or U200 (N_200,N_127,N_88);
xnor U201 (N_201,N_83,N_82);
nand U202 (N_202,N_21,N_33);
or U203 (N_203,N_111,In_172);
nand U204 (N_204,In_394,N_58);
nor U205 (N_205,N_90,N_46);
nor U206 (N_206,In_64,N_161);
and U207 (N_207,N_120,In_14);
nand U208 (N_208,N_7,N_128);
and U209 (N_209,In_206,In_76);
and U210 (N_210,In_127,N_56);
nor U211 (N_211,N_67,N_75);
and U212 (N_212,In_421,N_41);
nor U213 (N_213,N_118,In_221);
xnor U214 (N_214,In_473,In_296);
nand U215 (N_215,In_231,N_27);
nand U216 (N_216,N_122,N_129);
or U217 (N_217,N_152,N_153);
or U218 (N_218,N_177,N_60);
xnor U219 (N_219,N_194,N_132);
or U220 (N_220,N_74,N_32);
and U221 (N_221,N_186,In_427);
and U222 (N_222,N_106,N_179);
and U223 (N_223,N_101,N_57);
and U224 (N_224,N_143,N_49);
xor U225 (N_225,N_17,N_87);
and U226 (N_226,N_18,N_1);
nor U227 (N_227,In_432,N_43);
nand U228 (N_228,N_38,In_412);
xnor U229 (N_229,In_59,N_73);
or U230 (N_230,N_97,N_29);
nand U231 (N_231,In_154,In_210);
nor U232 (N_232,N_171,N_189);
and U233 (N_233,N_45,In_383);
nor U234 (N_234,N_37,N_137);
or U235 (N_235,N_191,In_319);
nand U236 (N_236,N_42,N_25);
nor U237 (N_237,N_113,N_104);
or U238 (N_238,In_270,N_183);
and U239 (N_239,N_8,In_12);
and U240 (N_240,In_320,N_64);
or U241 (N_241,N_110,N_176);
nand U242 (N_242,N_71,In_122);
nand U243 (N_243,N_135,N_94);
xnor U244 (N_244,N_63,N_3);
nand U245 (N_245,N_48,In_252);
nand U246 (N_246,In_375,In_386);
and U247 (N_247,N_156,In_423);
nor U248 (N_248,In_73,In_492);
nor U249 (N_249,In_93,N_154);
and U250 (N_250,In_49,N_198);
nand U251 (N_251,N_61,N_28);
nor U252 (N_252,N_100,In_323);
and U253 (N_253,N_35,N_170);
and U254 (N_254,N_15,N_172);
and U255 (N_255,N_117,N_187);
xor U256 (N_256,N_199,In_38);
xnor U257 (N_257,In_315,In_291);
or U258 (N_258,In_337,In_182);
nor U259 (N_259,N_193,N_14);
and U260 (N_260,N_138,N_31);
or U261 (N_261,N_51,N_24);
nand U262 (N_262,In_32,In_55);
nand U263 (N_263,In_195,In_286);
nor U264 (N_264,In_265,N_144);
nor U265 (N_265,N_99,In_282);
nor U266 (N_266,N_166,N_80);
or U267 (N_267,N_165,N_69);
and U268 (N_268,N_164,In_176);
or U269 (N_269,N_195,N_124);
nand U270 (N_270,In_254,In_96);
nand U271 (N_271,N_70,N_140);
or U272 (N_272,N_157,In_278);
or U273 (N_273,N_115,N_150);
nand U274 (N_274,N_91,N_96);
nor U275 (N_275,N_167,N_89);
xor U276 (N_276,In_45,N_185);
or U277 (N_277,N_148,N_178);
xnor U278 (N_278,N_62,N_40);
nand U279 (N_279,N_168,In_185);
and U280 (N_280,In_143,In_484);
xnor U281 (N_281,N_163,In_488);
or U282 (N_282,In_477,N_12);
or U283 (N_283,N_181,N_196);
and U284 (N_284,In_471,In_178);
xor U285 (N_285,N_162,In_322);
nand U286 (N_286,In_37,In_36);
nand U287 (N_287,N_2,N_182);
or U288 (N_288,N_16,N_76);
nor U289 (N_289,N_6,N_109);
xor U290 (N_290,In_234,N_95);
or U291 (N_291,In_366,N_10);
and U292 (N_292,N_44,N_54);
or U293 (N_293,N_9,N_126);
xnor U294 (N_294,In_61,In_448);
nand U295 (N_295,N_55,N_175);
or U296 (N_296,In_376,N_125);
nand U297 (N_297,N_119,In_184);
nor U298 (N_298,N_103,In_132);
nor U299 (N_299,In_490,N_19);
nor U300 (N_300,In_214,N_188);
and U301 (N_301,N_53,N_112);
xnor U302 (N_302,N_34,N_108);
and U303 (N_303,N_174,N_79);
xnor U304 (N_304,In_193,In_357);
and U305 (N_305,In_318,N_121);
and U306 (N_306,In_419,N_147);
nand U307 (N_307,In_345,N_151);
xnor U308 (N_308,N_0,In_183);
nand U309 (N_309,N_47,N_155);
or U310 (N_310,N_131,N_72);
and U311 (N_311,N_105,N_192);
xnor U312 (N_312,N_52,N_68);
and U313 (N_313,N_130,N_20);
xor U314 (N_314,N_141,N_5);
xnor U315 (N_315,N_98,N_85);
nand U316 (N_316,N_11,N_59);
xor U317 (N_317,In_236,N_65);
and U318 (N_318,N_116,N_26);
nor U319 (N_319,In_30,In_23);
and U320 (N_320,N_114,In_280);
nor U321 (N_321,In_374,N_77);
xor U322 (N_322,N_84,In_4);
and U323 (N_323,N_22,In_110);
or U324 (N_324,N_78,N_146);
and U325 (N_325,In_464,N_50);
and U326 (N_326,In_103,N_160);
nand U327 (N_327,N_36,N_134);
nor U328 (N_328,N_93,N_190);
or U329 (N_329,N_145,In_115);
nor U330 (N_330,N_142,In_274);
or U331 (N_331,In_106,N_92);
nor U332 (N_332,N_173,N_86);
or U333 (N_333,N_30,N_13);
xor U334 (N_334,N_81,N_169);
xnor U335 (N_335,In_39,In_20);
and U336 (N_336,N_197,N_66);
nand U337 (N_337,In_209,In_458);
and U338 (N_338,N_149,N_184);
or U339 (N_339,N_139,N_136);
nor U340 (N_340,N_123,In_155);
and U341 (N_341,In_332,In_13);
xnor U342 (N_342,In_324,N_107);
nand U343 (N_343,N_102,In_78);
and U344 (N_344,N_180,In_17);
or U345 (N_345,N_23,In_228);
nand U346 (N_346,N_159,N_39);
nand U347 (N_347,N_133,In_248);
nand U348 (N_348,In_212,In_267);
and U349 (N_349,N_4,N_158);
and U350 (N_350,In_473,N_170);
xor U351 (N_351,In_394,N_171);
and U352 (N_352,N_196,N_4);
or U353 (N_353,In_320,N_108);
xnor U354 (N_354,N_121,In_132);
or U355 (N_355,N_181,In_49);
nor U356 (N_356,In_386,N_9);
or U357 (N_357,In_195,In_248);
and U358 (N_358,In_357,N_6);
and U359 (N_359,In_59,N_175);
xnor U360 (N_360,N_35,N_96);
or U361 (N_361,N_80,N_55);
nand U362 (N_362,N_0,N_130);
nor U363 (N_363,In_221,N_73);
or U364 (N_364,N_139,N_117);
xor U365 (N_365,In_484,In_96);
xnor U366 (N_366,N_80,In_132);
nand U367 (N_367,N_0,N_158);
and U368 (N_368,N_90,N_104);
nor U369 (N_369,In_122,N_125);
xnor U370 (N_370,In_122,N_135);
and U371 (N_371,N_72,In_490);
or U372 (N_372,N_193,N_182);
or U373 (N_373,N_65,N_13);
xnor U374 (N_374,In_122,In_280);
nor U375 (N_375,N_86,In_23);
nand U376 (N_376,In_183,N_70);
nand U377 (N_377,N_79,N_109);
and U378 (N_378,In_228,N_31);
xnor U379 (N_379,In_488,In_183);
nand U380 (N_380,N_124,N_130);
xnor U381 (N_381,In_45,In_4);
or U382 (N_382,N_39,In_206);
nand U383 (N_383,N_133,N_6);
nor U384 (N_384,In_427,N_78);
nor U385 (N_385,In_178,N_123);
or U386 (N_386,In_115,N_132);
nand U387 (N_387,N_63,N_153);
and U388 (N_388,In_176,In_236);
or U389 (N_389,In_383,In_64);
xor U390 (N_390,In_110,In_214);
or U391 (N_391,In_73,In_337);
and U392 (N_392,N_42,N_181);
nor U393 (N_393,N_199,In_127);
nor U394 (N_394,N_34,N_68);
and U395 (N_395,N_121,N_84);
or U396 (N_396,N_73,In_323);
nor U397 (N_397,In_210,N_48);
xor U398 (N_398,N_47,In_458);
or U399 (N_399,In_143,N_36);
xnor U400 (N_400,N_397,N_219);
nand U401 (N_401,N_359,N_246);
or U402 (N_402,N_230,N_335);
or U403 (N_403,N_317,N_232);
nand U404 (N_404,N_269,N_255);
or U405 (N_405,N_346,N_340);
nand U406 (N_406,N_310,N_356);
xnor U407 (N_407,N_308,N_293);
nor U408 (N_408,N_378,N_316);
nand U409 (N_409,N_267,N_324);
or U410 (N_410,N_320,N_396);
or U411 (N_411,N_390,N_361);
xor U412 (N_412,N_315,N_279);
or U413 (N_413,N_253,N_264);
and U414 (N_414,N_341,N_223);
xnor U415 (N_415,N_290,N_212);
xnor U416 (N_416,N_278,N_399);
nor U417 (N_417,N_202,N_242);
nor U418 (N_418,N_234,N_348);
nand U419 (N_419,N_275,N_265);
xnor U420 (N_420,N_231,N_323);
and U421 (N_421,N_214,N_298);
or U422 (N_422,N_363,N_259);
nor U423 (N_423,N_371,N_209);
and U424 (N_424,N_254,N_235);
and U425 (N_425,N_225,N_244);
xor U426 (N_426,N_383,N_365);
xor U427 (N_427,N_252,N_273);
or U428 (N_428,N_307,N_206);
xnor U429 (N_429,N_301,N_398);
and U430 (N_430,N_328,N_380);
nand U431 (N_431,N_210,N_326);
and U432 (N_432,N_220,N_221);
and U433 (N_433,N_387,N_297);
or U434 (N_434,N_286,N_362);
or U435 (N_435,N_215,N_271);
or U436 (N_436,N_224,N_207);
nor U437 (N_437,N_337,N_395);
or U438 (N_438,N_236,N_276);
xnor U439 (N_439,N_353,N_249);
nor U440 (N_440,N_327,N_201);
nand U441 (N_441,N_374,N_218);
nor U442 (N_442,N_262,N_368);
or U443 (N_443,N_313,N_258);
or U444 (N_444,N_299,N_281);
nand U445 (N_445,N_302,N_243);
and U446 (N_446,N_248,N_217);
xnor U447 (N_447,N_304,N_237);
and U448 (N_448,N_332,N_343);
nor U449 (N_449,N_204,N_208);
xor U450 (N_450,N_355,N_291);
nor U451 (N_451,N_367,N_266);
or U452 (N_452,N_300,N_283);
xor U453 (N_453,N_285,N_330);
and U454 (N_454,N_222,N_280);
nand U455 (N_455,N_239,N_388);
or U456 (N_456,N_241,N_296);
nor U457 (N_457,N_311,N_385);
and U458 (N_458,N_288,N_268);
nor U459 (N_459,N_274,N_389);
or U460 (N_460,N_379,N_391);
and U461 (N_461,N_227,N_382);
and U462 (N_462,N_305,N_357);
and U463 (N_463,N_345,N_270);
nor U464 (N_464,N_303,N_229);
nand U465 (N_465,N_256,N_322);
xnor U466 (N_466,N_205,N_336);
nor U467 (N_467,N_257,N_384);
xnor U468 (N_468,N_375,N_247);
nor U469 (N_469,N_211,N_294);
and U470 (N_470,N_284,N_347);
nor U471 (N_471,N_344,N_372);
xnor U472 (N_472,N_312,N_350);
and U473 (N_473,N_360,N_366);
or U474 (N_474,N_376,N_203);
or U475 (N_475,N_216,N_245);
nor U476 (N_476,N_338,N_394);
and U477 (N_477,N_321,N_238);
and U478 (N_478,N_289,N_272);
or U479 (N_479,N_331,N_333);
or U480 (N_480,N_364,N_373);
nand U481 (N_481,N_319,N_261);
and U482 (N_482,N_213,N_349);
xor U483 (N_483,N_295,N_377);
nand U484 (N_484,N_306,N_200);
or U485 (N_485,N_318,N_352);
nand U486 (N_486,N_277,N_287);
or U487 (N_487,N_260,N_358);
and U488 (N_488,N_369,N_251);
nor U489 (N_489,N_325,N_351);
and U490 (N_490,N_370,N_240);
nor U491 (N_491,N_292,N_250);
and U492 (N_492,N_263,N_233);
or U493 (N_493,N_392,N_386);
and U494 (N_494,N_339,N_314);
xor U495 (N_495,N_309,N_282);
nand U496 (N_496,N_334,N_228);
nor U497 (N_497,N_354,N_393);
nand U498 (N_498,N_226,N_342);
and U499 (N_499,N_381,N_329);
xor U500 (N_500,N_334,N_390);
xnor U501 (N_501,N_250,N_319);
or U502 (N_502,N_380,N_258);
or U503 (N_503,N_243,N_206);
nor U504 (N_504,N_333,N_255);
nor U505 (N_505,N_398,N_220);
nand U506 (N_506,N_361,N_359);
or U507 (N_507,N_207,N_379);
xnor U508 (N_508,N_343,N_394);
and U509 (N_509,N_358,N_328);
nor U510 (N_510,N_380,N_398);
xor U511 (N_511,N_319,N_257);
xnor U512 (N_512,N_395,N_246);
nand U513 (N_513,N_395,N_346);
nor U514 (N_514,N_250,N_361);
and U515 (N_515,N_211,N_234);
xor U516 (N_516,N_346,N_236);
and U517 (N_517,N_375,N_305);
nor U518 (N_518,N_266,N_395);
xnor U519 (N_519,N_223,N_213);
and U520 (N_520,N_351,N_329);
and U521 (N_521,N_209,N_242);
or U522 (N_522,N_242,N_290);
and U523 (N_523,N_325,N_371);
and U524 (N_524,N_211,N_244);
xor U525 (N_525,N_208,N_220);
and U526 (N_526,N_256,N_337);
nor U527 (N_527,N_315,N_321);
xor U528 (N_528,N_285,N_382);
nor U529 (N_529,N_204,N_309);
xnor U530 (N_530,N_261,N_324);
nor U531 (N_531,N_287,N_214);
nand U532 (N_532,N_232,N_205);
and U533 (N_533,N_291,N_338);
and U534 (N_534,N_233,N_355);
nand U535 (N_535,N_381,N_316);
nand U536 (N_536,N_270,N_215);
nand U537 (N_537,N_357,N_260);
nor U538 (N_538,N_275,N_347);
nor U539 (N_539,N_234,N_355);
or U540 (N_540,N_383,N_299);
nor U541 (N_541,N_327,N_248);
nor U542 (N_542,N_361,N_268);
or U543 (N_543,N_257,N_267);
nor U544 (N_544,N_328,N_285);
nor U545 (N_545,N_274,N_357);
xor U546 (N_546,N_348,N_261);
and U547 (N_547,N_346,N_299);
and U548 (N_548,N_294,N_363);
or U549 (N_549,N_302,N_297);
nand U550 (N_550,N_338,N_383);
and U551 (N_551,N_376,N_333);
nand U552 (N_552,N_274,N_229);
nor U553 (N_553,N_379,N_335);
nand U554 (N_554,N_271,N_341);
nor U555 (N_555,N_310,N_316);
and U556 (N_556,N_294,N_373);
nand U557 (N_557,N_335,N_237);
and U558 (N_558,N_235,N_324);
and U559 (N_559,N_215,N_249);
nor U560 (N_560,N_239,N_227);
nor U561 (N_561,N_326,N_292);
or U562 (N_562,N_281,N_325);
nand U563 (N_563,N_305,N_393);
or U564 (N_564,N_224,N_294);
nand U565 (N_565,N_232,N_387);
or U566 (N_566,N_249,N_295);
nor U567 (N_567,N_362,N_374);
xnor U568 (N_568,N_225,N_342);
and U569 (N_569,N_376,N_307);
nand U570 (N_570,N_256,N_375);
and U571 (N_571,N_264,N_245);
or U572 (N_572,N_350,N_393);
nor U573 (N_573,N_293,N_397);
or U574 (N_574,N_385,N_289);
or U575 (N_575,N_378,N_321);
xor U576 (N_576,N_345,N_235);
xor U577 (N_577,N_309,N_391);
xor U578 (N_578,N_292,N_366);
xnor U579 (N_579,N_349,N_276);
xnor U580 (N_580,N_310,N_290);
nor U581 (N_581,N_380,N_353);
nor U582 (N_582,N_255,N_316);
or U583 (N_583,N_248,N_359);
xnor U584 (N_584,N_243,N_335);
xnor U585 (N_585,N_367,N_299);
xor U586 (N_586,N_341,N_399);
and U587 (N_587,N_247,N_280);
xnor U588 (N_588,N_201,N_272);
nand U589 (N_589,N_364,N_332);
nor U590 (N_590,N_209,N_276);
and U591 (N_591,N_292,N_396);
nand U592 (N_592,N_320,N_355);
or U593 (N_593,N_345,N_207);
and U594 (N_594,N_323,N_370);
nor U595 (N_595,N_352,N_214);
nand U596 (N_596,N_386,N_310);
nor U597 (N_597,N_234,N_354);
or U598 (N_598,N_339,N_236);
nor U599 (N_599,N_291,N_323);
and U600 (N_600,N_457,N_563);
and U601 (N_601,N_562,N_536);
and U602 (N_602,N_450,N_557);
xor U603 (N_603,N_595,N_447);
and U604 (N_604,N_555,N_469);
or U605 (N_605,N_516,N_463);
xnor U606 (N_606,N_464,N_565);
and U607 (N_607,N_404,N_494);
xor U608 (N_608,N_591,N_432);
and U609 (N_609,N_513,N_486);
nand U610 (N_610,N_476,N_575);
or U611 (N_611,N_521,N_512);
and U612 (N_612,N_519,N_431);
nor U613 (N_613,N_551,N_526);
nand U614 (N_614,N_539,N_462);
xnor U615 (N_615,N_472,N_449);
nand U616 (N_616,N_505,N_443);
and U617 (N_617,N_497,N_423);
xnor U618 (N_618,N_531,N_491);
or U619 (N_619,N_564,N_503);
nor U620 (N_620,N_540,N_502);
nand U621 (N_621,N_499,N_451);
nand U622 (N_622,N_584,N_461);
nor U623 (N_623,N_434,N_446);
and U624 (N_624,N_485,N_559);
xor U625 (N_625,N_573,N_506);
nand U626 (N_626,N_574,N_470);
and U627 (N_627,N_542,N_533);
nand U628 (N_628,N_546,N_422);
nand U629 (N_629,N_481,N_560);
nor U630 (N_630,N_527,N_593);
or U631 (N_631,N_545,N_419);
nor U632 (N_632,N_554,N_567);
nor U633 (N_633,N_571,N_406);
nor U634 (N_634,N_590,N_484);
nor U635 (N_635,N_430,N_458);
nand U636 (N_636,N_488,N_558);
nand U637 (N_637,N_568,N_493);
and U638 (N_638,N_475,N_489);
and U639 (N_639,N_599,N_410);
xor U640 (N_640,N_413,N_587);
nand U641 (N_641,N_570,N_433);
nor U642 (N_642,N_492,N_547);
or U643 (N_643,N_425,N_408);
xor U644 (N_644,N_468,N_466);
and U645 (N_645,N_411,N_594);
and U646 (N_646,N_455,N_509);
or U647 (N_647,N_403,N_498);
and U648 (N_648,N_482,N_460);
nor U649 (N_649,N_417,N_524);
xor U650 (N_650,N_578,N_483);
nand U651 (N_651,N_579,N_532);
nor U652 (N_652,N_517,N_566);
or U653 (N_653,N_454,N_550);
and U654 (N_654,N_523,N_474);
or U655 (N_655,N_589,N_445);
xnor U656 (N_656,N_427,N_514);
and U657 (N_657,N_522,N_543);
and U658 (N_658,N_416,N_437);
or U659 (N_659,N_597,N_452);
and U660 (N_660,N_473,N_538);
xor U661 (N_661,N_412,N_561);
or U662 (N_662,N_467,N_402);
xor U663 (N_663,N_400,N_401);
nand U664 (N_664,N_453,N_508);
xor U665 (N_665,N_448,N_577);
nand U666 (N_666,N_520,N_471);
and U667 (N_667,N_439,N_588);
xor U668 (N_668,N_572,N_480);
xnor U669 (N_669,N_465,N_511);
nor U670 (N_670,N_442,N_581);
and U671 (N_671,N_429,N_459);
and U672 (N_672,N_507,N_510);
nand U673 (N_673,N_528,N_501);
nor U674 (N_674,N_487,N_592);
nor U675 (N_675,N_549,N_421);
and U676 (N_676,N_435,N_418);
nor U677 (N_677,N_537,N_407);
nor U678 (N_678,N_426,N_585);
nor U679 (N_679,N_440,N_548);
or U680 (N_680,N_518,N_436);
nand U681 (N_681,N_553,N_534);
and U682 (N_682,N_569,N_456);
nand U683 (N_683,N_580,N_444);
and U684 (N_684,N_441,N_479);
nor U685 (N_685,N_541,N_428);
and U686 (N_686,N_535,N_525);
xnor U687 (N_687,N_409,N_495);
and U688 (N_688,N_582,N_477);
xor U689 (N_689,N_586,N_596);
or U690 (N_690,N_515,N_598);
and U691 (N_691,N_576,N_490);
nor U692 (N_692,N_478,N_544);
xnor U693 (N_693,N_583,N_530);
xor U694 (N_694,N_556,N_420);
or U695 (N_695,N_415,N_500);
xor U696 (N_696,N_504,N_529);
nor U697 (N_697,N_438,N_424);
and U698 (N_698,N_414,N_496);
nor U699 (N_699,N_552,N_405);
or U700 (N_700,N_535,N_586);
or U701 (N_701,N_503,N_514);
nor U702 (N_702,N_517,N_583);
nor U703 (N_703,N_569,N_467);
or U704 (N_704,N_562,N_483);
xnor U705 (N_705,N_527,N_567);
nor U706 (N_706,N_467,N_583);
xor U707 (N_707,N_417,N_505);
nand U708 (N_708,N_556,N_456);
nand U709 (N_709,N_427,N_556);
xnor U710 (N_710,N_426,N_474);
and U711 (N_711,N_473,N_557);
nor U712 (N_712,N_473,N_475);
xnor U713 (N_713,N_426,N_495);
or U714 (N_714,N_404,N_496);
nor U715 (N_715,N_512,N_548);
nand U716 (N_716,N_484,N_428);
nand U717 (N_717,N_523,N_479);
nand U718 (N_718,N_598,N_457);
and U719 (N_719,N_510,N_485);
or U720 (N_720,N_554,N_452);
nand U721 (N_721,N_566,N_565);
and U722 (N_722,N_450,N_597);
nand U723 (N_723,N_572,N_502);
xor U724 (N_724,N_573,N_481);
or U725 (N_725,N_431,N_522);
xor U726 (N_726,N_556,N_466);
nand U727 (N_727,N_439,N_535);
xnor U728 (N_728,N_403,N_495);
nor U729 (N_729,N_463,N_507);
nand U730 (N_730,N_432,N_568);
nor U731 (N_731,N_436,N_421);
nand U732 (N_732,N_421,N_495);
xnor U733 (N_733,N_483,N_527);
xnor U734 (N_734,N_525,N_509);
or U735 (N_735,N_425,N_585);
xor U736 (N_736,N_421,N_596);
nor U737 (N_737,N_560,N_500);
xor U738 (N_738,N_597,N_580);
xor U739 (N_739,N_547,N_465);
nor U740 (N_740,N_450,N_479);
or U741 (N_741,N_475,N_514);
or U742 (N_742,N_531,N_565);
nand U743 (N_743,N_542,N_477);
or U744 (N_744,N_577,N_403);
nand U745 (N_745,N_475,N_465);
xor U746 (N_746,N_498,N_437);
nor U747 (N_747,N_455,N_477);
and U748 (N_748,N_536,N_429);
xor U749 (N_749,N_503,N_480);
or U750 (N_750,N_562,N_464);
xnor U751 (N_751,N_482,N_496);
nand U752 (N_752,N_435,N_568);
xor U753 (N_753,N_567,N_437);
nand U754 (N_754,N_412,N_422);
or U755 (N_755,N_448,N_486);
and U756 (N_756,N_453,N_470);
and U757 (N_757,N_586,N_471);
nor U758 (N_758,N_531,N_452);
xor U759 (N_759,N_412,N_585);
and U760 (N_760,N_558,N_460);
nand U761 (N_761,N_441,N_581);
xnor U762 (N_762,N_476,N_431);
nand U763 (N_763,N_599,N_564);
nand U764 (N_764,N_572,N_526);
nand U765 (N_765,N_549,N_528);
xor U766 (N_766,N_516,N_417);
and U767 (N_767,N_519,N_567);
and U768 (N_768,N_563,N_586);
and U769 (N_769,N_440,N_499);
or U770 (N_770,N_587,N_523);
xnor U771 (N_771,N_455,N_430);
or U772 (N_772,N_464,N_575);
nor U773 (N_773,N_419,N_404);
nor U774 (N_774,N_438,N_531);
or U775 (N_775,N_558,N_474);
xnor U776 (N_776,N_441,N_460);
and U777 (N_777,N_528,N_568);
or U778 (N_778,N_484,N_586);
and U779 (N_779,N_458,N_528);
nand U780 (N_780,N_418,N_553);
or U781 (N_781,N_485,N_411);
or U782 (N_782,N_496,N_451);
nand U783 (N_783,N_408,N_517);
or U784 (N_784,N_404,N_565);
nor U785 (N_785,N_436,N_574);
xnor U786 (N_786,N_567,N_560);
nand U787 (N_787,N_488,N_466);
nor U788 (N_788,N_524,N_588);
or U789 (N_789,N_420,N_529);
or U790 (N_790,N_540,N_583);
and U791 (N_791,N_502,N_568);
and U792 (N_792,N_593,N_563);
and U793 (N_793,N_448,N_569);
and U794 (N_794,N_457,N_514);
xor U795 (N_795,N_555,N_592);
or U796 (N_796,N_402,N_473);
xnor U797 (N_797,N_587,N_535);
nor U798 (N_798,N_583,N_500);
nor U799 (N_799,N_411,N_582);
or U800 (N_800,N_604,N_649);
or U801 (N_801,N_639,N_626);
xnor U802 (N_802,N_719,N_627);
xor U803 (N_803,N_684,N_710);
and U804 (N_804,N_711,N_721);
nor U805 (N_805,N_751,N_686);
nand U806 (N_806,N_635,N_747);
xor U807 (N_807,N_652,N_718);
nor U808 (N_808,N_630,N_621);
or U809 (N_809,N_727,N_674);
or U810 (N_810,N_605,N_760);
xnor U811 (N_811,N_603,N_645);
and U812 (N_812,N_632,N_682);
nor U813 (N_813,N_778,N_799);
and U814 (N_814,N_772,N_690);
nor U815 (N_815,N_651,N_646);
xnor U816 (N_816,N_687,N_717);
and U817 (N_817,N_636,N_714);
nor U818 (N_818,N_601,N_625);
or U819 (N_819,N_709,N_666);
nor U820 (N_820,N_609,N_620);
nand U821 (N_821,N_607,N_697);
nand U822 (N_822,N_768,N_771);
and U823 (N_823,N_704,N_654);
or U824 (N_824,N_624,N_776);
and U825 (N_825,N_758,N_733);
nor U826 (N_826,N_715,N_696);
xor U827 (N_827,N_629,N_694);
and U828 (N_828,N_740,N_613);
and U829 (N_829,N_611,N_642);
and U830 (N_830,N_700,N_689);
or U831 (N_831,N_648,N_769);
xnor U832 (N_832,N_765,N_600);
xor U833 (N_833,N_670,N_790);
and U834 (N_834,N_617,N_643);
nor U835 (N_835,N_728,N_671);
nand U836 (N_836,N_789,N_680);
nand U837 (N_837,N_614,N_702);
nand U838 (N_838,N_698,N_623);
and U839 (N_839,N_631,N_742);
nor U840 (N_840,N_754,N_779);
or U841 (N_841,N_663,N_783);
xor U842 (N_842,N_762,N_657);
nand U843 (N_843,N_693,N_734);
or U844 (N_844,N_798,N_707);
and U845 (N_845,N_679,N_766);
or U846 (N_846,N_659,N_767);
or U847 (N_847,N_781,N_640);
nand U848 (N_848,N_763,N_622);
nor U849 (N_849,N_616,N_720);
xnor U850 (N_850,N_761,N_786);
or U851 (N_851,N_729,N_793);
or U852 (N_852,N_699,N_644);
nor U853 (N_853,N_775,N_759);
nand U854 (N_854,N_750,N_658);
xor U855 (N_855,N_724,N_665);
nor U856 (N_856,N_764,N_730);
and U857 (N_857,N_712,N_661);
nand U858 (N_858,N_777,N_726);
xor U859 (N_859,N_664,N_692);
xor U860 (N_860,N_749,N_606);
nand U861 (N_861,N_637,N_773);
and U862 (N_862,N_695,N_703);
nand U863 (N_863,N_675,N_770);
nand U864 (N_864,N_673,N_784);
xnor U865 (N_865,N_797,N_746);
nor U866 (N_866,N_676,N_701);
and U867 (N_867,N_787,N_745);
or U868 (N_868,N_685,N_757);
nand U869 (N_869,N_756,N_708);
xor U870 (N_870,N_633,N_780);
or U871 (N_871,N_634,N_653);
nor U872 (N_872,N_656,N_788);
nand U873 (N_873,N_610,N_796);
xnor U874 (N_874,N_608,N_736);
nand U875 (N_875,N_792,N_641);
and U876 (N_876,N_737,N_638);
or U877 (N_877,N_713,N_619);
xor U878 (N_878,N_755,N_739);
nand U879 (N_879,N_735,N_743);
and U880 (N_880,N_774,N_794);
nor U881 (N_881,N_785,N_612);
and U882 (N_882,N_691,N_723);
nor U883 (N_883,N_677,N_602);
nor U884 (N_884,N_722,N_782);
nor U885 (N_885,N_615,N_662);
and U886 (N_886,N_795,N_748);
xor U887 (N_887,N_725,N_705);
xnor U888 (N_888,N_706,N_752);
or U889 (N_889,N_647,N_738);
and U890 (N_890,N_753,N_731);
nand U891 (N_891,N_688,N_683);
or U892 (N_892,N_628,N_681);
xor U893 (N_893,N_650,N_741);
xor U894 (N_894,N_678,N_669);
nand U895 (N_895,N_667,N_744);
nand U896 (N_896,N_655,N_716);
xnor U897 (N_897,N_672,N_791);
and U898 (N_898,N_660,N_732);
and U899 (N_899,N_618,N_668);
xnor U900 (N_900,N_717,N_702);
and U901 (N_901,N_654,N_768);
or U902 (N_902,N_686,N_780);
nor U903 (N_903,N_626,N_798);
or U904 (N_904,N_792,N_771);
nor U905 (N_905,N_605,N_658);
nor U906 (N_906,N_691,N_656);
xnor U907 (N_907,N_744,N_665);
nor U908 (N_908,N_603,N_731);
nand U909 (N_909,N_614,N_751);
or U910 (N_910,N_729,N_768);
nand U911 (N_911,N_636,N_644);
or U912 (N_912,N_636,N_745);
xor U913 (N_913,N_740,N_610);
nor U914 (N_914,N_650,N_707);
nor U915 (N_915,N_626,N_661);
nand U916 (N_916,N_732,N_685);
nand U917 (N_917,N_755,N_721);
nand U918 (N_918,N_729,N_638);
nand U919 (N_919,N_615,N_665);
nor U920 (N_920,N_695,N_772);
and U921 (N_921,N_602,N_718);
nand U922 (N_922,N_748,N_651);
nand U923 (N_923,N_653,N_658);
nand U924 (N_924,N_720,N_769);
nand U925 (N_925,N_786,N_660);
or U926 (N_926,N_684,N_731);
xnor U927 (N_927,N_780,N_672);
or U928 (N_928,N_766,N_618);
nor U929 (N_929,N_652,N_621);
xor U930 (N_930,N_632,N_755);
nand U931 (N_931,N_792,N_756);
xor U932 (N_932,N_773,N_715);
and U933 (N_933,N_615,N_795);
nand U934 (N_934,N_773,N_731);
and U935 (N_935,N_620,N_671);
or U936 (N_936,N_655,N_745);
xor U937 (N_937,N_771,N_655);
nand U938 (N_938,N_705,N_661);
or U939 (N_939,N_674,N_661);
nor U940 (N_940,N_758,N_790);
nor U941 (N_941,N_699,N_739);
xnor U942 (N_942,N_794,N_662);
nor U943 (N_943,N_797,N_702);
xnor U944 (N_944,N_682,N_640);
or U945 (N_945,N_755,N_744);
or U946 (N_946,N_756,N_787);
and U947 (N_947,N_643,N_603);
or U948 (N_948,N_780,N_764);
and U949 (N_949,N_740,N_794);
nand U950 (N_950,N_728,N_663);
nor U951 (N_951,N_712,N_771);
nor U952 (N_952,N_607,N_757);
and U953 (N_953,N_694,N_677);
and U954 (N_954,N_763,N_724);
or U955 (N_955,N_676,N_620);
nand U956 (N_956,N_601,N_789);
and U957 (N_957,N_644,N_609);
and U958 (N_958,N_652,N_793);
nor U959 (N_959,N_731,N_620);
nand U960 (N_960,N_759,N_612);
nand U961 (N_961,N_630,N_775);
or U962 (N_962,N_761,N_700);
xnor U963 (N_963,N_790,N_794);
or U964 (N_964,N_769,N_733);
nor U965 (N_965,N_614,N_631);
or U966 (N_966,N_710,N_678);
and U967 (N_967,N_725,N_626);
nor U968 (N_968,N_658,N_681);
xnor U969 (N_969,N_790,N_750);
nand U970 (N_970,N_735,N_637);
and U971 (N_971,N_728,N_618);
xor U972 (N_972,N_688,N_725);
and U973 (N_973,N_706,N_605);
nor U974 (N_974,N_676,N_690);
nor U975 (N_975,N_797,N_775);
nand U976 (N_976,N_769,N_647);
and U977 (N_977,N_796,N_793);
nand U978 (N_978,N_794,N_622);
xnor U979 (N_979,N_621,N_725);
and U980 (N_980,N_722,N_675);
nor U981 (N_981,N_722,N_756);
nor U982 (N_982,N_785,N_761);
nor U983 (N_983,N_624,N_685);
xnor U984 (N_984,N_757,N_651);
or U985 (N_985,N_745,N_703);
nand U986 (N_986,N_624,N_698);
and U987 (N_987,N_693,N_740);
nand U988 (N_988,N_682,N_742);
and U989 (N_989,N_736,N_640);
nor U990 (N_990,N_737,N_682);
and U991 (N_991,N_787,N_717);
and U992 (N_992,N_782,N_612);
or U993 (N_993,N_728,N_710);
and U994 (N_994,N_732,N_650);
nor U995 (N_995,N_755,N_643);
nand U996 (N_996,N_723,N_708);
and U997 (N_997,N_674,N_731);
xnor U998 (N_998,N_754,N_726);
nand U999 (N_999,N_789,N_646);
or U1000 (N_1000,N_811,N_855);
and U1001 (N_1001,N_828,N_950);
nor U1002 (N_1002,N_841,N_952);
or U1003 (N_1003,N_998,N_884);
or U1004 (N_1004,N_853,N_906);
nand U1005 (N_1005,N_809,N_901);
xnor U1006 (N_1006,N_885,N_951);
or U1007 (N_1007,N_890,N_991);
xor U1008 (N_1008,N_942,N_963);
nand U1009 (N_1009,N_891,N_915);
nor U1010 (N_1010,N_807,N_983);
nor U1011 (N_1011,N_817,N_808);
or U1012 (N_1012,N_824,N_994);
or U1013 (N_1013,N_815,N_843);
and U1014 (N_1014,N_837,N_802);
or U1015 (N_1015,N_813,N_989);
or U1016 (N_1016,N_956,N_936);
xnor U1017 (N_1017,N_996,N_872);
and U1018 (N_1018,N_973,N_875);
xnor U1019 (N_1019,N_964,N_909);
xor U1020 (N_1020,N_858,N_982);
or U1021 (N_1021,N_836,N_866);
xor U1022 (N_1022,N_854,N_831);
xnor U1023 (N_1023,N_948,N_887);
xor U1024 (N_1024,N_870,N_834);
or U1025 (N_1025,N_900,N_864);
or U1026 (N_1026,N_993,N_894);
or U1027 (N_1027,N_877,N_842);
and U1028 (N_1028,N_911,N_937);
nand U1029 (N_1029,N_908,N_981);
and U1030 (N_1030,N_878,N_932);
and U1031 (N_1031,N_905,N_988);
xor U1032 (N_1032,N_869,N_886);
xnor U1033 (N_1033,N_959,N_880);
and U1034 (N_1034,N_962,N_957);
nand U1035 (N_1035,N_926,N_997);
nor U1036 (N_1036,N_992,N_873);
nor U1037 (N_1037,N_918,N_897);
nand U1038 (N_1038,N_883,N_966);
nor U1039 (N_1039,N_907,N_979);
or U1040 (N_1040,N_969,N_844);
and U1041 (N_1041,N_949,N_984);
and U1042 (N_1042,N_889,N_960);
and U1043 (N_1043,N_987,N_925);
and U1044 (N_1044,N_941,N_999);
xor U1045 (N_1045,N_975,N_840);
or U1046 (N_1046,N_835,N_803);
nor U1047 (N_1047,N_972,N_946);
or U1048 (N_1048,N_939,N_851);
and U1049 (N_1049,N_862,N_839);
or U1050 (N_1050,N_893,N_967);
xor U1051 (N_1051,N_825,N_895);
nor U1052 (N_1052,N_871,N_856);
xnor U1053 (N_1053,N_974,N_954);
and U1054 (N_1054,N_913,N_977);
or U1055 (N_1055,N_899,N_976);
and U1056 (N_1056,N_971,N_921);
nor U1057 (N_1057,N_929,N_985);
xor U1058 (N_1058,N_814,N_879);
or U1059 (N_1059,N_916,N_859);
and U1060 (N_1060,N_865,N_953);
xor U1061 (N_1061,N_848,N_849);
and U1062 (N_1062,N_904,N_945);
nand U1063 (N_1063,N_930,N_898);
xor U1064 (N_1064,N_830,N_892);
nand U1065 (N_1065,N_846,N_923);
xor U1066 (N_1066,N_876,N_838);
xnor U1067 (N_1067,N_933,N_882);
xnor U1068 (N_1068,N_990,N_812);
nor U1069 (N_1069,N_938,N_819);
and U1070 (N_1070,N_832,N_968);
and U1071 (N_1071,N_917,N_896);
or U1072 (N_1072,N_850,N_910);
xnor U1073 (N_1073,N_881,N_804);
nand U1074 (N_1074,N_903,N_829);
xor U1075 (N_1075,N_940,N_995);
and U1076 (N_1076,N_931,N_800);
nand U1077 (N_1077,N_818,N_970);
xnor U1078 (N_1078,N_826,N_861);
nor U1079 (N_1079,N_833,N_863);
and U1080 (N_1080,N_822,N_944);
or U1081 (N_1081,N_806,N_927);
and U1082 (N_1082,N_943,N_847);
or U1083 (N_1083,N_857,N_821);
nor U1084 (N_1084,N_978,N_888);
or U1085 (N_1085,N_852,N_955);
xor U1086 (N_1086,N_919,N_823);
or U1087 (N_1087,N_935,N_827);
and U1088 (N_1088,N_914,N_868);
or U1089 (N_1089,N_874,N_947);
xnor U1090 (N_1090,N_920,N_986);
or U1091 (N_1091,N_867,N_860);
nand U1092 (N_1092,N_928,N_980);
nor U1093 (N_1093,N_912,N_810);
xnor U1094 (N_1094,N_922,N_805);
or U1095 (N_1095,N_801,N_961);
nand U1096 (N_1096,N_924,N_902);
and U1097 (N_1097,N_934,N_845);
nand U1098 (N_1098,N_816,N_965);
or U1099 (N_1099,N_820,N_958);
or U1100 (N_1100,N_833,N_812);
nand U1101 (N_1101,N_856,N_852);
nor U1102 (N_1102,N_934,N_854);
or U1103 (N_1103,N_993,N_918);
nand U1104 (N_1104,N_932,N_928);
and U1105 (N_1105,N_952,N_969);
xor U1106 (N_1106,N_810,N_915);
xnor U1107 (N_1107,N_816,N_828);
or U1108 (N_1108,N_837,N_906);
nand U1109 (N_1109,N_862,N_944);
nand U1110 (N_1110,N_916,N_810);
xnor U1111 (N_1111,N_800,N_916);
or U1112 (N_1112,N_864,N_807);
or U1113 (N_1113,N_930,N_890);
nor U1114 (N_1114,N_927,N_895);
and U1115 (N_1115,N_881,N_883);
xor U1116 (N_1116,N_978,N_819);
nor U1117 (N_1117,N_915,N_852);
and U1118 (N_1118,N_896,N_821);
xor U1119 (N_1119,N_996,N_904);
nand U1120 (N_1120,N_807,N_977);
nand U1121 (N_1121,N_810,N_909);
nor U1122 (N_1122,N_860,N_832);
nand U1123 (N_1123,N_864,N_840);
and U1124 (N_1124,N_953,N_990);
nand U1125 (N_1125,N_879,N_980);
nor U1126 (N_1126,N_821,N_906);
nand U1127 (N_1127,N_997,N_859);
or U1128 (N_1128,N_812,N_927);
or U1129 (N_1129,N_939,N_910);
and U1130 (N_1130,N_866,N_910);
and U1131 (N_1131,N_827,N_943);
or U1132 (N_1132,N_993,N_890);
xor U1133 (N_1133,N_871,N_980);
xnor U1134 (N_1134,N_981,N_800);
nand U1135 (N_1135,N_991,N_809);
or U1136 (N_1136,N_940,N_919);
xor U1137 (N_1137,N_891,N_992);
and U1138 (N_1138,N_932,N_982);
nand U1139 (N_1139,N_849,N_934);
nand U1140 (N_1140,N_953,N_975);
xor U1141 (N_1141,N_881,N_935);
or U1142 (N_1142,N_886,N_953);
or U1143 (N_1143,N_859,N_927);
or U1144 (N_1144,N_879,N_851);
and U1145 (N_1145,N_817,N_802);
nand U1146 (N_1146,N_974,N_903);
and U1147 (N_1147,N_859,N_894);
nor U1148 (N_1148,N_813,N_925);
nand U1149 (N_1149,N_865,N_895);
xnor U1150 (N_1150,N_839,N_899);
nand U1151 (N_1151,N_943,N_912);
and U1152 (N_1152,N_877,N_999);
and U1153 (N_1153,N_928,N_961);
nand U1154 (N_1154,N_824,N_874);
or U1155 (N_1155,N_864,N_841);
nor U1156 (N_1156,N_803,N_982);
or U1157 (N_1157,N_874,N_867);
and U1158 (N_1158,N_976,N_857);
xor U1159 (N_1159,N_890,N_997);
xnor U1160 (N_1160,N_864,N_814);
xor U1161 (N_1161,N_844,N_954);
nor U1162 (N_1162,N_843,N_976);
nand U1163 (N_1163,N_990,N_833);
or U1164 (N_1164,N_808,N_803);
nand U1165 (N_1165,N_981,N_933);
xnor U1166 (N_1166,N_960,N_829);
nor U1167 (N_1167,N_962,N_851);
xor U1168 (N_1168,N_904,N_813);
nand U1169 (N_1169,N_888,N_899);
and U1170 (N_1170,N_904,N_868);
xor U1171 (N_1171,N_881,N_877);
nand U1172 (N_1172,N_961,N_902);
or U1173 (N_1173,N_862,N_865);
or U1174 (N_1174,N_812,N_933);
and U1175 (N_1175,N_823,N_993);
or U1176 (N_1176,N_810,N_817);
and U1177 (N_1177,N_857,N_907);
nand U1178 (N_1178,N_908,N_801);
nor U1179 (N_1179,N_807,N_870);
or U1180 (N_1180,N_849,N_827);
or U1181 (N_1181,N_940,N_804);
and U1182 (N_1182,N_811,N_902);
or U1183 (N_1183,N_930,N_997);
or U1184 (N_1184,N_819,N_855);
xor U1185 (N_1185,N_921,N_970);
and U1186 (N_1186,N_945,N_847);
and U1187 (N_1187,N_845,N_969);
nor U1188 (N_1188,N_842,N_807);
nor U1189 (N_1189,N_966,N_832);
xnor U1190 (N_1190,N_902,N_870);
xor U1191 (N_1191,N_995,N_833);
nor U1192 (N_1192,N_962,N_816);
xor U1193 (N_1193,N_933,N_986);
or U1194 (N_1194,N_880,N_812);
and U1195 (N_1195,N_847,N_864);
and U1196 (N_1196,N_938,N_810);
and U1197 (N_1197,N_907,N_839);
nand U1198 (N_1198,N_930,N_842);
xnor U1199 (N_1199,N_965,N_958);
and U1200 (N_1200,N_1005,N_1167);
nand U1201 (N_1201,N_1094,N_1082);
xnor U1202 (N_1202,N_1161,N_1027);
and U1203 (N_1203,N_1089,N_1095);
nand U1204 (N_1204,N_1121,N_1189);
nor U1205 (N_1205,N_1063,N_1130);
nor U1206 (N_1206,N_1012,N_1080);
xnor U1207 (N_1207,N_1026,N_1060);
nor U1208 (N_1208,N_1004,N_1133);
nor U1209 (N_1209,N_1062,N_1152);
and U1210 (N_1210,N_1081,N_1172);
xnor U1211 (N_1211,N_1144,N_1074);
and U1212 (N_1212,N_1156,N_1091);
nor U1213 (N_1213,N_1165,N_1170);
xor U1214 (N_1214,N_1149,N_1131);
nor U1215 (N_1215,N_1146,N_1096);
or U1216 (N_1216,N_1021,N_1070);
nand U1217 (N_1217,N_1101,N_1104);
nand U1218 (N_1218,N_1051,N_1097);
xor U1219 (N_1219,N_1187,N_1196);
and U1220 (N_1220,N_1056,N_1134);
nor U1221 (N_1221,N_1046,N_1160);
nor U1222 (N_1222,N_1129,N_1043);
nor U1223 (N_1223,N_1117,N_1092);
and U1224 (N_1224,N_1183,N_1000);
nand U1225 (N_1225,N_1015,N_1166);
nand U1226 (N_1226,N_1078,N_1035);
and U1227 (N_1227,N_1020,N_1148);
and U1228 (N_1228,N_1181,N_1164);
nand U1229 (N_1229,N_1052,N_1143);
and U1230 (N_1230,N_1186,N_1023);
and U1231 (N_1231,N_1112,N_1184);
nand U1232 (N_1232,N_1190,N_1169);
nor U1233 (N_1233,N_1029,N_1139);
nor U1234 (N_1234,N_1028,N_1055);
and U1235 (N_1235,N_1113,N_1107);
nor U1236 (N_1236,N_1102,N_1039);
xnor U1237 (N_1237,N_1177,N_1013);
or U1238 (N_1238,N_1114,N_1014);
nor U1239 (N_1239,N_1158,N_1150);
xnor U1240 (N_1240,N_1022,N_1175);
and U1241 (N_1241,N_1120,N_1067);
nand U1242 (N_1242,N_1198,N_1058);
xnor U1243 (N_1243,N_1025,N_1006);
nand U1244 (N_1244,N_1191,N_1194);
xnor U1245 (N_1245,N_1118,N_1088);
xnor U1246 (N_1246,N_1066,N_1093);
nor U1247 (N_1247,N_1009,N_1098);
nor U1248 (N_1248,N_1197,N_1003);
or U1249 (N_1249,N_1122,N_1071);
xor U1250 (N_1250,N_1064,N_1072);
or U1251 (N_1251,N_1044,N_1192);
nor U1252 (N_1252,N_1145,N_1157);
nand U1253 (N_1253,N_1036,N_1171);
xor U1254 (N_1254,N_1077,N_1049);
and U1255 (N_1255,N_1059,N_1135);
or U1256 (N_1256,N_1011,N_1193);
nor U1257 (N_1257,N_1109,N_1075);
or U1258 (N_1258,N_1178,N_1034);
xnor U1259 (N_1259,N_1085,N_1084);
xnor U1260 (N_1260,N_1155,N_1017);
xor U1261 (N_1261,N_1111,N_1147);
xor U1262 (N_1262,N_1176,N_1045);
or U1263 (N_1263,N_1151,N_1108);
nor U1264 (N_1264,N_1116,N_1179);
xnor U1265 (N_1265,N_1105,N_1128);
nor U1266 (N_1266,N_1119,N_1032);
or U1267 (N_1267,N_1068,N_1076);
nand U1268 (N_1268,N_1168,N_1086);
nor U1269 (N_1269,N_1061,N_1053);
nor U1270 (N_1270,N_1069,N_1001);
xor U1271 (N_1271,N_1138,N_1031);
and U1272 (N_1272,N_1030,N_1037);
nor U1273 (N_1273,N_1123,N_1048);
and U1274 (N_1274,N_1174,N_1136);
or U1275 (N_1275,N_1008,N_1195);
xor U1276 (N_1276,N_1162,N_1038);
nand U1277 (N_1277,N_1154,N_1173);
nor U1278 (N_1278,N_1033,N_1040);
or U1279 (N_1279,N_1159,N_1050);
xor U1280 (N_1280,N_1137,N_1057);
xnor U1281 (N_1281,N_1103,N_1110);
and U1282 (N_1282,N_1132,N_1007);
nor U1283 (N_1283,N_1087,N_1054);
xor U1284 (N_1284,N_1106,N_1019);
and U1285 (N_1285,N_1100,N_1199);
nand U1286 (N_1286,N_1024,N_1126);
nand U1287 (N_1287,N_1041,N_1163);
nor U1288 (N_1288,N_1180,N_1185);
or U1289 (N_1289,N_1083,N_1016);
nand U1290 (N_1290,N_1124,N_1099);
nor U1291 (N_1291,N_1188,N_1141);
nand U1292 (N_1292,N_1182,N_1073);
or U1293 (N_1293,N_1065,N_1153);
and U1294 (N_1294,N_1018,N_1140);
nand U1295 (N_1295,N_1142,N_1115);
xor U1296 (N_1296,N_1079,N_1002);
nor U1297 (N_1297,N_1010,N_1090);
nand U1298 (N_1298,N_1042,N_1047);
nor U1299 (N_1299,N_1127,N_1125);
nand U1300 (N_1300,N_1056,N_1065);
or U1301 (N_1301,N_1063,N_1016);
and U1302 (N_1302,N_1044,N_1061);
nand U1303 (N_1303,N_1104,N_1183);
xor U1304 (N_1304,N_1167,N_1120);
nand U1305 (N_1305,N_1049,N_1162);
nand U1306 (N_1306,N_1050,N_1109);
or U1307 (N_1307,N_1156,N_1074);
xor U1308 (N_1308,N_1055,N_1112);
nor U1309 (N_1309,N_1071,N_1188);
or U1310 (N_1310,N_1184,N_1100);
and U1311 (N_1311,N_1116,N_1071);
nor U1312 (N_1312,N_1000,N_1006);
and U1313 (N_1313,N_1021,N_1029);
xnor U1314 (N_1314,N_1016,N_1103);
and U1315 (N_1315,N_1182,N_1181);
or U1316 (N_1316,N_1194,N_1199);
nand U1317 (N_1317,N_1089,N_1144);
or U1318 (N_1318,N_1123,N_1076);
nand U1319 (N_1319,N_1011,N_1149);
and U1320 (N_1320,N_1180,N_1057);
xor U1321 (N_1321,N_1032,N_1012);
nand U1322 (N_1322,N_1168,N_1087);
xnor U1323 (N_1323,N_1045,N_1169);
or U1324 (N_1324,N_1168,N_1164);
and U1325 (N_1325,N_1109,N_1184);
nor U1326 (N_1326,N_1124,N_1173);
nor U1327 (N_1327,N_1151,N_1195);
or U1328 (N_1328,N_1117,N_1168);
xor U1329 (N_1329,N_1129,N_1127);
and U1330 (N_1330,N_1003,N_1112);
nor U1331 (N_1331,N_1182,N_1107);
nand U1332 (N_1332,N_1180,N_1122);
and U1333 (N_1333,N_1184,N_1165);
nand U1334 (N_1334,N_1007,N_1042);
nand U1335 (N_1335,N_1028,N_1129);
or U1336 (N_1336,N_1007,N_1061);
and U1337 (N_1337,N_1007,N_1050);
or U1338 (N_1338,N_1099,N_1122);
xnor U1339 (N_1339,N_1110,N_1152);
nor U1340 (N_1340,N_1140,N_1175);
or U1341 (N_1341,N_1186,N_1181);
nand U1342 (N_1342,N_1120,N_1156);
xnor U1343 (N_1343,N_1123,N_1065);
and U1344 (N_1344,N_1091,N_1161);
or U1345 (N_1345,N_1084,N_1094);
and U1346 (N_1346,N_1127,N_1134);
nor U1347 (N_1347,N_1111,N_1067);
nor U1348 (N_1348,N_1146,N_1100);
and U1349 (N_1349,N_1155,N_1083);
and U1350 (N_1350,N_1009,N_1104);
or U1351 (N_1351,N_1060,N_1178);
and U1352 (N_1352,N_1194,N_1195);
xor U1353 (N_1353,N_1121,N_1079);
nor U1354 (N_1354,N_1159,N_1180);
nor U1355 (N_1355,N_1103,N_1184);
nand U1356 (N_1356,N_1019,N_1159);
and U1357 (N_1357,N_1144,N_1184);
and U1358 (N_1358,N_1074,N_1158);
nand U1359 (N_1359,N_1151,N_1019);
xor U1360 (N_1360,N_1037,N_1034);
nand U1361 (N_1361,N_1097,N_1035);
nor U1362 (N_1362,N_1064,N_1065);
and U1363 (N_1363,N_1068,N_1065);
and U1364 (N_1364,N_1094,N_1135);
or U1365 (N_1365,N_1102,N_1168);
or U1366 (N_1366,N_1128,N_1190);
nand U1367 (N_1367,N_1174,N_1126);
xnor U1368 (N_1368,N_1133,N_1050);
and U1369 (N_1369,N_1191,N_1106);
or U1370 (N_1370,N_1023,N_1063);
xnor U1371 (N_1371,N_1181,N_1142);
nor U1372 (N_1372,N_1012,N_1064);
and U1373 (N_1373,N_1167,N_1140);
or U1374 (N_1374,N_1108,N_1185);
or U1375 (N_1375,N_1149,N_1017);
nand U1376 (N_1376,N_1057,N_1010);
nand U1377 (N_1377,N_1043,N_1166);
and U1378 (N_1378,N_1193,N_1115);
xor U1379 (N_1379,N_1197,N_1057);
and U1380 (N_1380,N_1039,N_1053);
and U1381 (N_1381,N_1155,N_1172);
xor U1382 (N_1382,N_1086,N_1050);
and U1383 (N_1383,N_1121,N_1145);
nand U1384 (N_1384,N_1158,N_1138);
nor U1385 (N_1385,N_1136,N_1114);
nor U1386 (N_1386,N_1091,N_1012);
or U1387 (N_1387,N_1083,N_1069);
and U1388 (N_1388,N_1069,N_1179);
nor U1389 (N_1389,N_1000,N_1177);
nand U1390 (N_1390,N_1089,N_1127);
xnor U1391 (N_1391,N_1174,N_1020);
nor U1392 (N_1392,N_1151,N_1115);
nand U1393 (N_1393,N_1080,N_1024);
nor U1394 (N_1394,N_1176,N_1065);
nor U1395 (N_1395,N_1137,N_1122);
nand U1396 (N_1396,N_1181,N_1024);
and U1397 (N_1397,N_1110,N_1049);
nand U1398 (N_1398,N_1089,N_1031);
xnor U1399 (N_1399,N_1148,N_1022);
xnor U1400 (N_1400,N_1377,N_1261);
nor U1401 (N_1401,N_1226,N_1315);
or U1402 (N_1402,N_1249,N_1236);
or U1403 (N_1403,N_1318,N_1216);
nand U1404 (N_1404,N_1365,N_1282);
xnor U1405 (N_1405,N_1334,N_1296);
nor U1406 (N_1406,N_1392,N_1397);
xor U1407 (N_1407,N_1386,N_1217);
nor U1408 (N_1408,N_1263,N_1258);
xnor U1409 (N_1409,N_1265,N_1248);
xor U1410 (N_1410,N_1266,N_1300);
nand U1411 (N_1411,N_1328,N_1389);
nor U1412 (N_1412,N_1227,N_1311);
xor U1413 (N_1413,N_1352,N_1280);
or U1414 (N_1414,N_1205,N_1277);
nor U1415 (N_1415,N_1239,N_1388);
nand U1416 (N_1416,N_1324,N_1350);
or U1417 (N_1417,N_1333,N_1380);
xnor U1418 (N_1418,N_1243,N_1246);
xor U1419 (N_1419,N_1294,N_1213);
or U1420 (N_1420,N_1381,N_1279);
nor U1421 (N_1421,N_1370,N_1343);
xnor U1422 (N_1422,N_1252,N_1271);
xnor U1423 (N_1423,N_1367,N_1379);
or U1424 (N_1424,N_1375,N_1251);
xor U1425 (N_1425,N_1222,N_1206);
nor U1426 (N_1426,N_1341,N_1245);
nand U1427 (N_1427,N_1382,N_1360);
or U1428 (N_1428,N_1387,N_1313);
xor U1429 (N_1429,N_1396,N_1284);
and U1430 (N_1430,N_1372,N_1208);
nand U1431 (N_1431,N_1207,N_1302);
xnor U1432 (N_1432,N_1260,N_1393);
nor U1433 (N_1433,N_1257,N_1209);
and U1434 (N_1434,N_1204,N_1356);
and U1435 (N_1435,N_1308,N_1273);
or U1436 (N_1436,N_1342,N_1347);
or U1437 (N_1437,N_1286,N_1288);
nor U1438 (N_1438,N_1369,N_1210);
and U1439 (N_1439,N_1354,N_1361);
nand U1440 (N_1440,N_1358,N_1384);
nor U1441 (N_1441,N_1353,N_1211);
or U1442 (N_1442,N_1346,N_1394);
nor U1443 (N_1443,N_1229,N_1297);
xnor U1444 (N_1444,N_1330,N_1378);
and U1445 (N_1445,N_1366,N_1221);
nand U1446 (N_1446,N_1274,N_1233);
nand U1447 (N_1447,N_1348,N_1224);
or U1448 (N_1448,N_1368,N_1267);
nor U1449 (N_1449,N_1326,N_1242);
or U1450 (N_1450,N_1281,N_1305);
or U1451 (N_1451,N_1268,N_1276);
nor U1452 (N_1452,N_1383,N_1295);
xnor U1453 (N_1453,N_1374,N_1241);
and U1454 (N_1454,N_1201,N_1390);
nor U1455 (N_1455,N_1344,N_1345);
nand U1456 (N_1456,N_1373,N_1359);
nor U1457 (N_1457,N_1218,N_1214);
and U1458 (N_1458,N_1304,N_1220);
nor U1459 (N_1459,N_1203,N_1234);
nor U1460 (N_1460,N_1320,N_1325);
xnor U1461 (N_1461,N_1329,N_1293);
nor U1462 (N_1462,N_1255,N_1272);
xnor U1463 (N_1463,N_1339,N_1307);
xor U1464 (N_1464,N_1225,N_1289);
nor U1465 (N_1465,N_1259,N_1336);
nor U1466 (N_1466,N_1362,N_1303);
nand U1467 (N_1467,N_1299,N_1310);
and U1468 (N_1468,N_1364,N_1250);
nor U1469 (N_1469,N_1254,N_1327);
or U1470 (N_1470,N_1301,N_1235);
and U1471 (N_1471,N_1290,N_1212);
nand U1472 (N_1472,N_1363,N_1285);
nand U1473 (N_1473,N_1244,N_1230);
or U1474 (N_1474,N_1237,N_1316);
and U1475 (N_1475,N_1283,N_1287);
nand U1476 (N_1476,N_1232,N_1298);
and U1477 (N_1477,N_1275,N_1291);
and U1478 (N_1478,N_1231,N_1371);
or U1479 (N_1479,N_1357,N_1385);
nand U1480 (N_1480,N_1238,N_1331);
nand U1481 (N_1481,N_1351,N_1323);
or U1482 (N_1482,N_1309,N_1337);
or U1483 (N_1483,N_1398,N_1335);
and U1484 (N_1484,N_1306,N_1332);
nor U1485 (N_1485,N_1256,N_1269);
nor U1486 (N_1486,N_1322,N_1202);
xor U1487 (N_1487,N_1215,N_1219);
nor U1488 (N_1488,N_1262,N_1228);
nand U1489 (N_1489,N_1355,N_1395);
nor U1490 (N_1490,N_1314,N_1223);
xnor U1491 (N_1491,N_1319,N_1264);
nand U1492 (N_1492,N_1391,N_1270);
and U1493 (N_1493,N_1292,N_1338);
nand U1494 (N_1494,N_1312,N_1399);
or U1495 (N_1495,N_1247,N_1349);
and U1496 (N_1496,N_1253,N_1200);
and U1497 (N_1497,N_1278,N_1240);
and U1498 (N_1498,N_1376,N_1340);
and U1499 (N_1499,N_1321,N_1317);
nor U1500 (N_1500,N_1230,N_1304);
nand U1501 (N_1501,N_1266,N_1231);
nor U1502 (N_1502,N_1245,N_1265);
nand U1503 (N_1503,N_1223,N_1263);
nand U1504 (N_1504,N_1372,N_1302);
or U1505 (N_1505,N_1202,N_1289);
nor U1506 (N_1506,N_1261,N_1270);
xor U1507 (N_1507,N_1243,N_1362);
and U1508 (N_1508,N_1257,N_1304);
nand U1509 (N_1509,N_1293,N_1220);
and U1510 (N_1510,N_1298,N_1252);
nor U1511 (N_1511,N_1307,N_1230);
xnor U1512 (N_1512,N_1328,N_1279);
and U1513 (N_1513,N_1356,N_1395);
nor U1514 (N_1514,N_1271,N_1317);
xor U1515 (N_1515,N_1281,N_1380);
xor U1516 (N_1516,N_1280,N_1300);
or U1517 (N_1517,N_1324,N_1362);
nor U1518 (N_1518,N_1297,N_1330);
nor U1519 (N_1519,N_1368,N_1280);
nand U1520 (N_1520,N_1240,N_1203);
or U1521 (N_1521,N_1274,N_1360);
and U1522 (N_1522,N_1213,N_1291);
xnor U1523 (N_1523,N_1386,N_1364);
or U1524 (N_1524,N_1395,N_1239);
and U1525 (N_1525,N_1272,N_1269);
xnor U1526 (N_1526,N_1278,N_1203);
and U1527 (N_1527,N_1244,N_1213);
nand U1528 (N_1528,N_1263,N_1207);
xnor U1529 (N_1529,N_1310,N_1287);
or U1530 (N_1530,N_1398,N_1372);
and U1531 (N_1531,N_1298,N_1376);
xnor U1532 (N_1532,N_1247,N_1378);
nand U1533 (N_1533,N_1381,N_1387);
and U1534 (N_1534,N_1340,N_1369);
nor U1535 (N_1535,N_1228,N_1275);
or U1536 (N_1536,N_1221,N_1395);
or U1537 (N_1537,N_1222,N_1374);
xnor U1538 (N_1538,N_1223,N_1384);
and U1539 (N_1539,N_1224,N_1318);
and U1540 (N_1540,N_1219,N_1338);
nand U1541 (N_1541,N_1298,N_1239);
xor U1542 (N_1542,N_1325,N_1230);
and U1543 (N_1543,N_1216,N_1326);
xor U1544 (N_1544,N_1333,N_1250);
and U1545 (N_1545,N_1275,N_1346);
xor U1546 (N_1546,N_1386,N_1228);
and U1547 (N_1547,N_1275,N_1384);
or U1548 (N_1548,N_1262,N_1312);
xnor U1549 (N_1549,N_1390,N_1200);
and U1550 (N_1550,N_1233,N_1311);
nand U1551 (N_1551,N_1289,N_1267);
nor U1552 (N_1552,N_1239,N_1260);
nor U1553 (N_1553,N_1319,N_1265);
xor U1554 (N_1554,N_1347,N_1274);
xor U1555 (N_1555,N_1271,N_1227);
nand U1556 (N_1556,N_1294,N_1375);
xor U1557 (N_1557,N_1372,N_1292);
and U1558 (N_1558,N_1351,N_1264);
nand U1559 (N_1559,N_1247,N_1301);
nand U1560 (N_1560,N_1324,N_1394);
nor U1561 (N_1561,N_1342,N_1252);
nand U1562 (N_1562,N_1336,N_1386);
and U1563 (N_1563,N_1306,N_1203);
or U1564 (N_1564,N_1395,N_1203);
and U1565 (N_1565,N_1279,N_1283);
nand U1566 (N_1566,N_1295,N_1238);
xor U1567 (N_1567,N_1284,N_1296);
or U1568 (N_1568,N_1253,N_1281);
nor U1569 (N_1569,N_1360,N_1293);
or U1570 (N_1570,N_1392,N_1300);
xnor U1571 (N_1571,N_1387,N_1388);
or U1572 (N_1572,N_1314,N_1383);
or U1573 (N_1573,N_1308,N_1288);
or U1574 (N_1574,N_1313,N_1312);
and U1575 (N_1575,N_1304,N_1349);
xnor U1576 (N_1576,N_1396,N_1205);
nor U1577 (N_1577,N_1299,N_1351);
or U1578 (N_1578,N_1273,N_1346);
or U1579 (N_1579,N_1248,N_1254);
or U1580 (N_1580,N_1346,N_1368);
xnor U1581 (N_1581,N_1365,N_1268);
and U1582 (N_1582,N_1336,N_1245);
or U1583 (N_1583,N_1250,N_1241);
nor U1584 (N_1584,N_1221,N_1354);
and U1585 (N_1585,N_1308,N_1272);
nor U1586 (N_1586,N_1393,N_1392);
nand U1587 (N_1587,N_1266,N_1382);
nand U1588 (N_1588,N_1377,N_1287);
or U1589 (N_1589,N_1336,N_1319);
or U1590 (N_1590,N_1283,N_1282);
or U1591 (N_1591,N_1245,N_1217);
nand U1592 (N_1592,N_1281,N_1221);
nor U1593 (N_1593,N_1287,N_1247);
and U1594 (N_1594,N_1388,N_1215);
and U1595 (N_1595,N_1330,N_1375);
xnor U1596 (N_1596,N_1318,N_1304);
and U1597 (N_1597,N_1301,N_1312);
xor U1598 (N_1598,N_1356,N_1245);
nand U1599 (N_1599,N_1368,N_1333);
xnor U1600 (N_1600,N_1452,N_1401);
or U1601 (N_1601,N_1432,N_1462);
nand U1602 (N_1602,N_1423,N_1559);
xor U1603 (N_1603,N_1438,N_1589);
xor U1604 (N_1604,N_1417,N_1428);
or U1605 (N_1605,N_1416,N_1588);
and U1606 (N_1606,N_1485,N_1480);
nor U1607 (N_1607,N_1457,N_1421);
xor U1608 (N_1608,N_1530,N_1464);
xor U1609 (N_1609,N_1435,N_1590);
and U1610 (N_1610,N_1562,N_1498);
xnor U1611 (N_1611,N_1422,N_1502);
xnor U1612 (N_1612,N_1578,N_1490);
nand U1613 (N_1613,N_1459,N_1534);
or U1614 (N_1614,N_1571,N_1404);
and U1615 (N_1615,N_1493,N_1440);
xor U1616 (N_1616,N_1447,N_1482);
xor U1617 (N_1617,N_1444,N_1439);
nor U1618 (N_1618,N_1536,N_1481);
or U1619 (N_1619,N_1551,N_1524);
nand U1620 (N_1620,N_1585,N_1516);
or U1621 (N_1621,N_1412,N_1577);
nor U1622 (N_1622,N_1595,N_1527);
and U1623 (N_1623,N_1594,N_1499);
xor U1624 (N_1624,N_1555,N_1424);
and U1625 (N_1625,N_1442,N_1494);
or U1626 (N_1626,N_1474,N_1514);
nand U1627 (N_1627,N_1575,N_1558);
and U1628 (N_1628,N_1572,N_1503);
and U1629 (N_1629,N_1596,N_1475);
or U1630 (N_1630,N_1426,N_1598);
nand U1631 (N_1631,N_1550,N_1574);
or U1632 (N_1632,N_1466,N_1402);
nor U1633 (N_1633,N_1519,N_1400);
or U1634 (N_1634,N_1495,N_1542);
nand U1635 (N_1635,N_1581,N_1454);
nand U1636 (N_1636,N_1528,N_1580);
nor U1637 (N_1637,N_1425,N_1413);
nand U1638 (N_1638,N_1545,N_1420);
and U1639 (N_1639,N_1518,N_1599);
nor U1640 (N_1640,N_1531,N_1418);
nand U1641 (N_1641,N_1556,N_1446);
or U1642 (N_1642,N_1484,N_1544);
xnor U1643 (N_1643,N_1549,N_1453);
nor U1644 (N_1644,N_1489,N_1411);
nor U1645 (N_1645,N_1586,N_1526);
xnor U1646 (N_1646,N_1525,N_1560);
or U1647 (N_1647,N_1557,N_1449);
xor U1648 (N_1648,N_1520,N_1523);
and U1649 (N_1649,N_1569,N_1521);
nor U1650 (N_1650,N_1451,N_1468);
nor U1651 (N_1651,N_1592,N_1513);
nor U1652 (N_1652,N_1419,N_1496);
nor U1653 (N_1653,N_1405,N_1456);
nor U1654 (N_1654,N_1504,N_1500);
nor U1655 (N_1655,N_1488,N_1492);
or U1656 (N_1656,N_1506,N_1477);
and U1657 (N_1657,N_1460,N_1529);
nand U1658 (N_1658,N_1441,N_1473);
or U1659 (N_1659,N_1448,N_1597);
nand U1660 (N_1660,N_1458,N_1443);
xnor U1661 (N_1661,N_1465,N_1497);
xnor U1662 (N_1662,N_1507,N_1517);
xnor U1663 (N_1663,N_1583,N_1430);
or U1664 (N_1664,N_1414,N_1433);
and U1665 (N_1665,N_1547,N_1509);
and U1666 (N_1666,N_1429,N_1537);
nand U1667 (N_1667,N_1427,N_1532);
nor U1668 (N_1668,N_1486,N_1570);
and U1669 (N_1669,N_1554,N_1478);
nor U1670 (N_1670,N_1501,N_1470);
and U1671 (N_1671,N_1469,N_1487);
nor U1672 (N_1672,N_1505,N_1471);
or U1673 (N_1673,N_1541,N_1543);
xnor U1674 (N_1674,N_1573,N_1552);
xnor U1675 (N_1675,N_1476,N_1450);
xor U1676 (N_1676,N_1510,N_1565);
and U1677 (N_1677,N_1540,N_1483);
nor U1678 (N_1678,N_1582,N_1437);
or U1679 (N_1679,N_1538,N_1522);
nor U1680 (N_1680,N_1436,N_1479);
nand U1681 (N_1681,N_1408,N_1568);
or U1682 (N_1682,N_1533,N_1584);
or U1683 (N_1683,N_1415,N_1406);
nor U1684 (N_1684,N_1431,N_1409);
and U1685 (N_1685,N_1512,N_1567);
nor U1686 (N_1686,N_1511,N_1566);
or U1687 (N_1687,N_1403,N_1515);
xor U1688 (N_1688,N_1539,N_1579);
nor U1689 (N_1689,N_1563,N_1410);
and U1690 (N_1690,N_1434,N_1491);
nand U1691 (N_1691,N_1508,N_1591);
nand U1692 (N_1692,N_1461,N_1553);
nor U1693 (N_1693,N_1564,N_1587);
xnor U1694 (N_1694,N_1407,N_1463);
or U1695 (N_1695,N_1535,N_1445);
xor U1696 (N_1696,N_1548,N_1561);
and U1697 (N_1697,N_1576,N_1593);
and U1698 (N_1698,N_1472,N_1455);
nand U1699 (N_1699,N_1546,N_1467);
nor U1700 (N_1700,N_1486,N_1572);
and U1701 (N_1701,N_1501,N_1519);
nor U1702 (N_1702,N_1529,N_1421);
and U1703 (N_1703,N_1500,N_1461);
or U1704 (N_1704,N_1473,N_1427);
or U1705 (N_1705,N_1512,N_1476);
nand U1706 (N_1706,N_1574,N_1442);
nand U1707 (N_1707,N_1578,N_1477);
or U1708 (N_1708,N_1440,N_1527);
xor U1709 (N_1709,N_1545,N_1560);
xnor U1710 (N_1710,N_1535,N_1408);
nand U1711 (N_1711,N_1422,N_1583);
nor U1712 (N_1712,N_1549,N_1410);
xnor U1713 (N_1713,N_1545,N_1513);
or U1714 (N_1714,N_1429,N_1436);
and U1715 (N_1715,N_1479,N_1503);
and U1716 (N_1716,N_1486,N_1442);
or U1717 (N_1717,N_1521,N_1486);
nor U1718 (N_1718,N_1465,N_1496);
and U1719 (N_1719,N_1453,N_1540);
nand U1720 (N_1720,N_1549,N_1522);
and U1721 (N_1721,N_1523,N_1488);
xor U1722 (N_1722,N_1475,N_1454);
xor U1723 (N_1723,N_1521,N_1497);
nor U1724 (N_1724,N_1432,N_1567);
and U1725 (N_1725,N_1532,N_1516);
xnor U1726 (N_1726,N_1412,N_1440);
nor U1727 (N_1727,N_1410,N_1445);
nand U1728 (N_1728,N_1567,N_1578);
nor U1729 (N_1729,N_1504,N_1511);
xnor U1730 (N_1730,N_1515,N_1565);
nand U1731 (N_1731,N_1406,N_1565);
or U1732 (N_1732,N_1516,N_1523);
and U1733 (N_1733,N_1536,N_1524);
nor U1734 (N_1734,N_1544,N_1562);
or U1735 (N_1735,N_1400,N_1554);
nor U1736 (N_1736,N_1539,N_1440);
xor U1737 (N_1737,N_1590,N_1432);
and U1738 (N_1738,N_1541,N_1516);
nor U1739 (N_1739,N_1437,N_1526);
xnor U1740 (N_1740,N_1576,N_1555);
nand U1741 (N_1741,N_1418,N_1480);
nand U1742 (N_1742,N_1499,N_1531);
and U1743 (N_1743,N_1409,N_1403);
or U1744 (N_1744,N_1497,N_1569);
nand U1745 (N_1745,N_1533,N_1510);
or U1746 (N_1746,N_1510,N_1465);
nand U1747 (N_1747,N_1532,N_1560);
and U1748 (N_1748,N_1475,N_1459);
and U1749 (N_1749,N_1561,N_1525);
or U1750 (N_1750,N_1480,N_1498);
and U1751 (N_1751,N_1575,N_1409);
or U1752 (N_1752,N_1524,N_1479);
or U1753 (N_1753,N_1494,N_1413);
nor U1754 (N_1754,N_1490,N_1420);
nand U1755 (N_1755,N_1479,N_1568);
xnor U1756 (N_1756,N_1450,N_1559);
nand U1757 (N_1757,N_1572,N_1448);
or U1758 (N_1758,N_1455,N_1490);
xor U1759 (N_1759,N_1512,N_1446);
nand U1760 (N_1760,N_1544,N_1487);
xor U1761 (N_1761,N_1480,N_1543);
and U1762 (N_1762,N_1544,N_1475);
nand U1763 (N_1763,N_1560,N_1499);
nand U1764 (N_1764,N_1427,N_1458);
xor U1765 (N_1765,N_1508,N_1420);
and U1766 (N_1766,N_1576,N_1557);
or U1767 (N_1767,N_1480,N_1502);
nor U1768 (N_1768,N_1483,N_1573);
nand U1769 (N_1769,N_1456,N_1566);
and U1770 (N_1770,N_1580,N_1511);
nor U1771 (N_1771,N_1581,N_1490);
xor U1772 (N_1772,N_1435,N_1527);
or U1773 (N_1773,N_1593,N_1507);
nand U1774 (N_1774,N_1413,N_1520);
nand U1775 (N_1775,N_1425,N_1434);
or U1776 (N_1776,N_1575,N_1403);
nor U1777 (N_1777,N_1549,N_1446);
xor U1778 (N_1778,N_1593,N_1449);
and U1779 (N_1779,N_1533,N_1566);
nor U1780 (N_1780,N_1540,N_1414);
and U1781 (N_1781,N_1551,N_1511);
nor U1782 (N_1782,N_1452,N_1538);
or U1783 (N_1783,N_1481,N_1426);
nor U1784 (N_1784,N_1551,N_1540);
xnor U1785 (N_1785,N_1544,N_1545);
nand U1786 (N_1786,N_1415,N_1426);
and U1787 (N_1787,N_1464,N_1458);
nand U1788 (N_1788,N_1579,N_1403);
nor U1789 (N_1789,N_1595,N_1487);
nor U1790 (N_1790,N_1551,N_1444);
nor U1791 (N_1791,N_1432,N_1508);
xor U1792 (N_1792,N_1466,N_1432);
nor U1793 (N_1793,N_1521,N_1570);
nand U1794 (N_1794,N_1507,N_1488);
or U1795 (N_1795,N_1446,N_1584);
nor U1796 (N_1796,N_1521,N_1560);
or U1797 (N_1797,N_1495,N_1425);
nor U1798 (N_1798,N_1583,N_1580);
and U1799 (N_1799,N_1502,N_1509);
xnor U1800 (N_1800,N_1728,N_1675);
or U1801 (N_1801,N_1706,N_1665);
nand U1802 (N_1802,N_1685,N_1699);
xnor U1803 (N_1803,N_1740,N_1792);
nor U1804 (N_1804,N_1631,N_1686);
nor U1805 (N_1805,N_1773,N_1739);
and U1806 (N_1806,N_1653,N_1781);
nand U1807 (N_1807,N_1679,N_1669);
xnor U1808 (N_1808,N_1649,N_1700);
nor U1809 (N_1809,N_1795,N_1698);
nor U1810 (N_1810,N_1661,N_1775);
xor U1811 (N_1811,N_1790,N_1786);
nor U1812 (N_1812,N_1610,N_1757);
nand U1813 (N_1813,N_1694,N_1751);
or U1814 (N_1814,N_1683,N_1633);
xnor U1815 (N_1815,N_1616,N_1601);
xnor U1816 (N_1816,N_1655,N_1704);
and U1817 (N_1817,N_1726,N_1767);
xnor U1818 (N_1818,N_1778,N_1624);
xnor U1819 (N_1819,N_1632,N_1684);
nor U1820 (N_1820,N_1738,N_1714);
xor U1821 (N_1821,N_1777,N_1771);
and U1822 (N_1822,N_1615,N_1617);
xor U1823 (N_1823,N_1712,N_1750);
and U1824 (N_1824,N_1769,N_1672);
nand U1825 (N_1825,N_1756,N_1676);
xnor U1826 (N_1826,N_1752,N_1637);
nand U1827 (N_1827,N_1693,N_1733);
nand U1828 (N_1828,N_1677,N_1611);
or U1829 (N_1829,N_1625,N_1731);
nor U1830 (N_1830,N_1747,N_1687);
and U1831 (N_1831,N_1697,N_1722);
xor U1832 (N_1832,N_1678,N_1622);
or U1833 (N_1833,N_1695,N_1734);
xor U1834 (N_1834,N_1788,N_1784);
and U1835 (N_1835,N_1707,N_1656);
nand U1836 (N_1836,N_1755,N_1674);
xor U1837 (N_1837,N_1780,N_1647);
nor U1838 (N_1838,N_1614,N_1662);
nand U1839 (N_1839,N_1754,N_1758);
xnor U1840 (N_1840,N_1668,N_1768);
or U1841 (N_1841,N_1713,N_1719);
and U1842 (N_1842,N_1783,N_1605);
nor U1843 (N_1843,N_1664,N_1671);
or U1844 (N_1844,N_1798,N_1621);
and U1845 (N_1845,N_1644,N_1708);
nand U1846 (N_1846,N_1660,N_1727);
nand U1847 (N_1847,N_1629,N_1689);
xnor U1848 (N_1848,N_1612,N_1741);
and U1849 (N_1849,N_1774,N_1702);
xnor U1850 (N_1850,N_1630,N_1794);
nand U1851 (N_1851,N_1760,N_1763);
or U1852 (N_1852,N_1652,N_1627);
nand U1853 (N_1853,N_1729,N_1721);
xnor U1854 (N_1854,N_1765,N_1746);
or U1855 (N_1855,N_1772,N_1716);
and U1856 (N_1856,N_1658,N_1688);
or U1857 (N_1857,N_1602,N_1648);
nand U1858 (N_1858,N_1723,N_1604);
nor U1859 (N_1859,N_1645,N_1659);
or U1860 (N_1860,N_1651,N_1737);
and U1861 (N_1861,N_1646,N_1638);
nand U1862 (N_1862,N_1618,N_1789);
nor U1863 (N_1863,N_1761,N_1782);
xnor U1864 (N_1864,N_1642,N_1636);
or U1865 (N_1865,N_1690,N_1635);
nor U1866 (N_1866,N_1681,N_1692);
nor U1867 (N_1867,N_1724,N_1701);
nand U1868 (N_1868,N_1753,N_1703);
xnor U1869 (N_1869,N_1626,N_1682);
nand U1870 (N_1870,N_1613,N_1634);
nand U1871 (N_1871,N_1623,N_1725);
or U1872 (N_1872,N_1667,N_1743);
and U1873 (N_1873,N_1791,N_1715);
and U1874 (N_1874,N_1654,N_1666);
or U1875 (N_1875,N_1641,N_1709);
nand U1876 (N_1876,N_1736,N_1787);
nand U1877 (N_1877,N_1785,N_1711);
nor U1878 (N_1878,N_1673,N_1797);
nand U1879 (N_1879,N_1744,N_1691);
and U1880 (N_1880,N_1770,N_1696);
or U1881 (N_1881,N_1639,N_1650);
nor U1882 (N_1882,N_1609,N_1643);
nand U1883 (N_1883,N_1759,N_1619);
or U1884 (N_1884,N_1749,N_1764);
or U1885 (N_1885,N_1670,N_1762);
nand U1886 (N_1886,N_1705,N_1628);
nand U1887 (N_1887,N_1796,N_1608);
nor U1888 (N_1888,N_1720,N_1640);
nand U1889 (N_1889,N_1793,N_1766);
and U1890 (N_1890,N_1607,N_1730);
xnor U1891 (N_1891,N_1799,N_1779);
or U1892 (N_1892,N_1606,N_1657);
nor U1893 (N_1893,N_1735,N_1680);
nor U1894 (N_1894,N_1600,N_1603);
and U1895 (N_1895,N_1732,N_1663);
or U1896 (N_1896,N_1748,N_1718);
or U1897 (N_1897,N_1742,N_1620);
nor U1898 (N_1898,N_1710,N_1745);
nand U1899 (N_1899,N_1776,N_1717);
and U1900 (N_1900,N_1608,N_1782);
nand U1901 (N_1901,N_1709,N_1683);
xor U1902 (N_1902,N_1724,N_1728);
xnor U1903 (N_1903,N_1677,N_1744);
nand U1904 (N_1904,N_1737,N_1799);
nand U1905 (N_1905,N_1728,N_1649);
nand U1906 (N_1906,N_1739,N_1790);
or U1907 (N_1907,N_1751,N_1632);
xor U1908 (N_1908,N_1645,N_1662);
and U1909 (N_1909,N_1729,N_1642);
xnor U1910 (N_1910,N_1686,N_1715);
and U1911 (N_1911,N_1603,N_1756);
nor U1912 (N_1912,N_1642,N_1747);
and U1913 (N_1913,N_1774,N_1667);
and U1914 (N_1914,N_1740,N_1608);
xnor U1915 (N_1915,N_1700,N_1704);
nand U1916 (N_1916,N_1747,N_1618);
xor U1917 (N_1917,N_1673,N_1688);
nand U1918 (N_1918,N_1741,N_1666);
xnor U1919 (N_1919,N_1610,N_1721);
nand U1920 (N_1920,N_1710,N_1637);
nand U1921 (N_1921,N_1789,N_1683);
and U1922 (N_1922,N_1678,N_1642);
nand U1923 (N_1923,N_1729,N_1754);
xnor U1924 (N_1924,N_1634,N_1687);
nor U1925 (N_1925,N_1731,N_1779);
nand U1926 (N_1926,N_1713,N_1683);
or U1927 (N_1927,N_1639,N_1688);
and U1928 (N_1928,N_1654,N_1693);
or U1929 (N_1929,N_1671,N_1750);
nand U1930 (N_1930,N_1796,N_1708);
or U1931 (N_1931,N_1630,N_1780);
or U1932 (N_1932,N_1704,N_1770);
or U1933 (N_1933,N_1695,N_1733);
nand U1934 (N_1934,N_1695,N_1675);
nor U1935 (N_1935,N_1759,N_1699);
and U1936 (N_1936,N_1728,N_1651);
nand U1937 (N_1937,N_1629,N_1663);
nor U1938 (N_1938,N_1607,N_1606);
xnor U1939 (N_1939,N_1729,N_1604);
xnor U1940 (N_1940,N_1734,N_1781);
and U1941 (N_1941,N_1666,N_1738);
xnor U1942 (N_1942,N_1607,N_1795);
nor U1943 (N_1943,N_1632,N_1771);
or U1944 (N_1944,N_1775,N_1794);
and U1945 (N_1945,N_1759,N_1774);
xor U1946 (N_1946,N_1734,N_1706);
and U1947 (N_1947,N_1782,N_1641);
xnor U1948 (N_1948,N_1776,N_1649);
xor U1949 (N_1949,N_1772,N_1650);
nand U1950 (N_1950,N_1768,N_1720);
and U1951 (N_1951,N_1699,N_1755);
nand U1952 (N_1952,N_1780,N_1709);
nor U1953 (N_1953,N_1600,N_1632);
xor U1954 (N_1954,N_1734,N_1668);
and U1955 (N_1955,N_1745,N_1766);
xnor U1956 (N_1956,N_1713,N_1631);
nor U1957 (N_1957,N_1680,N_1606);
nor U1958 (N_1958,N_1739,N_1686);
nor U1959 (N_1959,N_1724,N_1674);
xor U1960 (N_1960,N_1652,N_1611);
and U1961 (N_1961,N_1653,N_1695);
and U1962 (N_1962,N_1682,N_1728);
and U1963 (N_1963,N_1610,N_1797);
and U1964 (N_1964,N_1624,N_1687);
nor U1965 (N_1965,N_1679,N_1677);
or U1966 (N_1966,N_1630,N_1770);
xor U1967 (N_1967,N_1649,N_1640);
and U1968 (N_1968,N_1605,N_1697);
xor U1969 (N_1969,N_1775,N_1644);
and U1970 (N_1970,N_1755,N_1789);
or U1971 (N_1971,N_1746,N_1604);
nor U1972 (N_1972,N_1663,N_1651);
nand U1973 (N_1973,N_1668,N_1790);
nor U1974 (N_1974,N_1603,N_1777);
nor U1975 (N_1975,N_1638,N_1755);
nor U1976 (N_1976,N_1626,N_1638);
nor U1977 (N_1977,N_1648,N_1699);
and U1978 (N_1978,N_1766,N_1680);
xnor U1979 (N_1979,N_1734,N_1648);
or U1980 (N_1980,N_1634,N_1736);
nand U1981 (N_1981,N_1755,N_1662);
or U1982 (N_1982,N_1667,N_1770);
or U1983 (N_1983,N_1626,N_1767);
or U1984 (N_1984,N_1719,N_1675);
or U1985 (N_1985,N_1626,N_1644);
and U1986 (N_1986,N_1607,N_1601);
nand U1987 (N_1987,N_1764,N_1630);
xor U1988 (N_1988,N_1622,N_1649);
or U1989 (N_1989,N_1673,N_1744);
and U1990 (N_1990,N_1716,N_1673);
xor U1991 (N_1991,N_1656,N_1606);
xor U1992 (N_1992,N_1633,N_1762);
or U1993 (N_1993,N_1739,N_1786);
nor U1994 (N_1994,N_1683,N_1723);
and U1995 (N_1995,N_1769,N_1620);
nand U1996 (N_1996,N_1796,N_1799);
nand U1997 (N_1997,N_1682,N_1738);
or U1998 (N_1998,N_1747,N_1795);
and U1999 (N_1999,N_1794,N_1653);
nand U2000 (N_2000,N_1812,N_1921);
nor U2001 (N_2001,N_1804,N_1874);
xor U2002 (N_2002,N_1877,N_1820);
nand U2003 (N_2003,N_1816,N_1958);
xnor U2004 (N_2004,N_1805,N_1903);
or U2005 (N_2005,N_1953,N_1980);
and U2006 (N_2006,N_1934,N_1853);
xor U2007 (N_2007,N_1902,N_1869);
xnor U2008 (N_2008,N_1864,N_1872);
or U2009 (N_2009,N_1837,N_1847);
xnor U2010 (N_2010,N_1825,N_1937);
xor U2011 (N_2011,N_1875,N_1974);
nor U2012 (N_2012,N_1815,N_1987);
xnor U2013 (N_2013,N_1912,N_1807);
nand U2014 (N_2014,N_1915,N_1893);
and U2015 (N_2015,N_1997,N_1904);
nand U2016 (N_2016,N_1830,N_1965);
nand U2017 (N_2017,N_1906,N_1859);
and U2018 (N_2018,N_1894,N_1843);
nor U2019 (N_2019,N_1907,N_1854);
and U2020 (N_2020,N_1990,N_1986);
and U2021 (N_2021,N_1892,N_1914);
xnor U2022 (N_2022,N_1909,N_1982);
nand U2023 (N_2023,N_1861,N_1802);
or U2024 (N_2024,N_1927,N_1856);
xnor U2025 (N_2025,N_1828,N_1984);
xor U2026 (N_2026,N_1800,N_1901);
or U2027 (N_2027,N_1811,N_1832);
nor U2028 (N_2028,N_1842,N_1891);
nand U2029 (N_2029,N_1942,N_1882);
or U2030 (N_2030,N_1955,N_1846);
nand U2031 (N_2031,N_1951,N_1824);
or U2032 (N_2032,N_1885,N_1940);
or U2033 (N_2033,N_1826,N_1822);
xnor U2034 (N_2034,N_1976,N_1917);
and U2035 (N_2035,N_1808,N_1971);
nand U2036 (N_2036,N_1966,N_1989);
nand U2037 (N_2037,N_1857,N_1868);
or U2038 (N_2038,N_1881,N_1941);
xnor U2039 (N_2039,N_1886,N_1890);
nor U2040 (N_2040,N_1994,N_1862);
nor U2041 (N_2041,N_1968,N_1823);
and U2042 (N_2042,N_1961,N_1801);
and U2043 (N_2043,N_1817,N_1948);
or U2044 (N_2044,N_1988,N_1880);
nor U2045 (N_2045,N_1876,N_1991);
or U2046 (N_2046,N_1999,N_1919);
nor U2047 (N_2047,N_1946,N_1970);
nor U2048 (N_2048,N_1871,N_1863);
and U2049 (N_2049,N_1979,N_1878);
nor U2050 (N_2050,N_1900,N_1806);
or U2051 (N_2051,N_1962,N_1803);
xnor U2052 (N_2052,N_1889,N_1916);
and U2053 (N_2053,N_1848,N_1924);
nand U2054 (N_2054,N_1810,N_1908);
or U2055 (N_2055,N_1897,N_1985);
and U2056 (N_2056,N_1969,N_1867);
nor U2057 (N_2057,N_1935,N_1844);
or U2058 (N_2058,N_1967,N_1992);
or U2059 (N_2059,N_1933,N_1852);
nor U2060 (N_2060,N_1841,N_1838);
nor U2061 (N_2061,N_1855,N_1814);
and U2062 (N_2062,N_1920,N_1833);
and U2063 (N_2063,N_1998,N_1944);
nand U2064 (N_2064,N_1911,N_1932);
and U2065 (N_2065,N_1926,N_1959);
nor U2066 (N_2066,N_1952,N_1887);
nor U2067 (N_2067,N_1930,N_1983);
xor U2068 (N_2068,N_1960,N_1831);
or U2069 (N_2069,N_1829,N_1918);
nand U2070 (N_2070,N_1954,N_1827);
and U2071 (N_2071,N_1809,N_1905);
and U2072 (N_2072,N_1821,N_1884);
and U2073 (N_2073,N_1973,N_1981);
xor U2074 (N_2074,N_1923,N_1977);
and U2075 (N_2075,N_1896,N_1949);
and U2076 (N_2076,N_1925,N_1978);
nor U2077 (N_2077,N_1836,N_1964);
or U2078 (N_2078,N_1950,N_1834);
and U2079 (N_2079,N_1819,N_1860);
and U2080 (N_2080,N_1895,N_1913);
and U2081 (N_2081,N_1888,N_1845);
nand U2082 (N_2082,N_1850,N_1883);
nand U2083 (N_2083,N_1839,N_1972);
nor U2084 (N_2084,N_1870,N_1835);
and U2085 (N_2085,N_1865,N_1975);
nor U2086 (N_2086,N_1943,N_1858);
nor U2087 (N_2087,N_1993,N_1849);
xnor U2088 (N_2088,N_1818,N_1840);
xnor U2089 (N_2089,N_1873,N_1813);
or U2090 (N_2090,N_1957,N_1928);
or U2091 (N_2091,N_1910,N_1938);
nand U2092 (N_2092,N_1963,N_1936);
xor U2093 (N_2093,N_1851,N_1866);
or U2094 (N_2094,N_1995,N_1899);
and U2095 (N_2095,N_1931,N_1945);
nor U2096 (N_2096,N_1929,N_1996);
or U2097 (N_2097,N_1939,N_1879);
nor U2098 (N_2098,N_1956,N_1898);
or U2099 (N_2099,N_1922,N_1947);
and U2100 (N_2100,N_1829,N_1972);
and U2101 (N_2101,N_1866,N_1856);
nor U2102 (N_2102,N_1978,N_1801);
or U2103 (N_2103,N_1995,N_1802);
nor U2104 (N_2104,N_1980,N_1990);
xnor U2105 (N_2105,N_1914,N_1986);
and U2106 (N_2106,N_1999,N_1980);
or U2107 (N_2107,N_1906,N_1974);
xor U2108 (N_2108,N_1896,N_1907);
nor U2109 (N_2109,N_1838,N_1985);
or U2110 (N_2110,N_1996,N_1839);
xnor U2111 (N_2111,N_1835,N_1996);
and U2112 (N_2112,N_1964,N_1901);
nand U2113 (N_2113,N_1879,N_1824);
nor U2114 (N_2114,N_1979,N_1993);
nor U2115 (N_2115,N_1807,N_1901);
nand U2116 (N_2116,N_1964,N_1872);
nor U2117 (N_2117,N_1812,N_1936);
nand U2118 (N_2118,N_1896,N_1862);
or U2119 (N_2119,N_1862,N_1979);
and U2120 (N_2120,N_1910,N_1986);
and U2121 (N_2121,N_1975,N_1896);
nor U2122 (N_2122,N_1991,N_1823);
and U2123 (N_2123,N_1898,N_1933);
xnor U2124 (N_2124,N_1916,N_1803);
and U2125 (N_2125,N_1895,N_1831);
nor U2126 (N_2126,N_1980,N_1913);
nand U2127 (N_2127,N_1819,N_1980);
nor U2128 (N_2128,N_1956,N_1925);
nand U2129 (N_2129,N_1992,N_1870);
xor U2130 (N_2130,N_1844,N_1817);
and U2131 (N_2131,N_1835,N_1911);
and U2132 (N_2132,N_1916,N_1923);
xor U2133 (N_2133,N_1961,N_1941);
or U2134 (N_2134,N_1968,N_1882);
xnor U2135 (N_2135,N_1865,N_1987);
nand U2136 (N_2136,N_1955,N_1850);
or U2137 (N_2137,N_1904,N_1870);
nor U2138 (N_2138,N_1819,N_1932);
and U2139 (N_2139,N_1948,N_1912);
and U2140 (N_2140,N_1967,N_1827);
and U2141 (N_2141,N_1889,N_1883);
xor U2142 (N_2142,N_1892,N_1897);
nand U2143 (N_2143,N_1879,N_1915);
or U2144 (N_2144,N_1949,N_1921);
and U2145 (N_2145,N_1969,N_1967);
or U2146 (N_2146,N_1855,N_1897);
or U2147 (N_2147,N_1948,N_1921);
or U2148 (N_2148,N_1802,N_1887);
xnor U2149 (N_2149,N_1979,N_1884);
and U2150 (N_2150,N_1901,N_1937);
and U2151 (N_2151,N_1953,N_1909);
and U2152 (N_2152,N_1991,N_1866);
or U2153 (N_2153,N_1910,N_1896);
and U2154 (N_2154,N_1992,N_1842);
and U2155 (N_2155,N_1987,N_1940);
xnor U2156 (N_2156,N_1860,N_1801);
and U2157 (N_2157,N_1920,N_1883);
xor U2158 (N_2158,N_1839,N_1948);
xor U2159 (N_2159,N_1963,N_1867);
and U2160 (N_2160,N_1916,N_1896);
nor U2161 (N_2161,N_1808,N_1809);
nand U2162 (N_2162,N_1906,N_1864);
and U2163 (N_2163,N_1904,N_1896);
xor U2164 (N_2164,N_1998,N_1952);
nand U2165 (N_2165,N_1927,N_1953);
nor U2166 (N_2166,N_1927,N_1957);
nor U2167 (N_2167,N_1907,N_1960);
xor U2168 (N_2168,N_1833,N_1918);
or U2169 (N_2169,N_1995,N_1887);
xor U2170 (N_2170,N_1908,N_1889);
xor U2171 (N_2171,N_1877,N_1808);
nor U2172 (N_2172,N_1987,N_1989);
xnor U2173 (N_2173,N_1849,N_1923);
or U2174 (N_2174,N_1844,N_1983);
nand U2175 (N_2175,N_1805,N_1924);
nor U2176 (N_2176,N_1840,N_1983);
and U2177 (N_2177,N_1924,N_1974);
nor U2178 (N_2178,N_1865,N_1940);
nor U2179 (N_2179,N_1876,N_1961);
nor U2180 (N_2180,N_1864,N_1973);
nor U2181 (N_2181,N_1801,N_1852);
and U2182 (N_2182,N_1857,N_1811);
or U2183 (N_2183,N_1964,N_1994);
nor U2184 (N_2184,N_1889,N_1988);
xor U2185 (N_2185,N_1989,N_1975);
xnor U2186 (N_2186,N_1977,N_1903);
and U2187 (N_2187,N_1818,N_1864);
nor U2188 (N_2188,N_1981,N_1952);
or U2189 (N_2189,N_1830,N_1819);
nor U2190 (N_2190,N_1979,N_1956);
nand U2191 (N_2191,N_1890,N_1821);
or U2192 (N_2192,N_1898,N_1808);
and U2193 (N_2193,N_1826,N_1851);
and U2194 (N_2194,N_1875,N_1907);
or U2195 (N_2195,N_1891,N_1963);
nor U2196 (N_2196,N_1896,N_1997);
xor U2197 (N_2197,N_1899,N_1857);
nor U2198 (N_2198,N_1805,N_1951);
nand U2199 (N_2199,N_1964,N_1866);
nand U2200 (N_2200,N_2008,N_2136);
nand U2201 (N_2201,N_2106,N_2031);
nand U2202 (N_2202,N_2184,N_2076);
and U2203 (N_2203,N_2120,N_2004);
nor U2204 (N_2204,N_2045,N_2104);
or U2205 (N_2205,N_2020,N_2190);
xnor U2206 (N_2206,N_2152,N_2072);
nand U2207 (N_2207,N_2089,N_2035);
nand U2208 (N_2208,N_2118,N_2049);
xor U2209 (N_2209,N_2005,N_2092);
and U2210 (N_2210,N_2030,N_2175);
or U2211 (N_2211,N_2069,N_2119);
nand U2212 (N_2212,N_2047,N_2054);
or U2213 (N_2213,N_2042,N_2068);
and U2214 (N_2214,N_2151,N_2178);
nand U2215 (N_2215,N_2058,N_2032);
xnor U2216 (N_2216,N_2080,N_2150);
nor U2217 (N_2217,N_2098,N_2082);
nor U2218 (N_2218,N_2041,N_2037);
xor U2219 (N_2219,N_2064,N_2091);
nor U2220 (N_2220,N_2148,N_2133);
xnor U2221 (N_2221,N_2117,N_2022);
nor U2222 (N_2222,N_2075,N_2142);
nor U2223 (N_2223,N_2157,N_2000);
xnor U2224 (N_2224,N_2036,N_2100);
nand U2225 (N_2225,N_2132,N_2193);
nand U2226 (N_2226,N_2006,N_2027);
and U2227 (N_2227,N_2138,N_2172);
nand U2228 (N_2228,N_2182,N_2090);
nand U2229 (N_2229,N_2025,N_2083);
xnor U2230 (N_2230,N_2085,N_2097);
nand U2231 (N_2231,N_2026,N_2048);
nand U2232 (N_2232,N_2056,N_2194);
or U2233 (N_2233,N_2188,N_2122);
or U2234 (N_2234,N_2050,N_2198);
nand U2235 (N_2235,N_2125,N_2162);
or U2236 (N_2236,N_2010,N_2185);
or U2237 (N_2237,N_2060,N_2168);
xnor U2238 (N_2238,N_2009,N_2003);
and U2239 (N_2239,N_2167,N_2199);
and U2240 (N_2240,N_2023,N_2124);
xnor U2241 (N_2241,N_2158,N_2145);
or U2242 (N_2242,N_2176,N_2109);
xnor U2243 (N_2243,N_2177,N_2121);
and U2244 (N_2244,N_2012,N_2017);
or U2245 (N_2245,N_2134,N_2115);
nor U2246 (N_2246,N_2135,N_2123);
nand U2247 (N_2247,N_2081,N_2110);
nor U2248 (N_2248,N_2112,N_2161);
and U2249 (N_2249,N_2144,N_2087);
nor U2250 (N_2250,N_2019,N_2007);
nand U2251 (N_2251,N_2011,N_2166);
xnor U2252 (N_2252,N_2163,N_2086);
nand U2253 (N_2253,N_2102,N_2192);
and U2254 (N_2254,N_2015,N_2094);
xnor U2255 (N_2255,N_2062,N_2108);
xor U2256 (N_2256,N_2088,N_2130);
xor U2257 (N_2257,N_2016,N_2074);
nor U2258 (N_2258,N_2065,N_2055);
nor U2259 (N_2259,N_2093,N_2186);
or U2260 (N_2260,N_2155,N_2171);
nand U2261 (N_2261,N_2127,N_2195);
nor U2262 (N_2262,N_2160,N_2140);
nand U2263 (N_2263,N_2164,N_2073);
nor U2264 (N_2264,N_2105,N_2066);
and U2265 (N_2265,N_2107,N_2034);
nand U2266 (N_2266,N_2154,N_2173);
and U2267 (N_2267,N_2028,N_2053);
xnor U2268 (N_2268,N_2165,N_2040);
nand U2269 (N_2269,N_2116,N_2179);
nand U2270 (N_2270,N_2078,N_2099);
or U2271 (N_2271,N_2128,N_2039);
xor U2272 (N_2272,N_2191,N_2197);
nand U2273 (N_2273,N_2143,N_2029);
and U2274 (N_2274,N_2111,N_2113);
and U2275 (N_2275,N_2033,N_2187);
and U2276 (N_2276,N_2084,N_2057);
nand U2277 (N_2277,N_2024,N_2170);
nor U2278 (N_2278,N_2014,N_2181);
and U2279 (N_2279,N_2096,N_2070);
or U2280 (N_2280,N_2061,N_2103);
or U2281 (N_2281,N_2131,N_2051);
xnor U2282 (N_2282,N_2038,N_2169);
xnor U2283 (N_2283,N_2101,N_2044);
xor U2284 (N_2284,N_2059,N_2183);
and U2285 (N_2285,N_2002,N_2052);
nor U2286 (N_2286,N_2139,N_2137);
nand U2287 (N_2287,N_2071,N_2095);
xnor U2288 (N_2288,N_2180,N_2149);
and U2289 (N_2289,N_2189,N_2147);
and U2290 (N_2290,N_2079,N_2153);
or U2291 (N_2291,N_2156,N_2018);
xor U2292 (N_2292,N_2077,N_2159);
nor U2293 (N_2293,N_2046,N_2001);
nor U2294 (N_2294,N_2063,N_2174);
or U2295 (N_2295,N_2141,N_2126);
and U2296 (N_2296,N_2196,N_2013);
nor U2297 (N_2297,N_2021,N_2067);
and U2298 (N_2298,N_2043,N_2146);
nand U2299 (N_2299,N_2129,N_2114);
nor U2300 (N_2300,N_2036,N_2191);
and U2301 (N_2301,N_2113,N_2008);
and U2302 (N_2302,N_2163,N_2159);
nor U2303 (N_2303,N_2081,N_2129);
nand U2304 (N_2304,N_2136,N_2041);
xor U2305 (N_2305,N_2090,N_2116);
or U2306 (N_2306,N_2071,N_2184);
or U2307 (N_2307,N_2005,N_2011);
xnor U2308 (N_2308,N_2186,N_2119);
or U2309 (N_2309,N_2139,N_2197);
xnor U2310 (N_2310,N_2027,N_2077);
and U2311 (N_2311,N_2032,N_2013);
nor U2312 (N_2312,N_2029,N_2107);
and U2313 (N_2313,N_2182,N_2062);
nand U2314 (N_2314,N_2172,N_2055);
xor U2315 (N_2315,N_2047,N_2020);
nand U2316 (N_2316,N_2134,N_2060);
nor U2317 (N_2317,N_2044,N_2193);
nor U2318 (N_2318,N_2005,N_2181);
nand U2319 (N_2319,N_2173,N_2078);
nand U2320 (N_2320,N_2128,N_2129);
and U2321 (N_2321,N_2194,N_2143);
nor U2322 (N_2322,N_2095,N_2134);
nor U2323 (N_2323,N_2127,N_2108);
and U2324 (N_2324,N_2152,N_2145);
and U2325 (N_2325,N_2024,N_2061);
or U2326 (N_2326,N_2060,N_2146);
and U2327 (N_2327,N_2179,N_2110);
and U2328 (N_2328,N_2030,N_2157);
or U2329 (N_2329,N_2032,N_2022);
nor U2330 (N_2330,N_2183,N_2100);
nand U2331 (N_2331,N_2045,N_2152);
and U2332 (N_2332,N_2180,N_2147);
nand U2333 (N_2333,N_2109,N_2033);
or U2334 (N_2334,N_2103,N_2072);
nor U2335 (N_2335,N_2121,N_2087);
and U2336 (N_2336,N_2118,N_2061);
nor U2337 (N_2337,N_2188,N_2108);
nand U2338 (N_2338,N_2000,N_2181);
nand U2339 (N_2339,N_2110,N_2015);
nand U2340 (N_2340,N_2150,N_2002);
nor U2341 (N_2341,N_2134,N_2047);
nor U2342 (N_2342,N_2192,N_2104);
and U2343 (N_2343,N_2085,N_2040);
xnor U2344 (N_2344,N_2142,N_2117);
and U2345 (N_2345,N_2074,N_2100);
and U2346 (N_2346,N_2183,N_2036);
or U2347 (N_2347,N_2111,N_2178);
or U2348 (N_2348,N_2070,N_2012);
nand U2349 (N_2349,N_2009,N_2093);
and U2350 (N_2350,N_2008,N_2143);
nand U2351 (N_2351,N_2157,N_2086);
xor U2352 (N_2352,N_2014,N_2162);
or U2353 (N_2353,N_2030,N_2071);
xor U2354 (N_2354,N_2055,N_2103);
xnor U2355 (N_2355,N_2104,N_2179);
nand U2356 (N_2356,N_2096,N_2149);
xnor U2357 (N_2357,N_2043,N_2029);
and U2358 (N_2358,N_2123,N_2005);
or U2359 (N_2359,N_2114,N_2192);
nand U2360 (N_2360,N_2196,N_2009);
xor U2361 (N_2361,N_2100,N_2079);
nand U2362 (N_2362,N_2042,N_2164);
nand U2363 (N_2363,N_2178,N_2101);
nand U2364 (N_2364,N_2061,N_2071);
xor U2365 (N_2365,N_2191,N_2074);
nor U2366 (N_2366,N_2155,N_2069);
nand U2367 (N_2367,N_2121,N_2095);
nor U2368 (N_2368,N_2095,N_2109);
or U2369 (N_2369,N_2174,N_2109);
xnor U2370 (N_2370,N_2051,N_2138);
nand U2371 (N_2371,N_2178,N_2046);
or U2372 (N_2372,N_2084,N_2028);
and U2373 (N_2373,N_2143,N_2160);
or U2374 (N_2374,N_2196,N_2194);
or U2375 (N_2375,N_2040,N_2145);
xnor U2376 (N_2376,N_2030,N_2007);
nand U2377 (N_2377,N_2095,N_2011);
and U2378 (N_2378,N_2102,N_2112);
and U2379 (N_2379,N_2197,N_2104);
nor U2380 (N_2380,N_2066,N_2085);
xor U2381 (N_2381,N_2059,N_2069);
or U2382 (N_2382,N_2187,N_2119);
nor U2383 (N_2383,N_2030,N_2134);
nand U2384 (N_2384,N_2029,N_2180);
nor U2385 (N_2385,N_2148,N_2084);
xor U2386 (N_2386,N_2016,N_2160);
or U2387 (N_2387,N_2011,N_2001);
xnor U2388 (N_2388,N_2159,N_2064);
and U2389 (N_2389,N_2036,N_2174);
or U2390 (N_2390,N_2037,N_2103);
or U2391 (N_2391,N_2124,N_2010);
or U2392 (N_2392,N_2082,N_2051);
xnor U2393 (N_2393,N_2187,N_2159);
xor U2394 (N_2394,N_2110,N_2104);
xor U2395 (N_2395,N_2141,N_2023);
nor U2396 (N_2396,N_2135,N_2179);
and U2397 (N_2397,N_2031,N_2036);
nand U2398 (N_2398,N_2021,N_2080);
or U2399 (N_2399,N_2081,N_2097);
nor U2400 (N_2400,N_2364,N_2297);
or U2401 (N_2401,N_2271,N_2348);
or U2402 (N_2402,N_2340,N_2388);
xnor U2403 (N_2403,N_2344,N_2272);
or U2404 (N_2404,N_2200,N_2229);
nand U2405 (N_2405,N_2209,N_2208);
nand U2406 (N_2406,N_2284,N_2238);
xnor U2407 (N_2407,N_2249,N_2281);
xnor U2408 (N_2408,N_2204,N_2294);
xnor U2409 (N_2409,N_2338,N_2296);
nand U2410 (N_2410,N_2369,N_2223);
or U2411 (N_2411,N_2222,N_2334);
nand U2412 (N_2412,N_2362,N_2360);
or U2413 (N_2413,N_2361,N_2372);
nand U2414 (N_2414,N_2311,N_2299);
and U2415 (N_2415,N_2290,N_2381);
and U2416 (N_2416,N_2310,N_2258);
nand U2417 (N_2417,N_2260,N_2307);
nor U2418 (N_2418,N_2350,N_2315);
nand U2419 (N_2419,N_2206,N_2345);
or U2420 (N_2420,N_2225,N_2250);
xnor U2421 (N_2421,N_2373,N_2291);
nor U2422 (N_2422,N_2252,N_2327);
nand U2423 (N_2423,N_2283,N_2339);
and U2424 (N_2424,N_2328,N_2368);
xnor U2425 (N_2425,N_2216,N_2247);
and U2426 (N_2426,N_2226,N_2389);
nand U2427 (N_2427,N_2386,N_2363);
nor U2428 (N_2428,N_2275,N_2265);
or U2429 (N_2429,N_2262,N_2282);
and U2430 (N_2430,N_2205,N_2367);
xor U2431 (N_2431,N_2397,N_2277);
or U2432 (N_2432,N_2385,N_2399);
xor U2433 (N_2433,N_2246,N_2212);
and U2434 (N_2434,N_2341,N_2313);
and U2435 (N_2435,N_2248,N_2379);
nor U2436 (N_2436,N_2269,N_2286);
nor U2437 (N_2437,N_2211,N_2289);
nor U2438 (N_2438,N_2220,N_2357);
or U2439 (N_2439,N_2314,N_2263);
xor U2440 (N_2440,N_2215,N_2312);
nor U2441 (N_2441,N_2243,N_2221);
nand U2442 (N_2442,N_2330,N_2261);
xor U2443 (N_2443,N_2202,N_2394);
nor U2444 (N_2444,N_2255,N_2395);
nand U2445 (N_2445,N_2317,N_2266);
nor U2446 (N_2446,N_2321,N_2240);
and U2447 (N_2447,N_2234,N_2231);
nand U2448 (N_2448,N_2251,N_2320);
xor U2449 (N_2449,N_2359,N_2292);
nor U2450 (N_2450,N_2207,N_2319);
nor U2451 (N_2451,N_2336,N_2318);
or U2452 (N_2452,N_2356,N_2393);
nand U2453 (N_2453,N_2335,N_2259);
xor U2454 (N_2454,N_2264,N_2214);
xnor U2455 (N_2455,N_2387,N_2285);
xor U2456 (N_2456,N_2365,N_2309);
nor U2457 (N_2457,N_2337,N_2383);
nand U2458 (N_2458,N_2242,N_2280);
xnor U2459 (N_2459,N_2376,N_2322);
and U2460 (N_2460,N_2398,N_2352);
or U2461 (N_2461,N_2342,N_2274);
and U2462 (N_2462,N_2366,N_2382);
and U2463 (N_2463,N_2270,N_2232);
or U2464 (N_2464,N_2236,N_2257);
nand U2465 (N_2465,N_2324,N_2323);
nor U2466 (N_2466,N_2213,N_2377);
and U2467 (N_2467,N_2235,N_2233);
nor U2468 (N_2468,N_2391,N_2329);
and U2469 (N_2469,N_2332,N_2287);
or U2470 (N_2470,N_2227,N_2210);
and U2471 (N_2471,N_2370,N_2353);
and U2472 (N_2472,N_2304,N_2241);
nand U2473 (N_2473,N_2267,N_2331);
and U2474 (N_2474,N_2349,N_2203);
or U2475 (N_2475,N_2295,N_2347);
nand U2476 (N_2476,N_2201,N_2219);
and U2477 (N_2477,N_2228,N_2253);
nor U2478 (N_2478,N_2326,N_2279);
and U2479 (N_2479,N_2380,N_2374);
nor U2480 (N_2480,N_2298,N_2217);
or U2481 (N_2481,N_2333,N_2378);
nor U2482 (N_2482,N_2276,N_2375);
nor U2483 (N_2483,N_2300,N_2355);
nor U2484 (N_2484,N_2351,N_2371);
or U2485 (N_2485,N_2316,N_2256);
nand U2486 (N_2486,N_2230,N_2244);
or U2487 (N_2487,N_2346,N_2325);
or U2488 (N_2488,N_2305,N_2390);
nor U2489 (N_2489,N_2306,N_2384);
or U2490 (N_2490,N_2354,N_2245);
nand U2491 (N_2491,N_2288,N_2239);
nand U2492 (N_2492,N_2396,N_2293);
or U2493 (N_2493,N_2392,N_2303);
nand U2494 (N_2494,N_2301,N_2358);
nor U2495 (N_2495,N_2237,N_2268);
and U2496 (N_2496,N_2343,N_2224);
xor U2497 (N_2497,N_2302,N_2218);
xnor U2498 (N_2498,N_2278,N_2273);
nand U2499 (N_2499,N_2254,N_2308);
and U2500 (N_2500,N_2309,N_2202);
xor U2501 (N_2501,N_2364,N_2311);
nand U2502 (N_2502,N_2280,N_2258);
nor U2503 (N_2503,N_2200,N_2335);
nand U2504 (N_2504,N_2322,N_2243);
nor U2505 (N_2505,N_2259,N_2339);
and U2506 (N_2506,N_2297,N_2352);
xnor U2507 (N_2507,N_2392,N_2296);
nor U2508 (N_2508,N_2233,N_2256);
nand U2509 (N_2509,N_2278,N_2396);
and U2510 (N_2510,N_2386,N_2268);
nor U2511 (N_2511,N_2215,N_2362);
nor U2512 (N_2512,N_2210,N_2259);
nand U2513 (N_2513,N_2341,N_2265);
nand U2514 (N_2514,N_2303,N_2259);
xnor U2515 (N_2515,N_2382,N_2375);
nor U2516 (N_2516,N_2265,N_2365);
or U2517 (N_2517,N_2384,N_2213);
nor U2518 (N_2518,N_2319,N_2237);
nand U2519 (N_2519,N_2353,N_2240);
nor U2520 (N_2520,N_2359,N_2398);
or U2521 (N_2521,N_2291,N_2271);
and U2522 (N_2522,N_2217,N_2380);
nand U2523 (N_2523,N_2383,N_2280);
xor U2524 (N_2524,N_2261,N_2288);
and U2525 (N_2525,N_2277,N_2393);
xnor U2526 (N_2526,N_2316,N_2385);
xor U2527 (N_2527,N_2251,N_2399);
nand U2528 (N_2528,N_2311,N_2341);
nor U2529 (N_2529,N_2262,N_2237);
or U2530 (N_2530,N_2310,N_2343);
or U2531 (N_2531,N_2280,N_2376);
xnor U2532 (N_2532,N_2231,N_2287);
or U2533 (N_2533,N_2280,N_2221);
xnor U2534 (N_2534,N_2370,N_2341);
or U2535 (N_2535,N_2298,N_2339);
nand U2536 (N_2536,N_2393,N_2279);
and U2537 (N_2537,N_2232,N_2281);
nand U2538 (N_2538,N_2359,N_2217);
or U2539 (N_2539,N_2305,N_2295);
or U2540 (N_2540,N_2250,N_2224);
and U2541 (N_2541,N_2295,N_2372);
xor U2542 (N_2542,N_2313,N_2275);
and U2543 (N_2543,N_2220,N_2257);
nor U2544 (N_2544,N_2291,N_2233);
and U2545 (N_2545,N_2302,N_2382);
or U2546 (N_2546,N_2242,N_2299);
xor U2547 (N_2547,N_2326,N_2309);
nand U2548 (N_2548,N_2201,N_2251);
nor U2549 (N_2549,N_2300,N_2304);
and U2550 (N_2550,N_2256,N_2276);
xnor U2551 (N_2551,N_2286,N_2372);
nor U2552 (N_2552,N_2229,N_2272);
xor U2553 (N_2553,N_2339,N_2317);
or U2554 (N_2554,N_2319,N_2379);
nand U2555 (N_2555,N_2359,N_2206);
and U2556 (N_2556,N_2311,N_2317);
xor U2557 (N_2557,N_2369,N_2296);
or U2558 (N_2558,N_2212,N_2292);
nand U2559 (N_2559,N_2330,N_2371);
nor U2560 (N_2560,N_2240,N_2306);
and U2561 (N_2561,N_2224,N_2399);
and U2562 (N_2562,N_2299,N_2216);
nand U2563 (N_2563,N_2333,N_2328);
xnor U2564 (N_2564,N_2345,N_2252);
and U2565 (N_2565,N_2399,N_2339);
nor U2566 (N_2566,N_2224,N_2240);
xor U2567 (N_2567,N_2367,N_2308);
xor U2568 (N_2568,N_2276,N_2235);
and U2569 (N_2569,N_2375,N_2270);
or U2570 (N_2570,N_2247,N_2388);
nor U2571 (N_2571,N_2322,N_2340);
nand U2572 (N_2572,N_2215,N_2224);
and U2573 (N_2573,N_2291,N_2376);
nor U2574 (N_2574,N_2205,N_2308);
or U2575 (N_2575,N_2333,N_2316);
nand U2576 (N_2576,N_2214,N_2276);
nor U2577 (N_2577,N_2385,N_2294);
and U2578 (N_2578,N_2264,N_2369);
or U2579 (N_2579,N_2206,N_2220);
or U2580 (N_2580,N_2386,N_2374);
and U2581 (N_2581,N_2319,N_2249);
nand U2582 (N_2582,N_2316,N_2238);
or U2583 (N_2583,N_2398,N_2204);
nand U2584 (N_2584,N_2331,N_2366);
or U2585 (N_2585,N_2327,N_2232);
xnor U2586 (N_2586,N_2372,N_2377);
xor U2587 (N_2587,N_2375,N_2376);
nor U2588 (N_2588,N_2270,N_2311);
xnor U2589 (N_2589,N_2313,N_2286);
xor U2590 (N_2590,N_2254,N_2284);
xor U2591 (N_2591,N_2206,N_2270);
or U2592 (N_2592,N_2352,N_2388);
or U2593 (N_2593,N_2288,N_2355);
nor U2594 (N_2594,N_2311,N_2380);
nand U2595 (N_2595,N_2342,N_2388);
nand U2596 (N_2596,N_2304,N_2213);
xnor U2597 (N_2597,N_2253,N_2386);
and U2598 (N_2598,N_2338,N_2216);
xor U2599 (N_2599,N_2272,N_2376);
nor U2600 (N_2600,N_2545,N_2580);
nand U2601 (N_2601,N_2501,N_2564);
and U2602 (N_2602,N_2586,N_2410);
xor U2603 (N_2603,N_2595,N_2464);
nand U2604 (N_2604,N_2570,N_2444);
nand U2605 (N_2605,N_2423,N_2588);
nor U2606 (N_2606,N_2450,N_2548);
xnor U2607 (N_2607,N_2518,N_2406);
xor U2608 (N_2608,N_2524,N_2554);
nand U2609 (N_2609,N_2521,N_2476);
or U2610 (N_2610,N_2456,N_2500);
and U2611 (N_2611,N_2445,N_2573);
nand U2612 (N_2612,N_2407,N_2474);
and U2613 (N_2613,N_2590,N_2492);
nor U2614 (N_2614,N_2561,N_2491);
or U2615 (N_2615,N_2468,N_2473);
or U2616 (N_2616,N_2553,N_2490);
or U2617 (N_2617,N_2538,N_2598);
and U2618 (N_2618,N_2438,N_2514);
nand U2619 (N_2619,N_2462,N_2408);
nand U2620 (N_2620,N_2513,N_2503);
nor U2621 (N_2621,N_2466,N_2530);
and U2622 (N_2622,N_2584,N_2569);
nand U2623 (N_2623,N_2502,N_2405);
or U2624 (N_2624,N_2437,N_2576);
nand U2625 (N_2625,N_2589,N_2458);
nand U2626 (N_2626,N_2452,N_2451);
or U2627 (N_2627,N_2435,N_2540);
nor U2628 (N_2628,N_2532,N_2574);
xnor U2629 (N_2629,N_2411,N_2505);
or U2630 (N_2630,N_2594,N_2494);
nand U2631 (N_2631,N_2471,N_2443);
nor U2632 (N_2632,N_2403,N_2568);
nor U2633 (N_2633,N_2432,N_2495);
nor U2634 (N_2634,N_2425,N_2519);
xnor U2635 (N_2635,N_2424,N_2557);
or U2636 (N_2636,N_2575,N_2563);
nor U2637 (N_2637,N_2401,N_2577);
xnor U2638 (N_2638,N_2592,N_2489);
or U2639 (N_2639,N_2537,N_2566);
nor U2640 (N_2640,N_2463,N_2559);
and U2641 (N_2641,N_2525,N_2591);
nor U2642 (N_2642,N_2529,N_2552);
xor U2643 (N_2643,N_2597,N_2414);
nand U2644 (N_2644,N_2541,N_2431);
xnor U2645 (N_2645,N_2497,N_2507);
nand U2646 (N_2646,N_2496,N_2539);
nand U2647 (N_2647,N_2436,N_2565);
or U2648 (N_2648,N_2479,N_2511);
or U2649 (N_2649,N_2512,N_2404);
nand U2650 (N_2650,N_2421,N_2587);
xor U2651 (N_2651,N_2543,N_2417);
nand U2652 (N_2652,N_2482,N_2413);
nor U2653 (N_2653,N_2446,N_2430);
nor U2654 (N_2654,N_2434,N_2422);
or U2655 (N_2655,N_2428,N_2523);
xor U2656 (N_2656,N_2533,N_2493);
xor U2657 (N_2657,N_2429,N_2478);
nand U2658 (N_2658,N_2571,N_2506);
xnor U2659 (N_2659,N_2516,N_2499);
or U2660 (N_2660,N_2442,N_2467);
nand U2661 (N_2661,N_2420,N_2483);
xnor U2662 (N_2662,N_2572,N_2400);
or U2663 (N_2663,N_2440,N_2549);
or U2664 (N_2664,N_2498,N_2427);
nor U2665 (N_2665,N_2487,N_2527);
nand U2666 (N_2666,N_2415,N_2453);
and U2667 (N_2667,N_2412,N_2480);
nor U2668 (N_2668,N_2455,N_2509);
nand U2669 (N_2669,N_2581,N_2560);
nand U2670 (N_2670,N_2508,N_2599);
nand U2671 (N_2671,N_2486,N_2583);
xor U2672 (N_2672,N_2472,N_2504);
nor U2673 (N_2673,N_2550,N_2515);
and U2674 (N_2674,N_2593,N_2531);
xor U2675 (N_2675,N_2555,N_2542);
or U2676 (N_2676,N_2426,N_2433);
nor U2677 (N_2677,N_2461,N_2488);
nor U2678 (N_2678,N_2578,N_2510);
nand U2679 (N_2679,N_2562,N_2454);
nand U2680 (N_2680,N_2481,N_2579);
and U2681 (N_2681,N_2536,N_2544);
nor U2682 (N_2682,N_2522,N_2517);
xor U2683 (N_2683,N_2416,N_2465);
and U2684 (N_2684,N_2459,N_2556);
or U2685 (N_2685,N_2441,N_2485);
nand U2686 (N_2686,N_2567,N_2546);
nand U2687 (N_2687,N_2551,N_2520);
or U2688 (N_2688,N_2535,N_2460);
xnor U2689 (N_2689,N_2419,N_2558);
nor U2690 (N_2690,N_2477,N_2439);
xnor U2691 (N_2691,N_2409,N_2475);
and U2692 (N_2692,N_2534,N_2596);
and U2693 (N_2693,N_2547,N_2484);
or U2694 (N_2694,N_2418,N_2449);
nor U2695 (N_2695,N_2470,N_2448);
nand U2696 (N_2696,N_2457,N_2585);
and U2697 (N_2697,N_2402,N_2526);
and U2698 (N_2698,N_2469,N_2447);
nor U2699 (N_2699,N_2528,N_2582);
nand U2700 (N_2700,N_2486,N_2520);
nor U2701 (N_2701,N_2472,N_2579);
nor U2702 (N_2702,N_2479,N_2537);
xor U2703 (N_2703,N_2531,N_2515);
xnor U2704 (N_2704,N_2481,N_2441);
nor U2705 (N_2705,N_2464,N_2545);
and U2706 (N_2706,N_2490,N_2565);
and U2707 (N_2707,N_2552,N_2523);
xnor U2708 (N_2708,N_2445,N_2556);
nand U2709 (N_2709,N_2553,N_2586);
or U2710 (N_2710,N_2439,N_2531);
xnor U2711 (N_2711,N_2590,N_2508);
nand U2712 (N_2712,N_2541,N_2433);
or U2713 (N_2713,N_2403,N_2422);
or U2714 (N_2714,N_2519,N_2447);
nand U2715 (N_2715,N_2445,N_2468);
nor U2716 (N_2716,N_2435,N_2413);
and U2717 (N_2717,N_2542,N_2490);
xnor U2718 (N_2718,N_2544,N_2409);
nor U2719 (N_2719,N_2453,N_2525);
and U2720 (N_2720,N_2557,N_2590);
or U2721 (N_2721,N_2477,N_2562);
nor U2722 (N_2722,N_2401,N_2465);
and U2723 (N_2723,N_2465,N_2484);
nand U2724 (N_2724,N_2454,N_2435);
nor U2725 (N_2725,N_2574,N_2499);
nand U2726 (N_2726,N_2558,N_2466);
or U2727 (N_2727,N_2569,N_2542);
nand U2728 (N_2728,N_2572,N_2589);
nor U2729 (N_2729,N_2593,N_2407);
and U2730 (N_2730,N_2573,N_2509);
xnor U2731 (N_2731,N_2515,N_2539);
or U2732 (N_2732,N_2441,N_2555);
nor U2733 (N_2733,N_2483,N_2456);
nand U2734 (N_2734,N_2505,N_2593);
nand U2735 (N_2735,N_2480,N_2415);
and U2736 (N_2736,N_2486,N_2403);
xor U2737 (N_2737,N_2428,N_2444);
nand U2738 (N_2738,N_2483,N_2589);
and U2739 (N_2739,N_2451,N_2533);
and U2740 (N_2740,N_2555,N_2588);
and U2741 (N_2741,N_2501,N_2563);
nand U2742 (N_2742,N_2568,N_2510);
nor U2743 (N_2743,N_2539,N_2406);
and U2744 (N_2744,N_2464,N_2463);
and U2745 (N_2745,N_2465,N_2413);
or U2746 (N_2746,N_2570,N_2541);
xnor U2747 (N_2747,N_2560,N_2567);
nand U2748 (N_2748,N_2570,N_2558);
nand U2749 (N_2749,N_2594,N_2517);
nand U2750 (N_2750,N_2534,N_2429);
and U2751 (N_2751,N_2502,N_2445);
nand U2752 (N_2752,N_2534,N_2450);
nand U2753 (N_2753,N_2578,N_2531);
xnor U2754 (N_2754,N_2589,N_2509);
and U2755 (N_2755,N_2441,N_2572);
and U2756 (N_2756,N_2496,N_2492);
nor U2757 (N_2757,N_2416,N_2453);
xor U2758 (N_2758,N_2400,N_2547);
xor U2759 (N_2759,N_2494,N_2489);
nand U2760 (N_2760,N_2564,N_2565);
or U2761 (N_2761,N_2498,N_2597);
nand U2762 (N_2762,N_2594,N_2412);
nand U2763 (N_2763,N_2595,N_2546);
nand U2764 (N_2764,N_2583,N_2525);
or U2765 (N_2765,N_2572,N_2489);
nand U2766 (N_2766,N_2574,N_2520);
nor U2767 (N_2767,N_2537,N_2529);
nand U2768 (N_2768,N_2562,N_2447);
or U2769 (N_2769,N_2402,N_2482);
xnor U2770 (N_2770,N_2473,N_2493);
xor U2771 (N_2771,N_2595,N_2461);
nand U2772 (N_2772,N_2536,N_2522);
nor U2773 (N_2773,N_2456,N_2479);
nor U2774 (N_2774,N_2524,N_2535);
xnor U2775 (N_2775,N_2553,N_2545);
nor U2776 (N_2776,N_2488,N_2457);
nand U2777 (N_2777,N_2440,N_2465);
nand U2778 (N_2778,N_2403,N_2593);
or U2779 (N_2779,N_2434,N_2549);
and U2780 (N_2780,N_2558,N_2463);
or U2781 (N_2781,N_2422,N_2594);
nand U2782 (N_2782,N_2515,N_2424);
xor U2783 (N_2783,N_2514,N_2587);
or U2784 (N_2784,N_2476,N_2504);
and U2785 (N_2785,N_2550,N_2417);
xor U2786 (N_2786,N_2415,N_2587);
nand U2787 (N_2787,N_2522,N_2559);
or U2788 (N_2788,N_2570,N_2552);
nor U2789 (N_2789,N_2509,N_2567);
and U2790 (N_2790,N_2579,N_2463);
xnor U2791 (N_2791,N_2445,N_2402);
nand U2792 (N_2792,N_2562,N_2544);
xnor U2793 (N_2793,N_2426,N_2530);
nor U2794 (N_2794,N_2486,N_2413);
and U2795 (N_2795,N_2432,N_2501);
nor U2796 (N_2796,N_2582,N_2587);
or U2797 (N_2797,N_2500,N_2477);
xnor U2798 (N_2798,N_2547,N_2577);
nor U2799 (N_2799,N_2499,N_2423);
xnor U2800 (N_2800,N_2634,N_2601);
or U2801 (N_2801,N_2746,N_2777);
or U2802 (N_2802,N_2685,N_2769);
or U2803 (N_2803,N_2793,N_2714);
xor U2804 (N_2804,N_2704,N_2703);
nor U2805 (N_2805,N_2759,N_2682);
nand U2806 (N_2806,N_2605,N_2661);
xnor U2807 (N_2807,N_2699,N_2786);
or U2808 (N_2808,N_2772,N_2632);
nand U2809 (N_2809,N_2734,N_2787);
nand U2810 (N_2810,N_2628,N_2762);
nand U2811 (N_2811,N_2798,N_2768);
nand U2812 (N_2812,N_2783,N_2775);
or U2813 (N_2813,N_2707,N_2780);
nand U2814 (N_2814,N_2736,N_2720);
nand U2815 (N_2815,N_2669,N_2748);
nor U2816 (N_2816,N_2667,N_2701);
xor U2817 (N_2817,N_2664,N_2738);
or U2818 (N_2818,N_2675,N_2718);
and U2819 (N_2819,N_2790,N_2722);
or U2820 (N_2820,N_2670,N_2795);
xnor U2821 (N_2821,N_2668,N_2785);
nor U2822 (N_2822,N_2677,N_2717);
xnor U2823 (N_2823,N_2604,N_2732);
and U2824 (N_2824,N_2660,N_2648);
nand U2825 (N_2825,N_2650,N_2633);
or U2826 (N_2826,N_2615,N_2743);
or U2827 (N_2827,N_2635,N_2681);
nor U2828 (N_2828,N_2606,N_2709);
or U2829 (N_2829,N_2740,N_2691);
xor U2830 (N_2830,N_2629,N_2751);
nor U2831 (N_2831,N_2617,N_2774);
nand U2832 (N_2832,N_2758,N_2706);
and U2833 (N_2833,N_2612,N_2645);
and U2834 (N_2834,N_2610,N_2602);
nand U2835 (N_2835,N_2711,N_2725);
xnor U2836 (N_2836,N_2792,N_2698);
nor U2837 (N_2837,N_2656,N_2659);
or U2838 (N_2838,N_2726,N_2640);
nor U2839 (N_2839,N_2654,N_2733);
nand U2840 (N_2840,N_2766,N_2652);
and U2841 (N_2841,N_2694,N_2773);
xnor U2842 (N_2842,N_2686,N_2760);
nand U2843 (N_2843,N_2653,N_2765);
nor U2844 (N_2844,N_2679,N_2692);
nand U2845 (N_2845,N_2778,N_2754);
xor U2846 (N_2846,N_2716,N_2728);
and U2847 (N_2847,N_2781,N_2735);
xnor U2848 (N_2848,N_2770,N_2729);
nand U2849 (N_2849,N_2764,N_2776);
nor U2850 (N_2850,N_2646,N_2797);
nand U2851 (N_2851,N_2647,N_2688);
and U2852 (N_2852,N_2627,N_2641);
xor U2853 (N_2853,N_2672,N_2655);
xor U2854 (N_2854,N_2782,N_2731);
or U2855 (N_2855,N_2637,N_2621);
and U2856 (N_2856,N_2705,N_2613);
nor U2857 (N_2857,N_2695,N_2618);
nand U2858 (N_2858,N_2752,N_2708);
nor U2859 (N_2859,N_2649,N_2763);
and U2860 (N_2860,N_2724,N_2771);
or U2861 (N_2861,N_2642,N_2620);
nor U2862 (N_2862,N_2662,N_2689);
xnor U2863 (N_2863,N_2710,N_2609);
nand U2864 (N_2864,N_2611,N_2638);
and U2865 (N_2865,N_2631,N_2639);
nand U2866 (N_2866,N_2624,N_2794);
nand U2867 (N_2867,N_2799,N_2791);
nand U2868 (N_2868,N_2600,N_2619);
nand U2869 (N_2869,N_2678,N_2749);
or U2870 (N_2870,N_2614,N_2750);
nor U2871 (N_2871,N_2756,N_2788);
or U2872 (N_2872,N_2723,N_2630);
and U2873 (N_2873,N_2683,N_2713);
nand U2874 (N_2874,N_2666,N_2753);
xor U2875 (N_2875,N_2745,N_2644);
nor U2876 (N_2876,N_2684,N_2657);
xnor U2877 (N_2877,N_2623,N_2789);
nand U2878 (N_2878,N_2767,N_2779);
or U2879 (N_2879,N_2625,N_2700);
nand U2880 (N_2880,N_2676,N_2796);
or U2881 (N_2881,N_2730,N_2643);
nor U2882 (N_2882,N_2693,N_2680);
xnor U2883 (N_2883,N_2607,N_2626);
or U2884 (N_2884,N_2697,N_2742);
xnor U2885 (N_2885,N_2622,N_2715);
xor U2886 (N_2886,N_2658,N_2721);
or U2887 (N_2887,N_2757,N_2690);
and U2888 (N_2888,N_2741,N_2674);
or U2889 (N_2889,N_2737,N_2739);
nor U2890 (N_2890,N_2687,N_2636);
and U2891 (N_2891,N_2671,N_2651);
nor U2892 (N_2892,N_2727,N_2784);
nand U2893 (N_2893,N_2702,N_2744);
nor U2894 (N_2894,N_2747,N_2663);
and U2895 (N_2895,N_2608,N_2665);
and U2896 (N_2896,N_2696,N_2761);
nor U2897 (N_2897,N_2755,N_2603);
xnor U2898 (N_2898,N_2719,N_2616);
xnor U2899 (N_2899,N_2673,N_2712);
nor U2900 (N_2900,N_2745,N_2610);
nor U2901 (N_2901,N_2687,N_2624);
and U2902 (N_2902,N_2672,N_2661);
nor U2903 (N_2903,N_2717,N_2662);
nand U2904 (N_2904,N_2779,N_2612);
and U2905 (N_2905,N_2612,N_2725);
xnor U2906 (N_2906,N_2621,N_2726);
and U2907 (N_2907,N_2794,N_2661);
or U2908 (N_2908,N_2759,N_2663);
or U2909 (N_2909,N_2780,N_2708);
or U2910 (N_2910,N_2716,N_2718);
xor U2911 (N_2911,N_2708,N_2797);
and U2912 (N_2912,N_2798,N_2651);
and U2913 (N_2913,N_2784,N_2653);
and U2914 (N_2914,N_2608,N_2667);
or U2915 (N_2915,N_2633,N_2636);
nor U2916 (N_2916,N_2788,N_2777);
nor U2917 (N_2917,N_2700,N_2763);
and U2918 (N_2918,N_2691,N_2779);
xor U2919 (N_2919,N_2763,N_2648);
nand U2920 (N_2920,N_2693,N_2687);
nor U2921 (N_2921,N_2754,N_2794);
and U2922 (N_2922,N_2686,N_2721);
and U2923 (N_2923,N_2706,N_2697);
and U2924 (N_2924,N_2774,N_2764);
nand U2925 (N_2925,N_2760,N_2626);
nor U2926 (N_2926,N_2631,N_2772);
xor U2927 (N_2927,N_2747,N_2649);
nand U2928 (N_2928,N_2622,N_2664);
nor U2929 (N_2929,N_2684,N_2645);
nand U2930 (N_2930,N_2696,N_2746);
nand U2931 (N_2931,N_2664,N_2784);
and U2932 (N_2932,N_2607,N_2771);
nand U2933 (N_2933,N_2680,N_2688);
nand U2934 (N_2934,N_2620,N_2788);
or U2935 (N_2935,N_2744,N_2633);
nor U2936 (N_2936,N_2758,N_2742);
or U2937 (N_2937,N_2622,N_2767);
nor U2938 (N_2938,N_2606,N_2639);
nor U2939 (N_2939,N_2644,N_2787);
xor U2940 (N_2940,N_2669,N_2783);
or U2941 (N_2941,N_2659,N_2746);
nand U2942 (N_2942,N_2691,N_2643);
xor U2943 (N_2943,N_2702,N_2763);
nor U2944 (N_2944,N_2741,N_2736);
xor U2945 (N_2945,N_2720,N_2716);
nor U2946 (N_2946,N_2624,N_2709);
xor U2947 (N_2947,N_2616,N_2777);
and U2948 (N_2948,N_2773,N_2697);
or U2949 (N_2949,N_2652,N_2606);
xnor U2950 (N_2950,N_2692,N_2722);
xor U2951 (N_2951,N_2671,N_2760);
and U2952 (N_2952,N_2607,N_2710);
and U2953 (N_2953,N_2690,N_2675);
nor U2954 (N_2954,N_2676,N_2740);
nor U2955 (N_2955,N_2633,N_2620);
or U2956 (N_2956,N_2769,N_2602);
and U2957 (N_2957,N_2697,N_2654);
and U2958 (N_2958,N_2641,N_2600);
or U2959 (N_2959,N_2773,N_2757);
and U2960 (N_2960,N_2645,N_2767);
nand U2961 (N_2961,N_2769,N_2686);
xnor U2962 (N_2962,N_2759,N_2644);
and U2963 (N_2963,N_2621,N_2764);
xor U2964 (N_2964,N_2627,N_2673);
and U2965 (N_2965,N_2775,N_2704);
xor U2966 (N_2966,N_2605,N_2686);
and U2967 (N_2967,N_2627,N_2728);
nand U2968 (N_2968,N_2618,N_2629);
nand U2969 (N_2969,N_2751,N_2645);
xnor U2970 (N_2970,N_2699,N_2723);
nor U2971 (N_2971,N_2603,N_2662);
nor U2972 (N_2972,N_2760,N_2742);
xnor U2973 (N_2973,N_2658,N_2622);
xor U2974 (N_2974,N_2702,N_2651);
nor U2975 (N_2975,N_2696,N_2648);
xnor U2976 (N_2976,N_2706,N_2787);
nor U2977 (N_2977,N_2770,N_2731);
or U2978 (N_2978,N_2676,N_2674);
or U2979 (N_2979,N_2715,N_2667);
or U2980 (N_2980,N_2722,N_2783);
or U2981 (N_2981,N_2771,N_2601);
nand U2982 (N_2982,N_2698,N_2651);
or U2983 (N_2983,N_2746,N_2640);
and U2984 (N_2984,N_2744,N_2773);
and U2985 (N_2985,N_2785,N_2789);
nor U2986 (N_2986,N_2756,N_2703);
xnor U2987 (N_2987,N_2722,N_2799);
nor U2988 (N_2988,N_2615,N_2750);
and U2989 (N_2989,N_2636,N_2753);
nand U2990 (N_2990,N_2717,N_2678);
xnor U2991 (N_2991,N_2621,N_2755);
nor U2992 (N_2992,N_2749,N_2658);
nor U2993 (N_2993,N_2772,N_2724);
nand U2994 (N_2994,N_2714,N_2605);
and U2995 (N_2995,N_2752,N_2719);
xnor U2996 (N_2996,N_2603,N_2702);
or U2997 (N_2997,N_2795,N_2698);
xnor U2998 (N_2998,N_2717,N_2720);
or U2999 (N_2999,N_2736,N_2781);
xor UO_0 (O_0,N_2853,N_2960);
nand UO_1 (O_1,N_2871,N_2887);
nor UO_2 (O_2,N_2847,N_2836);
and UO_3 (O_3,N_2903,N_2838);
xor UO_4 (O_4,N_2910,N_2965);
nor UO_5 (O_5,N_2999,N_2899);
or UO_6 (O_6,N_2976,N_2907);
xnor UO_7 (O_7,N_2921,N_2914);
nand UO_8 (O_8,N_2818,N_2821);
or UO_9 (O_9,N_2876,N_2879);
nor UO_10 (O_10,N_2854,N_2890);
xnor UO_11 (O_11,N_2852,N_2917);
nor UO_12 (O_12,N_2866,N_2974);
xnor UO_13 (O_13,N_2932,N_2802);
and UO_14 (O_14,N_2982,N_2943);
or UO_15 (O_15,N_2955,N_2858);
xnor UO_16 (O_16,N_2830,N_2967);
nand UO_17 (O_17,N_2951,N_2908);
xnor UO_18 (O_18,N_2988,N_2979);
nor UO_19 (O_19,N_2807,N_2933);
or UO_20 (O_20,N_2940,N_2916);
nor UO_21 (O_21,N_2948,N_2983);
nand UO_22 (O_22,N_2884,N_2813);
or UO_23 (O_23,N_2808,N_2920);
and UO_24 (O_24,N_2843,N_2995);
nor UO_25 (O_25,N_2826,N_2975);
nor UO_26 (O_26,N_2942,N_2824);
xor UO_27 (O_27,N_2962,N_2895);
and UO_28 (O_28,N_2964,N_2936);
xnor UO_29 (O_29,N_2927,N_2883);
nand UO_30 (O_30,N_2810,N_2823);
and UO_31 (O_31,N_2819,N_2874);
or UO_32 (O_32,N_2850,N_2928);
xnor UO_33 (O_33,N_2905,N_2862);
or UO_34 (O_34,N_2877,N_2956);
nor UO_35 (O_35,N_2954,N_2941);
xnor UO_36 (O_36,N_2896,N_2841);
nor UO_37 (O_37,N_2885,N_2978);
or UO_38 (O_38,N_2844,N_2860);
and UO_39 (O_39,N_2882,N_2811);
nand UO_40 (O_40,N_2959,N_2912);
and UO_41 (O_41,N_2863,N_2909);
nor UO_42 (O_42,N_2919,N_2868);
and UO_43 (O_43,N_2981,N_2925);
or UO_44 (O_44,N_2831,N_2889);
xnor UO_45 (O_45,N_2873,N_2969);
nand UO_46 (O_46,N_2881,N_2953);
nand UO_47 (O_47,N_2865,N_2970);
nor UO_48 (O_48,N_2817,N_2875);
and UO_49 (O_49,N_2977,N_2918);
nand UO_50 (O_50,N_2856,N_2849);
xnor UO_51 (O_51,N_2901,N_2915);
nand UO_52 (O_52,N_2855,N_2958);
or UO_53 (O_53,N_2944,N_2991);
nand UO_54 (O_54,N_2878,N_2822);
nand UO_55 (O_55,N_2832,N_2846);
xnor UO_56 (O_56,N_2906,N_2900);
or UO_57 (O_57,N_2867,N_2806);
nor UO_58 (O_58,N_2893,N_2957);
nor UO_59 (O_59,N_2801,N_2851);
xor UO_60 (O_60,N_2987,N_2968);
or UO_61 (O_61,N_2859,N_2992);
nor UO_62 (O_62,N_2897,N_2805);
xnor UO_63 (O_63,N_2952,N_2946);
or UO_64 (O_64,N_2848,N_2994);
nand UO_65 (O_65,N_2803,N_2949);
nor UO_66 (O_66,N_2922,N_2997);
xnor UO_67 (O_67,N_2835,N_2809);
or UO_68 (O_68,N_2926,N_2986);
and UO_69 (O_69,N_2985,N_2869);
or UO_70 (O_70,N_2947,N_2834);
and UO_71 (O_71,N_2872,N_2935);
xnor UO_72 (O_72,N_2870,N_2989);
xnor UO_73 (O_73,N_2924,N_2894);
nor UO_74 (O_74,N_2934,N_2804);
and UO_75 (O_75,N_2996,N_2923);
xnor UO_76 (O_76,N_2845,N_2891);
xnor UO_77 (O_77,N_2837,N_2800);
xnor UO_78 (O_78,N_2828,N_2842);
or UO_79 (O_79,N_2950,N_2839);
or UO_80 (O_80,N_2880,N_2945);
xor UO_81 (O_81,N_2857,N_2888);
xor UO_82 (O_82,N_2902,N_2904);
or UO_83 (O_83,N_2833,N_2911);
xor UO_84 (O_84,N_2825,N_2966);
or UO_85 (O_85,N_2814,N_2892);
and UO_86 (O_86,N_2993,N_2930);
and UO_87 (O_87,N_2972,N_2939);
nor UO_88 (O_88,N_2980,N_2963);
or UO_89 (O_89,N_2829,N_2840);
and UO_90 (O_90,N_2998,N_2938);
and UO_91 (O_91,N_2815,N_2961);
and UO_92 (O_92,N_2990,N_2816);
xor UO_93 (O_93,N_2864,N_2861);
or UO_94 (O_94,N_2913,N_2973);
nand UO_95 (O_95,N_2812,N_2937);
and UO_96 (O_96,N_2827,N_2984);
or UO_97 (O_97,N_2820,N_2886);
nand UO_98 (O_98,N_2929,N_2971);
xnor UO_99 (O_99,N_2898,N_2931);
nand UO_100 (O_100,N_2847,N_2817);
or UO_101 (O_101,N_2968,N_2893);
xor UO_102 (O_102,N_2986,N_2848);
or UO_103 (O_103,N_2865,N_2851);
or UO_104 (O_104,N_2923,N_2890);
xnor UO_105 (O_105,N_2928,N_2963);
nor UO_106 (O_106,N_2837,N_2934);
nor UO_107 (O_107,N_2949,N_2823);
nor UO_108 (O_108,N_2884,N_2950);
or UO_109 (O_109,N_2903,N_2890);
nand UO_110 (O_110,N_2843,N_2850);
nand UO_111 (O_111,N_2858,N_2910);
nor UO_112 (O_112,N_2891,N_2896);
xnor UO_113 (O_113,N_2879,N_2919);
nor UO_114 (O_114,N_2823,N_2811);
or UO_115 (O_115,N_2829,N_2996);
xnor UO_116 (O_116,N_2988,N_2981);
nand UO_117 (O_117,N_2870,N_2953);
xor UO_118 (O_118,N_2934,N_2902);
nand UO_119 (O_119,N_2944,N_2927);
or UO_120 (O_120,N_2820,N_2973);
xor UO_121 (O_121,N_2960,N_2812);
or UO_122 (O_122,N_2864,N_2994);
and UO_123 (O_123,N_2927,N_2810);
nand UO_124 (O_124,N_2848,N_2893);
or UO_125 (O_125,N_2936,N_2860);
and UO_126 (O_126,N_2862,N_2824);
and UO_127 (O_127,N_2807,N_2900);
xor UO_128 (O_128,N_2933,N_2804);
or UO_129 (O_129,N_2948,N_2807);
or UO_130 (O_130,N_2819,N_2824);
or UO_131 (O_131,N_2917,N_2831);
nor UO_132 (O_132,N_2909,N_2845);
or UO_133 (O_133,N_2982,N_2961);
nand UO_134 (O_134,N_2959,N_2881);
nand UO_135 (O_135,N_2871,N_2862);
or UO_136 (O_136,N_2890,N_2906);
nor UO_137 (O_137,N_2904,N_2942);
and UO_138 (O_138,N_2852,N_2869);
nor UO_139 (O_139,N_2821,N_2867);
and UO_140 (O_140,N_2867,N_2970);
xnor UO_141 (O_141,N_2848,N_2922);
and UO_142 (O_142,N_2869,N_2902);
nand UO_143 (O_143,N_2821,N_2847);
or UO_144 (O_144,N_2988,N_2879);
xnor UO_145 (O_145,N_2873,N_2858);
nor UO_146 (O_146,N_2831,N_2962);
or UO_147 (O_147,N_2920,N_2951);
or UO_148 (O_148,N_2956,N_2922);
nand UO_149 (O_149,N_2956,N_2995);
xnor UO_150 (O_150,N_2888,N_2910);
and UO_151 (O_151,N_2957,N_2903);
nand UO_152 (O_152,N_2984,N_2920);
xnor UO_153 (O_153,N_2936,N_2993);
nand UO_154 (O_154,N_2834,N_2987);
xor UO_155 (O_155,N_2961,N_2994);
xnor UO_156 (O_156,N_2912,N_2816);
and UO_157 (O_157,N_2852,N_2826);
nand UO_158 (O_158,N_2822,N_2913);
nand UO_159 (O_159,N_2907,N_2886);
nor UO_160 (O_160,N_2873,N_2944);
or UO_161 (O_161,N_2959,N_2904);
xor UO_162 (O_162,N_2949,N_2937);
nand UO_163 (O_163,N_2932,N_2954);
xor UO_164 (O_164,N_2982,N_2817);
or UO_165 (O_165,N_2865,N_2859);
xnor UO_166 (O_166,N_2835,N_2962);
nand UO_167 (O_167,N_2920,N_2831);
xnor UO_168 (O_168,N_2912,N_2967);
nor UO_169 (O_169,N_2922,N_2969);
nor UO_170 (O_170,N_2935,N_2888);
nor UO_171 (O_171,N_2951,N_2837);
nor UO_172 (O_172,N_2900,N_2951);
nand UO_173 (O_173,N_2972,N_2951);
nor UO_174 (O_174,N_2805,N_2880);
xnor UO_175 (O_175,N_2857,N_2853);
nand UO_176 (O_176,N_2882,N_2969);
nor UO_177 (O_177,N_2894,N_2812);
xnor UO_178 (O_178,N_2946,N_2923);
or UO_179 (O_179,N_2823,N_2988);
and UO_180 (O_180,N_2850,N_2942);
or UO_181 (O_181,N_2819,N_2825);
xnor UO_182 (O_182,N_2896,N_2813);
or UO_183 (O_183,N_2872,N_2885);
nor UO_184 (O_184,N_2856,N_2886);
nor UO_185 (O_185,N_2847,N_2972);
nand UO_186 (O_186,N_2923,N_2917);
and UO_187 (O_187,N_2854,N_2974);
and UO_188 (O_188,N_2940,N_2802);
nand UO_189 (O_189,N_2840,N_2983);
nand UO_190 (O_190,N_2979,N_2885);
or UO_191 (O_191,N_2948,N_2886);
and UO_192 (O_192,N_2845,N_2988);
nand UO_193 (O_193,N_2835,N_2934);
nand UO_194 (O_194,N_2957,N_2933);
nand UO_195 (O_195,N_2814,N_2943);
nor UO_196 (O_196,N_2867,N_2822);
nor UO_197 (O_197,N_2808,N_2992);
nand UO_198 (O_198,N_2942,N_2988);
or UO_199 (O_199,N_2800,N_2921);
xnor UO_200 (O_200,N_2934,N_2912);
nand UO_201 (O_201,N_2907,N_2913);
nand UO_202 (O_202,N_2933,N_2827);
and UO_203 (O_203,N_2922,N_2952);
nor UO_204 (O_204,N_2944,N_2986);
and UO_205 (O_205,N_2847,N_2855);
xor UO_206 (O_206,N_2871,N_2964);
or UO_207 (O_207,N_2863,N_2826);
nand UO_208 (O_208,N_2873,N_2882);
and UO_209 (O_209,N_2850,N_2893);
nor UO_210 (O_210,N_2925,N_2951);
nand UO_211 (O_211,N_2918,N_2965);
nor UO_212 (O_212,N_2870,N_2925);
nand UO_213 (O_213,N_2953,N_2801);
and UO_214 (O_214,N_2818,N_2959);
or UO_215 (O_215,N_2931,N_2877);
nand UO_216 (O_216,N_2860,N_2887);
nor UO_217 (O_217,N_2839,N_2818);
xnor UO_218 (O_218,N_2852,N_2916);
nand UO_219 (O_219,N_2950,N_2920);
nand UO_220 (O_220,N_2859,N_2872);
nor UO_221 (O_221,N_2853,N_2802);
nor UO_222 (O_222,N_2945,N_2802);
xor UO_223 (O_223,N_2936,N_2904);
xnor UO_224 (O_224,N_2839,N_2880);
nand UO_225 (O_225,N_2823,N_2990);
nor UO_226 (O_226,N_2944,N_2865);
nand UO_227 (O_227,N_2995,N_2955);
nand UO_228 (O_228,N_2803,N_2965);
and UO_229 (O_229,N_2826,N_2878);
nor UO_230 (O_230,N_2983,N_2817);
xor UO_231 (O_231,N_2942,N_2830);
nand UO_232 (O_232,N_2897,N_2943);
or UO_233 (O_233,N_2953,N_2950);
nor UO_234 (O_234,N_2846,N_2974);
and UO_235 (O_235,N_2943,N_2993);
nor UO_236 (O_236,N_2932,N_2988);
nor UO_237 (O_237,N_2813,N_2886);
nand UO_238 (O_238,N_2902,N_2896);
and UO_239 (O_239,N_2894,N_2914);
nor UO_240 (O_240,N_2997,N_2832);
xor UO_241 (O_241,N_2942,N_2938);
xor UO_242 (O_242,N_2871,N_2943);
or UO_243 (O_243,N_2956,N_2854);
nor UO_244 (O_244,N_2969,N_2915);
xor UO_245 (O_245,N_2801,N_2962);
or UO_246 (O_246,N_2886,N_2878);
and UO_247 (O_247,N_2951,N_2856);
or UO_248 (O_248,N_2941,N_2911);
and UO_249 (O_249,N_2908,N_2914);
or UO_250 (O_250,N_2875,N_2874);
nor UO_251 (O_251,N_2861,N_2887);
and UO_252 (O_252,N_2995,N_2902);
and UO_253 (O_253,N_2836,N_2963);
xnor UO_254 (O_254,N_2948,N_2926);
nand UO_255 (O_255,N_2937,N_2950);
xor UO_256 (O_256,N_2879,N_2901);
nand UO_257 (O_257,N_2969,N_2948);
nand UO_258 (O_258,N_2925,N_2819);
or UO_259 (O_259,N_2856,N_2869);
and UO_260 (O_260,N_2814,N_2927);
nand UO_261 (O_261,N_2800,N_2934);
and UO_262 (O_262,N_2948,N_2868);
or UO_263 (O_263,N_2879,N_2836);
nor UO_264 (O_264,N_2852,N_2876);
xnor UO_265 (O_265,N_2862,N_2806);
or UO_266 (O_266,N_2892,N_2897);
or UO_267 (O_267,N_2830,N_2987);
and UO_268 (O_268,N_2916,N_2959);
or UO_269 (O_269,N_2823,N_2820);
xnor UO_270 (O_270,N_2869,N_2880);
and UO_271 (O_271,N_2843,N_2865);
nand UO_272 (O_272,N_2916,N_2946);
xor UO_273 (O_273,N_2871,N_2878);
nand UO_274 (O_274,N_2886,N_2824);
nand UO_275 (O_275,N_2811,N_2854);
and UO_276 (O_276,N_2819,N_2850);
and UO_277 (O_277,N_2999,N_2927);
nand UO_278 (O_278,N_2956,N_2812);
nand UO_279 (O_279,N_2829,N_2827);
xnor UO_280 (O_280,N_2966,N_2857);
xnor UO_281 (O_281,N_2950,N_2992);
xor UO_282 (O_282,N_2954,N_2863);
and UO_283 (O_283,N_2951,N_2826);
nand UO_284 (O_284,N_2866,N_2822);
xor UO_285 (O_285,N_2941,N_2900);
nand UO_286 (O_286,N_2844,N_2841);
xnor UO_287 (O_287,N_2909,N_2908);
and UO_288 (O_288,N_2869,N_2981);
xnor UO_289 (O_289,N_2848,N_2999);
nand UO_290 (O_290,N_2940,N_2988);
xnor UO_291 (O_291,N_2937,N_2894);
and UO_292 (O_292,N_2847,N_2908);
nor UO_293 (O_293,N_2812,N_2983);
and UO_294 (O_294,N_2975,N_2917);
nor UO_295 (O_295,N_2956,N_2903);
and UO_296 (O_296,N_2805,N_2993);
xor UO_297 (O_297,N_2891,N_2910);
and UO_298 (O_298,N_2943,N_2979);
nor UO_299 (O_299,N_2847,N_2985);
or UO_300 (O_300,N_2960,N_2991);
nand UO_301 (O_301,N_2873,N_2897);
and UO_302 (O_302,N_2902,N_2918);
xor UO_303 (O_303,N_2918,N_2883);
xnor UO_304 (O_304,N_2845,N_2837);
nand UO_305 (O_305,N_2933,N_2992);
nor UO_306 (O_306,N_2992,N_2892);
nand UO_307 (O_307,N_2959,N_2822);
xor UO_308 (O_308,N_2885,N_2841);
or UO_309 (O_309,N_2917,N_2899);
nand UO_310 (O_310,N_2916,N_2925);
or UO_311 (O_311,N_2875,N_2911);
and UO_312 (O_312,N_2823,N_2874);
xor UO_313 (O_313,N_2950,N_2893);
and UO_314 (O_314,N_2967,N_2813);
nor UO_315 (O_315,N_2903,N_2873);
nand UO_316 (O_316,N_2994,N_2957);
nand UO_317 (O_317,N_2877,N_2902);
xor UO_318 (O_318,N_2927,N_2916);
nand UO_319 (O_319,N_2808,N_2809);
nand UO_320 (O_320,N_2845,N_2821);
nor UO_321 (O_321,N_2832,N_2940);
or UO_322 (O_322,N_2869,N_2835);
nor UO_323 (O_323,N_2909,N_2970);
nor UO_324 (O_324,N_2834,N_2870);
nor UO_325 (O_325,N_2957,N_2825);
xor UO_326 (O_326,N_2813,N_2970);
or UO_327 (O_327,N_2964,N_2915);
or UO_328 (O_328,N_2887,N_2936);
and UO_329 (O_329,N_2932,N_2929);
nand UO_330 (O_330,N_2969,N_2810);
and UO_331 (O_331,N_2889,N_2877);
xor UO_332 (O_332,N_2968,N_2910);
and UO_333 (O_333,N_2851,N_2848);
xnor UO_334 (O_334,N_2926,N_2978);
and UO_335 (O_335,N_2877,N_2871);
nand UO_336 (O_336,N_2828,N_2952);
or UO_337 (O_337,N_2909,N_2981);
or UO_338 (O_338,N_2968,N_2941);
or UO_339 (O_339,N_2846,N_2884);
or UO_340 (O_340,N_2885,N_2984);
xor UO_341 (O_341,N_2901,N_2826);
and UO_342 (O_342,N_2889,N_2875);
and UO_343 (O_343,N_2997,N_2927);
nand UO_344 (O_344,N_2855,N_2920);
nand UO_345 (O_345,N_2814,N_2853);
nor UO_346 (O_346,N_2994,N_2914);
xnor UO_347 (O_347,N_2827,N_2972);
and UO_348 (O_348,N_2966,N_2800);
or UO_349 (O_349,N_2872,N_2933);
or UO_350 (O_350,N_2885,N_2983);
or UO_351 (O_351,N_2903,N_2885);
xor UO_352 (O_352,N_2987,N_2965);
or UO_353 (O_353,N_2872,N_2882);
nand UO_354 (O_354,N_2925,N_2977);
xnor UO_355 (O_355,N_2879,N_2953);
nand UO_356 (O_356,N_2847,N_2916);
xnor UO_357 (O_357,N_2959,N_2919);
and UO_358 (O_358,N_2922,N_2827);
nand UO_359 (O_359,N_2937,N_2891);
nand UO_360 (O_360,N_2924,N_2932);
and UO_361 (O_361,N_2820,N_2801);
and UO_362 (O_362,N_2889,N_2859);
and UO_363 (O_363,N_2998,N_2916);
and UO_364 (O_364,N_2982,N_2911);
nor UO_365 (O_365,N_2979,N_2831);
and UO_366 (O_366,N_2876,N_2973);
nor UO_367 (O_367,N_2805,N_2823);
nand UO_368 (O_368,N_2812,N_2837);
nor UO_369 (O_369,N_2863,N_2823);
nor UO_370 (O_370,N_2915,N_2851);
xnor UO_371 (O_371,N_2896,N_2940);
nand UO_372 (O_372,N_2978,N_2954);
and UO_373 (O_373,N_2926,N_2918);
xor UO_374 (O_374,N_2881,N_2900);
or UO_375 (O_375,N_2975,N_2967);
xnor UO_376 (O_376,N_2829,N_2912);
nor UO_377 (O_377,N_2921,N_2976);
or UO_378 (O_378,N_2884,N_2893);
and UO_379 (O_379,N_2925,N_2963);
nand UO_380 (O_380,N_2849,N_2976);
and UO_381 (O_381,N_2829,N_2943);
nor UO_382 (O_382,N_2930,N_2890);
xnor UO_383 (O_383,N_2830,N_2808);
or UO_384 (O_384,N_2890,N_2844);
xor UO_385 (O_385,N_2844,N_2971);
nor UO_386 (O_386,N_2900,N_2917);
nand UO_387 (O_387,N_2905,N_2912);
xnor UO_388 (O_388,N_2888,N_2816);
or UO_389 (O_389,N_2820,N_2819);
or UO_390 (O_390,N_2956,N_2804);
xor UO_391 (O_391,N_2970,N_2935);
or UO_392 (O_392,N_2910,N_2960);
xor UO_393 (O_393,N_2819,N_2993);
xor UO_394 (O_394,N_2919,N_2803);
xor UO_395 (O_395,N_2910,N_2915);
or UO_396 (O_396,N_2937,N_2828);
nor UO_397 (O_397,N_2956,N_2940);
nor UO_398 (O_398,N_2933,N_2937);
xor UO_399 (O_399,N_2874,N_2878);
nand UO_400 (O_400,N_2900,N_2929);
and UO_401 (O_401,N_2857,N_2814);
nand UO_402 (O_402,N_2835,N_2816);
xnor UO_403 (O_403,N_2990,N_2997);
or UO_404 (O_404,N_2978,N_2994);
nand UO_405 (O_405,N_2904,N_2873);
xnor UO_406 (O_406,N_2839,N_2929);
and UO_407 (O_407,N_2950,N_2918);
xor UO_408 (O_408,N_2984,N_2904);
nand UO_409 (O_409,N_2975,N_2828);
and UO_410 (O_410,N_2875,N_2879);
and UO_411 (O_411,N_2830,N_2921);
nand UO_412 (O_412,N_2837,N_2994);
and UO_413 (O_413,N_2920,N_2924);
nand UO_414 (O_414,N_2971,N_2957);
and UO_415 (O_415,N_2977,N_2984);
and UO_416 (O_416,N_2884,N_2985);
or UO_417 (O_417,N_2846,N_2879);
xor UO_418 (O_418,N_2952,N_2880);
nor UO_419 (O_419,N_2981,N_2815);
and UO_420 (O_420,N_2953,N_2947);
nor UO_421 (O_421,N_2990,N_2988);
or UO_422 (O_422,N_2987,N_2960);
nand UO_423 (O_423,N_2804,N_2955);
nor UO_424 (O_424,N_2940,N_2902);
or UO_425 (O_425,N_2921,N_2840);
and UO_426 (O_426,N_2983,N_2894);
nor UO_427 (O_427,N_2825,N_2896);
xnor UO_428 (O_428,N_2925,N_2905);
nand UO_429 (O_429,N_2812,N_2806);
or UO_430 (O_430,N_2987,N_2990);
xnor UO_431 (O_431,N_2866,N_2909);
nor UO_432 (O_432,N_2929,N_2847);
xnor UO_433 (O_433,N_2870,N_2979);
xnor UO_434 (O_434,N_2852,N_2959);
nand UO_435 (O_435,N_2955,N_2927);
nor UO_436 (O_436,N_2960,N_2984);
nor UO_437 (O_437,N_2818,N_2846);
xor UO_438 (O_438,N_2930,N_2923);
nor UO_439 (O_439,N_2839,N_2970);
and UO_440 (O_440,N_2848,N_2810);
nand UO_441 (O_441,N_2977,N_2953);
nand UO_442 (O_442,N_2968,N_2879);
and UO_443 (O_443,N_2836,N_2906);
or UO_444 (O_444,N_2838,N_2804);
and UO_445 (O_445,N_2975,N_2958);
or UO_446 (O_446,N_2863,N_2907);
nand UO_447 (O_447,N_2881,N_2822);
nand UO_448 (O_448,N_2973,N_2984);
and UO_449 (O_449,N_2978,N_2993);
nand UO_450 (O_450,N_2914,N_2827);
and UO_451 (O_451,N_2822,N_2897);
and UO_452 (O_452,N_2952,N_2953);
xor UO_453 (O_453,N_2834,N_2908);
or UO_454 (O_454,N_2815,N_2861);
or UO_455 (O_455,N_2913,N_2869);
nand UO_456 (O_456,N_2918,N_2898);
nor UO_457 (O_457,N_2973,N_2864);
nor UO_458 (O_458,N_2975,N_2968);
nor UO_459 (O_459,N_2897,N_2992);
nand UO_460 (O_460,N_2939,N_2936);
xnor UO_461 (O_461,N_2985,N_2863);
xor UO_462 (O_462,N_2988,N_2944);
or UO_463 (O_463,N_2903,N_2827);
or UO_464 (O_464,N_2872,N_2992);
xor UO_465 (O_465,N_2882,N_2823);
xnor UO_466 (O_466,N_2868,N_2844);
nor UO_467 (O_467,N_2856,N_2874);
xor UO_468 (O_468,N_2876,N_2832);
nor UO_469 (O_469,N_2830,N_2891);
nor UO_470 (O_470,N_2991,N_2906);
nor UO_471 (O_471,N_2924,N_2892);
and UO_472 (O_472,N_2879,N_2854);
and UO_473 (O_473,N_2809,N_2970);
and UO_474 (O_474,N_2971,N_2996);
nor UO_475 (O_475,N_2905,N_2959);
nor UO_476 (O_476,N_2877,N_2818);
xor UO_477 (O_477,N_2823,N_2927);
nor UO_478 (O_478,N_2850,N_2860);
nor UO_479 (O_479,N_2973,N_2988);
nand UO_480 (O_480,N_2977,N_2963);
nand UO_481 (O_481,N_2831,N_2983);
nand UO_482 (O_482,N_2903,N_2879);
and UO_483 (O_483,N_2993,N_2960);
or UO_484 (O_484,N_2918,N_2805);
xnor UO_485 (O_485,N_2875,N_2844);
nand UO_486 (O_486,N_2999,N_2869);
and UO_487 (O_487,N_2891,N_2801);
and UO_488 (O_488,N_2933,N_2841);
xnor UO_489 (O_489,N_2859,N_2987);
and UO_490 (O_490,N_2932,N_2916);
xnor UO_491 (O_491,N_2874,N_2966);
and UO_492 (O_492,N_2822,N_2864);
and UO_493 (O_493,N_2908,N_2906);
nor UO_494 (O_494,N_2823,N_2806);
or UO_495 (O_495,N_2967,N_2910);
or UO_496 (O_496,N_2898,N_2899);
nand UO_497 (O_497,N_2960,N_2809);
and UO_498 (O_498,N_2881,N_2859);
nand UO_499 (O_499,N_2959,N_2985);
endmodule