module basic_500_3000_500_40_levels_1xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_227,In_398);
and U1 (N_1,In_224,In_429);
nand U2 (N_2,In_469,In_131);
nor U3 (N_3,In_440,In_42);
or U4 (N_4,In_303,In_100);
and U5 (N_5,In_473,In_185);
nand U6 (N_6,In_156,In_324);
or U7 (N_7,In_233,In_372);
and U8 (N_8,In_310,In_433);
or U9 (N_9,In_408,In_265);
nand U10 (N_10,In_201,In_123);
nand U11 (N_11,In_132,In_441);
or U12 (N_12,In_226,In_490);
or U13 (N_13,In_105,In_190);
or U14 (N_14,In_427,In_395);
nor U15 (N_15,In_68,In_447);
or U16 (N_16,In_421,In_418);
nand U17 (N_17,In_382,In_24);
or U18 (N_18,In_450,In_376);
nor U19 (N_19,In_189,In_225);
and U20 (N_20,In_442,In_322);
xor U21 (N_21,In_195,In_352);
or U22 (N_22,In_448,In_45);
xor U23 (N_23,In_120,In_278);
and U24 (N_24,In_41,In_261);
or U25 (N_25,In_43,In_247);
nor U26 (N_26,In_26,In_173);
xnor U27 (N_27,In_309,In_221);
or U28 (N_28,In_357,In_426);
or U29 (N_29,In_101,In_254);
nor U30 (N_30,In_498,In_468);
and U31 (N_31,In_399,In_204);
nor U32 (N_32,In_35,In_170);
nor U33 (N_33,In_459,In_355);
nand U34 (N_34,In_83,In_428);
nand U35 (N_35,In_104,In_251);
or U36 (N_36,In_242,In_491);
or U37 (N_37,In_419,In_417);
or U38 (N_38,In_219,In_431);
nand U39 (N_39,In_283,In_229);
nor U40 (N_40,In_316,In_333);
nor U41 (N_41,In_400,In_342);
and U42 (N_42,In_177,In_200);
or U43 (N_43,In_55,In_5);
nand U44 (N_44,In_178,In_318);
nand U45 (N_45,In_16,In_307);
nand U46 (N_46,In_304,In_366);
nor U47 (N_47,In_102,In_438);
xor U48 (N_48,In_288,In_263);
or U49 (N_49,In_345,In_133);
and U50 (N_50,In_32,In_160);
and U51 (N_51,In_250,In_69);
and U52 (N_52,In_375,In_82);
nor U53 (N_53,In_205,In_191);
and U54 (N_54,In_404,In_332);
or U55 (N_55,In_302,In_339);
nor U56 (N_56,In_290,In_31);
or U57 (N_57,In_2,In_403);
nor U58 (N_58,In_208,In_381);
nor U59 (N_59,In_358,In_180);
nor U60 (N_60,In_327,In_449);
nor U61 (N_61,In_259,In_161);
nor U62 (N_62,In_60,In_434);
or U63 (N_63,In_108,In_262);
and U64 (N_64,In_58,In_480);
nor U65 (N_65,In_371,In_124);
or U66 (N_66,In_317,In_103);
nor U67 (N_67,In_377,In_413);
and U68 (N_68,In_112,In_174);
nor U69 (N_69,In_236,In_432);
or U70 (N_70,In_127,In_166);
or U71 (N_71,In_489,In_270);
or U72 (N_72,In_153,In_72);
and U73 (N_73,In_467,In_114);
or U74 (N_74,In_485,In_21);
nor U75 (N_75,In_171,In_274);
and U76 (N_76,In_269,In_228);
nor U77 (N_77,N_27,N_60);
or U78 (N_78,In_157,In_115);
nand U79 (N_79,In_57,In_154);
nand U80 (N_80,In_401,In_71);
or U81 (N_81,In_455,In_280);
nand U82 (N_82,In_186,In_70);
nand U83 (N_83,In_240,N_65);
and U84 (N_84,In_281,In_245);
nand U85 (N_85,In_194,In_458);
and U86 (N_86,In_465,In_353);
or U87 (N_87,In_336,In_407);
nand U88 (N_88,In_356,N_40);
or U89 (N_89,In_282,In_414);
or U90 (N_90,N_10,In_496);
and U91 (N_91,In_145,In_59);
nand U92 (N_92,In_135,In_152);
and U93 (N_93,In_392,In_17);
or U94 (N_94,In_143,In_367);
nor U95 (N_95,In_325,In_393);
and U96 (N_96,N_45,In_183);
nor U97 (N_97,In_239,In_477);
nor U98 (N_98,In_37,In_384);
and U99 (N_99,N_21,In_482);
and U100 (N_100,In_271,In_110);
or U101 (N_101,N_5,In_19);
nand U102 (N_102,In_284,In_319);
nand U103 (N_103,N_59,In_39);
or U104 (N_104,In_443,In_4);
and U105 (N_105,In_118,In_142);
nand U106 (N_106,In_292,In_475);
nor U107 (N_107,In_241,In_460);
nor U108 (N_108,N_72,In_217);
and U109 (N_109,In_248,In_78);
or U110 (N_110,In_215,In_40);
nor U111 (N_111,In_453,In_285);
nor U112 (N_112,N_0,In_331);
and U113 (N_113,In_264,In_46);
nand U114 (N_114,In_234,In_246);
nand U115 (N_115,In_207,In_326);
nor U116 (N_116,In_187,N_12);
and U117 (N_117,In_481,In_368);
xnor U118 (N_118,In_409,In_121);
and U119 (N_119,In_232,In_323);
nand U120 (N_120,N_22,N_74);
and U121 (N_121,In_80,In_230);
nand U122 (N_122,In_0,In_23);
or U123 (N_123,In_144,In_53);
nor U124 (N_124,N_57,In_10);
nor U125 (N_125,In_476,N_14);
nand U126 (N_126,In_18,In_54);
and U127 (N_127,In_463,In_391);
nor U128 (N_128,In_163,In_420);
or U129 (N_129,In_91,In_196);
and U130 (N_130,N_55,N_67);
nor U131 (N_131,In_430,In_125);
and U132 (N_132,In_328,In_62);
and U133 (N_133,In_47,In_478);
or U134 (N_134,In_38,N_43);
nor U135 (N_135,In_206,In_13);
nor U136 (N_136,N_71,N_64);
or U137 (N_137,In_79,N_17);
nor U138 (N_138,N_56,In_188);
or U139 (N_139,In_439,N_50);
nand U140 (N_140,In_335,In_343);
and U141 (N_141,In_360,N_26);
or U142 (N_142,In_126,In_97);
nand U143 (N_143,In_67,N_62);
or U144 (N_144,In_378,In_329);
nor U145 (N_145,In_51,In_406);
nor U146 (N_146,In_344,In_484);
and U147 (N_147,In_52,N_24);
and U148 (N_148,In_253,In_373);
and U149 (N_149,In_454,In_330);
nor U150 (N_150,N_93,In_84);
and U151 (N_151,N_75,In_486);
or U152 (N_152,In_425,N_38);
nand U153 (N_153,In_231,In_362);
nand U154 (N_154,In_499,In_483);
and U155 (N_155,In_117,N_61);
and U156 (N_156,In_193,In_155);
nand U157 (N_157,In_89,In_98);
nand U158 (N_158,In_348,In_140);
nand U159 (N_159,In_48,N_135);
nand U160 (N_160,In_122,N_39);
nor U161 (N_161,In_437,In_291);
nand U162 (N_162,In_176,In_275);
and U163 (N_163,N_63,In_15);
nand U164 (N_164,N_89,In_12);
nand U165 (N_165,In_338,N_23);
or U166 (N_166,In_149,N_123);
or U167 (N_167,In_181,In_172);
or U168 (N_168,In_95,In_296);
and U169 (N_169,In_349,In_396);
and U170 (N_170,N_102,In_151);
nand U171 (N_171,In_3,N_139);
nor U172 (N_172,In_92,N_107);
nor U173 (N_173,In_33,In_379);
and U174 (N_174,In_311,In_75);
nor U175 (N_175,N_118,In_457);
nand U176 (N_176,N_120,In_340);
or U177 (N_177,In_93,In_479);
and U178 (N_178,In_472,In_139);
nand U179 (N_179,In_88,In_297);
nand U180 (N_180,N_91,In_198);
and U181 (N_181,N_69,In_249);
and U182 (N_182,In_415,N_68);
nor U183 (N_183,In_64,N_36);
nand U184 (N_184,In_50,N_100);
nand U185 (N_185,In_272,N_70);
or U186 (N_186,N_142,In_308);
nor U187 (N_187,In_111,N_52);
and U188 (N_188,N_16,N_127);
or U189 (N_189,N_81,In_11);
and U190 (N_190,In_107,In_20);
or U191 (N_191,In_199,N_126);
and U192 (N_192,In_119,In_313);
nor U193 (N_193,In_222,In_351);
or U194 (N_194,N_9,N_20);
nor U195 (N_195,N_19,In_8);
nor U196 (N_196,In_446,In_492);
and U197 (N_197,In_87,N_131);
nor U198 (N_198,In_130,In_192);
nand U199 (N_199,In_273,In_106);
nand U200 (N_200,In_168,In_337);
or U201 (N_201,In_203,N_121);
or U202 (N_202,In_14,In_49);
or U203 (N_203,In_354,In_197);
nor U204 (N_204,In_63,N_99);
and U205 (N_205,N_94,N_146);
nor U206 (N_206,N_76,In_487);
nor U207 (N_207,In_364,In_27);
nand U208 (N_208,In_466,N_44);
and U209 (N_209,In_73,N_35);
and U210 (N_210,In_390,In_235);
nor U211 (N_211,In_306,In_294);
and U212 (N_212,In_394,N_2);
or U213 (N_213,N_11,In_445);
or U214 (N_214,In_212,In_169);
and U215 (N_215,N_105,In_471);
and U216 (N_216,In_369,N_148);
or U217 (N_217,In_286,In_138);
nor U218 (N_218,In_244,In_25);
and U219 (N_219,In_202,In_298);
or U220 (N_220,N_101,In_320);
nand U221 (N_221,In_334,In_86);
and U222 (N_222,N_78,In_451);
or U223 (N_223,In_387,N_66);
or U224 (N_224,In_300,In_1);
nand U225 (N_225,N_211,N_172);
nor U226 (N_226,In_30,N_196);
or U227 (N_227,In_488,N_164);
nand U228 (N_228,N_187,In_312);
nor U229 (N_229,In_293,N_109);
nand U230 (N_230,In_165,In_268);
or U231 (N_231,N_1,N_84);
nor U232 (N_232,N_180,N_179);
nor U233 (N_233,N_25,N_6);
nand U234 (N_234,In_494,N_28);
nand U235 (N_235,In_380,N_184);
nor U236 (N_236,N_186,In_223);
nand U237 (N_237,N_223,N_15);
and U238 (N_238,In_94,N_97);
nand U239 (N_239,N_160,In_44);
nand U240 (N_240,N_98,In_346);
and U241 (N_241,In_76,In_444);
and U242 (N_242,In_238,N_4);
or U243 (N_243,In_90,In_9);
or U244 (N_244,In_276,In_65);
or U245 (N_245,In_363,In_411);
or U246 (N_246,N_221,In_61);
nand U247 (N_247,In_159,N_159);
nand U248 (N_248,In_209,In_495);
or U249 (N_249,In_389,N_222);
and U250 (N_250,N_124,N_200);
or U251 (N_251,N_204,In_267);
or U252 (N_252,N_145,N_33);
or U253 (N_253,In_137,N_203);
or U254 (N_254,N_106,In_66);
nand U255 (N_255,N_58,N_217);
and U256 (N_256,N_155,N_46);
nand U257 (N_257,N_212,In_497);
and U258 (N_258,N_53,N_162);
nor U259 (N_259,In_164,In_109);
nand U260 (N_260,In_29,In_405);
and U261 (N_261,In_452,In_116);
nand U262 (N_262,In_218,In_81);
nand U263 (N_263,N_182,N_171);
and U264 (N_264,In_462,N_29);
and U265 (N_265,In_129,N_206);
nor U266 (N_266,N_178,In_162);
nand U267 (N_267,N_140,In_256);
and U268 (N_268,In_128,In_397);
or U269 (N_269,N_138,In_412);
nand U270 (N_270,N_152,N_119);
and U271 (N_271,N_83,N_87);
nand U272 (N_272,In_388,In_359);
and U273 (N_273,N_208,N_13);
nor U274 (N_274,In_22,N_197);
nor U275 (N_275,N_147,N_85);
nor U276 (N_276,N_190,N_137);
nor U277 (N_277,In_85,N_88);
nand U278 (N_278,N_30,N_80);
or U279 (N_279,In_252,N_134);
and U280 (N_280,N_167,In_28);
or U281 (N_281,In_167,N_112);
and U282 (N_282,N_173,In_279);
or U283 (N_283,In_182,In_260);
or U284 (N_284,In_258,In_148);
nand U285 (N_285,In_435,N_32);
and U286 (N_286,In_141,N_201);
xor U287 (N_287,N_210,In_146);
nand U288 (N_288,N_82,N_113);
or U289 (N_289,In_113,In_424);
nor U290 (N_290,In_365,In_402);
nor U291 (N_291,N_205,N_49);
and U292 (N_292,In_370,In_216);
xor U293 (N_293,In_179,In_347);
nand U294 (N_294,N_90,N_77);
nor U295 (N_295,In_383,In_211);
and U296 (N_296,N_166,N_170);
and U297 (N_297,In_257,In_464);
or U298 (N_298,N_96,N_18);
nor U299 (N_299,In_214,In_315);
nand U300 (N_300,N_225,N_267);
nand U301 (N_301,N_185,In_77);
nor U302 (N_302,In_287,N_115);
or U303 (N_303,N_247,N_286);
xnor U304 (N_304,N_193,N_285);
or U305 (N_305,In_314,In_96);
nor U306 (N_306,In_416,N_149);
nor U307 (N_307,N_255,N_296);
or U308 (N_308,In_305,N_275);
nor U309 (N_309,N_272,In_361);
nand U310 (N_310,N_293,N_227);
or U311 (N_311,N_284,N_48);
or U312 (N_312,N_228,N_128);
and U313 (N_313,N_133,N_188);
and U314 (N_314,N_161,N_224);
nor U315 (N_315,N_218,N_290);
and U316 (N_316,In_277,In_374);
xor U317 (N_317,N_283,N_175);
nor U318 (N_318,In_289,N_282);
or U319 (N_319,N_110,N_174);
or U320 (N_320,N_213,N_248);
or U321 (N_321,N_31,N_261);
and U322 (N_322,N_168,In_99);
nand U323 (N_323,N_238,N_111);
and U324 (N_324,N_114,N_158);
and U325 (N_325,In_461,N_181);
or U326 (N_326,N_288,N_258);
nand U327 (N_327,N_279,N_265);
nor U328 (N_328,N_271,N_220);
nor U329 (N_329,N_156,N_243);
nand U330 (N_330,N_299,In_213);
nor U331 (N_331,N_245,N_153);
or U332 (N_332,N_292,N_297);
and U333 (N_333,N_233,N_176);
or U334 (N_334,N_8,N_259);
and U335 (N_335,N_251,N_79);
and U336 (N_336,N_246,N_249);
or U337 (N_337,N_151,N_216);
nor U338 (N_338,N_154,N_287);
and U339 (N_339,In_36,In_474);
nand U340 (N_340,In_423,In_220);
and U341 (N_341,N_163,In_470);
nor U342 (N_342,N_250,N_150);
and U343 (N_343,N_268,N_215);
or U344 (N_344,N_130,N_294);
nand U345 (N_345,N_260,N_207);
nor U346 (N_346,In_56,N_143);
or U347 (N_347,In_7,N_191);
nor U348 (N_348,N_165,N_270);
or U349 (N_349,N_141,N_183);
nor U350 (N_350,N_298,N_189);
nand U351 (N_351,N_240,N_291);
nor U352 (N_352,N_276,N_209);
nor U353 (N_353,In_493,N_194);
nand U354 (N_354,N_232,In_237);
and U355 (N_355,N_34,In_266);
nor U356 (N_356,N_264,N_144);
nand U357 (N_357,In_299,N_236);
nand U358 (N_358,N_7,N_229);
or U359 (N_359,N_214,N_136);
nand U360 (N_360,N_256,In_210);
or U361 (N_361,N_37,N_177);
or U362 (N_362,N_103,N_95);
and U363 (N_363,N_241,In_301);
nor U364 (N_364,In_134,In_436);
or U365 (N_365,N_237,In_34);
nor U366 (N_366,N_239,N_280);
nor U367 (N_367,N_295,N_169);
and U368 (N_368,N_281,In_243);
nand U369 (N_369,N_92,N_73);
or U370 (N_370,In_321,In_74);
nor U371 (N_371,N_263,N_266);
or U372 (N_372,N_122,N_116);
nand U373 (N_373,N_257,In_385);
nor U374 (N_374,N_108,In_386);
nand U375 (N_375,N_370,N_367);
or U376 (N_376,N_344,N_309);
nand U377 (N_377,N_42,N_157);
nor U378 (N_378,N_315,N_350);
or U379 (N_379,N_368,In_295);
nor U380 (N_380,N_372,N_365);
or U381 (N_381,N_278,N_357);
nand U382 (N_382,N_342,N_289);
or U383 (N_383,N_349,N_198);
nand U384 (N_384,N_132,N_320);
or U385 (N_385,N_269,In_147);
or U386 (N_386,N_300,N_242);
nor U387 (N_387,N_333,N_324);
and U388 (N_388,In_341,N_303);
or U389 (N_389,N_369,N_202);
xnor U390 (N_390,N_317,N_319);
nand U391 (N_391,N_117,N_339);
nor U392 (N_392,N_353,N_231);
nor U393 (N_393,N_322,N_199);
or U394 (N_394,N_327,N_373);
and U395 (N_395,N_51,N_311);
and U396 (N_396,N_321,N_374);
and U397 (N_397,N_310,N_331);
nand U398 (N_398,N_341,N_104);
or U399 (N_399,N_336,N_307);
nand U400 (N_400,In_456,In_150);
nor U401 (N_401,In_422,N_371);
nor U402 (N_402,N_304,N_312);
and U403 (N_403,N_323,N_363);
or U404 (N_404,N_325,N_332);
nand U405 (N_405,N_219,N_306);
nor U406 (N_406,N_129,N_329);
and U407 (N_407,N_347,N_355);
or U408 (N_408,In_6,N_328);
and U409 (N_409,N_338,N_308);
and U410 (N_410,N_316,N_86);
nor U411 (N_411,N_340,N_348);
or U412 (N_412,N_366,N_273);
and U413 (N_413,N_314,N_244);
nand U414 (N_414,N_262,N_253);
and U415 (N_415,N_125,N_334);
or U416 (N_416,N_351,N_301);
nand U417 (N_417,N_364,N_345);
nor U418 (N_418,N_234,In_255);
nor U419 (N_419,N_47,N_326);
nor U420 (N_420,N_362,N_359);
nor U421 (N_421,N_226,N_354);
nand U422 (N_422,N_274,N_360);
nand U423 (N_423,In_410,N_305);
nand U424 (N_424,N_195,N_302);
and U425 (N_425,N_335,N_337);
or U426 (N_426,N_252,In_184);
nor U427 (N_427,N_330,N_192);
and U428 (N_428,In_175,In_350);
nor U429 (N_429,N_318,N_277);
nand U430 (N_430,N_358,N_41);
nor U431 (N_431,N_346,In_158);
or U432 (N_432,N_54,N_230);
nor U433 (N_433,N_3,N_313);
or U434 (N_434,In_136,N_254);
nor U435 (N_435,N_361,N_235);
or U436 (N_436,N_356,N_343);
nor U437 (N_437,N_352,N_308);
xnor U438 (N_438,N_198,N_315);
and U439 (N_439,N_355,N_345);
nor U440 (N_440,N_350,N_253);
nand U441 (N_441,N_305,N_350);
and U442 (N_442,N_340,N_117);
nor U443 (N_443,N_330,N_289);
and U444 (N_444,N_129,N_230);
or U445 (N_445,N_318,N_366);
nor U446 (N_446,N_289,N_348);
and U447 (N_447,N_117,N_373);
or U448 (N_448,N_278,N_311);
or U449 (N_449,N_198,N_157);
or U450 (N_450,N_391,N_413);
nor U451 (N_451,N_429,N_442);
nor U452 (N_452,N_408,N_401);
nand U453 (N_453,N_447,N_410);
nor U454 (N_454,N_440,N_431);
and U455 (N_455,N_377,N_448);
and U456 (N_456,N_418,N_376);
nor U457 (N_457,N_427,N_381);
and U458 (N_458,N_382,N_439);
nand U459 (N_459,N_394,N_436);
or U460 (N_460,N_428,N_411);
or U461 (N_461,N_425,N_390);
nor U462 (N_462,N_417,N_443);
or U463 (N_463,N_449,N_416);
and U464 (N_464,N_409,N_423);
nand U465 (N_465,N_446,N_434);
or U466 (N_466,N_397,N_385);
nand U467 (N_467,N_383,N_421);
nand U468 (N_468,N_445,N_414);
and U469 (N_469,N_396,N_402);
and U470 (N_470,N_437,N_404);
and U471 (N_471,N_426,N_392);
nand U472 (N_472,N_380,N_388);
nand U473 (N_473,N_384,N_400);
nand U474 (N_474,N_389,N_379);
or U475 (N_475,N_406,N_386);
or U476 (N_476,N_420,N_415);
nor U477 (N_477,N_430,N_438);
nor U478 (N_478,N_424,N_432);
nand U479 (N_479,N_435,N_412);
nor U480 (N_480,N_398,N_419);
and U481 (N_481,N_387,N_433);
or U482 (N_482,N_444,N_393);
nand U483 (N_483,N_407,N_403);
and U484 (N_484,N_399,N_395);
nor U485 (N_485,N_375,N_405);
nor U486 (N_486,N_441,N_378);
nand U487 (N_487,N_422,N_409);
and U488 (N_488,N_421,N_402);
nor U489 (N_489,N_444,N_438);
nand U490 (N_490,N_446,N_398);
and U491 (N_491,N_403,N_437);
nor U492 (N_492,N_410,N_415);
or U493 (N_493,N_388,N_422);
nand U494 (N_494,N_407,N_393);
nand U495 (N_495,N_400,N_394);
and U496 (N_496,N_399,N_380);
nand U497 (N_497,N_407,N_446);
nor U498 (N_498,N_427,N_426);
or U499 (N_499,N_445,N_427);
xor U500 (N_500,N_442,N_378);
and U501 (N_501,N_435,N_426);
nor U502 (N_502,N_414,N_438);
or U503 (N_503,N_411,N_429);
or U504 (N_504,N_401,N_395);
or U505 (N_505,N_400,N_397);
nor U506 (N_506,N_406,N_393);
and U507 (N_507,N_437,N_384);
xor U508 (N_508,N_431,N_419);
nor U509 (N_509,N_426,N_442);
nor U510 (N_510,N_423,N_386);
nor U511 (N_511,N_394,N_438);
or U512 (N_512,N_402,N_406);
nand U513 (N_513,N_398,N_399);
and U514 (N_514,N_399,N_377);
nor U515 (N_515,N_418,N_405);
nand U516 (N_516,N_401,N_416);
and U517 (N_517,N_383,N_395);
and U518 (N_518,N_379,N_404);
nand U519 (N_519,N_439,N_440);
nor U520 (N_520,N_414,N_399);
or U521 (N_521,N_399,N_415);
and U522 (N_522,N_378,N_433);
nand U523 (N_523,N_405,N_433);
nand U524 (N_524,N_406,N_436);
nor U525 (N_525,N_473,N_517);
nand U526 (N_526,N_523,N_480);
nor U527 (N_527,N_450,N_489);
and U528 (N_528,N_499,N_474);
and U529 (N_529,N_521,N_510);
xnor U530 (N_530,N_464,N_496);
and U531 (N_531,N_505,N_476);
nor U532 (N_532,N_519,N_492);
nor U533 (N_533,N_483,N_468);
nor U534 (N_534,N_479,N_455);
nor U535 (N_535,N_466,N_524);
nand U536 (N_536,N_472,N_513);
nand U537 (N_537,N_498,N_452);
nand U538 (N_538,N_509,N_502);
nor U539 (N_539,N_497,N_456);
nand U540 (N_540,N_462,N_485);
nand U541 (N_541,N_461,N_494);
or U542 (N_542,N_490,N_503);
and U543 (N_543,N_475,N_471);
nor U544 (N_544,N_514,N_465);
and U545 (N_545,N_457,N_454);
nor U546 (N_546,N_463,N_508);
nand U547 (N_547,N_478,N_484);
nor U548 (N_548,N_500,N_460);
or U549 (N_549,N_516,N_491);
nor U550 (N_550,N_470,N_459);
nand U551 (N_551,N_495,N_501);
nand U552 (N_552,N_488,N_467);
nand U553 (N_553,N_511,N_512);
nand U554 (N_554,N_518,N_482);
nand U555 (N_555,N_453,N_451);
nor U556 (N_556,N_469,N_522);
or U557 (N_557,N_520,N_506);
and U558 (N_558,N_515,N_458);
and U559 (N_559,N_493,N_507);
or U560 (N_560,N_481,N_477);
nand U561 (N_561,N_486,N_504);
nor U562 (N_562,N_487,N_485);
nor U563 (N_563,N_516,N_520);
and U564 (N_564,N_502,N_494);
or U565 (N_565,N_513,N_509);
nand U566 (N_566,N_457,N_465);
or U567 (N_567,N_509,N_505);
nand U568 (N_568,N_450,N_474);
nand U569 (N_569,N_478,N_485);
nor U570 (N_570,N_492,N_470);
nand U571 (N_571,N_492,N_474);
or U572 (N_572,N_484,N_522);
or U573 (N_573,N_470,N_471);
nor U574 (N_574,N_518,N_507);
and U575 (N_575,N_524,N_508);
nand U576 (N_576,N_480,N_466);
nor U577 (N_577,N_463,N_475);
nand U578 (N_578,N_472,N_475);
or U579 (N_579,N_458,N_475);
or U580 (N_580,N_503,N_512);
nor U581 (N_581,N_497,N_452);
or U582 (N_582,N_475,N_481);
nand U583 (N_583,N_482,N_462);
nor U584 (N_584,N_477,N_520);
nand U585 (N_585,N_492,N_477);
and U586 (N_586,N_513,N_521);
nor U587 (N_587,N_495,N_513);
nand U588 (N_588,N_513,N_499);
nand U589 (N_589,N_451,N_494);
or U590 (N_590,N_457,N_462);
or U591 (N_591,N_469,N_482);
or U592 (N_592,N_472,N_493);
nand U593 (N_593,N_497,N_509);
nand U594 (N_594,N_455,N_491);
and U595 (N_595,N_451,N_450);
or U596 (N_596,N_462,N_467);
nor U597 (N_597,N_520,N_507);
or U598 (N_598,N_515,N_522);
and U599 (N_599,N_477,N_460);
or U600 (N_600,N_544,N_526);
nor U601 (N_601,N_590,N_565);
and U602 (N_602,N_599,N_534);
and U603 (N_603,N_589,N_593);
and U604 (N_604,N_531,N_561);
or U605 (N_605,N_568,N_564);
nor U606 (N_606,N_556,N_532);
and U607 (N_607,N_555,N_560);
and U608 (N_608,N_582,N_525);
nor U609 (N_609,N_530,N_594);
or U610 (N_610,N_543,N_552);
nand U611 (N_611,N_559,N_537);
or U612 (N_612,N_587,N_569);
nand U613 (N_613,N_570,N_547);
nand U614 (N_614,N_592,N_540);
nor U615 (N_615,N_596,N_550);
nor U616 (N_616,N_539,N_538);
nor U617 (N_617,N_563,N_571);
nor U618 (N_618,N_567,N_533);
and U619 (N_619,N_584,N_529);
nand U620 (N_620,N_595,N_536);
nand U621 (N_621,N_580,N_583);
nand U622 (N_622,N_562,N_557);
nand U623 (N_623,N_574,N_573);
and U624 (N_624,N_542,N_591);
and U625 (N_625,N_554,N_551);
and U626 (N_626,N_578,N_546);
or U627 (N_627,N_553,N_575);
nand U628 (N_628,N_585,N_566);
and U629 (N_629,N_586,N_545);
nor U630 (N_630,N_579,N_558);
nor U631 (N_631,N_527,N_535);
nand U632 (N_632,N_548,N_588);
or U633 (N_633,N_528,N_541);
nand U634 (N_634,N_581,N_572);
or U635 (N_635,N_597,N_577);
nor U636 (N_636,N_549,N_598);
nand U637 (N_637,N_576,N_589);
or U638 (N_638,N_536,N_532);
or U639 (N_639,N_534,N_546);
nor U640 (N_640,N_589,N_580);
nor U641 (N_641,N_573,N_566);
nor U642 (N_642,N_568,N_576);
nor U643 (N_643,N_554,N_542);
nand U644 (N_644,N_548,N_541);
and U645 (N_645,N_562,N_555);
nand U646 (N_646,N_585,N_558);
nor U647 (N_647,N_583,N_568);
nor U648 (N_648,N_584,N_525);
and U649 (N_649,N_597,N_534);
or U650 (N_650,N_563,N_549);
and U651 (N_651,N_587,N_563);
nor U652 (N_652,N_590,N_597);
nor U653 (N_653,N_572,N_574);
and U654 (N_654,N_525,N_579);
nand U655 (N_655,N_570,N_529);
and U656 (N_656,N_564,N_588);
and U657 (N_657,N_568,N_536);
or U658 (N_658,N_571,N_539);
nand U659 (N_659,N_548,N_568);
nand U660 (N_660,N_533,N_562);
nor U661 (N_661,N_570,N_575);
nor U662 (N_662,N_568,N_579);
and U663 (N_663,N_556,N_576);
or U664 (N_664,N_570,N_569);
and U665 (N_665,N_578,N_548);
or U666 (N_666,N_554,N_548);
nand U667 (N_667,N_598,N_572);
nor U668 (N_668,N_562,N_556);
and U669 (N_669,N_577,N_575);
or U670 (N_670,N_566,N_533);
and U671 (N_671,N_585,N_584);
or U672 (N_672,N_539,N_567);
or U673 (N_673,N_587,N_549);
and U674 (N_674,N_593,N_570);
and U675 (N_675,N_611,N_659);
and U676 (N_676,N_612,N_640);
nor U677 (N_677,N_636,N_647);
nand U678 (N_678,N_652,N_623);
and U679 (N_679,N_672,N_641);
nand U680 (N_680,N_667,N_669);
and U681 (N_681,N_646,N_626);
and U682 (N_682,N_605,N_658);
nand U683 (N_683,N_657,N_614);
nand U684 (N_684,N_624,N_666);
or U685 (N_685,N_619,N_653);
nand U686 (N_686,N_638,N_649);
or U687 (N_687,N_637,N_627);
nor U688 (N_688,N_620,N_661);
nand U689 (N_689,N_643,N_645);
nand U690 (N_690,N_601,N_642);
nor U691 (N_691,N_603,N_664);
and U692 (N_692,N_662,N_655);
nor U693 (N_693,N_671,N_656);
nor U694 (N_694,N_670,N_608);
nor U695 (N_695,N_634,N_621);
nor U696 (N_696,N_668,N_628);
nor U697 (N_697,N_633,N_622);
nor U698 (N_698,N_663,N_609);
and U699 (N_699,N_632,N_604);
and U700 (N_700,N_618,N_629);
nor U701 (N_701,N_674,N_660);
and U702 (N_702,N_635,N_625);
nor U703 (N_703,N_648,N_651);
and U704 (N_704,N_600,N_631);
nor U705 (N_705,N_613,N_606);
nand U706 (N_706,N_665,N_650);
nand U707 (N_707,N_630,N_602);
nor U708 (N_708,N_673,N_654);
and U709 (N_709,N_639,N_616);
nand U710 (N_710,N_615,N_610);
nand U711 (N_711,N_644,N_617);
or U712 (N_712,N_607,N_665);
and U713 (N_713,N_661,N_608);
or U714 (N_714,N_635,N_604);
nor U715 (N_715,N_657,N_630);
and U716 (N_716,N_633,N_659);
and U717 (N_717,N_600,N_668);
nor U718 (N_718,N_661,N_633);
and U719 (N_719,N_648,N_629);
or U720 (N_720,N_608,N_605);
or U721 (N_721,N_603,N_644);
nand U722 (N_722,N_663,N_634);
or U723 (N_723,N_622,N_605);
nand U724 (N_724,N_616,N_652);
or U725 (N_725,N_674,N_624);
nand U726 (N_726,N_656,N_606);
and U727 (N_727,N_642,N_668);
or U728 (N_728,N_668,N_636);
and U729 (N_729,N_606,N_653);
nor U730 (N_730,N_629,N_649);
nand U731 (N_731,N_652,N_626);
or U732 (N_732,N_617,N_606);
or U733 (N_733,N_606,N_609);
nand U734 (N_734,N_642,N_623);
or U735 (N_735,N_668,N_631);
or U736 (N_736,N_611,N_670);
nand U737 (N_737,N_662,N_622);
or U738 (N_738,N_604,N_620);
or U739 (N_739,N_600,N_655);
nor U740 (N_740,N_665,N_614);
and U741 (N_741,N_662,N_637);
and U742 (N_742,N_641,N_604);
and U743 (N_743,N_651,N_674);
nand U744 (N_744,N_609,N_615);
nand U745 (N_745,N_633,N_652);
nand U746 (N_746,N_629,N_642);
nor U747 (N_747,N_638,N_626);
and U748 (N_748,N_651,N_662);
nand U749 (N_749,N_657,N_671);
and U750 (N_750,N_724,N_696);
nor U751 (N_751,N_746,N_688);
and U752 (N_752,N_719,N_697);
nor U753 (N_753,N_740,N_713);
and U754 (N_754,N_731,N_711);
nor U755 (N_755,N_698,N_732);
and U756 (N_756,N_705,N_747);
nand U757 (N_757,N_680,N_699);
nand U758 (N_758,N_707,N_725);
nand U759 (N_759,N_690,N_676);
or U760 (N_760,N_745,N_677);
nand U761 (N_761,N_714,N_728);
nand U762 (N_762,N_733,N_718);
nor U763 (N_763,N_727,N_693);
nor U764 (N_764,N_710,N_730);
and U765 (N_765,N_734,N_701);
or U766 (N_766,N_720,N_721);
nor U767 (N_767,N_739,N_679);
nor U768 (N_768,N_729,N_726);
nand U769 (N_769,N_738,N_689);
nand U770 (N_770,N_687,N_685);
nor U771 (N_771,N_700,N_735);
nand U772 (N_772,N_694,N_678);
nand U773 (N_773,N_704,N_692);
nor U774 (N_774,N_686,N_716);
nand U775 (N_775,N_675,N_712);
and U776 (N_776,N_708,N_743);
nor U777 (N_777,N_748,N_736);
and U778 (N_778,N_717,N_744);
nor U779 (N_779,N_742,N_695);
and U780 (N_780,N_706,N_722);
or U781 (N_781,N_715,N_741);
nand U782 (N_782,N_702,N_683);
nand U783 (N_783,N_709,N_737);
or U784 (N_784,N_749,N_684);
nor U785 (N_785,N_681,N_682);
and U786 (N_786,N_723,N_703);
or U787 (N_787,N_691,N_701);
nor U788 (N_788,N_719,N_705);
or U789 (N_789,N_738,N_675);
nand U790 (N_790,N_708,N_726);
nand U791 (N_791,N_698,N_701);
xnor U792 (N_792,N_734,N_682);
nor U793 (N_793,N_696,N_689);
and U794 (N_794,N_708,N_676);
nand U795 (N_795,N_715,N_709);
and U796 (N_796,N_699,N_733);
and U797 (N_797,N_706,N_697);
or U798 (N_798,N_723,N_740);
nor U799 (N_799,N_717,N_732);
and U800 (N_800,N_744,N_741);
nor U801 (N_801,N_743,N_745);
nand U802 (N_802,N_744,N_708);
and U803 (N_803,N_738,N_718);
or U804 (N_804,N_731,N_676);
or U805 (N_805,N_675,N_687);
nand U806 (N_806,N_693,N_706);
and U807 (N_807,N_733,N_726);
or U808 (N_808,N_721,N_708);
or U809 (N_809,N_699,N_731);
or U810 (N_810,N_710,N_709);
nor U811 (N_811,N_687,N_711);
and U812 (N_812,N_730,N_717);
or U813 (N_813,N_684,N_725);
nor U814 (N_814,N_716,N_706);
nand U815 (N_815,N_694,N_732);
and U816 (N_816,N_690,N_726);
or U817 (N_817,N_722,N_707);
xor U818 (N_818,N_747,N_734);
and U819 (N_819,N_700,N_685);
and U820 (N_820,N_722,N_740);
nor U821 (N_821,N_722,N_721);
or U822 (N_822,N_675,N_696);
nand U823 (N_823,N_678,N_693);
or U824 (N_824,N_705,N_714);
nand U825 (N_825,N_774,N_800);
or U826 (N_826,N_803,N_765);
or U827 (N_827,N_788,N_780);
and U828 (N_828,N_758,N_751);
nor U829 (N_829,N_815,N_791);
and U830 (N_830,N_822,N_753);
nor U831 (N_831,N_808,N_790);
nor U832 (N_832,N_811,N_755);
xnor U833 (N_833,N_775,N_817);
nand U834 (N_834,N_759,N_816);
or U835 (N_835,N_792,N_754);
or U836 (N_836,N_784,N_781);
or U837 (N_837,N_763,N_773);
nor U838 (N_838,N_812,N_750);
or U839 (N_839,N_799,N_783);
or U840 (N_840,N_818,N_761);
or U841 (N_841,N_764,N_809);
or U842 (N_842,N_821,N_807);
and U843 (N_843,N_776,N_824);
and U844 (N_844,N_785,N_793);
and U845 (N_845,N_806,N_768);
or U846 (N_846,N_805,N_752);
nand U847 (N_847,N_819,N_771);
or U848 (N_848,N_757,N_801);
and U849 (N_849,N_756,N_786);
nor U850 (N_850,N_770,N_767);
nor U851 (N_851,N_802,N_795);
nand U852 (N_852,N_762,N_777);
nand U853 (N_853,N_794,N_796);
or U854 (N_854,N_782,N_804);
nor U855 (N_855,N_760,N_766);
or U856 (N_856,N_798,N_779);
and U857 (N_857,N_823,N_814);
and U858 (N_858,N_789,N_797);
and U859 (N_859,N_778,N_772);
nor U860 (N_860,N_787,N_810);
and U861 (N_861,N_813,N_820);
and U862 (N_862,N_769,N_805);
xor U863 (N_863,N_786,N_809);
and U864 (N_864,N_789,N_773);
nor U865 (N_865,N_753,N_819);
or U866 (N_866,N_756,N_811);
nor U867 (N_867,N_809,N_819);
nand U868 (N_868,N_750,N_761);
nand U869 (N_869,N_801,N_817);
nand U870 (N_870,N_790,N_755);
nand U871 (N_871,N_774,N_824);
or U872 (N_872,N_796,N_820);
nand U873 (N_873,N_813,N_752);
nor U874 (N_874,N_775,N_753);
nor U875 (N_875,N_789,N_788);
and U876 (N_876,N_808,N_775);
or U877 (N_877,N_813,N_774);
nand U878 (N_878,N_763,N_813);
or U879 (N_879,N_763,N_752);
or U880 (N_880,N_819,N_814);
nand U881 (N_881,N_806,N_777);
or U882 (N_882,N_817,N_773);
xnor U883 (N_883,N_763,N_795);
nand U884 (N_884,N_791,N_812);
nand U885 (N_885,N_758,N_765);
or U886 (N_886,N_769,N_784);
nand U887 (N_887,N_774,N_793);
nor U888 (N_888,N_778,N_761);
and U889 (N_889,N_765,N_807);
or U890 (N_890,N_807,N_774);
nor U891 (N_891,N_822,N_812);
and U892 (N_892,N_763,N_755);
and U893 (N_893,N_801,N_758);
nor U894 (N_894,N_781,N_753);
or U895 (N_895,N_790,N_806);
and U896 (N_896,N_808,N_799);
and U897 (N_897,N_803,N_773);
nor U898 (N_898,N_774,N_752);
nor U899 (N_899,N_813,N_810);
and U900 (N_900,N_852,N_849);
and U901 (N_901,N_851,N_830);
or U902 (N_902,N_835,N_853);
and U903 (N_903,N_861,N_874);
and U904 (N_904,N_884,N_840);
nand U905 (N_905,N_841,N_896);
or U906 (N_906,N_858,N_836);
and U907 (N_907,N_854,N_863);
and U908 (N_908,N_856,N_869);
and U909 (N_909,N_890,N_831);
or U910 (N_910,N_879,N_889);
nand U911 (N_911,N_862,N_897);
nor U912 (N_912,N_825,N_898);
nor U913 (N_913,N_865,N_839);
and U914 (N_914,N_859,N_881);
nand U915 (N_915,N_838,N_883);
and U916 (N_916,N_895,N_891);
nor U917 (N_917,N_844,N_886);
nor U918 (N_918,N_847,N_866);
and U919 (N_919,N_892,N_877);
nor U920 (N_920,N_887,N_826);
or U921 (N_921,N_875,N_864);
nand U922 (N_922,N_885,N_893);
and U923 (N_923,N_850,N_843);
nor U924 (N_924,N_834,N_857);
nand U925 (N_925,N_827,N_876);
nand U926 (N_926,N_837,N_848);
nor U927 (N_927,N_878,N_828);
or U928 (N_928,N_842,N_833);
nand U929 (N_929,N_845,N_867);
nand U930 (N_930,N_872,N_832);
nor U931 (N_931,N_882,N_880);
or U932 (N_932,N_868,N_870);
nand U933 (N_933,N_873,N_855);
or U934 (N_934,N_888,N_829);
nor U935 (N_935,N_894,N_846);
nor U936 (N_936,N_860,N_899);
or U937 (N_937,N_871,N_860);
nand U938 (N_938,N_839,N_880);
nor U939 (N_939,N_867,N_881);
nor U940 (N_940,N_854,N_845);
nand U941 (N_941,N_851,N_863);
and U942 (N_942,N_826,N_841);
nand U943 (N_943,N_876,N_867);
xor U944 (N_944,N_877,N_879);
and U945 (N_945,N_868,N_877);
and U946 (N_946,N_839,N_849);
nand U947 (N_947,N_853,N_882);
or U948 (N_948,N_886,N_876);
and U949 (N_949,N_831,N_837);
nor U950 (N_950,N_862,N_836);
or U951 (N_951,N_832,N_849);
nand U952 (N_952,N_890,N_840);
nor U953 (N_953,N_870,N_845);
or U954 (N_954,N_866,N_858);
and U955 (N_955,N_888,N_884);
nand U956 (N_956,N_880,N_859);
nor U957 (N_957,N_829,N_893);
and U958 (N_958,N_882,N_886);
nor U959 (N_959,N_880,N_883);
and U960 (N_960,N_880,N_866);
nor U961 (N_961,N_884,N_865);
nor U962 (N_962,N_872,N_898);
or U963 (N_963,N_849,N_841);
nand U964 (N_964,N_895,N_835);
or U965 (N_965,N_834,N_876);
or U966 (N_966,N_898,N_868);
nand U967 (N_967,N_894,N_845);
nand U968 (N_968,N_829,N_891);
nor U969 (N_969,N_827,N_860);
nor U970 (N_970,N_847,N_898);
nor U971 (N_971,N_864,N_856);
or U972 (N_972,N_897,N_895);
nor U973 (N_973,N_844,N_827);
nand U974 (N_974,N_866,N_833);
nor U975 (N_975,N_931,N_951);
and U976 (N_976,N_953,N_947);
nand U977 (N_977,N_935,N_950);
and U978 (N_978,N_974,N_957);
and U979 (N_979,N_971,N_945);
nand U980 (N_980,N_913,N_907);
and U981 (N_981,N_970,N_962);
nand U982 (N_982,N_922,N_965);
nand U983 (N_983,N_926,N_900);
nor U984 (N_984,N_927,N_939);
and U985 (N_985,N_929,N_938);
and U986 (N_986,N_952,N_910);
nor U987 (N_987,N_920,N_967);
or U988 (N_988,N_912,N_937);
nand U989 (N_989,N_944,N_940);
nor U990 (N_990,N_905,N_930);
nand U991 (N_991,N_959,N_968);
nor U992 (N_992,N_972,N_936);
and U993 (N_993,N_919,N_955);
and U994 (N_994,N_925,N_973);
nor U995 (N_995,N_921,N_960);
or U996 (N_996,N_943,N_916);
and U997 (N_997,N_963,N_934);
nand U998 (N_998,N_958,N_956);
nor U999 (N_999,N_941,N_917);
nor U1000 (N_1000,N_928,N_903);
nor U1001 (N_1001,N_924,N_954);
nand U1002 (N_1002,N_933,N_948);
nand U1003 (N_1003,N_923,N_942);
or U1004 (N_1004,N_969,N_932);
and U1005 (N_1005,N_946,N_966);
nand U1006 (N_1006,N_902,N_915);
and U1007 (N_1007,N_949,N_904);
and U1008 (N_1008,N_914,N_964);
nor U1009 (N_1009,N_906,N_918);
nand U1010 (N_1010,N_908,N_909);
and U1011 (N_1011,N_901,N_911);
nor U1012 (N_1012,N_961,N_924);
nand U1013 (N_1013,N_970,N_920);
nand U1014 (N_1014,N_965,N_956);
nand U1015 (N_1015,N_940,N_906);
nor U1016 (N_1016,N_911,N_952);
nor U1017 (N_1017,N_967,N_936);
nor U1018 (N_1018,N_955,N_961);
and U1019 (N_1019,N_961,N_964);
nor U1020 (N_1020,N_950,N_965);
and U1021 (N_1021,N_930,N_941);
or U1022 (N_1022,N_943,N_906);
nand U1023 (N_1023,N_926,N_959);
or U1024 (N_1024,N_900,N_903);
nand U1025 (N_1025,N_927,N_918);
nor U1026 (N_1026,N_928,N_922);
nand U1027 (N_1027,N_906,N_932);
nand U1028 (N_1028,N_905,N_921);
and U1029 (N_1029,N_947,N_946);
or U1030 (N_1030,N_963,N_938);
nor U1031 (N_1031,N_908,N_914);
xnor U1032 (N_1032,N_966,N_945);
or U1033 (N_1033,N_952,N_955);
and U1034 (N_1034,N_920,N_937);
nor U1035 (N_1035,N_946,N_948);
nor U1036 (N_1036,N_900,N_972);
nand U1037 (N_1037,N_941,N_967);
nor U1038 (N_1038,N_937,N_917);
or U1039 (N_1039,N_955,N_968);
and U1040 (N_1040,N_922,N_908);
or U1041 (N_1041,N_953,N_945);
and U1042 (N_1042,N_965,N_921);
nor U1043 (N_1043,N_969,N_959);
nor U1044 (N_1044,N_921,N_939);
and U1045 (N_1045,N_958,N_902);
or U1046 (N_1046,N_959,N_913);
and U1047 (N_1047,N_903,N_953);
nor U1048 (N_1048,N_925,N_902);
nand U1049 (N_1049,N_949,N_901);
and U1050 (N_1050,N_982,N_994);
nand U1051 (N_1051,N_979,N_995);
nor U1052 (N_1052,N_1022,N_1019);
nand U1053 (N_1053,N_1042,N_992);
nand U1054 (N_1054,N_980,N_1023);
nand U1055 (N_1055,N_1027,N_1006);
or U1056 (N_1056,N_1005,N_1010);
nor U1057 (N_1057,N_1001,N_1036);
and U1058 (N_1058,N_1048,N_1020);
or U1059 (N_1059,N_1021,N_1029);
or U1060 (N_1060,N_978,N_1043);
nand U1061 (N_1061,N_989,N_993);
or U1062 (N_1062,N_1024,N_1011);
or U1063 (N_1063,N_1003,N_984);
nand U1064 (N_1064,N_975,N_1004);
nor U1065 (N_1065,N_997,N_1044);
nor U1066 (N_1066,N_991,N_987);
nor U1067 (N_1067,N_1013,N_981);
or U1068 (N_1068,N_1015,N_1017);
nand U1069 (N_1069,N_1032,N_1007);
or U1070 (N_1070,N_999,N_1012);
nor U1071 (N_1071,N_1014,N_1039);
nand U1072 (N_1072,N_1028,N_1026);
nand U1073 (N_1073,N_1009,N_998);
and U1074 (N_1074,N_1030,N_988);
nand U1075 (N_1075,N_1016,N_1037);
and U1076 (N_1076,N_1018,N_996);
and U1077 (N_1077,N_1041,N_1033);
and U1078 (N_1078,N_976,N_1031);
or U1079 (N_1079,N_986,N_1038);
and U1080 (N_1080,N_990,N_1047);
nor U1081 (N_1081,N_1008,N_977);
nor U1082 (N_1082,N_1002,N_1034);
and U1083 (N_1083,N_1040,N_1045);
and U1084 (N_1084,N_1049,N_1035);
and U1085 (N_1085,N_983,N_1046);
nor U1086 (N_1086,N_1000,N_1025);
or U1087 (N_1087,N_985,N_1034);
or U1088 (N_1088,N_996,N_1022);
nand U1089 (N_1089,N_979,N_980);
nor U1090 (N_1090,N_983,N_978);
nor U1091 (N_1091,N_1049,N_992);
and U1092 (N_1092,N_997,N_1026);
nor U1093 (N_1093,N_1009,N_979);
and U1094 (N_1094,N_1042,N_1014);
nor U1095 (N_1095,N_1001,N_1002);
nor U1096 (N_1096,N_1015,N_1023);
or U1097 (N_1097,N_1013,N_992);
or U1098 (N_1098,N_1044,N_1019);
nor U1099 (N_1099,N_1023,N_976);
nor U1100 (N_1100,N_1019,N_986);
nor U1101 (N_1101,N_1016,N_986);
xor U1102 (N_1102,N_1012,N_1004);
or U1103 (N_1103,N_1039,N_1030);
and U1104 (N_1104,N_1013,N_1040);
nand U1105 (N_1105,N_1000,N_976);
or U1106 (N_1106,N_1033,N_1011);
nand U1107 (N_1107,N_986,N_987);
nand U1108 (N_1108,N_1013,N_1031);
or U1109 (N_1109,N_1015,N_988);
and U1110 (N_1110,N_978,N_1001);
nor U1111 (N_1111,N_979,N_985);
nor U1112 (N_1112,N_1023,N_1026);
and U1113 (N_1113,N_1034,N_1011);
or U1114 (N_1114,N_987,N_993);
nand U1115 (N_1115,N_1001,N_1023);
or U1116 (N_1116,N_1032,N_1011);
and U1117 (N_1117,N_1019,N_989);
and U1118 (N_1118,N_1004,N_1030);
nor U1119 (N_1119,N_994,N_997);
nor U1120 (N_1120,N_1043,N_1049);
and U1121 (N_1121,N_976,N_1046);
nor U1122 (N_1122,N_998,N_1045);
nand U1123 (N_1123,N_1001,N_1020);
nor U1124 (N_1124,N_1024,N_982);
and U1125 (N_1125,N_1068,N_1124);
nand U1126 (N_1126,N_1092,N_1072);
and U1127 (N_1127,N_1069,N_1113);
nand U1128 (N_1128,N_1108,N_1104);
and U1129 (N_1129,N_1103,N_1074);
nor U1130 (N_1130,N_1089,N_1051);
and U1131 (N_1131,N_1073,N_1061);
nor U1132 (N_1132,N_1081,N_1058);
nand U1133 (N_1133,N_1088,N_1098);
nand U1134 (N_1134,N_1080,N_1071);
or U1135 (N_1135,N_1115,N_1075);
nor U1136 (N_1136,N_1059,N_1105);
nand U1137 (N_1137,N_1120,N_1078);
nand U1138 (N_1138,N_1091,N_1065);
or U1139 (N_1139,N_1063,N_1090);
or U1140 (N_1140,N_1116,N_1070);
or U1141 (N_1141,N_1099,N_1094);
or U1142 (N_1142,N_1112,N_1076);
nand U1143 (N_1143,N_1083,N_1060);
nor U1144 (N_1144,N_1097,N_1117);
or U1145 (N_1145,N_1064,N_1085);
or U1146 (N_1146,N_1119,N_1050);
and U1147 (N_1147,N_1086,N_1122);
nor U1148 (N_1148,N_1077,N_1109);
or U1149 (N_1149,N_1062,N_1067);
and U1150 (N_1150,N_1095,N_1118);
and U1151 (N_1151,N_1110,N_1123);
and U1152 (N_1152,N_1053,N_1096);
and U1153 (N_1153,N_1093,N_1106);
nor U1154 (N_1154,N_1079,N_1082);
nor U1155 (N_1155,N_1052,N_1055);
nand U1156 (N_1156,N_1101,N_1057);
and U1157 (N_1157,N_1111,N_1087);
nor U1158 (N_1158,N_1084,N_1102);
nand U1159 (N_1159,N_1114,N_1056);
nor U1160 (N_1160,N_1121,N_1107);
nor U1161 (N_1161,N_1100,N_1066);
nor U1162 (N_1162,N_1054,N_1122);
nand U1163 (N_1163,N_1090,N_1104);
or U1164 (N_1164,N_1081,N_1100);
nor U1165 (N_1165,N_1090,N_1081);
nand U1166 (N_1166,N_1121,N_1072);
and U1167 (N_1167,N_1095,N_1069);
nor U1168 (N_1168,N_1072,N_1054);
nand U1169 (N_1169,N_1054,N_1104);
nand U1170 (N_1170,N_1103,N_1113);
or U1171 (N_1171,N_1070,N_1064);
nor U1172 (N_1172,N_1052,N_1075);
nor U1173 (N_1173,N_1112,N_1066);
or U1174 (N_1174,N_1109,N_1092);
or U1175 (N_1175,N_1102,N_1104);
or U1176 (N_1176,N_1086,N_1070);
and U1177 (N_1177,N_1105,N_1107);
and U1178 (N_1178,N_1082,N_1060);
nor U1179 (N_1179,N_1092,N_1060);
nor U1180 (N_1180,N_1120,N_1097);
nor U1181 (N_1181,N_1059,N_1066);
nand U1182 (N_1182,N_1124,N_1122);
nor U1183 (N_1183,N_1120,N_1071);
nand U1184 (N_1184,N_1113,N_1082);
nand U1185 (N_1185,N_1123,N_1098);
or U1186 (N_1186,N_1051,N_1072);
or U1187 (N_1187,N_1121,N_1102);
or U1188 (N_1188,N_1051,N_1100);
nand U1189 (N_1189,N_1066,N_1093);
nor U1190 (N_1190,N_1058,N_1070);
nand U1191 (N_1191,N_1060,N_1096);
nor U1192 (N_1192,N_1064,N_1055);
or U1193 (N_1193,N_1114,N_1092);
nand U1194 (N_1194,N_1080,N_1110);
nand U1195 (N_1195,N_1099,N_1058);
and U1196 (N_1196,N_1123,N_1116);
nor U1197 (N_1197,N_1121,N_1114);
and U1198 (N_1198,N_1076,N_1118);
nor U1199 (N_1199,N_1094,N_1065);
and U1200 (N_1200,N_1152,N_1138);
and U1201 (N_1201,N_1181,N_1192);
nor U1202 (N_1202,N_1127,N_1170);
nor U1203 (N_1203,N_1153,N_1149);
or U1204 (N_1204,N_1156,N_1165);
or U1205 (N_1205,N_1185,N_1144);
or U1206 (N_1206,N_1128,N_1133);
or U1207 (N_1207,N_1199,N_1196);
or U1208 (N_1208,N_1174,N_1168);
and U1209 (N_1209,N_1183,N_1132);
and U1210 (N_1210,N_1147,N_1178);
nor U1211 (N_1211,N_1151,N_1136);
nand U1212 (N_1212,N_1190,N_1158);
nor U1213 (N_1213,N_1145,N_1131);
and U1214 (N_1214,N_1126,N_1135);
nand U1215 (N_1215,N_1125,N_1177);
nor U1216 (N_1216,N_1141,N_1173);
or U1217 (N_1217,N_1142,N_1163);
nor U1218 (N_1218,N_1195,N_1197);
and U1219 (N_1219,N_1179,N_1188);
and U1220 (N_1220,N_1159,N_1129);
or U1221 (N_1221,N_1180,N_1193);
nor U1222 (N_1222,N_1171,N_1150);
and U1223 (N_1223,N_1155,N_1137);
or U1224 (N_1224,N_1164,N_1160);
or U1225 (N_1225,N_1161,N_1194);
nand U1226 (N_1226,N_1176,N_1172);
nor U1227 (N_1227,N_1187,N_1169);
xor U1228 (N_1228,N_1186,N_1134);
and U1229 (N_1229,N_1154,N_1143);
nor U1230 (N_1230,N_1175,N_1184);
or U1231 (N_1231,N_1157,N_1198);
nor U1232 (N_1232,N_1191,N_1148);
and U1233 (N_1233,N_1182,N_1162);
nor U1234 (N_1234,N_1189,N_1167);
or U1235 (N_1235,N_1146,N_1139);
or U1236 (N_1236,N_1130,N_1166);
or U1237 (N_1237,N_1140,N_1195);
and U1238 (N_1238,N_1137,N_1147);
nor U1239 (N_1239,N_1144,N_1159);
nor U1240 (N_1240,N_1184,N_1177);
or U1241 (N_1241,N_1198,N_1189);
nand U1242 (N_1242,N_1126,N_1163);
or U1243 (N_1243,N_1127,N_1190);
nand U1244 (N_1244,N_1181,N_1133);
nor U1245 (N_1245,N_1156,N_1194);
or U1246 (N_1246,N_1125,N_1131);
or U1247 (N_1247,N_1130,N_1192);
or U1248 (N_1248,N_1172,N_1170);
nor U1249 (N_1249,N_1129,N_1171);
and U1250 (N_1250,N_1197,N_1199);
or U1251 (N_1251,N_1183,N_1151);
nor U1252 (N_1252,N_1192,N_1160);
nand U1253 (N_1253,N_1167,N_1193);
nor U1254 (N_1254,N_1154,N_1187);
or U1255 (N_1255,N_1180,N_1185);
or U1256 (N_1256,N_1148,N_1149);
nand U1257 (N_1257,N_1152,N_1180);
nand U1258 (N_1258,N_1163,N_1130);
nor U1259 (N_1259,N_1166,N_1156);
nor U1260 (N_1260,N_1152,N_1196);
nand U1261 (N_1261,N_1170,N_1159);
nor U1262 (N_1262,N_1167,N_1132);
or U1263 (N_1263,N_1131,N_1141);
and U1264 (N_1264,N_1181,N_1186);
or U1265 (N_1265,N_1186,N_1195);
nand U1266 (N_1266,N_1171,N_1131);
and U1267 (N_1267,N_1157,N_1129);
or U1268 (N_1268,N_1150,N_1125);
and U1269 (N_1269,N_1162,N_1193);
or U1270 (N_1270,N_1173,N_1143);
nand U1271 (N_1271,N_1185,N_1167);
and U1272 (N_1272,N_1178,N_1150);
nand U1273 (N_1273,N_1190,N_1184);
or U1274 (N_1274,N_1126,N_1198);
nand U1275 (N_1275,N_1217,N_1224);
nor U1276 (N_1276,N_1274,N_1202);
nand U1277 (N_1277,N_1266,N_1213);
and U1278 (N_1278,N_1200,N_1260);
or U1279 (N_1279,N_1259,N_1226);
or U1280 (N_1280,N_1215,N_1245);
nand U1281 (N_1281,N_1242,N_1243);
nand U1282 (N_1282,N_1210,N_1252);
and U1283 (N_1283,N_1256,N_1253);
or U1284 (N_1284,N_1262,N_1227);
or U1285 (N_1285,N_1247,N_1244);
or U1286 (N_1286,N_1235,N_1208);
or U1287 (N_1287,N_1236,N_1269);
or U1288 (N_1288,N_1239,N_1212);
or U1289 (N_1289,N_1232,N_1214);
and U1290 (N_1290,N_1258,N_1268);
nor U1291 (N_1291,N_1203,N_1251);
or U1292 (N_1292,N_1229,N_1267);
nor U1293 (N_1293,N_1237,N_1264);
and U1294 (N_1294,N_1248,N_1206);
and U1295 (N_1295,N_1230,N_1233);
nor U1296 (N_1296,N_1211,N_1270);
or U1297 (N_1297,N_1255,N_1228);
nor U1298 (N_1298,N_1234,N_1231);
nor U1299 (N_1299,N_1263,N_1254);
nand U1300 (N_1300,N_1218,N_1225);
nor U1301 (N_1301,N_1238,N_1222);
nand U1302 (N_1302,N_1257,N_1219);
nand U1303 (N_1303,N_1216,N_1221);
xnor U1304 (N_1304,N_1250,N_1246);
and U1305 (N_1305,N_1265,N_1209);
nor U1306 (N_1306,N_1271,N_1261);
nand U1307 (N_1307,N_1204,N_1273);
nand U1308 (N_1308,N_1201,N_1207);
and U1309 (N_1309,N_1249,N_1223);
or U1310 (N_1310,N_1205,N_1272);
and U1311 (N_1311,N_1240,N_1220);
nand U1312 (N_1312,N_1241,N_1242);
nand U1313 (N_1313,N_1270,N_1259);
or U1314 (N_1314,N_1248,N_1259);
nor U1315 (N_1315,N_1230,N_1270);
nor U1316 (N_1316,N_1256,N_1204);
nor U1317 (N_1317,N_1230,N_1261);
and U1318 (N_1318,N_1220,N_1235);
and U1319 (N_1319,N_1250,N_1260);
nor U1320 (N_1320,N_1223,N_1267);
nor U1321 (N_1321,N_1236,N_1232);
or U1322 (N_1322,N_1236,N_1201);
or U1323 (N_1323,N_1274,N_1210);
or U1324 (N_1324,N_1205,N_1268);
nor U1325 (N_1325,N_1221,N_1266);
and U1326 (N_1326,N_1201,N_1242);
or U1327 (N_1327,N_1273,N_1268);
nor U1328 (N_1328,N_1220,N_1221);
or U1329 (N_1329,N_1210,N_1226);
nor U1330 (N_1330,N_1226,N_1213);
nor U1331 (N_1331,N_1258,N_1207);
or U1332 (N_1332,N_1238,N_1251);
or U1333 (N_1333,N_1243,N_1227);
nand U1334 (N_1334,N_1240,N_1267);
nand U1335 (N_1335,N_1246,N_1254);
or U1336 (N_1336,N_1203,N_1265);
and U1337 (N_1337,N_1253,N_1237);
and U1338 (N_1338,N_1231,N_1244);
nand U1339 (N_1339,N_1261,N_1265);
nor U1340 (N_1340,N_1231,N_1230);
or U1341 (N_1341,N_1211,N_1242);
or U1342 (N_1342,N_1271,N_1202);
nand U1343 (N_1343,N_1209,N_1205);
nor U1344 (N_1344,N_1255,N_1263);
and U1345 (N_1345,N_1270,N_1268);
nand U1346 (N_1346,N_1211,N_1241);
nand U1347 (N_1347,N_1215,N_1272);
and U1348 (N_1348,N_1266,N_1200);
and U1349 (N_1349,N_1273,N_1207);
nor U1350 (N_1350,N_1287,N_1333);
nor U1351 (N_1351,N_1327,N_1323);
and U1352 (N_1352,N_1309,N_1291);
nor U1353 (N_1353,N_1296,N_1302);
nor U1354 (N_1354,N_1278,N_1311);
nor U1355 (N_1355,N_1321,N_1344);
nand U1356 (N_1356,N_1301,N_1328);
nand U1357 (N_1357,N_1322,N_1275);
or U1358 (N_1358,N_1303,N_1337);
and U1359 (N_1359,N_1294,N_1332);
or U1360 (N_1360,N_1293,N_1339);
nand U1361 (N_1361,N_1312,N_1343);
and U1362 (N_1362,N_1326,N_1324);
nand U1363 (N_1363,N_1276,N_1280);
or U1364 (N_1364,N_1330,N_1315);
or U1365 (N_1365,N_1320,N_1283);
or U1366 (N_1366,N_1347,N_1314);
or U1367 (N_1367,N_1308,N_1286);
nand U1368 (N_1368,N_1299,N_1288);
and U1369 (N_1369,N_1349,N_1348);
nand U1370 (N_1370,N_1298,N_1319);
and U1371 (N_1371,N_1346,N_1279);
or U1372 (N_1372,N_1305,N_1310);
nand U1373 (N_1373,N_1325,N_1329);
and U1374 (N_1374,N_1292,N_1306);
and U1375 (N_1375,N_1331,N_1289);
or U1376 (N_1376,N_1316,N_1297);
or U1377 (N_1377,N_1342,N_1285);
or U1378 (N_1378,N_1317,N_1336);
nand U1379 (N_1379,N_1338,N_1345);
nor U1380 (N_1380,N_1334,N_1341);
nor U1381 (N_1381,N_1295,N_1281);
and U1382 (N_1382,N_1277,N_1304);
nor U1383 (N_1383,N_1340,N_1284);
nand U1384 (N_1384,N_1300,N_1290);
nand U1385 (N_1385,N_1335,N_1318);
and U1386 (N_1386,N_1307,N_1313);
nand U1387 (N_1387,N_1282,N_1290);
or U1388 (N_1388,N_1280,N_1329);
and U1389 (N_1389,N_1299,N_1316);
nor U1390 (N_1390,N_1293,N_1292);
nor U1391 (N_1391,N_1323,N_1340);
nor U1392 (N_1392,N_1288,N_1347);
or U1393 (N_1393,N_1278,N_1280);
and U1394 (N_1394,N_1319,N_1325);
and U1395 (N_1395,N_1313,N_1324);
or U1396 (N_1396,N_1312,N_1335);
nor U1397 (N_1397,N_1292,N_1302);
and U1398 (N_1398,N_1341,N_1346);
nand U1399 (N_1399,N_1298,N_1280);
nand U1400 (N_1400,N_1338,N_1339);
or U1401 (N_1401,N_1312,N_1275);
nor U1402 (N_1402,N_1332,N_1328);
nand U1403 (N_1403,N_1330,N_1325);
and U1404 (N_1404,N_1346,N_1327);
and U1405 (N_1405,N_1283,N_1307);
nand U1406 (N_1406,N_1321,N_1300);
nor U1407 (N_1407,N_1341,N_1326);
nor U1408 (N_1408,N_1302,N_1339);
nor U1409 (N_1409,N_1279,N_1327);
nor U1410 (N_1410,N_1312,N_1303);
and U1411 (N_1411,N_1309,N_1343);
and U1412 (N_1412,N_1288,N_1292);
and U1413 (N_1413,N_1333,N_1338);
or U1414 (N_1414,N_1330,N_1301);
or U1415 (N_1415,N_1327,N_1345);
and U1416 (N_1416,N_1322,N_1326);
xnor U1417 (N_1417,N_1314,N_1276);
or U1418 (N_1418,N_1299,N_1329);
and U1419 (N_1419,N_1284,N_1312);
and U1420 (N_1420,N_1320,N_1332);
or U1421 (N_1421,N_1281,N_1342);
or U1422 (N_1422,N_1295,N_1293);
nor U1423 (N_1423,N_1320,N_1291);
nor U1424 (N_1424,N_1326,N_1289);
and U1425 (N_1425,N_1376,N_1389);
nor U1426 (N_1426,N_1367,N_1355);
nor U1427 (N_1427,N_1419,N_1396);
or U1428 (N_1428,N_1393,N_1360);
nand U1429 (N_1429,N_1411,N_1399);
or U1430 (N_1430,N_1363,N_1382);
or U1431 (N_1431,N_1370,N_1416);
or U1432 (N_1432,N_1383,N_1405);
nand U1433 (N_1433,N_1352,N_1421);
nor U1434 (N_1434,N_1354,N_1398);
nand U1435 (N_1435,N_1410,N_1372);
nor U1436 (N_1436,N_1409,N_1423);
nor U1437 (N_1437,N_1353,N_1414);
nand U1438 (N_1438,N_1381,N_1359);
nand U1439 (N_1439,N_1385,N_1412);
nand U1440 (N_1440,N_1418,N_1361);
nand U1441 (N_1441,N_1395,N_1366);
and U1442 (N_1442,N_1386,N_1388);
nor U1443 (N_1443,N_1424,N_1407);
nor U1444 (N_1444,N_1401,N_1377);
or U1445 (N_1445,N_1394,N_1375);
nor U1446 (N_1446,N_1368,N_1415);
and U1447 (N_1447,N_1379,N_1357);
nor U1448 (N_1448,N_1373,N_1408);
nand U1449 (N_1449,N_1391,N_1400);
nor U1450 (N_1450,N_1397,N_1403);
xor U1451 (N_1451,N_1374,N_1417);
or U1452 (N_1452,N_1369,N_1371);
nand U1453 (N_1453,N_1406,N_1378);
and U1454 (N_1454,N_1420,N_1380);
or U1455 (N_1455,N_1413,N_1350);
nor U1456 (N_1456,N_1392,N_1351);
nand U1457 (N_1457,N_1404,N_1384);
or U1458 (N_1458,N_1362,N_1364);
nand U1459 (N_1459,N_1387,N_1356);
and U1460 (N_1460,N_1422,N_1390);
nand U1461 (N_1461,N_1402,N_1358);
nand U1462 (N_1462,N_1365,N_1408);
nand U1463 (N_1463,N_1414,N_1358);
nand U1464 (N_1464,N_1397,N_1358);
or U1465 (N_1465,N_1357,N_1350);
or U1466 (N_1466,N_1423,N_1353);
nor U1467 (N_1467,N_1388,N_1383);
nor U1468 (N_1468,N_1396,N_1403);
and U1469 (N_1469,N_1397,N_1356);
nand U1470 (N_1470,N_1408,N_1378);
and U1471 (N_1471,N_1392,N_1374);
nand U1472 (N_1472,N_1421,N_1403);
nor U1473 (N_1473,N_1389,N_1352);
nor U1474 (N_1474,N_1384,N_1356);
and U1475 (N_1475,N_1396,N_1353);
nor U1476 (N_1476,N_1399,N_1367);
nand U1477 (N_1477,N_1393,N_1361);
or U1478 (N_1478,N_1378,N_1399);
and U1479 (N_1479,N_1362,N_1405);
nor U1480 (N_1480,N_1411,N_1353);
nand U1481 (N_1481,N_1359,N_1369);
and U1482 (N_1482,N_1408,N_1404);
nor U1483 (N_1483,N_1374,N_1361);
nand U1484 (N_1484,N_1422,N_1367);
nand U1485 (N_1485,N_1407,N_1398);
and U1486 (N_1486,N_1417,N_1376);
and U1487 (N_1487,N_1370,N_1373);
nand U1488 (N_1488,N_1357,N_1383);
and U1489 (N_1489,N_1378,N_1404);
nand U1490 (N_1490,N_1390,N_1379);
or U1491 (N_1491,N_1355,N_1397);
nand U1492 (N_1492,N_1360,N_1406);
nor U1493 (N_1493,N_1393,N_1396);
nor U1494 (N_1494,N_1367,N_1381);
and U1495 (N_1495,N_1368,N_1377);
nor U1496 (N_1496,N_1376,N_1354);
nor U1497 (N_1497,N_1391,N_1389);
and U1498 (N_1498,N_1383,N_1411);
nand U1499 (N_1499,N_1361,N_1406);
and U1500 (N_1500,N_1452,N_1455);
or U1501 (N_1501,N_1428,N_1499);
nor U1502 (N_1502,N_1438,N_1462);
nand U1503 (N_1503,N_1433,N_1478);
or U1504 (N_1504,N_1484,N_1457);
nor U1505 (N_1505,N_1430,N_1432);
nor U1506 (N_1506,N_1439,N_1483);
nand U1507 (N_1507,N_1445,N_1450);
and U1508 (N_1508,N_1481,N_1498);
nand U1509 (N_1509,N_1443,N_1431);
nand U1510 (N_1510,N_1464,N_1461);
nand U1511 (N_1511,N_1477,N_1425);
nand U1512 (N_1512,N_1471,N_1492);
and U1513 (N_1513,N_1434,N_1479);
nand U1514 (N_1514,N_1465,N_1447);
nand U1515 (N_1515,N_1426,N_1482);
or U1516 (N_1516,N_1460,N_1444);
and U1517 (N_1517,N_1449,N_1473);
or U1518 (N_1518,N_1436,N_1485);
nand U1519 (N_1519,N_1480,N_1442);
and U1520 (N_1520,N_1441,N_1491);
or U1521 (N_1521,N_1437,N_1497);
nand U1522 (N_1522,N_1458,N_1470);
or U1523 (N_1523,N_1493,N_1495);
nor U1524 (N_1524,N_1469,N_1440);
and U1525 (N_1525,N_1456,N_1466);
or U1526 (N_1526,N_1496,N_1474);
nor U1527 (N_1527,N_1453,N_1476);
nand U1528 (N_1528,N_1468,N_1475);
xnor U1529 (N_1529,N_1494,N_1490);
and U1530 (N_1530,N_1459,N_1435);
nand U1531 (N_1531,N_1467,N_1429);
nand U1532 (N_1532,N_1486,N_1454);
or U1533 (N_1533,N_1488,N_1451);
nor U1534 (N_1534,N_1487,N_1489);
nand U1535 (N_1535,N_1463,N_1446);
or U1536 (N_1536,N_1427,N_1472);
nor U1537 (N_1537,N_1448,N_1436);
or U1538 (N_1538,N_1439,N_1497);
or U1539 (N_1539,N_1443,N_1430);
nor U1540 (N_1540,N_1427,N_1436);
nand U1541 (N_1541,N_1494,N_1469);
or U1542 (N_1542,N_1498,N_1486);
xnor U1543 (N_1543,N_1438,N_1432);
and U1544 (N_1544,N_1428,N_1442);
or U1545 (N_1545,N_1455,N_1494);
and U1546 (N_1546,N_1429,N_1470);
nand U1547 (N_1547,N_1434,N_1457);
or U1548 (N_1548,N_1433,N_1427);
nand U1549 (N_1549,N_1429,N_1456);
and U1550 (N_1550,N_1467,N_1455);
or U1551 (N_1551,N_1471,N_1447);
and U1552 (N_1552,N_1433,N_1447);
and U1553 (N_1553,N_1481,N_1462);
nand U1554 (N_1554,N_1437,N_1449);
nand U1555 (N_1555,N_1476,N_1440);
nor U1556 (N_1556,N_1432,N_1433);
and U1557 (N_1557,N_1495,N_1478);
or U1558 (N_1558,N_1462,N_1492);
and U1559 (N_1559,N_1494,N_1442);
or U1560 (N_1560,N_1455,N_1453);
nor U1561 (N_1561,N_1447,N_1439);
nor U1562 (N_1562,N_1472,N_1445);
nor U1563 (N_1563,N_1487,N_1499);
nor U1564 (N_1564,N_1496,N_1430);
and U1565 (N_1565,N_1492,N_1444);
or U1566 (N_1566,N_1471,N_1460);
nor U1567 (N_1567,N_1460,N_1432);
nor U1568 (N_1568,N_1497,N_1452);
nor U1569 (N_1569,N_1480,N_1430);
nand U1570 (N_1570,N_1431,N_1488);
nor U1571 (N_1571,N_1451,N_1427);
nor U1572 (N_1572,N_1431,N_1450);
nand U1573 (N_1573,N_1438,N_1465);
or U1574 (N_1574,N_1478,N_1455);
nor U1575 (N_1575,N_1543,N_1514);
nor U1576 (N_1576,N_1537,N_1541);
or U1577 (N_1577,N_1521,N_1550);
nor U1578 (N_1578,N_1569,N_1508);
and U1579 (N_1579,N_1532,N_1562);
nor U1580 (N_1580,N_1566,N_1552);
nor U1581 (N_1581,N_1561,N_1564);
nand U1582 (N_1582,N_1542,N_1555);
or U1583 (N_1583,N_1529,N_1500);
nor U1584 (N_1584,N_1571,N_1505);
or U1585 (N_1585,N_1524,N_1570);
or U1586 (N_1586,N_1517,N_1553);
and U1587 (N_1587,N_1506,N_1557);
or U1588 (N_1588,N_1530,N_1559);
and U1589 (N_1589,N_1560,N_1522);
nor U1590 (N_1590,N_1503,N_1545);
nor U1591 (N_1591,N_1515,N_1533);
nor U1592 (N_1592,N_1540,N_1527);
nor U1593 (N_1593,N_1520,N_1504);
nor U1594 (N_1594,N_1546,N_1534);
or U1595 (N_1595,N_1554,N_1516);
nand U1596 (N_1596,N_1544,N_1501);
and U1597 (N_1597,N_1519,N_1509);
nand U1598 (N_1598,N_1573,N_1572);
or U1599 (N_1599,N_1535,N_1525);
nor U1600 (N_1600,N_1538,N_1563);
nand U1601 (N_1601,N_1548,N_1531);
or U1602 (N_1602,N_1511,N_1507);
and U1603 (N_1603,N_1567,N_1526);
nand U1604 (N_1604,N_1547,N_1558);
and U1605 (N_1605,N_1513,N_1510);
and U1606 (N_1606,N_1518,N_1574);
nand U1607 (N_1607,N_1556,N_1502);
and U1608 (N_1608,N_1523,N_1551);
nand U1609 (N_1609,N_1539,N_1536);
nand U1610 (N_1610,N_1549,N_1528);
nand U1611 (N_1611,N_1512,N_1565);
or U1612 (N_1612,N_1568,N_1537);
and U1613 (N_1613,N_1519,N_1542);
or U1614 (N_1614,N_1539,N_1557);
nand U1615 (N_1615,N_1546,N_1502);
or U1616 (N_1616,N_1537,N_1556);
nor U1617 (N_1617,N_1516,N_1525);
or U1618 (N_1618,N_1523,N_1550);
nand U1619 (N_1619,N_1534,N_1519);
nor U1620 (N_1620,N_1518,N_1548);
nand U1621 (N_1621,N_1528,N_1530);
nor U1622 (N_1622,N_1550,N_1548);
and U1623 (N_1623,N_1550,N_1559);
nor U1624 (N_1624,N_1512,N_1513);
or U1625 (N_1625,N_1509,N_1525);
nor U1626 (N_1626,N_1502,N_1537);
or U1627 (N_1627,N_1534,N_1526);
nor U1628 (N_1628,N_1523,N_1538);
and U1629 (N_1629,N_1567,N_1512);
and U1630 (N_1630,N_1533,N_1512);
nor U1631 (N_1631,N_1507,N_1517);
or U1632 (N_1632,N_1546,N_1572);
nor U1633 (N_1633,N_1573,N_1530);
and U1634 (N_1634,N_1568,N_1536);
nor U1635 (N_1635,N_1547,N_1548);
or U1636 (N_1636,N_1527,N_1550);
and U1637 (N_1637,N_1572,N_1543);
and U1638 (N_1638,N_1516,N_1569);
and U1639 (N_1639,N_1502,N_1504);
or U1640 (N_1640,N_1545,N_1511);
nand U1641 (N_1641,N_1544,N_1526);
or U1642 (N_1642,N_1567,N_1520);
xor U1643 (N_1643,N_1552,N_1543);
nor U1644 (N_1644,N_1548,N_1552);
nand U1645 (N_1645,N_1522,N_1535);
nor U1646 (N_1646,N_1570,N_1561);
nor U1647 (N_1647,N_1522,N_1516);
nand U1648 (N_1648,N_1522,N_1561);
nand U1649 (N_1649,N_1564,N_1520);
and U1650 (N_1650,N_1631,N_1644);
or U1651 (N_1651,N_1615,N_1617);
or U1652 (N_1652,N_1639,N_1575);
or U1653 (N_1653,N_1621,N_1590);
nor U1654 (N_1654,N_1589,N_1637);
or U1655 (N_1655,N_1606,N_1580);
nor U1656 (N_1656,N_1649,N_1586);
or U1657 (N_1657,N_1636,N_1635);
nor U1658 (N_1658,N_1600,N_1638);
nand U1659 (N_1659,N_1612,N_1581);
or U1660 (N_1660,N_1611,N_1576);
nand U1661 (N_1661,N_1629,N_1595);
nand U1662 (N_1662,N_1607,N_1609);
nor U1663 (N_1663,N_1632,N_1646);
nor U1664 (N_1664,N_1630,N_1613);
and U1665 (N_1665,N_1588,N_1587);
nor U1666 (N_1666,N_1608,N_1624);
nand U1667 (N_1667,N_1594,N_1596);
nand U1668 (N_1668,N_1599,N_1578);
or U1669 (N_1669,N_1625,N_1614);
or U1670 (N_1670,N_1620,N_1601);
and U1671 (N_1671,N_1642,N_1605);
nor U1672 (N_1672,N_1641,N_1640);
nor U1673 (N_1673,N_1623,N_1633);
and U1674 (N_1674,N_1592,N_1598);
or U1675 (N_1675,N_1622,N_1579);
or U1676 (N_1676,N_1584,N_1619);
nor U1677 (N_1677,N_1582,N_1593);
nor U1678 (N_1678,N_1648,N_1585);
and U1679 (N_1679,N_1645,N_1597);
nor U1680 (N_1680,N_1627,N_1583);
nand U1681 (N_1681,N_1591,N_1628);
and U1682 (N_1682,N_1616,N_1634);
and U1683 (N_1683,N_1602,N_1577);
nor U1684 (N_1684,N_1604,N_1603);
nand U1685 (N_1685,N_1647,N_1626);
nand U1686 (N_1686,N_1610,N_1643);
nor U1687 (N_1687,N_1618,N_1593);
nand U1688 (N_1688,N_1642,N_1625);
or U1689 (N_1689,N_1589,N_1587);
and U1690 (N_1690,N_1593,N_1599);
or U1691 (N_1691,N_1639,N_1584);
nor U1692 (N_1692,N_1609,N_1589);
or U1693 (N_1693,N_1604,N_1598);
or U1694 (N_1694,N_1610,N_1589);
and U1695 (N_1695,N_1635,N_1605);
or U1696 (N_1696,N_1649,N_1580);
and U1697 (N_1697,N_1632,N_1620);
nor U1698 (N_1698,N_1633,N_1579);
and U1699 (N_1699,N_1630,N_1645);
xor U1700 (N_1700,N_1644,N_1630);
nor U1701 (N_1701,N_1639,N_1641);
or U1702 (N_1702,N_1629,N_1592);
nor U1703 (N_1703,N_1630,N_1592);
or U1704 (N_1704,N_1595,N_1604);
and U1705 (N_1705,N_1617,N_1621);
or U1706 (N_1706,N_1632,N_1590);
or U1707 (N_1707,N_1575,N_1633);
nor U1708 (N_1708,N_1592,N_1581);
nor U1709 (N_1709,N_1588,N_1589);
nor U1710 (N_1710,N_1636,N_1633);
or U1711 (N_1711,N_1586,N_1634);
xnor U1712 (N_1712,N_1645,N_1576);
and U1713 (N_1713,N_1618,N_1581);
and U1714 (N_1714,N_1585,N_1581);
nor U1715 (N_1715,N_1604,N_1637);
nand U1716 (N_1716,N_1619,N_1641);
or U1717 (N_1717,N_1629,N_1577);
nor U1718 (N_1718,N_1591,N_1579);
nand U1719 (N_1719,N_1595,N_1599);
nor U1720 (N_1720,N_1634,N_1587);
nand U1721 (N_1721,N_1591,N_1609);
nor U1722 (N_1722,N_1634,N_1603);
nand U1723 (N_1723,N_1577,N_1596);
or U1724 (N_1724,N_1587,N_1603);
or U1725 (N_1725,N_1722,N_1683);
and U1726 (N_1726,N_1721,N_1714);
or U1727 (N_1727,N_1658,N_1681);
nor U1728 (N_1728,N_1663,N_1709);
xnor U1729 (N_1729,N_1675,N_1720);
or U1730 (N_1730,N_1716,N_1673);
nand U1731 (N_1731,N_1678,N_1655);
and U1732 (N_1732,N_1704,N_1657);
nor U1733 (N_1733,N_1687,N_1688);
nand U1734 (N_1734,N_1659,N_1689);
and U1735 (N_1735,N_1672,N_1711);
nand U1736 (N_1736,N_1702,N_1696);
or U1737 (N_1737,N_1706,N_1699);
nand U1738 (N_1738,N_1718,N_1667);
and U1739 (N_1739,N_1693,N_1669);
nor U1740 (N_1740,N_1707,N_1692);
nor U1741 (N_1741,N_1694,N_1705);
or U1742 (N_1742,N_1710,N_1682);
nor U1743 (N_1743,N_1713,N_1679);
and U1744 (N_1744,N_1690,N_1674);
or U1745 (N_1745,N_1654,N_1651);
nand U1746 (N_1746,N_1680,N_1712);
or U1747 (N_1747,N_1671,N_1650);
nand U1748 (N_1748,N_1700,N_1715);
or U1749 (N_1749,N_1717,N_1676);
nand U1750 (N_1750,N_1684,N_1668);
nand U1751 (N_1751,N_1665,N_1666);
nand U1752 (N_1752,N_1685,N_1701);
and U1753 (N_1753,N_1691,N_1724);
nor U1754 (N_1754,N_1697,N_1695);
xnor U1755 (N_1755,N_1719,N_1670);
nor U1756 (N_1756,N_1686,N_1653);
nor U1757 (N_1757,N_1656,N_1723);
or U1758 (N_1758,N_1664,N_1703);
nor U1759 (N_1759,N_1652,N_1661);
nor U1760 (N_1760,N_1708,N_1662);
nand U1761 (N_1761,N_1660,N_1698);
and U1762 (N_1762,N_1677,N_1723);
nand U1763 (N_1763,N_1704,N_1663);
or U1764 (N_1764,N_1688,N_1659);
nand U1765 (N_1765,N_1667,N_1700);
or U1766 (N_1766,N_1668,N_1670);
nor U1767 (N_1767,N_1664,N_1656);
and U1768 (N_1768,N_1723,N_1679);
nor U1769 (N_1769,N_1682,N_1680);
nand U1770 (N_1770,N_1696,N_1700);
nand U1771 (N_1771,N_1688,N_1680);
and U1772 (N_1772,N_1680,N_1655);
nand U1773 (N_1773,N_1719,N_1710);
or U1774 (N_1774,N_1659,N_1699);
or U1775 (N_1775,N_1656,N_1721);
and U1776 (N_1776,N_1724,N_1697);
nand U1777 (N_1777,N_1673,N_1667);
or U1778 (N_1778,N_1689,N_1680);
nor U1779 (N_1779,N_1688,N_1672);
and U1780 (N_1780,N_1675,N_1677);
nor U1781 (N_1781,N_1704,N_1670);
and U1782 (N_1782,N_1700,N_1716);
or U1783 (N_1783,N_1692,N_1689);
nand U1784 (N_1784,N_1685,N_1712);
nand U1785 (N_1785,N_1678,N_1716);
nand U1786 (N_1786,N_1705,N_1654);
or U1787 (N_1787,N_1680,N_1686);
or U1788 (N_1788,N_1694,N_1673);
or U1789 (N_1789,N_1674,N_1652);
nand U1790 (N_1790,N_1669,N_1697);
nor U1791 (N_1791,N_1709,N_1700);
or U1792 (N_1792,N_1672,N_1682);
and U1793 (N_1793,N_1667,N_1693);
nand U1794 (N_1794,N_1696,N_1712);
nor U1795 (N_1795,N_1654,N_1684);
or U1796 (N_1796,N_1724,N_1707);
nor U1797 (N_1797,N_1666,N_1674);
and U1798 (N_1798,N_1709,N_1666);
and U1799 (N_1799,N_1686,N_1650);
nor U1800 (N_1800,N_1751,N_1767);
nor U1801 (N_1801,N_1780,N_1736);
or U1802 (N_1802,N_1779,N_1788);
and U1803 (N_1803,N_1755,N_1789);
and U1804 (N_1804,N_1733,N_1745);
nand U1805 (N_1805,N_1783,N_1749);
or U1806 (N_1806,N_1746,N_1738);
nand U1807 (N_1807,N_1762,N_1758);
nor U1808 (N_1808,N_1790,N_1765);
nor U1809 (N_1809,N_1782,N_1792);
nor U1810 (N_1810,N_1768,N_1781);
and U1811 (N_1811,N_1770,N_1798);
or U1812 (N_1812,N_1771,N_1743);
nor U1813 (N_1813,N_1747,N_1754);
or U1814 (N_1814,N_1763,N_1761);
nand U1815 (N_1815,N_1730,N_1752);
or U1816 (N_1816,N_1795,N_1793);
nor U1817 (N_1817,N_1744,N_1799);
nor U1818 (N_1818,N_1772,N_1791);
and U1819 (N_1819,N_1740,N_1750);
and U1820 (N_1820,N_1737,N_1784);
and U1821 (N_1821,N_1766,N_1753);
or U1822 (N_1822,N_1748,N_1794);
and U1823 (N_1823,N_1777,N_1726);
or U1824 (N_1824,N_1760,N_1773);
nand U1825 (N_1825,N_1786,N_1797);
or U1826 (N_1826,N_1742,N_1739);
and U1827 (N_1827,N_1734,N_1796);
or U1828 (N_1828,N_1775,N_1759);
nand U1829 (N_1829,N_1728,N_1727);
and U1830 (N_1830,N_1787,N_1725);
nor U1831 (N_1831,N_1731,N_1776);
or U1832 (N_1832,N_1778,N_1729);
nand U1833 (N_1833,N_1785,N_1764);
nor U1834 (N_1834,N_1769,N_1756);
or U1835 (N_1835,N_1741,N_1757);
or U1836 (N_1836,N_1732,N_1774);
nor U1837 (N_1837,N_1735,N_1745);
nand U1838 (N_1838,N_1746,N_1787);
nand U1839 (N_1839,N_1763,N_1736);
nor U1840 (N_1840,N_1798,N_1772);
nor U1841 (N_1841,N_1782,N_1785);
and U1842 (N_1842,N_1731,N_1732);
nand U1843 (N_1843,N_1727,N_1784);
nand U1844 (N_1844,N_1773,N_1751);
and U1845 (N_1845,N_1731,N_1764);
or U1846 (N_1846,N_1729,N_1738);
nor U1847 (N_1847,N_1769,N_1790);
and U1848 (N_1848,N_1731,N_1744);
and U1849 (N_1849,N_1770,N_1759);
or U1850 (N_1850,N_1793,N_1745);
nand U1851 (N_1851,N_1757,N_1791);
nor U1852 (N_1852,N_1759,N_1761);
xor U1853 (N_1853,N_1777,N_1742);
nand U1854 (N_1854,N_1788,N_1757);
or U1855 (N_1855,N_1772,N_1794);
and U1856 (N_1856,N_1799,N_1774);
and U1857 (N_1857,N_1730,N_1727);
and U1858 (N_1858,N_1758,N_1751);
nand U1859 (N_1859,N_1765,N_1779);
or U1860 (N_1860,N_1735,N_1795);
or U1861 (N_1861,N_1792,N_1737);
or U1862 (N_1862,N_1785,N_1735);
or U1863 (N_1863,N_1783,N_1797);
nor U1864 (N_1864,N_1796,N_1789);
or U1865 (N_1865,N_1790,N_1782);
and U1866 (N_1866,N_1758,N_1733);
nand U1867 (N_1867,N_1769,N_1734);
and U1868 (N_1868,N_1780,N_1779);
nand U1869 (N_1869,N_1796,N_1752);
or U1870 (N_1870,N_1781,N_1792);
nor U1871 (N_1871,N_1778,N_1794);
and U1872 (N_1872,N_1775,N_1788);
nand U1873 (N_1873,N_1735,N_1740);
or U1874 (N_1874,N_1751,N_1730);
nor U1875 (N_1875,N_1864,N_1844);
nor U1876 (N_1876,N_1867,N_1805);
or U1877 (N_1877,N_1810,N_1824);
and U1878 (N_1878,N_1817,N_1804);
nand U1879 (N_1879,N_1830,N_1865);
nand U1880 (N_1880,N_1872,N_1852);
or U1881 (N_1881,N_1838,N_1871);
and U1882 (N_1882,N_1851,N_1858);
and U1883 (N_1883,N_1869,N_1808);
and U1884 (N_1884,N_1859,N_1842);
nand U1885 (N_1885,N_1835,N_1821);
and U1886 (N_1886,N_1823,N_1801);
or U1887 (N_1887,N_1803,N_1863);
nand U1888 (N_1888,N_1857,N_1822);
and U1889 (N_1889,N_1828,N_1820);
and U1890 (N_1890,N_1839,N_1802);
nand U1891 (N_1891,N_1846,N_1816);
nor U1892 (N_1892,N_1848,N_1850);
and U1893 (N_1893,N_1831,N_1836);
nor U1894 (N_1894,N_1837,N_1870);
nor U1895 (N_1895,N_1826,N_1855);
nand U1896 (N_1896,N_1833,N_1840);
or U1897 (N_1897,N_1849,N_1847);
and U1898 (N_1898,N_1809,N_1800);
nor U1899 (N_1899,N_1829,N_1827);
nand U1900 (N_1900,N_1819,N_1866);
and U1901 (N_1901,N_1825,N_1841);
nand U1902 (N_1902,N_1807,N_1853);
and U1903 (N_1903,N_1818,N_1873);
nor U1904 (N_1904,N_1813,N_1856);
nor U1905 (N_1905,N_1860,N_1834);
nand U1906 (N_1906,N_1868,N_1812);
or U1907 (N_1907,N_1815,N_1806);
nand U1908 (N_1908,N_1862,N_1874);
nor U1909 (N_1909,N_1811,N_1832);
and U1910 (N_1910,N_1814,N_1861);
and U1911 (N_1911,N_1845,N_1854);
or U1912 (N_1912,N_1843,N_1813);
nor U1913 (N_1913,N_1849,N_1824);
nand U1914 (N_1914,N_1824,N_1822);
and U1915 (N_1915,N_1821,N_1837);
nand U1916 (N_1916,N_1804,N_1854);
nand U1917 (N_1917,N_1867,N_1841);
and U1918 (N_1918,N_1810,N_1873);
and U1919 (N_1919,N_1832,N_1854);
nand U1920 (N_1920,N_1873,N_1849);
and U1921 (N_1921,N_1810,N_1839);
nand U1922 (N_1922,N_1820,N_1868);
nand U1923 (N_1923,N_1843,N_1817);
and U1924 (N_1924,N_1861,N_1869);
nor U1925 (N_1925,N_1801,N_1825);
nand U1926 (N_1926,N_1846,N_1860);
and U1927 (N_1927,N_1821,N_1868);
or U1928 (N_1928,N_1856,N_1848);
nand U1929 (N_1929,N_1826,N_1808);
nor U1930 (N_1930,N_1805,N_1838);
nor U1931 (N_1931,N_1815,N_1801);
or U1932 (N_1932,N_1853,N_1809);
nand U1933 (N_1933,N_1857,N_1827);
or U1934 (N_1934,N_1820,N_1806);
or U1935 (N_1935,N_1853,N_1806);
or U1936 (N_1936,N_1869,N_1864);
nand U1937 (N_1937,N_1813,N_1857);
or U1938 (N_1938,N_1870,N_1826);
nor U1939 (N_1939,N_1855,N_1863);
or U1940 (N_1940,N_1869,N_1805);
nand U1941 (N_1941,N_1814,N_1822);
nor U1942 (N_1942,N_1800,N_1857);
or U1943 (N_1943,N_1818,N_1817);
nand U1944 (N_1944,N_1831,N_1856);
nor U1945 (N_1945,N_1805,N_1821);
nand U1946 (N_1946,N_1847,N_1841);
nor U1947 (N_1947,N_1834,N_1818);
nand U1948 (N_1948,N_1825,N_1843);
nor U1949 (N_1949,N_1853,N_1863);
nand U1950 (N_1950,N_1940,N_1944);
and U1951 (N_1951,N_1928,N_1933);
or U1952 (N_1952,N_1878,N_1947);
nor U1953 (N_1953,N_1922,N_1886);
and U1954 (N_1954,N_1916,N_1925);
nand U1955 (N_1955,N_1924,N_1901);
nor U1956 (N_1956,N_1929,N_1879);
nor U1957 (N_1957,N_1949,N_1895);
nor U1958 (N_1958,N_1926,N_1918);
and U1959 (N_1959,N_1875,N_1939);
nand U1960 (N_1960,N_1883,N_1907);
or U1961 (N_1961,N_1911,N_1876);
nand U1962 (N_1962,N_1936,N_1881);
nor U1963 (N_1963,N_1885,N_1904);
nor U1964 (N_1964,N_1896,N_1931);
nand U1965 (N_1965,N_1880,N_1914);
or U1966 (N_1966,N_1934,N_1905);
and U1967 (N_1967,N_1902,N_1898);
and U1968 (N_1968,N_1908,N_1891);
and U1969 (N_1969,N_1892,N_1913);
nor U1970 (N_1970,N_1909,N_1943);
nand U1971 (N_1971,N_1877,N_1919);
and U1972 (N_1972,N_1948,N_1946);
or U1973 (N_1973,N_1889,N_1882);
or U1974 (N_1974,N_1912,N_1887);
nor U1975 (N_1975,N_1903,N_1945);
nor U1976 (N_1976,N_1897,N_1921);
nor U1977 (N_1977,N_1894,N_1927);
nor U1978 (N_1978,N_1937,N_1917);
or U1979 (N_1979,N_1910,N_1941);
nor U1980 (N_1980,N_1900,N_1920);
or U1981 (N_1981,N_1906,N_1938);
and U1982 (N_1982,N_1893,N_1915);
nand U1983 (N_1983,N_1942,N_1935);
and U1984 (N_1984,N_1890,N_1932);
or U1985 (N_1985,N_1899,N_1888);
or U1986 (N_1986,N_1930,N_1884);
nor U1987 (N_1987,N_1923,N_1924);
and U1988 (N_1988,N_1925,N_1941);
nor U1989 (N_1989,N_1892,N_1915);
or U1990 (N_1990,N_1905,N_1941);
and U1991 (N_1991,N_1880,N_1900);
and U1992 (N_1992,N_1928,N_1941);
nor U1993 (N_1993,N_1948,N_1880);
and U1994 (N_1994,N_1897,N_1914);
nand U1995 (N_1995,N_1904,N_1948);
or U1996 (N_1996,N_1932,N_1948);
and U1997 (N_1997,N_1911,N_1899);
nor U1998 (N_1998,N_1897,N_1901);
and U1999 (N_1999,N_1889,N_1921);
nand U2000 (N_2000,N_1916,N_1880);
and U2001 (N_2001,N_1928,N_1927);
and U2002 (N_2002,N_1891,N_1895);
or U2003 (N_2003,N_1892,N_1943);
nand U2004 (N_2004,N_1885,N_1888);
and U2005 (N_2005,N_1907,N_1936);
or U2006 (N_2006,N_1934,N_1918);
or U2007 (N_2007,N_1887,N_1907);
or U2008 (N_2008,N_1933,N_1922);
nand U2009 (N_2009,N_1931,N_1917);
nor U2010 (N_2010,N_1918,N_1875);
nand U2011 (N_2011,N_1926,N_1897);
or U2012 (N_2012,N_1897,N_1929);
or U2013 (N_2013,N_1917,N_1895);
nor U2014 (N_2014,N_1880,N_1879);
nand U2015 (N_2015,N_1946,N_1930);
nand U2016 (N_2016,N_1928,N_1913);
or U2017 (N_2017,N_1926,N_1933);
nand U2018 (N_2018,N_1947,N_1894);
and U2019 (N_2019,N_1888,N_1895);
nor U2020 (N_2020,N_1886,N_1949);
and U2021 (N_2021,N_1876,N_1891);
or U2022 (N_2022,N_1914,N_1878);
or U2023 (N_2023,N_1946,N_1881);
nand U2024 (N_2024,N_1888,N_1908);
nand U2025 (N_2025,N_2009,N_1993);
nand U2026 (N_2026,N_1996,N_2016);
and U2027 (N_2027,N_1989,N_1995);
and U2028 (N_2028,N_2022,N_1984);
and U2029 (N_2029,N_1961,N_1974);
and U2030 (N_2030,N_2019,N_2024);
nor U2031 (N_2031,N_1972,N_2011);
or U2032 (N_2032,N_1978,N_1990);
and U2033 (N_2033,N_1960,N_1980);
nand U2034 (N_2034,N_1977,N_2000);
nand U2035 (N_2035,N_1983,N_1997);
or U2036 (N_2036,N_2010,N_1967);
nor U2037 (N_2037,N_1957,N_2023);
nor U2038 (N_2038,N_1988,N_1981);
and U2039 (N_2039,N_2002,N_1985);
and U2040 (N_2040,N_2015,N_1965);
nand U2041 (N_2041,N_1950,N_1951);
or U2042 (N_2042,N_1982,N_2018);
or U2043 (N_2043,N_1959,N_1964);
and U2044 (N_2044,N_1962,N_1952);
or U2045 (N_2045,N_1954,N_2014);
nand U2046 (N_2046,N_2012,N_2003);
nand U2047 (N_2047,N_1973,N_2006);
nand U2048 (N_2048,N_2007,N_2008);
xnor U2049 (N_2049,N_2021,N_2017);
nor U2050 (N_2050,N_1968,N_2020);
nor U2051 (N_2051,N_1987,N_2001);
nor U2052 (N_2052,N_1958,N_1971);
or U2053 (N_2053,N_2013,N_1956);
nor U2054 (N_2054,N_1998,N_2005);
and U2055 (N_2055,N_1969,N_1975);
or U2056 (N_2056,N_1976,N_1986);
nor U2057 (N_2057,N_1970,N_1955);
nand U2058 (N_2058,N_1953,N_1994);
and U2059 (N_2059,N_1966,N_1991);
and U2060 (N_2060,N_1979,N_1999);
or U2061 (N_2061,N_2004,N_1963);
and U2062 (N_2062,N_1992,N_1997);
or U2063 (N_2063,N_1976,N_2012);
nor U2064 (N_2064,N_1962,N_1956);
nor U2065 (N_2065,N_1994,N_2017);
and U2066 (N_2066,N_2015,N_1971);
nor U2067 (N_2067,N_1984,N_1968);
and U2068 (N_2068,N_1951,N_1955);
and U2069 (N_2069,N_1964,N_2013);
nand U2070 (N_2070,N_1990,N_2022);
and U2071 (N_2071,N_2017,N_1991);
nand U2072 (N_2072,N_2003,N_2005);
or U2073 (N_2073,N_1992,N_1985);
or U2074 (N_2074,N_1995,N_2007);
nand U2075 (N_2075,N_1997,N_1971);
or U2076 (N_2076,N_1970,N_1969);
or U2077 (N_2077,N_1960,N_1952);
and U2078 (N_2078,N_1989,N_1980);
nand U2079 (N_2079,N_2006,N_1951);
or U2080 (N_2080,N_1971,N_2003);
nand U2081 (N_2081,N_1977,N_1983);
or U2082 (N_2082,N_2017,N_1970);
and U2083 (N_2083,N_2012,N_2008);
nand U2084 (N_2084,N_2014,N_2003);
nor U2085 (N_2085,N_1999,N_1983);
and U2086 (N_2086,N_1966,N_2008);
nand U2087 (N_2087,N_1996,N_1967);
or U2088 (N_2088,N_2012,N_1980);
xnor U2089 (N_2089,N_2007,N_1998);
nor U2090 (N_2090,N_2007,N_1950);
nor U2091 (N_2091,N_1958,N_2006);
and U2092 (N_2092,N_2021,N_1999);
and U2093 (N_2093,N_2018,N_1957);
nor U2094 (N_2094,N_1984,N_1995);
and U2095 (N_2095,N_1962,N_1954);
or U2096 (N_2096,N_2016,N_2006);
or U2097 (N_2097,N_1951,N_1997);
nor U2098 (N_2098,N_1984,N_1990);
or U2099 (N_2099,N_2023,N_1956);
nor U2100 (N_2100,N_2062,N_2055);
and U2101 (N_2101,N_2045,N_2040);
or U2102 (N_2102,N_2077,N_2068);
nand U2103 (N_2103,N_2047,N_2048);
and U2104 (N_2104,N_2098,N_2035);
or U2105 (N_2105,N_2075,N_2026);
nand U2106 (N_2106,N_2060,N_2041);
nand U2107 (N_2107,N_2092,N_2063);
or U2108 (N_2108,N_2037,N_2072);
or U2109 (N_2109,N_2029,N_2057);
or U2110 (N_2110,N_2043,N_2085);
nor U2111 (N_2111,N_2086,N_2074);
nor U2112 (N_2112,N_2039,N_2088);
nand U2113 (N_2113,N_2097,N_2051);
or U2114 (N_2114,N_2090,N_2089);
or U2115 (N_2115,N_2065,N_2078);
nand U2116 (N_2116,N_2094,N_2069);
and U2117 (N_2117,N_2064,N_2032);
or U2118 (N_2118,N_2099,N_2030);
nand U2119 (N_2119,N_2087,N_2054);
nand U2120 (N_2120,N_2096,N_2053);
nand U2121 (N_2121,N_2059,N_2083);
and U2122 (N_2122,N_2084,N_2058);
nand U2123 (N_2123,N_2025,N_2076);
and U2124 (N_2124,N_2044,N_2034);
or U2125 (N_2125,N_2079,N_2038);
and U2126 (N_2126,N_2049,N_2071);
and U2127 (N_2127,N_2027,N_2091);
nand U2128 (N_2128,N_2061,N_2080);
nand U2129 (N_2129,N_2042,N_2081);
nand U2130 (N_2130,N_2050,N_2070);
or U2131 (N_2131,N_2052,N_2093);
nor U2132 (N_2132,N_2082,N_2066);
nand U2133 (N_2133,N_2031,N_2095);
nand U2134 (N_2134,N_2033,N_2067);
or U2135 (N_2135,N_2046,N_2028);
and U2136 (N_2136,N_2036,N_2056);
and U2137 (N_2137,N_2073,N_2045);
and U2138 (N_2138,N_2094,N_2048);
nor U2139 (N_2139,N_2077,N_2089);
nand U2140 (N_2140,N_2047,N_2080);
nand U2141 (N_2141,N_2040,N_2068);
and U2142 (N_2142,N_2091,N_2094);
and U2143 (N_2143,N_2077,N_2070);
xor U2144 (N_2144,N_2054,N_2031);
and U2145 (N_2145,N_2074,N_2043);
or U2146 (N_2146,N_2081,N_2052);
and U2147 (N_2147,N_2070,N_2041);
and U2148 (N_2148,N_2075,N_2090);
and U2149 (N_2149,N_2040,N_2050);
nand U2150 (N_2150,N_2068,N_2061);
nand U2151 (N_2151,N_2092,N_2033);
and U2152 (N_2152,N_2035,N_2076);
and U2153 (N_2153,N_2066,N_2063);
nand U2154 (N_2154,N_2050,N_2045);
and U2155 (N_2155,N_2043,N_2090);
or U2156 (N_2156,N_2084,N_2059);
nor U2157 (N_2157,N_2055,N_2035);
nor U2158 (N_2158,N_2090,N_2095);
nand U2159 (N_2159,N_2078,N_2038);
and U2160 (N_2160,N_2063,N_2095);
and U2161 (N_2161,N_2093,N_2071);
and U2162 (N_2162,N_2049,N_2087);
nand U2163 (N_2163,N_2066,N_2050);
and U2164 (N_2164,N_2075,N_2028);
xnor U2165 (N_2165,N_2045,N_2098);
and U2166 (N_2166,N_2032,N_2093);
and U2167 (N_2167,N_2047,N_2050);
or U2168 (N_2168,N_2041,N_2089);
or U2169 (N_2169,N_2029,N_2063);
and U2170 (N_2170,N_2074,N_2097);
and U2171 (N_2171,N_2071,N_2099);
or U2172 (N_2172,N_2094,N_2082);
and U2173 (N_2173,N_2076,N_2087);
and U2174 (N_2174,N_2067,N_2065);
nand U2175 (N_2175,N_2131,N_2166);
and U2176 (N_2176,N_2104,N_2158);
and U2177 (N_2177,N_2163,N_2133);
nor U2178 (N_2178,N_2100,N_2113);
or U2179 (N_2179,N_2140,N_2149);
nor U2180 (N_2180,N_2142,N_2109);
nand U2181 (N_2181,N_2108,N_2112);
nor U2182 (N_2182,N_2107,N_2122);
nor U2183 (N_2183,N_2156,N_2171);
or U2184 (N_2184,N_2119,N_2162);
nand U2185 (N_2185,N_2124,N_2159);
nand U2186 (N_2186,N_2111,N_2164);
nand U2187 (N_2187,N_2139,N_2168);
xor U2188 (N_2188,N_2121,N_2141);
nand U2189 (N_2189,N_2157,N_2127);
and U2190 (N_2190,N_2170,N_2103);
nand U2191 (N_2191,N_2129,N_2155);
nand U2192 (N_2192,N_2172,N_2105);
nor U2193 (N_2193,N_2134,N_2130);
and U2194 (N_2194,N_2146,N_2123);
or U2195 (N_2195,N_2114,N_2143);
nand U2196 (N_2196,N_2151,N_2154);
and U2197 (N_2197,N_2118,N_2102);
or U2198 (N_2198,N_2138,N_2167);
nand U2199 (N_2199,N_2117,N_2115);
or U2200 (N_2200,N_2147,N_2153);
nor U2201 (N_2201,N_2125,N_2126);
or U2202 (N_2202,N_2101,N_2136);
nand U2203 (N_2203,N_2144,N_2116);
or U2204 (N_2204,N_2150,N_2174);
or U2205 (N_2205,N_2128,N_2173);
nor U2206 (N_2206,N_2148,N_2161);
nand U2207 (N_2207,N_2152,N_2165);
xor U2208 (N_2208,N_2106,N_2145);
or U2209 (N_2209,N_2137,N_2110);
or U2210 (N_2210,N_2120,N_2132);
or U2211 (N_2211,N_2135,N_2169);
or U2212 (N_2212,N_2160,N_2129);
nor U2213 (N_2213,N_2134,N_2108);
and U2214 (N_2214,N_2130,N_2170);
nor U2215 (N_2215,N_2101,N_2151);
and U2216 (N_2216,N_2112,N_2104);
and U2217 (N_2217,N_2169,N_2161);
or U2218 (N_2218,N_2111,N_2146);
nor U2219 (N_2219,N_2103,N_2149);
nand U2220 (N_2220,N_2113,N_2102);
xnor U2221 (N_2221,N_2126,N_2101);
or U2222 (N_2222,N_2144,N_2135);
nor U2223 (N_2223,N_2160,N_2125);
nor U2224 (N_2224,N_2140,N_2105);
nand U2225 (N_2225,N_2132,N_2125);
nor U2226 (N_2226,N_2104,N_2129);
nor U2227 (N_2227,N_2148,N_2118);
and U2228 (N_2228,N_2122,N_2113);
nand U2229 (N_2229,N_2174,N_2127);
nor U2230 (N_2230,N_2158,N_2107);
nor U2231 (N_2231,N_2108,N_2131);
nor U2232 (N_2232,N_2105,N_2145);
and U2233 (N_2233,N_2108,N_2145);
nand U2234 (N_2234,N_2140,N_2102);
and U2235 (N_2235,N_2161,N_2147);
or U2236 (N_2236,N_2116,N_2102);
or U2237 (N_2237,N_2122,N_2127);
nor U2238 (N_2238,N_2163,N_2116);
nand U2239 (N_2239,N_2145,N_2150);
nor U2240 (N_2240,N_2166,N_2129);
or U2241 (N_2241,N_2172,N_2120);
nor U2242 (N_2242,N_2149,N_2115);
nor U2243 (N_2243,N_2137,N_2114);
and U2244 (N_2244,N_2141,N_2171);
nand U2245 (N_2245,N_2143,N_2109);
nor U2246 (N_2246,N_2166,N_2124);
nor U2247 (N_2247,N_2100,N_2128);
or U2248 (N_2248,N_2144,N_2140);
or U2249 (N_2249,N_2171,N_2142);
nor U2250 (N_2250,N_2215,N_2231);
and U2251 (N_2251,N_2182,N_2206);
and U2252 (N_2252,N_2208,N_2233);
and U2253 (N_2253,N_2235,N_2177);
and U2254 (N_2254,N_2236,N_2227);
nor U2255 (N_2255,N_2213,N_2230);
or U2256 (N_2256,N_2245,N_2205);
nor U2257 (N_2257,N_2237,N_2232);
nand U2258 (N_2258,N_2176,N_2200);
nand U2259 (N_2259,N_2229,N_2218);
nand U2260 (N_2260,N_2247,N_2226);
nand U2261 (N_2261,N_2241,N_2195);
nor U2262 (N_2262,N_2202,N_2246);
nor U2263 (N_2263,N_2225,N_2201);
or U2264 (N_2264,N_2219,N_2197);
or U2265 (N_2265,N_2224,N_2216);
and U2266 (N_2266,N_2187,N_2199);
or U2267 (N_2267,N_2234,N_2196);
or U2268 (N_2268,N_2239,N_2217);
nor U2269 (N_2269,N_2228,N_2242);
nor U2270 (N_2270,N_2248,N_2175);
nor U2271 (N_2271,N_2179,N_2178);
nand U2272 (N_2272,N_2193,N_2183);
or U2273 (N_2273,N_2204,N_2222);
and U2274 (N_2274,N_2184,N_2189);
nor U2275 (N_2275,N_2192,N_2180);
and U2276 (N_2276,N_2244,N_2181);
and U2277 (N_2277,N_2190,N_2220);
or U2278 (N_2278,N_2186,N_2214);
nor U2279 (N_2279,N_2188,N_2249);
and U2280 (N_2280,N_2221,N_2240);
or U2281 (N_2281,N_2209,N_2210);
nand U2282 (N_2282,N_2185,N_2238);
nand U2283 (N_2283,N_2243,N_2223);
and U2284 (N_2284,N_2207,N_2191);
nor U2285 (N_2285,N_2198,N_2212);
or U2286 (N_2286,N_2194,N_2211);
or U2287 (N_2287,N_2203,N_2230);
or U2288 (N_2288,N_2240,N_2179);
nand U2289 (N_2289,N_2245,N_2210);
and U2290 (N_2290,N_2179,N_2206);
and U2291 (N_2291,N_2206,N_2242);
or U2292 (N_2292,N_2247,N_2223);
or U2293 (N_2293,N_2193,N_2231);
nand U2294 (N_2294,N_2231,N_2216);
nor U2295 (N_2295,N_2238,N_2190);
and U2296 (N_2296,N_2213,N_2229);
nor U2297 (N_2297,N_2177,N_2239);
or U2298 (N_2298,N_2217,N_2178);
or U2299 (N_2299,N_2198,N_2203);
and U2300 (N_2300,N_2194,N_2220);
and U2301 (N_2301,N_2239,N_2197);
and U2302 (N_2302,N_2230,N_2183);
or U2303 (N_2303,N_2197,N_2204);
nand U2304 (N_2304,N_2219,N_2224);
nor U2305 (N_2305,N_2190,N_2188);
nor U2306 (N_2306,N_2217,N_2249);
and U2307 (N_2307,N_2212,N_2245);
or U2308 (N_2308,N_2177,N_2189);
nor U2309 (N_2309,N_2203,N_2219);
nand U2310 (N_2310,N_2176,N_2221);
and U2311 (N_2311,N_2179,N_2218);
or U2312 (N_2312,N_2190,N_2186);
and U2313 (N_2313,N_2222,N_2206);
nor U2314 (N_2314,N_2236,N_2241);
and U2315 (N_2315,N_2188,N_2176);
and U2316 (N_2316,N_2220,N_2211);
or U2317 (N_2317,N_2242,N_2226);
nor U2318 (N_2318,N_2212,N_2248);
or U2319 (N_2319,N_2221,N_2224);
and U2320 (N_2320,N_2232,N_2196);
and U2321 (N_2321,N_2198,N_2233);
nor U2322 (N_2322,N_2199,N_2210);
nand U2323 (N_2323,N_2185,N_2246);
and U2324 (N_2324,N_2246,N_2233);
and U2325 (N_2325,N_2257,N_2321);
nand U2326 (N_2326,N_2260,N_2290);
or U2327 (N_2327,N_2322,N_2270);
or U2328 (N_2328,N_2288,N_2317);
and U2329 (N_2329,N_2273,N_2279);
nand U2330 (N_2330,N_2289,N_2301);
or U2331 (N_2331,N_2266,N_2298);
nand U2332 (N_2332,N_2271,N_2254);
nor U2333 (N_2333,N_2315,N_2280);
nand U2334 (N_2334,N_2305,N_2312);
and U2335 (N_2335,N_2293,N_2284);
nand U2336 (N_2336,N_2275,N_2306);
nand U2337 (N_2337,N_2318,N_2250);
or U2338 (N_2338,N_2292,N_2311);
and U2339 (N_2339,N_2324,N_2302);
nor U2340 (N_2340,N_2303,N_2309);
or U2341 (N_2341,N_2320,N_2308);
nor U2342 (N_2342,N_2296,N_2262);
nor U2343 (N_2343,N_2251,N_2272);
nor U2344 (N_2344,N_2300,N_2252);
or U2345 (N_2345,N_2263,N_2299);
nand U2346 (N_2346,N_2310,N_2268);
and U2347 (N_2347,N_2287,N_2261);
nor U2348 (N_2348,N_2286,N_2253);
nand U2349 (N_2349,N_2276,N_2269);
nor U2350 (N_2350,N_2278,N_2291);
nor U2351 (N_2351,N_2264,N_2319);
nand U2352 (N_2352,N_2285,N_2316);
or U2353 (N_2353,N_2265,N_2255);
nand U2354 (N_2354,N_2313,N_2282);
nand U2355 (N_2355,N_2274,N_2281);
nand U2356 (N_2356,N_2277,N_2258);
or U2357 (N_2357,N_2283,N_2323);
nand U2358 (N_2358,N_2307,N_2267);
or U2359 (N_2359,N_2297,N_2256);
nor U2360 (N_2360,N_2295,N_2259);
and U2361 (N_2361,N_2294,N_2314);
or U2362 (N_2362,N_2304,N_2268);
and U2363 (N_2363,N_2317,N_2278);
nand U2364 (N_2364,N_2290,N_2317);
or U2365 (N_2365,N_2308,N_2319);
or U2366 (N_2366,N_2304,N_2292);
and U2367 (N_2367,N_2317,N_2271);
or U2368 (N_2368,N_2323,N_2287);
nand U2369 (N_2369,N_2319,N_2252);
nor U2370 (N_2370,N_2301,N_2298);
or U2371 (N_2371,N_2289,N_2291);
nor U2372 (N_2372,N_2324,N_2312);
or U2373 (N_2373,N_2288,N_2261);
and U2374 (N_2374,N_2284,N_2290);
xnor U2375 (N_2375,N_2269,N_2307);
or U2376 (N_2376,N_2292,N_2309);
nand U2377 (N_2377,N_2273,N_2284);
and U2378 (N_2378,N_2282,N_2274);
or U2379 (N_2379,N_2278,N_2264);
xnor U2380 (N_2380,N_2263,N_2277);
and U2381 (N_2381,N_2301,N_2320);
nor U2382 (N_2382,N_2282,N_2308);
and U2383 (N_2383,N_2291,N_2265);
or U2384 (N_2384,N_2281,N_2286);
nor U2385 (N_2385,N_2308,N_2278);
and U2386 (N_2386,N_2314,N_2285);
or U2387 (N_2387,N_2281,N_2259);
nand U2388 (N_2388,N_2291,N_2266);
nand U2389 (N_2389,N_2282,N_2281);
nand U2390 (N_2390,N_2316,N_2281);
nor U2391 (N_2391,N_2269,N_2317);
and U2392 (N_2392,N_2272,N_2307);
nor U2393 (N_2393,N_2272,N_2312);
nor U2394 (N_2394,N_2276,N_2258);
or U2395 (N_2395,N_2264,N_2301);
and U2396 (N_2396,N_2309,N_2288);
or U2397 (N_2397,N_2309,N_2306);
nand U2398 (N_2398,N_2305,N_2293);
or U2399 (N_2399,N_2290,N_2287);
nand U2400 (N_2400,N_2375,N_2385);
nand U2401 (N_2401,N_2333,N_2389);
and U2402 (N_2402,N_2395,N_2390);
or U2403 (N_2403,N_2360,N_2370);
nor U2404 (N_2404,N_2338,N_2373);
nor U2405 (N_2405,N_2368,N_2352);
and U2406 (N_2406,N_2386,N_2380);
and U2407 (N_2407,N_2356,N_2359);
nor U2408 (N_2408,N_2398,N_2354);
and U2409 (N_2409,N_2353,N_2345);
nand U2410 (N_2410,N_2342,N_2328);
and U2411 (N_2411,N_2393,N_2343);
or U2412 (N_2412,N_2340,N_2376);
nor U2413 (N_2413,N_2364,N_2326);
nand U2414 (N_2414,N_2388,N_2337);
and U2415 (N_2415,N_2378,N_2365);
nor U2416 (N_2416,N_2355,N_2377);
or U2417 (N_2417,N_2329,N_2361);
nor U2418 (N_2418,N_2341,N_2383);
nor U2419 (N_2419,N_2397,N_2384);
nor U2420 (N_2420,N_2379,N_2346);
and U2421 (N_2421,N_2387,N_2348);
or U2422 (N_2422,N_2339,N_2349);
nor U2423 (N_2423,N_2381,N_2350);
nor U2424 (N_2424,N_2367,N_2331);
nand U2425 (N_2425,N_2347,N_2363);
nor U2426 (N_2426,N_2327,N_2351);
nor U2427 (N_2427,N_2392,N_2332);
nand U2428 (N_2428,N_2372,N_2336);
nor U2429 (N_2429,N_2335,N_2330);
or U2430 (N_2430,N_2394,N_2357);
xor U2431 (N_2431,N_2382,N_2344);
or U2432 (N_2432,N_2334,N_2371);
nor U2433 (N_2433,N_2369,N_2391);
and U2434 (N_2434,N_2374,N_2366);
nor U2435 (N_2435,N_2358,N_2399);
nor U2436 (N_2436,N_2325,N_2362);
and U2437 (N_2437,N_2396,N_2346);
and U2438 (N_2438,N_2370,N_2329);
and U2439 (N_2439,N_2389,N_2399);
and U2440 (N_2440,N_2332,N_2361);
nand U2441 (N_2441,N_2366,N_2337);
and U2442 (N_2442,N_2386,N_2345);
or U2443 (N_2443,N_2337,N_2368);
nor U2444 (N_2444,N_2342,N_2341);
or U2445 (N_2445,N_2383,N_2396);
or U2446 (N_2446,N_2388,N_2333);
nor U2447 (N_2447,N_2333,N_2367);
nand U2448 (N_2448,N_2329,N_2346);
nand U2449 (N_2449,N_2363,N_2382);
nand U2450 (N_2450,N_2363,N_2362);
and U2451 (N_2451,N_2374,N_2387);
nor U2452 (N_2452,N_2344,N_2347);
nand U2453 (N_2453,N_2338,N_2350);
nor U2454 (N_2454,N_2399,N_2393);
nor U2455 (N_2455,N_2357,N_2368);
nor U2456 (N_2456,N_2332,N_2347);
nand U2457 (N_2457,N_2353,N_2350);
or U2458 (N_2458,N_2385,N_2389);
or U2459 (N_2459,N_2396,N_2344);
nor U2460 (N_2460,N_2340,N_2379);
and U2461 (N_2461,N_2392,N_2383);
nor U2462 (N_2462,N_2331,N_2360);
or U2463 (N_2463,N_2390,N_2326);
nand U2464 (N_2464,N_2333,N_2386);
and U2465 (N_2465,N_2375,N_2351);
or U2466 (N_2466,N_2376,N_2395);
nand U2467 (N_2467,N_2370,N_2374);
and U2468 (N_2468,N_2335,N_2385);
or U2469 (N_2469,N_2348,N_2372);
and U2470 (N_2470,N_2338,N_2333);
or U2471 (N_2471,N_2363,N_2375);
nand U2472 (N_2472,N_2351,N_2361);
or U2473 (N_2473,N_2333,N_2390);
and U2474 (N_2474,N_2350,N_2343);
nand U2475 (N_2475,N_2444,N_2430);
or U2476 (N_2476,N_2433,N_2426);
nor U2477 (N_2477,N_2472,N_2402);
nand U2478 (N_2478,N_2417,N_2454);
nor U2479 (N_2479,N_2460,N_2459);
nand U2480 (N_2480,N_2465,N_2400);
and U2481 (N_2481,N_2453,N_2445);
nor U2482 (N_2482,N_2446,N_2405);
and U2483 (N_2483,N_2415,N_2467);
nand U2484 (N_2484,N_2428,N_2423);
and U2485 (N_2485,N_2421,N_2469);
and U2486 (N_2486,N_2447,N_2422);
nand U2487 (N_2487,N_2407,N_2438);
nand U2488 (N_2488,N_2439,N_2424);
or U2489 (N_2489,N_2466,N_2436);
and U2490 (N_2490,N_2456,N_2408);
or U2491 (N_2491,N_2470,N_2471);
or U2492 (N_2492,N_2449,N_2440);
and U2493 (N_2493,N_2410,N_2435);
and U2494 (N_2494,N_2443,N_2427);
nor U2495 (N_2495,N_2437,N_2455);
nor U2496 (N_2496,N_2418,N_2419);
or U2497 (N_2497,N_2463,N_2413);
or U2498 (N_2498,N_2425,N_2432);
nor U2499 (N_2499,N_2429,N_2403);
or U2500 (N_2500,N_2411,N_2404);
and U2501 (N_2501,N_2450,N_2461);
and U2502 (N_2502,N_2431,N_2412);
and U2503 (N_2503,N_2409,N_2434);
and U2504 (N_2504,N_2468,N_2406);
or U2505 (N_2505,N_2442,N_2457);
nand U2506 (N_2506,N_2420,N_2401);
and U2507 (N_2507,N_2474,N_2451);
nand U2508 (N_2508,N_2414,N_2448);
nor U2509 (N_2509,N_2416,N_2462);
and U2510 (N_2510,N_2458,N_2441);
or U2511 (N_2511,N_2473,N_2452);
or U2512 (N_2512,N_2464,N_2459);
and U2513 (N_2513,N_2453,N_2450);
nand U2514 (N_2514,N_2470,N_2442);
or U2515 (N_2515,N_2452,N_2453);
and U2516 (N_2516,N_2465,N_2461);
nand U2517 (N_2517,N_2471,N_2448);
and U2518 (N_2518,N_2457,N_2436);
nor U2519 (N_2519,N_2437,N_2452);
or U2520 (N_2520,N_2412,N_2446);
and U2521 (N_2521,N_2458,N_2451);
or U2522 (N_2522,N_2449,N_2427);
or U2523 (N_2523,N_2456,N_2469);
nand U2524 (N_2524,N_2409,N_2470);
or U2525 (N_2525,N_2450,N_2409);
or U2526 (N_2526,N_2427,N_2435);
or U2527 (N_2527,N_2473,N_2455);
nor U2528 (N_2528,N_2431,N_2411);
nor U2529 (N_2529,N_2423,N_2447);
nor U2530 (N_2530,N_2418,N_2442);
nand U2531 (N_2531,N_2418,N_2468);
and U2532 (N_2532,N_2446,N_2458);
and U2533 (N_2533,N_2429,N_2469);
or U2534 (N_2534,N_2461,N_2413);
nand U2535 (N_2535,N_2442,N_2431);
nor U2536 (N_2536,N_2404,N_2463);
nand U2537 (N_2537,N_2400,N_2432);
or U2538 (N_2538,N_2430,N_2410);
xor U2539 (N_2539,N_2429,N_2434);
or U2540 (N_2540,N_2445,N_2457);
and U2541 (N_2541,N_2410,N_2470);
or U2542 (N_2542,N_2462,N_2425);
or U2543 (N_2543,N_2425,N_2469);
nand U2544 (N_2544,N_2439,N_2441);
and U2545 (N_2545,N_2435,N_2434);
nor U2546 (N_2546,N_2445,N_2454);
or U2547 (N_2547,N_2420,N_2465);
nor U2548 (N_2548,N_2426,N_2410);
or U2549 (N_2549,N_2445,N_2432);
or U2550 (N_2550,N_2531,N_2498);
or U2551 (N_2551,N_2514,N_2483);
nor U2552 (N_2552,N_2523,N_2505);
nor U2553 (N_2553,N_2522,N_2539);
and U2554 (N_2554,N_2548,N_2536);
or U2555 (N_2555,N_2485,N_2532);
nor U2556 (N_2556,N_2544,N_2530);
nor U2557 (N_2557,N_2549,N_2497);
and U2558 (N_2558,N_2494,N_2510);
and U2559 (N_2559,N_2501,N_2487);
nor U2560 (N_2560,N_2534,N_2518);
nand U2561 (N_2561,N_2540,N_2529);
or U2562 (N_2562,N_2499,N_2538);
or U2563 (N_2563,N_2496,N_2517);
or U2564 (N_2564,N_2527,N_2503);
nor U2565 (N_2565,N_2525,N_2486);
and U2566 (N_2566,N_2515,N_2528);
nor U2567 (N_2567,N_2526,N_2512);
and U2568 (N_2568,N_2542,N_2546);
nor U2569 (N_2569,N_2484,N_2533);
nor U2570 (N_2570,N_2490,N_2478);
and U2571 (N_2571,N_2506,N_2492);
nor U2572 (N_2572,N_2502,N_2516);
and U2573 (N_2573,N_2535,N_2475);
and U2574 (N_2574,N_2489,N_2488);
and U2575 (N_2575,N_2477,N_2481);
nor U2576 (N_2576,N_2479,N_2480);
nor U2577 (N_2577,N_2476,N_2508);
nor U2578 (N_2578,N_2524,N_2500);
nor U2579 (N_2579,N_2521,N_2491);
and U2580 (N_2580,N_2482,N_2495);
nand U2581 (N_2581,N_2519,N_2541);
and U2582 (N_2582,N_2543,N_2545);
nor U2583 (N_2583,N_2547,N_2511);
or U2584 (N_2584,N_2520,N_2509);
nor U2585 (N_2585,N_2504,N_2493);
nor U2586 (N_2586,N_2537,N_2507);
and U2587 (N_2587,N_2513,N_2507);
nand U2588 (N_2588,N_2532,N_2498);
xnor U2589 (N_2589,N_2476,N_2506);
nand U2590 (N_2590,N_2478,N_2518);
and U2591 (N_2591,N_2489,N_2497);
and U2592 (N_2592,N_2497,N_2506);
nor U2593 (N_2593,N_2542,N_2489);
or U2594 (N_2594,N_2538,N_2490);
xnor U2595 (N_2595,N_2516,N_2523);
nand U2596 (N_2596,N_2498,N_2476);
nand U2597 (N_2597,N_2516,N_2479);
nor U2598 (N_2598,N_2539,N_2499);
nor U2599 (N_2599,N_2507,N_2502);
or U2600 (N_2600,N_2547,N_2538);
nor U2601 (N_2601,N_2477,N_2527);
and U2602 (N_2602,N_2498,N_2521);
nand U2603 (N_2603,N_2533,N_2482);
nor U2604 (N_2604,N_2484,N_2525);
or U2605 (N_2605,N_2505,N_2511);
nand U2606 (N_2606,N_2502,N_2478);
or U2607 (N_2607,N_2491,N_2477);
nand U2608 (N_2608,N_2500,N_2520);
and U2609 (N_2609,N_2507,N_2481);
nand U2610 (N_2610,N_2502,N_2537);
and U2611 (N_2611,N_2514,N_2508);
or U2612 (N_2612,N_2477,N_2532);
or U2613 (N_2613,N_2516,N_2505);
or U2614 (N_2614,N_2501,N_2549);
nand U2615 (N_2615,N_2478,N_2528);
nor U2616 (N_2616,N_2546,N_2515);
nand U2617 (N_2617,N_2530,N_2522);
and U2618 (N_2618,N_2545,N_2533);
and U2619 (N_2619,N_2497,N_2487);
and U2620 (N_2620,N_2512,N_2485);
and U2621 (N_2621,N_2506,N_2498);
xor U2622 (N_2622,N_2524,N_2491);
or U2623 (N_2623,N_2487,N_2549);
nand U2624 (N_2624,N_2516,N_2512);
and U2625 (N_2625,N_2601,N_2613);
nand U2626 (N_2626,N_2604,N_2574);
and U2627 (N_2627,N_2571,N_2578);
nand U2628 (N_2628,N_2610,N_2553);
or U2629 (N_2629,N_2554,N_2612);
nor U2630 (N_2630,N_2569,N_2570);
and U2631 (N_2631,N_2581,N_2592);
and U2632 (N_2632,N_2596,N_2566);
nor U2633 (N_2633,N_2579,N_2583);
or U2634 (N_2634,N_2588,N_2597);
nor U2635 (N_2635,N_2600,N_2615);
nand U2636 (N_2636,N_2593,N_2564);
or U2637 (N_2637,N_2611,N_2557);
nand U2638 (N_2638,N_2576,N_2614);
nand U2639 (N_2639,N_2552,N_2619);
or U2640 (N_2640,N_2608,N_2594);
or U2641 (N_2641,N_2621,N_2602);
and U2642 (N_2642,N_2584,N_2609);
or U2643 (N_2643,N_2567,N_2573);
or U2644 (N_2644,N_2616,N_2590);
and U2645 (N_2645,N_2559,N_2568);
and U2646 (N_2646,N_2551,N_2580);
nor U2647 (N_2647,N_2562,N_2587);
or U2648 (N_2648,N_2617,N_2577);
nor U2649 (N_2649,N_2624,N_2605);
nor U2650 (N_2650,N_2565,N_2555);
or U2651 (N_2651,N_2620,N_2575);
nand U2652 (N_2652,N_2623,N_2599);
nand U2653 (N_2653,N_2622,N_2595);
nor U2654 (N_2654,N_2550,N_2560);
nand U2655 (N_2655,N_2572,N_2556);
and U2656 (N_2656,N_2561,N_2586);
and U2657 (N_2657,N_2582,N_2618);
or U2658 (N_2658,N_2606,N_2598);
or U2659 (N_2659,N_2585,N_2563);
or U2660 (N_2660,N_2558,N_2603);
and U2661 (N_2661,N_2591,N_2607);
nor U2662 (N_2662,N_2589,N_2602);
nor U2663 (N_2663,N_2599,N_2552);
or U2664 (N_2664,N_2616,N_2569);
nand U2665 (N_2665,N_2612,N_2594);
nor U2666 (N_2666,N_2583,N_2582);
nor U2667 (N_2667,N_2622,N_2593);
nand U2668 (N_2668,N_2604,N_2597);
nand U2669 (N_2669,N_2566,N_2567);
nor U2670 (N_2670,N_2554,N_2568);
and U2671 (N_2671,N_2606,N_2567);
nand U2672 (N_2672,N_2596,N_2578);
nor U2673 (N_2673,N_2582,N_2575);
nand U2674 (N_2674,N_2596,N_2575);
nor U2675 (N_2675,N_2575,N_2601);
or U2676 (N_2676,N_2617,N_2584);
or U2677 (N_2677,N_2585,N_2579);
or U2678 (N_2678,N_2583,N_2595);
or U2679 (N_2679,N_2566,N_2569);
or U2680 (N_2680,N_2619,N_2599);
and U2681 (N_2681,N_2577,N_2610);
nor U2682 (N_2682,N_2581,N_2565);
or U2683 (N_2683,N_2562,N_2601);
and U2684 (N_2684,N_2585,N_2555);
and U2685 (N_2685,N_2607,N_2615);
nand U2686 (N_2686,N_2561,N_2585);
nor U2687 (N_2687,N_2572,N_2598);
nand U2688 (N_2688,N_2572,N_2582);
and U2689 (N_2689,N_2579,N_2561);
nor U2690 (N_2690,N_2608,N_2620);
nor U2691 (N_2691,N_2580,N_2609);
and U2692 (N_2692,N_2551,N_2574);
or U2693 (N_2693,N_2582,N_2585);
nor U2694 (N_2694,N_2593,N_2623);
and U2695 (N_2695,N_2555,N_2597);
or U2696 (N_2696,N_2611,N_2560);
or U2697 (N_2697,N_2594,N_2610);
xor U2698 (N_2698,N_2569,N_2601);
and U2699 (N_2699,N_2588,N_2562);
nor U2700 (N_2700,N_2629,N_2665);
nor U2701 (N_2701,N_2637,N_2675);
and U2702 (N_2702,N_2663,N_2682);
or U2703 (N_2703,N_2680,N_2631);
and U2704 (N_2704,N_2686,N_2681);
nor U2705 (N_2705,N_2633,N_2690);
or U2706 (N_2706,N_2661,N_2687);
nor U2707 (N_2707,N_2669,N_2655);
or U2708 (N_2708,N_2652,N_2668);
and U2709 (N_2709,N_2667,N_2676);
or U2710 (N_2710,N_2648,N_2626);
nor U2711 (N_2711,N_2645,N_2638);
nor U2712 (N_2712,N_2664,N_2674);
nand U2713 (N_2713,N_2679,N_2688);
and U2714 (N_2714,N_2630,N_2653);
nand U2715 (N_2715,N_2698,N_2694);
or U2716 (N_2716,N_2695,N_2697);
and U2717 (N_2717,N_2658,N_2625);
nor U2718 (N_2718,N_2699,N_2639);
nor U2719 (N_2719,N_2660,N_2670);
nand U2720 (N_2720,N_2689,N_2632);
or U2721 (N_2721,N_2642,N_2671);
or U2722 (N_2722,N_2692,N_2659);
or U2723 (N_2723,N_2643,N_2678);
or U2724 (N_2724,N_2628,N_2657);
or U2725 (N_2725,N_2673,N_2662);
nor U2726 (N_2726,N_2634,N_2656);
nand U2727 (N_2727,N_2693,N_2691);
nand U2728 (N_2728,N_2640,N_2644);
nor U2729 (N_2729,N_2684,N_2627);
nor U2730 (N_2730,N_2666,N_2654);
nand U2731 (N_2731,N_2646,N_2649);
and U2732 (N_2732,N_2677,N_2651);
nand U2733 (N_2733,N_2672,N_2636);
and U2734 (N_2734,N_2685,N_2635);
or U2735 (N_2735,N_2641,N_2650);
or U2736 (N_2736,N_2696,N_2647);
nor U2737 (N_2737,N_2683,N_2674);
nor U2738 (N_2738,N_2646,N_2647);
nor U2739 (N_2739,N_2687,N_2698);
and U2740 (N_2740,N_2683,N_2678);
or U2741 (N_2741,N_2662,N_2648);
nor U2742 (N_2742,N_2650,N_2693);
nor U2743 (N_2743,N_2666,N_2628);
and U2744 (N_2744,N_2692,N_2691);
or U2745 (N_2745,N_2647,N_2629);
and U2746 (N_2746,N_2634,N_2625);
nor U2747 (N_2747,N_2648,N_2656);
or U2748 (N_2748,N_2688,N_2644);
or U2749 (N_2749,N_2641,N_2671);
nor U2750 (N_2750,N_2660,N_2682);
or U2751 (N_2751,N_2631,N_2699);
nor U2752 (N_2752,N_2641,N_2687);
nor U2753 (N_2753,N_2688,N_2672);
nor U2754 (N_2754,N_2653,N_2626);
or U2755 (N_2755,N_2686,N_2689);
nor U2756 (N_2756,N_2628,N_2633);
nand U2757 (N_2757,N_2685,N_2667);
nand U2758 (N_2758,N_2633,N_2677);
and U2759 (N_2759,N_2637,N_2673);
nand U2760 (N_2760,N_2651,N_2656);
and U2761 (N_2761,N_2693,N_2678);
nor U2762 (N_2762,N_2645,N_2654);
or U2763 (N_2763,N_2634,N_2676);
nand U2764 (N_2764,N_2625,N_2639);
nand U2765 (N_2765,N_2685,N_2679);
nand U2766 (N_2766,N_2645,N_2673);
nand U2767 (N_2767,N_2667,N_2627);
nand U2768 (N_2768,N_2628,N_2691);
nor U2769 (N_2769,N_2676,N_2646);
nand U2770 (N_2770,N_2630,N_2629);
or U2771 (N_2771,N_2628,N_2625);
and U2772 (N_2772,N_2674,N_2647);
and U2773 (N_2773,N_2685,N_2657);
nor U2774 (N_2774,N_2630,N_2658);
and U2775 (N_2775,N_2726,N_2751);
and U2776 (N_2776,N_2711,N_2744);
or U2777 (N_2777,N_2708,N_2717);
nor U2778 (N_2778,N_2739,N_2704);
nor U2779 (N_2779,N_2705,N_2700);
and U2780 (N_2780,N_2764,N_2719);
or U2781 (N_2781,N_2724,N_2723);
or U2782 (N_2782,N_2727,N_2740);
nor U2783 (N_2783,N_2743,N_2773);
or U2784 (N_2784,N_2734,N_2768);
nor U2785 (N_2785,N_2748,N_2772);
nor U2786 (N_2786,N_2750,N_2712);
nand U2787 (N_2787,N_2756,N_2732);
and U2788 (N_2788,N_2747,N_2753);
nor U2789 (N_2789,N_2725,N_2718);
or U2790 (N_2790,N_2701,N_2755);
and U2791 (N_2791,N_2728,N_2749);
and U2792 (N_2792,N_2702,N_2735);
nand U2793 (N_2793,N_2730,N_2742);
and U2794 (N_2794,N_2738,N_2709);
nor U2795 (N_2795,N_2741,N_2731);
nand U2796 (N_2796,N_2771,N_2745);
nor U2797 (N_2797,N_2757,N_2713);
nand U2798 (N_2798,N_2769,N_2761);
or U2799 (N_2799,N_2716,N_2703);
nand U2800 (N_2800,N_2707,N_2754);
nor U2801 (N_2801,N_2765,N_2733);
nor U2802 (N_2802,N_2762,N_2729);
or U2803 (N_2803,N_2752,N_2722);
or U2804 (N_2804,N_2715,N_2763);
nor U2805 (N_2805,N_2766,N_2706);
or U2806 (N_2806,N_2737,N_2720);
nand U2807 (N_2807,N_2767,N_2759);
nor U2808 (N_2808,N_2774,N_2714);
nand U2809 (N_2809,N_2760,N_2721);
nand U2810 (N_2810,N_2736,N_2758);
and U2811 (N_2811,N_2710,N_2770);
nand U2812 (N_2812,N_2746,N_2736);
nor U2813 (N_2813,N_2771,N_2727);
and U2814 (N_2814,N_2726,N_2761);
xnor U2815 (N_2815,N_2725,N_2757);
or U2816 (N_2816,N_2743,N_2701);
or U2817 (N_2817,N_2707,N_2718);
nor U2818 (N_2818,N_2722,N_2728);
or U2819 (N_2819,N_2760,N_2756);
and U2820 (N_2820,N_2701,N_2708);
nor U2821 (N_2821,N_2735,N_2750);
and U2822 (N_2822,N_2741,N_2745);
or U2823 (N_2823,N_2731,N_2746);
nor U2824 (N_2824,N_2712,N_2735);
nor U2825 (N_2825,N_2714,N_2710);
nor U2826 (N_2826,N_2739,N_2735);
or U2827 (N_2827,N_2765,N_2771);
and U2828 (N_2828,N_2769,N_2725);
or U2829 (N_2829,N_2725,N_2713);
nand U2830 (N_2830,N_2705,N_2747);
or U2831 (N_2831,N_2768,N_2730);
nor U2832 (N_2832,N_2769,N_2726);
nor U2833 (N_2833,N_2757,N_2771);
nand U2834 (N_2834,N_2771,N_2733);
and U2835 (N_2835,N_2702,N_2732);
nand U2836 (N_2836,N_2730,N_2735);
nand U2837 (N_2837,N_2759,N_2751);
or U2838 (N_2838,N_2748,N_2745);
or U2839 (N_2839,N_2763,N_2738);
and U2840 (N_2840,N_2755,N_2718);
nor U2841 (N_2841,N_2730,N_2761);
nand U2842 (N_2842,N_2751,N_2716);
and U2843 (N_2843,N_2735,N_2707);
and U2844 (N_2844,N_2749,N_2733);
and U2845 (N_2845,N_2767,N_2700);
nand U2846 (N_2846,N_2713,N_2728);
or U2847 (N_2847,N_2745,N_2713);
and U2848 (N_2848,N_2706,N_2729);
nor U2849 (N_2849,N_2703,N_2729);
nand U2850 (N_2850,N_2814,N_2801);
nand U2851 (N_2851,N_2812,N_2834);
nor U2852 (N_2852,N_2776,N_2775);
or U2853 (N_2853,N_2789,N_2793);
or U2854 (N_2854,N_2807,N_2795);
nand U2855 (N_2855,N_2839,N_2778);
nand U2856 (N_2856,N_2813,N_2797);
nand U2857 (N_2857,N_2818,N_2830);
nor U2858 (N_2858,N_2802,N_2785);
or U2859 (N_2859,N_2788,N_2835);
and U2860 (N_2860,N_2819,N_2840);
or U2861 (N_2861,N_2846,N_2821);
and U2862 (N_2862,N_2787,N_2845);
nor U2863 (N_2863,N_2796,N_2794);
xnor U2864 (N_2864,N_2843,N_2826);
or U2865 (N_2865,N_2791,N_2780);
nor U2866 (N_2866,N_2833,N_2825);
and U2867 (N_2867,N_2828,N_2810);
or U2868 (N_2868,N_2798,N_2824);
and U2869 (N_2869,N_2790,N_2786);
nand U2870 (N_2870,N_2827,N_2783);
nand U2871 (N_2871,N_2837,N_2809);
or U2872 (N_2872,N_2847,N_2784);
and U2873 (N_2873,N_2808,N_2838);
nor U2874 (N_2874,N_2842,N_2831);
nor U2875 (N_2875,N_2803,N_2829);
or U2876 (N_2876,N_2799,N_2806);
nand U2877 (N_2877,N_2782,N_2848);
or U2878 (N_2878,N_2844,N_2841);
xnor U2879 (N_2879,N_2836,N_2779);
and U2880 (N_2880,N_2811,N_2822);
nand U2881 (N_2881,N_2832,N_2777);
and U2882 (N_2882,N_2820,N_2805);
or U2883 (N_2883,N_2817,N_2849);
or U2884 (N_2884,N_2804,N_2792);
and U2885 (N_2885,N_2800,N_2781);
and U2886 (N_2886,N_2823,N_2816);
nor U2887 (N_2887,N_2815,N_2797);
and U2888 (N_2888,N_2779,N_2819);
nor U2889 (N_2889,N_2792,N_2840);
nand U2890 (N_2890,N_2834,N_2840);
nand U2891 (N_2891,N_2789,N_2831);
or U2892 (N_2892,N_2790,N_2785);
nor U2893 (N_2893,N_2847,N_2824);
nand U2894 (N_2894,N_2802,N_2827);
or U2895 (N_2895,N_2816,N_2809);
nand U2896 (N_2896,N_2834,N_2807);
nor U2897 (N_2897,N_2778,N_2825);
nand U2898 (N_2898,N_2811,N_2839);
and U2899 (N_2899,N_2842,N_2791);
nand U2900 (N_2900,N_2812,N_2801);
and U2901 (N_2901,N_2816,N_2782);
or U2902 (N_2902,N_2775,N_2785);
and U2903 (N_2903,N_2797,N_2835);
or U2904 (N_2904,N_2780,N_2801);
or U2905 (N_2905,N_2805,N_2785);
nand U2906 (N_2906,N_2787,N_2808);
and U2907 (N_2907,N_2834,N_2829);
nand U2908 (N_2908,N_2845,N_2784);
nand U2909 (N_2909,N_2827,N_2816);
or U2910 (N_2910,N_2800,N_2827);
and U2911 (N_2911,N_2780,N_2790);
and U2912 (N_2912,N_2799,N_2835);
nand U2913 (N_2913,N_2835,N_2778);
or U2914 (N_2914,N_2840,N_2832);
or U2915 (N_2915,N_2836,N_2803);
nor U2916 (N_2916,N_2834,N_2777);
and U2917 (N_2917,N_2801,N_2811);
and U2918 (N_2918,N_2818,N_2833);
nand U2919 (N_2919,N_2840,N_2802);
or U2920 (N_2920,N_2801,N_2795);
nor U2921 (N_2921,N_2814,N_2815);
and U2922 (N_2922,N_2846,N_2848);
xnor U2923 (N_2923,N_2812,N_2846);
and U2924 (N_2924,N_2789,N_2829);
nor U2925 (N_2925,N_2921,N_2854);
nand U2926 (N_2926,N_2868,N_2891);
or U2927 (N_2927,N_2855,N_2910);
nand U2928 (N_2928,N_2870,N_2886);
xor U2929 (N_2929,N_2916,N_2889);
nand U2930 (N_2930,N_2904,N_2894);
or U2931 (N_2931,N_2874,N_2873);
nand U2932 (N_2932,N_2917,N_2876);
and U2933 (N_2933,N_2899,N_2901);
and U2934 (N_2934,N_2900,N_2875);
or U2935 (N_2935,N_2853,N_2865);
nor U2936 (N_2936,N_2919,N_2863);
or U2937 (N_2937,N_2903,N_2914);
nor U2938 (N_2938,N_2915,N_2907);
and U2939 (N_2939,N_2882,N_2906);
nand U2940 (N_2940,N_2869,N_2883);
nor U2941 (N_2941,N_2866,N_2893);
or U2942 (N_2942,N_2892,N_2872);
nand U2943 (N_2943,N_2871,N_2922);
nand U2944 (N_2944,N_2890,N_2905);
or U2945 (N_2945,N_2858,N_2908);
or U2946 (N_2946,N_2920,N_2911);
and U2947 (N_2947,N_2881,N_2867);
and U2948 (N_2948,N_2850,N_2909);
or U2949 (N_2949,N_2896,N_2884);
or U2950 (N_2950,N_2898,N_2913);
and U2951 (N_2951,N_2878,N_2862);
and U2952 (N_2952,N_2924,N_2859);
nor U2953 (N_2953,N_2860,N_2888);
or U2954 (N_2954,N_2885,N_2877);
nor U2955 (N_2955,N_2861,N_2902);
or U2956 (N_2956,N_2879,N_2923);
nor U2957 (N_2957,N_2887,N_2912);
or U2958 (N_2958,N_2895,N_2918);
or U2959 (N_2959,N_2864,N_2856);
nor U2960 (N_2960,N_2857,N_2880);
nand U2961 (N_2961,N_2851,N_2852);
and U2962 (N_2962,N_2897,N_2885);
or U2963 (N_2963,N_2872,N_2865);
or U2964 (N_2964,N_2921,N_2920);
nor U2965 (N_2965,N_2863,N_2923);
xnor U2966 (N_2966,N_2920,N_2874);
and U2967 (N_2967,N_2898,N_2883);
nand U2968 (N_2968,N_2893,N_2881);
nand U2969 (N_2969,N_2882,N_2915);
and U2970 (N_2970,N_2924,N_2921);
or U2971 (N_2971,N_2911,N_2919);
nor U2972 (N_2972,N_2853,N_2913);
nor U2973 (N_2973,N_2902,N_2883);
nor U2974 (N_2974,N_2871,N_2923);
or U2975 (N_2975,N_2903,N_2858);
nor U2976 (N_2976,N_2898,N_2917);
nand U2977 (N_2977,N_2921,N_2864);
nor U2978 (N_2978,N_2923,N_2899);
or U2979 (N_2979,N_2891,N_2919);
nand U2980 (N_2980,N_2866,N_2857);
nor U2981 (N_2981,N_2872,N_2915);
and U2982 (N_2982,N_2859,N_2904);
or U2983 (N_2983,N_2884,N_2865);
nor U2984 (N_2984,N_2898,N_2894);
nand U2985 (N_2985,N_2864,N_2913);
or U2986 (N_2986,N_2919,N_2913);
or U2987 (N_2987,N_2882,N_2909);
nor U2988 (N_2988,N_2863,N_2852);
nor U2989 (N_2989,N_2873,N_2858);
or U2990 (N_2990,N_2886,N_2920);
nor U2991 (N_2991,N_2891,N_2920);
nor U2992 (N_2992,N_2866,N_2908);
or U2993 (N_2993,N_2922,N_2920);
nor U2994 (N_2994,N_2850,N_2912);
nand U2995 (N_2995,N_2871,N_2877);
nand U2996 (N_2996,N_2899,N_2915);
or U2997 (N_2997,N_2891,N_2892);
or U2998 (N_2998,N_2880,N_2921);
nor U2999 (N_2999,N_2875,N_2924);
and UO_0 (O_0,N_2986,N_2997);
nor UO_1 (O_1,N_2998,N_2983);
nand UO_2 (O_2,N_2966,N_2937);
nor UO_3 (O_3,N_2991,N_2979);
or UO_4 (O_4,N_2933,N_2955);
and UO_5 (O_5,N_2930,N_2947);
or UO_6 (O_6,N_2952,N_2945);
and UO_7 (O_7,N_2973,N_2963);
nor UO_8 (O_8,N_2974,N_2985);
or UO_9 (O_9,N_2988,N_2925);
nand UO_10 (O_10,N_2962,N_2940);
nand UO_11 (O_11,N_2942,N_2982);
and UO_12 (O_12,N_2938,N_2968);
nor UO_13 (O_13,N_2999,N_2992);
nand UO_14 (O_14,N_2990,N_2967);
or UO_15 (O_15,N_2993,N_2995);
and UO_16 (O_16,N_2981,N_2965);
nor UO_17 (O_17,N_2958,N_2987);
or UO_18 (O_18,N_2977,N_2994);
or UO_19 (O_19,N_2957,N_2961);
and UO_20 (O_20,N_2939,N_2941);
or UO_21 (O_21,N_2956,N_2976);
nand UO_22 (O_22,N_2954,N_2934);
and UO_23 (O_23,N_2946,N_2948);
or UO_24 (O_24,N_2926,N_2996);
nand UO_25 (O_25,N_2969,N_2960);
nor UO_26 (O_26,N_2964,N_2950);
and UO_27 (O_27,N_2936,N_2989);
nand UO_28 (O_28,N_2951,N_2928);
xor UO_29 (O_29,N_2949,N_2931);
or UO_30 (O_30,N_2944,N_2935);
and UO_31 (O_31,N_2970,N_2980);
or UO_32 (O_32,N_2972,N_2959);
nor UO_33 (O_33,N_2971,N_2932);
nor UO_34 (O_34,N_2929,N_2953);
and UO_35 (O_35,N_2978,N_2927);
and UO_36 (O_36,N_2975,N_2943);
or UO_37 (O_37,N_2984,N_2953);
nand UO_38 (O_38,N_2962,N_2977);
or UO_39 (O_39,N_2965,N_2931);
and UO_40 (O_40,N_2961,N_2973);
nor UO_41 (O_41,N_2928,N_2999);
or UO_42 (O_42,N_2994,N_2971);
or UO_43 (O_43,N_2942,N_2959);
and UO_44 (O_44,N_2991,N_2925);
nand UO_45 (O_45,N_2935,N_2973);
and UO_46 (O_46,N_2926,N_2942);
or UO_47 (O_47,N_2962,N_2948);
nor UO_48 (O_48,N_2981,N_2958);
nor UO_49 (O_49,N_2952,N_2994);
and UO_50 (O_50,N_2966,N_2968);
and UO_51 (O_51,N_2974,N_2969);
nor UO_52 (O_52,N_2937,N_2925);
nand UO_53 (O_53,N_2925,N_2978);
nor UO_54 (O_54,N_2934,N_2952);
and UO_55 (O_55,N_2932,N_2970);
and UO_56 (O_56,N_2993,N_2936);
and UO_57 (O_57,N_2969,N_2929);
and UO_58 (O_58,N_2931,N_2941);
or UO_59 (O_59,N_2981,N_2968);
or UO_60 (O_60,N_2970,N_2977);
and UO_61 (O_61,N_2962,N_2932);
nand UO_62 (O_62,N_2944,N_2961);
nand UO_63 (O_63,N_2951,N_2958);
nor UO_64 (O_64,N_2964,N_2947);
or UO_65 (O_65,N_2986,N_2925);
nor UO_66 (O_66,N_2960,N_2999);
nand UO_67 (O_67,N_2990,N_2980);
or UO_68 (O_68,N_2961,N_2971);
or UO_69 (O_69,N_2981,N_2982);
or UO_70 (O_70,N_2928,N_2939);
and UO_71 (O_71,N_2932,N_2985);
nor UO_72 (O_72,N_2999,N_2929);
or UO_73 (O_73,N_2991,N_2944);
nor UO_74 (O_74,N_2995,N_2929);
or UO_75 (O_75,N_2926,N_2983);
nor UO_76 (O_76,N_2947,N_2971);
and UO_77 (O_77,N_2980,N_2941);
nor UO_78 (O_78,N_2958,N_2989);
or UO_79 (O_79,N_2966,N_2976);
and UO_80 (O_80,N_2987,N_2947);
or UO_81 (O_81,N_2945,N_2964);
or UO_82 (O_82,N_2979,N_2975);
nor UO_83 (O_83,N_2966,N_2925);
and UO_84 (O_84,N_2974,N_2956);
and UO_85 (O_85,N_2954,N_2983);
nor UO_86 (O_86,N_2934,N_2937);
nor UO_87 (O_87,N_2967,N_2982);
and UO_88 (O_88,N_2983,N_2935);
or UO_89 (O_89,N_2948,N_2925);
or UO_90 (O_90,N_2988,N_2939);
or UO_91 (O_91,N_2968,N_2953);
and UO_92 (O_92,N_2983,N_2936);
nor UO_93 (O_93,N_2947,N_2959);
nand UO_94 (O_94,N_2981,N_2947);
or UO_95 (O_95,N_2926,N_2936);
nand UO_96 (O_96,N_2972,N_2935);
nor UO_97 (O_97,N_2967,N_2963);
or UO_98 (O_98,N_2964,N_2948);
nand UO_99 (O_99,N_2942,N_2990);
or UO_100 (O_100,N_2995,N_2961);
or UO_101 (O_101,N_2968,N_2967);
nand UO_102 (O_102,N_2945,N_2939);
nand UO_103 (O_103,N_2970,N_2979);
nor UO_104 (O_104,N_2972,N_2987);
and UO_105 (O_105,N_2972,N_2976);
xnor UO_106 (O_106,N_2946,N_2944);
and UO_107 (O_107,N_2992,N_2955);
or UO_108 (O_108,N_2978,N_2988);
or UO_109 (O_109,N_2949,N_2986);
and UO_110 (O_110,N_2989,N_2926);
nor UO_111 (O_111,N_2925,N_2994);
nand UO_112 (O_112,N_2965,N_2954);
nor UO_113 (O_113,N_2941,N_2995);
and UO_114 (O_114,N_2961,N_2956);
nor UO_115 (O_115,N_2950,N_2953);
and UO_116 (O_116,N_2988,N_2941);
nor UO_117 (O_117,N_2935,N_2968);
xor UO_118 (O_118,N_2991,N_2977);
nand UO_119 (O_119,N_2932,N_2934);
and UO_120 (O_120,N_2943,N_2994);
and UO_121 (O_121,N_2964,N_2963);
or UO_122 (O_122,N_2976,N_2938);
xnor UO_123 (O_123,N_2993,N_2972);
nand UO_124 (O_124,N_2926,N_2994);
xnor UO_125 (O_125,N_2974,N_2977);
or UO_126 (O_126,N_2975,N_2977);
or UO_127 (O_127,N_2975,N_2953);
and UO_128 (O_128,N_2926,N_2981);
and UO_129 (O_129,N_2930,N_2958);
nand UO_130 (O_130,N_2973,N_2997);
nor UO_131 (O_131,N_2937,N_2979);
nand UO_132 (O_132,N_2972,N_2946);
or UO_133 (O_133,N_2975,N_2994);
or UO_134 (O_134,N_2953,N_2927);
or UO_135 (O_135,N_2969,N_2975);
or UO_136 (O_136,N_2980,N_2961);
and UO_137 (O_137,N_2962,N_2976);
or UO_138 (O_138,N_2986,N_2935);
or UO_139 (O_139,N_2994,N_2929);
or UO_140 (O_140,N_2943,N_2968);
nand UO_141 (O_141,N_2961,N_2952);
xor UO_142 (O_142,N_2942,N_2979);
or UO_143 (O_143,N_2937,N_2990);
or UO_144 (O_144,N_2925,N_2949);
and UO_145 (O_145,N_2938,N_2973);
nor UO_146 (O_146,N_2981,N_2995);
nand UO_147 (O_147,N_2933,N_2969);
xnor UO_148 (O_148,N_2940,N_2933);
and UO_149 (O_149,N_2990,N_2965);
and UO_150 (O_150,N_2939,N_2957);
or UO_151 (O_151,N_2949,N_2943);
and UO_152 (O_152,N_2967,N_2930);
nor UO_153 (O_153,N_2950,N_2961);
nand UO_154 (O_154,N_2947,N_2936);
nand UO_155 (O_155,N_2962,N_2943);
or UO_156 (O_156,N_2938,N_2950);
nand UO_157 (O_157,N_2962,N_2927);
nand UO_158 (O_158,N_2949,N_2948);
nor UO_159 (O_159,N_2993,N_2971);
nor UO_160 (O_160,N_2928,N_2954);
or UO_161 (O_161,N_2979,N_2971);
and UO_162 (O_162,N_2977,N_2986);
nor UO_163 (O_163,N_2988,N_2933);
nand UO_164 (O_164,N_2943,N_2969);
or UO_165 (O_165,N_2948,N_2978);
nor UO_166 (O_166,N_2968,N_2942);
and UO_167 (O_167,N_2951,N_2934);
and UO_168 (O_168,N_2994,N_2935);
and UO_169 (O_169,N_2931,N_2944);
and UO_170 (O_170,N_2984,N_2981);
nand UO_171 (O_171,N_2944,N_2998);
or UO_172 (O_172,N_2968,N_2949);
or UO_173 (O_173,N_2983,N_2933);
xnor UO_174 (O_174,N_2928,N_2986);
and UO_175 (O_175,N_2932,N_2946);
or UO_176 (O_176,N_2997,N_2971);
nor UO_177 (O_177,N_2971,N_2928);
or UO_178 (O_178,N_2984,N_2949);
nor UO_179 (O_179,N_2951,N_2996);
and UO_180 (O_180,N_2995,N_2939);
nand UO_181 (O_181,N_2951,N_2956);
nor UO_182 (O_182,N_2975,N_2932);
nand UO_183 (O_183,N_2970,N_2933);
nor UO_184 (O_184,N_2948,N_2944);
nand UO_185 (O_185,N_2932,N_2928);
nand UO_186 (O_186,N_2999,N_2926);
nor UO_187 (O_187,N_2946,N_2987);
nand UO_188 (O_188,N_2989,N_2953);
nand UO_189 (O_189,N_2981,N_2959);
xor UO_190 (O_190,N_2942,N_2957);
nor UO_191 (O_191,N_2936,N_2938);
nand UO_192 (O_192,N_2937,N_2961);
and UO_193 (O_193,N_2935,N_2939);
nor UO_194 (O_194,N_2952,N_2993);
nor UO_195 (O_195,N_2961,N_2931);
and UO_196 (O_196,N_2954,N_2985);
xnor UO_197 (O_197,N_2942,N_2977);
xor UO_198 (O_198,N_2947,N_2939);
xnor UO_199 (O_199,N_2939,N_2966);
nor UO_200 (O_200,N_2977,N_2953);
nor UO_201 (O_201,N_2928,N_2978);
nand UO_202 (O_202,N_2948,N_2966);
nand UO_203 (O_203,N_2941,N_2932);
or UO_204 (O_204,N_2958,N_2932);
nor UO_205 (O_205,N_2989,N_2948);
nor UO_206 (O_206,N_2928,N_2953);
or UO_207 (O_207,N_2983,N_2979);
or UO_208 (O_208,N_2931,N_2980);
or UO_209 (O_209,N_2958,N_2997);
and UO_210 (O_210,N_2971,N_2953);
and UO_211 (O_211,N_2952,N_2968);
nor UO_212 (O_212,N_2954,N_2940);
nand UO_213 (O_213,N_2999,N_2937);
or UO_214 (O_214,N_2941,N_2991);
nor UO_215 (O_215,N_2930,N_2950);
or UO_216 (O_216,N_2943,N_2948);
or UO_217 (O_217,N_2971,N_2933);
nor UO_218 (O_218,N_2993,N_2939);
or UO_219 (O_219,N_2977,N_2996);
or UO_220 (O_220,N_2984,N_2994);
or UO_221 (O_221,N_2965,N_2982);
nand UO_222 (O_222,N_2992,N_2991);
nor UO_223 (O_223,N_2940,N_2980);
nand UO_224 (O_224,N_2953,N_2962);
and UO_225 (O_225,N_2990,N_2987);
and UO_226 (O_226,N_2975,N_2937);
nand UO_227 (O_227,N_2999,N_2949);
or UO_228 (O_228,N_2941,N_2964);
nor UO_229 (O_229,N_2944,N_2997);
nand UO_230 (O_230,N_2940,N_2974);
nand UO_231 (O_231,N_2951,N_2959);
nand UO_232 (O_232,N_2984,N_2929);
nand UO_233 (O_233,N_2987,N_2963);
nand UO_234 (O_234,N_2942,N_2969);
or UO_235 (O_235,N_2956,N_2944);
nand UO_236 (O_236,N_2972,N_2930);
nor UO_237 (O_237,N_2969,N_2938);
and UO_238 (O_238,N_2972,N_2951);
and UO_239 (O_239,N_2974,N_2995);
or UO_240 (O_240,N_2938,N_2930);
or UO_241 (O_241,N_2979,N_2963);
nand UO_242 (O_242,N_2935,N_2933);
or UO_243 (O_243,N_2948,N_2993);
and UO_244 (O_244,N_2958,N_2995);
or UO_245 (O_245,N_2927,N_2982);
nor UO_246 (O_246,N_2970,N_2935);
nor UO_247 (O_247,N_2968,N_2947);
and UO_248 (O_248,N_2969,N_2993);
nand UO_249 (O_249,N_2998,N_2993);
or UO_250 (O_250,N_2925,N_2927);
and UO_251 (O_251,N_2961,N_2993);
and UO_252 (O_252,N_2967,N_2984);
nor UO_253 (O_253,N_2947,N_2977);
and UO_254 (O_254,N_2998,N_2994);
and UO_255 (O_255,N_2984,N_2952);
nand UO_256 (O_256,N_2945,N_2936);
and UO_257 (O_257,N_2933,N_2944);
and UO_258 (O_258,N_2992,N_2943);
nor UO_259 (O_259,N_2960,N_2996);
and UO_260 (O_260,N_2993,N_2963);
nor UO_261 (O_261,N_2971,N_2974);
and UO_262 (O_262,N_2953,N_2957);
nor UO_263 (O_263,N_2939,N_2933);
nor UO_264 (O_264,N_2999,N_2939);
nor UO_265 (O_265,N_2970,N_2928);
nor UO_266 (O_266,N_2950,N_2968);
and UO_267 (O_267,N_2960,N_2978);
and UO_268 (O_268,N_2996,N_2994);
nor UO_269 (O_269,N_2997,N_2962);
and UO_270 (O_270,N_2968,N_2936);
and UO_271 (O_271,N_2929,N_2970);
nand UO_272 (O_272,N_2927,N_2932);
and UO_273 (O_273,N_2975,N_2976);
nand UO_274 (O_274,N_2925,N_2977);
nand UO_275 (O_275,N_2952,N_2971);
and UO_276 (O_276,N_2984,N_2976);
or UO_277 (O_277,N_2935,N_2993);
nand UO_278 (O_278,N_2977,N_2930);
or UO_279 (O_279,N_2981,N_2974);
nor UO_280 (O_280,N_2980,N_2971);
nor UO_281 (O_281,N_2967,N_2970);
nand UO_282 (O_282,N_2969,N_2947);
and UO_283 (O_283,N_2927,N_2944);
or UO_284 (O_284,N_2925,N_2942);
nor UO_285 (O_285,N_2963,N_2985);
and UO_286 (O_286,N_2956,N_2926);
nand UO_287 (O_287,N_2942,N_2935);
and UO_288 (O_288,N_2971,N_2970);
nand UO_289 (O_289,N_2954,N_2961);
or UO_290 (O_290,N_2945,N_2940);
nand UO_291 (O_291,N_2960,N_2967);
or UO_292 (O_292,N_2934,N_2945);
and UO_293 (O_293,N_2989,N_2998);
xnor UO_294 (O_294,N_2969,N_2999);
or UO_295 (O_295,N_2991,N_2975);
xnor UO_296 (O_296,N_2932,N_2947);
nor UO_297 (O_297,N_2996,N_2998);
or UO_298 (O_298,N_2969,N_2973);
nor UO_299 (O_299,N_2937,N_2971);
nor UO_300 (O_300,N_2956,N_2995);
and UO_301 (O_301,N_2967,N_2965);
and UO_302 (O_302,N_2947,N_2951);
and UO_303 (O_303,N_2943,N_2935);
nor UO_304 (O_304,N_2989,N_2935);
and UO_305 (O_305,N_2968,N_2996);
and UO_306 (O_306,N_2939,N_2989);
nor UO_307 (O_307,N_2949,N_2954);
nand UO_308 (O_308,N_2990,N_2997);
nor UO_309 (O_309,N_2981,N_2938);
nor UO_310 (O_310,N_2958,N_2934);
or UO_311 (O_311,N_2983,N_2942);
or UO_312 (O_312,N_2992,N_2989);
and UO_313 (O_313,N_2981,N_2954);
nor UO_314 (O_314,N_2927,N_2992);
nand UO_315 (O_315,N_2949,N_2995);
nand UO_316 (O_316,N_2952,N_2949);
nand UO_317 (O_317,N_2998,N_2949);
nor UO_318 (O_318,N_2947,N_2978);
nor UO_319 (O_319,N_2989,N_2943);
and UO_320 (O_320,N_2961,N_2939);
nand UO_321 (O_321,N_2991,N_2982);
nor UO_322 (O_322,N_2932,N_2999);
or UO_323 (O_323,N_2973,N_2929);
nor UO_324 (O_324,N_2952,N_2937);
nand UO_325 (O_325,N_2959,N_2950);
nor UO_326 (O_326,N_2925,N_2951);
and UO_327 (O_327,N_2967,N_2949);
nor UO_328 (O_328,N_2976,N_2970);
or UO_329 (O_329,N_2982,N_2937);
nand UO_330 (O_330,N_2970,N_2948);
or UO_331 (O_331,N_2978,N_2985);
and UO_332 (O_332,N_2991,N_2933);
or UO_333 (O_333,N_2945,N_2970);
nand UO_334 (O_334,N_2952,N_2931);
nor UO_335 (O_335,N_2935,N_2952);
or UO_336 (O_336,N_2978,N_2991);
nor UO_337 (O_337,N_2953,N_2958);
nor UO_338 (O_338,N_2932,N_2937);
and UO_339 (O_339,N_2948,N_2955);
or UO_340 (O_340,N_2959,N_2976);
nand UO_341 (O_341,N_2930,N_2975);
or UO_342 (O_342,N_2996,N_2946);
and UO_343 (O_343,N_2956,N_2950);
or UO_344 (O_344,N_2932,N_2979);
nor UO_345 (O_345,N_2968,N_2984);
nor UO_346 (O_346,N_2939,N_2967);
or UO_347 (O_347,N_2997,N_2964);
nand UO_348 (O_348,N_2968,N_2992);
or UO_349 (O_349,N_2977,N_2954);
and UO_350 (O_350,N_2937,N_2950);
nor UO_351 (O_351,N_2982,N_2961);
or UO_352 (O_352,N_2999,N_2971);
nand UO_353 (O_353,N_2953,N_2933);
and UO_354 (O_354,N_2925,N_2934);
and UO_355 (O_355,N_2979,N_2962);
nor UO_356 (O_356,N_2976,N_2937);
nand UO_357 (O_357,N_2925,N_2975);
nor UO_358 (O_358,N_2961,N_2997);
and UO_359 (O_359,N_2951,N_2980);
nor UO_360 (O_360,N_2985,N_2958);
nor UO_361 (O_361,N_2950,N_2963);
and UO_362 (O_362,N_2969,N_2941);
and UO_363 (O_363,N_2954,N_2948);
nor UO_364 (O_364,N_2979,N_2948);
nor UO_365 (O_365,N_2930,N_2962);
nor UO_366 (O_366,N_2980,N_2933);
or UO_367 (O_367,N_2958,N_2931);
nor UO_368 (O_368,N_2935,N_2945);
and UO_369 (O_369,N_2945,N_2983);
nand UO_370 (O_370,N_2927,N_2963);
or UO_371 (O_371,N_2979,N_2926);
nor UO_372 (O_372,N_2991,N_2999);
and UO_373 (O_373,N_2929,N_2927);
nand UO_374 (O_374,N_2984,N_2971);
or UO_375 (O_375,N_2966,N_2956);
and UO_376 (O_376,N_2992,N_2986);
nor UO_377 (O_377,N_2992,N_2959);
nand UO_378 (O_378,N_2952,N_2982);
or UO_379 (O_379,N_2985,N_2980);
or UO_380 (O_380,N_2979,N_2928);
and UO_381 (O_381,N_2981,N_2936);
nor UO_382 (O_382,N_2985,N_2966);
nor UO_383 (O_383,N_2939,N_2959);
or UO_384 (O_384,N_2927,N_2995);
nand UO_385 (O_385,N_2953,N_2985);
or UO_386 (O_386,N_2931,N_2929);
or UO_387 (O_387,N_2959,N_2966);
nand UO_388 (O_388,N_2943,N_2977);
or UO_389 (O_389,N_2977,N_2961);
nand UO_390 (O_390,N_2928,N_2925);
and UO_391 (O_391,N_2929,N_2981);
nand UO_392 (O_392,N_2935,N_2951);
nand UO_393 (O_393,N_2980,N_2942);
nand UO_394 (O_394,N_2945,N_2967);
nand UO_395 (O_395,N_2937,N_2970);
nand UO_396 (O_396,N_2927,N_2958);
or UO_397 (O_397,N_2955,N_2974);
nor UO_398 (O_398,N_2988,N_2981);
nand UO_399 (O_399,N_2940,N_2928);
and UO_400 (O_400,N_2968,N_2970);
or UO_401 (O_401,N_2938,N_2975);
and UO_402 (O_402,N_2960,N_2941);
and UO_403 (O_403,N_2936,N_2997);
nor UO_404 (O_404,N_2948,N_2956);
and UO_405 (O_405,N_2960,N_2934);
nand UO_406 (O_406,N_2960,N_2933);
nand UO_407 (O_407,N_2969,N_2968);
or UO_408 (O_408,N_2983,N_2968);
and UO_409 (O_409,N_2954,N_2970);
or UO_410 (O_410,N_2988,N_2944);
nand UO_411 (O_411,N_2946,N_2962);
nand UO_412 (O_412,N_2951,N_2929);
and UO_413 (O_413,N_2996,N_2997);
nand UO_414 (O_414,N_2973,N_2995);
and UO_415 (O_415,N_2955,N_2975);
nand UO_416 (O_416,N_2985,N_2987);
or UO_417 (O_417,N_2975,N_2949);
or UO_418 (O_418,N_2968,N_2954);
nor UO_419 (O_419,N_2930,N_2987);
or UO_420 (O_420,N_2960,N_2994);
nor UO_421 (O_421,N_2937,N_2962);
nor UO_422 (O_422,N_2949,N_2997);
and UO_423 (O_423,N_2932,N_2952);
and UO_424 (O_424,N_2967,N_2996);
nor UO_425 (O_425,N_2971,N_2969);
nand UO_426 (O_426,N_2952,N_2986);
xor UO_427 (O_427,N_2947,N_2931);
and UO_428 (O_428,N_2977,N_2931);
and UO_429 (O_429,N_2974,N_2970);
and UO_430 (O_430,N_2990,N_2996);
or UO_431 (O_431,N_2926,N_2945);
nand UO_432 (O_432,N_2957,N_2950);
or UO_433 (O_433,N_2977,N_2959);
nand UO_434 (O_434,N_2990,N_2983);
nand UO_435 (O_435,N_2942,N_2939);
xnor UO_436 (O_436,N_2962,N_2973);
and UO_437 (O_437,N_2972,N_2966);
nand UO_438 (O_438,N_2966,N_2928);
nor UO_439 (O_439,N_2965,N_2980);
nand UO_440 (O_440,N_2948,N_2936);
nor UO_441 (O_441,N_2955,N_2980);
and UO_442 (O_442,N_2926,N_2950);
and UO_443 (O_443,N_2983,N_2966);
nor UO_444 (O_444,N_2990,N_2977);
and UO_445 (O_445,N_2995,N_2954);
nand UO_446 (O_446,N_2987,N_2961);
nor UO_447 (O_447,N_2996,N_2983);
nor UO_448 (O_448,N_2941,N_2943);
and UO_449 (O_449,N_2949,N_2944);
or UO_450 (O_450,N_2925,N_2941);
and UO_451 (O_451,N_2954,N_2964);
or UO_452 (O_452,N_2932,N_2977);
nand UO_453 (O_453,N_2961,N_2946);
nor UO_454 (O_454,N_2990,N_2953);
and UO_455 (O_455,N_2940,N_2989);
and UO_456 (O_456,N_2957,N_2980);
and UO_457 (O_457,N_2976,N_2949);
nand UO_458 (O_458,N_2989,N_2933);
or UO_459 (O_459,N_2998,N_2979);
nor UO_460 (O_460,N_2932,N_2936);
or UO_461 (O_461,N_2952,N_2995);
or UO_462 (O_462,N_2994,N_2999);
and UO_463 (O_463,N_2989,N_2956);
and UO_464 (O_464,N_2991,N_2947);
or UO_465 (O_465,N_2969,N_2940);
nor UO_466 (O_466,N_2989,N_2934);
nand UO_467 (O_467,N_2968,N_2944);
nand UO_468 (O_468,N_2986,N_2942);
or UO_469 (O_469,N_2938,N_2998);
nand UO_470 (O_470,N_2933,N_2982);
nor UO_471 (O_471,N_2997,N_2987);
nor UO_472 (O_472,N_2970,N_2952);
nand UO_473 (O_473,N_2934,N_2990);
nand UO_474 (O_474,N_2962,N_2971);
or UO_475 (O_475,N_2987,N_2951);
and UO_476 (O_476,N_2956,N_2960);
nor UO_477 (O_477,N_2984,N_2982);
and UO_478 (O_478,N_2988,N_2984);
nor UO_479 (O_479,N_2980,N_2946);
or UO_480 (O_480,N_2972,N_2944);
nor UO_481 (O_481,N_2997,N_2974);
nand UO_482 (O_482,N_2935,N_2971);
and UO_483 (O_483,N_2986,N_2954);
nand UO_484 (O_484,N_2974,N_2962);
nor UO_485 (O_485,N_2991,N_2931);
nor UO_486 (O_486,N_2937,N_2929);
nor UO_487 (O_487,N_2991,N_2949);
nor UO_488 (O_488,N_2992,N_2941);
nand UO_489 (O_489,N_2974,N_2967);
nand UO_490 (O_490,N_2926,N_2995);
nor UO_491 (O_491,N_2952,N_2962);
or UO_492 (O_492,N_2940,N_2999);
or UO_493 (O_493,N_2940,N_2936);
or UO_494 (O_494,N_2951,N_2938);
and UO_495 (O_495,N_2933,N_2932);
nor UO_496 (O_496,N_2927,N_2936);
or UO_497 (O_497,N_2996,N_2945);
and UO_498 (O_498,N_2929,N_2948);
nor UO_499 (O_499,N_2948,N_2952);
endmodule