module basic_750_5000_1000_25_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_676,In_571);
or U1 (N_1,In_215,In_635);
xor U2 (N_2,In_550,In_5);
and U3 (N_3,In_167,In_4);
or U4 (N_4,In_429,In_278);
nand U5 (N_5,In_648,In_30);
nand U6 (N_6,In_272,In_68);
nand U7 (N_7,In_316,In_664);
nand U8 (N_8,In_131,In_470);
nor U9 (N_9,In_465,In_224);
or U10 (N_10,In_112,In_424);
nor U11 (N_11,In_148,In_62);
nand U12 (N_12,In_232,In_641);
xnor U13 (N_13,In_417,In_307);
and U14 (N_14,In_458,In_715);
xnor U15 (N_15,In_669,In_729);
nand U16 (N_16,In_306,In_168);
and U17 (N_17,In_59,In_710);
xnor U18 (N_18,In_717,In_361);
and U19 (N_19,In_41,In_88);
nor U20 (N_20,In_238,In_241);
xor U21 (N_21,In_13,In_651);
nand U22 (N_22,In_313,In_746);
nand U23 (N_23,In_7,In_244);
nand U24 (N_24,In_478,In_166);
xnor U25 (N_25,In_616,In_356);
and U26 (N_26,In_666,In_340);
xor U27 (N_27,In_357,In_187);
nor U28 (N_28,In_693,In_358);
or U29 (N_29,In_198,In_509);
nand U30 (N_30,In_622,In_559);
and U31 (N_31,In_573,In_591);
or U32 (N_32,In_654,In_44);
nand U33 (N_33,In_450,In_656);
and U34 (N_34,In_599,In_481);
nor U35 (N_35,In_541,In_47);
or U36 (N_36,In_464,In_468);
nor U37 (N_37,In_94,In_703);
and U38 (N_38,In_526,In_264);
nand U39 (N_39,In_551,In_691);
and U40 (N_40,In_512,In_300);
xnor U41 (N_41,In_497,In_701);
nand U42 (N_42,In_297,In_189);
and U43 (N_43,In_386,In_359);
nor U44 (N_44,In_546,In_365);
nor U45 (N_45,In_394,In_197);
nor U46 (N_46,In_443,In_519);
nand U47 (N_47,In_565,In_250);
and U48 (N_48,In_243,In_154);
nand U49 (N_49,In_524,In_677);
xnor U50 (N_50,In_183,In_364);
and U51 (N_51,In_720,In_118);
nor U52 (N_52,In_370,In_706);
nand U53 (N_53,In_130,In_477);
nor U54 (N_54,In_496,In_403);
nand U55 (N_55,In_9,In_523);
and U56 (N_56,In_96,In_678);
or U57 (N_57,In_466,In_220);
or U58 (N_58,In_423,In_704);
xnor U59 (N_59,In_158,In_646);
and U60 (N_60,In_248,In_554);
xor U61 (N_61,In_325,In_687);
nor U62 (N_62,In_146,In_1);
and U63 (N_63,In_291,In_170);
and U64 (N_64,In_536,In_54);
and U65 (N_65,In_375,In_682);
nor U66 (N_66,In_352,In_191);
nor U67 (N_67,In_199,In_14);
nor U68 (N_68,In_90,In_501);
xnor U69 (N_69,In_303,In_111);
and U70 (N_70,In_585,In_226);
or U71 (N_71,In_63,In_418);
and U72 (N_72,In_553,In_110);
nand U73 (N_73,In_169,In_462);
nor U74 (N_74,In_650,In_506);
nor U75 (N_75,In_177,In_201);
nand U76 (N_76,In_208,In_725);
or U77 (N_77,In_567,In_731);
nor U78 (N_78,In_204,In_611);
and U79 (N_79,In_607,In_58);
xnor U80 (N_80,In_415,In_552);
and U81 (N_81,In_507,In_737);
and U82 (N_82,In_285,In_147);
or U83 (N_83,In_51,In_91);
and U84 (N_84,In_564,In_637);
or U85 (N_85,In_320,In_430);
xor U86 (N_86,In_437,In_293);
or U87 (N_87,In_164,In_271);
or U88 (N_88,In_301,In_712);
and U89 (N_89,In_270,In_134);
or U90 (N_90,In_463,In_511);
or U91 (N_91,In_193,In_685);
nand U92 (N_92,In_3,In_378);
or U93 (N_93,In_239,In_86);
xor U94 (N_94,In_499,In_684);
nor U95 (N_95,In_249,In_192);
nor U96 (N_96,In_350,In_342);
nand U97 (N_97,In_435,In_459);
nor U98 (N_98,In_49,In_558);
nor U99 (N_99,In_395,In_494);
nand U100 (N_100,In_389,In_184);
nand U101 (N_101,In_80,In_502);
or U102 (N_102,In_143,In_413);
nor U103 (N_103,In_317,In_655);
nor U104 (N_104,In_12,In_500);
xnor U105 (N_105,In_521,In_730);
nand U106 (N_106,In_602,In_173);
or U107 (N_107,In_438,In_535);
xor U108 (N_108,In_679,In_322);
or U109 (N_109,In_310,In_736);
and U110 (N_110,In_222,In_348);
nor U111 (N_111,In_630,In_686);
xor U112 (N_112,In_613,In_406);
nor U113 (N_113,In_246,In_23);
and U114 (N_114,In_331,In_245);
nor U115 (N_115,In_127,In_747);
and U116 (N_116,In_453,In_488);
or U117 (N_117,In_699,In_416);
and U118 (N_118,In_104,In_163);
and U119 (N_119,In_733,In_83);
nor U120 (N_120,In_537,In_402);
nand U121 (N_121,In_469,In_330);
or U122 (N_122,In_289,In_405);
nand U123 (N_123,In_89,In_434);
and U124 (N_124,In_588,In_381);
and U125 (N_125,In_321,In_475);
and U126 (N_126,In_67,In_76);
xor U127 (N_127,In_16,In_610);
or U128 (N_128,In_516,In_456);
nand U129 (N_129,In_21,In_446);
nand U130 (N_130,In_431,In_547);
and U131 (N_131,In_142,In_741);
nor U132 (N_132,In_263,In_145);
or U133 (N_133,In_85,In_476);
and U134 (N_134,In_606,In_25);
nand U135 (N_135,In_344,In_576);
nand U136 (N_136,In_336,In_619);
nor U137 (N_137,In_714,In_149);
nand U138 (N_138,In_625,In_695);
nor U139 (N_139,In_670,In_689);
or U140 (N_140,In_188,In_633);
nand U141 (N_141,In_195,In_367);
and U142 (N_142,In_11,In_18);
nor U143 (N_143,In_445,In_461);
and U144 (N_144,In_2,In_583);
and U145 (N_145,In_345,In_319);
nor U146 (N_146,In_108,In_745);
nor U147 (N_147,In_572,In_493);
and U148 (N_148,In_99,In_24);
nor U149 (N_149,In_627,In_78);
or U150 (N_150,In_608,In_377);
and U151 (N_151,In_34,In_179);
or U152 (N_152,In_581,In_103);
nor U153 (N_153,In_578,In_335);
nor U154 (N_154,In_411,In_95);
nand U155 (N_155,In_209,In_376);
nand U156 (N_156,In_71,In_570);
nand U157 (N_157,In_19,In_236);
nand U158 (N_158,In_267,In_257);
xor U159 (N_159,In_557,In_174);
nor U160 (N_160,In_160,In_180);
nor U161 (N_161,In_140,In_455);
or U162 (N_162,In_93,In_735);
or U163 (N_163,In_665,In_522);
nor U164 (N_164,In_626,In_290);
and U165 (N_165,In_337,In_29);
nand U166 (N_166,In_657,In_436);
nand U167 (N_167,In_634,In_661);
and U168 (N_168,In_514,In_483);
nand U169 (N_169,In_603,In_694);
xnor U170 (N_170,In_675,In_548);
xnor U171 (N_171,In_360,In_46);
nand U172 (N_172,In_298,In_314);
and U173 (N_173,In_474,In_202);
or U174 (N_174,In_8,In_732);
nor U175 (N_175,In_296,In_543);
nor U176 (N_176,In_50,In_498);
nor U177 (N_177,In_433,In_568);
nor U178 (N_178,In_329,In_440);
or U179 (N_179,In_39,In_491);
and U180 (N_180,In_407,In_273);
or U181 (N_181,In_722,In_719);
and U182 (N_182,In_172,In_17);
or U183 (N_183,In_495,In_141);
nand U184 (N_184,In_667,In_98);
nand U185 (N_185,In_744,In_258);
nand U186 (N_186,In_266,In_74);
and U187 (N_187,In_596,In_35);
or U188 (N_188,In_0,In_346);
and U189 (N_189,In_390,In_72);
nand U190 (N_190,In_409,In_604);
and U191 (N_191,In_587,In_520);
or U192 (N_192,In_617,In_323);
and U193 (N_193,In_471,In_408);
nor U194 (N_194,In_420,In_620);
nand U195 (N_195,In_186,In_31);
xnor U196 (N_196,In_157,In_454);
nand U197 (N_197,In_539,In_55);
nand U198 (N_198,In_117,In_441);
or U199 (N_199,In_339,In_137);
and U200 (N_200,In_57,In_73);
nor U201 (N_201,N_88,N_193);
and U202 (N_202,In_178,In_489);
nor U203 (N_203,N_5,N_98);
nand U204 (N_204,N_40,In_40);
nor U205 (N_205,In_529,In_518);
nor U206 (N_206,In_341,N_126);
nor U207 (N_207,N_138,N_183);
or U208 (N_208,In_309,N_170);
or U209 (N_209,In_6,N_52);
and U210 (N_210,N_157,In_38);
nor U211 (N_211,In_354,N_107);
or U212 (N_212,N_140,In_305);
nor U213 (N_213,In_242,In_702);
nor U214 (N_214,In_205,In_451);
and U215 (N_215,N_28,N_16);
or U216 (N_216,In_439,N_11);
or U217 (N_217,In_254,In_738);
nand U218 (N_218,N_179,N_62);
nand U219 (N_219,In_234,N_131);
and U220 (N_220,In_302,In_334);
nand U221 (N_221,In_697,N_120);
nor U222 (N_222,N_108,In_743);
nor U223 (N_223,In_680,In_632);
nand U224 (N_224,In_614,N_26);
or U225 (N_225,N_111,N_12);
or U226 (N_226,In_176,In_504);
nor U227 (N_227,N_0,In_288);
xnor U228 (N_228,N_154,N_191);
nand U229 (N_229,In_60,In_230);
or U230 (N_230,N_160,N_151);
and U231 (N_231,In_211,In_333);
nand U232 (N_232,In_448,N_90);
or U233 (N_233,In_284,In_82);
nand U234 (N_234,In_582,In_505);
nand U235 (N_235,In_369,In_105);
nor U236 (N_236,N_83,In_229);
nand U237 (N_237,N_48,N_94);
nand U238 (N_238,In_527,N_162);
xor U239 (N_239,N_172,In_414);
nor U240 (N_240,N_185,In_724);
or U241 (N_241,In_276,N_114);
or U242 (N_242,In_629,In_77);
or U243 (N_243,N_6,In_223);
nand U244 (N_244,N_13,In_592);
xor U245 (N_245,N_18,N_164);
nand U246 (N_246,In_315,In_421);
and U247 (N_247,In_533,In_327);
nand U248 (N_248,In_708,In_412);
and U249 (N_249,N_63,In_705);
or U250 (N_250,In_312,N_129);
or U251 (N_251,In_612,N_50);
nor U252 (N_252,N_34,In_318);
and U253 (N_253,In_27,In_396);
or U254 (N_254,N_125,In_388);
or U255 (N_255,In_624,N_144);
xor U256 (N_256,In_525,N_124);
and U257 (N_257,In_721,In_363);
nand U258 (N_258,In_97,In_61);
nor U259 (N_259,In_126,N_77);
xor U260 (N_260,In_472,N_44);
xor U261 (N_261,N_137,In_740);
or U262 (N_262,In_718,N_195);
or U263 (N_263,In_742,In_674);
xnor U264 (N_264,N_155,In_283);
and U265 (N_265,In_566,N_93);
nor U266 (N_266,N_30,In_124);
or U267 (N_267,In_100,In_269);
nand U268 (N_268,N_2,N_78);
nor U269 (N_269,In_253,In_113);
xnor U270 (N_270,N_169,N_141);
and U271 (N_271,In_393,N_103);
or U272 (N_272,N_122,In_136);
and U273 (N_273,In_473,In_398);
nor U274 (N_274,In_125,In_534);
or U275 (N_275,In_683,N_106);
nand U276 (N_276,N_112,N_142);
nor U277 (N_277,N_92,In_700);
xor U278 (N_278,N_69,In_653);
or U279 (N_279,In_139,In_45);
xor U280 (N_280,In_260,In_123);
nand U281 (N_281,In_159,N_113);
or U282 (N_282,In_332,N_187);
and U283 (N_283,In_428,N_59);
nor U284 (N_284,In_452,In_399);
xor U285 (N_285,N_60,In_508);
nor U286 (N_286,In_544,In_643);
or U287 (N_287,In_373,In_70);
or U288 (N_288,In_165,In_503);
and U289 (N_289,In_304,In_748);
nor U290 (N_290,In_419,N_128);
xor U291 (N_291,In_349,In_640);
nand U292 (N_292,In_153,In_383);
xor U293 (N_293,N_81,In_150);
and U294 (N_294,In_15,N_163);
nand U295 (N_295,N_89,In_102);
nor U296 (N_296,In_107,N_117);
or U297 (N_297,N_53,In_101);
nand U298 (N_298,In_133,In_10);
nand U299 (N_299,In_218,In_392);
xor U300 (N_300,N_184,N_25);
nand U301 (N_301,In_295,N_175);
nor U302 (N_302,In_577,In_618);
xnor U303 (N_303,In_181,N_10);
and U304 (N_304,In_580,N_1);
xor U305 (N_305,In_628,In_379);
xor U306 (N_306,In_135,N_84);
nor U307 (N_307,N_105,In_482);
and U308 (N_308,In_644,In_155);
nand U309 (N_309,In_530,In_156);
xnor U310 (N_310,N_97,In_410);
and U311 (N_311,In_696,In_277);
or U312 (N_312,In_513,N_136);
nor U313 (N_313,N_66,N_38);
and U314 (N_314,N_190,In_56);
xor U315 (N_315,In_274,In_353);
xor U316 (N_316,In_515,N_182);
and U317 (N_317,N_71,In_87);
nand U318 (N_318,In_203,In_328);
and U319 (N_319,In_749,In_479);
or U320 (N_320,In_69,In_698);
nand U321 (N_321,In_609,In_540);
or U322 (N_322,In_492,N_165);
nand U323 (N_323,In_151,In_586);
and U324 (N_324,In_185,N_51);
xor U325 (N_325,N_196,N_54);
and U326 (N_326,N_20,N_116);
nand U327 (N_327,In_484,In_563);
and U328 (N_328,N_64,In_510);
and U329 (N_329,N_4,In_621);
nand U330 (N_330,In_681,In_728);
nand U331 (N_331,N_3,N_58);
or U332 (N_332,N_197,In_639);
nand U333 (N_333,N_194,N_14);
xor U334 (N_334,N_41,In_560);
xnor U335 (N_335,In_32,N_121);
nand U336 (N_336,In_196,N_177);
and U337 (N_337,In_216,In_33);
nand U338 (N_338,In_182,N_161);
and U339 (N_339,In_555,In_561);
nor U340 (N_340,In_672,In_132);
or U341 (N_341,In_597,In_457);
nand U342 (N_342,In_391,N_146);
nor U343 (N_343,In_668,In_542);
nand U344 (N_344,N_57,In_268);
or U345 (N_345,In_549,In_144);
nand U346 (N_346,N_159,N_133);
nor U347 (N_347,N_27,N_168);
nand U348 (N_348,In_265,In_449);
and U349 (N_349,N_86,N_167);
xnor U350 (N_350,In_275,In_401);
nand U351 (N_351,In_486,N_186);
and U352 (N_352,In_240,N_152);
nand U353 (N_353,In_707,N_8);
and U354 (N_354,N_82,In_338);
and U355 (N_355,In_114,In_279);
nand U356 (N_356,In_255,In_129);
and U357 (N_357,In_64,In_531);
and U358 (N_358,In_380,N_95);
or U359 (N_359,N_35,N_143);
or U360 (N_360,In_404,N_171);
xor U361 (N_361,In_311,N_127);
or U362 (N_362,N_181,In_42);
or U363 (N_363,In_237,In_711);
nor U364 (N_364,In_119,N_153);
or U365 (N_365,N_99,In_233);
xor U366 (N_366,In_84,In_256);
nor U367 (N_367,In_281,In_623);
nor U368 (N_368,N_115,In_221);
or U369 (N_369,In_92,In_53);
or U370 (N_370,In_447,N_46);
xnor U371 (N_371,N_189,In_723);
or U372 (N_372,In_528,In_326);
nor U373 (N_373,In_190,In_649);
or U374 (N_374,In_36,In_716);
and U375 (N_375,N_32,N_139);
nor U376 (N_376,In_688,N_47);
or U377 (N_377,N_29,In_645);
nor U378 (N_378,In_261,N_73);
and U379 (N_379,In_589,N_72);
nor U380 (N_380,In_467,In_574);
xnor U381 (N_381,In_690,N_100);
and U382 (N_382,In_442,N_36);
or U383 (N_383,In_374,In_287);
or U384 (N_384,In_210,N_118);
nand U385 (N_385,In_262,In_658);
nand U386 (N_386,In_299,N_101);
nor U387 (N_387,In_231,In_372);
and U388 (N_388,In_308,In_175);
xnor U389 (N_389,In_400,In_487);
nor U390 (N_390,In_225,N_33);
nor U391 (N_391,In_385,In_324);
nand U392 (N_392,In_286,In_194);
xor U393 (N_393,In_426,N_166);
xnor U394 (N_394,In_638,In_671);
and U395 (N_395,In_425,In_259);
nor U396 (N_396,N_96,In_663);
and U397 (N_397,In_252,In_590);
and U398 (N_398,N_65,N_199);
or U399 (N_399,In_593,In_26);
nor U400 (N_400,N_320,N_282);
and U401 (N_401,N_273,In_162);
and U402 (N_402,N_298,N_377);
nor U403 (N_403,N_352,In_66);
and U404 (N_404,N_269,N_333);
and U405 (N_405,N_79,N_286);
nand U406 (N_406,N_109,N_200);
and U407 (N_407,In_251,In_20);
or U408 (N_408,N_240,N_319);
or U409 (N_409,N_332,N_102);
nor U410 (N_410,N_267,N_387);
and U411 (N_411,N_307,In_485);
nand U412 (N_412,In_642,N_216);
nand U413 (N_413,N_272,In_605);
and U414 (N_414,In_43,In_79);
or U415 (N_415,N_245,N_209);
nand U416 (N_416,N_328,N_336);
or U417 (N_417,N_388,N_55);
nand U418 (N_418,N_366,In_615);
nor U419 (N_419,In_517,N_359);
and U420 (N_420,In_652,N_304);
nor U421 (N_421,In_206,In_292);
xnor U422 (N_422,In_444,N_394);
and U423 (N_423,In_739,N_296);
nor U424 (N_424,N_250,In_115);
nand U425 (N_425,N_221,N_174);
and U426 (N_426,In_247,In_545);
nand U427 (N_427,N_241,N_277);
nor U428 (N_428,N_293,N_295);
or U429 (N_429,N_331,N_284);
nand U430 (N_430,In_432,In_171);
and U431 (N_431,In_351,N_288);
xor U432 (N_432,In_227,N_373);
nor U433 (N_433,N_61,N_357);
nand U434 (N_434,In_152,In_212);
or U435 (N_435,In_480,N_299);
and U436 (N_436,N_346,N_188);
nor U437 (N_437,N_258,N_268);
nand U438 (N_438,In_662,N_110);
nand U439 (N_439,N_202,N_334);
or U440 (N_440,In_427,N_39);
nor U441 (N_441,N_369,In_384);
xnor U442 (N_442,N_397,N_351);
and U443 (N_443,N_180,N_212);
nor U444 (N_444,N_224,N_342);
nand U445 (N_445,In_347,N_370);
nand U446 (N_446,N_274,In_120);
nand U447 (N_447,N_297,N_104);
nor U448 (N_448,N_70,N_379);
nor U449 (N_449,N_178,In_343);
nand U450 (N_450,In_709,N_231);
nor U451 (N_451,In_600,N_270);
nor U452 (N_452,In_595,N_24);
nand U453 (N_453,N_214,N_263);
or U454 (N_454,In_598,In_575);
nor U455 (N_455,N_257,N_132);
or U456 (N_456,N_21,N_364);
nand U457 (N_457,N_374,N_156);
nand U458 (N_458,N_31,N_244);
and U459 (N_459,N_49,N_375);
nor U460 (N_460,N_391,N_262);
nand U461 (N_461,N_278,N_134);
or U462 (N_462,In_200,N_259);
or U463 (N_463,N_340,N_210);
and U464 (N_464,N_243,N_148);
and U465 (N_465,In_368,In_579);
nand U466 (N_466,N_264,N_42);
nand U467 (N_467,N_343,N_205);
or U468 (N_468,N_313,N_43);
nor U469 (N_469,N_7,In_109);
or U470 (N_470,N_316,N_362);
nand U471 (N_471,N_389,N_367);
xor U472 (N_472,In_673,N_252);
and U473 (N_473,In_569,N_225);
and U474 (N_474,N_337,N_384);
xor U475 (N_475,In_294,N_291);
and U476 (N_476,In_52,N_234);
or U477 (N_477,In_116,N_253);
nor U478 (N_478,N_358,N_37);
or U479 (N_479,N_119,In_460);
or U480 (N_480,N_198,N_15);
or U481 (N_481,In_371,N_354);
nor U482 (N_482,In_355,N_325);
or U483 (N_483,N_398,N_355);
or U484 (N_484,N_87,N_217);
nor U485 (N_485,N_9,In_106);
nor U486 (N_486,N_235,N_238);
nor U487 (N_487,N_67,N_17);
and U488 (N_488,N_266,N_327);
and U489 (N_489,In_538,In_659);
nand U490 (N_490,In_490,N_380);
or U491 (N_491,In_48,In_734);
nand U492 (N_492,N_360,N_91);
nor U493 (N_493,N_356,In_228);
and U494 (N_494,N_306,N_247);
xnor U495 (N_495,N_289,N_361);
and U496 (N_496,N_372,N_345);
nand U497 (N_497,N_329,In_207);
xor U498 (N_498,In_219,In_562);
or U499 (N_499,N_222,N_211);
nor U500 (N_500,N_283,N_149);
or U501 (N_501,In_362,N_204);
nor U502 (N_502,N_368,N_378);
nand U503 (N_503,N_308,In_65);
or U504 (N_504,In_584,N_22);
or U505 (N_505,N_135,N_19);
or U506 (N_506,N_321,N_386);
and U507 (N_507,In_556,In_161);
and U508 (N_508,N_80,N_309);
or U509 (N_509,N_310,N_363);
nand U510 (N_510,In_121,N_323);
xnor U511 (N_511,N_371,N_335);
nor U512 (N_512,N_385,In_217);
or U513 (N_513,N_23,N_287);
and U514 (N_514,In_636,N_349);
or U515 (N_515,In_660,N_381);
or U516 (N_516,N_203,In_601);
and U517 (N_517,In_235,In_81);
nor U518 (N_518,N_207,N_348);
and U519 (N_519,In_422,N_317);
nand U520 (N_520,N_312,N_242);
xnor U521 (N_521,N_292,N_227);
and U522 (N_522,N_256,N_130);
and U523 (N_523,In_727,N_326);
nor U524 (N_524,In_280,N_285);
and U525 (N_525,N_215,N_281);
nor U526 (N_526,In_213,N_383);
nor U527 (N_527,In_532,N_353);
and U528 (N_528,N_395,N_300);
and U529 (N_529,N_338,N_341);
or U530 (N_530,In_726,N_213);
xor U531 (N_531,In_382,N_176);
and U532 (N_532,In_713,N_249);
and U533 (N_533,N_392,In_594);
nand U534 (N_534,N_260,N_158);
nor U535 (N_535,In_214,N_314);
nor U536 (N_536,N_76,N_279);
or U537 (N_537,In_37,N_233);
nand U538 (N_538,N_330,N_344);
xnor U539 (N_539,N_251,N_232);
xor U540 (N_540,N_305,N_315);
nand U541 (N_541,N_301,In_387);
or U542 (N_542,N_201,In_22);
nand U543 (N_543,N_236,N_218);
xnor U544 (N_544,N_280,N_322);
nor U545 (N_545,N_75,N_271);
and U546 (N_546,N_350,N_230);
nand U547 (N_547,N_74,In_397);
xnor U548 (N_548,N_290,N_147);
nand U549 (N_549,N_254,N_220);
or U550 (N_550,N_390,N_246);
and U551 (N_551,In_647,In_138);
or U552 (N_552,N_56,N_339);
nand U553 (N_553,N_85,N_192);
or U554 (N_554,In_282,N_265);
nand U555 (N_555,N_68,In_75);
nor U556 (N_556,N_324,In_631);
and U557 (N_557,N_294,N_239);
and U558 (N_558,N_208,N_318);
nand U559 (N_559,N_276,N_248);
or U560 (N_560,N_311,N_223);
and U561 (N_561,N_219,N_229);
nor U562 (N_562,N_303,N_123);
xnor U563 (N_563,In_692,N_226);
and U564 (N_564,N_302,In_366);
nand U565 (N_565,N_206,In_122);
nor U566 (N_566,N_150,N_275);
xnor U567 (N_567,N_228,N_347);
nor U568 (N_568,N_173,N_382);
or U569 (N_569,In_128,N_45);
nand U570 (N_570,N_255,N_396);
or U571 (N_571,N_145,N_393);
nand U572 (N_572,N_261,N_365);
nand U573 (N_573,N_237,N_376);
or U574 (N_574,In_28,N_399);
and U575 (N_575,N_218,N_23);
nor U576 (N_576,N_355,In_162);
xnor U577 (N_577,In_212,In_20);
or U578 (N_578,N_336,In_713);
and U579 (N_579,N_56,N_24);
nand U580 (N_580,In_647,In_235);
or U581 (N_581,N_148,N_330);
or U582 (N_582,N_399,N_245);
or U583 (N_583,In_713,N_262);
nor U584 (N_584,N_321,N_355);
nand U585 (N_585,N_272,N_370);
nor U586 (N_586,In_162,In_709);
xnor U587 (N_587,N_7,N_247);
and U588 (N_588,N_340,In_662);
nand U589 (N_589,N_265,In_615);
or U590 (N_590,N_281,N_352);
and U591 (N_591,N_279,N_256);
nor U592 (N_592,N_341,N_362);
and U593 (N_593,N_206,N_260);
nor U594 (N_594,In_444,N_206);
and U595 (N_595,N_148,N_247);
and U596 (N_596,In_739,In_594);
xnor U597 (N_597,N_7,In_427);
or U598 (N_598,N_345,N_322);
nand U599 (N_599,N_224,N_180);
nand U600 (N_600,N_492,N_566);
or U601 (N_601,N_483,N_543);
and U602 (N_602,N_565,N_529);
or U603 (N_603,N_490,N_421);
and U604 (N_604,N_514,N_509);
and U605 (N_605,N_540,N_520);
and U606 (N_606,N_451,N_555);
and U607 (N_607,N_536,N_595);
nor U608 (N_608,N_557,N_573);
nor U609 (N_609,N_474,N_587);
xor U610 (N_610,N_570,N_531);
nor U611 (N_611,N_592,N_479);
and U612 (N_612,N_433,N_465);
and U613 (N_613,N_586,N_477);
nand U614 (N_614,N_491,N_581);
nor U615 (N_615,N_548,N_589);
nand U616 (N_616,N_480,N_471);
nand U617 (N_617,N_410,N_445);
or U618 (N_618,N_554,N_537);
and U619 (N_619,N_512,N_559);
nor U620 (N_620,N_460,N_524);
nand U621 (N_621,N_528,N_505);
and U622 (N_622,N_434,N_582);
nand U623 (N_623,N_473,N_584);
nand U624 (N_624,N_456,N_486);
or U625 (N_625,N_447,N_533);
xor U626 (N_626,N_549,N_521);
nor U627 (N_627,N_562,N_443);
nand U628 (N_628,N_527,N_596);
and U629 (N_629,N_412,N_499);
and U630 (N_630,N_428,N_437);
or U631 (N_631,N_576,N_551);
or U632 (N_632,N_523,N_510);
or U633 (N_633,N_449,N_422);
xnor U634 (N_634,N_405,N_487);
and U635 (N_635,N_511,N_401);
and U636 (N_636,N_470,N_475);
xor U637 (N_637,N_454,N_530);
nand U638 (N_638,N_442,N_575);
nand U639 (N_639,N_438,N_419);
nand U640 (N_640,N_518,N_571);
nand U641 (N_641,N_457,N_538);
and U642 (N_642,N_455,N_556);
or U643 (N_643,N_481,N_502);
or U644 (N_644,N_564,N_568);
nand U645 (N_645,N_503,N_439);
xnor U646 (N_646,N_448,N_542);
and U647 (N_647,N_591,N_496);
nor U648 (N_648,N_513,N_574);
nor U649 (N_649,N_462,N_408);
nor U650 (N_650,N_464,N_482);
nand U651 (N_651,N_500,N_497);
and U652 (N_652,N_418,N_588);
and U653 (N_653,N_558,N_569);
nand U654 (N_654,N_466,N_535);
nor U655 (N_655,N_544,N_590);
or U656 (N_656,N_450,N_485);
nand U657 (N_657,N_440,N_446);
and U658 (N_658,N_467,N_534);
or U659 (N_659,N_453,N_539);
or U660 (N_660,N_488,N_472);
xor U661 (N_661,N_572,N_407);
nand U662 (N_662,N_478,N_425);
nor U663 (N_663,N_426,N_522);
and U664 (N_664,N_493,N_409);
nand U665 (N_665,N_414,N_452);
nand U666 (N_666,N_515,N_431);
or U667 (N_667,N_420,N_406);
nor U668 (N_668,N_517,N_411);
nor U669 (N_669,N_532,N_583);
nor U670 (N_670,N_599,N_550);
nor U671 (N_671,N_416,N_494);
nand U672 (N_672,N_506,N_468);
and U673 (N_673,N_444,N_525);
nand U674 (N_674,N_553,N_507);
nor U675 (N_675,N_541,N_516);
nand U676 (N_676,N_546,N_597);
nand U677 (N_677,N_489,N_417);
nand U678 (N_678,N_501,N_578);
nand U679 (N_679,N_561,N_580);
or U680 (N_680,N_560,N_435);
nand U681 (N_681,N_427,N_476);
or U682 (N_682,N_461,N_423);
nand U683 (N_683,N_413,N_436);
and U684 (N_684,N_459,N_547);
nor U685 (N_685,N_484,N_415);
nand U686 (N_686,N_526,N_429);
nand U687 (N_687,N_545,N_577);
nor U688 (N_688,N_504,N_430);
and U689 (N_689,N_403,N_404);
xnor U690 (N_690,N_469,N_441);
nand U691 (N_691,N_508,N_594);
nor U692 (N_692,N_585,N_400);
or U693 (N_693,N_463,N_424);
nor U694 (N_694,N_593,N_579);
xor U695 (N_695,N_552,N_519);
or U696 (N_696,N_498,N_567);
and U697 (N_697,N_495,N_432);
or U698 (N_698,N_402,N_563);
or U699 (N_699,N_458,N_598);
and U700 (N_700,N_427,N_464);
or U701 (N_701,N_554,N_573);
nand U702 (N_702,N_448,N_480);
nand U703 (N_703,N_496,N_526);
nor U704 (N_704,N_479,N_429);
nand U705 (N_705,N_466,N_481);
and U706 (N_706,N_514,N_595);
nor U707 (N_707,N_462,N_516);
nand U708 (N_708,N_532,N_513);
and U709 (N_709,N_409,N_544);
and U710 (N_710,N_511,N_454);
or U711 (N_711,N_540,N_466);
nand U712 (N_712,N_433,N_406);
and U713 (N_713,N_575,N_567);
nor U714 (N_714,N_565,N_566);
or U715 (N_715,N_461,N_598);
nand U716 (N_716,N_522,N_561);
nor U717 (N_717,N_545,N_566);
nand U718 (N_718,N_589,N_405);
nand U719 (N_719,N_516,N_547);
nor U720 (N_720,N_472,N_543);
and U721 (N_721,N_442,N_447);
or U722 (N_722,N_553,N_526);
nand U723 (N_723,N_522,N_498);
nor U724 (N_724,N_427,N_499);
or U725 (N_725,N_535,N_587);
or U726 (N_726,N_541,N_424);
xor U727 (N_727,N_501,N_472);
and U728 (N_728,N_592,N_434);
nor U729 (N_729,N_571,N_433);
xor U730 (N_730,N_519,N_561);
and U731 (N_731,N_512,N_473);
and U732 (N_732,N_547,N_438);
or U733 (N_733,N_470,N_532);
nand U734 (N_734,N_515,N_419);
nor U735 (N_735,N_597,N_403);
and U736 (N_736,N_482,N_489);
or U737 (N_737,N_581,N_549);
nand U738 (N_738,N_490,N_541);
and U739 (N_739,N_446,N_433);
and U740 (N_740,N_451,N_589);
and U741 (N_741,N_445,N_579);
or U742 (N_742,N_510,N_456);
xnor U743 (N_743,N_565,N_592);
nor U744 (N_744,N_588,N_569);
nand U745 (N_745,N_536,N_549);
and U746 (N_746,N_486,N_516);
nand U747 (N_747,N_513,N_565);
or U748 (N_748,N_495,N_408);
and U749 (N_749,N_587,N_457);
or U750 (N_750,N_455,N_451);
nand U751 (N_751,N_570,N_400);
nor U752 (N_752,N_491,N_541);
or U753 (N_753,N_534,N_482);
or U754 (N_754,N_436,N_565);
or U755 (N_755,N_418,N_502);
and U756 (N_756,N_448,N_578);
and U757 (N_757,N_459,N_597);
and U758 (N_758,N_409,N_516);
xor U759 (N_759,N_510,N_552);
nand U760 (N_760,N_455,N_467);
nor U761 (N_761,N_529,N_588);
nand U762 (N_762,N_425,N_567);
or U763 (N_763,N_546,N_518);
nand U764 (N_764,N_483,N_548);
and U765 (N_765,N_549,N_414);
xnor U766 (N_766,N_461,N_452);
and U767 (N_767,N_599,N_401);
and U768 (N_768,N_522,N_558);
and U769 (N_769,N_463,N_492);
and U770 (N_770,N_571,N_484);
or U771 (N_771,N_425,N_406);
and U772 (N_772,N_422,N_465);
or U773 (N_773,N_562,N_524);
or U774 (N_774,N_570,N_431);
and U775 (N_775,N_461,N_589);
or U776 (N_776,N_509,N_567);
and U777 (N_777,N_441,N_553);
or U778 (N_778,N_486,N_457);
and U779 (N_779,N_577,N_443);
and U780 (N_780,N_509,N_555);
nand U781 (N_781,N_400,N_458);
nand U782 (N_782,N_531,N_576);
nand U783 (N_783,N_572,N_439);
nor U784 (N_784,N_556,N_444);
or U785 (N_785,N_455,N_595);
nor U786 (N_786,N_505,N_595);
or U787 (N_787,N_479,N_596);
nor U788 (N_788,N_585,N_466);
or U789 (N_789,N_500,N_432);
nand U790 (N_790,N_522,N_583);
nand U791 (N_791,N_403,N_493);
or U792 (N_792,N_559,N_474);
and U793 (N_793,N_475,N_593);
nor U794 (N_794,N_521,N_555);
nand U795 (N_795,N_550,N_450);
xnor U796 (N_796,N_578,N_446);
or U797 (N_797,N_454,N_467);
nand U798 (N_798,N_490,N_572);
or U799 (N_799,N_461,N_446);
and U800 (N_800,N_629,N_790);
nor U801 (N_801,N_788,N_634);
xnor U802 (N_802,N_749,N_721);
or U803 (N_803,N_650,N_679);
and U804 (N_804,N_697,N_600);
or U805 (N_805,N_663,N_777);
nand U806 (N_806,N_793,N_762);
nand U807 (N_807,N_739,N_646);
and U808 (N_808,N_640,N_628);
xnor U809 (N_809,N_602,N_607);
nand U810 (N_810,N_604,N_741);
nand U811 (N_811,N_661,N_794);
nor U812 (N_812,N_619,N_700);
nand U813 (N_813,N_752,N_738);
nor U814 (N_814,N_753,N_680);
or U815 (N_815,N_651,N_649);
and U816 (N_816,N_787,N_674);
nor U817 (N_817,N_765,N_667);
nor U818 (N_818,N_638,N_760);
nand U819 (N_819,N_695,N_785);
or U820 (N_820,N_745,N_726);
nand U821 (N_821,N_611,N_740);
or U822 (N_822,N_672,N_789);
nor U823 (N_823,N_690,N_660);
nand U824 (N_824,N_758,N_761);
and U825 (N_825,N_678,N_795);
nor U826 (N_826,N_747,N_691);
nand U827 (N_827,N_731,N_792);
nand U828 (N_828,N_624,N_734);
and U829 (N_829,N_706,N_673);
nor U830 (N_830,N_653,N_621);
or U831 (N_831,N_648,N_767);
and U832 (N_832,N_799,N_684);
or U833 (N_833,N_720,N_724);
and U834 (N_834,N_776,N_623);
nor U835 (N_835,N_756,N_633);
and U836 (N_836,N_616,N_727);
or U837 (N_837,N_773,N_698);
or U838 (N_838,N_750,N_748);
nand U839 (N_839,N_718,N_658);
nor U840 (N_840,N_774,N_682);
or U841 (N_841,N_780,N_620);
nor U842 (N_842,N_654,N_635);
nor U843 (N_843,N_713,N_707);
and U844 (N_844,N_610,N_668);
nand U845 (N_845,N_641,N_693);
nor U846 (N_846,N_603,N_732);
nand U847 (N_847,N_609,N_755);
nor U848 (N_848,N_683,N_671);
nor U849 (N_849,N_696,N_716);
or U850 (N_850,N_772,N_681);
nor U851 (N_851,N_730,N_647);
and U852 (N_852,N_659,N_770);
nor U853 (N_853,N_708,N_639);
nand U854 (N_854,N_786,N_798);
nor U855 (N_855,N_686,N_797);
or U856 (N_856,N_665,N_782);
and U857 (N_857,N_630,N_605);
and U858 (N_858,N_735,N_746);
nor U859 (N_859,N_759,N_645);
or U860 (N_860,N_796,N_615);
xor U861 (N_861,N_625,N_687);
and U862 (N_862,N_652,N_717);
or U863 (N_863,N_675,N_703);
and U864 (N_864,N_757,N_676);
and U865 (N_865,N_781,N_608);
nand U866 (N_866,N_606,N_689);
nand U867 (N_867,N_617,N_666);
or U868 (N_868,N_733,N_725);
and U869 (N_869,N_669,N_688);
nand U870 (N_870,N_775,N_715);
and U871 (N_871,N_737,N_627);
nand U872 (N_872,N_601,N_723);
and U873 (N_873,N_743,N_614);
and U874 (N_874,N_685,N_771);
nand U875 (N_875,N_764,N_712);
nand U876 (N_876,N_692,N_714);
and U877 (N_877,N_636,N_736);
nor U878 (N_878,N_766,N_783);
nor U879 (N_879,N_632,N_694);
nand U880 (N_880,N_699,N_618);
nor U881 (N_881,N_779,N_631);
nand U882 (N_882,N_670,N_742);
nor U883 (N_883,N_763,N_709);
or U884 (N_884,N_768,N_642);
nor U885 (N_885,N_719,N_644);
nor U886 (N_886,N_677,N_729);
nor U887 (N_887,N_613,N_751);
or U888 (N_888,N_702,N_769);
and U889 (N_889,N_722,N_791);
nand U890 (N_890,N_612,N_656);
nand U891 (N_891,N_710,N_622);
and U892 (N_892,N_705,N_626);
or U893 (N_893,N_637,N_701);
nor U894 (N_894,N_744,N_664);
nand U895 (N_895,N_662,N_778);
or U896 (N_896,N_655,N_704);
or U897 (N_897,N_728,N_784);
or U898 (N_898,N_754,N_711);
nor U899 (N_899,N_657,N_643);
or U900 (N_900,N_717,N_751);
or U901 (N_901,N_722,N_756);
nand U902 (N_902,N_611,N_644);
xor U903 (N_903,N_698,N_787);
or U904 (N_904,N_761,N_753);
nor U905 (N_905,N_654,N_734);
nand U906 (N_906,N_630,N_796);
or U907 (N_907,N_760,N_601);
or U908 (N_908,N_605,N_736);
nand U909 (N_909,N_632,N_768);
or U910 (N_910,N_647,N_609);
and U911 (N_911,N_618,N_622);
or U912 (N_912,N_759,N_660);
and U913 (N_913,N_606,N_640);
or U914 (N_914,N_693,N_654);
nor U915 (N_915,N_645,N_627);
and U916 (N_916,N_621,N_648);
and U917 (N_917,N_769,N_771);
and U918 (N_918,N_652,N_687);
nor U919 (N_919,N_600,N_625);
nand U920 (N_920,N_670,N_663);
or U921 (N_921,N_785,N_698);
and U922 (N_922,N_617,N_729);
and U923 (N_923,N_756,N_753);
or U924 (N_924,N_639,N_684);
nand U925 (N_925,N_621,N_600);
xor U926 (N_926,N_673,N_781);
nor U927 (N_927,N_780,N_651);
xnor U928 (N_928,N_620,N_749);
nand U929 (N_929,N_767,N_718);
nor U930 (N_930,N_741,N_726);
nor U931 (N_931,N_642,N_783);
or U932 (N_932,N_705,N_728);
or U933 (N_933,N_751,N_769);
nand U934 (N_934,N_682,N_607);
or U935 (N_935,N_764,N_740);
nand U936 (N_936,N_753,N_769);
and U937 (N_937,N_618,N_644);
xor U938 (N_938,N_630,N_774);
nor U939 (N_939,N_679,N_760);
and U940 (N_940,N_682,N_678);
or U941 (N_941,N_791,N_710);
nor U942 (N_942,N_724,N_746);
nand U943 (N_943,N_762,N_771);
or U944 (N_944,N_771,N_759);
nor U945 (N_945,N_732,N_651);
nor U946 (N_946,N_744,N_740);
xor U947 (N_947,N_740,N_674);
nand U948 (N_948,N_645,N_621);
nor U949 (N_949,N_763,N_735);
and U950 (N_950,N_647,N_706);
and U951 (N_951,N_732,N_783);
nor U952 (N_952,N_645,N_669);
and U953 (N_953,N_741,N_668);
xnor U954 (N_954,N_733,N_710);
nor U955 (N_955,N_696,N_724);
nor U956 (N_956,N_658,N_601);
nand U957 (N_957,N_660,N_641);
nor U958 (N_958,N_771,N_647);
nor U959 (N_959,N_789,N_669);
or U960 (N_960,N_730,N_791);
nor U961 (N_961,N_607,N_611);
or U962 (N_962,N_717,N_631);
nor U963 (N_963,N_741,N_772);
nor U964 (N_964,N_694,N_656);
nor U965 (N_965,N_713,N_617);
and U966 (N_966,N_644,N_676);
or U967 (N_967,N_700,N_784);
nand U968 (N_968,N_644,N_774);
nand U969 (N_969,N_756,N_698);
nor U970 (N_970,N_656,N_710);
nand U971 (N_971,N_745,N_695);
or U972 (N_972,N_686,N_643);
or U973 (N_973,N_652,N_738);
and U974 (N_974,N_615,N_751);
nor U975 (N_975,N_698,N_701);
nand U976 (N_976,N_750,N_754);
and U977 (N_977,N_611,N_639);
nor U978 (N_978,N_633,N_693);
nand U979 (N_979,N_784,N_720);
nand U980 (N_980,N_726,N_606);
or U981 (N_981,N_700,N_748);
or U982 (N_982,N_775,N_661);
or U983 (N_983,N_639,N_648);
or U984 (N_984,N_698,N_681);
nand U985 (N_985,N_631,N_630);
nor U986 (N_986,N_687,N_736);
or U987 (N_987,N_783,N_717);
xor U988 (N_988,N_775,N_631);
nor U989 (N_989,N_666,N_656);
nand U990 (N_990,N_627,N_753);
xor U991 (N_991,N_701,N_622);
nand U992 (N_992,N_683,N_789);
nand U993 (N_993,N_613,N_677);
and U994 (N_994,N_668,N_648);
nor U995 (N_995,N_706,N_642);
nand U996 (N_996,N_738,N_796);
and U997 (N_997,N_676,N_765);
xor U998 (N_998,N_686,N_710);
nand U999 (N_999,N_745,N_676);
and U1000 (N_1000,N_986,N_869);
nor U1001 (N_1001,N_962,N_877);
nor U1002 (N_1002,N_904,N_938);
or U1003 (N_1003,N_893,N_910);
xor U1004 (N_1004,N_996,N_822);
nand U1005 (N_1005,N_914,N_955);
nor U1006 (N_1006,N_879,N_800);
and U1007 (N_1007,N_944,N_876);
nor U1008 (N_1008,N_923,N_857);
nand U1009 (N_1009,N_834,N_946);
nor U1010 (N_1010,N_858,N_999);
and U1011 (N_1011,N_807,N_801);
xnor U1012 (N_1012,N_990,N_929);
and U1013 (N_1013,N_838,N_920);
nor U1014 (N_1014,N_868,N_878);
nand U1015 (N_1015,N_915,N_837);
nor U1016 (N_1016,N_802,N_865);
nor U1017 (N_1017,N_917,N_899);
and U1018 (N_1018,N_926,N_847);
nand U1019 (N_1019,N_934,N_855);
and U1020 (N_1020,N_909,N_974);
nor U1021 (N_1021,N_989,N_921);
and U1022 (N_1022,N_911,N_981);
nand U1023 (N_1023,N_805,N_852);
or U1024 (N_1024,N_866,N_939);
nor U1025 (N_1025,N_845,N_827);
or U1026 (N_1026,N_988,N_951);
xnor U1027 (N_1027,N_928,N_843);
or U1028 (N_1028,N_810,N_985);
xor U1029 (N_1029,N_896,N_861);
and U1030 (N_1030,N_961,N_821);
and U1031 (N_1031,N_913,N_916);
or U1032 (N_1032,N_970,N_823);
and U1033 (N_1033,N_842,N_975);
xor U1034 (N_1034,N_969,N_846);
nor U1035 (N_1035,N_856,N_979);
nand U1036 (N_1036,N_952,N_824);
xor U1037 (N_1037,N_832,N_968);
and U1038 (N_1038,N_967,N_884);
nand U1039 (N_1039,N_947,N_991);
or U1040 (N_1040,N_987,N_978);
and U1041 (N_1041,N_849,N_883);
and U1042 (N_1042,N_966,N_922);
or U1043 (N_1043,N_851,N_965);
or U1044 (N_1044,N_871,N_853);
or U1045 (N_1045,N_958,N_905);
nand U1046 (N_1046,N_907,N_841);
nor U1047 (N_1047,N_873,N_903);
nand U1048 (N_1048,N_806,N_937);
xnor U1049 (N_1049,N_924,N_976);
and U1050 (N_1050,N_840,N_954);
nand U1051 (N_1051,N_820,N_956);
nand U1052 (N_1052,N_992,N_862);
and U1053 (N_1053,N_918,N_828);
or U1054 (N_1054,N_943,N_892);
or U1055 (N_1055,N_948,N_894);
xor U1056 (N_1056,N_900,N_912);
nor U1057 (N_1057,N_908,N_812);
and U1058 (N_1058,N_964,N_864);
nand U1059 (N_1059,N_835,N_995);
or U1060 (N_1060,N_818,N_932);
and U1061 (N_1061,N_872,N_859);
nor U1062 (N_1062,N_931,N_942);
nand U1063 (N_1063,N_870,N_880);
nor U1064 (N_1064,N_973,N_998);
nor U1065 (N_1065,N_933,N_949);
and U1066 (N_1066,N_960,N_889);
nand U1067 (N_1067,N_839,N_953);
or U1068 (N_1068,N_919,N_885);
nand U1069 (N_1069,N_829,N_980);
or U1070 (N_1070,N_814,N_819);
and U1071 (N_1071,N_863,N_850);
nor U1072 (N_1072,N_936,N_815);
nand U1073 (N_1073,N_887,N_886);
nor U1074 (N_1074,N_809,N_895);
and U1075 (N_1075,N_959,N_994);
nand U1076 (N_1076,N_888,N_930);
nand U1077 (N_1077,N_890,N_804);
or U1078 (N_1078,N_963,N_831);
nand U1079 (N_1079,N_816,N_830);
nor U1080 (N_1080,N_882,N_902);
xnor U1081 (N_1081,N_950,N_941);
nor U1082 (N_1082,N_935,N_833);
nor U1083 (N_1083,N_867,N_925);
and U1084 (N_1084,N_997,N_875);
or U1085 (N_1085,N_844,N_874);
nand U1086 (N_1086,N_891,N_993);
or U1087 (N_1087,N_897,N_813);
nor U1088 (N_1088,N_881,N_898);
or U1089 (N_1089,N_836,N_971);
or U1090 (N_1090,N_972,N_906);
nor U1091 (N_1091,N_826,N_803);
or U1092 (N_1092,N_854,N_945);
or U1093 (N_1093,N_811,N_860);
and U1094 (N_1094,N_982,N_977);
nand U1095 (N_1095,N_848,N_984);
nor U1096 (N_1096,N_901,N_983);
or U1097 (N_1097,N_817,N_927);
nor U1098 (N_1098,N_957,N_940);
xnor U1099 (N_1099,N_808,N_825);
nor U1100 (N_1100,N_975,N_988);
and U1101 (N_1101,N_940,N_999);
and U1102 (N_1102,N_971,N_993);
and U1103 (N_1103,N_898,N_821);
nor U1104 (N_1104,N_808,N_899);
and U1105 (N_1105,N_857,N_910);
nand U1106 (N_1106,N_927,N_877);
and U1107 (N_1107,N_896,N_887);
nand U1108 (N_1108,N_975,N_889);
nand U1109 (N_1109,N_893,N_955);
xor U1110 (N_1110,N_922,N_802);
or U1111 (N_1111,N_938,N_942);
nor U1112 (N_1112,N_865,N_822);
nand U1113 (N_1113,N_999,N_883);
or U1114 (N_1114,N_915,N_806);
nand U1115 (N_1115,N_822,N_831);
or U1116 (N_1116,N_928,N_938);
nand U1117 (N_1117,N_845,N_941);
xor U1118 (N_1118,N_815,N_953);
or U1119 (N_1119,N_991,N_851);
nor U1120 (N_1120,N_834,N_925);
nor U1121 (N_1121,N_827,N_994);
or U1122 (N_1122,N_959,N_903);
and U1123 (N_1123,N_946,N_902);
and U1124 (N_1124,N_889,N_821);
xnor U1125 (N_1125,N_885,N_991);
nand U1126 (N_1126,N_961,N_886);
nor U1127 (N_1127,N_837,N_979);
or U1128 (N_1128,N_959,N_925);
nor U1129 (N_1129,N_841,N_878);
or U1130 (N_1130,N_801,N_901);
nand U1131 (N_1131,N_861,N_962);
nor U1132 (N_1132,N_877,N_800);
nor U1133 (N_1133,N_997,N_962);
or U1134 (N_1134,N_991,N_842);
nor U1135 (N_1135,N_947,N_896);
nand U1136 (N_1136,N_916,N_926);
nor U1137 (N_1137,N_965,N_949);
nand U1138 (N_1138,N_865,N_956);
nor U1139 (N_1139,N_840,N_962);
xnor U1140 (N_1140,N_913,N_970);
nand U1141 (N_1141,N_916,N_839);
nor U1142 (N_1142,N_917,N_827);
nor U1143 (N_1143,N_842,N_962);
and U1144 (N_1144,N_863,N_985);
nor U1145 (N_1145,N_827,N_975);
or U1146 (N_1146,N_885,N_990);
or U1147 (N_1147,N_846,N_891);
nor U1148 (N_1148,N_869,N_924);
nor U1149 (N_1149,N_937,N_963);
and U1150 (N_1150,N_945,N_918);
and U1151 (N_1151,N_934,N_880);
nand U1152 (N_1152,N_882,N_949);
nand U1153 (N_1153,N_846,N_868);
or U1154 (N_1154,N_960,N_983);
or U1155 (N_1155,N_968,N_871);
nor U1156 (N_1156,N_930,N_887);
or U1157 (N_1157,N_960,N_973);
nor U1158 (N_1158,N_913,N_902);
and U1159 (N_1159,N_988,N_962);
nand U1160 (N_1160,N_827,N_800);
or U1161 (N_1161,N_914,N_874);
nand U1162 (N_1162,N_832,N_837);
or U1163 (N_1163,N_992,N_965);
nand U1164 (N_1164,N_988,N_999);
or U1165 (N_1165,N_937,N_830);
nand U1166 (N_1166,N_978,N_813);
nand U1167 (N_1167,N_806,N_825);
nand U1168 (N_1168,N_918,N_930);
nor U1169 (N_1169,N_811,N_931);
or U1170 (N_1170,N_816,N_896);
nand U1171 (N_1171,N_830,N_916);
nor U1172 (N_1172,N_912,N_965);
and U1173 (N_1173,N_940,N_873);
nand U1174 (N_1174,N_885,N_889);
nand U1175 (N_1175,N_997,N_955);
and U1176 (N_1176,N_808,N_835);
and U1177 (N_1177,N_994,N_848);
nand U1178 (N_1178,N_903,N_823);
nand U1179 (N_1179,N_845,N_948);
nor U1180 (N_1180,N_850,N_931);
or U1181 (N_1181,N_858,N_855);
nand U1182 (N_1182,N_874,N_809);
nand U1183 (N_1183,N_912,N_931);
and U1184 (N_1184,N_846,N_895);
nand U1185 (N_1185,N_957,N_894);
nor U1186 (N_1186,N_903,N_836);
nor U1187 (N_1187,N_986,N_823);
xnor U1188 (N_1188,N_861,N_869);
and U1189 (N_1189,N_821,N_920);
nand U1190 (N_1190,N_812,N_972);
nand U1191 (N_1191,N_936,N_939);
nand U1192 (N_1192,N_903,N_868);
and U1193 (N_1193,N_991,N_987);
nand U1194 (N_1194,N_871,N_860);
or U1195 (N_1195,N_801,N_848);
nor U1196 (N_1196,N_862,N_934);
nor U1197 (N_1197,N_857,N_845);
nor U1198 (N_1198,N_936,N_949);
or U1199 (N_1199,N_992,N_807);
or U1200 (N_1200,N_1001,N_1186);
nor U1201 (N_1201,N_1041,N_1088);
nand U1202 (N_1202,N_1010,N_1195);
xnor U1203 (N_1203,N_1199,N_1026);
or U1204 (N_1204,N_1087,N_1050);
nor U1205 (N_1205,N_1078,N_1058);
and U1206 (N_1206,N_1125,N_1081);
xor U1207 (N_1207,N_1163,N_1039);
and U1208 (N_1208,N_1159,N_1169);
nor U1209 (N_1209,N_1123,N_1036);
nand U1210 (N_1210,N_1177,N_1133);
or U1211 (N_1211,N_1022,N_1120);
and U1212 (N_1212,N_1170,N_1023);
or U1213 (N_1213,N_1111,N_1134);
and U1214 (N_1214,N_1063,N_1082);
nand U1215 (N_1215,N_1046,N_1066);
nand U1216 (N_1216,N_1126,N_1034);
nand U1217 (N_1217,N_1052,N_1196);
or U1218 (N_1218,N_1083,N_1065);
and U1219 (N_1219,N_1187,N_1074);
xnor U1220 (N_1220,N_1136,N_1172);
nand U1221 (N_1221,N_1119,N_1184);
or U1222 (N_1222,N_1140,N_1130);
or U1223 (N_1223,N_1104,N_1102);
nand U1224 (N_1224,N_1093,N_1038);
nand U1225 (N_1225,N_1020,N_1072);
and U1226 (N_1226,N_1189,N_1002);
nand U1227 (N_1227,N_1100,N_1122);
nand U1228 (N_1228,N_1030,N_1137);
or U1229 (N_1229,N_1028,N_1037);
and U1230 (N_1230,N_1105,N_1094);
and U1231 (N_1231,N_1147,N_1181);
or U1232 (N_1232,N_1194,N_1054);
or U1233 (N_1233,N_1179,N_1060);
or U1234 (N_1234,N_1173,N_1185);
or U1235 (N_1235,N_1043,N_1131);
nand U1236 (N_1236,N_1151,N_1166);
nor U1237 (N_1237,N_1068,N_1071);
and U1238 (N_1238,N_1069,N_1005);
and U1239 (N_1239,N_1096,N_1162);
or U1240 (N_1240,N_1141,N_1183);
nand U1241 (N_1241,N_1009,N_1124);
nor U1242 (N_1242,N_1138,N_1029);
or U1243 (N_1243,N_1011,N_1110);
or U1244 (N_1244,N_1097,N_1175);
or U1245 (N_1245,N_1193,N_1064);
xnor U1246 (N_1246,N_1116,N_1171);
or U1247 (N_1247,N_1145,N_1040);
or U1248 (N_1248,N_1129,N_1047);
and U1249 (N_1249,N_1000,N_1101);
and U1250 (N_1250,N_1032,N_1154);
nor U1251 (N_1251,N_1118,N_1008);
xnor U1252 (N_1252,N_1062,N_1055);
xnor U1253 (N_1253,N_1053,N_1167);
and U1254 (N_1254,N_1027,N_1085);
nor U1255 (N_1255,N_1025,N_1033);
and U1256 (N_1256,N_1076,N_1049);
and U1257 (N_1257,N_1044,N_1017);
nand U1258 (N_1258,N_1059,N_1098);
or U1259 (N_1259,N_1095,N_1198);
or U1260 (N_1260,N_1155,N_1135);
or U1261 (N_1261,N_1070,N_1168);
nand U1262 (N_1262,N_1178,N_1152);
and U1263 (N_1263,N_1157,N_1143);
or U1264 (N_1264,N_1042,N_1018);
or U1265 (N_1265,N_1114,N_1158);
or U1266 (N_1266,N_1190,N_1015);
xnor U1267 (N_1267,N_1014,N_1075);
or U1268 (N_1268,N_1144,N_1089);
nand U1269 (N_1269,N_1021,N_1176);
nor U1270 (N_1270,N_1139,N_1192);
and U1271 (N_1271,N_1079,N_1128);
nand U1272 (N_1272,N_1077,N_1103);
xnor U1273 (N_1273,N_1045,N_1091);
and U1274 (N_1274,N_1117,N_1153);
xor U1275 (N_1275,N_1121,N_1084);
xnor U1276 (N_1276,N_1056,N_1188);
nand U1277 (N_1277,N_1197,N_1156);
nand U1278 (N_1278,N_1019,N_1003);
nand U1279 (N_1279,N_1149,N_1007);
and U1280 (N_1280,N_1092,N_1006);
or U1281 (N_1281,N_1182,N_1067);
nor U1282 (N_1282,N_1024,N_1180);
xor U1283 (N_1283,N_1150,N_1012);
nand U1284 (N_1284,N_1061,N_1161);
xor U1285 (N_1285,N_1112,N_1016);
and U1286 (N_1286,N_1115,N_1107);
or U1287 (N_1287,N_1127,N_1004);
xnor U1288 (N_1288,N_1132,N_1160);
nor U1289 (N_1289,N_1109,N_1148);
and U1290 (N_1290,N_1099,N_1165);
nor U1291 (N_1291,N_1191,N_1106);
nor U1292 (N_1292,N_1080,N_1090);
and U1293 (N_1293,N_1164,N_1142);
and U1294 (N_1294,N_1035,N_1174);
nand U1295 (N_1295,N_1073,N_1031);
and U1296 (N_1296,N_1108,N_1051);
and U1297 (N_1297,N_1113,N_1086);
nand U1298 (N_1298,N_1057,N_1048);
nor U1299 (N_1299,N_1013,N_1146);
and U1300 (N_1300,N_1125,N_1176);
xnor U1301 (N_1301,N_1175,N_1158);
xor U1302 (N_1302,N_1090,N_1052);
and U1303 (N_1303,N_1166,N_1161);
nor U1304 (N_1304,N_1184,N_1071);
xor U1305 (N_1305,N_1013,N_1136);
nand U1306 (N_1306,N_1158,N_1124);
or U1307 (N_1307,N_1136,N_1129);
and U1308 (N_1308,N_1008,N_1158);
or U1309 (N_1309,N_1089,N_1083);
nand U1310 (N_1310,N_1006,N_1098);
nand U1311 (N_1311,N_1092,N_1015);
nand U1312 (N_1312,N_1127,N_1052);
and U1313 (N_1313,N_1123,N_1090);
xor U1314 (N_1314,N_1090,N_1021);
and U1315 (N_1315,N_1138,N_1003);
xnor U1316 (N_1316,N_1050,N_1047);
nand U1317 (N_1317,N_1026,N_1054);
and U1318 (N_1318,N_1066,N_1089);
nor U1319 (N_1319,N_1120,N_1197);
nor U1320 (N_1320,N_1020,N_1077);
nor U1321 (N_1321,N_1086,N_1081);
and U1322 (N_1322,N_1038,N_1112);
xnor U1323 (N_1323,N_1078,N_1009);
and U1324 (N_1324,N_1184,N_1151);
xnor U1325 (N_1325,N_1142,N_1102);
nor U1326 (N_1326,N_1146,N_1020);
and U1327 (N_1327,N_1126,N_1131);
and U1328 (N_1328,N_1161,N_1125);
nand U1329 (N_1329,N_1056,N_1059);
or U1330 (N_1330,N_1136,N_1143);
or U1331 (N_1331,N_1113,N_1127);
nand U1332 (N_1332,N_1022,N_1072);
nand U1333 (N_1333,N_1017,N_1184);
and U1334 (N_1334,N_1054,N_1136);
nor U1335 (N_1335,N_1182,N_1063);
or U1336 (N_1336,N_1171,N_1127);
nand U1337 (N_1337,N_1053,N_1137);
nor U1338 (N_1338,N_1107,N_1166);
or U1339 (N_1339,N_1139,N_1170);
nor U1340 (N_1340,N_1016,N_1157);
and U1341 (N_1341,N_1006,N_1129);
nand U1342 (N_1342,N_1129,N_1037);
xor U1343 (N_1343,N_1190,N_1103);
and U1344 (N_1344,N_1043,N_1159);
nor U1345 (N_1345,N_1017,N_1013);
or U1346 (N_1346,N_1085,N_1099);
nand U1347 (N_1347,N_1167,N_1159);
or U1348 (N_1348,N_1016,N_1038);
nand U1349 (N_1349,N_1073,N_1196);
or U1350 (N_1350,N_1121,N_1040);
xnor U1351 (N_1351,N_1184,N_1016);
nor U1352 (N_1352,N_1042,N_1170);
and U1353 (N_1353,N_1070,N_1182);
or U1354 (N_1354,N_1038,N_1074);
and U1355 (N_1355,N_1180,N_1008);
nand U1356 (N_1356,N_1154,N_1143);
and U1357 (N_1357,N_1091,N_1129);
or U1358 (N_1358,N_1127,N_1169);
or U1359 (N_1359,N_1033,N_1030);
nand U1360 (N_1360,N_1107,N_1012);
nand U1361 (N_1361,N_1115,N_1189);
nor U1362 (N_1362,N_1112,N_1155);
xor U1363 (N_1363,N_1173,N_1121);
or U1364 (N_1364,N_1029,N_1051);
or U1365 (N_1365,N_1052,N_1179);
or U1366 (N_1366,N_1115,N_1166);
or U1367 (N_1367,N_1002,N_1016);
nand U1368 (N_1368,N_1012,N_1092);
nor U1369 (N_1369,N_1155,N_1160);
or U1370 (N_1370,N_1079,N_1163);
nor U1371 (N_1371,N_1150,N_1168);
nor U1372 (N_1372,N_1090,N_1199);
nor U1373 (N_1373,N_1038,N_1051);
or U1374 (N_1374,N_1145,N_1048);
or U1375 (N_1375,N_1152,N_1138);
and U1376 (N_1376,N_1089,N_1056);
nand U1377 (N_1377,N_1089,N_1124);
xnor U1378 (N_1378,N_1011,N_1191);
nor U1379 (N_1379,N_1151,N_1128);
or U1380 (N_1380,N_1185,N_1098);
and U1381 (N_1381,N_1038,N_1026);
nand U1382 (N_1382,N_1199,N_1008);
xnor U1383 (N_1383,N_1098,N_1064);
or U1384 (N_1384,N_1099,N_1134);
xor U1385 (N_1385,N_1032,N_1133);
nor U1386 (N_1386,N_1101,N_1157);
nor U1387 (N_1387,N_1066,N_1026);
nor U1388 (N_1388,N_1045,N_1009);
nand U1389 (N_1389,N_1198,N_1119);
xor U1390 (N_1390,N_1063,N_1168);
xor U1391 (N_1391,N_1005,N_1017);
nor U1392 (N_1392,N_1007,N_1183);
nor U1393 (N_1393,N_1097,N_1046);
nand U1394 (N_1394,N_1044,N_1106);
and U1395 (N_1395,N_1054,N_1148);
nor U1396 (N_1396,N_1069,N_1042);
nand U1397 (N_1397,N_1014,N_1159);
nand U1398 (N_1398,N_1117,N_1063);
nor U1399 (N_1399,N_1138,N_1119);
or U1400 (N_1400,N_1210,N_1388);
nand U1401 (N_1401,N_1353,N_1330);
or U1402 (N_1402,N_1366,N_1286);
xnor U1403 (N_1403,N_1242,N_1371);
and U1404 (N_1404,N_1253,N_1361);
nand U1405 (N_1405,N_1230,N_1274);
and U1406 (N_1406,N_1298,N_1305);
nand U1407 (N_1407,N_1394,N_1200);
or U1408 (N_1408,N_1204,N_1225);
or U1409 (N_1409,N_1382,N_1291);
and U1410 (N_1410,N_1288,N_1212);
nand U1411 (N_1411,N_1339,N_1297);
nor U1412 (N_1412,N_1292,N_1333);
or U1413 (N_1413,N_1293,N_1229);
nand U1414 (N_1414,N_1316,N_1273);
and U1415 (N_1415,N_1217,N_1215);
nor U1416 (N_1416,N_1250,N_1270);
xor U1417 (N_1417,N_1331,N_1369);
or U1418 (N_1418,N_1240,N_1268);
nand U1419 (N_1419,N_1251,N_1266);
and U1420 (N_1420,N_1348,N_1214);
xor U1421 (N_1421,N_1290,N_1231);
xnor U1422 (N_1422,N_1243,N_1258);
nor U1423 (N_1423,N_1314,N_1289);
xor U1424 (N_1424,N_1208,N_1319);
nor U1425 (N_1425,N_1301,N_1205);
nand U1426 (N_1426,N_1271,N_1350);
or U1427 (N_1427,N_1201,N_1381);
nor U1428 (N_1428,N_1279,N_1356);
or U1429 (N_1429,N_1307,N_1387);
and U1430 (N_1430,N_1312,N_1328);
and U1431 (N_1431,N_1284,N_1375);
nand U1432 (N_1432,N_1216,N_1222);
nor U1433 (N_1433,N_1396,N_1347);
xor U1434 (N_1434,N_1213,N_1302);
nor U1435 (N_1435,N_1317,N_1265);
nor U1436 (N_1436,N_1372,N_1327);
nor U1437 (N_1437,N_1376,N_1378);
and U1438 (N_1438,N_1337,N_1323);
nand U1439 (N_1439,N_1238,N_1300);
nor U1440 (N_1440,N_1232,N_1247);
and U1441 (N_1441,N_1219,N_1257);
and U1442 (N_1442,N_1335,N_1227);
or U1443 (N_1443,N_1248,N_1338);
nand U1444 (N_1444,N_1324,N_1278);
nand U1445 (N_1445,N_1373,N_1367);
and U1446 (N_1446,N_1392,N_1264);
xnor U1447 (N_1447,N_1377,N_1267);
nor U1448 (N_1448,N_1282,N_1263);
nor U1449 (N_1449,N_1340,N_1395);
or U1450 (N_1450,N_1386,N_1246);
nand U1451 (N_1451,N_1342,N_1351);
and U1452 (N_1452,N_1295,N_1383);
xnor U1453 (N_1453,N_1315,N_1393);
or U1454 (N_1454,N_1203,N_1304);
and U1455 (N_1455,N_1309,N_1255);
and U1456 (N_1456,N_1277,N_1202);
nand U1457 (N_1457,N_1385,N_1344);
nor U1458 (N_1458,N_1241,N_1397);
nor U1459 (N_1459,N_1233,N_1236);
nand U1460 (N_1460,N_1218,N_1234);
or U1461 (N_1461,N_1354,N_1380);
nand U1462 (N_1462,N_1363,N_1237);
nor U1463 (N_1463,N_1334,N_1310);
and U1464 (N_1464,N_1318,N_1332);
xnor U1465 (N_1465,N_1303,N_1220);
or U1466 (N_1466,N_1352,N_1357);
or U1467 (N_1467,N_1343,N_1209);
xor U1468 (N_1468,N_1249,N_1223);
or U1469 (N_1469,N_1374,N_1281);
nand U1470 (N_1470,N_1311,N_1325);
and U1471 (N_1471,N_1262,N_1245);
nand U1472 (N_1472,N_1260,N_1321);
nor U1473 (N_1473,N_1287,N_1364);
nand U1474 (N_1474,N_1384,N_1391);
nor U1475 (N_1475,N_1239,N_1320);
nand U1476 (N_1476,N_1256,N_1365);
and U1477 (N_1477,N_1329,N_1399);
nor U1478 (N_1478,N_1313,N_1360);
nor U1479 (N_1479,N_1276,N_1306);
and U1480 (N_1480,N_1349,N_1390);
or U1481 (N_1481,N_1206,N_1252);
nor U1482 (N_1482,N_1299,N_1368);
or U1483 (N_1483,N_1275,N_1261);
xnor U1484 (N_1484,N_1221,N_1355);
or U1485 (N_1485,N_1254,N_1336);
nor U1486 (N_1486,N_1226,N_1294);
or U1487 (N_1487,N_1283,N_1207);
or U1488 (N_1488,N_1296,N_1228);
and U1489 (N_1489,N_1359,N_1280);
or U1490 (N_1490,N_1259,N_1398);
xnor U1491 (N_1491,N_1379,N_1322);
nand U1492 (N_1492,N_1211,N_1285);
and U1493 (N_1493,N_1346,N_1389);
and U1494 (N_1494,N_1345,N_1358);
xor U1495 (N_1495,N_1235,N_1224);
nor U1496 (N_1496,N_1326,N_1269);
nor U1497 (N_1497,N_1308,N_1370);
or U1498 (N_1498,N_1362,N_1244);
and U1499 (N_1499,N_1341,N_1272);
and U1500 (N_1500,N_1244,N_1245);
nor U1501 (N_1501,N_1343,N_1297);
nand U1502 (N_1502,N_1353,N_1240);
or U1503 (N_1503,N_1212,N_1314);
or U1504 (N_1504,N_1342,N_1212);
nand U1505 (N_1505,N_1211,N_1204);
nor U1506 (N_1506,N_1318,N_1327);
nand U1507 (N_1507,N_1253,N_1393);
or U1508 (N_1508,N_1332,N_1275);
or U1509 (N_1509,N_1285,N_1391);
nand U1510 (N_1510,N_1322,N_1257);
nor U1511 (N_1511,N_1393,N_1314);
nand U1512 (N_1512,N_1330,N_1201);
and U1513 (N_1513,N_1339,N_1248);
nand U1514 (N_1514,N_1349,N_1388);
nor U1515 (N_1515,N_1274,N_1349);
nor U1516 (N_1516,N_1399,N_1391);
nand U1517 (N_1517,N_1245,N_1337);
nand U1518 (N_1518,N_1256,N_1265);
and U1519 (N_1519,N_1207,N_1210);
or U1520 (N_1520,N_1385,N_1355);
and U1521 (N_1521,N_1320,N_1310);
nor U1522 (N_1522,N_1303,N_1257);
nand U1523 (N_1523,N_1264,N_1379);
nor U1524 (N_1524,N_1243,N_1256);
nand U1525 (N_1525,N_1354,N_1294);
nor U1526 (N_1526,N_1382,N_1266);
or U1527 (N_1527,N_1283,N_1320);
nor U1528 (N_1528,N_1367,N_1229);
and U1529 (N_1529,N_1383,N_1261);
nand U1530 (N_1530,N_1218,N_1335);
and U1531 (N_1531,N_1372,N_1206);
and U1532 (N_1532,N_1392,N_1395);
nand U1533 (N_1533,N_1395,N_1282);
and U1534 (N_1534,N_1281,N_1326);
and U1535 (N_1535,N_1348,N_1296);
and U1536 (N_1536,N_1216,N_1380);
nor U1537 (N_1537,N_1273,N_1238);
xnor U1538 (N_1538,N_1285,N_1222);
xor U1539 (N_1539,N_1320,N_1242);
nand U1540 (N_1540,N_1370,N_1331);
nand U1541 (N_1541,N_1225,N_1280);
or U1542 (N_1542,N_1201,N_1364);
nor U1543 (N_1543,N_1323,N_1203);
xor U1544 (N_1544,N_1267,N_1238);
nand U1545 (N_1545,N_1374,N_1309);
and U1546 (N_1546,N_1335,N_1298);
or U1547 (N_1547,N_1375,N_1287);
or U1548 (N_1548,N_1280,N_1367);
and U1549 (N_1549,N_1343,N_1306);
or U1550 (N_1550,N_1360,N_1257);
or U1551 (N_1551,N_1320,N_1326);
and U1552 (N_1552,N_1252,N_1250);
and U1553 (N_1553,N_1372,N_1383);
nand U1554 (N_1554,N_1297,N_1236);
or U1555 (N_1555,N_1376,N_1249);
xor U1556 (N_1556,N_1231,N_1368);
nor U1557 (N_1557,N_1223,N_1283);
nand U1558 (N_1558,N_1325,N_1375);
nand U1559 (N_1559,N_1387,N_1399);
nor U1560 (N_1560,N_1304,N_1229);
nand U1561 (N_1561,N_1231,N_1289);
or U1562 (N_1562,N_1313,N_1332);
nor U1563 (N_1563,N_1383,N_1247);
or U1564 (N_1564,N_1232,N_1395);
nor U1565 (N_1565,N_1301,N_1350);
nand U1566 (N_1566,N_1371,N_1387);
or U1567 (N_1567,N_1285,N_1348);
nand U1568 (N_1568,N_1378,N_1328);
nor U1569 (N_1569,N_1303,N_1360);
nand U1570 (N_1570,N_1388,N_1259);
and U1571 (N_1571,N_1293,N_1370);
nor U1572 (N_1572,N_1216,N_1254);
and U1573 (N_1573,N_1289,N_1228);
nor U1574 (N_1574,N_1265,N_1328);
and U1575 (N_1575,N_1263,N_1274);
nor U1576 (N_1576,N_1297,N_1309);
nor U1577 (N_1577,N_1398,N_1339);
and U1578 (N_1578,N_1251,N_1368);
nand U1579 (N_1579,N_1311,N_1323);
nor U1580 (N_1580,N_1288,N_1388);
and U1581 (N_1581,N_1230,N_1352);
nor U1582 (N_1582,N_1380,N_1361);
nand U1583 (N_1583,N_1272,N_1263);
nand U1584 (N_1584,N_1297,N_1229);
or U1585 (N_1585,N_1269,N_1235);
nor U1586 (N_1586,N_1209,N_1334);
xor U1587 (N_1587,N_1212,N_1348);
nand U1588 (N_1588,N_1225,N_1312);
or U1589 (N_1589,N_1345,N_1224);
and U1590 (N_1590,N_1367,N_1318);
nand U1591 (N_1591,N_1366,N_1276);
nand U1592 (N_1592,N_1306,N_1323);
xnor U1593 (N_1593,N_1235,N_1292);
nand U1594 (N_1594,N_1361,N_1240);
nor U1595 (N_1595,N_1373,N_1344);
xnor U1596 (N_1596,N_1255,N_1319);
nand U1597 (N_1597,N_1359,N_1326);
nand U1598 (N_1598,N_1241,N_1333);
nor U1599 (N_1599,N_1256,N_1390);
and U1600 (N_1600,N_1535,N_1486);
nand U1601 (N_1601,N_1495,N_1460);
nand U1602 (N_1602,N_1430,N_1477);
nand U1603 (N_1603,N_1435,N_1407);
or U1604 (N_1604,N_1511,N_1421);
and U1605 (N_1605,N_1413,N_1493);
or U1606 (N_1606,N_1573,N_1464);
nand U1607 (N_1607,N_1497,N_1592);
nand U1608 (N_1608,N_1414,N_1499);
and U1609 (N_1609,N_1594,N_1523);
and U1610 (N_1610,N_1540,N_1510);
nor U1611 (N_1611,N_1527,N_1491);
nor U1612 (N_1612,N_1564,N_1474);
and U1613 (N_1613,N_1480,N_1580);
xor U1614 (N_1614,N_1508,N_1530);
nand U1615 (N_1615,N_1526,N_1471);
nand U1616 (N_1616,N_1468,N_1431);
or U1617 (N_1617,N_1403,N_1498);
nand U1618 (N_1618,N_1465,N_1574);
or U1619 (N_1619,N_1475,N_1507);
or U1620 (N_1620,N_1448,N_1541);
nand U1621 (N_1621,N_1583,N_1452);
nand U1622 (N_1622,N_1536,N_1406);
and U1623 (N_1623,N_1418,N_1555);
nand U1624 (N_1624,N_1449,N_1445);
xor U1625 (N_1625,N_1416,N_1588);
xor U1626 (N_1626,N_1405,N_1590);
nand U1627 (N_1627,N_1542,N_1479);
xnor U1628 (N_1628,N_1504,N_1482);
nor U1629 (N_1629,N_1478,N_1593);
and U1630 (N_1630,N_1457,N_1500);
nand U1631 (N_1631,N_1562,N_1550);
and U1632 (N_1632,N_1549,N_1556);
nor U1633 (N_1633,N_1489,N_1424);
nor U1634 (N_1634,N_1463,N_1488);
and U1635 (N_1635,N_1447,N_1476);
and U1636 (N_1636,N_1534,N_1568);
nand U1637 (N_1637,N_1567,N_1554);
xor U1638 (N_1638,N_1422,N_1432);
nand U1639 (N_1639,N_1492,N_1485);
nand U1640 (N_1640,N_1505,N_1553);
nand U1641 (N_1641,N_1538,N_1563);
nor U1642 (N_1642,N_1533,N_1557);
and U1643 (N_1643,N_1579,N_1454);
and U1644 (N_1644,N_1446,N_1461);
xor U1645 (N_1645,N_1515,N_1569);
nand U1646 (N_1646,N_1455,N_1419);
nand U1647 (N_1647,N_1521,N_1524);
or U1648 (N_1648,N_1427,N_1501);
and U1649 (N_1649,N_1441,N_1514);
and U1650 (N_1650,N_1467,N_1575);
nand U1651 (N_1651,N_1528,N_1494);
nand U1652 (N_1652,N_1428,N_1577);
nor U1653 (N_1653,N_1581,N_1599);
or U1654 (N_1654,N_1423,N_1437);
and U1655 (N_1655,N_1596,N_1543);
nand U1656 (N_1656,N_1525,N_1576);
nor U1657 (N_1657,N_1412,N_1444);
and U1658 (N_1658,N_1560,N_1509);
nand U1659 (N_1659,N_1484,N_1539);
nand U1660 (N_1660,N_1566,N_1496);
and U1661 (N_1661,N_1531,N_1582);
and U1662 (N_1662,N_1439,N_1451);
nor U1663 (N_1663,N_1544,N_1597);
and U1664 (N_1664,N_1410,N_1547);
or U1665 (N_1665,N_1462,N_1506);
nand U1666 (N_1666,N_1522,N_1402);
and U1667 (N_1667,N_1561,N_1470);
and U1668 (N_1668,N_1529,N_1595);
nand U1669 (N_1669,N_1589,N_1584);
or U1670 (N_1670,N_1436,N_1442);
xor U1671 (N_1671,N_1516,N_1572);
and U1672 (N_1672,N_1466,N_1585);
nand U1673 (N_1673,N_1425,N_1415);
or U1674 (N_1674,N_1537,N_1552);
xor U1675 (N_1675,N_1559,N_1490);
and U1676 (N_1676,N_1481,N_1456);
nor U1677 (N_1677,N_1591,N_1426);
nand U1678 (N_1678,N_1571,N_1503);
nor U1679 (N_1679,N_1532,N_1517);
or U1680 (N_1680,N_1586,N_1400);
nor U1681 (N_1681,N_1408,N_1411);
nand U1682 (N_1682,N_1519,N_1401);
and U1683 (N_1683,N_1458,N_1459);
nand U1684 (N_1684,N_1429,N_1518);
nor U1685 (N_1685,N_1440,N_1558);
nand U1686 (N_1686,N_1443,N_1551);
and U1687 (N_1687,N_1404,N_1578);
or U1688 (N_1688,N_1450,N_1420);
and U1689 (N_1689,N_1433,N_1565);
nand U1690 (N_1690,N_1472,N_1598);
nand U1691 (N_1691,N_1545,N_1434);
nand U1692 (N_1692,N_1409,N_1548);
and U1693 (N_1693,N_1483,N_1570);
and U1694 (N_1694,N_1513,N_1520);
nand U1695 (N_1695,N_1546,N_1502);
xor U1696 (N_1696,N_1469,N_1487);
nor U1697 (N_1697,N_1587,N_1473);
and U1698 (N_1698,N_1453,N_1512);
nor U1699 (N_1699,N_1417,N_1438);
nand U1700 (N_1700,N_1511,N_1468);
or U1701 (N_1701,N_1576,N_1505);
and U1702 (N_1702,N_1519,N_1597);
nand U1703 (N_1703,N_1517,N_1573);
nand U1704 (N_1704,N_1492,N_1574);
nand U1705 (N_1705,N_1476,N_1514);
nor U1706 (N_1706,N_1529,N_1547);
and U1707 (N_1707,N_1444,N_1502);
nor U1708 (N_1708,N_1482,N_1507);
or U1709 (N_1709,N_1516,N_1589);
nand U1710 (N_1710,N_1455,N_1558);
nand U1711 (N_1711,N_1541,N_1487);
nand U1712 (N_1712,N_1459,N_1582);
nor U1713 (N_1713,N_1521,N_1405);
nor U1714 (N_1714,N_1539,N_1425);
and U1715 (N_1715,N_1490,N_1567);
or U1716 (N_1716,N_1590,N_1486);
nor U1717 (N_1717,N_1556,N_1550);
or U1718 (N_1718,N_1516,N_1462);
xor U1719 (N_1719,N_1422,N_1511);
and U1720 (N_1720,N_1436,N_1560);
and U1721 (N_1721,N_1533,N_1586);
xnor U1722 (N_1722,N_1424,N_1599);
nor U1723 (N_1723,N_1530,N_1589);
or U1724 (N_1724,N_1426,N_1531);
nand U1725 (N_1725,N_1404,N_1456);
nand U1726 (N_1726,N_1567,N_1594);
xor U1727 (N_1727,N_1470,N_1585);
or U1728 (N_1728,N_1476,N_1550);
xnor U1729 (N_1729,N_1450,N_1518);
nand U1730 (N_1730,N_1537,N_1503);
nor U1731 (N_1731,N_1448,N_1499);
and U1732 (N_1732,N_1506,N_1477);
and U1733 (N_1733,N_1490,N_1430);
nor U1734 (N_1734,N_1519,N_1405);
and U1735 (N_1735,N_1437,N_1510);
nand U1736 (N_1736,N_1512,N_1563);
and U1737 (N_1737,N_1502,N_1449);
and U1738 (N_1738,N_1549,N_1585);
nor U1739 (N_1739,N_1423,N_1561);
nand U1740 (N_1740,N_1511,N_1501);
nor U1741 (N_1741,N_1416,N_1471);
and U1742 (N_1742,N_1456,N_1402);
nand U1743 (N_1743,N_1499,N_1583);
xor U1744 (N_1744,N_1567,N_1597);
and U1745 (N_1745,N_1497,N_1488);
xor U1746 (N_1746,N_1446,N_1491);
nor U1747 (N_1747,N_1466,N_1419);
and U1748 (N_1748,N_1433,N_1400);
and U1749 (N_1749,N_1529,N_1467);
or U1750 (N_1750,N_1497,N_1475);
nor U1751 (N_1751,N_1593,N_1437);
and U1752 (N_1752,N_1583,N_1455);
and U1753 (N_1753,N_1438,N_1511);
nand U1754 (N_1754,N_1400,N_1436);
nand U1755 (N_1755,N_1513,N_1445);
nand U1756 (N_1756,N_1598,N_1581);
nand U1757 (N_1757,N_1517,N_1599);
and U1758 (N_1758,N_1514,N_1439);
and U1759 (N_1759,N_1443,N_1407);
nor U1760 (N_1760,N_1562,N_1582);
xnor U1761 (N_1761,N_1541,N_1561);
xnor U1762 (N_1762,N_1528,N_1531);
nor U1763 (N_1763,N_1466,N_1530);
or U1764 (N_1764,N_1464,N_1512);
nand U1765 (N_1765,N_1535,N_1595);
xor U1766 (N_1766,N_1486,N_1542);
and U1767 (N_1767,N_1461,N_1533);
and U1768 (N_1768,N_1584,N_1511);
and U1769 (N_1769,N_1486,N_1461);
and U1770 (N_1770,N_1405,N_1585);
nand U1771 (N_1771,N_1501,N_1588);
and U1772 (N_1772,N_1434,N_1445);
or U1773 (N_1773,N_1485,N_1532);
or U1774 (N_1774,N_1579,N_1411);
xor U1775 (N_1775,N_1547,N_1519);
nand U1776 (N_1776,N_1531,N_1465);
nand U1777 (N_1777,N_1450,N_1539);
nand U1778 (N_1778,N_1434,N_1485);
xnor U1779 (N_1779,N_1438,N_1542);
and U1780 (N_1780,N_1574,N_1570);
or U1781 (N_1781,N_1586,N_1525);
nand U1782 (N_1782,N_1523,N_1589);
and U1783 (N_1783,N_1566,N_1558);
nor U1784 (N_1784,N_1488,N_1437);
nor U1785 (N_1785,N_1452,N_1465);
and U1786 (N_1786,N_1574,N_1550);
xor U1787 (N_1787,N_1451,N_1445);
nand U1788 (N_1788,N_1541,N_1405);
nor U1789 (N_1789,N_1510,N_1499);
and U1790 (N_1790,N_1471,N_1591);
nor U1791 (N_1791,N_1464,N_1451);
nand U1792 (N_1792,N_1496,N_1569);
nand U1793 (N_1793,N_1525,N_1470);
and U1794 (N_1794,N_1558,N_1418);
nand U1795 (N_1795,N_1570,N_1567);
and U1796 (N_1796,N_1465,N_1584);
or U1797 (N_1797,N_1591,N_1586);
xor U1798 (N_1798,N_1476,N_1546);
nor U1799 (N_1799,N_1532,N_1548);
nor U1800 (N_1800,N_1750,N_1649);
nand U1801 (N_1801,N_1616,N_1703);
and U1802 (N_1802,N_1610,N_1661);
or U1803 (N_1803,N_1617,N_1658);
nand U1804 (N_1804,N_1612,N_1692);
nand U1805 (N_1805,N_1621,N_1728);
nand U1806 (N_1806,N_1682,N_1717);
nor U1807 (N_1807,N_1638,N_1714);
nand U1808 (N_1808,N_1761,N_1643);
nor U1809 (N_1809,N_1758,N_1746);
and U1810 (N_1810,N_1716,N_1735);
nand U1811 (N_1811,N_1672,N_1653);
and U1812 (N_1812,N_1640,N_1744);
and U1813 (N_1813,N_1600,N_1702);
and U1814 (N_1814,N_1724,N_1655);
or U1815 (N_1815,N_1727,N_1693);
or U1816 (N_1816,N_1722,N_1700);
and U1817 (N_1817,N_1681,N_1689);
nand U1818 (N_1818,N_1764,N_1632);
and U1819 (N_1819,N_1776,N_1601);
or U1820 (N_1820,N_1603,N_1797);
nand U1821 (N_1821,N_1705,N_1721);
nor U1822 (N_1822,N_1633,N_1747);
nor U1823 (N_1823,N_1790,N_1707);
nand U1824 (N_1824,N_1699,N_1711);
and U1825 (N_1825,N_1737,N_1696);
nand U1826 (N_1826,N_1765,N_1652);
or U1827 (N_1827,N_1626,N_1697);
and U1828 (N_1828,N_1730,N_1629);
and U1829 (N_1829,N_1627,N_1794);
nand U1830 (N_1830,N_1745,N_1767);
or U1831 (N_1831,N_1656,N_1679);
and U1832 (N_1832,N_1650,N_1720);
and U1833 (N_1833,N_1671,N_1694);
or U1834 (N_1834,N_1718,N_1607);
nand U1835 (N_1835,N_1686,N_1662);
nand U1836 (N_1836,N_1732,N_1795);
or U1837 (N_1837,N_1788,N_1611);
xor U1838 (N_1838,N_1754,N_1783);
and U1839 (N_1839,N_1787,N_1622);
or U1840 (N_1840,N_1615,N_1753);
or U1841 (N_1841,N_1719,N_1775);
nor U1842 (N_1842,N_1614,N_1784);
nand U1843 (N_1843,N_1698,N_1796);
and U1844 (N_1844,N_1789,N_1709);
and U1845 (N_1845,N_1676,N_1663);
or U1846 (N_1846,N_1646,N_1706);
or U1847 (N_1847,N_1779,N_1624);
nand U1848 (N_1848,N_1602,N_1618);
and U1849 (N_1849,N_1736,N_1659);
and U1850 (N_1850,N_1799,N_1741);
nand U1851 (N_1851,N_1628,N_1680);
or U1852 (N_1852,N_1791,N_1773);
and U1853 (N_1853,N_1670,N_1778);
and U1854 (N_1854,N_1613,N_1757);
and U1855 (N_1855,N_1708,N_1623);
or U1856 (N_1856,N_1620,N_1704);
and U1857 (N_1857,N_1723,N_1738);
xor U1858 (N_1858,N_1664,N_1654);
nor U1859 (N_1859,N_1760,N_1635);
nor U1860 (N_1860,N_1740,N_1798);
nor U1861 (N_1861,N_1685,N_1637);
or U1862 (N_1862,N_1726,N_1641);
or U1863 (N_1863,N_1763,N_1642);
or U1864 (N_1864,N_1665,N_1648);
or U1865 (N_1865,N_1668,N_1725);
or U1866 (N_1866,N_1781,N_1608);
or U1867 (N_1867,N_1606,N_1712);
and U1868 (N_1868,N_1634,N_1675);
and U1869 (N_1869,N_1645,N_1770);
and U1870 (N_1870,N_1678,N_1625);
nand U1871 (N_1871,N_1793,N_1639);
or U1872 (N_1872,N_1762,N_1710);
nand U1873 (N_1873,N_1691,N_1631);
xor U1874 (N_1874,N_1739,N_1690);
and U1875 (N_1875,N_1669,N_1743);
nand U1876 (N_1876,N_1666,N_1752);
nor U1877 (N_1877,N_1772,N_1701);
xnor U1878 (N_1878,N_1636,N_1715);
or U1879 (N_1879,N_1657,N_1609);
or U1880 (N_1880,N_1673,N_1604);
nor U1881 (N_1881,N_1683,N_1786);
nor U1882 (N_1882,N_1713,N_1687);
nand U1883 (N_1883,N_1688,N_1684);
and U1884 (N_1884,N_1729,N_1768);
nor U1885 (N_1885,N_1674,N_1667);
xor U1886 (N_1886,N_1660,N_1751);
nor U1887 (N_1887,N_1644,N_1777);
nor U1888 (N_1888,N_1605,N_1677);
nand U1889 (N_1889,N_1792,N_1766);
or U1890 (N_1890,N_1749,N_1733);
and U1891 (N_1891,N_1782,N_1651);
nand U1892 (N_1892,N_1647,N_1756);
nor U1893 (N_1893,N_1731,N_1748);
nor U1894 (N_1894,N_1774,N_1742);
and U1895 (N_1895,N_1759,N_1734);
nand U1896 (N_1896,N_1769,N_1695);
nor U1897 (N_1897,N_1780,N_1630);
or U1898 (N_1898,N_1771,N_1785);
xor U1899 (N_1899,N_1755,N_1619);
or U1900 (N_1900,N_1776,N_1785);
or U1901 (N_1901,N_1767,N_1627);
nor U1902 (N_1902,N_1613,N_1624);
nand U1903 (N_1903,N_1680,N_1645);
nand U1904 (N_1904,N_1791,N_1674);
and U1905 (N_1905,N_1655,N_1786);
nand U1906 (N_1906,N_1698,N_1799);
or U1907 (N_1907,N_1630,N_1711);
and U1908 (N_1908,N_1737,N_1728);
or U1909 (N_1909,N_1733,N_1663);
or U1910 (N_1910,N_1742,N_1718);
nand U1911 (N_1911,N_1610,N_1679);
xor U1912 (N_1912,N_1620,N_1753);
and U1913 (N_1913,N_1774,N_1677);
nand U1914 (N_1914,N_1677,N_1798);
nand U1915 (N_1915,N_1671,N_1634);
and U1916 (N_1916,N_1778,N_1634);
nand U1917 (N_1917,N_1772,N_1784);
or U1918 (N_1918,N_1782,N_1797);
or U1919 (N_1919,N_1722,N_1749);
nand U1920 (N_1920,N_1681,N_1643);
and U1921 (N_1921,N_1723,N_1686);
nor U1922 (N_1922,N_1700,N_1778);
or U1923 (N_1923,N_1679,N_1702);
nand U1924 (N_1924,N_1766,N_1718);
nor U1925 (N_1925,N_1781,N_1707);
or U1926 (N_1926,N_1795,N_1765);
nand U1927 (N_1927,N_1706,N_1602);
nand U1928 (N_1928,N_1708,N_1658);
or U1929 (N_1929,N_1647,N_1720);
and U1930 (N_1930,N_1609,N_1775);
nor U1931 (N_1931,N_1661,N_1611);
nor U1932 (N_1932,N_1624,N_1660);
nor U1933 (N_1933,N_1683,N_1633);
nor U1934 (N_1934,N_1750,N_1671);
or U1935 (N_1935,N_1751,N_1733);
or U1936 (N_1936,N_1681,N_1757);
and U1937 (N_1937,N_1649,N_1748);
and U1938 (N_1938,N_1752,N_1613);
xor U1939 (N_1939,N_1688,N_1639);
or U1940 (N_1940,N_1600,N_1668);
and U1941 (N_1941,N_1716,N_1660);
or U1942 (N_1942,N_1764,N_1707);
and U1943 (N_1943,N_1610,N_1736);
nor U1944 (N_1944,N_1646,N_1745);
xor U1945 (N_1945,N_1654,N_1650);
nand U1946 (N_1946,N_1695,N_1780);
nor U1947 (N_1947,N_1677,N_1737);
and U1948 (N_1948,N_1639,N_1767);
and U1949 (N_1949,N_1705,N_1707);
xor U1950 (N_1950,N_1678,N_1605);
nor U1951 (N_1951,N_1673,N_1749);
nand U1952 (N_1952,N_1746,N_1708);
nand U1953 (N_1953,N_1789,N_1671);
nand U1954 (N_1954,N_1692,N_1794);
and U1955 (N_1955,N_1670,N_1666);
nor U1956 (N_1956,N_1791,N_1783);
and U1957 (N_1957,N_1634,N_1667);
nor U1958 (N_1958,N_1646,N_1695);
nand U1959 (N_1959,N_1745,N_1735);
nor U1960 (N_1960,N_1699,N_1759);
or U1961 (N_1961,N_1718,N_1786);
nand U1962 (N_1962,N_1752,N_1629);
nor U1963 (N_1963,N_1784,N_1714);
nand U1964 (N_1964,N_1677,N_1607);
nand U1965 (N_1965,N_1660,N_1691);
nand U1966 (N_1966,N_1798,N_1708);
nor U1967 (N_1967,N_1633,N_1711);
or U1968 (N_1968,N_1649,N_1629);
and U1969 (N_1969,N_1754,N_1729);
nand U1970 (N_1970,N_1746,N_1667);
nor U1971 (N_1971,N_1729,N_1755);
xor U1972 (N_1972,N_1774,N_1664);
or U1973 (N_1973,N_1601,N_1766);
and U1974 (N_1974,N_1635,N_1765);
nand U1975 (N_1975,N_1705,N_1600);
and U1976 (N_1976,N_1606,N_1750);
nand U1977 (N_1977,N_1694,N_1765);
nand U1978 (N_1978,N_1717,N_1728);
and U1979 (N_1979,N_1763,N_1738);
xnor U1980 (N_1980,N_1636,N_1743);
or U1981 (N_1981,N_1755,N_1659);
nand U1982 (N_1982,N_1626,N_1724);
or U1983 (N_1983,N_1755,N_1718);
and U1984 (N_1984,N_1746,N_1786);
nand U1985 (N_1985,N_1716,N_1601);
and U1986 (N_1986,N_1624,N_1641);
or U1987 (N_1987,N_1706,N_1749);
and U1988 (N_1988,N_1696,N_1628);
nand U1989 (N_1989,N_1608,N_1643);
nor U1990 (N_1990,N_1630,N_1737);
xor U1991 (N_1991,N_1642,N_1710);
nand U1992 (N_1992,N_1786,N_1764);
xor U1993 (N_1993,N_1678,N_1763);
nand U1994 (N_1994,N_1635,N_1637);
nand U1995 (N_1995,N_1706,N_1670);
or U1996 (N_1996,N_1761,N_1625);
nand U1997 (N_1997,N_1605,N_1719);
or U1998 (N_1998,N_1755,N_1719);
nand U1999 (N_1999,N_1701,N_1775);
nand U2000 (N_2000,N_1982,N_1814);
nand U2001 (N_2001,N_1826,N_1876);
and U2002 (N_2002,N_1924,N_1855);
or U2003 (N_2003,N_1950,N_1811);
xnor U2004 (N_2004,N_1909,N_1887);
and U2005 (N_2005,N_1917,N_1904);
nor U2006 (N_2006,N_1945,N_1864);
nand U2007 (N_2007,N_1978,N_1852);
nand U2008 (N_2008,N_1821,N_1988);
and U2009 (N_2009,N_1835,N_1949);
xor U2010 (N_2010,N_1856,N_1804);
nor U2011 (N_2011,N_1812,N_1873);
xor U2012 (N_2012,N_1891,N_1997);
or U2013 (N_2013,N_1933,N_1823);
and U2014 (N_2014,N_1942,N_1952);
nor U2015 (N_2015,N_1889,N_1888);
and U2016 (N_2016,N_1871,N_1987);
and U2017 (N_2017,N_1870,N_1931);
nor U2018 (N_2018,N_1866,N_1934);
nand U2019 (N_2019,N_1863,N_1808);
nand U2020 (N_2020,N_1854,N_1807);
and U2021 (N_2021,N_1972,N_1970);
or U2022 (N_2022,N_1968,N_1913);
nor U2023 (N_2023,N_1953,N_1869);
or U2024 (N_2024,N_1928,N_1960);
nor U2025 (N_2025,N_1885,N_1989);
and U2026 (N_2026,N_1974,N_1940);
and U2027 (N_2027,N_1976,N_1813);
nand U2028 (N_2028,N_1892,N_1925);
or U2029 (N_2029,N_1882,N_1877);
nor U2030 (N_2030,N_1963,N_1837);
xnor U2031 (N_2031,N_1958,N_1943);
or U2032 (N_2032,N_1944,N_1858);
or U2033 (N_2033,N_1985,N_1966);
and U2034 (N_2034,N_1916,N_1860);
nor U2035 (N_2035,N_1906,N_1810);
nand U2036 (N_2036,N_1842,N_1859);
xnor U2037 (N_2037,N_1971,N_1959);
and U2038 (N_2038,N_1907,N_1938);
or U2039 (N_2039,N_1926,N_1818);
nor U2040 (N_2040,N_1845,N_1896);
nand U2041 (N_2041,N_1956,N_1836);
nand U2042 (N_2042,N_1946,N_1922);
nor U2043 (N_2043,N_1912,N_1830);
and U2044 (N_2044,N_1822,N_1857);
and U2045 (N_2045,N_1880,N_1851);
nand U2046 (N_2046,N_1827,N_1941);
nand U2047 (N_2047,N_1905,N_1990);
or U2048 (N_2048,N_1894,N_1805);
xor U2049 (N_2049,N_1999,N_1964);
nand U2050 (N_2050,N_1948,N_1802);
or U2051 (N_2051,N_1967,N_1868);
nor U2052 (N_2052,N_1824,N_1996);
or U2053 (N_2053,N_1803,N_1923);
or U2054 (N_2054,N_1844,N_1914);
xor U2055 (N_2055,N_1874,N_1815);
nand U2056 (N_2056,N_1881,N_1910);
nor U2057 (N_2057,N_1919,N_1834);
xor U2058 (N_2058,N_1861,N_1902);
nand U2059 (N_2059,N_1800,N_1862);
and U2060 (N_2060,N_1825,N_1962);
and U2061 (N_2061,N_1979,N_1981);
and U2062 (N_2062,N_1937,N_1901);
and U2063 (N_2063,N_1995,N_1927);
and U2064 (N_2064,N_1975,N_1932);
nand U2065 (N_2065,N_1961,N_1977);
and U2066 (N_2066,N_1838,N_1947);
and U2067 (N_2067,N_1936,N_1930);
nor U2068 (N_2068,N_1893,N_1983);
nor U2069 (N_2069,N_1897,N_1839);
and U2070 (N_2070,N_1991,N_1890);
xor U2071 (N_2071,N_1899,N_1921);
and U2072 (N_2072,N_1957,N_1867);
and U2073 (N_2073,N_1820,N_1955);
nand U2074 (N_2074,N_1850,N_1898);
xnor U2075 (N_2075,N_1915,N_1833);
nor U2076 (N_2076,N_1843,N_1828);
nand U2077 (N_2077,N_1986,N_1816);
nor U2078 (N_2078,N_1900,N_1992);
and U2079 (N_2079,N_1875,N_1969);
xnor U2080 (N_2080,N_1929,N_1809);
and U2081 (N_2081,N_1819,N_1984);
nand U2082 (N_2082,N_1883,N_1951);
or U2083 (N_2083,N_1806,N_1878);
xor U2084 (N_2084,N_1998,N_1848);
nor U2085 (N_2085,N_1832,N_1965);
nand U2086 (N_2086,N_1884,N_1920);
or U2087 (N_2087,N_1841,N_1817);
or U2088 (N_2088,N_1853,N_1879);
or U2089 (N_2089,N_1886,N_1973);
and U2090 (N_2090,N_1829,N_1849);
nand U2091 (N_2091,N_1939,N_1801);
nand U2092 (N_2092,N_1872,N_1911);
and U2093 (N_2093,N_1994,N_1846);
or U2094 (N_2094,N_1993,N_1903);
or U2095 (N_2095,N_1840,N_1918);
nand U2096 (N_2096,N_1935,N_1831);
nor U2097 (N_2097,N_1847,N_1865);
or U2098 (N_2098,N_1908,N_1954);
xor U2099 (N_2099,N_1980,N_1895);
nand U2100 (N_2100,N_1934,N_1872);
and U2101 (N_2101,N_1862,N_1925);
nand U2102 (N_2102,N_1823,N_1932);
and U2103 (N_2103,N_1847,N_1955);
nor U2104 (N_2104,N_1880,N_1815);
nand U2105 (N_2105,N_1827,N_1911);
xnor U2106 (N_2106,N_1979,N_1990);
nand U2107 (N_2107,N_1805,N_1965);
xor U2108 (N_2108,N_1892,N_1997);
nand U2109 (N_2109,N_1948,N_1984);
or U2110 (N_2110,N_1802,N_1911);
or U2111 (N_2111,N_1828,N_1896);
nand U2112 (N_2112,N_1896,N_1971);
or U2113 (N_2113,N_1854,N_1814);
nor U2114 (N_2114,N_1978,N_1905);
or U2115 (N_2115,N_1832,N_1996);
xor U2116 (N_2116,N_1897,N_1830);
or U2117 (N_2117,N_1881,N_1987);
xnor U2118 (N_2118,N_1899,N_1906);
xor U2119 (N_2119,N_1892,N_1973);
nand U2120 (N_2120,N_1810,N_1836);
and U2121 (N_2121,N_1874,N_1853);
nand U2122 (N_2122,N_1841,N_1934);
and U2123 (N_2123,N_1957,N_1994);
and U2124 (N_2124,N_1858,N_1965);
nor U2125 (N_2125,N_1921,N_1862);
or U2126 (N_2126,N_1834,N_1992);
or U2127 (N_2127,N_1940,N_1995);
nor U2128 (N_2128,N_1853,N_1983);
nor U2129 (N_2129,N_1887,N_1973);
and U2130 (N_2130,N_1817,N_1963);
nor U2131 (N_2131,N_1975,N_1985);
nand U2132 (N_2132,N_1985,N_1814);
or U2133 (N_2133,N_1860,N_1848);
nor U2134 (N_2134,N_1850,N_1870);
and U2135 (N_2135,N_1876,N_1881);
or U2136 (N_2136,N_1850,N_1922);
and U2137 (N_2137,N_1881,N_1994);
nor U2138 (N_2138,N_1878,N_1894);
or U2139 (N_2139,N_1861,N_1921);
or U2140 (N_2140,N_1899,N_1806);
or U2141 (N_2141,N_1806,N_1926);
nand U2142 (N_2142,N_1970,N_1917);
xnor U2143 (N_2143,N_1977,N_1979);
or U2144 (N_2144,N_1833,N_1884);
nor U2145 (N_2145,N_1932,N_1826);
and U2146 (N_2146,N_1911,N_1992);
xnor U2147 (N_2147,N_1964,N_1904);
and U2148 (N_2148,N_1808,N_1993);
or U2149 (N_2149,N_1906,N_1813);
and U2150 (N_2150,N_1921,N_1935);
and U2151 (N_2151,N_1866,N_1851);
nor U2152 (N_2152,N_1957,N_1924);
xnor U2153 (N_2153,N_1864,N_1902);
or U2154 (N_2154,N_1834,N_1940);
nand U2155 (N_2155,N_1800,N_1950);
or U2156 (N_2156,N_1994,N_1823);
nor U2157 (N_2157,N_1921,N_1801);
or U2158 (N_2158,N_1875,N_1924);
nand U2159 (N_2159,N_1837,N_1847);
or U2160 (N_2160,N_1824,N_1815);
and U2161 (N_2161,N_1821,N_1956);
or U2162 (N_2162,N_1951,N_1847);
and U2163 (N_2163,N_1954,N_1898);
and U2164 (N_2164,N_1807,N_1834);
nand U2165 (N_2165,N_1934,N_1806);
and U2166 (N_2166,N_1984,N_1908);
nand U2167 (N_2167,N_1932,N_1868);
nand U2168 (N_2168,N_1994,N_1909);
xor U2169 (N_2169,N_1974,N_1807);
nor U2170 (N_2170,N_1819,N_1910);
nand U2171 (N_2171,N_1954,N_1819);
or U2172 (N_2172,N_1931,N_1989);
and U2173 (N_2173,N_1913,N_1834);
or U2174 (N_2174,N_1989,N_1971);
and U2175 (N_2175,N_1914,N_1837);
nand U2176 (N_2176,N_1941,N_1962);
nand U2177 (N_2177,N_1889,N_1860);
nand U2178 (N_2178,N_1899,N_1960);
nand U2179 (N_2179,N_1827,N_1819);
and U2180 (N_2180,N_1896,N_1998);
nand U2181 (N_2181,N_1974,N_1913);
and U2182 (N_2182,N_1969,N_1898);
or U2183 (N_2183,N_1832,N_1807);
xnor U2184 (N_2184,N_1922,N_1812);
nor U2185 (N_2185,N_1998,N_1828);
and U2186 (N_2186,N_1973,N_1846);
nor U2187 (N_2187,N_1883,N_1847);
nand U2188 (N_2188,N_1927,N_1813);
xnor U2189 (N_2189,N_1800,N_1998);
or U2190 (N_2190,N_1943,N_1955);
nor U2191 (N_2191,N_1893,N_1997);
or U2192 (N_2192,N_1811,N_1968);
and U2193 (N_2193,N_1978,N_1898);
xor U2194 (N_2194,N_1830,N_1833);
or U2195 (N_2195,N_1831,N_1872);
nor U2196 (N_2196,N_1812,N_1975);
or U2197 (N_2197,N_1991,N_1843);
or U2198 (N_2198,N_1959,N_1933);
nor U2199 (N_2199,N_1841,N_1992);
and U2200 (N_2200,N_2139,N_2126);
nand U2201 (N_2201,N_2000,N_2098);
nand U2202 (N_2202,N_2152,N_2196);
nand U2203 (N_2203,N_2052,N_2107);
nor U2204 (N_2204,N_2013,N_2124);
and U2205 (N_2205,N_2031,N_2004);
nor U2206 (N_2206,N_2072,N_2096);
nor U2207 (N_2207,N_2050,N_2033);
and U2208 (N_2208,N_2009,N_2164);
and U2209 (N_2209,N_2112,N_2066);
or U2210 (N_2210,N_2039,N_2155);
nor U2211 (N_2211,N_2058,N_2060);
nand U2212 (N_2212,N_2083,N_2153);
nor U2213 (N_2213,N_2119,N_2195);
or U2214 (N_2214,N_2006,N_2190);
or U2215 (N_2215,N_2169,N_2117);
and U2216 (N_2216,N_2014,N_2010);
and U2217 (N_2217,N_2192,N_2175);
or U2218 (N_2218,N_2108,N_2015);
nor U2219 (N_2219,N_2061,N_2043);
or U2220 (N_2220,N_2162,N_2046);
and U2221 (N_2221,N_2178,N_2054);
or U2222 (N_2222,N_2069,N_2145);
xnor U2223 (N_2223,N_2021,N_2005);
nor U2224 (N_2224,N_2084,N_2064);
nor U2225 (N_2225,N_2129,N_2148);
xnor U2226 (N_2226,N_2103,N_2104);
nand U2227 (N_2227,N_2076,N_2095);
or U2228 (N_2228,N_2194,N_2048);
nand U2229 (N_2229,N_2197,N_2147);
nor U2230 (N_2230,N_2174,N_2041);
nand U2231 (N_2231,N_2156,N_2063);
or U2232 (N_2232,N_2193,N_2020);
and U2233 (N_2233,N_2062,N_2167);
or U2234 (N_2234,N_2057,N_2089);
and U2235 (N_2235,N_2105,N_2172);
or U2236 (N_2236,N_2027,N_2132);
or U2237 (N_2237,N_2093,N_2055);
and U2238 (N_2238,N_2091,N_2179);
or U2239 (N_2239,N_2019,N_2012);
nand U2240 (N_2240,N_2073,N_2077);
xnor U2241 (N_2241,N_2199,N_2036);
and U2242 (N_2242,N_2128,N_2051);
nand U2243 (N_2243,N_2163,N_2151);
xnor U2244 (N_2244,N_2047,N_2102);
and U2245 (N_2245,N_2059,N_2053);
or U2246 (N_2246,N_2184,N_2024);
nor U2247 (N_2247,N_2100,N_2088);
or U2248 (N_2248,N_2113,N_2092);
nor U2249 (N_2249,N_2008,N_2186);
nor U2250 (N_2250,N_2028,N_2165);
nand U2251 (N_2251,N_2017,N_2142);
nor U2252 (N_2252,N_2122,N_2016);
or U2253 (N_2253,N_2011,N_2110);
nand U2254 (N_2254,N_2181,N_2029);
nand U2255 (N_2255,N_2114,N_2131);
or U2256 (N_2256,N_2187,N_2166);
and U2257 (N_2257,N_2168,N_2143);
or U2258 (N_2258,N_2159,N_2030);
nor U2259 (N_2259,N_2198,N_2101);
nand U2260 (N_2260,N_2171,N_2087);
and U2261 (N_2261,N_2135,N_2133);
and U2262 (N_2262,N_2044,N_2111);
or U2263 (N_2263,N_2160,N_2079);
nand U2264 (N_2264,N_2042,N_2075);
or U2265 (N_2265,N_2086,N_2136);
nor U2266 (N_2266,N_2018,N_2183);
nand U2267 (N_2267,N_2090,N_2078);
xor U2268 (N_2268,N_2177,N_2049);
and U2269 (N_2269,N_2134,N_2189);
nand U2270 (N_2270,N_2116,N_2068);
or U2271 (N_2271,N_2034,N_2170);
xor U2272 (N_2272,N_2121,N_2023);
or U2273 (N_2273,N_2106,N_2045);
nand U2274 (N_2274,N_2118,N_2188);
or U2275 (N_2275,N_2115,N_2074);
or U2276 (N_2276,N_2003,N_2040);
xnor U2277 (N_2277,N_2022,N_2094);
nand U2278 (N_2278,N_2070,N_2085);
nand U2279 (N_2279,N_2099,N_2158);
and U2280 (N_2280,N_2056,N_2120);
and U2281 (N_2281,N_2149,N_2154);
nor U2282 (N_2282,N_2026,N_2125);
xor U2283 (N_2283,N_2130,N_2180);
nor U2284 (N_2284,N_2191,N_2071);
or U2285 (N_2285,N_2065,N_2150);
or U2286 (N_2286,N_2185,N_2138);
xnor U2287 (N_2287,N_2080,N_2067);
or U2288 (N_2288,N_2037,N_2176);
and U2289 (N_2289,N_2137,N_2140);
nor U2290 (N_2290,N_2141,N_2146);
xnor U2291 (N_2291,N_2025,N_2173);
nor U2292 (N_2292,N_2127,N_2001);
nand U2293 (N_2293,N_2082,N_2157);
nor U2294 (N_2294,N_2032,N_2002);
and U2295 (N_2295,N_2144,N_2081);
xor U2296 (N_2296,N_2035,N_2161);
and U2297 (N_2297,N_2123,N_2038);
nand U2298 (N_2298,N_2182,N_2109);
and U2299 (N_2299,N_2007,N_2097);
xnor U2300 (N_2300,N_2116,N_2006);
or U2301 (N_2301,N_2138,N_2069);
or U2302 (N_2302,N_2199,N_2094);
and U2303 (N_2303,N_2157,N_2168);
nor U2304 (N_2304,N_2121,N_2119);
or U2305 (N_2305,N_2031,N_2002);
xor U2306 (N_2306,N_2075,N_2089);
or U2307 (N_2307,N_2058,N_2172);
or U2308 (N_2308,N_2065,N_2066);
and U2309 (N_2309,N_2160,N_2042);
nor U2310 (N_2310,N_2153,N_2114);
nand U2311 (N_2311,N_2110,N_2149);
or U2312 (N_2312,N_2020,N_2131);
or U2313 (N_2313,N_2018,N_2054);
and U2314 (N_2314,N_2034,N_2181);
and U2315 (N_2315,N_2058,N_2166);
nand U2316 (N_2316,N_2162,N_2026);
nor U2317 (N_2317,N_2081,N_2047);
and U2318 (N_2318,N_2023,N_2092);
nand U2319 (N_2319,N_2146,N_2099);
nand U2320 (N_2320,N_2173,N_2164);
or U2321 (N_2321,N_2129,N_2025);
nand U2322 (N_2322,N_2039,N_2168);
nor U2323 (N_2323,N_2182,N_2158);
nor U2324 (N_2324,N_2166,N_2034);
nand U2325 (N_2325,N_2003,N_2055);
and U2326 (N_2326,N_2029,N_2089);
xnor U2327 (N_2327,N_2015,N_2065);
nor U2328 (N_2328,N_2082,N_2198);
nor U2329 (N_2329,N_2073,N_2078);
or U2330 (N_2330,N_2163,N_2196);
nand U2331 (N_2331,N_2076,N_2058);
nand U2332 (N_2332,N_2074,N_2177);
and U2333 (N_2333,N_2147,N_2015);
nor U2334 (N_2334,N_2104,N_2013);
nor U2335 (N_2335,N_2002,N_2072);
and U2336 (N_2336,N_2051,N_2170);
and U2337 (N_2337,N_2055,N_2108);
and U2338 (N_2338,N_2126,N_2026);
and U2339 (N_2339,N_2181,N_2060);
or U2340 (N_2340,N_2093,N_2194);
xor U2341 (N_2341,N_2168,N_2199);
nand U2342 (N_2342,N_2055,N_2068);
nand U2343 (N_2343,N_2038,N_2071);
nand U2344 (N_2344,N_2196,N_2012);
nand U2345 (N_2345,N_2158,N_2009);
or U2346 (N_2346,N_2106,N_2159);
xor U2347 (N_2347,N_2048,N_2172);
and U2348 (N_2348,N_2041,N_2034);
nand U2349 (N_2349,N_2180,N_2115);
nor U2350 (N_2350,N_2015,N_2150);
and U2351 (N_2351,N_2073,N_2035);
nor U2352 (N_2352,N_2072,N_2118);
and U2353 (N_2353,N_2074,N_2187);
and U2354 (N_2354,N_2121,N_2015);
nand U2355 (N_2355,N_2047,N_2011);
xor U2356 (N_2356,N_2115,N_2187);
or U2357 (N_2357,N_2153,N_2162);
nor U2358 (N_2358,N_2129,N_2020);
or U2359 (N_2359,N_2006,N_2097);
and U2360 (N_2360,N_2165,N_2056);
or U2361 (N_2361,N_2082,N_2134);
xnor U2362 (N_2362,N_2133,N_2054);
or U2363 (N_2363,N_2077,N_2006);
nand U2364 (N_2364,N_2021,N_2085);
nand U2365 (N_2365,N_2018,N_2149);
and U2366 (N_2366,N_2028,N_2033);
nand U2367 (N_2367,N_2094,N_2128);
nand U2368 (N_2368,N_2082,N_2050);
and U2369 (N_2369,N_2030,N_2161);
nor U2370 (N_2370,N_2044,N_2014);
or U2371 (N_2371,N_2153,N_2168);
and U2372 (N_2372,N_2014,N_2141);
or U2373 (N_2373,N_2030,N_2073);
nand U2374 (N_2374,N_2072,N_2043);
and U2375 (N_2375,N_2143,N_2003);
and U2376 (N_2376,N_2172,N_2022);
nand U2377 (N_2377,N_2046,N_2131);
nand U2378 (N_2378,N_2102,N_2068);
and U2379 (N_2379,N_2130,N_2033);
nand U2380 (N_2380,N_2196,N_2106);
nor U2381 (N_2381,N_2015,N_2177);
or U2382 (N_2382,N_2184,N_2003);
and U2383 (N_2383,N_2174,N_2003);
and U2384 (N_2384,N_2144,N_2115);
or U2385 (N_2385,N_2030,N_2052);
nor U2386 (N_2386,N_2087,N_2090);
xor U2387 (N_2387,N_2017,N_2050);
and U2388 (N_2388,N_2183,N_2099);
nor U2389 (N_2389,N_2119,N_2097);
nand U2390 (N_2390,N_2117,N_2005);
nand U2391 (N_2391,N_2188,N_2034);
or U2392 (N_2392,N_2058,N_2167);
xnor U2393 (N_2393,N_2006,N_2108);
nand U2394 (N_2394,N_2163,N_2029);
nand U2395 (N_2395,N_2072,N_2144);
and U2396 (N_2396,N_2091,N_2181);
nand U2397 (N_2397,N_2167,N_2146);
xor U2398 (N_2398,N_2188,N_2068);
nand U2399 (N_2399,N_2099,N_2057);
nor U2400 (N_2400,N_2290,N_2330);
and U2401 (N_2401,N_2349,N_2397);
nand U2402 (N_2402,N_2331,N_2313);
nand U2403 (N_2403,N_2222,N_2283);
or U2404 (N_2404,N_2207,N_2308);
xor U2405 (N_2405,N_2210,N_2260);
nand U2406 (N_2406,N_2277,N_2220);
or U2407 (N_2407,N_2304,N_2205);
or U2408 (N_2408,N_2269,N_2365);
and U2409 (N_2409,N_2390,N_2318);
nor U2410 (N_2410,N_2257,N_2327);
or U2411 (N_2411,N_2340,N_2356);
nor U2412 (N_2412,N_2375,N_2240);
and U2413 (N_2413,N_2353,N_2237);
and U2414 (N_2414,N_2300,N_2326);
or U2415 (N_2415,N_2249,N_2266);
nor U2416 (N_2416,N_2368,N_2263);
or U2417 (N_2417,N_2296,N_2206);
nand U2418 (N_2418,N_2204,N_2273);
nand U2419 (N_2419,N_2264,N_2270);
and U2420 (N_2420,N_2344,N_2218);
xor U2421 (N_2421,N_2208,N_2399);
and U2422 (N_2422,N_2246,N_2377);
and U2423 (N_2423,N_2234,N_2373);
nor U2424 (N_2424,N_2248,N_2236);
nor U2425 (N_2425,N_2374,N_2291);
nand U2426 (N_2426,N_2329,N_2392);
xnor U2427 (N_2427,N_2200,N_2298);
nor U2428 (N_2428,N_2303,N_2201);
xor U2429 (N_2429,N_2345,N_2293);
or U2430 (N_2430,N_2267,N_2226);
or U2431 (N_2431,N_2342,N_2328);
nor U2432 (N_2432,N_2364,N_2287);
and U2433 (N_2433,N_2359,N_2216);
or U2434 (N_2434,N_2350,N_2292);
or U2435 (N_2435,N_2255,N_2295);
nand U2436 (N_2436,N_2280,N_2363);
and U2437 (N_2437,N_2385,N_2332);
xor U2438 (N_2438,N_2317,N_2343);
and U2439 (N_2439,N_2275,N_2341);
xnor U2440 (N_2440,N_2243,N_2379);
nor U2441 (N_2441,N_2235,N_2337);
and U2442 (N_2442,N_2288,N_2241);
nor U2443 (N_2443,N_2217,N_2302);
nor U2444 (N_2444,N_2211,N_2372);
nand U2445 (N_2445,N_2299,N_2225);
and U2446 (N_2446,N_2361,N_2247);
nand U2447 (N_2447,N_2209,N_2360);
nand U2448 (N_2448,N_2378,N_2384);
or U2449 (N_2449,N_2321,N_2314);
nor U2450 (N_2450,N_2219,N_2258);
nor U2451 (N_2451,N_2398,N_2396);
and U2452 (N_2452,N_2347,N_2370);
nand U2453 (N_2453,N_2371,N_2355);
and U2454 (N_2454,N_2366,N_2256);
nand U2455 (N_2455,N_2346,N_2307);
and U2456 (N_2456,N_2339,N_2245);
nor U2457 (N_2457,N_2393,N_2362);
nor U2458 (N_2458,N_2367,N_2212);
nand U2459 (N_2459,N_2272,N_2244);
or U2460 (N_2460,N_2358,N_2271);
or U2461 (N_2461,N_2278,N_2369);
and U2462 (N_2462,N_2315,N_2386);
nor U2463 (N_2463,N_2215,N_2228);
or U2464 (N_2464,N_2253,N_2305);
nand U2465 (N_2465,N_2325,N_2297);
or U2466 (N_2466,N_2352,N_2333);
or U2467 (N_2467,N_2306,N_2282);
xnor U2468 (N_2468,N_2354,N_2261);
nor U2469 (N_2469,N_2281,N_2224);
nand U2470 (N_2470,N_2227,N_2391);
nor U2471 (N_2471,N_2323,N_2250);
nand U2472 (N_2472,N_2229,N_2316);
nand U2473 (N_2473,N_2338,N_2223);
nor U2474 (N_2474,N_2294,N_2262);
or U2475 (N_2475,N_2380,N_2231);
and U2476 (N_2476,N_2289,N_2202);
or U2477 (N_2477,N_2381,N_2251);
or U2478 (N_2478,N_2351,N_2311);
or U2479 (N_2479,N_2312,N_2230);
nor U2480 (N_2480,N_2335,N_2336);
xor U2481 (N_2481,N_2395,N_2238);
and U2482 (N_2482,N_2286,N_2274);
nand U2483 (N_2483,N_2334,N_2221);
nand U2484 (N_2484,N_2265,N_2276);
nand U2485 (N_2485,N_2383,N_2232);
or U2486 (N_2486,N_2239,N_2310);
nor U2487 (N_2487,N_2254,N_2309);
and U2488 (N_2488,N_2319,N_2279);
or U2489 (N_2489,N_2242,N_2214);
nand U2490 (N_2490,N_2382,N_2284);
nand U2491 (N_2491,N_2357,N_2389);
nor U2492 (N_2492,N_2387,N_2252);
nor U2493 (N_2493,N_2233,N_2388);
and U2494 (N_2494,N_2285,N_2394);
nor U2495 (N_2495,N_2268,N_2322);
and U2496 (N_2496,N_2259,N_2320);
nand U2497 (N_2497,N_2301,N_2203);
and U2498 (N_2498,N_2324,N_2376);
and U2499 (N_2499,N_2213,N_2348);
or U2500 (N_2500,N_2220,N_2248);
and U2501 (N_2501,N_2258,N_2337);
nand U2502 (N_2502,N_2282,N_2307);
nor U2503 (N_2503,N_2393,N_2361);
nand U2504 (N_2504,N_2273,N_2266);
and U2505 (N_2505,N_2221,N_2313);
and U2506 (N_2506,N_2294,N_2267);
nand U2507 (N_2507,N_2313,N_2266);
and U2508 (N_2508,N_2273,N_2316);
nand U2509 (N_2509,N_2215,N_2280);
or U2510 (N_2510,N_2397,N_2265);
nand U2511 (N_2511,N_2305,N_2256);
nor U2512 (N_2512,N_2233,N_2339);
nor U2513 (N_2513,N_2262,N_2388);
and U2514 (N_2514,N_2226,N_2234);
or U2515 (N_2515,N_2252,N_2396);
nand U2516 (N_2516,N_2328,N_2242);
nor U2517 (N_2517,N_2298,N_2279);
xnor U2518 (N_2518,N_2226,N_2366);
xnor U2519 (N_2519,N_2256,N_2354);
nand U2520 (N_2520,N_2399,N_2312);
or U2521 (N_2521,N_2325,N_2380);
or U2522 (N_2522,N_2247,N_2232);
nand U2523 (N_2523,N_2350,N_2345);
nand U2524 (N_2524,N_2222,N_2270);
nor U2525 (N_2525,N_2241,N_2352);
or U2526 (N_2526,N_2377,N_2364);
xnor U2527 (N_2527,N_2244,N_2358);
nor U2528 (N_2528,N_2214,N_2329);
nand U2529 (N_2529,N_2249,N_2324);
and U2530 (N_2530,N_2306,N_2393);
or U2531 (N_2531,N_2282,N_2259);
and U2532 (N_2532,N_2335,N_2218);
xor U2533 (N_2533,N_2243,N_2343);
nand U2534 (N_2534,N_2324,N_2374);
or U2535 (N_2535,N_2262,N_2254);
nor U2536 (N_2536,N_2336,N_2368);
or U2537 (N_2537,N_2221,N_2394);
nand U2538 (N_2538,N_2206,N_2278);
nor U2539 (N_2539,N_2225,N_2234);
xor U2540 (N_2540,N_2255,N_2265);
nand U2541 (N_2541,N_2264,N_2283);
xor U2542 (N_2542,N_2357,N_2337);
nand U2543 (N_2543,N_2389,N_2392);
nor U2544 (N_2544,N_2343,N_2388);
and U2545 (N_2545,N_2359,N_2307);
nor U2546 (N_2546,N_2305,N_2206);
nor U2547 (N_2547,N_2348,N_2302);
or U2548 (N_2548,N_2320,N_2385);
and U2549 (N_2549,N_2346,N_2381);
nor U2550 (N_2550,N_2259,N_2305);
and U2551 (N_2551,N_2358,N_2321);
and U2552 (N_2552,N_2342,N_2305);
and U2553 (N_2553,N_2214,N_2259);
nand U2554 (N_2554,N_2399,N_2213);
or U2555 (N_2555,N_2358,N_2324);
or U2556 (N_2556,N_2283,N_2286);
nand U2557 (N_2557,N_2387,N_2280);
nor U2558 (N_2558,N_2269,N_2344);
nand U2559 (N_2559,N_2383,N_2267);
nor U2560 (N_2560,N_2386,N_2247);
or U2561 (N_2561,N_2365,N_2225);
nor U2562 (N_2562,N_2367,N_2225);
or U2563 (N_2563,N_2212,N_2310);
nand U2564 (N_2564,N_2307,N_2397);
nand U2565 (N_2565,N_2270,N_2368);
nand U2566 (N_2566,N_2226,N_2311);
nand U2567 (N_2567,N_2273,N_2396);
nor U2568 (N_2568,N_2392,N_2368);
and U2569 (N_2569,N_2343,N_2380);
nand U2570 (N_2570,N_2318,N_2323);
and U2571 (N_2571,N_2202,N_2218);
and U2572 (N_2572,N_2335,N_2312);
and U2573 (N_2573,N_2336,N_2399);
nand U2574 (N_2574,N_2293,N_2346);
nor U2575 (N_2575,N_2298,N_2325);
and U2576 (N_2576,N_2273,N_2382);
nand U2577 (N_2577,N_2210,N_2304);
and U2578 (N_2578,N_2365,N_2305);
nand U2579 (N_2579,N_2214,N_2240);
xnor U2580 (N_2580,N_2247,N_2284);
or U2581 (N_2581,N_2204,N_2321);
and U2582 (N_2582,N_2249,N_2360);
or U2583 (N_2583,N_2255,N_2396);
xnor U2584 (N_2584,N_2233,N_2208);
nand U2585 (N_2585,N_2245,N_2314);
nor U2586 (N_2586,N_2361,N_2204);
or U2587 (N_2587,N_2319,N_2328);
and U2588 (N_2588,N_2333,N_2234);
or U2589 (N_2589,N_2318,N_2289);
or U2590 (N_2590,N_2351,N_2384);
xnor U2591 (N_2591,N_2222,N_2332);
or U2592 (N_2592,N_2328,N_2389);
nand U2593 (N_2593,N_2359,N_2379);
or U2594 (N_2594,N_2265,N_2339);
or U2595 (N_2595,N_2388,N_2361);
nor U2596 (N_2596,N_2341,N_2354);
nor U2597 (N_2597,N_2251,N_2220);
or U2598 (N_2598,N_2290,N_2214);
and U2599 (N_2599,N_2336,N_2354);
xnor U2600 (N_2600,N_2438,N_2507);
nor U2601 (N_2601,N_2532,N_2582);
nor U2602 (N_2602,N_2501,N_2569);
nand U2603 (N_2603,N_2468,N_2451);
nor U2604 (N_2604,N_2543,N_2425);
nand U2605 (N_2605,N_2594,N_2530);
or U2606 (N_2606,N_2473,N_2573);
nor U2607 (N_2607,N_2457,N_2553);
nand U2608 (N_2608,N_2505,N_2443);
xnor U2609 (N_2609,N_2570,N_2434);
xor U2610 (N_2610,N_2424,N_2470);
or U2611 (N_2611,N_2433,N_2598);
nand U2612 (N_2612,N_2466,N_2493);
and U2613 (N_2613,N_2441,N_2566);
or U2614 (N_2614,N_2583,N_2549);
nor U2615 (N_2615,N_2508,N_2565);
xnor U2616 (N_2616,N_2419,N_2580);
nand U2617 (N_2617,N_2414,N_2528);
and U2618 (N_2618,N_2430,N_2588);
nand U2619 (N_2619,N_2427,N_2435);
nand U2620 (N_2620,N_2579,N_2442);
and U2621 (N_2621,N_2599,N_2568);
nand U2622 (N_2622,N_2411,N_2485);
xor U2623 (N_2623,N_2597,N_2416);
and U2624 (N_2624,N_2546,N_2450);
and U2625 (N_2625,N_2449,N_2480);
nand U2626 (N_2626,N_2403,N_2500);
nand U2627 (N_2627,N_2408,N_2593);
nor U2628 (N_2628,N_2455,N_2524);
and U2629 (N_2629,N_2556,N_2544);
xnor U2630 (N_2630,N_2539,N_2538);
nor U2631 (N_2631,N_2478,N_2542);
and U2632 (N_2632,N_2495,N_2469);
xor U2633 (N_2633,N_2572,N_2558);
nor U2634 (N_2634,N_2577,N_2479);
and U2635 (N_2635,N_2429,N_2477);
or U2636 (N_2636,N_2595,N_2475);
nor U2637 (N_2637,N_2465,N_2482);
and U2638 (N_2638,N_2488,N_2412);
nand U2639 (N_2639,N_2550,N_2422);
or U2640 (N_2640,N_2581,N_2406);
xnor U2641 (N_2641,N_2489,N_2513);
or U2642 (N_2642,N_2520,N_2446);
nand U2643 (N_2643,N_2436,N_2563);
and U2644 (N_2644,N_2592,N_2540);
nor U2645 (N_2645,N_2561,N_2481);
and U2646 (N_2646,N_2452,N_2440);
xnor U2647 (N_2647,N_2491,N_2444);
nor U2648 (N_2648,N_2448,N_2418);
nand U2649 (N_2649,N_2459,N_2576);
and U2650 (N_2650,N_2548,N_2494);
nand U2651 (N_2651,N_2584,N_2511);
and U2652 (N_2652,N_2552,N_2401);
nor U2653 (N_2653,N_2596,N_2555);
and U2654 (N_2654,N_2447,N_2486);
nand U2655 (N_2655,N_2487,N_2562);
or U2656 (N_2656,N_2409,N_2463);
or U2657 (N_2657,N_2510,N_2504);
nor U2658 (N_2658,N_2464,N_2483);
nor U2659 (N_2659,N_2560,N_2490);
nor U2660 (N_2660,N_2506,N_2521);
or U2661 (N_2661,N_2462,N_2502);
or U2662 (N_2662,N_2474,N_2499);
xnor U2663 (N_2663,N_2526,N_2571);
xor U2664 (N_2664,N_2534,N_2535);
or U2665 (N_2665,N_2512,N_2426);
or U2666 (N_2666,N_2590,N_2407);
or U2667 (N_2667,N_2527,N_2589);
or U2668 (N_2668,N_2415,N_2554);
xnor U2669 (N_2669,N_2410,N_2536);
nor U2670 (N_2670,N_2458,N_2472);
nand U2671 (N_2671,N_2456,N_2547);
nand U2672 (N_2672,N_2551,N_2522);
nand U2673 (N_2673,N_2575,N_2585);
or U2674 (N_2674,N_2564,N_2467);
nor U2675 (N_2675,N_2461,N_2454);
or U2676 (N_2676,N_2517,N_2586);
nor U2677 (N_2677,N_2533,N_2417);
or U2678 (N_2678,N_2537,N_2405);
or U2679 (N_2679,N_2439,N_2545);
or U2680 (N_2680,N_2587,N_2503);
nand U2681 (N_2681,N_2428,N_2431);
nand U2682 (N_2682,N_2567,N_2420);
or U2683 (N_2683,N_2529,N_2423);
nor U2684 (N_2684,N_2496,N_2492);
nand U2685 (N_2685,N_2484,N_2531);
xor U2686 (N_2686,N_2578,N_2432);
nand U2687 (N_2687,N_2413,N_2402);
nor U2688 (N_2688,N_2460,N_2525);
nor U2689 (N_2689,N_2421,N_2559);
nand U2690 (N_2690,N_2476,N_2541);
or U2691 (N_2691,N_2514,N_2518);
and U2692 (N_2692,N_2404,N_2498);
nor U2693 (N_2693,N_2471,N_2400);
or U2694 (N_2694,N_2453,N_2591);
xor U2695 (N_2695,N_2445,N_2519);
nand U2696 (N_2696,N_2509,N_2515);
and U2697 (N_2697,N_2516,N_2574);
and U2698 (N_2698,N_2557,N_2497);
nand U2699 (N_2699,N_2437,N_2523);
nor U2700 (N_2700,N_2462,N_2412);
xnor U2701 (N_2701,N_2516,N_2545);
nand U2702 (N_2702,N_2437,N_2548);
or U2703 (N_2703,N_2459,N_2451);
xor U2704 (N_2704,N_2524,N_2508);
nand U2705 (N_2705,N_2596,N_2574);
nand U2706 (N_2706,N_2559,N_2571);
and U2707 (N_2707,N_2432,N_2494);
nand U2708 (N_2708,N_2589,N_2480);
nor U2709 (N_2709,N_2465,N_2531);
nor U2710 (N_2710,N_2456,N_2581);
nor U2711 (N_2711,N_2519,N_2575);
or U2712 (N_2712,N_2464,N_2442);
and U2713 (N_2713,N_2506,N_2543);
or U2714 (N_2714,N_2585,N_2531);
nor U2715 (N_2715,N_2476,N_2558);
nor U2716 (N_2716,N_2422,N_2449);
xnor U2717 (N_2717,N_2435,N_2409);
or U2718 (N_2718,N_2511,N_2462);
xor U2719 (N_2719,N_2524,N_2576);
or U2720 (N_2720,N_2422,N_2423);
nand U2721 (N_2721,N_2547,N_2515);
or U2722 (N_2722,N_2503,N_2598);
nand U2723 (N_2723,N_2429,N_2427);
or U2724 (N_2724,N_2440,N_2432);
nand U2725 (N_2725,N_2527,N_2472);
nor U2726 (N_2726,N_2428,N_2538);
nor U2727 (N_2727,N_2426,N_2454);
nor U2728 (N_2728,N_2462,N_2456);
nand U2729 (N_2729,N_2593,N_2487);
and U2730 (N_2730,N_2443,N_2514);
or U2731 (N_2731,N_2409,N_2565);
and U2732 (N_2732,N_2586,N_2403);
and U2733 (N_2733,N_2526,N_2438);
and U2734 (N_2734,N_2523,N_2580);
and U2735 (N_2735,N_2429,N_2470);
and U2736 (N_2736,N_2508,N_2518);
nor U2737 (N_2737,N_2552,N_2430);
and U2738 (N_2738,N_2419,N_2575);
and U2739 (N_2739,N_2441,N_2426);
nand U2740 (N_2740,N_2437,N_2469);
nand U2741 (N_2741,N_2595,N_2504);
xnor U2742 (N_2742,N_2560,N_2564);
or U2743 (N_2743,N_2428,N_2415);
nor U2744 (N_2744,N_2496,N_2403);
nor U2745 (N_2745,N_2401,N_2569);
nor U2746 (N_2746,N_2528,N_2417);
nor U2747 (N_2747,N_2464,N_2596);
and U2748 (N_2748,N_2424,N_2403);
nand U2749 (N_2749,N_2411,N_2508);
xor U2750 (N_2750,N_2596,N_2452);
and U2751 (N_2751,N_2539,N_2590);
or U2752 (N_2752,N_2571,N_2509);
or U2753 (N_2753,N_2520,N_2596);
nand U2754 (N_2754,N_2511,N_2404);
and U2755 (N_2755,N_2539,N_2471);
xor U2756 (N_2756,N_2538,N_2578);
or U2757 (N_2757,N_2585,N_2456);
nand U2758 (N_2758,N_2557,N_2458);
or U2759 (N_2759,N_2569,N_2498);
nand U2760 (N_2760,N_2458,N_2429);
or U2761 (N_2761,N_2521,N_2525);
nor U2762 (N_2762,N_2583,N_2512);
xnor U2763 (N_2763,N_2443,N_2408);
and U2764 (N_2764,N_2544,N_2448);
nand U2765 (N_2765,N_2427,N_2490);
and U2766 (N_2766,N_2554,N_2555);
nor U2767 (N_2767,N_2517,N_2481);
nand U2768 (N_2768,N_2483,N_2466);
nand U2769 (N_2769,N_2500,N_2462);
nand U2770 (N_2770,N_2475,N_2559);
and U2771 (N_2771,N_2552,N_2420);
nor U2772 (N_2772,N_2510,N_2523);
or U2773 (N_2773,N_2412,N_2451);
nor U2774 (N_2774,N_2596,N_2560);
nor U2775 (N_2775,N_2473,N_2512);
nor U2776 (N_2776,N_2513,N_2505);
nor U2777 (N_2777,N_2575,N_2565);
nor U2778 (N_2778,N_2491,N_2513);
and U2779 (N_2779,N_2584,N_2492);
nor U2780 (N_2780,N_2474,N_2479);
or U2781 (N_2781,N_2509,N_2484);
nor U2782 (N_2782,N_2456,N_2468);
and U2783 (N_2783,N_2551,N_2581);
nand U2784 (N_2784,N_2497,N_2590);
and U2785 (N_2785,N_2512,N_2403);
xnor U2786 (N_2786,N_2568,N_2547);
nand U2787 (N_2787,N_2405,N_2593);
nand U2788 (N_2788,N_2566,N_2461);
nand U2789 (N_2789,N_2439,N_2552);
or U2790 (N_2790,N_2474,N_2573);
or U2791 (N_2791,N_2401,N_2550);
xnor U2792 (N_2792,N_2513,N_2533);
and U2793 (N_2793,N_2440,N_2555);
and U2794 (N_2794,N_2541,N_2420);
and U2795 (N_2795,N_2434,N_2482);
nand U2796 (N_2796,N_2548,N_2404);
nor U2797 (N_2797,N_2507,N_2482);
xnor U2798 (N_2798,N_2494,N_2561);
nor U2799 (N_2799,N_2488,N_2464);
and U2800 (N_2800,N_2796,N_2649);
nand U2801 (N_2801,N_2731,N_2757);
nor U2802 (N_2802,N_2615,N_2738);
nand U2803 (N_2803,N_2620,N_2618);
or U2804 (N_2804,N_2621,N_2631);
nand U2805 (N_2805,N_2634,N_2650);
and U2806 (N_2806,N_2767,N_2775);
nand U2807 (N_2807,N_2698,N_2668);
nand U2808 (N_2808,N_2611,N_2712);
xnor U2809 (N_2809,N_2776,N_2779);
or U2810 (N_2810,N_2659,N_2714);
and U2811 (N_2811,N_2748,N_2743);
and U2812 (N_2812,N_2610,N_2752);
xor U2813 (N_2813,N_2685,N_2740);
nand U2814 (N_2814,N_2773,N_2768);
nand U2815 (N_2815,N_2763,N_2687);
nor U2816 (N_2816,N_2682,N_2706);
nand U2817 (N_2817,N_2730,N_2795);
nor U2818 (N_2818,N_2629,N_2672);
nor U2819 (N_2819,N_2751,N_2747);
or U2820 (N_2820,N_2749,N_2710);
nand U2821 (N_2821,N_2616,N_2742);
and U2822 (N_2822,N_2691,N_2644);
nand U2823 (N_2823,N_2741,N_2703);
nand U2824 (N_2824,N_2626,N_2681);
or U2825 (N_2825,N_2673,N_2732);
and U2826 (N_2826,N_2784,N_2619);
nor U2827 (N_2827,N_2717,N_2766);
and U2828 (N_2828,N_2613,N_2765);
nor U2829 (N_2829,N_2666,N_2771);
nor U2830 (N_2830,N_2720,N_2728);
or U2831 (N_2831,N_2657,N_2725);
xnor U2832 (N_2832,N_2676,N_2762);
or U2833 (N_2833,N_2708,N_2637);
and U2834 (N_2834,N_2652,N_2722);
xnor U2835 (N_2835,N_2697,N_2608);
or U2836 (N_2836,N_2647,N_2716);
and U2837 (N_2837,N_2758,N_2769);
or U2838 (N_2838,N_2683,N_2674);
and U2839 (N_2839,N_2760,N_2684);
nor U2840 (N_2840,N_2656,N_2664);
nand U2841 (N_2841,N_2739,N_2600);
nor U2842 (N_2842,N_2799,N_2635);
or U2843 (N_2843,N_2654,N_2617);
and U2844 (N_2844,N_2721,N_2680);
or U2845 (N_2845,N_2638,N_2701);
nor U2846 (N_2846,N_2797,N_2604);
or U2847 (N_2847,N_2601,N_2783);
nor U2848 (N_2848,N_2753,N_2718);
or U2849 (N_2849,N_2602,N_2792);
and U2850 (N_2850,N_2793,N_2715);
nor U2851 (N_2851,N_2780,N_2606);
and U2852 (N_2852,N_2736,N_2671);
and U2853 (N_2853,N_2678,N_2605);
nand U2854 (N_2854,N_2729,N_2625);
nor U2855 (N_2855,N_2726,N_2607);
nor U2856 (N_2856,N_2632,N_2677);
nand U2857 (N_2857,N_2623,N_2642);
nand U2858 (N_2858,N_2764,N_2707);
xor U2859 (N_2859,N_2778,N_2653);
nand U2860 (N_2860,N_2646,N_2639);
or U2861 (N_2861,N_2786,N_2609);
xnor U2862 (N_2862,N_2648,N_2755);
nor U2863 (N_2863,N_2614,N_2719);
and U2864 (N_2864,N_2737,N_2651);
and U2865 (N_2865,N_2787,N_2643);
nand U2866 (N_2866,N_2688,N_2612);
xor U2867 (N_2867,N_2774,N_2700);
nor U2868 (N_2868,N_2754,N_2794);
nor U2869 (N_2869,N_2696,N_2663);
nor U2870 (N_2870,N_2636,N_2798);
nand U2871 (N_2871,N_2735,N_2624);
and U2872 (N_2872,N_2746,N_2693);
and U2873 (N_2873,N_2675,N_2781);
nand U2874 (N_2874,N_2713,N_2761);
and U2875 (N_2875,N_2689,N_2658);
or U2876 (N_2876,N_2733,N_2744);
and U2877 (N_2877,N_2782,N_2694);
nor U2878 (N_2878,N_2645,N_2690);
and U2879 (N_2879,N_2692,N_2777);
nor U2880 (N_2880,N_2756,N_2723);
nand U2881 (N_2881,N_2695,N_2670);
and U2882 (N_2882,N_2770,N_2750);
nand U2883 (N_2883,N_2791,N_2603);
nor U2884 (N_2884,N_2702,N_2727);
or U2885 (N_2885,N_2655,N_2667);
and U2886 (N_2886,N_2679,N_2711);
or U2887 (N_2887,N_2661,N_2633);
nand U2888 (N_2888,N_2704,N_2686);
nor U2889 (N_2889,N_2745,N_2724);
and U2890 (N_2890,N_2705,N_2660);
nor U2891 (N_2891,N_2699,N_2628);
and U2892 (N_2892,N_2789,N_2785);
nor U2893 (N_2893,N_2669,N_2759);
nor U2894 (N_2894,N_2790,N_2622);
xnor U2895 (N_2895,N_2641,N_2772);
and U2896 (N_2896,N_2734,N_2630);
nand U2897 (N_2897,N_2662,N_2788);
xor U2898 (N_2898,N_2709,N_2627);
or U2899 (N_2899,N_2665,N_2640);
and U2900 (N_2900,N_2762,N_2685);
and U2901 (N_2901,N_2729,N_2605);
xnor U2902 (N_2902,N_2763,N_2652);
nor U2903 (N_2903,N_2692,N_2720);
or U2904 (N_2904,N_2696,N_2745);
and U2905 (N_2905,N_2764,N_2771);
nand U2906 (N_2906,N_2740,N_2751);
nand U2907 (N_2907,N_2707,N_2759);
nor U2908 (N_2908,N_2609,N_2730);
or U2909 (N_2909,N_2762,N_2601);
xnor U2910 (N_2910,N_2628,N_2706);
or U2911 (N_2911,N_2717,N_2705);
nor U2912 (N_2912,N_2667,N_2763);
or U2913 (N_2913,N_2734,N_2635);
nand U2914 (N_2914,N_2624,N_2748);
or U2915 (N_2915,N_2655,N_2689);
or U2916 (N_2916,N_2603,N_2725);
and U2917 (N_2917,N_2760,N_2722);
or U2918 (N_2918,N_2648,N_2698);
nor U2919 (N_2919,N_2689,N_2683);
and U2920 (N_2920,N_2740,N_2621);
and U2921 (N_2921,N_2615,N_2607);
nand U2922 (N_2922,N_2665,N_2600);
or U2923 (N_2923,N_2641,N_2609);
nand U2924 (N_2924,N_2603,N_2712);
nor U2925 (N_2925,N_2663,N_2697);
nor U2926 (N_2926,N_2751,N_2626);
and U2927 (N_2927,N_2687,N_2742);
nor U2928 (N_2928,N_2705,N_2752);
and U2929 (N_2929,N_2664,N_2731);
nor U2930 (N_2930,N_2716,N_2642);
or U2931 (N_2931,N_2799,N_2756);
nor U2932 (N_2932,N_2790,N_2755);
or U2933 (N_2933,N_2633,N_2734);
nand U2934 (N_2934,N_2621,N_2772);
and U2935 (N_2935,N_2691,N_2662);
and U2936 (N_2936,N_2613,N_2641);
and U2937 (N_2937,N_2682,N_2710);
nand U2938 (N_2938,N_2651,N_2611);
xnor U2939 (N_2939,N_2689,N_2648);
or U2940 (N_2940,N_2639,N_2700);
nor U2941 (N_2941,N_2794,N_2610);
nand U2942 (N_2942,N_2609,N_2670);
nor U2943 (N_2943,N_2654,N_2619);
nor U2944 (N_2944,N_2735,N_2699);
and U2945 (N_2945,N_2764,N_2659);
and U2946 (N_2946,N_2727,N_2641);
nand U2947 (N_2947,N_2751,N_2605);
and U2948 (N_2948,N_2691,N_2719);
or U2949 (N_2949,N_2780,N_2797);
xnor U2950 (N_2950,N_2645,N_2733);
or U2951 (N_2951,N_2759,N_2629);
nor U2952 (N_2952,N_2785,N_2624);
or U2953 (N_2953,N_2699,N_2622);
and U2954 (N_2954,N_2664,N_2701);
nand U2955 (N_2955,N_2649,N_2721);
or U2956 (N_2956,N_2707,N_2632);
or U2957 (N_2957,N_2621,N_2617);
or U2958 (N_2958,N_2670,N_2781);
nor U2959 (N_2959,N_2636,N_2621);
xnor U2960 (N_2960,N_2677,N_2742);
or U2961 (N_2961,N_2756,N_2782);
and U2962 (N_2962,N_2766,N_2692);
nor U2963 (N_2963,N_2725,N_2619);
nor U2964 (N_2964,N_2752,N_2692);
and U2965 (N_2965,N_2645,N_2624);
nand U2966 (N_2966,N_2712,N_2663);
nand U2967 (N_2967,N_2633,N_2614);
nand U2968 (N_2968,N_2609,N_2651);
or U2969 (N_2969,N_2774,N_2754);
nand U2970 (N_2970,N_2750,N_2764);
and U2971 (N_2971,N_2707,N_2692);
nand U2972 (N_2972,N_2710,N_2730);
and U2973 (N_2973,N_2722,N_2726);
and U2974 (N_2974,N_2751,N_2614);
xnor U2975 (N_2975,N_2738,N_2705);
nor U2976 (N_2976,N_2601,N_2702);
nor U2977 (N_2977,N_2625,N_2773);
nand U2978 (N_2978,N_2637,N_2736);
nor U2979 (N_2979,N_2724,N_2693);
and U2980 (N_2980,N_2691,N_2772);
and U2981 (N_2981,N_2719,N_2647);
and U2982 (N_2982,N_2769,N_2620);
nor U2983 (N_2983,N_2639,N_2752);
nor U2984 (N_2984,N_2724,N_2668);
and U2985 (N_2985,N_2617,N_2773);
or U2986 (N_2986,N_2654,N_2764);
or U2987 (N_2987,N_2737,N_2726);
or U2988 (N_2988,N_2722,N_2731);
nor U2989 (N_2989,N_2786,N_2615);
or U2990 (N_2990,N_2683,N_2717);
nor U2991 (N_2991,N_2603,N_2600);
nand U2992 (N_2992,N_2781,N_2770);
and U2993 (N_2993,N_2789,N_2660);
nand U2994 (N_2994,N_2714,N_2752);
and U2995 (N_2995,N_2618,N_2782);
xnor U2996 (N_2996,N_2755,N_2704);
xnor U2997 (N_2997,N_2765,N_2630);
or U2998 (N_2998,N_2600,N_2764);
or U2999 (N_2999,N_2720,N_2730);
or U3000 (N_3000,N_2823,N_2805);
nor U3001 (N_3001,N_2835,N_2990);
and U3002 (N_3002,N_2883,N_2846);
or U3003 (N_3003,N_2837,N_2917);
and U3004 (N_3004,N_2953,N_2886);
and U3005 (N_3005,N_2811,N_2919);
nand U3006 (N_3006,N_2803,N_2848);
and U3007 (N_3007,N_2908,N_2885);
nor U3008 (N_3008,N_2854,N_2964);
and U3009 (N_3009,N_2844,N_2926);
and U3010 (N_3010,N_2963,N_2996);
or U3011 (N_3011,N_2954,N_2988);
nand U3012 (N_3012,N_2952,N_2967);
nor U3013 (N_3013,N_2842,N_2915);
nand U3014 (N_3014,N_2891,N_2861);
and U3015 (N_3015,N_2934,N_2874);
xnor U3016 (N_3016,N_2975,N_2950);
and U3017 (N_3017,N_2881,N_2914);
nand U3018 (N_3018,N_2977,N_2984);
nor U3019 (N_3019,N_2997,N_2993);
nor U3020 (N_3020,N_2920,N_2927);
nand U3021 (N_3021,N_2966,N_2860);
nor U3022 (N_3022,N_2804,N_2892);
and U3023 (N_3023,N_2935,N_2956);
nor U3024 (N_3024,N_2822,N_2949);
nor U3025 (N_3025,N_2991,N_2970);
nand U3026 (N_3026,N_2870,N_2928);
nand U3027 (N_3027,N_2900,N_2815);
or U3028 (N_3028,N_2962,N_2916);
and U3029 (N_3029,N_2974,N_2839);
xnor U3030 (N_3030,N_2913,N_2851);
nor U3031 (N_3031,N_2933,N_2901);
and U3032 (N_3032,N_2938,N_2961);
nor U3033 (N_3033,N_2945,N_2955);
nor U3034 (N_3034,N_2878,N_2871);
and U3035 (N_3035,N_2862,N_2931);
and U3036 (N_3036,N_2865,N_2880);
nor U3037 (N_3037,N_2807,N_2976);
nor U3038 (N_3038,N_2906,N_2944);
nor U3039 (N_3039,N_2838,N_2867);
or U3040 (N_3040,N_2922,N_2825);
nor U3041 (N_3041,N_2969,N_2866);
nor U3042 (N_3042,N_2899,N_2951);
nor U3043 (N_3043,N_2818,N_2802);
nor U3044 (N_3044,N_2985,N_2830);
nor U3045 (N_3045,N_2946,N_2882);
or U3046 (N_3046,N_2813,N_2889);
and U3047 (N_3047,N_2849,N_2918);
and U3048 (N_3048,N_2968,N_2986);
nand U3049 (N_3049,N_2869,N_2828);
nor U3050 (N_3050,N_2824,N_2868);
or U3051 (N_3051,N_2832,N_2864);
xor U3052 (N_3052,N_2834,N_2887);
nor U3053 (N_3053,N_2987,N_2929);
nand U3054 (N_3054,N_2841,N_2937);
and U3055 (N_3055,N_2808,N_2924);
and U3056 (N_3056,N_2942,N_2909);
xor U3057 (N_3057,N_2820,N_2912);
and U3058 (N_3058,N_2816,N_2959);
nand U3059 (N_3059,N_2983,N_2859);
nand U3060 (N_3060,N_2814,N_2905);
and U3061 (N_3061,N_2980,N_2806);
nand U3062 (N_3062,N_2957,N_2958);
xor U3063 (N_3063,N_2831,N_2819);
or U3064 (N_3064,N_2890,N_2932);
nor U3065 (N_3065,N_2856,N_2836);
and U3066 (N_3066,N_2877,N_2829);
or U3067 (N_3067,N_2876,N_2873);
and U3068 (N_3068,N_2893,N_2972);
xor U3069 (N_3069,N_2897,N_2872);
nand U3070 (N_3070,N_2939,N_2936);
xor U3071 (N_3071,N_2941,N_2904);
and U3072 (N_3072,N_2810,N_2812);
nand U3073 (N_3073,N_2978,N_2995);
nor U3074 (N_3074,N_2894,N_2884);
nor U3075 (N_3075,N_2847,N_2801);
and U3076 (N_3076,N_2843,N_2960);
xor U3077 (N_3077,N_2895,N_2999);
and U3078 (N_3078,N_2857,N_2947);
or U3079 (N_3079,N_2875,N_2826);
nor U3080 (N_3080,N_2982,N_2940);
and U3081 (N_3081,N_2923,N_2992);
nand U3082 (N_3082,N_2800,N_2948);
nor U3083 (N_3083,N_2821,N_2853);
nor U3084 (N_3084,N_2817,N_2898);
and U3085 (N_3085,N_2907,N_2902);
nand U3086 (N_3086,N_2998,N_2971);
nand U3087 (N_3087,N_2903,N_2855);
xnor U3088 (N_3088,N_2852,N_2911);
nand U3089 (N_3089,N_2827,N_2809);
or U3090 (N_3090,N_2943,N_2979);
or U3091 (N_3091,N_2863,N_2973);
xor U3092 (N_3092,N_2833,N_2845);
and U3093 (N_3093,N_2930,N_2981);
and U3094 (N_3094,N_2840,N_2888);
nand U3095 (N_3095,N_2910,N_2896);
or U3096 (N_3096,N_2850,N_2879);
or U3097 (N_3097,N_2989,N_2921);
nand U3098 (N_3098,N_2858,N_2965);
and U3099 (N_3099,N_2994,N_2925);
and U3100 (N_3100,N_2916,N_2988);
and U3101 (N_3101,N_2872,N_2986);
and U3102 (N_3102,N_2850,N_2838);
and U3103 (N_3103,N_2886,N_2902);
and U3104 (N_3104,N_2938,N_2927);
nand U3105 (N_3105,N_2863,N_2982);
or U3106 (N_3106,N_2844,N_2870);
or U3107 (N_3107,N_2825,N_2819);
nand U3108 (N_3108,N_2885,N_2805);
xor U3109 (N_3109,N_2838,N_2861);
xor U3110 (N_3110,N_2941,N_2817);
nand U3111 (N_3111,N_2862,N_2869);
and U3112 (N_3112,N_2861,N_2856);
or U3113 (N_3113,N_2870,N_2956);
or U3114 (N_3114,N_2878,N_2893);
and U3115 (N_3115,N_2896,N_2972);
xor U3116 (N_3116,N_2832,N_2829);
and U3117 (N_3117,N_2897,N_2977);
or U3118 (N_3118,N_2986,N_2887);
nor U3119 (N_3119,N_2962,N_2857);
and U3120 (N_3120,N_2855,N_2993);
or U3121 (N_3121,N_2944,N_2810);
or U3122 (N_3122,N_2838,N_2988);
nor U3123 (N_3123,N_2864,N_2964);
nor U3124 (N_3124,N_2976,N_2984);
nor U3125 (N_3125,N_2850,N_2925);
or U3126 (N_3126,N_2914,N_2888);
nor U3127 (N_3127,N_2995,N_2937);
nand U3128 (N_3128,N_2847,N_2911);
or U3129 (N_3129,N_2894,N_2915);
nor U3130 (N_3130,N_2902,N_2819);
nor U3131 (N_3131,N_2965,N_2944);
nand U3132 (N_3132,N_2909,N_2893);
xor U3133 (N_3133,N_2862,N_2913);
and U3134 (N_3134,N_2859,N_2815);
nand U3135 (N_3135,N_2954,N_2979);
xnor U3136 (N_3136,N_2907,N_2837);
or U3137 (N_3137,N_2942,N_2954);
xor U3138 (N_3138,N_2846,N_2808);
and U3139 (N_3139,N_2950,N_2873);
or U3140 (N_3140,N_2929,N_2984);
nand U3141 (N_3141,N_2903,N_2960);
or U3142 (N_3142,N_2867,N_2965);
nor U3143 (N_3143,N_2804,N_2926);
or U3144 (N_3144,N_2942,N_2989);
or U3145 (N_3145,N_2932,N_2810);
nor U3146 (N_3146,N_2936,N_2804);
or U3147 (N_3147,N_2827,N_2911);
nand U3148 (N_3148,N_2977,N_2930);
nand U3149 (N_3149,N_2853,N_2949);
nor U3150 (N_3150,N_2933,N_2939);
nor U3151 (N_3151,N_2975,N_2974);
or U3152 (N_3152,N_2996,N_2991);
and U3153 (N_3153,N_2909,N_2948);
xnor U3154 (N_3154,N_2844,N_2986);
and U3155 (N_3155,N_2818,N_2803);
or U3156 (N_3156,N_2976,N_2839);
nor U3157 (N_3157,N_2913,N_2949);
nor U3158 (N_3158,N_2860,N_2956);
and U3159 (N_3159,N_2957,N_2886);
and U3160 (N_3160,N_2848,N_2975);
or U3161 (N_3161,N_2973,N_2926);
or U3162 (N_3162,N_2901,N_2803);
and U3163 (N_3163,N_2979,N_2813);
nor U3164 (N_3164,N_2861,N_2839);
nand U3165 (N_3165,N_2818,N_2916);
nand U3166 (N_3166,N_2986,N_2851);
and U3167 (N_3167,N_2816,N_2923);
nand U3168 (N_3168,N_2855,N_2859);
and U3169 (N_3169,N_2823,N_2916);
or U3170 (N_3170,N_2852,N_2924);
nand U3171 (N_3171,N_2836,N_2999);
nand U3172 (N_3172,N_2831,N_2931);
xor U3173 (N_3173,N_2870,N_2863);
nor U3174 (N_3174,N_2973,N_2840);
and U3175 (N_3175,N_2806,N_2862);
nand U3176 (N_3176,N_2827,N_2995);
and U3177 (N_3177,N_2918,N_2995);
and U3178 (N_3178,N_2952,N_2824);
nor U3179 (N_3179,N_2879,N_2842);
nand U3180 (N_3180,N_2850,N_2962);
nand U3181 (N_3181,N_2873,N_2988);
nor U3182 (N_3182,N_2874,N_2892);
xnor U3183 (N_3183,N_2886,N_2952);
nor U3184 (N_3184,N_2962,N_2987);
or U3185 (N_3185,N_2845,N_2916);
or U3186 (N_3186,N_2900,N_2990);
xor U3187 (N_3187,N_2897,N_2856);
nand U3188 (N_3188,N_2995,N_2852);
or U3189 (N_3189,N_2970,N_2851);
nor U3190 (N_3190,N_2972,N_2927);
nor U3191 (N_3191,N_2857,N_2996);
nor U3192 (N_3192,N_2855,N_2973);
nor U3193 (N_3193,N_2912,N_2953);
xor U3194 (N_3194,N_2992,N_2968);
nand U3195 (N_3195,N_2992,N_2940);
and U3196 (N_3196,N_2819,N_2946);
and U3197 (N_3197,N_2950,N_2958);
nor U3198 (N_3198,N_2888,N_2996);
and U3199 (N_3199,N_2900,N_2851);
xnor U3200 (N_3200,N_3172,N_3034);
nor U3201 (N_3201,N_3111,N_3165);
nor U3202 (N_3202,N_3198,N_3013);
nand U3203 (N_3203,N_3050,N_3178);
nor U3204 (N_3204,N_3011,N_3115);
or U3205 (N_3205,N_3098,N_3109);
and U3206 (N_3206,N_3191,N_3048);
nor U3207 (N_3207,N_3058,N_3009);
or U3208 (N_3208,N_3040,N_3148);
or U3209 (N_3209,N_3061,N_3126);
xnor U3210 (N_3210,N_3072,N_3157);
nor U3211 (N_3211,N_3195,N_3056);
and U3212 (N_3212,N_3146,N_3010);
and U3213 (N_3213,N_3099,N_3085);
or U3214 (N_3214,N_3192,N_3140);
nor U3215 (N_3215,N_3182,N_3166);
and U3216 (N_3216,N_3156,N_3064);
and U3217 (N_3217,N_3110,N_3149);
or U3218 (N_3218,N_3093,N_3119);
and U3219 (N_3219,N_3167,N_3032);
nor U3220 (N_3220,N_3043,N_3152);
nand U3221 (N_3221,N_3068,N_3047);
or U3222 (N_3222,N_3125,N_3012);
nand U3223 (N_3223,N_3090,N_3150);
and U3224 (N_3224,N_3071,N_3184);
nor U3225 (N_3225,N_3174,N_3170);
and U3226 (N_3226,N_3031,N_3075);
nand U3227 (N_3227,N_3024,N_3091);
or U3228 (N_3228,N_3015,N_3067);
or U3229 (N_3229,N_3089,N_3036);
and U3230 (N_3230,N_3168,N_3066);
and U3231 (N_3231,N_3122,N_3073);
or U3232 (N_3232,N_3005,N_3100);
xnor U3233 (N_3233,N_3028,N_3135);
nand U3234 (N_3234,N_3095,N_3147);
xnor U3235 (N_3235,N_3088,N_3196);
nand U3236 (N_3236,N_3180,N_3059);
or U3237 (N_3237,N_3092,N_3141);
or U3238 (N_3238,N_3051,N_3133);
and U3239 (N_3239,N_3083,N_3124);
and U3240 (N_3240,N_3029,N_3153);
or U3241 (N_3241,N_3118,N_3128);
nand U3242 (N_3242,N_3103,N_3132);
nand U3243 (N_3243,N_3094,N_3155);
or U3244 (N_3244,N_3022,N_3181);
nor U3245 (N_3245,N_3096,N_3004);
nand U3246 (N_3246,N_3069,N_3020);
and U3247 (N_3247,N_3016,N_3163);
or U3248 (N_3248,N_3079,N_3164);
and U3249 (N_3249,N_3074,N_3065);
nand U3250 (N_3250,N_3023,N_3038);
nand U3251 (N_3251,N_3042,N_3199);
xor U3252 (N_3252,N_3021,N_3188);
or U3253 (N_3253,N_3120,N_3113);
nor U3254 (N_3254,N_3101,N_3002);
and U3255 (N_3255,N_3026,N_3112);
nor U3256 (N_3256,N_3078,N_3117);
and U3257 (N_3257,N_3003,N_3070);
and U3258 (N_3258,N_3000,N_3169);
xor U3259 (N_3259,N_3197,N_3076);
or U3260 (N_3260,N_3045,N_3171);
or U3261 (N_3261,N_3097,N_3080);
nand U3262 (N_3262,N_3054,N_3130);
nand U3263 (N_3263,N_3162,N_3131);
or U3264 (N_3264,N_3173,N_3137);
nor U3265 (N_3265,N_3055,N_3134);
and U3266 (N_3266,N_3186,N_3087);
nand U3267 (N_3267,N_3121,N_3189);
nand U3268 (N_3268,N_3030,N_3107);
or U3269 (N_3269,N_3060,N_3114);
or U3270 (N_3270,N_3193,N_3136);
or U3271 (N_3271,N_3006,N_3063);
or U3272 (N_3272,N_3175,N_3102);
and U3273 (N_3273,N_3052,N_3187);
and U3274 (N_3274,N_3129,N_3144);
nand U3275 (N_3275,N_3154,N_3033);
or U3276 (N_3276,N_3084,N_3108);
nand U3277 (N_3277,N_3046,N_3106);
nor U3278 (N_3278,N_3158,N_3159);
nand U3279 (N_3279,N_3185,N_3027);
nor U3280 (N_3280,N_3086,N_3044);
and U3281 (N_3281,N_3142,N_3019);
nor U3282 (N_3282,N_3053,N_3105);
and U3283 (N_3283,N_3062,N_3057);
and U3284 (N_3284,N_3041,N_3183);
nor U3285 (N_3285,N_3160,N_3025);
or U3286 (N_3286,N_3081,N_3104);
and U3287 (N_3287,N_3179,N_3161);
nor U3288 (N_3288,N_3037,N_3035);
nand U3289 (N_3289,N_3008,N_3138);
nor U3290 (N_3290,N_3001,N_3116);
nor U3291 (N_3291,N_3123,N_3194);
nor U3292 (N_3292,N_3139,N_3176);
nand U3293 (N_3293,N_3007,N_3049);
and U3294 (N_3294,N_3127,N_3014);
or U3295 (N_3295,N_3177,N_3190);
nand U3296 (N_3296,N_3143,N_3077);
and U3297 (N_3297,N_3039,N_3082);
and U3298 (N_3298,N_3017,N_3151);
nor U3299 (N_3299,N_3018,N_3145);
or U3300 (N_3300,N_3081,N_3098);
or U3301 (N_3301,N_3076,N_3168);
and U3302 (N_3302,N_3107,N_3130);
nand U3303 (N_3303,N_3195,N_3188);
or U3304 (N_3304,N_3062,N_3004);
and U3305 (N_3305,N_3025,N_3152);
nor U3306 (N_3306,N_3197,N_3143);
nor U3307 (N_3307,N_3167,N_3184);
and U3308 (N_3308,N_3006,N_3071);
and U3309 (N_3309,N_3176,N_3026);
and U3310 (N_3310,N_3138,N_3129);
nor U3311 (N_3311,N_3077,N_3052);
and U3312 (N_3312,N_3181,N_3033);
nand U3313 (N_3313,N_3117,N_3130);
nor U3314 (N_3314,N_3041,N_3179);
xnor U3315 (N_3315,N_3059,N_3025);
and U3316 (N_3316,N_3099,N_3142);
nand U3317 (N_3317,N_3119,N_3044);
nand U3318 (N_3318,N_3148,N_3069);
nand U3319 (N_3319,N_3061,N_3088);
nor U3320 (N_3320,N_3015,N_3135);
xor U3321 (N_3321,N_3158,N_3048);
and U3322 (N_3322,N_3039,N_3049);
or U3323 (N_3323,N_3151,N_3199);
nor U3324 (N_3324,N_3071,N_3187);
or U3325 (N_3325,N_3189,N_3034);
nor U3326 (N_3326,N_3171,N_3141);
or U3327 (N_3327,N_3052,N_3015);
or U3328 (N_3328,N_3181,N_3152);
nand U3329 (N_3329,N_3094,N_3105);
nand U3330 (N_3330,N_3135,N_3009);
and U3331 (N_3331,N_3191,N_3139);
nor U3332 (N_3332,N_3140,N_3033);
or U3333 (N_3333,N_3094,N_3096);
and U3334 (N_3334,N_3042,N_3016);
nor U3335 (N_3335,N_3041,N_3126);
xnor U3336 (N_3336,N_3040,N_3103);
and U3337 (N_3337,N_3032,N_3040);
xor U3338 (N_3338,N_3048,N_3188);
nand U3339 (N_3339,N_3026,N_3013);
or U3340 (N_3340,N_3002,N_3165);
and U3341 (N_3341,N_3131,N_3120);
nand U3342 (N_3342,N_3140,N_3170);
nand U3343 (N_3343,N_3008,N_3061);
nor U3344 (N_3344,N_3151,N_3148);
nand U3345 (N_3345,N_3009,N_3044);
and U3346 (N_3346,N_3198,N_3094);
or U3347 (N_3347,N_3055,N_3159);
nand U3348 (N_3348,N_3169,N_3124);
or U3349 (N_3349,N_3036,N_3003);
nor U3350 (N_3350,N_3112,N_3129);
and U3351 (N_3351,N_3027,N_3090);
nand U3352 (N_3352,N_3034,N_3100);
xor U3353 (N_3353,N_3178,N_3016);
or U3354 (N_3354,N_3005,N_3185);
and U3355 (N_3355,N_3094,N_3059);
and U3356 (N_3356,N_3098,N_3159);
nor U3357 (N_3357,N_3044,N_3091);
nand U3358 (N_3358,N_3069,N_3089);
nor U3359 (N_3359,N_3124,N_3050);
and U3360 (N_3360,N_3065,N_3133);
xnor U3361 (N_3361,N_3155,N_3139);
xnor U3362 (N_3362,N_3157,N_3070);
and U3363 (N_3363,N_3136,N_3179);
nand U3364 (N_3364,N_3041,N_3077);
nand U3365 (N_3365,N_3094,N_3029);
or U3366 (N_3366,N_3042,N_3158);
or U3367 (N_3367,N_3190,N_3182);
nand U3368 (N_3368,N_3065,N_3004);
nand U3369 (N_3369,N_3086,N_3091);
or U3370 (N_3370,N_3079,N_3006);
xor U3371 (N_3371,N_3049,N_3005);
nor U3372 (N_3372,N_3147,N_3055);
nor U3373 (N_3373,N_3002,N_3162);
nand U3374 (N_3374,N_3135,N_3012);
nor U3375 (N_3375,N_3003,N_3154);
nor U3376 (N_3376,N_3183,N_3150);
xnor U3377 (N_3377,N_3108,N_3167);
or U3378 (N_3378,N_3075,N_3183);
and U3379 (N_3379,N_3179,N_3165);
and U3380 (N_3380,N_3157,N_3074);
nor U3381 (N_3381,N_3124,N_3187);
xor U3382 (N_3382,N_3179,N_3172);
and U3383 (N_3383,N_3099,N_3048);
xor U3384 (N_3384,N_3131,N_3155);
nor U3385 (N_3385,N_3057,N_3021);
nand U3386 (N_3386,N_3033,N_3187);
nor U3387 (N_3387,N_3104,N_3118);
and U3388 (N_3388,N_3043,N_3192);
and U3389 (N_3389,N_3165,N_3008);
and U3390 (N_3390,N_3084,N_3100);
nand U3391 (N_3391,N_3089,N_3128);
and U3392 (N_3392,N_3064,N_3138);
and U3393 (N_3393,N_3070,N_3014);
nand U3394 (N_3394,N_3037,N_3011);
or U3395 (N_3395,N_3034,N_3060);
nor U3396 (N_3396,N_3037,N_3185);
and U3397 (N_3397,N_3036,N_3171);
xnor U3398 (N_3398,N_3120,N_3016);
xor U3399 (N_3399,N_3132,N_3151);
and U3400 (N_3400,N_3349,N_3376);
or U3401 (N_3401,N_3285,N_3244);
or U3402 (N_3402,N_3364,N_3211);
nor U3403 (N_3403,N_3226,N_3321);
nor U3404 (N_3404,N_3287,N_3350);
or U3405 (N_3405,N_3311,N_3390);
nor U3406 (N_3406,N_3227,N_3373);
and U3407 (N_3407,N_3240,N_3296);
and U3408 (N_3408,N_3222,N_3213);
nand U3409 (N_3409,N_3223,N_3243);
or U3410 (N_3410,N_3308,N_3345);
nand U3411 (N_3411,N_3314,N_3295);
or U3412 (N_3412,N_3256,N_3306);
nand U3413 (N_3413,N_3216,N_3327);
nor U3414 (N_3414,N_3207,N_3262);
nor U3415 (N_3415,N_3247,N_3333);
nor U3416 (N_3416,N_3309,N_3371);
nor U3417 (N_3417,N_3369,N_3331);
xor U3418 (N_3418,N_3312,N_3206);
nor U3419 (N_3419,N_3283,N_3250);
nand U3420 (N_3420,N_3377,N_3200);
or U3421 (N_3421,N_3361,N_3355);
nor U3422 (N_3422,N_3375,N_3284);
nor U3423 (N_3423,N_3342,N_3265);
and U3424 (N_3424,N_3278,N_3334);
nor U3425 (N_3425,N_3394,N_3238);
nor U3426 (N_3426,N_3239,N_3292);
or U3427 (N_3427,N_3365,N_3270);
nor U3428 (N_3428,N_3391,N_3362);
or U3429 (N_3429,N_3347,N_3228);
and U3430 (N_3430,N_3358,N_3305);
nor U3431 (N_3431,N_3225,N_3298);
nor U3432 (N_3432,N_3388,N_3279);
and U3433 (N_3433,N_3242,N_3351);
nand U3434 (N_3434,N_3263,N_3387);
and U3435 (N_3435,N_3363,N_3352);
and U3436 (N_3436,N_3268,N_3325);
or U3437 (N_3437,N_3368,N_3360);
or U3438 (N_3438,N_3232,N_3335);
and U3439 (N_3439,N_3251,N_3230);
nand U3440 (N_3440,N_3380,N_3217);
and U3441 (N_3441,N_3307,N_3348);
and U3442 (N_3442,N_3214,N_3304);
or U3443 (N_3443,N_3288,N_3259);
nor U3444 (N_3444,N_3276,N_3337);
nand U3445 (N_3445,N_3385,N_3316);
nor U3446 (N_3446,N_3356,N_3392);
nand U3447 (N_3447,N_3313,N_3264);
nand U3448 (N_3448,N_3303,N_3341);
xor U3449 (N_3449,N_3282,N_3310);
and U3450 (N_3450,N_3281,N_3249);
or U3451 (N_3451,N_3220,N_3389);
xnor U3452 (N_3452,N_3209,N_3398);
or U3453 (N_3453,N_3353,N_3234);
nor U3454 (N_3454,N_3378,N_3383);
xnor U3455 (N_3455,N_3324,N_3267);
nor U3456 (N_3456,N_3202,N_3332);
or U3457 (N_3457,N_3315,N_3293);
and U3458 (N_3458,N_3374,N_3215);
xor U3459 (N_3459,N_3253,N_3260);
or U3460 (N_3460,N_3255,N_3326);
nand U3461 (N_3461,N_3218,N_3396);
or U3462 (N_3462,N_3329,N_3271);
xnor U3463 (N_3463,N_3367,N_3302);
nor U3464 (N_3464,N_3366,N_3246);
nor U3465 (N_3465,N_3343,N_3346);
nand U3466 (N_3466,N_3294,N_3340);
xor U3467 (N_3467,N_3274,N_3272);
xor U3468 (N_3468,N_3208,N_3245);
xor U3469 (N_3469,N_3338,N_3275);
and U3470 (N_3470,N_3339,N_3258);
and U3471 (N_3471,N_3317,N_3322);
or U3472 (N_3472,N_3205,N_3229);
and U3473 (N_3473,N_3203,N_3235);
and U3474 (N_3474,N_3384,N_3241);
nor U3475 (N_3475,N_3289,N_3393);
and U3476 (N_3476,N_3233,N_3397);
nor U3477 (N_3477,N_3237,N_3204);
and U3478 (N_3478,N_3254,N_3359);
nor U3479 (N_3479,N_3219,N_3210);
and U3480 (N_3480,N_3286,N_3212);
nand U3481 (N_3481,N_3299,N_3330);
and U3482 (N_3482,N_3323,N_3297);
nand U3483 (N_3483,N_3291,N_3382);
nand U3484 (N_3484,N_3252,N_3320);
nand U3485 (N_3485,N_3221,N_3319);
or U3486 (N_3486,N_3300,N_3301);
or U3487 (N_3487,N_3261,N_3224);
or U3488 (N_3488,N_3370,N_3266);
or U3489 (N_3489,N_3395,N_3236);
nor U3490 (N_3490,N_3248,N_3290);
nand U3491 (N_3491,N_3328,N_3357);
xnor U3492 (N_3492,N_3280,N_3231);
and U3493 (N_3493,N_3257,N_3269);
nor U3494 (N_3494,N_3318,N_3372);
xor U3495 (N_3495,N_3344,N_3336);
and U3496 (N_3496,N_3386,N_3277);
nand U3497 (N_3497,N_3354,N_3201);
and U3498 (N_3498,N_3399,N_3381);
nand U3499 (N_3499,N_3273,N_3379);
nand U3500 (N_3500,N_3204,N_3267);
nand U3501 (N_3501,N_3344,N_3393);
nor U3502 (N_3502,N_3290,N_3220);
or U3503 (N_3503,N_3389,N_3350);
nand U3504 (N_3504,N_3223,N_3308);
or U3505 (N_3505,N_3382,N_3395);
nand U3506 (N_3506,N_3320,N_3394);
xnor U3507 (N_3507,N_3208,N_3379);
nand U3508 (N_3508,N_3338,N_3253);
and U3509 (N_3509,N_3203,N_3255);
and U3510 (N_3510,N_3264,N_3352);
nand U3511 (N_3511,N_3246,N_3356);
or U3512 (N_3512,N_3398,N_3292);
nand U3513 (N_3513,N_3294,N_3369);
nand U3514 (N_3514,N_3220,N_3323);
nand U3515 (N_3515,N_3206,N_3317);
nor U3516 (N_3516,N_3291,N_3241);
and U3517 (N_3517,N_3294,N_3287);
xor U3518 (N_3518,N_3220,N_3279);
xor U3519 (N_3519,N_3260,N_3342);
nand U3520 (N_3520,N_3209,N_3321);
nand U3521 (N_3521,N_3359,N_3351);
nor U3522 (N_3522,N_3292,N_3382);
nor U3523 (N_3523,N_3303,N_3274);
and U3524 (N_3524,N_3222,N_3353);
nand U3525 (N_3525,N_3237,N_3289);
and U3526 (N_3526,N_3252,N_3340);
and U3527 (N_3527,N_3396,N_3226);
and U3528 (N_3528,N_3352,N_3242);
or U3529 (N_3529,N_3381,N_3289);
or U3530 (N_3530,N_3384,N_3367);
and U3531 (N_3531,N_3256,N_3361);
xnor U3532 (N_3532,N_3340,N_3315);
and U3533 (N_3533,N_3345,N_3357);
and U3534 (N_3534,N_3272,N_3339);
or U3535 (N_3535,N_3388,N_3311);
nand U3536 (N_3536,N_3222,N_3380);
and U3537 (N_3537,N_3204,N_3276);
and U3538 (N_3538,N_3333,N_3246);
nand U3539 (N_3539,N_3299,N_3393);
and U3540 (N_3540,N_3285,N_3364);
nand U3541 (N_3541,N_3253,N_3395);
xnor U3542 (N_3542,N_3334,N_3210);
and U3543 (N_3543,N_3230,N_3267);
or U3544 (N_3544,N_3228,N_3289);
and U3545 (N_3545,N_3244,N_3328);
nand U3546 (N_3546,N_3341,N_3338);
nor U3547 (N_3547,N_3219,N_3355);
or U3548 (N_3548,N_3354,N_3212);
nand U3549 (N_3549,N_3227,N_3319);
nand U3550 (N_3550,N_3336,N_3386);
nor U3551 (N_3551,N_3235,N_3257);
nor U3552 (N_3552,N_3249,N_3303);
and U3553 (N_3553,N_3343,N_3202);
and U3554 (N_3554,N_3357,N_3351);
xor U3555 (N_3555,N_3258,N_3381);
nand U3556 (N_3556,N_3204,N_3366);
nand U3557 (N_3557,N_3208,N_3263);
or U3558 (N_3558,N_3251,N_3222);
or U3559 (N_3559,N_3265,N_3260);
nand U3560 (N_3560,N_3258,N_3296);
nand U3561 (N_3561,N_3332,N_3364);
nand U3562 (N_3562,N_3334,N_3245);
nand U3563 (N_3563,N_3259,N_3375);
nand U3564 (N_3564,N_3234,N_3270);
and U3565 (N_3565,N_3262,N_3339);
nand U3566 (N_3566,N_3351,N_3220);
nand U3567 (N_3567,N_3385,N_3282);
and U3568 (N_3568,N_3210,N_3369);
and U3569 (N_3569,N_3267,N_3272);
nor U3570 (N_3570,N_3297,N_3308);
nor U3571 (N_3571,N_3293,N_3341);
and U3572 (N_3572,N_3341,N_3379);
and U3573 (N_3573,N_3302,N_3289);
nor U3574 (N_3574,N_3383,N_3291);
nor U3575 (N_3575,N_3276,N_3226);
nand U3576 (N_3576,N_3358,N_3213);
nand U3577 (N_3577,N_3346,N_3344);
nand U3578 (N_3578,N_3246,N_3279);
nand U3579 (N_3579,N_3215,N_3322);
or U3580 (N_3580,N_3303,N_3206);
or U3581 (N_3581,N_3219,N_3299);
and U3582 (N_3582,N_3300,N_3279);
nand U3583 (N_3583,N_3255,N_3220);
and U3584 (N_3584,N_3247,N_3223);
nor U3585 (N_3585,N_3202,N_3372);
xnor U3586 (N_3586,N_3220,N_3207);
or U3587 (N_3587,N_3388,N_3211);
nor U3588 (N_3588,N_3261,N_3363);
and U3589 (N_3589,N_3255,N_3376);
nor U3590 (N_3590,N_3225,N_3237);
nor U3591 (N_3591,N_3238,N_3321);
nand U3592 (N_3592,N_3261,N_3294);
xor U3593 (N_3593,N_3360,N_3349);
xor U3594 (N_3594,N_3350,N_3275);
nand U3595 (N_3595,N_3331,N_3230);
and U3596 (N_3596,N_3358,N_3373);
nand U3597 (N_3597,N_3223,N_3250);
nor U3598 (N_3598,N_3305,N_3391);
nand U3599 (N_3599,N_3245,N_3236);
and U3600 (N_3600,N_3545,N_3579);
nand U3601 (N_3601,N_3598,N_3462);
or U3602 (N_3602,N_3552,N_3493);
and U3603 (N_3603,N_3433,N_3408);
nor U3604 (N_3604,N_3485,N_3540);
nor U3605 (N_3605,N_3528,N_3582);
nand U3606 (N_3606,N_3599,N_3498);
or U3607 (N_3607,N_3567,N_3430);
nor U3608 (N_3608,N_3595,N_3483);
nand U3609 (N_3609,N_3526,N_3541);
nand U3610 (N_3610,N_3401,N_3409);
or U3611 (N_3611,N_3469,N_3536);
or U3612 (N_3612,N_3417,N_3527);
nor U3613 (N_3613,N_3578,N_3491);
nand U3614 (N_3614,N_3407,N_3502);
and U3615 (N_3615,N_3454,N_3476);
nand U3616 (N_3616,N_3439,N_3431);
nand U3617 (N_3617,N_3500,N_3412);
nor U3618 (N_3618,N_3529,N_3486);
nor U3619 (N_3619,N_3435,N_3563);
and U3620 (N_3620,N_3413,N_3560);
nand U3621 (N_3621,N_3518,N_3474);
xnor U3622 (N_3622,N_3496,N_3591);
xor U3623 (N_3623,N_3434,N_3423);
and U3624 (N_3624,N_3586,N_3447);
nor U3625 (N_3625,N_3571,N_3521);
nor U3626 (N_3626,N_3451,N_3425);
nand U3627 (N_3627,N_3555,N_3585);
nor U3628 (N_3628,N_3534,N_3446);
nor U3629 (N_3629,N_3482,N_3458);
and U3630 (N_3630,N_3584,N_3488);
and U3631 (N_3631,N_3468,N_3480);
or U3632 (N_3632,N_3524,N_3597);
and U3633 (N_3633,N_3479,N_3547);
and U3634 (N_3634,N_3514,N_3421);
nand U3635 (N_3635,N_3569,N_3470);
and U3636 (N_3636,N_3539,N_3420);
xnor U3637 (N_3637,N_3410,N_3424);
nand U3638 (N_3638,N_3588,N_3465);
nand U3639 (N_3639,N_3592,N_3506);
or U3640 (N_3640,N_3453,N_3419);
and U3641 (N_3641,N_3472,N_3583);
nand U3642 (N_3642,N_3437,N_3531);
and U3643 (N_3643,N_3427,N_3554);
xnor U3644 (N_3644,N_3556,N_3492);
and U3645 (N_3645,N_3415,N_3487);
or U3646 (N_3646,N_3504,N_3450);
or U3647 (N_3647,N_3484,N_3573);
xor U3648 (N_3648,N_3537,N_3444);
or U3649 (N_3649,N_3510,N_3495);
and U3650 (N_3650,N_3519,N_3463);
xnor U3651 (N_3651,N_3575,N_3516);
nor U3652 (N_3652,N_3473,N_3589);
nand U3653 (N_3653,N_3576,N_3557);
nand U3654 (N_3654,N_3549,N_3402);
or U3655 (N_3655,N_3490,N_3406);
xnor U3656 (N_3656,N_3416,N_3455);
nand U3657 (N_3657,N_3544,N_3565);
or U3658 (N_3658,N_3561,N_3497);
and U3659 (N_3659,N_3440,N_3543);
nand U3660 (N_3660,N_3511,N_3559);
nor U3661 (N_3661,N_3580,N_3509);
or U3662 (N_3662,N_3457,N_3570);
nand U3663 (N_3663,N_3404,N_3452);
and U3664 (N_3664,N_3553,N_3535);
or U3665 (N_3665,N_3525,N_3577);
xnor U3666 (N_3666,N_3477,N_3596);
xnor U3667 (N_3667,N_3558,N_3581);
and U3668 (N_3668,N_3587,N_3520);
nor U3669 (N_3669,N_3530,N_3508);
xor U3670 (N_3670,N_3568,N_3478);
nand U3671 (N_3671,N_3438,N_3443);
nand U3672 (N_3672,N_3441,N_3512);
or U3673 (N_3673,N_3499,N_3405);
and U3674 (N_3674,N_3467,N_3436);
nand U3675 (N_3675,N_3501,N_3503);
nand U3676 (N_3676,N_3551,N_3566);
and U3677 (N_3677,N_3426,N_3411);
and U3678 (N_3678,N_3532,N_3445);
or U3679 (N_3679,N_3429,N_3459);
nor U3680 (N_3680,N_3505,N_3400);
or U3681 (N_3681,N_3550,N_3522);
nand U3682 (N_3682,N_3517,N_3449);
xnor U3683 (N_3683,N_3572,N_3515);
nor U3684 (N_3684,N_3538,N_3466);
nand U3685 (N_3685,N_3456,N_3594);
nor U3686 (N_3686,N_3418,N_3432);
and U3687 (N_3687,N_3590,N_3414);
nand U3688 (N_3688,N_3464,N_3513);
nor U3689 (N_3689,N_3475,N_3593);
nor U3690 (N_3690,N_3494,N_3533);
xnor U3691 (N_3691,N_3562,N_3481);
and U3692 (N_3692,N_3542,N_3507);
nor U3693 (N_3693,N_3460,N_3489);
nor U3694 (N_3694,N_3442,N_3548);
nand U3695 (N_3695,N_3461,N_3422);
and U3696 (N_3696,N_3523,N_3564);
or U3697 (N_3697,N_3471,N_3428);
nand U3698 (N_3698,N_3403,N_3546);
nor U3699 (N_3699,N_3574,N_3448);
nor U3700 (N_3700,N_3418,N_3490);
nand U3701 (N_3701,N_3437,N_3562);
nand U3702 (N_3702,N_3591,N_3572);
or U3703 (N_3703,N_3490,N_3493);
nor U3704 (N_3704,N_3558,N_3445);
nand U3705 (N_3705,N_3565,N_3570);
and U3706 (N_3706,N_3542,N_3509);
or U3707 (N_3707,N_3400,N_3405);
or U3708 (N_3708,N_3470,N_3454);
and U3709 (N_3709,N_3586,N_3593);
nor U3710 (N_3710,N_3422,N_3479);
nand U3711 (N_3711,N_3510,N_3453);
nand U3712 (N_3712,N_3402,N_3474);
or U3713 (N_3713,N_3476,N_3464);
nor U3714 (N_3714,N_3524,N_3581);
and U3715 (N_3715,N_3461,N_3531);
or U3716 (N_3716,N_3496,N_3436);
nand U3717 (N_3717,N_3434,N_3410);
nor U3718 (N_3718,N_3565,N_3591);
nor U3719 (N_3719,N_3520,N_3567);
nand U3720 (N_3720,N_3468,N_3562);
and U3721 (N_3721,N_3426,N_3580);
and U3722 (N_3722,N_3564,N_3444);
and U3723 (N_3723,N_3541,N_3487);
and U3724 (N_3724,N_3588,N_3474);
xor U3725 (N_3725,N_3449,N_3438);
xor U3726 (N_3726,N_3595,N_3554);
and U3727 (N_3727,N_3406,N_3435);
nor U3728 (N_3728,N_3448,N_3521);
and U3729 (N_3729,N_3540,N_3462);
nor U3730 (N_3730,N_3540,N_3486);
nor U3731 (N_3731,N_3515,N_3596);
and U3732 (N_3732,N_3504,N_3410);
nor U3733 (N_3733,N_3537,N_3504);
nor U3734 (N_3734,N_3535,N_3588);
nor U3735 (N_3735,N_3530,N_3525);
nor U3736 (N_3736,N_3483,N_3442);
and U3737 (N_3737,N_3479,N_3578);
or U3738 (N_3738,N_3486,N_3597);
and U3739 (N_3739,N_3507,N_3552);
nor U3740 (N_3740,N_3444,N_3535);
nor U3741 (N_3741,N_3408,N_3401);
nand U3742 (N_3742,N_3416,N_3579);
or U3743 (N_3743,N_3434,N_3512);
or U3744 (N_3744,N_3419,N_3448);
and U3745 (N_3745,N_3546,N_3545);
and U3746 (N_3746,N_3480,N_3464);
and U3747 (N_3747,N_3510,N_3432);
nand U3748 (N_3748,N_3525,N_3571);
or U3749 (N_3749,N_3516,N_3467);
nor U3750 (N_3750,N_3501,N_3414);
and U3751 (N_3751,N_3448,N_3452);
or U3752 (N_3752,N_3514,N_3439);
and U3753 (N_3753,N_3455,N_3584);
or U3754 (N_3754,N_3561,N_3400);
nand U3755 (N_3755,N_3439,N_3558);
and U3756 (N_3756,N_3578,N_3599);
nand U3757 (N_3757,N_3574,N_3562);
or U3758 (N_3758,N_3474,N_3423);
nor U3759 (N_3759,N_3529,N_3421);
and U3760 (N_3760,N_3523,N_3590);
and U3761 (N_3761,N_3581,N_3484);
nor U3762 (N_3762,N_3459,N_3476);
nand U3763 (N_3763,N_3584,N_3429);
nand U3764 (N_3764,N_3562,N_3535);
nand U3765 (N_3765,N_3429,N_3597);
and U3766 (N_3766,N_3491,N_3550);
xnor U3767 (N_3767,N_3513,N_3550);
or U3768 (N_3768,N_3544,N_3555);
or U3769 (N_3769,N_3470,N_3576);
xnor U3770 (N_3770,N_3521,N_3482);
and U3771 (N_3771,N_3483,N_3437);
nor U3772 (N_3772,N_3477,N_3550);
nand U3773 (N_3773,N_3559,N_3480);
or U3774 (N_3774,N_3530,N_3543);
and U3775 (N_3775,N_3534,N_3481);
xor U3776 (N_3776,N_3557,N_3567);
or U3777 (N_3777,N_3452,N_3456);
nand U3778 (N_3778,N_3577,N_3448);
or U3779 (N_3779,N_3583,N_3517);
nand U3780 (N_3780,N_3422,N_3493);
nand U3781 (N_3781,N_3446,N_3502);
nor U3782 (N_3782,N_3473,N_3415);
or U3783 (N_3783,N_3469,N_3595);
and U3784 (N_3784,N_3535,N_3499);
nand U3785 (N_3785,N_3429,N_3490);
nand U3786 (N_3786,N_3581,N_3580);
nand U3787 (N_3787,N_3438,N_3558);
nor U3788 (N_3788,N_3430,N_3466);
and U3789 (N_3789,N_3474,N_3432);
xor U3790 (N_3790,N_3502,N_3404);
nand U3791 (N_3791,N_3462,N_3474);
nor U3792 (N_3792,N_3559,N_3437);
or U3793 (N_3793,N_3525,N_3472);
or U3794 (N_3794,N_3559,N_3537);
nor U3795 (N_3795,N_3544,N_3401);
and U3796 (N_3796,N_3486,N_3444);
nor U3797 (N_3797,N_3419,N_3526);
nand U3798 (N_3798,N_3417,N_3413);
nor U3799 (N_3799,N_3522,N_3495);
and U3800 (N_3800,N_3711,N_3748);
nor U3801 (N_3801,N_3641,N_3710);
nand U3802 (N_3802,N_3760,N_3714);
nor U3803 (N_3803,N_3619,N_3709);
or U3804 (N_3804,N_3729,N_3643);
or U3805 (N_3805,N_3642,N_3614);
or U3806 (N_3806,N_3617,N_3741);
or U3807 (N_3807,N_3670,N_3751);
xnor U3808 (N_3808,N_3633,N_3661);
nor U3809 (N_3809,N_3693,N_3708);
nor U3810 (N_3810,N_3679,N_3790);
or U3811 (N_3811,N_3684,N_3724);
nor U3812 (N_3812,N_3668,N_3785);
nand U3813 (N_3813,N_3607,N_3777);
xnor U3814 (N_3814,N_3783,N_3782);
nand U3815 (N_3815,N_3610,N_3773);
nand U3816 (N_3816,N_3772,N_3667);
nor U3817 (N_3817,N_3701,N_3658);
nand U3818 (N_3818,N_3734,N_3771);
nor U3819 (N_3819,N_3722,N_3675);
and U3820 (N_3820,N_3739,N_3742);
nand U3821 (N_3821,N_3789,N_3750);
or U3822 (N_3822,N_3612,N_3743);
nor U3823 (N_3823,N_3707,N_3753);
nor U3824 (N_3824,N_3629,N_3705);
or U3825 (N_3825,N_3616,N_3737);
nor U3826 (N_3826,N_3627,N_3792);
or U3827 (N_3827,N_3674,N_3779);
nand U3828 (N_3828,N_3600,N_3728);
nand U3829 (N_3829,N_3637,N_3695);
nor U3830 (N_3830,N_3796,N_3632);
and U3831 (N_3831,N_3780,N_3654);
and U3832 (N_3832,N_3699,N_3788);
nor U3833 (N_3833,N_3700,N_3769);
nor U3834 (N_3834,N_3645,N_3656);
nor U3835 (N_3835,N_3636,N_3770);
nand U3836 (N_3836,N_3676,N_3786);
and U3837 (N_3837,N_3752,N_3669);
nand U3838 (N_3838,N_3683,N_3652);
nand U3839 (N_3839,N_3744,N_3687);
nand U3840 (N_3840,N_3758,N_3625);
nand U3841 (N_3841,N_3601,N_3733);
or U3842 (N_3842,N_3776,N_3746);
xnor U3843 (N_3843,N_3762,N_3621);
and U3844 (N_3844,N_3798,N_3749);
nor U3845 (N_3845,N_3678,N_3720);
or U3846 (N_3846,N_3606,N_3723);
nand U3847 (N_3847,N_3694,N_3639);
nand U3848 (N_3848,N_3623,N_3774);
or U3849 (N_3849,N_3657,N_3756);
nand U3850 (N_3850,N_3725,N_3673);
nand U3851 (N_3851,N_3680,N_3635);
or U3852 (N_3852,N_3763,N_3795);
nand U3853 (N_3853,N_3712,N_3640);
or U3854 (N_3854,N_3787,N_3799);
nor U3855 (N_3855,N_3791,N_3630);
and U3856 (N_3856,N_3618,N_3747);
nand U3857 (N_3857,N_3745,N_3653);
and U3858 (N_3858,N_3682,N_3647);
and U3859 (N_3859,N_3650,N_3626);
nor U3860 (N_3860,N_3784,N_3648);
or U3861 (N_3861,N_3721,N_3624);
nor U3862 (N_3862,N_3688,N_3740);
nor U3863 (N_3863,N_3697,N_3690);
and U3864 (N_3864,N_3761,N_3768);
or U3865 (N_3865,N_3759,N_3660);
and U3866 (N_3866,N_3691,N_3730);
xor U3867 (N_3867,N_3704,N_3732);
nand U3868 (N_3868,N_3608,N_3738);
nand U3869 (N_3869,N_3696,N_3659);
or U3870 (N_3870,N_3628,N_3764);
or U3871 (N_3871,N_3655,N_3726);
nand U3872 (N_3872,N_3775,N_3681);
nand U3873 (N_3873,N_3649,N_3703);
xnor U3874 (N_3874,N_3755,N_3731);
and U3875 (N_3875,N_3757,N_3797);
xor U3876 (N_3876,N_3677,N_3646);
or U3877 (N_3877,N_3727,N_3794);
and U3878 (N_3878,N_3644,N_3717);
or U3879 (N_3879,N_3613,N_3615);
or U3880 (N_3880,N_3793,N_3716);
nor U3881 (N_3881,N_3651,N_3778);
or U3882 (N_3882,N_3718,N_3754);
nand U3883 (N_3883,N_3686,N_3672);
nand U3884 (N_3884,N_3664,N_3634);
nor U3885 (N_3885,N_3765,N_3631);
and U3886 (N_3886,N_3604,N_3620);
or U3887 (N_3887,N_3766,N_3663);
nand U3888 (N_3888,N_3609,N_3736);
xor U3889 (N_3889,N_3662,N_3685);
or U3890 (N_3890,N_3689,N_3715);
nand U3891 (N_3891,N_3692,N_3735);
or U3892 (N_3892,N_3781,N_3713);
or U3893 (N_3893,N_3702,N_3611);
nand U3894 (N_3894,N_3602,N_3605);
and U3895 (N_3895,N_3767,N_3665);
nand U3896 (N_3896,N_3706,N_3603);
or U3897 (N_3897,N_3666,N_3638);
nand U3898 (N_3898,N_3698,N_3719);
or U3899 (N_3899,N_3671,N_3622);
nor U3900 (N_3900,N_3673,N_3787);
nand U3901 (N_3901,N_3625,N_3684);
and U3902 (N_3902,N_3702,N_3642);
or U3903 (N_3903,N_3609,N_3681);
nand U3904 (N_3904,N_3779,N_3723);
nand U3905 (N_3905,N_3611,N_3674);
and U3906 (N_3906,N_3790,N_3639);
and U3907 (N_3907,N_3742,N_3701);
nand U3908 (N_3908,N_3703,N_3616);
nor U3909 (N_3909,N_3699,N_3653);
nor U3910 (N_3910,N_3696,N_3646);
nand U3911 (N_3911,N_3613,N_3634);
nor U3912 (N_3912,N_3712,N_3767);
nand U3913 (N_3913,N_3607,N_3654);
or U3914 (N_3914,N_3659,N_3654);
and U3915 (N_3915,N_3621,N_3787);
nor U3916 (N_3916,N_3621,N_3701);
nand U3917 (N_3917,N_3731,N_3637);
nand U3918 (N_3918,N_3670,N_3665);
nand U3919 (N_3919,N_3733,N_3776);
or U3920 (N_3920,N_3799,N_3788);
or U3921 (N_3921,N_3651,N_3650);
nor U3922 (N_3922,N_3709,N_3659);
or U3923 (N_3923,N_3763,N_3652);
or U3924 (N_3924,N_3723,N_3757);
nand U3925 (N_3925,N_3617,N_3797);
nand U3926 (N_3926,N_3693,N_3629);
nor U3927 (N_3927,N_3643,N_3718);
xnor U3928 (N_3928,N_3737,N_3633);
nand U3929 (N_3929,N_3731,N_3642);
nand U3930 (N_3930,N_3663,N_3670);
or U3931 (N_3931,N_3739,N_3791);
nor U3932 (N_3932,N_3628,N_3798);
xnor U3933 (N_3933,N_3767,N_3683);
or U3934 (N_3934,N_3776,N_3649);
xor U3935 (N_3935,N_3628,N_3637);
and U3936 (N_3936,N_3680,N_3666);
nand U3937 (N_3937,N_3679,N_3650);
nor U3938 (N_3938,N_3640,N_3642);
nor U3939 (N_3939,N_3710,N_3709);
nor U3940 (N_3940,N_3744,N_3686);
or U3941 (N_3941,N_3761,N_3726);
nand U3942 (N_3942,N_3763,N_3689);
nand U3943 (N_3943,N_3798,N_3690);
nand U3944 (N_3944,N_3661,N_3763);
nand U3945 (N_3945,N_3758,N_3728);
nor U3946 (N_3946,N_3747,N_3791);
and U3947 (N_3947,N_3750,N_3765);
or U3948 (N_3948,N_3648,N_3723);
or U3949 (N_3949,N_3735,N_3623);
nand U3950 (N_3950,N_3648,N_3711);
nor U3951 (N_3951,N_3645,N_3707);
nand U3952 (N_3952,N_3762,N_3742);
xnor U3953 (N_3953,N_3650,N_3676);
xnor U3954 (N_3954,N_3610,N_3604);
nand U3955 (N_3955,N_3779,N_3697);
and U3956 (N_3956,N_3712,N_3678);
and U3957 (N_3957,N_3642,N_3675);
and U3958 (N_3958,N_3776,N_3695);
nand U3959 (N_3959,N_3684,N_3708);
and U3960 (N_3960,N_3650,N_3742);
and U3961 (N_3961,N_3669,N_3753);
nor U3962 (N_3962,N_3719,N_3797);
nor U3963 (N_3963,N_3778,N_3722);
nor U3964 (N_3964,N_3704,N_3760);
nand U3965 (N_3965,N_3655,N_3657);
and U3966 (N_3966,N_3762,N_3618);
nand U3967 (N_3967,N_3721,N_3760);
nand U3968 (N_3968,N_3685,N_3688);
and U3969 (N_3969,N_3648,N_3652);
nor U3970 (N_3970,N_3684,N_3750);
and U3971 (N_3971,N_3735,N_3755);
nor U3972 (N_3972,N_3730,N_3630);
and U3973 (N_3973,N_3604,N_3625);
nand U3974 (N_3974,N_3642,N_3645);
or U3975 (N_3975,N_3750,N_3625);
or U3976 (N_3976,N_3688,N_3777);
or U3977 (N_3977,N_3643,N_3721);
and U3978 (N_3978,N_3648,N_3754);
or U3979 (N_3979,N_3789,N_3682);
and U3980 (N_3980,N_3790,N_3601);
nor U3981 (N_3981,N_3643,N_3755);
nor U3982 (N_3982,N_3664,N_3604);
nand U3983 (N_3983,N_3755,N_3637);
and U3984 (N_3984,N_3664,N_3684);
or U3985 (N_3985,N_3797,N_3751);
nor U3986 (N_3986,N_3723,N_3671);
xor U3987 (N_3987,N_3640,N_3763);
or U3988 (N_3988,N_3690,N_3662);
nand U3989 (N_3989,N_3725,N_3666);
and U3990 (N_3990,N_3725,N_3702);
nand U3991 (N_3991,N_3691,N_3646);
nor U3992 (N_3992,N_3750,N_3680);
or U3993 (N_3993,N_3671,N_3673);
nand U3994 (N_3994,N_3766,N_3626);
xor U3995 (N_3995,N_3773,N_3759);
nand U3996 (N_3996,N_3654,N_3670);
nand U3997 (N_3997,N_3683,N_3681);
xor U3998 (N_3998,N_3603,N_3636);
or U3999 (N_3999,N_3698,N_3641);
nand U4000 (N_4000,N_3912,N_3867);
and U4001 (N_4001,N_3918,N_3891);
or U4002 (N_4002,N_3995,N_3846);
nand U4003 (N_4003,N_3884,N_3914);
or U4004 (N_4004,N_3893,N_3938);
and U4005 (N_4005,N_3848,N_3942);
or U4006 (N_4006,N_3871,N_3864);
or U4007 (N_4007,N_3982,N_3911);
xnor U4008 (N_4008,N_3989,N_3837);
nor U4009 (N_4009,N_3929,N_3850);
nor U4010 (N_4010,N_3983,N_3957);
or U4011 (N_4011,N_3817,N_3879);
nand U4012 (N_4012,N_3882,N_3999);
or U4013 (N_4013,N_3908,N_3892);
and U4014 (N_4014,N_3840,N_3830);
nand U4015 (N_4015,N_3889,N_3845);
nand U4016 (N_4016,N_3826,N_3812);
and U4017 (N_4017,N_3964,N_3880);
nand U4018 (N_4018,N_3854,N_3800);
xor U4019 (N_4019,N_3819,N_3910);
nand U4020 (N_4020,N_3906,N_3838);
or U4021 (N_4021,N_3897,N_3927);
or U4022 (N_4022,N_3921,N_3990);
nand U4023 (N_4023,N_3959,N_3919);
nand U4024 (N_4024,N_3898,N_3954);
xnor U4025 (N_4025,N_3976,N_3886);
nor U4026 (N_4026,N_3814,N_3847);
nor U4027 (N_4027,N_3857,N_3907);
nand U4028 (N_4028,N_3988,N_3941);
nand U4029 (N_4029,N_3993,N_3809);
or U4030 (N_4030,N_3978,N_3934);
or U4031 (N_4031,N_3831,N_3955);
nor U4032 (N_4032,N_3804,N_3943);
nand U4033 (N_4033,N_3870,N_3841);
or U4034 (N_4034,N_3902,N_3947);
nand U4035 (N_4035,N_3913,N_3909);
and U4036 (N_4036,N_3924,N_3997);
nor U4037 (N_4037,N_3931,N_3876);
nand U4038 (N_4038,N_3869,N_3971);
nor U4039 (N_4039,N_3935,N_3904);
nand U4040 (N_4040,N_3899,N_3951);
and U4041 (N_4041,N_3881,N_3915);
nor U4042 (N_4042,N_3962,N_3963);
or U4043 (N_4043,N_3885,N_3808);
nor U4044 (N_4044,N_3832,N_3949);
or U4045 (N_4045,N_3820,N_3900);
and U4046 (N_4046,N_3994,N_3868);
nor U4047 (N_4047,N_3825,N_3984);
and U4048 (N_4048,N_3928,N_3952);
or U4049 (N_4049,N_3968,N_3950);
or U4050 (N_4050,N_3839,N_3862);
or U4051 (N_4051,N_3828,N_3945);
or U4052 (N_4052,N_3888,N_3816);
or U4053 (N_4053,N_3946,N_3925);
nand U4054 (N_4054,N_3975,N_3866);
and U4055 (N_4055,N_3961,N_3834);
xnor U4056 (N_4056,N_3930,N_3822);
xor U4057 (N_4057,N_3933,N_3821);
and U4058 (N_4058,N_3851,N_3855);
and U4059 (N_4059,N_3979,N_3827);
and U4060 (N_4060,N_3944,N_3977);
nand U4061 (N_4061,N_3901,N_3966);
or U4062 (N_4062,N_3823,N_3998);
and U4063 (N_4063,N_3940,N_3872);
or U4064 (N_4064,N_3920,N_3874);
nor U4065 (N_4065,N_3926,N_3953);
and U4066 (N_4066,N_3985,N_3960);
nand U4067 (N_4067,N_3980,N_3923);
nand U4068 (N_4068,N_3860,N_3844);
nor U4069 (N_4069,N_3970,N_3829);
nor U4070 (N_4070,N_3937,N_3895);
nand U4071 (N_4071,N_3936,N_3818);
nand U4072 (N_4072,N_3996,N_3878);
nor U4073 (N_4073,N_3981,N_3967);
nor U4074 (N_4074,N_3852,N_3903);
nor U4075 (N_4075,N_3849,N_3917);
xnor U4076 (N_4076,N_3807,N_3810);
nand U4077 (N_4077,N_3861,N_3805);
nor U4078 (N_4078,N_3875,N_3815);
xnor U4079 (N_4079,N_3890,N_3973);
or U4080 (N_4080,N_3922,N_3965);
or U4081 (N_4081,N_3992,N_3905);
nor U4082 (N_4082,N_3858,N_3932);
nand U4083 (N_4083,N_3877,N_3894);
and U4084 (N_4084,N_3813,N_3916);
and U4085 (N_4085,N_3833,N_3991);
or U4086 (N_4086,N_3948,N_3873);
xnor U4087 (N_4087,N_3843,N_3863);
and U4088 (N_4088,N_3883,N_3986);
or U4089 (N_4089,N_3939,N_3972);
xor U4090 (N_4090,N_3801,N_3856);
nand U4091 (N_4091,N_3956,N_3887);
and U4092 (N_4092,N_3836,N_3842);
and U4093 (N_4093,N_3803,N_3987);
and U4094 (N_4094,N_3865,N_3811);
and U4095 (N_4095,N_3806,N_3802);
nor U4096 (N_4096,N_3974,N_3853);
and U4097 (N_4097,N_3859,N_3958);
nor U4098 (N_4098,N_3835,N_3824);
nand U4099 (N_4099,N_3896,N_3969);
and U4100 (N_4100,N_3986,N_3805);
or U4101 (N_4101,N_3947,N_3960);
or U4102 (N_4102,N_3837,N_3893);
nand U4103 (N_4103,N_3968,N_3952);
nor U4104 (N_4104,N_3879,N_3954);
nor U4105 (N_4105,N_3925,N_3966);
and U4106 (N_4106,N_3935,N_3834);
or U4107 (N_4107,N_3938,N_3880);
nand U4108 (N_4108,N_3939,N_3883);
nor U4109 (N_4109,N_3971,N_3824);
nand U4110 (N_4110,N_3979,N_3973);
or U4111 (N_4111,N_3904,N_3810);
nand U4112 (N_4112,N_3975,N_3890);
and U4113 (N_4113,N_3949,N_3897);
and U4114 (N_4114,N_3926,N_3860);
xnor U4115 (N_4115,N_3817,N_3993);
nand U4116 (N_4116,N_3879,N_3938);
nor U4117 (N_4117,N_3913,N_3855);
xor U4118 (N_4118,N_3916,N_3858);
nand U4119 (N_4119,N_3855,N_3962);
or U4120 (N_4120,N_3812,N_3970);
nand U4121 (N_4121,N_3812,N_3991);
nor U4122 (N_4122,N_3844,N_3970);
and U4123 (N_4123,N_3847,N_3804);
and U4124 (N_4124,N_3841,N_3963);
nor U4125 (N_4125,N_3813,N_3823);
and U4126 (N_4126,N_3825,N_3813);
and U4127 (N_4127,N_3917,N_3898);
nor U4128 (N_4128,N_3996,N_3844);
or U4129 (N_4129,N_3852,N_3921);
nand U4130 (N_4130,N_3810,N_3901);
nand U4131 (N_4131,N_3846,N_3878);
or U4132 (N_4132,N_3927,N_3885);
nor U4133 (N_4133,N_3916,N_3946);
nor U4134 (N_4134,N_3872,N_3889);
and U4135 (N_4135,N_3877,N_3870);
and U4136 (N_4136,N_3802,N_3924);
nand U4137 (N_4137,N_3800,N_3902);
nor U4138 (N_4138,N_3830,N_3993);
nor U4139 (N_4139,N_3815,N_3990);
or U4140 (N_4140,N_3908,N_3939);
and U4141 (N_4141,N_3924,N_3899);
or U4142 (N_4142,N_3955,N_3859);
xor U4143 (N_4143,N_3877,N_3804);
nor U4144 (N_4144,N_3892,N_3903);
or U4145 (N_4145,N_3840,N_3887);
or U4146 (N_4146,N_3921,N_3915);
nor U4147 (N_4147,N_3986,N_3839);
nand U4148 (N_4148,N_3996,N_3924);
nor U4149 (N_4149,N_3948,N_3818);
or U4150 (N_4150,N_3810,N_3962);
and U4151 (N_4151,N_3853,N_3800);
and U4152 (N_4152,N_3938,N_3892);
or U4153 (N_4153,N_3897,N_3806);
nor U4154 (N_4154,N_3932,N_3839);
or U4155 (N_4155,N_3808,N_3930);
and U4156 (N_4156,N_3862,N_3894);
or U4157 (N_4157,N_3820,N_3957);
nor U4158 (N_4158,N_3954,N_3950);
nor U4159 (N_4159,N_3826,N_3828);
nand U4160 (N_4160,N_3909,N_3894);
nor U4161 (N_4161,N_3838,N_3913);
and U4162 (N_4162,N_3952,N_3860);
nand U4163 (N_4163,N_3896,N_3859);
nor U4164 (N_4164,N_3901,N_3984);
nor U4165 (N_4165,N_3910,N_3855);
xnor U4166 (N_4166,N_3863,N_3832);
or U4167 (N_4167,N_3882,N_3862);
nand U4168 (N_4168,N_3831,N_3895);
nand U4169 (N_4169,N_3853,N_3871);
or U4170 (N_4170,N_3816,N_3891);
nand U4171 (N_4171,N_3904,N_3864);
nor U4172 (N_4172,N_3805,N_3977);
or U4173 (N_4173,N_3954,N_3861);
nand U4174 (N_4174,N_3818,N_3997);
nand U4175 (N_4175,N_3838,N_3988);
nand U4176 (N_4176,N_3925,N_3858);
xor U4177 (N_4177,N_3869,N_3831);
and U4178 (N_4178,N_3976,N_3905);
nor U4179 (N_4179,N_3963,N_3856);
nor U4180 (N_4180,N_3940,N_3898);
nand U4181 (N_4181,N_3870,N_3829);
xor U4182 (N_4182,N_3922,N_3860);
nand U4183 (N_4183,N_3984,N_3905);
nor U4184 (N_4184,N_3942,N_3833);
and U4185 (N_4185,N_3886,N_3837);
or U4186 (N_4186,N_3858,N_3989);
and U4187 (N_4187,N_3938,N_3870);
and U4188 (N_4188,N_3801,N_3806);
nand U4189 (N_4189,N_3998,N_3832);
nand U4190 (N_4190,N_3985,N_3833);
or U4191 (N_4191,N_3841,N_3831);
nor U4192 (N_4192,N_3823,N_3859);
xnor U4193 (N_4193,N_3883,N_3897);
and U4194 (N_4194,N_3836,N_3872);
or U4195 (N_4195,N_3983,N_3967);
or U4196 (N_4196,N_3943,N_3999);
nor U4197 (N_4197,N_3918,N_3970);
nor U4198 (N_4198,N_3911,N_3833);
or U4199 (N_4199,N_3971,N_3990);
and U4200 (N_4200,N_4065,N_4105);
nand U4201 (N_4201,N_4097,N_4093);
or U4202 (N_4202,N_4124,N_4165);
nor U4203 (N_4203,N_4012,N_4008);
and U4204 (N_4204,N_4128,N_4166);
nor U4205 (N_4205,N_4111,N_4048);
xor U4206 (N_4206,N_4024,N_4138);
or U4207 (N_4207,N_4196,N_4122);
and U4208 (N_4208,N_4149,N_4033);
nand U4209 (N_4209,N_4009,N_4064);
nor U4210 (N_4210,N_4058,N_4068);
or U4211 (N_4211,N_4055,N_4119);
nor U4212 (N_4212,N_4140,N_4132);
nor U4213 (N_4213,N_4028,N_4017);
nor U4214 (N_4214,N_4034,N_4173);
or U4215 (N_4215,N_4102,N_4154);
nand U4216 (N_4216,N_4164,N_4103);
nand U4217 (N_4217,N_4115,N_4148);
and U4218 (N_4218,N_4189,N_4010);
and U4219 (N_4219,N_4063,N_4133);
or U4220 (N_4220,N_4100,N_4042);
nand U4221 (N_4221,N_4142,N_4180);
nand U4222 (N_4222,N_4083,N_4167);
or U4223 (N_4223,N_4002,N_4080);
nor U4224 (N_4224,N_4062,N_4059);
nand U4225 (N_4225,N_4151,N_4157);
nand U4226 (N_4226,N_4090,N_4091);
nand U4227 (N_4227,N_4060,N_4169);
xnor U4228 (N_4228,N_4141,N_4031);
and U4229 (N_4229,N_4185,N_4073);
nand U4230 (N_4230,N_4075,N_4135);
or U4231 (N_4231,N_4161,N_4013);
nor U4232 (N_4232,N_4172,N_4179);
nor U4233 (N_4233,N_4194,N_4035);
and U4234 (N_4234,N_4095,N_4120);
or U4235 (N_4235,N_4158,N_4022);
or U4236 (N_4236,N_4054,N_4011);
and U4237 (N_4237,N_4087,N_4107);
nor U4238 (N_4238,N_4192,N_4050);
xor U4239 (N_4239,N_4066,N_4136);
nor U4240 (N_4240,N_4076,N_4078);
nor U4241 (N_4241,N_4026,N_4197);
and U4242 (N_4242,N_4004,N_4145);
xnor U4243 (N_4243,N_4146,N_4153);
nand U4244 (N_4244,N_4003,N_4082);
or U4245 (N_4245,N_4067,N_4199);
or U4246 (N_4246,N_4096,N_4036);
or U4247 (N_4247,N_4110,N_4047);
and U4248 (N_4248,N_4195,N_4121);
and U4249 (N_4249,N_4014,N_4190);
nor U4250 (N_4250,N_4046,N_4040);
nand U4251 (N_4251,N_4021,N_4018);
and U4252 (N_4252,N_4170,N_4049);
nor U4253 (N_4253,N_4000,N_4101);
nand U4254 (N_4254,N_4099,N_4051);
and U4255 (N_4255,N_4016,N_4134);
and U4256 (N_4256,N_4043,N_4162);
xnor U4257 (N_4257,N_4094,N_4104);
nor U4258 (N_4258,N_4116,N_4030);
or U4259 (N_4259,N_4125,N_4081);
nor U4260 (N_4260,N_4108,N_4184);
nand U4261 (N_4261,N_4041,N_4126);
and U4262 (N_4262,N_4032,N_4057);
nor U4263 (N_4263,N_4181,N_4117);
nand U4264 (N_4264,N_4175,N_4071);
and U4265 (N_4265,N_4176,N_4006);
or U4266 (N_4266,N_4156,N_4160);
nand U4267 (N_4267,N_4025,N_4056);
nand U4268 (N_4268,N_4143,N_4088);
nand U4269 (N_4269,N_4045,N_4037);
or U4270 (N_4270,N_4113,N_4178);
and U4271 (N_4271,N_4001,N_4144);
nand U4272 (N_4272,N_4044,N_4147);
nor U4273 (N_4273,N_4069,N_4077);
nor U4274 (N_4274,N_4061,N_4005);
nor U4275 (N_4275,N_4152,N_4007);
and U4276 (N_4276,N_4070,N_4130);
or U4277 (N_4277,N_4177,N_4131);
and U4278 (N_4278,N_4053,N_4193);
and U4279 (N_4279,N_4139,N_4155);
nand U4280 (N_4280,N_4086,N_4191);
nor U4281 (N_4281,N_4137,N_4098);
and U4282 (N_4282,N_4015,N_4187);
nor U4283 (N_4283,N_4198,N_4038);
and U4284 (N_4284,N_4039,N_4027);
or U4285 (N_4285,N_4072,N_4074);
xnor U4286 (N_4286,N_4183,N_4186);
and U4287 (N_4287,N_4085,N_4118);
nor U4288 (N_4288,N_4163,N_4052);
nand U4289 (N_4289,N_4127,N_4109);
and U4290 (N_4290,N_4129,N_4019);
or U4291 (N_4291,N_4159,N_4171);
nor U4292 (N_4292,N_4150,N_4188);
nand U4293 (N_4293,N_4123,N_4092);
and U4294 (N_4294,N_4174,N_4112);
and U4295 (N_4295,N_4020,N_4168);
nand U4296 (N_4296,N_4089,N_4106);
and U4297 (N_4297,N_4084,N_4023);
xnor U4298 (N_4298,N_4182,N_4079);
nand U4299 (N_4299,N_4029,N_4114);
nor U4300 (N_4300,N_4144,N_4155);
xnor U4301 (N_4301,N_4161,N_4037);
nand U4302 (N_4302,N_4052,N_4178);
or U4303 (N_4303,N_4100,N_4046);
or U4304 (N_4304,N_4096,N_4131);
and U4305 (N_4305,N_4094,N_4120);
and U4306 (N_4306,N_4010,N_4181);
or U4307 (N_4307,N_4028,N_4174);
xnor U4308 (N_4308,N_4022,N_4021);
and U4309 (N_4309,N_4085,N_4129);
nand U4310 (N_4310,N_4108,N_4093);
and U4311 (N_4311,N_4103,N_4163);
and U4312 (N_4312,N_4128,N_4035);
xor U4313 (N_4313,N_4104,N_4128);
or U4314 (N_4314,N_4025,N_4181);
nor U4315 (N_4315,N_4150,N_4069);
and U4316 (N_4316,N_4083,N_4126);
or U4317 (N_4317,N_4062,N_4186);
or U4318 (N_4318,N_4092,N_4144);
and U4319 (N_4319,N_4108,N_4160);
nor U4320 (N_4320,N_4149,N_4130);
nor U4321 (N_4321,N_4027,N_4012);
or U4322 (N_4322,N_4090,N_4088);
and U4323 (N_4323,N_4014,N_4018);
nor U4324 (N_4324,N_4036,N_4124);
or U4325 (N_4325,N_4121,N_4173);
nor U4326 (N_4326,N_4182,N_4032);
nor U4327 (N_4327,N_4143,N_4124);
or U4328 (N_4328,N_4131,N_4013);
and U4329 (N_4329,N_4144,N_4076);
nand U4330 (N_4330,N_4072,N_4193);
and U4331 (N_4331,N_4196,N_4121);
nor U4332 (N_4332,N_4109,N_4082);
nand U4333 (N_4333,N_4068,N_4118);
nand U4334 (N_4334,N_4154,N_4131);
nand U4335 (N_4335,N_4012,N_4024);
or U4336 (N_4336,N_4084,N_4019);
nor U4337 (N_4337,N_4193,N_4017);
nor U4338 (N_4338,N_4020,N_4191);
nand U4339 (N_4339,N_4163,N_4058);
nor U4340 (N_4340,N_4108,N_4012);
nor U4341 (N_4341,N_4126,N_4144);
and U4342 (N_4342,N_4160,N_4161);
and U4343 (N_4343,N_4067,N_4089);
and U4344 (N_4344,N_4100,N_4001);
nand U4345 (N_4345,N_4056,N_4081);
or U4346 (N_4346,N_4018,N_4182);
nand U4347 (N_4347,N_4162,N_4149);
or U4348 (N_4348,N_4040,N_4074);
nand U4349 (N_4349,N_4178,N_4050);
and U4350 (N_4350,N_4048,N_4050);
or U4351 (N_4351,N_4038,N_4086);
or U4352 (N_4352,N_4062,N_4073);
nand U4353 (N_4353,N_4082,N_4149);
nor U4354 (N_4354,N_4122,N_4162);
nor U4355 (N_4355,N_4138,N_4140);
nor U4356 (N_4356,N_4170,N_4032);
and U4357 (N_4357,N_4022,N_4172);
nor U4358 (N_4358,N_4025,N_4094);
nand U4359 (N_4359,N_4150,N_4005);
and U4360 (N_4360,N_4041,N_4181);
xnor U4361 (N_4361,N_4050,N_4076);
xnor U4362 (N_4362,N_4034,N_4108);
nand U4363 (N_4363,N_4128,N_4016);
or U4364 (N_4364,N_4102,N_4140);
nor U4365 (N_4365,N_4088,N_4135);
or U4366 (N_4366,N_4120,N_4151);
xnor U4367 (N_4367,N_4021,N_4019);
nand U4368 (N_4368,N_4174,N_4007);
or U4369 (N_4369,N_4147,N_4139);
nand U4370 (N_4370,N_4074,N_4071);
or U4371 (N_4371,N_4098,N_4167);
or U4372 (N_4372,N_4197,N_4172);
nor U4373 (N_4373,N_4081,N_4015);
and U4374 (N_4374,N_4083,N_4084);
or U4375 (N_4375,N_4123,N_4190);
nand U4376 (N_4376,N_4113,N_4037);
nand U4377 (N_4377,N_4160,N_4056);
or U4378 (N_4378,N_4001,N_4022);
and U4379 (N_4379,N_4094,N_4186);
and U4380 (N_4380,N_4059,N_4065);
nor U4381 (N_4381,N_4147,N_4122);
nor U4382 (N_4382,N_4063,N_4032);
and U4383 (N_4383,N_4118,N_4060);
nor U4384 (N_4384,N_4044,N_4112);
nand U4385 (N_4385,N_4152,N_4050);
nor U4386 (N_4386,N_4095,N_4185);
nor U4387 (N_4387,N_4073,N_4183);
nand U4388 (N_4388,N_4006,N_4136);
nand U4389 (N_4389,N_4142,N_4169);
nor U4390 (N_4390,N_4117,N_4095);
xnor U4391 (N_4391,N_4107,N_4114);
nor U4392 (N_4392,N_4085,N_4020);
nand U4393 (N_4393,N_4043,N_4186);
nand U4394 (N_4394,N_4069,N_4148);
nand U4395 (N_4395,N_4137,N_4032);
and U4396 (N_4396,N_4092,N_4063);
nor U4397 (N_4397,N_4050,N_4137);
and U4398 (N_4398,N_4030,N_4003);
nand U4399 (N_4399,N_4001,N_4040);
nor U4400 (N_4400,N_4379,N_4347);
xor U4401 (N_4401,N_4350,N_4295);
nor U4402 (N_4402,N_4290,N_4258);
or U4403 (N_4403,N_4275,N_4324);
nand U4404 (N_4404,N_4376,N_4255);
and U4405 (N_4405,N_4213,N_4368);
nor U4406 (N_4406,N_4367,N_4221);
or U4407 (N_4407,N_4325,N_4242);
nand U4408 (N_4408,N_4340,N_4253);
and U4409 (N_4409,N_4264,N_4285);
or U4410 (N_4410,N_4202,N_4338);
nand U4411 (N_4411,N_4215,N_4280);
xnor U4412 (N_4412,N_4320,N_4303);
and U4413 (N_4413,N_4297,N_4336);
nor U4414 (N_4414,N_4286,N_4262);
xnor U4415 (N_4415,N_4276,N_4267);
nor U4416 (N_4416,N_4212,N_4227);
or U4417 (N_4417,N_4344,N_4391);
nand U4418 (N_4418,N_4229,N_4223);
or U4419 (N_4419,N_4389,N_4399);
xnor U4420 (N_4420,N_4291,N_4312);
nand U4421 (N_4421,N_4374,N_4300);
nor U4422 (N_4422,N_4385,N_4284);
and U4423 (N_4423,N_4259,N_4270);
and U4424 (N_4424,N_4304,N_4266);
and U4425 (N_4425,N_4332,N_4355);
and U4426 (N_4426,N_4279,N_4386);
nor U4427 (N_4427,N_4217,N_4211);
or U4428 (N_4428,N_4366,N_4306);
nor U4429 (N_4429,N_4214,N_4283);
nor U4430 (N_4430,N_4346,N_4319);
nor U4431 (N_4431,N_4268,N_4354);
nand U4432 (N_4432,N_4226,N_4220);
and U4433 (N_4433,N_4353,N_4390);
nor U4434 (N_4434,N_4233,N_4236);
nand U4435 (N_4435,N_4205,N_4360);
nand U4436 (N_4436,N_4231,N_4370);
nand U4437 (N_4437,N_4362,N_4373);
nor U4438 (N_4438,N_4398,N_4357);
nand U4439 (N_4439,N_4250,N_4210);
and U4440 (N_4440,N_4252,N_4382);
and U4441 (N_4441,N_4311,N_4200);
xor U4442 (N_4442,N_4341,N_4307);
or U4443 (N_4443,N_4292,N_4239);
nand U4444 (N_4444,N_4396,N_4343);
or U4445 (N_4445,N_4281,N_4310);
nor U4446 (N_4446,N_4287,N_4257);
or U4447 (N_4447,N_4260,N_4241);
nand U4448 (N_4448,N_4321,N_4216);
nor U4449 (N_4449,N_4372,N_4269);
nor U4450 (N_4450,N_4247,N_4378);
nand U4451 (N_4451,N_4203,N_4331);
nor U4452 (N_4452,N_4380,N_4228);
nand U4453 (N_4453,N_4327,N_4309);
nand U4454 (N_4454,N_4371,N_4298);
nor U4455 (N_4455,N_4333,N_4206);
nor U4456 (N_4456,N_4289,N_4274);
and U4457 (N_4457,N_4294,N_4238);
xnor U4458 (N_4458,N_4265,N_4271);
or U4459 (N_4459,N_4356,N_4335);
nor U4460 (N_4460,N_4358,N_4234);
and U4461 (N_4461,N_4256,N_4393);
nor U4462 (N_4462,N_4384,N_4245);
nand U4463 (N_4463,N_4388,N_4337);
nand U4464 (N_4464,N_4244,N_4278);
nor U4465 (N_4465,N_4375,N_4282);
and U4466 (N_4466,N_4272,N_4313);
nor U4467 (N_4467,N_4249,N_4235);
nor U4468 (N_4468,N_4383,N_4251);
and U4469 (N_4469,N_4322,N_4369);
nand U4470 (N_4470,N_4316,N_4394);
or U4471 (N_4471,N_4326,N_4334);
nor U4472 (N_4472,N_4293,N_4365);
and U4473 (N_4473,N_4273,N_4329);
or U4474 (N_4474,N_4222,N_4208);
nor U4475 (N_4475,N_4330,N_4345);
and U4476 (N_4476,N_4387,N_4288);
nand U4477 (N_4477,N_4392,N_4315);
nor U4478 (N_4478,N_4302,N_4230);
nor U4479 (N_4479,N_4240,N_4348);
nand U4480 (N_4480,N_4209,N_4248);
nand U4481 (N_4481,N_4381,N_4377);
and U4482 (N_4482,N_4263,N_4296);
nor U4483 (N_4483,N_4301,N_4232);
nand U4484 (N_4484,N_4395,N_4299);
or U4485 (N_4485,N_4219,N_4397);
nand U4486 (N_4486,N_4218,N_4361);
or U4487 (N_4487,N_4237,N_4359);
xor U4488 (N_4488,N_4243,N_4254);
or U4489 (N_4489,N_4261,N_4207);
xor U4490 (N_4490,N_4339,N_4328);
or U4491 (N_4491,N_4364,N_4246);
nand U4492 (N_4492,N_4342,N_4318);
or U4493 (N_4493,N_4224,N_4363);
or U4494 (N_4494,N_4225,N_4308);
and U4495 (N_4495,N_4204,N_4314);
nor U4496 (N_4496,N_4349,N_4277);
or U4497 (N_4497,N_4323,N_4317);
nand U4498 (N_4498,N_4305,N_4352);
nor U4499 (N_4499,N_4351,N_4201);
and U4500 (N_4500,N_4269,N_4249);
nor U4501 (N_4501,N_4365,N_4274);
or U4502 (N_4502,N_4209,N_4222);
xor U4503 (N_4503,N_4399,N_4356);
nand U4504 (N_4504,N_4223,N_4393);
or U4505 (N_4505,N_4353,N_4332);
nor U4506 (N_4506,N_4340,N_4352);
or U4507 (N_4507,N_4307,N_4210);
and U4508 (N_4508,N_4278,N_4245);
and U4509 (N_4509,N_4285,N_4210);
nand U4510 (N_4510,N_4379,N_4230);
or U4511 (N_4511,N_4298,N_4251);
xor U4512 (N_4512,N_4239,N_4202);
nand U4513 (N_4513,N_4292,N_4393);
or U4514 (N_4514,N_4204,N_4389);
xnor U4515 (N_4515,N_4208,N_4202);
nand U4516 (N_4516,N_4388,N_4381);
and U4517 (N_4517,N_4369,N_4326);
nand U4518 (N_4518,N_4354,N_4312);
or U4519 (N_4519,N_4371,N_4348);
nand U4520 (N_4520,N_4288,N_4217);
or U4521 (N_4521,N_4370,N_4316);
or U4522 (N_4522,N_4317,N_4242);
nand U4523 (N_4523,N_4369,N_4246);
and U4524 (N_4524,N_4240,N_4296);
and U4525 (N_4525,N_4362,N_4338);
or U4526 (N_4526,N_4394,N_4256);
nor U4527 (N_4527,N_4208,N_4308);
nand U4528 (N_4528,N_4347,N_4373);
or U4529 (N_4529,N_4207,N_4237);
nand U4530 (N_4530,N_4364,N_4310);
xor U4531 (N_4531,N_4301,N_4392);
and U4532 (N_4532,N_4217,N_4277);
or U4533 (N_4533,N_4358,N_4287);
nor U4534 (N_4534,N_4264,N_4317);
nor U4535 (N_4535,N_4251,N_4363);
or U4536 (N_4536,N_4239,N_4358);
xnor U4537 (N_4537,N_4257,N_4335);
nand U4538 (N_4538,N_4214,N_4271);
nor U4539 (N_4539,N_4337,N_4258);
and U4540 (N_4540,N_4381,N_4257);
nor U4541 (N_4541,N_4377,N_4266);
or U4542 (N_4542,N_4398,N_4307);
nor U4543 (N_4543,N_4202,N_4230);
nand U4544 (N_4544,N_4319,N_4344);
and U4545 (N_4545,N_4378,N_4315);
xnor U4546 (N_4546,N_4265,N_4319);
or U4547 (N_4547,N_4205,N_4234);
and U4548 (N_4548,N_4321,N_4329);
or U4549 (N_4549,N_4256,N_4345);
nand U4550 (N_4550,N_4374,N_4217);
xor U4551 (N_4551,N_4204,N_4277);
xnor U4552 (N_4552,N_4342,N_4324);
nor U4553 (N_4553,N_4231,N_4325);
or U4554 (N_4554,N_4391,N_4287);
nor U4555 (N_4555,N_4330,N_4207);
nor U4556 (N_4556,N_4376,N_4248);
and U4557 (N_4557,N_4393,N_4310);
or U4558 (N_4558,N_4367,N_4284);
nor U4559 (N_4559,N_4384,N_4376);
nor U4560 (N_4560,N_4344,N_4262);
or U4561 (N_4561,N_4312,N_4308);
nor U4562 (N_4562,N_4257,N_4375);
nor U4563 (N_4563,N_4391,N_4211);
nand U4564 (N_4564,N_4271,N_4377);
nor U4565 (N_4565,N_4293,N_4276);
and U4566 (N_4566,N_4318,N_4286);
or U4567 (N_4567,N_4355,N_4388);
nand U4568 (N_4568,N_4360,N_4255);
nand U4569 (N_4569,N_4274,N_4270);
nor U4570 (N_4570,N_4353,N_4319);
nor U4571 (N_4571,N_4310,N_4293);
or U4572 (N_4572,N_4381,N_4339);
xnor U4573 (N_4573,N_4374,N_4228);
xnor U4574 (N_4574,N_4278,N_4230);
nor U4575 (N_4575,N_4237,N_4384);
and U4576 (N_4576,N_4335,N_4212);
and U4577 (N_4577,N_4231,N_4380);
nor U4578 (N_4578,N_4393,N_4327);
nor U4579 (N_4579,N_4243,N_4201);
nor U4580 (N_4580,N_4250,N_4389);
nor U4581 (N_4581,N_4324,N_4303);
xor U4582 (N_4582,N_4360,N_4350);
nor U4583 (N_4583,N_4202,N_4363);
and U4584 (N_4584,N_4246,N_4343);
and U4585 (N_4585,N_4251,N_4266);
and U4586 (N_4586,N_4373,N_4207);
nor U4587 (N_4587,N_4275,N_4246);
xnor U4588 (N_4588,N_4266,N_4314);
or U4589 (N_4589,N_4292,N_4281);
nor U4590 (N_4590,N_4392,N_4240);
nor U4591 (N_4591,N_4225,N_4302);
nand U4592 (N_4592,N_4220,N_4295);
and U4593 (N_4593,N_4233,N_4378);
and U4594 (N_4594,N_4241,N_4351);
xnor U4595 (N_4595,N_4350,N_4320);
and U4596 (N_4596,N_4381,N_4217);
and U4597 (N_4597,N_4312,N_4329);
xor U4598 (N_4598,N_4381,N_4247);
nor U4599 (N_4599,N_4378,N_4284);
or U4600 (N_4600,N_4519,N_4558);
xor U4601 (N_4601,N_4506,N_4594);
nand U4602 (N_4602,N_4433,N_4553);
nand U4603 (N_4603,N_4539,N_4442);
or U4604 (N_4604,N_4522,N_4480);
and U4605 (N_4605,N_4491,N_4550);
nor U4606 (N_4606,N_4475,N_4444);
nand U4607 (N_4607,N_4570,N_4422);
or U4608 (N_4608,N_4572,N_4410);
nand U4609 (N_4609,N_4488,N_4441);
nand U4610 (N_4610,N_4530,N_4520);
nor U4611 (N_4611,N_4469,N_4404);
nand U4612 (N_4612,N_4541,N_4402);
or U4613 (N_4613,N_4406,N_4481);
nor U4614 (N_4614,N_4516,N_4489);
nand U4615 (N_4615,N_4436,N_4582);
or U4616 (N_4616,N_4494,N_4577);
nand U4617 (N_4617,N_4545,N_4512);
nor U4618 (N_4618,N_4587,N_4598);
nand U4619 (N_4619,N_4551,N_4467);
nor U4620 (N_4620,N_4499,N_4592);
nor U4621 (N_4621,N_4543,N_4571);
nor U4622 (N_4622,N_4439,N_4403);
nand U4623 (N_4623,N_4446,N_4400);
nand U4624 (N_4624,N_4560,N_4524);
or U4625 (N_4625,N_4596,N_4401);
and U4626 (N_4626,N_4584,N_4454);
or U4627 (N_4627,N_4409,N_4595);
and U4628 (N_4628,N_4473,N_4492);
xnor U4629 (N_4629,N_4430,N_4464);
nand U4630 (N_4630,N_4471,N_4424);
nand U4631 (N_4631,N_4534,N_4423);
and U4632 (N_4632,N_4503,N_4450);
nand U4633 (N_4633,N_4413,N_4426);
nand U4634 (N_4634,N_4452,N_4498);
or U4635 (N_4635,N_4557,N_4527);
nor U4636 (N_4636,N_4579,N_4559);
or U4637 (N_4637,N_4508,N_4420);
nor U4638 (N_4638,N_4448,N_4418);
or U4639 (N_4639,N_4578,N_4497);
nand U4640 (N_4640,N_4537,N_4591);
or U4641 (N_4641,N_4501,N_4563);
nand U4642 (N_4642,N_4581,N_4461);
and U4643 (N_4643,N_4573,N_4419);
or U4644 (N_4644,N_4474,N_4484);
or U4645 (N_4645,N_4496,N_4432);
nor U4646 (N_4646,N_4569,N_4477);
and U4647 (N_4647,N_4412,N_4451);
nand U4648 (N_4648,N_4447,N_4472);
or U4649 (N_4649,N_4405,N_4590);
or U4650 (N_4650,N_4565,N_4556);
nor U4651 (N_4651,N_4415,N_4478);
nor U4652 (N_4652,N_4542,N_4533);
nand U4653 (N_4653,N_4504,N_4438);
nand U4654 (N_4654,N_4547,N_4548);
or U4655 (N_4655,N_4407,N_4487);
nor U4656 (N_4656,N_4549,N_4588);
and U4657 (N_4657,N_4515,N_4417);
or U4658 (N_4658,N_4445,N_4483);
or U4659 (N_4659,N_4552,N_4535);
nor U4660 (N_4660,N_4463,N_4513);
or U4661 (N_4661,N_4583,N_4589);
xor U4662 (N_4662,N_4470,N_4546);
nand U4663 (N_4663,N_4526,N_4544);
xor U4664 (N_4664,N_4599,N_4453);
or U4665 (N_4665,N_4465,N_4505);
nand U4666 (N_4666,N_4455,N_4528);
or U4667 (N_4667,N_4562,N_4434);
or U4668 (N_4668,N_4490,N_4493);
nor U4669 (N_4669,N_4460,N_4532);
and U4670 (N_4670,N_4437,N_4421);
and U4671 (N_4671,N_4459,N_4525);
and U4672 (N_4672,N_4479,N_4427);
nor U4673 (N_4673,N_4456,N_4574);
or U4674 (N_4674,N_4408,N_4538);
nand U4675 (N_4675,N_4443,N_4575);
and U4676 (N_4676,N_4568,N_4428);
nand U4677 (N_4677,N_4540,N_4531);
and U4678 (N_4678,N_4425,N_4567);
or U4679 (N_4679,N_4486,N_4485);
nor U4680 (N_4680,N_4509,N_4435);
nor U4681 (N_4681,N_4466,N_4523);
and U4682 (N_4682,N_4458,N_4536);
nand U4683 (N_4683,N_4482,N_4580);
or U4684 (N_4684,N_4449,N_4431);
nor U4685 (N_4685,N_4554,N_4521);
nor U4686 (N_4686,N_4510,N_4593);
nor U4687 (N_4687,N_4416,N_4514);
or U4688 (N_4688,N_4411,N_4462);
and U4689 (N_4689,N_4566,N_4555);
nand U4690 (N_4690,N_4476,N_4529);
nor U4691 (N_4691,N_4440,N_4517);
and U4692 (N_4692,N_4518,N_4564);
nand U4693 (N_4693,N_4597,N_4457);
xor U4694 (N_4694,N_4500,N_4511);
nand U4695 (N_4695,N_4429,N_4585);
nor U4696 (N_4696,N_4502,N_4468);
or U4697 (N_4697,N_4495,N_4586);
xor U4698 (N_4698,N_4414,N_4507);
and U4699 (N_4699,N_4576,N_4561);
or U4700 (N_4700,N_4429,N_4460);
nor U4701 (N_4701,N_4429,N_4443);
nand U4702 (N_4702,N_4594,N_4543);
or U4703 (N_4703,N_4434,N_4511);
xnor U4704 (N_4704,N_4510,N_4578);
nor U4705 (N_4705,N_4466,N_4532);
nor U4706 (N_4706,N_4536,N_4525);
nand U4707 (N_4707,N_4502,N_4557);
and U4708 (N_4708,N_4573,N_4447);
nor U4709 (N_4709,N_4473,N_4531);
or U4710 (N_4710,N_4537,N_4403);
nor U4711 (N_4711,N_4599,N_4451);
nand U4712 (N_4712,N_4587,N_4464);
or U4713 (N_4713,N_4440,N_4484);
and U4714 (N_4714,N_4434,N_4420);
nor U4715 (N_4715,N_4448,N_4558);
nand U4716 (N_4716,N_4436,N_4496);
nand U4717 (N_4717,N_4522,N_4573);
nand U4718 (N_4718,N_4558,N_4575);
nand U4719 (N_4719,N_4458,N_4443);
and U4720 (N_4720,N_4568,N_4442);
nand U4721 (N_4721,N_4564,N_4591);
xor U4722 (N_4722,N_4567,N_4440);
xnor U4723 (N_4723,N_4571,N_4527);
nor U4724 (N_4724,N_4495,N_4503);
and U4725 (N_4725,N_4507,N_4505);
and U4726 (N_4726,N_4566,N_4582);
and U4727 (N_4727,N_4593,N_4486);
nor U4728 (N_4728,N_4441,N_4426);
nand U4729 (N_4729,N_4499,N_4585);
xor U4730 (N_4730,N_4586,N_4461);
nor U4731 (N_4731,N_4436,N_4589);
nand U4732 (N_4732,N_4536,N_4584);
nor U4733 (N_4733,N_4513,N_4589);
or U4734 (N_4734,N_4571,N_4536);
nand U4735 (N_4735,N_4522,N_4552);
or U4736 (N_4736,N_4423,N_4495);
nor U4737 (N_4737,N_4502,N_4551);
nand U4738 (N_4738,N_4487,N_4579);
or U4739 (N_4739,N_4427,N_4598);
or U4740 (N_4740,N_4403,N_4492);
and U4741 (N_4741,N_4446,N_4444);
or U4742 (N_4742,N_4438,N_4458);
or U4743 (N_4743,N_4497,N_4503);
nor U4744 (N_4744,N_4517,N_4582);
nor U4745 (N_4745,N_4513,N_4429);
nand U4746 (N_4746,N_4547,N_4546);
nor U4747 (N_4747,N_4405,N_4458);
nand U4748 (N_4748,N_4575,N_4507);
nand U4749 (N_4749,N_4401,N_4487);
or U4750 (N_4750,N_4579,N_4523);
and U4751 (N_4751,N_4463,N_4595);
nor U4752 (N_4752,N_4434,N_4446);
nand U4753 (N_4753,N_4456,N_4438);
nand U4754 (N_4754,N_4582,N_4493);
or U4755 (N_4755,N_4462,N_4421);
or U4756 (N_4756,N_4447,N_4508);
nor U4757 (N_4757,N_4533,N_4502);
and U4758 (N_4758,N_4482,N_4426);
nand U4759 (N_4759,N_4552,N_4438);
nand U4760 (N_4760,N_4497,N_4428);
nand U4761 (N_4761,N_4463,N_4483);
nand U4762 (N_4762,N_4575,N_4589);
nand U4763 (N_4763,N_4495,N_4560);
nor U4764 (N_4764,N_4509,N_4453);
nor U4765 (N_4765,N_4406,N_4536);
and U4766 (N_4766,N_4537,N_4551);
or U4767 (N_4767,N_4571,N_4595);
or U4768 (N_4768,N_4581,N_4553);
or U4769 (N_4769,N_4504,N_4547);
nor U4770 (N_4770,N_4472,N_4409);
nand U4771 (N_4771,N_4515,N_4534);
xnor U4772 (N_4772,N_4474,N_4557);
nand U4773 (N_4773,N_4485,N_4475);
or U4774 (N_4774,N_4511,N_4533);
nor U4775 (N_4775,N_4524,N_4443);
nand U4776 (N_4776,N_4414,N_4544);
and U4777 (N_4777,N_4448,N_4436);
or U4778 (N_4778,N_4407,N_4560);
nand U4779 (N_4779,N_4497,N_4523);
xor U4780 (N_4780,N_4564,N_4409);
or U4781 (N_4781,N_4556,N_4448);
nand U4782 (N_4782,N_4565,N_4497);
xor U4783 (N_4783,N_4409,N_4438);
nand U4784 (N_4784,N_4449,N_4416);
or U4785 (N_4785,N_4578,N_4565);
and U4786 (N_4786,N_4524,N_4465);
xor U4787 (N_4787,N_4527,N_4541);
nand U4788 (N_4788,N_4539,N_4425);
or U4789 (N_4789,N_4448,N_4461);
and U4790 (N_4790,N_4402,N_4413);
nor U4791 (N_4791,N_4481,N_4497);
or U4792 (N_4792,N_4535,N_4523);
nand U4793 (N_4793,N_4493,N_4543);
or U4794 (N_4794,N_4575,N_4520);
nor U4795 (N_4795,N_4461,N_4440);
nand U4796 (N_4796,N_4564,N_4461);
and U4797 (N_4797,N_4404,N_4436);
and U4798 (N_4798,N_4586,N_4548);
or U4799 (N_4799,N_4426,N_4476);
or U4800 (N_4800,N_4680,N_4778);
nand U4801 (N_4801,N_4718,N_4753);
nand U4802 (N_4802,N_4758,N_4624);
nor U4803 (N_4803,N_4695,N_4641);
or U4804 (N_4804,N_4616,N_4623);
and U4805 (N_4805,N_4627,N_4713);
xnor U4806 (N_4806,N_4667,N_4781);
xor U4807 (N_4807,N_4744,N_4653);
nor U4808 (N_4808,N_4606,N_4772);
nor U4809 (N_4809,N_4746,N_4619);
and U4810 (N_4810,N_4661,N_4603);
or U4811 (N_4811,N_4711,N_4687);
nor U4812 (N_4812,N_4712,N_4604);
nor U4813 (N_4813,N_4688,N_4782);
nand U4814 (N_4814,N_4662,N_4708);
and U4815 (N_4815,N_4791,N_4632);
or U4816 (N_4816,N_4634,N_4762);
and U4817 (N_4817,N_4664,N_4609);
nand U4818 (N_4818,N_4621,N_4716);
nor U4819 (N_4819,N_4767,N_4790);
xor U4820 (N_4820,N_4613,N_4656);
nor U4821 (N_4821,N_4673,N_4777);
xnor U4822 (N_4822,N_4608,N_4635);
nor U4823 (N_4823,N_4757,N_4703);
xor U4824 (N_4824,N_4660,N_4764);
nor U4825 (N_4825,N_4614,N_4639);
nor U4826 (N_4826,N_4618,N_4721);
or U4827 (N_4827,N_4691,N_4780);
nor U4828 (N_4828,N_4717,N_4737);
nand U4829 (N_4829,N_4643,N_4732);
or U4830 (N_4830,N_4665,N_4766);
xor U4831 (N_4831,N_4788,N_4797);
nor U4832 (N_4832,N_4724,N_4785);
nand U4833 (N_4833,N_4645,N_4742);
nor U4834 (N_4834,N_4622,N_4647);
or U4835 (N_4835,N_4773,N_4607);
nand U4836 (N_4836,N_4676,N_4658);
or U4837 (N_4837,N_4686,N_4625);
and U4838 (N_4838,N_4776,N_4784);
and U4839 (N_4839,N_4699,N_4786);
or U4840 (N_4840,N_4646,N_4705);
nand U4841 (N_4841,N_4605,N_4749);
and U4842 (N_4842,N_4675,N_4770);
nand U4843 (N_4843,N_4640,N_4734);
xnor U4844 (N_4844,N_4650,N_4668);
and U4845 (N_4845,N_4689,N_4638);
and U4846 (N_4846,N_4697,N_4710);
nand U4847 (N_4847,N_4630,N_4652);
nand U4848 (N_4848,N_4736,N_4700);
xor U4849 (N_4849,N_4725,N_4759);
nand U4850 (N_4850,N_4774,N_4733);
and U4851 (N_4851,N_4681,N_4731);
nand U4852 (N_4852,N_4765,N_4756);
or U4853 (N_4853,N_4769,N_4701);
xor U4854 (N_4854,N_4657,N_4706);
and U4855 (N_4855,N_4729,N_4796);
nor U4856 (N_4856,N_4644,N_4611);
or U4857 (N_4857,N_4768,N_4620);
xnor U4858 (N_4858,N_4669,N_4692);
nand U4859 (N_4859,N_4649,N_4787);
and U4860 (N_4860,N_4671,N_4636);
nor U4861 (N_4861,N_4637,N_4685);
nor U4862 (N_4862,N_4722,N_4694);
nor U4863 (N_4863,N_4779,N_4763);
or U4864 (N_4864,N_4743,N_4684);
nand U4865 (N_4865,N_4799,N_4750);
xnor U4866 (N_4866,N_4683,N_4654);
and U4867 (N_4867,N_4792,N_4789);
nor U4868 (N_4868,N_4704,N_4720);
or U4869 (N_4869,N_4723,N_4693);
and U4870 (N_4870,N_4715,N_4748);
nor U4871 (N_4871,N_4615,N_4601);
or U4872 (N_4872,N_4666,N_4670);
and U4873 (N_4873,N_4730,N_4682);
nand U4874 (N_4874,N_4678,N_4727);
and U4875 (N_4875,N_4752,N_4775);
and U4876 (N_4876,N_4663,N_4655);
nor U4877 (N_4877,N_4761,N_4677);
and U4878 (N_4878,N_4709,N_4600);
or U4879 (N_4879,N_4651,N_4751);
and U4880 (N_4880,N_4795,N_4633);
or U4881 (N_4881,N_4745,N_4794);
nand U4882 (N_4882,N_4719,N_4726);
nand U4883 (N_4883,N_4771,N_4798);
xnor U4884 (N_4884,N_4747,N_4642);
or U4885 (N_4885,N_4659,N_4738);
and U4886 (N_4886,N_4612,N_4610);
and U4887 (N_4887,N_4631,N_4755);
and U4888 (N_4888,N_4628,N_4793);
or U4889 (N_4889,N_4617,N_4648);
or U4890 (N_4890,N_4754,N_4602);
or U4891 (N_4891,N_4741,N_4740);
and U4892 (N_4892,N_4626,N_4735);
and U4893 (N_4893,N_4679,N_4760);
nor U4894 (N_4894,N_4783,N_4739);
xor U4895 (N_4895,N_4707,N_4690);
nor U4896 (N_4896,N_4714,N_4702);
xor U4897 (N_4897,N_4674,N_4696);
and U4898 (N_4898,N_4698,N_4672);
nor U4899 (N_4899,N_4728,N_4629);
or U4900 (N_4900,N_4666,N_4624);
nand U4901 (N_4901,N_4626,N_4617);
nor U4902 (N_4902,N_4727,N_4770);
and U4903 (N_4903,N_4607,N_4715);
nand U4904 (N_4904,N_4670,N_4658);
xnor U4905 (N_4905,N_4716,N_4759);
nor U4906 (N_4906,N_4613,N_4669);
and U4907 (N_4907,N_4630,N_4745);
nand U4908 (N_4908,N_4690,N_4657);
or U4909 (N_4909,N_4623,N_4703);
nand U4910 (N_4910,N_4761,N_4620);
nor U4911 (N_4911,N_4695,N_4783);
nor U4912 (N_4912,N_4609,N_4788);
nor U4913 (N_4913,N_4620,N_4712);
or U4914 (N_4914,N_4782,N_4754);
nor U4915 (N_4915,N_4632,N_4798);
and U4916 (N_4916,N_4743,N_4637);
nand U4917 (N_4917,N_4697,N_4695);
nor U4918 (N_4918,N_4603,N_4731);
nand U4919 (N_4919,N_4634,N_4746);
nand U4920 (N_4920,N_4695,N_4768);
nand U4921 (N_4921,N_4715,N_4709);
nand U4922 (N_4922,N_4635,N_4743);
nor U4923 (N_4923,N_4726,N_4708);
nand U4924 (N_4924,N_4648,N_4688);
nor U4925 (N_4925,N_4734,N_4794);
nor U4926 (N_4926,N_4679,N_4754);
or U4927 (N_4927,N_4705,N_4790);
or U4928 (N_4928,N_4791,N_4798);
nor U4929 (N_4929,N_4611,N_4704);
nand U4930 (N_4930,N_4702,N_4620);
nand U4931 (N_4931,N_4662,N_4741);
and U4932 (N_4932,N_4639,N_4765);
nand U4933 (N_4933,N_4619,N_4658);
nor U4934 (N_4934,N_4711,N_4638);
and U4935 (N_4935,N_4785,N_4786);
nand U4936 (N_4936,N_4686,N_4723);
and U4937 (N_4937,N_4623,N_4749);
nor U4938 (N_4938,N_4789,N_4779);
xor U4939 (N_4939,N_4761,N_4686);
nor U4940 (N_4940,N_4616,N_4703);
nand U4941 (N_4941,N_4661,N_4663);
xor U4942 (N_4942,N_4706,N_4679);
nand U4943 (N_4943,N_4680,N_4695);
nand U4944 (N_4944,N_4753,N_4779);
xor U4945 (N_4945,N_4667,N_4747);
nand U4946 (N_4946,N_4681,N_4730);
xnor U4947 (N_4947,N_4712,N_4656);
nor U4948 (N_4948,N_4733,N_4628);
or U4949 (N_4949,N_4778,N_4772);
or U4950 (N_4950,N_4705,N_4752);
nor U4951 (N_4951,N_4732,N_4714);
nor U4952 (N_4952,N_4726,N_4700);
and U4953 (N_4953,N_4779,N_4736);
nor U4954 (N_4954,N_4721,N_4770);
nor U4955 (N_4955,N_4740,N_4771);
nand U4956 (N_4956,N_4661,N_4627);
nor U4957 (N_4957,N_4762,N_4661);
and U4958 (N_4958,N_4743,N_4740);
nand U4959 (N_4959,N_4672,N_4727);
nand U4960 (N_4960,N_4763,N_4688);
nand U4961 (N_4961,N_4613,N_4768);
nand U4962 (N_4962,N_4654,N_4796);
nor U4963 (N_4963,N_4783,N_4666);
nand U4964 (N_4964,N_4679,N_4748);
nor U4965 (N_4965,N_4687,N_4692);
or U4966 (N_4966,N_4687,N_4707);
nand U4967 (N_4967,N_4712,N_4636);
xor U4968 (N_4968,N_4762,N_4639);
or U4969 (N_4969,N_4658,N_4629);
nor U4970 (N_4970,N_4670,N_4604);
nand U4971 (N_4971,N_4694,N_4695);
and U4972 (N_4972,N_4645,N_4677);
nor U4973 (N_4973,N_4670,N_4724);
nor U4974 (N_4974,N_4633,N_4743);
and U4975 (N_4975,N_4764,N_4684);
nand U4976 (N_4976,N_4722,N_4624);
nor U4977 (N_4977,N_4602,N_4737);
nand U4978 (N_4978,N_4664,N_4641);
and U4979 (N_4979,N_4786,N_4722);
nand U4980 (N_4980,N_4789,N_4780);
nand U4981 (N_4981,N_4774,N_4681);
nand U4982 (N_4982,N_4701,N_4717);
and U4983 (N_4983,N_4658,N_4665);
nor U4984 (N_4984,N_4758,N_4611);
and U4985 (N_4985,N_4749,N_4635);
and U4986 (N_4986,N_4671,N_4696);
or U4987 (N_4987,N_4653,N_4671);
nand U4988 (N_4988,N_4603,N_4610);
nand U4989 (N_4989,N_4637,N_4699);
or U4990 (N_4990,N_4740,N_4756);
nand U4991 (N_4991,N_4679,N_4607);
xor U4992 (N_4992,N_4647,N_4620);
nand U4993 (N_4993,N_4775,N_4613);
and U4994 (N_4994,N_4612,N_4616);
nor U4995 (N_4995,N_4757,N_4797);
or U4996 (N_4996,N_4752,N_4724);
nand U4997 (N_4997,N_4621,N_4748);
nand U4998 (N_4998,N_4740,N_4664);
and U4999 (N_4999,N_4651,N_4719);
or UO_0 (O_0,N_4866,N_4889);
or UO_1 (O_1,N_4938,N_4806);
nor UO_2 (O_2,N_4928,N_4812);
nor UO_3 (O_3,N_4958,N_4808);
or UO_4 (O_4,N_4851,N_4945);
xor UO_5 (O_5,N_4983,N_4902);
and UO_6 (O_6,N_4814,N_4877);
xor UO_7 (O_7,N_4936,N_4848);
or UO_8 (O_8,N_4834,N_4916);
and UO_9 (O_9,N_4886,N_4996);
or UO_10 (O_10,N_4910,N_4833);
or UO_11 (O_11,N_4872,N_4839);
and UO_12 (O_12,N_4852,N_4860);
and UO_13 (O_13,N_4980,N_4962);
or UO_14 (O_14,N_4899,N_4894);
nand UO_15 (O_15,N_4967,N_4920);
or UO_16 (O_16,N_4989,N_4895);
and UO_17 (O_17,N_4842,N_4977);
nand UO_18 (O_18,N_4929,N_4971);
and UO_19 (O_19,N_4898,N_4979);
nand UO_20 (O_20,N_4992,N_4932);
or UO_21 (O_21,N_4825,N_4914);
or UO_22 (O_22,N_4884,N_4931);
and UO_23 (O_23,N_4862,N_4816);
and UO_24 (O_24,N_4951,N_4933);
nand UO_25 (O_25,N_4818,N_4876);
nand UO_26 (O_26,N_4952,N_4935);
and UO_27 (O_27,N_4937,N_4800);
nand UO_28 (O_28,N_4900,N_4982);
nor UO_29 (O_29,N_4828,N_4912);
nor UO_30 (O_30,N_4970,N_4981);
or UO_31 (O_31,N_4999,N_4969);
and UO_32 (O_32,N_4864,N_4875);
nor UO_33 (O_33,N_4925,N_4998);
nand UO_34 (O_34,N_4888,N_4819);
nor UO_35 (O_35,N_4890,N_4811);
xor UO_36 (O_36,N_4802,N_4924);
and UO_37 (O_37,N_4896,N_4950);
or UO_38 (O_38,N_4861,N_4904);
and UO_39 (O_39,N_4955,N_4879);
or UO_40 (O_40,N_4949,N_4960);
or UO_41 (O_41,N_4843,N_4984);
or UO_42 (O_42,N_4942,N_4850);
xor UO_43 (O_43,N_4817,N_4887);
nor UO_44 (O_44,N_4838,N_4934);
and UO_45 (O_45,N_4966,N_4845);
and UO_46 (O_46,N_4805,N_4882);
xor UO_47 (O_47,N_4873,N_4885);
xnor UO_48 (O_48,N_4832,N_4804);
nand UO_49 (O_49,N_4993,N_4892);
or UO_50 (O_50,N_4810,N_4959);
nor UO_51 (O_51,N_4847,N_4987);
and UO_52 (O_52,N_4823,N_4893);
nand UO_53 (O_53,N_4827,N_4881);
or UO_54 (O_54,N_4853,N_4880);
and UO_55 (O_55,N_4849,N_4922);
and UO_56 (O_56,N_4995,N_4918);
nor UO_57 (O_57,N_4939,N_4891);
and UO_58 (O_58,N_4907,N_4988);
xor UO_59 (O_59,N_4921,N_4871);
and UO_60 (O_60,N_4826,N_4997);
or UO_61 (O_61,N_4868,N_4854);
and UO_62 (O_62,N_4829,N_4813);
and UO_63 (O_63,N_4883,N_4926);
nor UO_64 (O_64,N_4857,N_4968);
and UO_65 (O_65,N_4975,N_4822);
or UO_66 (O_66,N_4897,N_4836);
xnor UO_67 (O_67,N_4953,N_4944);
nor UO_68 (O_68,N_4903,N_4954);
xor UO_69 (O_69,N_4863,N_4809);
nor UO_70 (O_70,N_4911,N_4986);
and UO_71 (O_71,N_4840,N_4985);
or UO_72 (O_72,N_4824,N_4948);
nand UO_73 (O_73,N_4961,N_4923);
and UO_74 (O_74,N_4919,N_4940);
nor UO_75 (O_75,N_4867,N_4913);
and UO_76 (O_76,N_4909,N_4835);
nor UO_77 (O_77,N_4801,N_4869);
nand UO_78 (O_78,N_4815,N_4973);
or UO_79 (O_79,N_4941,N_4870);
nand UO_80 (O_80,N_4855,N_4901);
nand UO_81 (O_81,N_4859,N_4878);
xor UO_82 (O_82,N_4991,N_4957);
nor UO_83 (O_83,N_4831,N_4874);
nor UO_84 (O_84,N_4820,N_4963);
xnor UO_85 (O_85,N_4964,N_4927);
and UO_86 (O_86,N_4807,N_4841);
nor UO_87 (O_87,N_4858,N_4947);
and UO_88 (O_88,N_4803,N_4976);
nor UO_89 (O_89,N_4908,N_4830);
nor UO_90 (O_90,N_4994,N_4917);
nand UO_91 (O_91,N_4837,N_4906);
nand UO_92 (O_92,N_4965,N_4946);
nand UO_93 (O_93,N_4865,N_4844);
and UO_94 (O_94,N_4990,N_4956);
or UO_95 (O_95,N_4915,N_4978);
xor UO_96 (O_96,N_4974,N_4905);
nor UO_97 (O_97,N_4943,N_4856);
and UO_98 (O_98,N_4821,N_4930);
and UO_99 (O_99,N_4846,N_4972);
nand UO_100 (O_100,N_4994,N_4887);
or UO_101 (O_101,N_4879,N_4858);
nor UO_102 (O_102,N_4978,N_4948);
nor UO_103 (O_103,N_4989,N_4911);
or UO_104 (O_104,N_4960,N_4847);
and UO_105 (O_105,N_4984,N_4855);
or UO_106 (O_106,N_4862,N_4894);
xor UO_107 (O_107,N_4825,N_4888);
xnor UO_108 (O_108,N_4951,N_4927);
nor UO_109 (O_109,N_4872,N_4992);
xor UO_110 (O_110,N_4960,N_4946);
nor UO_111 (O_111,N_4840,N_4983);
nand UO_112 (O_112,N_4977,N_4937);
nand UO_113 (O_113,N_4867,N_4817);
xor UO_114 (O_114,N_4944,N_4823);
nor UO_115 (O_115,N_4936,N_4905);
nand UO_116 (O_116,N_4859,N_4998);
or UO_117 (O_117,N_4945,N_4975);
nand UO_118 (O_118,N_4959,N_4998);
or UO_119 (O_119,N_4802,N_4904);
or UO_120 (O_120,N_4830,N_4847);
nand UO_121 (O_121,N_4816,N_4832);
and UO_122 (O_122,N_4833,N_4815);
nand UO_123 (O_123,N_4929,N_4926);
xor UO_124 (O_124,N_4931,N_4812);
and UO_125 (O_125,N_4898,N_4813);
or UO_126 (O_126,N_4938,N_4829);
nor UO_127 (O_127,N_4944,N_4969);
nor UO_128 (O_128,N_4841,N_4984);
or UO_129 (O_129,N_4893,N_4800);
nor UO_130 (O_130,N_4980,N_4890);
or UO_131 (O_131,N_4915,N_4837);
nor UO_132 (O_132,N_4849,N_4874);
nand UO_133 (O_133,N_4908,N_4970);
or UO_134 (O_134,N_4913,N_4849);
and UO_135 (O_135,N_4933,N_4993);
nand UO_136 (O_136,N_4948,N_4971);
and UO_137 (O_137,N_4932,N_4889);
nor UO_138 (O_138,N_4827,N_4993);
or UO_139 (O_139,N_4930,N_4927);
nand UO_140 (O_140,N_4974,N_4978);
or UO_141 (O_141,N_4929,N_4853);
or UO_142 (O_142,N_4807,N_4937);
or UO_143 (O_143,N_4856,N_4874);
or UO_144 (O_144,N_4912,N_4928);
or UO_145 (O_145,N_4958,N_4997);
nor UO_146 (O_146,N_4922,N_4841);
nand UO_147 (O_147,N_4995,N_4947);
nand UO_148 (O_148,N_4899,N_4912);
nor UO_149 (O_149,N_4865,N_4990);
and UO_150 (O_150,N_4938,N_4988);
nand UO_151 (O_151,N_4817,N_4908);
and UO_152 (O_152,N_4814,N_4985);
or UO_153 (O_153,N_4981,N_4813);
nor UO_154 (O_154,N_4876,N_4971);
nor UO_155 (O_155,N_4984,N_4898);
nor UO_156 (O_156,N_4924,N_4947);
nand UO_157 (O_157,N_4872,N_4804);
nand UO_158 (O_158,N_4897,N_4983);
nand UO_159 (O_159,N_4833,N_4931);
nand UO_160 (O_160,N_4912,N_4955);
nand UO_161 (O_161,N_4892,N_4888);
nand UO_162 (O_162,N_4917,N_4878);
nor UO_163 (O_163,N_4939,N_4828);
and UO_164 (O_164,N_4954,N_4825);
nor UO_165 (O_165,N_4858,N_4827);
nand UO_166 (O_166,N_4816,N_4950);
nor UO_167 (O_167,N_4906,N_4875);
nor UO_168 (O_168,N_4824,N_4871);
or UO_169 (O_169,N_4860,N_4899);
nand UO_170 (O_170,N_4878,N_4909);
and UO_171 (O_171,N_4973,N_4971);
nand UO_172 (O_172,N_4938,N_4856);
nand UO_173 (O_173,N_4998,N_4962);
or UO_174 (O_174,N_4882,N_4899);
and UO_175 (O_175,N_4976,N_4806);
nand UO_176 (O_176,N_4894,N_4916);
or UO_177 (O_177,N_4988,N_4829);
nand UO_178 (O_178,N_4834,N_4938);
nor UO_179 (O_179,N_4992,N_4919);
or UO_180 (O_180,N_4802,N_4818);
or UO_181 (O_181,N_4840,N_4914);
xnor UO_182 (O_182,N_4909,N_4973);
nor UO_183 (O_183,N_4815,N_4910);
or UO_184 (O_184,N_4953,N_4836);
and UO_185 (O_185,N_4954,N_4881);
or UO_186 (O_186,N_4810,N_4838);
or UO_187 (O_187,N_4831,N_4926);
and UO_188 (O_188,N_4871,N_4893);
or UO_189 (O_189,N_4893,N_4846);
nand UO_190 (O_190,N_4949,N_4809);
and UO_191 (O_191,N_4802,N_4826);
xor UO_192 (O_192,N_4853,N_4935);
nand UO_193 (O_193,N_4970,N_4870);
nor UO_194 (O_194,N_4956,N_4843);
nand UO_195 (O_195,N_4932,N_4833);
nor UO_196 (O_196,N_4813,N_4858);
nor UO_197 (O_197,N_4914,N_4856);
nor UO_198 (O_198,N_4871,N_4887);
nand UO_199 (O_199,N_4827,N_4937);
nand UO_200 (O_200,N_4972,N_4935);
nor UO_201 (O_201,N_4942,N_4998);
nand UO_202 (O_202,N_4931,N_4915);
nand UO_203 (O_203,N_4874,N_4840);
or UO_204 (O_204,N_4883,N_4864);
and UO_205 (O_205,N_4838,N_4845);
xor UO_206 (O_206,N_4917,N_4857);
nor UO_207 (O_207,N_4824,N_4881);
or UO_208 (O_208,N_4889,N_4800);
nand UO_209 (O_209,N_4886,N_4893);
or UO_210 (O_210,N_4972,N_4954);
nand UO_211 (O_211,N_4882,N_4890);
nand UO_212 (O_212,N_4914,N_4868);
xor UO_213 (O_213,N_4937,N_4983);
and UO_214 (O_214,N_4937,N_4861);
or UO_215 (O_215,N_4922,N_4929);
or UO_216 (O_216,N_4928,N_4801);
and UO_217 (O_217,N_4925,N_4906);
or UO_218 (O_218,N_4961,N_4944);
xor UO_219 (O_219,N_4959,N_4856);
and UO_220 (O_220,N_4816,N_4873);
or UO_221 (O_221,N_4880,N_4941);
or UO_222 (O_222,N_4985,N_4823);
nand UO_223 (O_223,N_4835,N_4900);
or UO_224 (O_224,N_4895,N_4898);
and UO_225 (O_225,N_4824,N_4982);
nor UO_226 (O_226,N_4995,N_4937);
nand UO_227 (O_227,N_4879,N_4893);
nor UO_228 (O_228,N_4912,N_4917);
nand UO_229 (O_229,N_4918,N_4929);
or UO_230 (O_230,N_4910,N_4873);
and UO_231 (O_231,N_4929,N_4849);
nand UO_232 (O_232,N_4827,N_4818);
nor UO_233 (O_233,N_4903,N_4983);
or UO_234 (O_234,N_4951,N_4964);
nor UO_235 (O_235,N_4867,N_4964);
and UO_236 (O_236,N_4908,N_4900);
or UO_237 (O_237,N_4859,N_4922);
and UO_238 (O_238,N_4887,N_4972);
nand UO_239 (O_239,N_4947,N_4976);
and UO_240 (O_240,N_4951,N_4868);
or UO_241 (O_241,N_4868,N_4830);
and UO_242 (O_242,N_4963,N_4979);
nand UO_243 (O_243,N_4827,N_4891);
or UO_244 (O_244,N_4814,N_4854);
xor UO_245 (O_245,N_4943,N_4873);
or UO_246 (O_246,N_4945,N_4901);
nand UO_247 (O_247,N_4958,N_4908);
and UO_248 (O_248,N_4936,N_4857);
nor UO_249 (O_249,N_4919,N_4988);
and UO_250 (O_250,N_4893,N_4801);
nor UO_251 (O_251,N_4972,N_4965);
or UO_252 (O_252,N_4977,N_4818);
or UO_253 (O_253,N_4885,N_4887);
and UO_254 (O_254,N_4940,N_4826);
and UO_255 (O_255,N_4918,N_4899);
and UO_256 (O_256,N_4984,N_4818);
nor UO_257 (O_257,N_4904,N_4983);
nor UO_258 (O_258,N_4830,N_4826);
or UO_259 (O_259,N_4988,N_4989);
or UO_260 (O_260,N_4821,N_4949);
nand UO_261 (O_261,N_4816,N_4895);
or UO_262 (O_262,N_4806,N_4913);
xor UO_263 (O_263,N_4847,N_4878);
nor UO_264 (O_264,N_4882,N_4802);
or UO_265 (O_265,N_4962,N_4862);
nand UO_266 (O_266,N_4826,N_4967);
nand UO_267 (O_267,N_4909,N_4858);
or UO_268 (O_268,N_4873,N_4826);
and UO_269 (O_269,N_4971,N_4950);
nand UO_270 (O_270,N_4983,N_4915);
nor UO_271 (O_271,N_4892,N_4878);
nor UO_272 (O_272,N_4919,N_4948);
and UO_273 (O_273,N_4841,N_4889);
nor UO_274 (O_274,N_4842,N_4829);
nand UO_275 (O_275,N_4903,N_4833);
and UO_276 (O_276,N_4934,N_4875);
nand UO_277 (O_277,N_4932,N_4893);
xor UO_278 (O_278,N_4959,N_4874);
nand UO_279 (O_279,N_4883,N_4870);
nor UO_280 (O_280,N_4979,N_4901);
nor UO_281 (O_281,N_4805,N_4920);
or UO_282 (O_282,N_4941,N_4898);
and UO_283 (O_283,N_4812,N_4815);
or UO_284 (O_284,N_4890,N_4866);
nor UO_285 (O_285,N_4966,N_4915);
or UO_286 (O_286,N_4824,N_4819);
nand UO_287 (O_287,N_4951,N_4961);
and UO_288 (O_288,N_4858,N_4973);
and UO_289 (O_289,N_4922,N_4924);
and UO_290 (O_290,N_4821,N_4864);
nor UO_291 (O_291,N_4849,N_4911);
nand UO_292 (O_292,N_4885,N_4870);
nor UO_293 (O_293,N_4836,N_4972);
and UO_294 (O_294,N_4936,N_4822);
nand UO_295 (O_295,N_4830,N_4861);
nand UO_296 (O_296,N_4874,N_4860);
nor UO_297 (O_297,N_4917,N_4979);
and UO_298 (O_298,N_4806,N_4980);
nand UO_299 (O_299,N_4868,N_4877);
nor UO_300 (O_300,N_4844,N_4944);
nor UO_301 (O_301,N_4849,N_4841);
or UO_302 (O_302,N_4975,N_4839);
nor UO_303 (O_303,N_4838,N_4818);
nor UO_304 (O_304,N_4847,N_4889);
and UO_305 (O_305,N_4832,N_4913);
nor UO_306 (O_306,N_4987,N_4850);
or UO_307 (O_307,N_4853,N_4997);
and UO_308 (O_308,N_4880,N_4966);
or UO_309 (O_309,N_4829,N_4991);
and UO_310 (O_310,N_4857,N_4912);
nand UO_311 (O_311,N_4819,N_4890);
and UO_312 (O_312,N_4830,N_4910);
xnor UO_313 (O_313,N_4967,N_4912);
nand UO_314 (O_314,N_4878,N_4829);
or UO_315 (O_315,N_4858,N_4960);
xor UO_316 (O_316,N_4824,N_4802);
or UO_317 (O_317,N_4969,N_4806);
or UO_318 (O_318,N_4929,N_4823);
nand UO_319 (O_319,N_4977,N_4884);
and UO_320 (O_320,N_4836,N_4868);
and UO_321 (O_321,N_4977,N_4869);
xnor UO_322 (O_322,N_4879,N_4975);
nor UO_323 (O_323,N_4814,N_4941);
nand UO_324 (O_324,N_4850,N_4817);
nand UO_325 (O_325,N_4892,N_4862);
and UO_326 (O_326,N_4963,N_4801);
and UO_327 (O_327,N_4865,N_4868);
and UO_328 (O_328,N_4979,N_4964);
nor UO_329 (O_329,N_4914,N_4983);
or UO_330 (O_330,N_4913,N_4902);
and UO_331 (O_331,N_4889,N_4931);
nor UO_332 (O_332,N_4975,N_4859);
nand UO_333 (O_333,N_4926,N_4974);
nor UO_334 (O_334,N_4918,N_4969);
and UO_335 (O_335,N_4928,N_4826);
and UO_336 (O_336,N_4878,N_4879);
nand UO_337 (O_337,N_4861,N_4973);
nor UO_338 (O_338,N_4944,N_4841);
nand UO_339 (O_339,N_4891,N_4866);
and UO_340 (O_340,N_4932,N_4896);
and UO_341 (O_341,N_4837,N_4937);
xnor UO_342 (O_342,N_4834,N_4974);
or UO_343 (O_343,N_4992,N_4959);
and UO_344 (O_344,N_4945,N_4848);
nand UO_345 (O_345,N_4810,N_4852);
nor UO_346 (O_346,N_4980,N_4963);
and UO_347 (O_347,N_4958,N_4816);
and UO_348 (O_348,N_4986,N_4810);
and UO_349 (O_349,N_4982,N_4817);
or UO_350 (O_350,N_4853,N_4963);
nor UO_351 (O_351,N_4987,N_4873);
or UO_352 (O_352,N_4939,N_4917);
nand UO_353 (O_353,N_4950,N_4866);
and UO_354 (O_354,N_4975,N_4914);
or UO_355 (O_355,N_4947,N_4816);
nor UO_356 (O_356,N_4914,N_4978);
xor UO_357 (O_357,N_4907,N_4824);
nand UO_358 (O_358,N_4943,N_4894);
or UO_359 (O_359,N_4953,N_4862);
or UO_360 (O_360,N_4885,N_4926);
nor UO_361 (O_361,N_4882,N_4841);
nand UO_362 (O_362,N_4814,N_4871);
xnor UO_363 (O_363,N_4875,N_4971);
nand UO_364 (O_364,N_4997,N_4900);
and UO_365 (O_365,N_4906,N_4881);
nor UO_366 (O_366,N_4967,N_4980);
and UO_367 (O_367,N_4967,N_4844);
and UO_368 (O_368,N_4857,N_4812);
xor UO_369 (O_369,N_4805,N_4807);
xnor UO_370 (O_370,N_4894,N_4905);
nand UO_371 (O_371,N_4973,N_4820);
nor UO_372 (O_372,N_4968,N_4926);
or UO_373 (O_373,N_4872,N_4917);
and UO_374 (O_374,N_4878,N_4854);
xnor UO_375 (O_375,N_4970,N_4883);
or UO_376 (O_376,N_4966,N_4968);
or UO_377 (O_377,N_4959,N_4818);
or UO_378 (O_378,N_4814,N_4956);
or UO_379 (O_379,N_4911,N_4865);
nand UO_380 (O_380,N_4889,N_4974);
nand UO_381 (O_381,N_4824,N_4854);
and UO_382 (O_382,N_4867,N_4888);
or UO_383 (O_383,N_4820,N_4900);
and UO_384 (O_384,N_4947,N_4971);
xor UO_385 (O_385,N_4963,N_4873);
nor UO_386 (O_386,N_4988,N_4846);
or UO_387 (O_387,N_4842,N_4819);
nor UO_388 (O_388,N_4972,N_4971);
nand UO_389 (O_389,N_4810,N_4851);
and UO_390 (O_390,N_4993,N_4918);
or UO_391 (O_391,N_4863,N_4936);
nor UO_392 (O_392,N_4900,N_4839);
or UO_393 (O_393,N_4901,N_4875);
nand UO_394 (O_394,N_4815,N_4929);
nand UO_395 (O_395,N_4823,N_4973);
nand UO_396 (O_396,N_4839,N_4989);
xor UO_397 (O_397,N_4893,N_4847);
and UO_398 (O_398,N_4930,N_4858);
xor UO_399 (O_399,N_4963,N_4915);
nand UO_400 (O_400,N_4976,N_4998);
or UO_401 (O_401,N_4902,N_4917);
nand UO_402 (O_402,N_4986,N_4922);
or UO_403 (O_403,N_4919,N_4862);
and UO_404 (O_404,N_4895,N_4837);
nand UO_405 (O_405,N_4948,N_4853);
or UO_406 (O_406,N_4918,N_4852);
and UO_407 (O_407,N_4972,N_4823);
and UO_408 (O_408,N_4974,N_4821);
nor UO_409 (O_409,N_4930,N_4899);
nor UO_410 (O_410,N_4849,N_4960);
or UO_411 (O_411,N_4987,N_4825);
or UO_412 (O_412,N_4989,N_4959);
nand UO_413 (O_413,N_4895,N_4825);
nand UO_414 (O_414,N_4948,N_4964);
or UO_415 (O_415,N_4943,N_4868);
and UO_416 (O_416,N_4980,N_4995);
or UO_417 (O_417,N_4942,N_4967);
and UO_418 (O_418,N_4920,N_4808);
or UO_419 (O_419,N_4988,N_4960);
and UO_420 (O_420,N_4841,N_4976);
nand UO_421 (O_421,N_4913,N_4921);
nand UO_422 (O_422,N_4870,N_4835);
or UO_423 (O_423,N_4858,N_4840);
nand UO_424 (O_424,N_4887,N_4971);
or UO_425 (O_425,N_4810,N_4925);
nand UO_426 (O_426,N_4882,N_4931);
nand UO_427 (O_427,N_4924,N_4823);
or UO_428 (O_428,N_4985,N_4878);
nor UO_429 (O_429,N_4830,N_4860);
or UO_430 (O_430,N_4983,N_4860);
xor UO_431 (O_431,N_4985,N_4868);
nor UO_432 (O_432,N_4812,N_4818);
or UO_433 (O_433,N_4965,N_4987);
and UO_434 (O_434,N_4965,N_4833);
or UO_435 (O_435,N_4844,N_4949);
nor UO_436 (O_436,N_4993,N_4927);
and UO_437 (O_437,N_4945,N_4928);
nor UO_438 (O_438,N_4819,N_4910);
xnor UO_439 (O_439,N_4857,N_4937);
nand UO_440 (O_440,N_4951,N_4944);
xor UO_441 (O_441,N_4801,N_4823);
nand UO_442 (O_442,N_4982,N_4892);
xor UO_443 (O_443,N_4898,N_4986);
nand UO_444 (O_444,N_4901,N_4908);
and UO_445 (O_445,N_4973,N_4988);
or UO_446 (O_446,N_4864,N_4887);
nand UO_447 (O_447,N_4973,N_4991);
nand UO_448 (O_448,N_4999,N_4978);
nor UO_449 (O_449,N_4855,N_4831);
nand UO_450 (O_450,N_4896,N_4834);
nand UO_451 (O_451,N_4825,N_4810);
nor UO_452 (O_452,N_4929,N_4870);
or UO_453 (O_453,N_4807,N_4834);
and UO_454 (O_454,N_4915,N_4808);
or UO_455 (O_455,N_4946,N_4987);
and UO_456 (O_456,N_4942,N_4886);
nor UO_457 (O_457,N_4975,N_4994);
nor UO_458 (O_458,N_4916,N_4819);
and UO_459 (O_459,N_4979,N_4992);
nor UO_460 (O_460,N_4866,N_4807);
or UO_461 (O_461,N_4918,N_4990);
or UO_462 (O_462,N_4896,N_4900);
and UO_463 (O_463,N_4938,N_4893);
or UO_464 (O_464,N_4979,N_4944);
or UO_465 (O_465,N_4926,N_4835);
xnor UO_466 (O_466,N_4884,N_4957);
and UO_467 (O_467,N_4963,N_4957);
and UO_468 (O_468,N_4822,N_4925);
or UO_469 (O_469,N_4967,N_4806);
nand UO_470 (O_470,N_4881,N_4909);
nand UO_471 (O_471,N_4800,N_4971);
or UO_472 (O_472,N_4853,N_4824);
or UO_473 (O_473,N_4887,N_4862);
nor UO_474 (O_474,N_4853,N_4945);
and UO_475 (O_475,N_4800,N_4970);
nor UO_476 (O_476,N_4912,N_4869);
and UO_477 (O_477,N_4860,N_4999);
xnor UO_478 (O_478,N_4807,N_4924);
and UO_479 (O_479,N_4826,N_4958);
or UO_480 (O_480,N_4965,N_4804);
nand UO_481 (O_481,N_4838,N_4974);
nor UO_482 (O_482,N_4848,N_4917);
xnor UO_483 (O_483,N_4954,N_4818);
xor UO_484 (O_484,N_4970,N_4967);
nand UO_485 (O_485,N_4940,N_4996);
nor UO_486 (O_486,N_4827,N_4913);
and UO_487 (O_487,N_4834,N_4847);
or UO_488 (O_488,N_4855,N_4883);
nand UO_489 (O_489,N_4977,N_4914);
nand UO_490 (O_490,N_4848,N_4832);
nor UO_491 (O_491,N_4996,N_4910);
and UO_492 (O_492,N_4912,N_4831);
nor UO_493 (O_493,N_4884,N_4954);
and UO_494 (O_494,N_4872,N_4842);
nor UO_495 (O_495,N_4856,N_4953);
nor UO_496 (O_496,N_4882,N_4804);
or UO_497 (O_497,N_4938,N_4892);
or UO_498 (O_498,N_4946,N_4970);
or UO_499 (O_499,N_4886,N_4960);
or UO_500 (O_500,N_4939,N_4958);
nand UO_501 (O_501,N_4833,N_4941);
nor UO_502 (O_502,N_4965,N_4840);
xor UO_503 (O_503,N_4914,N_4812);
and UO_504 (O_504,N_4819,N_4802);
or UO_505 (O_505,N_4954,N_4976);
and UO_506 (O_506,N_4914,N_4851);
nor UO_507 (O_507,N_4972,N_4834);
and UO_508 (O_508,N_4954,N_4955);
nand UO_509 (O_509,N_4862,N_4847);
or UO_510 (O_510,N_4873,N_4957);
nand UO_511 (O_511,N_4916,N_4990);
nor UO_512 (O_512,N_4937,N_4930);
nand UO_513 (O_513,N_4964,N_4802);
nand UO_514 (O_514,N_4906,N_4917);
and UO_515 (O_515,N_4959,N_4854);
nand UO_516 (O_516,N_4818,N_4951);
nand UO_517 (O_517,N_4911,N_4803);
and UO_518 (O_518,N_4819,N_4817);
nand UO_519 (O_519,N_4987,N_4881);
or UO_520 (O_520,N_4828,N_4879);
xnor UO_521 (O_521,N_4819,N_4874);
or UO_522 (O_522,N_4920,N_4883);
or UO_523 (O_523,N_4907,N_4982);
or UO_524 (O_524,N_4915,N_4932);
or UO_525 (O_525,N_4888,N_4826);
and UO_526 (O_526,N_4939,N_4818);
or UO_527 (O_527,N_4951,N_4939);
nor UO_528 (O_528,N_4846,N_4872);
nand UO_529 (O_529,N_4945,N_4973);
nor UO_530 (O_530,N_4904,N_4944);
nand UO_531 (O_531,N_4972,N_4973);
nor UO_532 (O_532,N_4844,N_4883);
and UO_533 (O_533,N_4930,N_4850);
nand UO_534 (O_534,N_4827,N_4996);
or UO_535 (O_535,N_4964,N_4842);
nand UO_536 (O_536,N_4871,N_4936);
nand UO_537 (O_537,N_4968,N_4855);
xor UO_538 (O_538,N_4912,N_4904);
and UO_539 (O_539,N_4975,N_4974);
xnor UO_540 (O_540,N_4869,N_4984);
nand UO_541 (O_541,N_4981,N_4851);
and UO_542 (O_542,N_4834,N_4983);
nor UO_543 (O_543,N_4884,N_4944);
nor UO_544 (O_544,N_4801,N_4955);
and UO_545 (O_545,N_4926,N_4873);
or UO_546 (O_546,N_4976,N_4823);
and UO_547 (O_547,N_4863,N_4829);
nand UO_548 (O_548,N_4899,N_4909);
nor UO_549 (O_549,N_4997,N_4830);
or UO_550 (O_550,N_4803,N_4892);
and UO_551 (O_551,N_4904,N_4892);
nand UO_552 (O_552,N_4968,N_4835);
or UO_553 (O_553,N_4830,N_4835);
nand UO_554 (O_554,N_4979,N_4878);
nor UO_555 (O_555,N_4905,N_4928);
or UO_556 (O_556,N_4872,N_4900);
nand UO_557 (O_557,N_4849,N_4992);
or UO_558 (O_558,N_4980,N_4924);
nand UO_559 (O_559,N_4804,N_4888);
or UO_560 (O_560,N_4904,N_4952);
or UO_561 (O_561,N_4937,N_4815);
and UO_562 (O_562,N_4840,N_4938);
xnor UO_563 (O_563,N_4850,N_4857);
nor UO_564 (O_564,N_4909,N_4931);
or UO_565 (O_565,N_4975,N_4986);
or UO_566 (O_566,N_4898,N_4881);
nor UO_567 (O_567,N_4915,N_4959);
and UO_568 (O_568,N_4821,N_4882);
nand UO_569 (O_569,N_4970,N_4937);
and UO_570 (O_570,N_4893,N_4906);
xor UO_571 (O_571,N_4858,N_4819);
or UO_572 (O_572,N_4840,N_4986);
nor UO_573 (O_573,N_4841,N_4817);
and UO_574 (O_574,N_4906,N_4829);
or UO_575 (O_575,N_4819,N_4866);
and UO_576 (O_576,N_4951,N_4943);
nand UO_577 (O_577,N_4904,N_4888);
nand UO_578 (O_578,N_4896,N_4830);
nor UO_579 (O_579,N_4879,N_4921);
and UO_580 (O_580,N_4930,N_4886);
and UO_581 (O_581,N_4896,N_4962);
nand UO_582 (O_582,N_4828,N_4846);
nand UO_583 (O_583,N_4860,N_4801);
or UO_584 (O_584,N_4829,N_4861);
nand UO_585 (O_585,N_4883,N_4826);
or UO_586 (O_586,N_4809,N_4864);
nand UO_587 (O_587,N_4855,N_4820);
nand UO_588 (O_588,N_4912,N_4833);
xnor UO_589 (O_589,N_4981,N_4807);
nor UO_590 (O_590,N_4835,N_4851);
nand UO_591 (O_591,N_4853,N_4827);
nand UO_592 (O_592,N_4871,N_4984);
and UO_593 (O_593,N_4941,N_4984);
nand UO_594 (O_594,N_4923,N_4850);
and UO_595 (O_595,N_4839,N_4866);
and UO_596 (O_596,N_4820,N_4847);
or UO_597 (O_597,N_4896,N_4996);
or UO_598 (O_598,N_4915,N_4961);
nand UO_599 (O_599,N_4982,N_4917);
xnor UO_600 (O_600,N_4869,N_4887);
nand UO_601 (O_601,N_4955,N_4953);
and UO_602 (O_602,N_4812,N_4840);
and UO_603 (O_603,N_4902,N_4824);
nand UO_604 (O_604,N_4801,N_4910);
nor UO_605 (O_605,N_4880,N_4864);
and UO_606 (O_606,N_4901,N_4808);
nand UO_607 (O_607,N_4863,N_4877);
and UO_608 (O_608,N_4846,N_4907);
nand UO_609 (O_609,N_4921,N_4856);
or UO_610 (O_610,N_4821,N_4991);
nand UO_611 (O_611,N_4983,N_4991);
and UO_612 (O_612,N_4846,N_4878);
nor UO_613 (O_613,N_4806,N_4919);
or UO_614 (O_614,N_4938,N_4823);
and UO_615 (O_615,N_4872,N_4897);
nand UO_616 (O_616,N_4918,N_4823);
xnor UO_617 (O_617,N_4853,N_4966);
or UO_618 (O_618,N_4815,N_4950);
or UO_619 (O_619,N_4958,N_4850);
or UO_620 (O_620,N_4879,N_4968);
nor UO_621 (O_621,N_4812,N_4839);
nor UO_622 (O_622,N_4912,N_4888);
or UO_623 (O_623,N_4872,N_4990);
and UO_624 (O_624,N_4883,N_4984);
nor UO_625 (O_625,N_4892,N_4830);
nor UO_626 (O_626,N_4805,N_4921);
xnor UO_627 (O_627,N_4957,N_4942);
xor UO_628 (O_628,N_4902,N_4872);
nor UO_629 (O_629,N_4984,N_4908);
nor UO_630 (O_630,N_4984,N_4987);
or UO_631 (O_631,N_4988,N_4954);
nor UO_632 (O_632,N_4845,N_4988);
or UO_633 (O_633,N_4920,N_4904);
nand UO_634 (O_634,N_4895,N_4887);
or UO_635 (O_635,N_4938,N_4996);
xor UO_636 (O_636,N_4907,N_4916);
or UO_637 (O_637,N_4899,N_4891);
nand UO_638 (O_638,N_4860,N_4826);
xnor UO_639 (O_639,N_4999,N_4881);
nor UO_640 (O_640,N_4900,N_4892);
and UO_641 (O_641,N_4868,N_4883);
or UO_642 (O_642,N_4970,N_4933);
nand UO_643 (O_643,N_4891,N_4859);
and UO_644 (O_644,N_4827,N_4941);
xor UO_645 (O_645,N_4862,N_4844);
nor UO_646 (O_646,N_4915,N_4842);
and UO_647 (O_647,N_4960,N_4834);
nor UO_648 (O_648,N_4979,N_4981);
nor UO_649 (O_649,N_4843,N_4973);
and UO_650 (O_650,N_4844,N_4881);
nor UO_651 (O_651,N_4916,N_4912);
or UO_652 (O_652,N_4968,N_4832);
xnor UO_653 (O_653,N_4868,N_4850);
or UO_654 (O_654,N_4939,N_4843);
and UO_655 (O_655,N_4950,N_4999);
or UO_656 (O_656,N_4844,N_4907);
xor UO_657 (O_657,N_4860,N_4949);
xnor UO_658 (O_658,N_4881,N_4921);
nor UO_659 (O_659,N_4830,N_4924);
and UO_660 (O_660,N_4830,N_4972);
and UO_661 (O_661,N_4949,N_4934);
or UO_662 (O_662,N_4978,N_4805);
nor UO_663 (O_663,N_4992,N_4936);
nor UO_664 (O_664,N_4810,N_4862);
and UO_665 (O_665,N_4955,N_4924);
nand UO_666 (O_666,N_4915,N_4935);
xor UO_667 (O_667,N_4857,N_4886);
nor UO_668 (O_668,N_4936,N_4907);
and UO_669 (O_669,N_4911,N_4984);
nand UO_670 (O_670,N_4980,N_4880);
nand UO_671 (O_671,N_4865,N_4851);
and UO_672 (O_672,N_4944,N_4882);
and UO_673 (O_673,N_4926,N_4844);
and UO_674 (O_674,N_4975,N_4875);
nor UO_675 (O_675,N_4969,N_4832);
xnor UO_676 (O_676,N_4816,N_4831);
and UO_677 (O_677,N_4887,N_4955);
nand UO_678 (O_678,N_4854,N_4800);
or UO_679 (O_679,N_4832,N_4907);
or UO_680 (O_680,N_4938,N_4965);
and UO_681 (O_681,N_4806,N_4954);
or UO_682 (O_682,N_4881,N_4943);
nor UO_683 (O_683,N_4887,N_4897);
xnor UO_684 (O_684,N_4905,N_4912);
nor UO_685 (O_685,N_4850,N_4882);
nand UO_686 (O_686,N_4814,N_4816);
nand UO_687 (O_687,N_4984,N_4980);
and UO_688 (O_688,N_4940,N_4832);
or UO_689 (O_689,N_4951,N_4984);
nor UO_690 (O_690,N_4964,N_4993);
and UO_691 (O_691,N_4877,N_4906);
or UO_692 (O_692,N_4831,N_4911);
nand UO_693 (O_693,N_4941,N_4852);
or UO_694 (O_694,N_4801,N_4810);
and UO_695 (O_695,N_4947,N_4999);
and UO_696 (O_696,N_4872,N_4820);
or UO_697 (O_697,N_4886,N_4999);
nand UO_698 (O_698,N_4983,N_4960);
nand UO_699 (O_699,N_4942,N_4904);
xnor UO_700 (O_700,N_4835,N_4981);
or UO_701 (O_701,N_4925,N_4893);
and UO_702 (O_702,N_4849,N_4816);
and UO_703 (O_703,N_4860,N_4867);
and UO_704 (O_704,N_4905,N_4840);
or UO_705 (O_705,N_4900,N_4957);
and UO_706 (O_706,N_4963,N_4897);
nand UO_707 (O_707,N_4816,N_4982);
nand UO_708 (O_708,N_4824,N_4815);
xnor UO_709 (O_709,N_4945,N_4963);
nand UO_710 (O_710,N_4812,N_4897);
xor UO_711 (O_711,N_4870,N_4892);
and UO_712 (O_712,N_4925,N_4828);
and UO_713 (O_713,N_4802,N_4811);
and UO_714 (O_714,N_4995,N_4800);
nand UO_715 (O_715,N_4871,N_4905);
nand UO_716 (O_716,N_4864,N_4800);
or UO_717 (O_717,N_4848,N_4889);
xnor UO_718 (O_718,N_4906,N_4846);
and UO_719 (O_719,N_4968,N_4823);
and UO_720 (O_720,N_4810,N_4908);
or UO_721 (O_721,N_4965,N_4883);
nand UO_722 (O_722,N_4889,N_4992);
or UO_723 (O_723,N_4820,N_4806);
and UO_724 (O_724,N_4961,N_4959);
and UO_725 (O_725,N_4999,N_4889);
and UO_726 (O_726,N_4817,N_4959);
or UO_727 (O_727,N_4828,N_4979);
nand UO_728 (O_728,N_4819,N_4886);
xor UO_729 (O_729,N_4896,N_4886);
nor UO_730 (O_730,N_4897,N_4883);
or UO_731 (O_731,N_4958,N_4992);
nand UO_732 (O_732,N_4898,N_4951);
and UO_733 (O_733,N_4858,N_4820);
nor UO_734 (O_734,N_4997,N_4991);
and UO_735 (O_735,N_4846,N_4865);
and UO_736 (O_736,N_4839,N_4873);
and UO_737 (O_737,N_4811,N_4861);
or UO_738 (O_738,N_4937,N_4891);
nand UO_739 (O_739,N_4955,N_4921);
nand UO_740 (O_740,N_4981,N_4867);
nor UO_741 (O_741,N_4816,N_4912);
nand UO_742 (O_742,N_4885,N_4803);
or UO_743 (O_743,N_4937,N_4940);
nand UO_744 (O_744,N_4902,N_4986);
nor UO_745 (O_745,N_4984,N_4804);
xnor UO_746 (O_746,N_4823,N_4821);
and UO_747 (O_747,N_4991,N_4809);
and UO_748 (O_748,N_4872,N_4918);
nor UO_749 (O_749,N_4839,N_4874);
and UO_750 (O_750,N_4841,N_4906);
or UO_751 (O_751,N_4833,N_4831);
and UO_752 (O_752,N_4804,N_4880);
nand UO_753 (O_753,N_4861,N_4879);
and UO_754 (O_754,N_4876,N_4930);
nor UO_755 (O_755,N_4921,N_4938);
and UO_756 (O_756,N_4816,N_4900);
nor UO_757 (O_757,N_4894,N_4908);
or UO_758 (O_758,N_4904,N_4899);
and UO_759 (O_759,N_4804,N_4810);
and UO_760 (O_760,N_4880,N_4828);
and UO_761 (O_761,N_4870,N_4926);
or UO_762 (O_762,N_4900,N_4966);
nand UO_763 (O_763,N_4949,N_4933);
xor UO_764 (O_764,N_4972,N_4889);
or UO_765 (O_765,N_4807,N_4929);
and UO_766 (O_766,N_4824,N_4961);
and UO_767 (O_767,N_4910,N_4957);
or UO_768 (O_768,N_4957,N_4806);
nor UO_769 (O_769,N_4850,N_4810);
or UO_770 (O_770,N_4935,N_4969);
or UO_771 (O_771,N_4836,N_4932);
nand UO_772 (O_772,N_4952,N_4802);
and UO_773 (O_773,N_4811,N_4940);
nand UO_774 (O_774,N_4823,N_4989);
and UO_775 (O_775,N_4919,N_4822);
and UO_776 (O_776,N_4900,N_4834);
or UO_777 (O_777,N_4981,N_4985);
nor UO_778 (O_778,N_4860,N_4908);
nand UO_779 (O_779,N_4954,N_4897);
nand UO_780 (O_780,N_4901,N_4887);
and UO_781 (O_781,N_4816,N_4930);
nand UO_782 (O_782,N_4896,N_4926);
and UO_783 (O_783,N_4972,N_4816);
or UO_784 (O_784,N_4917,N_4924);
and UO_785 (O_785,N_4965,N_4976);
or UO_786 (O_786,N_4880,N_4810);
or UO_787 (O_787,N_4959,N_4835);
and UO_788 (O_788,N_4942,N_4883);
nand UO_789 (O_789,N_4948,N_4838);
nor UO_790 (O_790,N_4890,N_4902);
xor UO_791 (O_791,N_4985,N_4897);
or UO_792 (O_792,N_4990,N_4984);
or UO_793 (O_793,N_4975,N_4969);
or UO_794 (O_794,N_4833,N_4971);
or UO_795 (O_795,N_4866,N_4885);
nand UO_796 (O_796,N_4980,N_4966);
nand UO_797 (O_797,N_4974,N_4912);
nand UO_798 (O_798,N_4828,N_4981);
nor UO_799 (O_799,N_4911,N_4822);
nand UO_800 (O_800,N_4950,N_4814);
and UO_801 (O_801,N_4879,N_4870);
or UO_802 (O_802,N_4912,N_4924);
xor UO_803 (O_803,N_4987,N_4812);
and UO_804 (O_804,N_4809,N_4822);
xnor UO_805 (O_805,N_4850,N_4906);
xor UO_806 (O_806,N_4987,N_4852);
nand UO_807 (O_807,N_4841,N_4926);
and UO_808 (O_808,N_4851,N_4891);
or UO_809 (O_809,N_4826,N_4984);
or UO_810 (O_810,N_4999,N_4898);
nand UO_811 (O_811,N_4843,N_4979);
nor UO_812 (O_812,N_4845,N_4813);
or UO_813 (O_813,N_4965,N_4827);
and UO_814 (O_814,N_4932,N_4938);
nand UO_815 (O_815,N_4917,N_4897);
nand UO_816 (O_816,N_4884,N_4864);
nor UO_817 (O_817,N_4939,N_4935);
nor UO_818 (O_818,N_4898,N_4802);
or UO_819 (O_819,N_4805,N_4813);
and UO_820 (O_820,N_4830,N_4978);
nand UO_821 (O_821,N_4855,N_4993);
nor UO_822 (O_822,N_4923,N_4910);
or UO_823 (O_823,N_4997,N_4999);
xnor UO_824 (O_824,N_4855,N_4895);
and UO_825 (O_825,N_4904,N_4808);
nand UO_826 (O_826,N_4949,N_4825);
or UO_827 (O_827,N_4920,N_4923);
nor UO_828 (O_828,N_4863,N_4873);
or UO_829 (O_829,N_4947,N_4930);
and UO_830 (O_830,N_4813,N_4871);
nor UO_831 (O_831,N_4829,N_4913);
and UO_832 (O_832,N_4830,N_4862);
and UO_833 (O_833,N_4836,N_4983);
or UO_834 (O_834,N_4953,N_4977);
and UO_835 (O_835,N_4969,N_4991);
or UO_836 (O_836,N_4969,N_4847);
and UO_837 (O_837,N_4826,N_4938);
nand UO_838 (O_838,N_4903,N_4999);
or UO_839 (O_839,N_4861,N_4985);
nand UO_840 (O_840,N_4827,N_4862);
xnor UO_841 (O_841,N_4995,N_4825);
nor UO_842 (O_842,N_4956,N_4819);
nor UO_843 (O_843,N_4933,N_4889);
nor UO_844 (O_844,N_4808,N_4928);
nor UO_845 (O_845,N_4908,N_4867);
and UO_846 (O_846,N_4847,N_4981);
and UO_847 (O_847,N_4834,N_4977);
nor UO_848 (O_848,N_4918,N_4907);
nand UO_849 (O_849,N_4928,N_4880);
or UO_850 (O_850,N_4855,N_4991);
nor UO_851 (O_851,N_4936,N_4969);
or UO_852 (O_852,N_4802,N_4969);
or UO_853 (O_853,N_4951,N_4901);
or UO_854 (O_854,N_4825,N_4920);
nand UO_855 (O_855,N_4971,N_4933);
and UO_856 (O_856,N_4880,N_4803);
and UO_857 (O_857,N_4862,N_4943);
nor UO_858 (O_858,N_4923,N_4835);
nor UO_859 (O_859,N_4873,N_4905);
nand UO_860 (O_860,N_4879,N_4938);
or UO_861 (O_861,N_4959,N_4964);
and UO_862 (O_862,N_4916,N_4843);
nand UO_863 (O_863,N_4852,N_4812);
nor UO_864 (O_864,N_4970,N_4887);
nor UO_865 (O_865,N_4906,N_4979);
or UO_866 (O_866,N_4851,N_4827);
nor UO_867 (O_867,N_4818,N_4875);
nor UO_868 (O_868,N_4926,N_4807);
and UO_869 (O_869,N_4955,N_4985);
nand UO_870 (O_870,N_4895,N_4818);
nor UO_871 (O_871,N_4987,N_4836);
and UO_872 (O_872,N_4902,N_4800);
nor UO_873 (O_873,N_4830,N_4932);
or UO_874 (O_874,N_4833,N_4845);
nand UO_875 (O_875,N_4852,N_4831);
nor UO_876 (O_876,N_4931,N_4860);
xor UO_877 (O_877,N_4843,N_4835);
xnor UO_878 (O_878,N_4848,N_4913);
and UO_879 (O_879,N_4904,N_4853);
and UO_880 (O_880,N_4952,N_4843);
and UO_881 (O_881,N_4823,N_4886);
nand UO_882 (O_882,N_4851,N_4935);
nor UO_883 (O_883,N_4919,N_4885);
nand UO_884 (O_884,N_4945,N_4989);
xor UO_885 (O_885,N_4951,N_4875);
or UO_886 (O_886,N_4924,N_4984);
nand UO_887 (O_887,N_4959,N_4907);
nor UO_888 (O_888,N_4882,N_4855);
nor UO_889 (O_889,N_4922,N_4897);
or UO_890 (O_890,N_4854,N_4950);
and UO_891 (O_891,N_4967,N_4934);
and UO_892 (O_892,N_4855,N_4953);
nand UO_893 (O_893,N_4807,N_4923);
xnor UO_894 (O_894,N_4864,N_4903);
nor UO_895 (O_895,N_4911,N_4842);
nor UO_896 (O_896,N_4960,N_4833);
and UO_897 (O_897,N_4988,N_4975);
or UO_898 (O_898,N_4915,N_4912);
or UO_899 (O_899,N_4849,N_4846);
and UO_900 (O_900,N_4992,N_4978);
nand UO_901 (O_901,N_4955,N_4891);
nand UO_902 (O_902,N_4965,N_4830);
nor UO_903 (O_903,N_4817,N_4949);
nor UO_904 (O_904,N_4841,N_4913);
nand UO_905 (O_905,N_4819,N_4880);
or UO_906 (O_906,N_4843,N_4894);
nand UO_907 (O_907,N_4850,N_4951);
and UO_908 (O_908,N_4964,N_4962);
nor UO_909 (O_909,N_4813,N_4925);
nand UO_910 (O_910,N_4916,N_4928);
and UO_911 (O_911,N_4975,N_4869);
nand UO_912 (O_912,N_4844,N_4810);
nor UO_913 (O_913,N_4918,N_4986);
nand UO_914 (O_914,N_4908,N_4866);
nand UO_915 (O_915,N_4885,N_4978);
nor UO_916 (O_916,N_4956,N_4817);
nor UO_917 (O_917,N_4980,N_4976);
xor UO_918 (O_918,N_4872,N_4921);
xor UO_919 (O_919,N_4819,N_4941);
nand UO_920 (O_920,N_4980,N_4946);
or UO_921 (O_921,N_4973,N_4875);
nand UO_922 (O_922,N_4943,N_4920);
and UO_923 (O_923,N_4936,N_4816);
nor UO_924 (O_924,N_4912,N_4847);
or UO_925 (O_925,N_4876,N_4906);
nor UO_926 (O_926,N_4958,N_4923);
or UO_927 (O_927,N_4869,N_4937);
nor UO_928 (O_928,N_4978,N_4823);
and UO_929 (O_929,N_4816,N_4837);
nor UO_930 (O_930,N_4817,N_4963);
or UO_931 (O_931,N_4859,N_4886);
nor UO_932 (O_932,N_4911,N_4971);
and UO_933 (O_933,N_4977,N_4895);
nor UO_934 (O_934,N_4954,N_4826);
nand UO_935 (O_935,N_4926,N_4979);
nand UO_936 (O_936,N_4951,N_4893);
or UO_937 (O_937,N_4850,N_4824);
or UO_938 (O_938,N_4832,N_4952);
xor UO_939 (O_939,N_4901,N_4856);
and UO_940 (O_940,N_4975,N_4846);
and UO_941 (O_941,N_4908,N_4990);
and UO_942 (O_942,N_4888,N_4910);
or UO_943 (O_943,N_4979,N_4850);
or UO_944 (O_944,N_4809,N_4941);
or UO_945 (O_945,N_4928,N_4825);
and UO_946 (O_946,N_4961,N_4880);
or UO_947 (O_947,N_4812,N_4929);
nor UO_948 (O_948,N_4905,N_4935);
and UO_949 (O_949,N_4941,N_4849);
nor UO_950 (O_950,N_4852,N_4811);
xnor UO_951 (O_951,N_4978,N_4951);
nand UO_952 (O_952,N_4971,N_4970);
and UO_953 (O_953,N_4879,N_4827);
or UO_954 (O_954,N_4908,N_4853);
nor UO_955 (O_955,N_4909,N_4868);
and UO_956 (O_956,N_4959,N_4884);
nand UO_957 (O_957,N_4986,N_4977);
nand UO_958 (O_958,N_4811,N_4943);
xor UO_959 (O_959,N_4999,N_4826);
xor UO_960 (O_960,N_4906,N_4937);
or UO_961 (O_961,N_4859,N_4864);
xor UO_962 (O_962,N_4831,N_4929);
nand UO_963 (O_963,N_4896,N_4893);
nand UO_964 (O_964,N_4883,N_4976);
and UO_965 (O_965,N_4875,N_4916);
and UO_966 (O_966,N_4940,N_4873);
nor UO_967 (O_967,N_4835,N_4956);
and UO_968 (O_968,N_4996,N_4818);
nor UO_969 (O_969,N_4991,N_4880);
nor UO_970 (O_970,N_4916,N_4943);
xnor UO_971 (O_971,N_4971,N_4846);
nor UO_972 (O_972,N_4924,N_4800);
and UO_973 (O_973,N_4805,N_4938);
nor UO_974 (O_974,N_4935,N_4872);
or UO_975 (O_975,N_4982,N_4906);
xor UO_976 (O_976,N_4895,N_4824);
and UO_977 (O_977,N_4819,N_4844);
xor UO_978 (O_978,N_4840,N_4898);
nand UO_979 (O_979,N_4846,N_4899);
or UO_980 (O_980,N_4969,N_4977);
or UO_981 (O_981,N_4855,N_4916);
nand UO_982 (O_982,N_4890,N_4843);
nand UO_983 (O_983,N_4902,N_4972);
nand UO_984 (O_984,N_4845,N_4884);
or UO_985 (O_985,N_4975,N_4930);
and UO_986 (O_986,N_4992,N_4802);
and UO_987 (O_987,N_4837,N_4880);
or UO_988 (O_988,N_4932,N_4936);
nand UO_989 (O_989,N_4986,N_4940);
nand UO_990 (O_990,N_4903,N_4845);
or UO_991 (O_991,N_4825,N_4982);
nor UO_992 (O_992,N_4963,N_4986);
or UO_993 (O_993,N_4877,N_4840);
nor UO_994 (O_994,N_4836,N_4952);
nand UO_995 (O_995,N_4915,N_4997);
nor UO_996 (O_996,N_4895,N_4806);
nor UO_997 (O_997,N_4908,N_4864);
or UO_998 (O_998,N_4942,N_4819);
or UO_999 (O_999,N_4850,N_4843);
endmodule