module basic_500_3000_500_4_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_219,In_86);
xor U1 (N_1,In_170,In_171);
nand U2 (N_2,In_81,In_338);
nor U3 (N_3,In_6,In_388);
xor U4 (N_4,In_372,In_497);
nand U5 (N_5,In_400,In_64);
nand U6 (N_6,In_441,In_138);
nor U7 (N_7,In_387,In_154);
nand U8 (N_8,In_285,In_176);
xor U9 (N_9,In_455,In_325);
or U10 (N_10,In_131,In_365);
and U11 (N_11,In_10,In_8);
or U12 (N_12,In_269,In_357);
nor U13 (N_13,In_286,In_102);
nand U14 (N_14,In_168,In_11);
and U15 (N_15,In_222,In_209);
nor U16 (N_16,In_129,In_311);
nand U17 (N_17,In_144,In_471);
and U18 (N_18,In_345,In_248);
and U19 (N_19,In_386,In_197);
nor U20 (N_20,In_192,In_330);
or U21 (N_21,In_73,In_94);
xnor U22 (N_22,In_57,In_213);
and U23 (N_23,In_373,In_195);
or U24 (N_24,In_243,In_320);
or U25 (N_25,In_297,In_448);
xnor U26 (N_26,In_40,In_169);
xnor U27 (N_27,In_273,In_340);
nor U28 (N_28,In_250,In_165);
nor U29 (N_29,In_278,In_63);
xnor U30 (N_30,In_95,In_415);
or U31 (N_31,In_466,In_424);
or U32 (N_32,In_156,In_324);
or U33 (N_33,In_389,In_290);
xnor U34 (N_34,In_465,In_488);
nand U35 (N_35,In_1,In_299);
xnor U36 (N_36,In_339,In_2);
or U37 (N_37,In_283,In_158);
or U38 (N_38,In_353,In_454);
nand U39 (N_39,In_97,In_118);
nor U40 (N_40,In_348,In_364);
nand U41 (N_41,In_85,In_490);
xnor U42 (N_42,In_337,In_15);
nand U43 (N_43,In_152,In_346);
and U44 (N_44,In_136,In_91);
and U45 (N_45,In_434,In_208);
nor U46 (N_46,In_280,In_382);
and U47 (N_47,In_238,In_287);
or U48 (N_48,In_23,In_361);
or U49 (N_49,In_438,In_240);
nor U50 (N_50,In_89,In_350);
and U51 (N_51,In_113,In_453);
xnor U52 (N_52,In_31,In_431);
nand U53 (N_53,In_189,In_385);
and U54 (N_54,In_360,In_141);
or U55 (N_55,In_482,In_459);
nand U56 (N_56,In_174,In_26);
or U57 (N_57,In_32,In_38);
or U58 (N_58,In_492,In_125);
nor U59 (N_59,In_146,In_318);
nand U60 (N_60,In_225,In_114);
nor U61 (N_61,In_428,In_155);
and U62 (N_62,In_90,In_496);
nand U63 (N_63,In_254,In_202);
xor U64 (N_64,In_39,In_147);
nor U65 (N_65,In_148,In_442);
nor U66 (N_66,In_474,In_47);
nor U67 (N_67,In_145,In_333);
nor U68 (N_68,In_468,In_443);
and U69 (N_69,In_321,In_264);
nand U70 (N_70,In_36,In_51);
nor U71 (N_71,In_205,In_157);
nor U72 (N_72,In_216,In_263);
xor U73 (N_73,In_328,In_368);
or U74 (N_74,In_383,In_7);
nor U75 (N_75,In_93,In_245);
or U76 (N_76,In_162,In_435);
or U77 (N_77,In_25,In_275);
or U78 (N_78,In_303,In_377);
nand U79 (N_79,In_122,In_82);
nand U80 (N_80,In_104,In_288);
xnor U81 (N_81,In_425,In_463);
xor U82 (N_82,In_418,In_249);
nand U83 (N_83,In_449,In_207);
nor U84 (N_84,In_127,In_187);
nand U85 (N_85,In_369,In_326);
or U86 (N_86,In_322,In_67);
nor U87 (N_87,In_109,In_251);
or U88 (N_88,In_87,In_198);
or U89 (N_89,In_394,In_457);
xor U90 (N_90,In_160,In_37);
nand U91 (N_91,In_69,In_88);
xor U92 (N_92,In_83,In_246);
xnor U93 (N_93,In_396,In_317);
nor U94 (N_94,In_21,In_419);
xor U95 (N_95,In_414,In_342);
and U96 (N_96,In_312,In_49);
nand U97 (N_97,In_422,In_413);
or U98 (N_98,In_110,In_301);
xnor U99 (N_99,In_472,In_451);
nor U100 (N_100,In_112,In_117);
and U101 (N_101,In_478,In_105);
and U102 (N_102,In_409,In_267);
or U103 (N_103,In_341,In_226);
xor U104 (N_104,In_257,In_177);
or U105 (N_105,In_116,In_479);
xnor U106 (N_106,In_436,In_65);
xor U107 (N_107,In_352,In_244);
or U108 (N_108,In_355,In_420);
xnor U109 (N_109,In_439,In_61);
or U110 (N_110,In_334,In_16);
and U111 (N_111,In_281,In_60);
and U112 (N_112,In_390,In_447);
xor U113 (N_113,In_62,In_41);
xor U114 (N_114,In_124,In_370);
and U115 (N_115,In_253,In_261);
nand U116 (N_116,In_14,In_193);
nor U117 (N_117,In_430,In_445);
nand U118 (N_118,In_232,In_13);
xnor U119 (N_119,In_315,In_358);
and U120 (N_120,In_467,In_179);
xor U121 (N_121,In_211,In_9);
nor U122 (N_122,In_384,In_234);
or U123 (N_123,In_399,In_48);
nor U124 (N_124,In_164,In_371);
nand U125 (N_125,In_42,In_18);
xor U126 (N_126,In_103,In_456);
and U127 (N_127,In_276,In_221);
nor U128 (N_128,In_450,In_485);
and U129 (N_129,In_293,In_402);
nor U130 (N_130,In_172,In_461);
nor U131 (N_131,In_499,In_247);
and U132 (N_132,In_210,In_231);
nor U133 (N_133,In_282,In_52);
or U134 (N_134,In_423,In_133);
and U135 (N_135,In_200,In_440);
nand U136 (N_136,In_71,In_329);
nand U137 (N_137,In_185,In_421);
and U138 (N_138,In_66,In_199);
and U139 (N_139,In_309,In_188);
and U140 (N_140,In_151,In_397);
and U141 (N_141,In_363,In_217);
nand U142 (N_142,In_433,In_153);
nor U143 (N_143,In_239,In_314);
nand U144 (N_144,In_218,In_374);
nor U145 (N_145,In_405,In_274);
nand U146 (N_146,In_182,In_284);
or U147 (N_147,In_135,In_108);
and U148 (N_148,In_470,In_412);
and U149 (N_149,In_142,In_59);
or U150 (N_150,In_493,In_224);
and U151 (N_151,In_469,In_101);
xnor U152 (N_152,In_120,In_391);
nand U153 (N_153,In_180,In_194);
and U154 (N_154,In_3,In_375);
or U155 (N_155,In_308,In_427);
nand U156 (N_156,In_173,In_491);
and U157 (N_157,In_53,In_143);
nor U158 (N_158,In_34,In_432);
and U159 (N_159,In_178,In_410);
or U160 (N_160,In_483,In_55);
xnor U161 (N_161,In_111,In_305);
nand U162 (N_162,In_163,In_4);
nand U163 (N_163,In_75,In_126);
nand U164 (N_164,In_139,In_296);
and U165 (N_165,In_79,In_395);
xor U166 (N_166,In_304,In_184);
xnor U167 (N_167,In_68,In_356);
and U168 (N_168,In_460,In_130);
and U169 (N_169,In_306,In_429);
nor U170 (N_170,In_476,In_331);
xor U171 (N_171,In_181,In_19);
or U172 (N_172,In_262,In_190);
or U173 (N_173,In_35,In_268);
and U174 (N_174,In_475,In_236);
or U175 (N_175,In_50,In_452);
xor U176 (N_176,In_401,In_323);
nand U177 (N_177,In_140,In_359);
nand U178 (N_178,In_45,In_201);
nand U179 (N_179,In_256,In_367);
nand U180 (N_180,In_327,In_426);
or U181 (N_181,In_332,In_347);
and U182 (N_182,In_313,In_406);
and U183 (N_183,In_242,In_404);
nor U184 (N_184,In_498,In_223);
or U185 (N_185,In_307,In_235);
nand U186 (N_186,In_0,In_310);
xor U187 (N_187,In_149,In_458);
nor U188 (N_188,In_366,In_80);
and U189 (N_189,In_381,In_107);
or U190 (N_190,In_228,In_20);
nor U191 (N_191,In_44,In_408);
and U192 (N_192,In_84,In_183);
nand U193 (N_193,In_398,In_203);
xnor U194 (N_194,In_487,In_335);
xnor U195 (N_195,In_128,In_464);
or U196 (N_196,In_123,In_486);
or U197 (N_197,In_46,In_417);
or U198 (N_198,In_289,In_106);
xnor U199 (N_199,In_255,In_54);
or U200 (N_200,In_56,In_237);
xnor U201 (N_201,In_76,In_252);
and U202 (N_202,In_258,In_379);
and U203 (N_203,In_119,In_494);
or U204 (N_204,In_392,In_477);
or U205 (N_205,In_266,In_351);
xnor U206 (N_206,In_473,In_70);
or U207 (N_207,In_393,In_444);
nand U208 (N_208,In_462,In_206);
and U209 (N_209,In_29,In_298);
and U210 (N_210,In_319,In_437);
or U211 (N_211,In_416,In_362);
or U212 (N_212,In_300,In_166);
xnor U213 (N_213,In_92,In_186);
nand U214 (N_214,In_17,In_354);
and U215 (N_215,In_227,In_411);
or U216 (N_216,In_33,In_272);
nor U217 (N_217,In_196,In_100);
or U218 (N_218,In_380,In_271);
nor U219 (N_219,In_407,In_43);
nand U220 (N_220,In_96,In_220);
nor U221 (N_221,In_233,In_489);
nand U222 (N_222,In_291,In_403);
nand U223 (N_223,In_74,In_167);
and U224 (N_224,In_58,In_24);
nand U225 (N_225,In_77,In_27);
nor U226 (N_226,In_343,In_98);
xor U227 (N_227,In_72,In_12);
and U228 (N_228,In_121,In_265);
or U229 (N_229,In_294,In_191);
or U230 (N_230,In_161,In_99);
nand U231 (N_231,In_5,In_241);
nor U232 (N_232,In_378,In_260);
xnor U233 (N_233,In_349,In_481);
or U234 (N_234,In_484,In_279);
nor U235 (N_235,In_175,In_480);
and U236 (N_236,In_295,In_230);
nand U237 (N_237,In_292,In_316);
nor U238 (N_238,In_446,In_376);
xor U239 (N_239,In_259,In_336);
nor U240 (N_240,In_215,In_214);
nand U241 (N_241,In_302,In_229);
or U242 (N_242,In_204,In_495);
nand U243 (N_243,In_134,In_22);
nor U244 (N_244,In_78,In_150);
and U245 (N_245,In_159,In_132);
and U246 (N_246,In_30,In_270);
or U247 (N_247,In_277,In_212);
or U248 (N_248,In_115,In_28);
or U249 (N_249,In_344,In_137);
xnor U250 (N_250,In_247,In_192);
or U251 (N_251,In_94,In_109);
nand U252 (N_252,In_110,In_328);
xnor U253 (N_253,In_282,In_449);
nor U254 (N_254,In_316,In_13);
nand U255 (N_255,In_324,In_257);
nand U256 (N_256,In_408,In_110);
nor U257 (N_257,In_182,In_116);
xor U258 (N_258,In_495,In_283);
and U259 (N_259,In_138,In_398);
nand U260 (N_260,In_192,In_388);
xor U261 (N_261,In_16,In_87);
xnor U262 (N_262,In_67,In_224);
or U263 (N_263,In_498,In_25);
xor U264 (N_264,In_404,In_71);
or U265 (N_265,In_300,In_214);
and U266 (N_266,In_120,In_50);
xnor U267 (N_267,In_412,In_320);
or U268 (N_268,In_250,In_62);
nor U269 (N_269,In_16,In_252);
and U270 (N_270,In_210,In_221);
and U271 (N_271,In_499,In_394);
and U272 (N_272,In_401,In_213);
xnor U273 (N_273,In_17,In_70);
or U274 (N_274,In_242,In_229);
nor U275 (N_275,In_222,In_381);
nand U276 (N_276,In_153,In_374);
and U277 (N_277,In_206,In_255);
and U278 (N_278,In_283,In_67);
or U279 (N_279,In_162,In_248);
or U280 (N_280,In_444,In_132);
xor U281 (N_281,In_164,In_413);
nand U282 (N_282,In_247,In_281);
xor U283 (N_283,In_174,In_198);
or U284 (N_284,In_269,In_71);
xor U285 (N_285,In_265,In_225);
nor U286 (N_286,In_163,In_347);
nor U287 (N_287,In_485,In_402);
or U288 (N_288,In_227,In_283);
xnor U289 (N_289,In_245,In_453);
xnor U290 (N_290,In_165,In_191);
nor U291 (N_291,In_349,In_199);
nor U292 (N_292,In_147,In_393);
nor U293 (N_293,In_413,In_469);
xor U294 (N_294,In_385,In_281);
or U295 (N_295,In_455,In_321);
and U296 (N_296,In_375,In_162);
nand U297 (N_297,In_142,In_214);
and U298 (N_298,In_161,In_338);
nand U299 (N_299,In_313,In_65);
xnor U300 (N_300,In_39,In_3);
nand U301 (N_301,In_120,In_32);
or U302 (N_302,In_484,In_311);
xor U303 (N_303,In_110,In_154);
nor U304 (N_304,In_445,In_160);
nand U305 (N_305,In_362,In_344);
xor U306 (N_306,In_265,In_204);
xnor U307 (N_307,In_230,In_175);
or U308 (N_308,In_299,In_341);
nand U309 (N_309,In_206,In_239);
or U310 (N_310,In_397,In_59);
or U311 (N_311,In_220,In_285);
xnor U312 (N_312,In_366,In_125);
xor U313 (N_313,In_482,In_498);
xor U314 (N_314,In_238,In_498);
and U315 (N_315,In_288,In_355);
nand U316 (N_316,In_37,In_141);
nor U317 (N_317,In_267,In_31);
xnor U318 (N_318,In_80,In_5);
nand U319 (N_319,In_186,In_90);
or U320 (N_320,In_171,In_362);
nor U321 (N_321,In_351,In_473);
and U322 (N_322,In_288,In_59);
nor U323 (N_323,In_366,In_152);
nand U324 (N_324,In_321,In_470);
and U325 (N_325,In_388,In_368);
and U326 (N_326,In_171,In_145);
nor U327 (N_327,In_109,In_289);
and U328 (N_328,In_24,In_339);
xnor U329 (N_329,In_299,In_477);
nand U330 (N_330,In_286,In_193);
nand U331 (N_331,In_490,In_143);
nor U332 (N_332,In_235,In_141);
xnor U333 (N_333,In_44,In_207);
nand U334 (N_334,In_76,In_366);
nor U335 (N_335,In_104,In_25);
or U336 (N_336,In_395,In_171);
or U337 (N_337,In_234,In_341);
and U338 (N_338,In_356,In_377);
or U339 (N_339,In_456,In_71);
or U340 (N_340,In_393,In_432);
or U341 (N_341,In_346,In_376);
or U342 (N_342,In_102,In_128);
or U343 (N_343,In_145,In_337);
xnor U344 (N_344,In_23,In_255);
nand U345 (N_345,In_439,In_476);
xor U346 (N_346,In_37,In_442);
xnor U347 (N_347,In_186,In_484);
nor U348 (N_348,In_288,In_127);
or U349 (N_349,In_202,In_122);
xor U350 (N_350,In_31,In_258);
nand U351 (N_351,In_146,In_331);
or U352 (N_352,In_303,In_428);
or U353 (N_353,In_467,In_271);
nor U354 (N_354,In_250,In_4);
and U355 (N_355,In_0,In_271);
nand U356 (N_356,In_13,In_18);
xnor U357 (N_357,In_314,In_3);
and U358 (N_358,In_119,In_475);
and U359 (N_359,In_255,In_338);
or U360 (N_360,In_301,In_242);
or U361 (N_361,In_239,In_213);
xnor U362 (N_362,In_379,In_427);
nand U363 (N_363,In_468,In_223);
and U364 (N_364,In_364,In_399);
and U365 (N_365,In_200,In_88);
xnor U366 (N_366,In_473,In_440);
nor U367 (N_367,In_370,In_354);
nor U368 (N_368,In_48,In_59);
and U369 (N_369,In_257,In_393);
or U370 (N_370,In_337,In_130);
and U371 (N_371,In_166,In_207);
or U372 (N_372,In_97,In_421);
and U373 (N_373,In_242,In_386);
nor U374 (N_374,In_83,In_468);
or U375 (N_375,In_272,In_257);
nor U376 (N_376,In_327,In_78);
xor U377 (N_377,In_138,In_192);
nand U378 (N_378,In_23,In_237);
xor U379 (N_379,In_412,In_68);
xnor U380 (N_380,In_247,In_482);
nand U381 (N_381,In_259,In_370);
xnor U382 (N_382,In_213,In_314);
nand U383 (N_383,In_42,In_375);
nand U384 (N_384,In_336,In_376);
xnor U385 (N_385,In_368,In_66);
xnor U386 (N_386,In_456,In_211);
xnor U387 (N_387,In_210,In_296);
or U388 (N_388,In_230,In_360);
nor U389 (N_389,In_280,In_290);
nand U390 (N_390,In_338,In_306);
or U391 (N_391,In_21,In_93);
nand U392 (N_392,In_57,In_414);
xnor U393 (N_393,In_268,In_323);
nor U394 (N_394,In_0,In_263);
nor U395 (N_395,In_138,In_448);
or U396 (N_396,In_195,In_29);
nor U397 (N_397,In_406,In_176);
xor U398 (N_398,In_300,In_305);
xor U399 (N_399,In_478,In_455);
nor U400 (N_400,In_377,In_133);
and U401 (N_401,In_290,In_378);
and U402 (N_402,In_254,In_371);
nor U403 (N_403,In_173,In_352);
nor U404 (N_404,In_243,In_491);
nor U405 (N_405,In_382,In_169);
or U406 (N_406,In_249,In_231);
xnor U407 (N_407,In_424,In_266);
nand U408 (N_408,In_307,In_267);
and U409 (N_409,In_218,In_8);
nand U410 (N_410,In_59,In_46);
nor U411 (N_411,In_312,In_239);
nand U412 (N_412,In_190,In_72);
xor U413 (N_413,In_141,In_186);
and U414 (N_414,In_97,In_206);
xnor U415 (N_415,In_441,In_328);
and U416 (N_416,In_310,In_24);
or U417 (N_417,In_333,In_155);
or U418 (N_418,In_42,In_276);
nand U419 (N_419,In_475,In_308);
and U420 (N_420,In_414,In_41);
or U421 (N_421,In_319,In_294);
nand U422 (N_422,In_51,In_55);
or U423 (N_423,In_81,In_393);
nand U424 (N_424,In_257,In_300);
xor U425 (N_425,In_399,In_335);
and U426 (N_426,In_155,In_106);
xnor U427 (N_427,In_371,In_253);
xnor U428 (N_428,In_410,In_164);
xor U429 (N_429,In_386,In_345);
xnor U430 (N_430,In_70,In_109);
nand U431 (N_431,In_187,In_369);
or U432 (N_432,In_203,In_207);
nor U433 (N_433,In_350,In_477);
nand U434 (N_434,In_290,In_250);
xnor U435 (N_435,In_359,In_54);
or U436 (N_436,In_179,In_43);
xnor U437 (N_437,In_14,In_494);
nand U438 (N_438,In_73,In_404);
or U439 (N_439,In_450,In_289);
xor U440 (N_440,In_249,In_122);
xor U441 (N_441,In_468,In_463);
nand U442 (N_442,In_428,In_184);
xor U443 (N_443,In_481,In_92);
nand U444 (N_444,In_182,In_489);
nand U445 (N_445,In_481,In_131);
and U446 (N_446,In_305,In_179);
and U447 (N_447,In_389,In_1);
and U448 (N_448,In_239,In_177);
nor U449 (N_449,In_306,In_74);
and U450 (N_450,In_3,In_434);
nor U451 (N_451,In_177,In_418);
nor U452 (N_452,In_221,In_226);
and U453 (N_453,In_118,In_100);
and U454 (N_454,In_297,In_296);
nand U455 (N_455,In_152,In_194);
and U456 (N_456,In_146,In_425);
nor U457 (N_457,In_407,In_86);
nor U458 (N_458,In_229,In_108);
and U459 (N_459,In_186,In_32);
nand U460 (N_460,In_13,In_230);
xor U461 (N_461,In_287,In_347);
xnor U462 (N_462,In_376,In_183);
nor U463 (N_463,In_375,In_468);
nand U464 (N_464,In_357,In_328);
and U465 (N_465,In_192,In_442);
or U466 (N_466,In_107,In_4);
nor U467 (N_467,In_340,In_11);
xnor U468 (N_468,In_384,In_275);
nor U469 (N_469,In_228,In_458);
nand U470 (N_470,In_217,In_294);
nand U471 (N_471,In_366,In_453);
xor U472 (N_472,In_71,In_20);
nor U473 (N_473,In_139,In_171);
or U474 (N_474,In_80,In_285);
nor U475 (N_475,In_63,In_80);
nor U476 (N_476,In_241,In_109);
nand U477 (N_477,In_19,In_433);
xnor U478 (N_478,In_232,In_97);
xnor U479 (N_479,In_297,In_470);
or U480 (N_480,In_363,In_93);
nand U481 (N_481,In_54,In_425);
or U482 (N_482,In_494,In_184);
xor U483 (N_483,In_357,In_167);
nand U484 (N_484,In_94,In_204);
nor U485 (N_485,In_398,In_295);
nor U486 (N_486,In_455,In_305);
xnor U487 (N_487,In_442,In_220);
and U488 (N_488,In_104,In_230);
nand U489 (N_489,In_83,In_261);
and U490 (N_490,In_259,In_3);
and U491 (N_491,In_361,In_250);
nor U492 (N_492,In_181,In_315);
xor U493 (N_493,In_32,In_247);
nor U494 (N_494,In_302,In_279);
nor U495 (N_495,In_57,In_347);
nor U496 (N_496,In_342,In_278);
nor U497 (N_497,In_6,In_373);
and U498 (N_498,In_228,In_334);
nand U499 (N_499,In_284,In_174);
or U500 (N_500,In_372,In_294);
or U501 (N_501,In_257,In_113);
nand U502 (N_502,In_475,In_268);
nand U503 (N_503,In_429,In_249);
nand U504 (N_504,In_168,In_337);
nand U505 (N_505,In_326,In_459);
or U506 (N_506,In_23,In_317);
nand U507 (N_507,In_200,In_140);
nand U508 (N_508,In_359,In_248);
or U509 (N_509,In_361,In_282);
and U510 (N_510,In_197,In_246);
and U511 (N_511,In_5,In_86);
nor U512 (N_512,In_234,In_342);
nor U513 (N_513,In_46,In_325);
nand U514 (N_514,In_305,In_435);
and U515 (N_515,In_155,In_315);
and U516 (N_516,In_315,In_451);
nor U517 (N_517,In_72,In_208);
nand U518 (N_518,In_364,In_94);
nand U519 (N_519,In_190,In_403);
and U520 (N_520,In_433,In_239);
or U521 (N_521,In_50,In_218);
or U522 (N_522,In_228,In_408);
xor U523 (N_523,In_329,In_92);
or U524 (N_524,In_211,In_122);
or U525 (N_525,In_344,In_54);
or U526 (N_526,In_128,In_39);
xnor U527 (N_527,In_44,In_393);
nor U528 (N_528,In_23,In_450);
or U529 (N_529,In_248,In_319);
xnor U530 (N_530,In_351,In_333);
nand U531 (N_531,In_438,In_302);
nand U532 (N_532,In_362,In_441);
xnor U533 (N_533,In_277,In_440);
nand U534 (N_534,In_147,In_188);
nor U535 (N_535,In_475,In_255);
and U536 (N_536,In_25,In_105);
nand U537 (N_537,In_364,In_313);
or U538 (N_538,In_312,In_370);
and U539 (N_539,In_487,In_291);
and U540 (N_540,In_202,In_35);
xor U541 (N_541,In_232,In_429);
and U542 (N_542,In_3,In_152);
xor U543 (N_543,In_169,In_130);
or U544 (N_544,In_134,In_21);
and U545 (N_545,In_463,In_428);
xnor U546 (N_546,In_392,In_291);
nor U547 (N_547,In_364,In_61);
and U548 (N_548,In_222,In_393);
and U549 (N_549,In_155,In_186);
nor U550 (N_550,In_400,In_114);
nand U551 (N_551,In_214,In_149);
or U552 (N_552,In_267,In_136);
xnor U553 (N_553,In_20,In_138);
and U554 (N_554,In_356,In_95);
nor U555 (N_555,In_364,In_13);
xor U556 (N_556,In_334,In_18);
nor U557 (N_557,In_95,In_13);
or U558 (N_558,In_381,In_345);
nand U559 (N_559,In_166,In_477);
xnor U560 (N_560,In_73,In_176);
nand U561 (N_561,In_153,In_209);
nor U562 (N_562,In_172,In_138);
xnor U563 (N_563,In_131,In_262);
nand U564 (N_564,In_55,In_259);
and U565 (N_565,In_21,In_214);
nand U566 (N_566,In_412,In_351);
nor U567 (N_567,In_330,In_468);
and U568 (N_568,In_270,In_361);
nand U569 (N_569,In_344,In_152);
or U570 (N_570,In_437,In_114);
nand U571 (N_571,In_61,In_409);
nor U572 (N_572,In_44,In_228);
nor U573 (N_573,In_275,In_303);
xor U574 (N_574,In_470,In_426);
nor U575 (N_575,In_87,In_220);
xor U576 (N_576,In_309,In_231);
or U577 (N_577,In_82,In_257);
xor U578 (N_578,In_328,In_93);
xnor U579 (N_579,In_32,In_438);
nand U580 (N_580,In_100,In_105);
xnor U581 (N_581,In_104,In_429);
and U582 (N_582,In_4,In_192);
nand U583 (N_583,In_380,In_95);
or U584 (N_584,In_454,In_347);
nor U585 (N_585,In_498,In_258);
nor U586 (N_586,In_163,In_432);
nor U587 (N_587,In_161,In_408);
and U588 (N_588,In_253,In_356);
nand U589 (N_589,In_379,In_203);
xnor U590 (N_590,In_223,In_315);
nor U591 (N_591,In_417,In_194);
or U592 (N_592,In_53,In_7);
nor U593 (N_593,In_346,In_478);
xnor U594 (N_594,In_402,In_164);
xnor U595 (N_595,In_28,In_4);
and U596 (N_596,In_285,In_89);
nand U597 (N_597,In_288,In_124);
or U598 (N_598,In_93,In_171);
and U599 (N_599,In_218,In_95);
and U600 (N_600,In_138,In_228);
nand U601 (N_601,In_79,In_472);
xnor U602 (N_602,In_109,In_153);
and U603 (N_603,In_113,In_30);
nand U604 (N_604,In_383,In_165);
and U605 (N_605,In_109,In_172);
or U606 (N_606,In_259,In_356);
and U607 (N_607,In_176,In_471);
nand U608 (N_608,In_98,In_324);
nand U609 (N_609,In_184,In_25);
and U610 (N_610,In_489,In_159);
and U611 (N_611,In_431,In_312);
nand U612 (N_612,In_328,In_490);
nand U613 (N_613,In_158,In_356);
nor U614 (N_614,In_117,In_103);
xor U615 (N_615,In_401,In_276);
xnor U616 (N_616,In_416,In_344);
and U617 (N_617,In_333,In_191);
and U618 (N_618,In_235,In_99);
nand U619 (N_619,In_123,In_214);
or U620 (N_620,In_75,In_31);
and U621 (N_621,In_335,In_18);
nand U622 (N_622,In_335,In_370);
nand U623 (N_623,In_375,In_374);
nand U624 (N_624,In_185,In_306);
nor U625 (N_625,In_375,In_169);
or U626 (N_626,In_235,In_181);
or U627 (N_627,In_164,In_206);
nand U628 (N_628,In_347,In_493);
xor U629 (N_629,In_61,In_129);
and U630 (N_630,In_20,In_15);
nand U631 (N_631,In_17,In_297);
nand U632 (N_632,In_433,In_233);
and U633 (N_633,In_356,In_495);
and U634 (N_634,In_336,In_473);
nand U635 (N_635,In_343,In_151);
nand U636 (N_636,In_275,In_456);
and U637 (N_637,In_235,In_190);
nand U638 (N_638,In_454,In_271);
nand U639 (N_639,In_374,In_344);
or U640 (N_640,In_281,In_328);
and U641 (N_641,In_398,In_290);
or U642 (N_642,In_359,In_123);
xor U643 (N_643,In_34,In_376);
or U644 (N_644,In_140,In_129);
or U645 (N_645,In_417,In_347);
nand U646 (N_646,In_206,In_321);
and U647 (N_647,In_324,In_153);
xor U648 (N_648,In_37,In_237);
and U649 (N_649,In_410,In_278);
xor U650 (N_650,In_220,In_13);
xor U651 (N_651,In_113,In_249);
nor U652 (N_652,In_356,In_339);
and U653 (N_653,In_283,In_155);
nor U654 (N_654,In_363,In_407);
xor U655 (N_655,In_278,In_30);
xor U656 (N_656,In_363,In_354);
and U657 (N_657,In_140,In_378);
and U658 (N_658,In_196,In_183);
and U659 (N_659,In_66,In_374);
xor U660 (N_660,In_113,In_340);
xnor U661 (N_661,In_286,In_263);
nor U662 (N_662,In_367,In_348);
and U663 (N_663,In_126,In_70);
nand U664 (N_664,In_222,In_338);
xnor U665 (N_665,In_163,In_433);
and U666 (N_666,In_297,In_220);
and U667 (N_667,In_260,In_306);
and U668 (N_668,In_329,In_220);
nor U669 (N_669,In_447,In_124);
xor U670 (N_670,In_16,In_437);
or U671 (N_671,In_433,In_360);
xor U672 (N_672,In_6,In_287);
xnor U673 (N_673,In_237,In_97);
and U674 (N_674,In_137,In_330);
xor U675 (N_675,In_7,In_337);
nor U676 (N_676,In_484,In_496);
and U677 (N_677,In_403,In_353);
xor U678 (N_678,In_5,In_462);
nor U679 (N_679,In_12,In_497);
nand U680 (N_680,In_119,In_237);
or U681 (N_681,In_167,In_313);
or U682 (N_682,In_178,In_437);
and U683 (N_683,In_284,In_83);
or U684 (N_684,In_242,In_69);
or U685 (N_685,In_327,In_392);
nor U686 (N_686,In_354,In_308);
nor U687 (N_687,In_45,In_240);
or U688 (N_688,In_476,In_123);
nand U689 (N_689,In_219,In_98);
nor U690 (N_690,In_140,In_29);
xnor U691 (N_691,In_91,In_95);
nor U692 (N_692,In_449,In_350);
nand U693 (N_693,In_112,In_488);
nand U694 (N_694,In_79,In_189);
nor U695 (N_695,In_180,In_267);
nor U696 (N_696,In_55,In_240);
or U697 (N_697,In_417,In_76);
xnor U698 (N_698,In_268,In_206);
and U699 (N_699,In_89,In_373);
nor U700 (N_700,In_157,In_216);
nand U701 (N_701,In_145,In_16);
xnor U702 (N_702,In_125,In_65);
and U703 (N_703,In_206,In_223);
xor U704 (N_704,In_59,In_94);
nand U705 (N_705,In_345,In_371);
and U706 (N_706,In_5,In_93);
xor U707 (N_707,In_69,In_487);
or U708 (N_708,In_290,In_17);
xor U709 (N_709,In_146,In_354);
and U710 (N_710,In_465,In_416);
nor U711 (N_711,In_269,In_235);
xor U712 (N_712,In_304,In_116);
or U713 (N_713,In_10,In_254);
xor U714 (N_714,In_116,In_270);
and U715 (N_715,In_291,In_428);
or U716 (N_716,In_339,In_195);
or U717 (N_717,In_141,In_171);
and U718 (N_718,In_499,In_10);
nand U719 (N_719,In_410,In_323);
nor U720 (N_720,In_232,In_268);
xor U721 (N_721,In_416,In_458);
xor U722 (N_722,In_79,In_70);
and U723 (N_723,In_275,In_431);
nor U724 (N_724,In_413,In_431);
xor U725 (N_725,In_495,In_423);
and U726 (N_726,In_409,In_249);
xnor U727 (N_727,In_219,In_13);
nand U728 (N_728,In_164,In_286);
nor U729 (N_729,In_364,In_85);
nor U730 (N_730,In_178,In_252);
and U731 (N_731,In_325,In_264);
and U732 (N_732,In_115,In_130);
or U733 (N_733,In_14,In_269);
nor U734 (N_734,In_333,In_158);
xor U735 (N_735,In_70,In_232);
nand U736 (N_736,In_167,In_434);
or U737 (N_737,In_89,In_15);
nand U738 (N_738,In_470,In_73);
xor U739 (N_739,In_264,In_45);
xor U740 (N_740,In_193,In_47);
and U741 (N_741,In_18,In_208);
nand U742 (N_742,In_25,In_367);
nor U743 (N_743,In_475,In_174);
or U744 (N_744,In_135,In_218);
or U745 (N_745,In_234,In_71);
xnor U746 (N_746,In_5,In_197);
nor U747 (N_747,In_361,In_232);
xnor U748 (N_748,In_17,In_391);
nor U749 (N_749,In_206,In_229);
nor U750 (N_750,N_222,N_720);
nor U751 (N_751,N_267,N_130);
xor U752 (N_752,N_213,N_573);
xnor U753 (N_753,N_671,N_735);
xor U754 (N_754,N_27,N_476);
xor U755 (N_755,N_269,N_627);
or U756 (N_756,N_379,N_400);
nand U757 (N_757,N_40,N_74);
or U758 (N_758,N_164,N_180);
and U759 (N_759,N_740,N_746);
nand U760 (N_760,N_188,N_570);
xor U761 (N_761,N_734,N_230);
or U762 (N_762,N_274,N_246);
nor U763 (N_763,N_549,N_647);
and U764 (N_764,N_457,N_625);
nand U765 (N_765,N_727,N_435);
and U766 (N_766,N_628,N_724);
xnor U767 (N_767,N_508,N_108);
and U768 (N_768,N_626,N_373);
nand U769 (N_769,N_516,N_713);
nand U770 (N_770,N_646,N_490);
and U771 (N_771,N_449,N_429);
nand U772 (N_772,N_126,N_521);
xnor U773 (N_773,N_183,N_389);
nand U774 (N_774,N_434,N_640);
and U775 (N_775,N_420,N_357);
nand U776 (N_776,N_600,N_633);
xor U777 (N_777,N_321,N_387);
and U778 (N_778,N_263,N_468);
or U779 (N_779,N_107,N_422);
nor U780 (N_780,N_191,N_169);
xnor U781 (N_781,N_660,N_150);
or U782 (N_782,N_90,N_425);
nand U783 (N_783,N_316,N_220);
or U784 (N_784,N_391,N_704);
nor U785 (N_785,N_441,N_326);
nor U786 (N_786,N_271,N_374);
or U787 (N_787,N_731,N_201);
or U788 (N_788,N_437,N_63);
nor U789 (N_789,N_284,N_385);
nor U790 (N_790,N_162,N_466);
nand U791 (N_791,N_665,N_125);
xor U792 (N_792,N_629,N_716);
or U793 (N_793,N_670,N_75);
and U794 (N_794,N_370,N_632);
and U795 (N_795,N_683,N_433);
nand U796 (N_796,N_312,N_555);
and U797 (N_797,N_708,N_14);
or U798 (N_798,N_428,N_289);
or U799 (N_799,N_645,N_705);
xor U800 (N_800,N_648,N_149);
or U801 (N_801,N_743,N_382);
nand U802 (N_802,N_539,N_639);
nor U803 (N_803,N_66,N_657);
and U804 (N_804,N_736,N_693);
xor U805 (N_805,N_447,N_403);
and U806 (N_806,N_28,N_182);
nand U807 (N_807,N_21,N_679);
nor U808 (N_808,N_455,N_86);
nor U809 (N_809,N_733,N_376);
xnor U810 (N_810,N_452,N_300);
or U811 (N_811,N_189,N_674);
nor U812 (N_812,N_275,N_745);
or U813 (N_813,N_407,N_232);
and U814 (N_814,N_446,N_318);
and U815 (N_815,N_116,N_694);
and U816 (N_816,N_340,N_637);
or U817 (N_817,N_5,N_0);
xor U818 (N_818,N_60,N_586);
or U819 (N_819,N_609,N_245);
or U820 (N_820,N_748,N_358);
or U821 (N_821,N_73,N_545);
xor U822 (N_822,N_236,N_620);
xnor U823 (N_823,N_22,N_459);
nor U824 (N_824,N_239,N_285);
or U825 (N_825,N_596,N_479);
or U826 (N_826,N_268,N_592);
nand U827 (N_827,N_322,N_95);
or U828 (N_828,N_112,N_439);
nand U829 (N_829,N_484,N_525);
or U830 (N_830,N_590,N_481);
nor U831 (N_831,N_579,N_546);
or U832 (N_832,N_352,N_383);
xnor U833 (N_833,N_1,N_44);
or U834 (N_834,N_401,N_91);
xnor U835 (N_835,N_210,N_578);
or U836 (N_836,N_386,N_438);
nor U837 (N_837,N_390,N_166);
and U838 (N_838,N_522,N_652);
xnor U839 (N_839,N_356,N_121);
xnor U840 (N_840,N_360,N_281);
or U841 (N_841,N_412,N_717);
and U842 (N_842,N_601,N_491);
or U843 (N_843,N_461,N_682);
nor U844 (N_844,N_39,N_749);
nand U845 (N_845,N_675,N_470);
or U846 (N_846,N_698,N_124);
and U847 (N_847,N_410,N_686);
and U848 (N_848,N_738,N_494);
nand U849 (N_849,N_336,N_97);
or U850 (N_850,N_132,N_584);
xor U851 (N_851,N_314,N_529);
nor U852 (N_852,N_242,N_260);
and U853 (N_853,N_313,N_524);
nor U854 (N_854,N_141,N_54);
xor U855 (N_855,N_688,N_31);
or U856 (N_856,N_547,N_576);
xnor U857 (N_857,N_496,N_170);
and U858 (N_858,N_581,N_719);
or U859 (N_859,N_582,N_131);
and U860 (N_860,N_254,N_26);
or U861 (N_861,N_598,N_709);
nor U862 (N_862,N_78,N_741);
nand U863 (N_863,N_544,N_493);
xor U864 (N_864,N_324,N_474);
xnor U865 (N_865,N_402,N_71);
xnor U866 (N_866,N_585,N_695);
xor U867 (N_867,N_37,N_380);
and U868 (N_868,N_610,N_46);
xnor U869 (N_869,N_540,N_597);
xor U870 (N_870,N_365,N_145);
and U871 (N_871,N_50,N_42);
and U872 (N_872,N_594,N_472);
xnor U873 (N_873,N_565,N_175);
or U874 (N_874,N_621,N_566);
xnor U875 (N_875,N_553,N_375);
nand U876 (N_876,N_122,N_485);
xnor U877 (N_877,N_513,N_61);
xnor U878 (N_878,N_424,N_681);
and U879 (N_879,N_371,N_292);
and U880 (N_880,N_413,N_241);
xor U881 (N_881,N_554,N_193);
nor U882 (N_882,N_649,N_173);
xnor U883 (N_883,N_426,N_15);
and U884 (N_884,N_2,N_52);
nor U885 (N_885,N_510,N_266);
nor U886 (N_886,N_622,N_378);
nor U887 (N_887,N_687,N_286);
or U888 (N_888,N_408,N_115);
or U889 (N_889,N_317,N_663);
xnor U890 (N_890,N_226,N_742);
nor U891 (N_891,N_451,N_673);
nor U892 (N_892,N_415,N_293);
nand U893 (N_893,N_345,N_443);
or U894 (N_894,N_248,N_616);
and U895 (N_895,N_467,N_41);
or U896 (N_896,N_344,N_589);
nand U897 (N_897,N_482,N_168);
nand U898 (N_898,N_250,N_432);
nor U899 (N_899,N_18,N_299);
and U900 (N_900,N_45,N_49);
and U901 (N_901,N_158,N_302);
or U902 (N_902,N_187,N_475);
and U903 (N_903,N_635,N_612);
nand U904 (N_904,N_348,N_153);
or U905 (N_905,N_197,N_89);
nor U906 (N_906,N_367,N_53);
xnor U907 (N_907,N_165,N_702);
nand U908 (N_908,N_445,N_676);
nor U909 (N_909,N_231,N_473);
nand U910 (N_910,N_76,N_247);
and U911 (N_911,N_557,N_331);
xor U912 (N_912,N_611,N_176);
xor U913 (N_913,N_337,N_329);
nor U914 (N_914,N_478,N_243);
or U915 (N_915,N_689,N_83);
nand U916 (N_916,N_159,N_283);
nand U917 (N_917,N_70,N_151);
nor U918 (N_918,N_414,N_580);
or U919 (N_919,N_67,N_192);
or U920 (N_920,N_335,N_364);
or U921 (N_921,N_349,N_330);
and U922 (N_922,N_261,N_362);
nor U923 (N_923,N_699,N_664);
nand U924 (N_924,N_543,N_462);
xor U925 (N_925,N_138,N_65);
and U926 (N_926,N_186,N_377);
nor U927 (N_927,N_181,N_661);
and U928 (N_928,N_258,N_531);
nand U929 (N_929,N_99,N_471);
nand U930 (N_930,N_23,N_120);
nor U931 (N_931,N_214,N_558);
nand U932 (N_932,N_282,N_103);
xnor U933 (N_933,N_7,N_556);
or U934 (N_934,N_307,N_87);
xor U935 (N_935,N_77,N_477);
and U936 (N_936,N_217,N_142);
and U937 (N_937,N_667,N_505);
and U938 (N_938,N_572,N_134);
and U939 (N_939,N_397,N_119);
nor U940 (N_940,N_235,N_604);
and U941 (N_941,N_228,N_690);
nand U942 (N_942,N_684,N_599);
nand U943 (N_943,N_118,N_262);
nand U944 (N_944,N_721,N_533);
or U945 (N_945,N_587,N_700);
and U946 (N_946,N_36,N_714);
and U947 (N_947,N_630,N_677);
nor U948 (N_948,N_642,N_225);
xor U949 (N_949,N_11,N_515);
nor U950 (N_950,N_227,N_588);
nand U951 (N_951,N_233,N_517);
and U952 (N_952,N_562,N_221);
xnor U953 (N_953,N_301,N_644);
nand U954 (N_954,N_519,N_306);
nand U955 (N_955,N_305,N_106);
nor U956 (N_956,N_59,N_272);
xor U957 (N_957,N_623,N_614);
nand U958 (N_958,N_526,N_489);
xor U959 (N_959,N_707,N_501);
nor U960 (N_960,N_259,N_550);
nor U961 (N_961,N_495,N_33);
nand U962 (N_962,N_35,N_315);
or U963 (N_963,N_499,N_659);
nor U964 (N_964,N_295,N_507);
nand U965 (N_965,N_398,N_416);
nor U966 (N_966,N_480,N_334);
and U967 (N_967,N_64,N_123);
or U968 (N_968,N_653,N_57);
and U969 (N_969,N_678,N_725);
nor U970 (N_970,N_19,N_185);
xor U971 (N_971,N_528,N_464);
and U972 (N_972,N_602,N_190);
nand U973 (N_973,N_229,N_163);
or U974 (N_974,N_409,N_363);
nand U975 (N_975,N_339,N_105);
nor U976 (N_976,N_114,N_101);
nor U977 (N_977,N_148,N_288);
xnor U978 (N_978,N_34,N_366);
or U979 (N_979,N_171,N_656);
or U980 (N_980,N_442,N_174);
nor U981 (N_981,N_133,N_668);
xnor U982 (N_982,N_146,N_732);
nand U983 (N_983,N_606,N_591);
nand U984 (N_984,N_706,N_483);
or U985 (N_985,N_448,N_654);
nand U986 (N_986,N_223,N_583);
nor U987 (N_987,N_79,N_351);
xnor U988 (N_988,N_160,N_179);
and U989 (N_989,N_184,N_4);
xor U990 (N_990,N_692,N_207);
xnor U991 (N_991,N_739,N_712);
xor U992 (N_992,N_718,N_701);
nor U993 (N_993,N_215,N_372);
nor U994 (N_994,N_427,N_279);
and U995 (N_995,N_251,N_58);
and U996 (N_996,N_498,N_615);
or U997 (N_997,N_518,N_541);
and U998 (N_998,N_619,N_111);
and U999 (N_999,N_651,N_234);
nor U1000 (N_1000,N_384,N_744);
nand U1001 (N_1001,N_634,N_393);
and U1002 (N_1002,N_30,N_287);
xnor U1003 (N_1003,N_156,N_25);
nand U1004 (N_1004,N_641,N_728);
and U1005 (N_1005,N_135,N_104);
nand U1006 (N_1006,N_723,N_394);
or U1007 (N_1007,N_430,N_294);
and U1008 (N_1008,N_548,N_444);
or U1009 (N_1009,N_298,N_147);
nand U1010 (N_1010,N_617,N_527);
and U1011 (N_1011,N_24,N_280);
or U1012 (N_1012,N_198,N_535);
xnor U1013 (N_1013,N_310,N_152);
and U1014 (N_1014,N_80,N_249);
nand U1015 (N_1015,N_55,N_325);
and U1016 (N_1016,N_206,N_199);
or U1017 (N_1017,N_423,N_488);
and U1018 (N_1018,N_208,N_341);
and U1019 (N_1019,N_569,N_405);
nand U1020 (N_1020,N_143,N_304);
nor U1021 (N_1021,N_320,N_436);
or U1022 (N_1022,N_368,N_418);
nand U1023 (N_1023,N_219,N_154);
and U1024 (N_1024,N_560,N_512);
and U1025 (N_1025,N_511,N_563);
or U1026 (N_1026,N_13,N_722);
xnor U1027 (N_1027,N_38,N_711);
nor U1028 (N_1028,N_82,N_85);
nor U1029 (N_1029,N_458,N_297);
and U1030 (N_1030,N_296,N_195);
nand U1031 (N_1031,N_456,N_685);
nand U1032 (N_1032,N_68,N_534);
or U1033 (N_1033,N_669,N_244);
nor U1034 (N_1034,N_202,N_369);
xnor U1035 (N_1035,N_463,N_20);
and U1036 (N_1036,N_178,N_561);
nand U1037 (N_1037,N_672,N_605);
nor U1038 (N_1038,N_167,N_290);
nor U1039 (N_1039,N_200,N_577);
nand U1040 (N_1040,N_574,N_551);
nor U1041 (N_1041,N_381,N_638);
and U1042 (N_1042,N_662,N_559);
or U1043 (N_1043,N_608,N_666);
or U1044 (N_1044,N_431,N_278);
or U1045 (N_1045,N_353,N_388);
xnor U1046 (N_1046,N_238,N_308);
or U1047 (N_1047,N_16,N_117);
nand U1048 (N_1048,N_504,N_161);
nand U1049 (N_1049,N_177,N_155);
and U1050 (N_1050,N_273,N_658);
and U1051 (N_1051,N_710,N_697);
xor U1052 (N_1052,N_136,N_139);
or U1053 (N_1053,N_726,N_696);
xnor U1054 (N_1054,N_252,N_417);
or U1055 (N_1055,N_8,N_575);
nand U1056 (N_1056,N_264,N_691);
nor U1057 (N_1057,N_538,N_32);
or U1058 (N_1058,N_276,N_514);
and U1059 (N_1059,N_311,N_440);
xnor U1060 (N_1060,N_81,N_359);
or U1061 (N_1061,N_327,N_595);
xor U1062 (N_1062,N_17,N_350);
xor U1063 (N_1063,N_343,N_624);
or U1064 (N_1064,N_487,N_94);
xor U1065 (N_1065,N_98,N_137);
nor U1066 (N_1066,N_460,N_421);
nor U1067 (N_1067,N_607,N_29);
and U1068 (N_1068,N_6,N_631);
nor U1069 (N_1069,N_399,N_224);
xnor U1070 (N_1070,N_93,N_354);
or U1071 (N_1071,N_205,N_500);
nor U1072 (N_1072,N_568,N_395);
or U1073 (N_1073,N_536,N_9);
xor U1074 (N_1074,N_12,N_747);
xor U1075 (N_1075,N_564,N_237);
nor U1076 (N_1076,N_532,N_503);
nor U1077 (N_1077,N_506,N_453);
and U1078 (N_1078,N_255,N_392);
nor U1079 (N_1079,N_129,N_567);
or U1080 (N_1080,N_328,N_265);
nand U1081 (N_1081,N_465,N_454);
nand U1082 (N_1082,N_730,N_257);
or U1083 (N_1083,N_277,N_613);
xor U1084 (N_1084,N_338,N_530);
nor U1085 (N_1085,N_486,N_212);
or U1086 (N_1086,N_10,N_361);
or U1087 (N_1087,N_319,N_643);
and U1088 (N_1088,N_253,N_419);
and U1089 (N_1089,N_323,N_650);
nor U1090 (N_1090,N_469,N_303);
nand U1091 (N_1091,N_537,N_404);
nand U1092 (N_1092,N_332,N_396);
nor U1093 (N_1093,N_92,N_571);
and U1094 (N_1094,N_204,N_128);
xnor U1095 (N_1095,N_203,N_100);
nor U1096 (N_1096,N_144,N_256);
or U1097 (N_1097,N_109,N_96);
nand U1098 (N_1098,N_655,N_406);
or U1099 (N_1099,N_291,N_211);
nand U1100 (N_1100,N_240,N_110);
nand U1101 (N_1101,N_69,N_603);
xnor U1102 (N_1102,N_209,N_333);
nand U1103 (N_1103,N_270,N_157);
or U1104 (N_1104,N_715,N_342);
or U1105 (N_1105,N_520,N_127);
nand U1106 (N_1106,N_680,N_51);
and U1107 (N_1107,N_196,N_48);
xnor U1108 (N_1108,N_346,N_703);
xnor U1109 (N_1109,N_3,N_737);
or U1110 (N_1110,N_218,N_216);
nor U1111 (N_1111,N_194,N_411);
nand U1112 (N_1112,N_552,N_618);
nor U1113 (N_1113,N_43,N_172);
nor U1114 (N_1114,N_47,N_84);
xor U1115 (N_1115,N_502,N_72);
or U1116 (N_1116,N_309,N_593);
or U1117 (N_1117,N_542,N_102);
and U1118 (N_1118,N_523,N_62);
nand U1119 (N_1119,N_140,N_450);
or U1120 (N_1120,N_347,N_509);
and U1121 (N_1121,N_56,N_88);
nand U1122 (N_1122,N_497,N_729);
xor U1123 (N_1123,N_492,N_636);
and U1124 (N_1124,N_355,N_113);
or U1125 (N_1125,N_460,N_386);
xor U1126 (N_1126,N_506,N_57);
or U1127 (N_1127,N_105,N_325);
nor U1128 (N_1128,N_267,N_395);
xnor U1129 (N_1129,N_217,N_186);
xor U1130 (N_1130,N_243,N_624);
and U1131 (N_1131,N_165,N_399);
xnor U1132 (N_1132,N_230,N_386);
xnor U1133 (N_1133,N_276,N_308);
and U1134 (N_1134,N_194,N_353);
xnor U1135 (N_1135,N_109,N_409);
nand U1136 (N_1136,N_704,N_208);
nor U1137 (N_1137,N_399,N_27);
nand U1138 (N_1138,N_459,N_658);
xnor U1139 (N_1139,N_192,N_201);
and U1140 (N_1140,N_411,N_223);
xnor U1141 (N_1141,N_220,N_85);
xnor U1142 (N_1142,N_27,N_236);
xnor U1143 (N_1143,N_693,N_200);
nand U1144 (N_1144,N_514,N_280);
or U1145 (N_1145,N_536,N_231);
xnor U1146 (N_1146,N_361,N_347);
xor U1147 (N_1147,N_435,N_177);
and U1148 (N_1148,N_288,N_346);
xor U1149 (N_1149,N_48,N_283);
or U1150 (N_1150,N_128,N_194);
or U1151 (N_1151,N_445,N_19);
nor U1152 (N_1152,N_373,N_743);
xor U1153 (N_1153,N_612,N_142);
or U1154 (N_1154,N_622,N_483);
nor U1155 (N_1155,N_126,N_613);
nand U1156 (N_1156,N_243,N_202);
nor U1157 (N_1157,N_361,N_704);
xor U1158 (N_1158,N_148,N_507);
nor U1159 (N_1159,N_573,N_129);
nor U1160 (N_1160,N_494,N_105);
nor U1161 (N_1161,N_309,N_412);
nor U1162 (N_1162,N_697,N_73);
xor U1163 (N_1163,N_443,N_734);
nor U1164 (N_1164,N_715,N_204);
or U1165 (N_1165,N_593,N_209);
nor U1166 (N_1166,N_118,N_173);
and U1167 (N_1167,N_605,N_283);
and U1168 (N_1168,N_386,N_737);
nand U1169 (N_1169,N_53,N_191);
and U1170 (N_1170,N_150,N_419);
nand U1171 (N_1171,N_516,N_204);
and U1172 (N_1172,N_690,N_343);
or U1173 (N_1173,N_354,N_10);
nand U1174 (N_1174,N_69,N_257);
or U1175 (N_1175,N_518,N_381);
nand U1176 (N_1176,N_6,N_21);
and U1177 (N_1177,N_267,N_122);
xor U1178 (N_1178,N_299,N_405);
xor U1179 (N_1179,N_546,N_430);
nor U1180 (N_1180,N_619,N_391);
and U1181 (N_1181,N_8,N_337);
nor U1182 (N_1182,N_304,N_22);
and U1183 (N_1183,N_460,N_596);
and U1184 (N_1184,N_57,N_130);
or U1185 (N_1185,N_698,N_672);
nor U1186 (N_1186,N_744,N_380);
nor U1187 (N_1187,N_138,N_439);
or U1188 (N_1188,N_39,N_297);
nor U1189 (N_1189,N_312,N_603);
xor U1190 (N_1190,N_206,N_673);
nand U1191 (N_1191,N_648,N_675);
nor U1192 (N_1192,N_372,N_444);
and U1193 (N_1193,N_640,N_310);
and U1194 (N_1194,N_273,N_108);
nand U1195 (N_1195,N_515,N_162);
or U1196 (N_1196,N_645,N_293);
or U1197 (N_1197,N_639,N_522);
nor U1198 (N_1198,N_430,N_41);
or U1199 (N_1199,N_351,N_269);
nand U1200 (N_1200,N_513,N_707);
nor U1201 (N_1201,N_56,N_114);
and U1202 (N_1202,N_8,N_728);
nor U1203 (N_1203,N_324,N_423);
nand U1204 (N_1204,N_707,N_540);
and U1205 (N_1205,N_206,N_124);
and U1206 (N_1206,N_156,N_620);
and U1207 (N_1207,N_390,N_283);
nor U1208 (N_1208,N_603,N_21);
xor U1209 (N_1209,N_231,N_70);
nand U1210 (N_1210,N_23,N_72);
nor U1211 (N_1211,N_554,N_271);
and U1212 (N_1212,N_323,N_172);
nor U1213 (N_1213,N_55,N_50);
xnor U1214 (N_1214,N_32,N_308);
nor U1215 (N_1215,N_653,N_384);
or U1216 (N_1216,N_593,N_524);
nor U1217 (N_1217,N_399,N_226);
or U1218 (N_1218,N_80,N_559);
nand U1219 (N_1219,N_549,N_411);
nand U1220 (N_1220,N_53,N_139);
and U1221 (N_1221,N_230,N_469);
or U1222 (N_1222,N_72,N_321);
or U1223 (N_1223,N_629,N_176);
nor U1224 (N_1224,N_455,N_265);
and U1225 (N_1225,N_110,N_127);
xnor U1226 (N_1226,N_487,N_525);
or U1227 (N_1227,N_264,N_229);
nor U1228 (N_1228,N_324,N_410);
nor U1229 (N_1229,N_23,N_495);
and U1230 (N_1230,N_658,N_122);
nand U1231 (N_1231,N_472,N_239);
xor U1232 (N_1232,N_306,N_241);
xnor U1233 (N_1233,N_561,N_281);
or U1234 (N_1234,N_708,N_138);
and U1235 (N_1235,N_529,N_624);
xnor U1236 (N_1236,N_720,N_130);
nor U1237 (N_1237,N_656,N_2);
xor U1238 (N_1238,N_574,N_282);
nor U1239 (N_1239,N_544,N_540);
or U1240 (N_1240,N_19,N_618);
nand U1241 (N_1241,N_457,N_295);
xor U1242 (N_1242,N_743,N_409);
nor U1243 (N_1243,N_283,N_588);
and U1244 (N_1244,N_352,N_728);
and U1245 (N_1245,N_268,N_610);
nand U1246 (N_1246,N_258,N_556);
xnor U1247 (N_1247,N_347,N_128);
and U1248 (N_1248,N_342,N_714);
xnor U1249 (N_1249,N_422,N_129);
and U1250 (N_1250,N_725,N_28);
nand U1251 (N_1251,N_582,N_684);
and U1252 (N_1252,N_477,N_15);
xor U1253 (N_1253,N_347,N_13);
and U1254 (N_1254,N_336,N_302);
and U1255 (N_1255,N_300,N_744);
nand U1256 (N_1256,N_180,N_192);
nand U1257 (N_1257,N_258,N_364);
nor U1258 (N_1258,N_119,N_587);
and U1259 (N_1259,N_282,N_727);
and U1260 (N_1260,N_427,N_362);
nand U1261 (N_1261,N_218,N_572);
xnor U1262 (N_1262,N_556,N_618);
nor U1263 (N_1263,N_67,N_22);
and U1264 (N_1264,N_213,N_640);
or U1265 (N_1265,N_45,N_706);
nand U1266 (N_1266,N_106,N_297);
and U1267 (N_1267,N_534,N_78);
nand U1268 (N_1268,N_649,N_729);
xnor U1269 (N_1269,N_82,N_188);
or U1270 (N_1270,N_741,N_604);
nor U1271 (N_1271,N_415,N_569);
nand U1272 (N_1272,N_294,N_531);
and U1273 (N_1273,N_106,N_454);
nor U1274 (N_1274,N_538,N_338);
nor U1275 (N_1275,N_501,N_89);
nand U1276 (N_1276,N_368,N_532);
xor U1277 (N_1277,N_483,N_678);
xor U1278 (N_1278,N_694,N_422);
nand U1279 (N_1279,N_279,N_104);
nand U1280 (N_1280,N_295,N_709);
nand U1281 (N_1281,N_407,N_277);
nor U1282 (N_1282,N_133,N_172);
xor U1283 (N_1283,N_383,N_686);
or U1284 (N_1284,N_114,N_660);
or U1285 (N_1285,N_271,N_645);
nor U1286 (N_1286,N_599,N_483);
xor U1287 (N_1287,N_438,N_446);
nand U1288 (N_1288,N_36,N_511);
nand U1289 (N_1289,N_565,N_642);
nand U1290 (N_1290,N_281,N_647);
nand U1291 (N_1291,N_533,N_619);
nor U1292 (N_1292,N_402,N_125);
nor U1293 (N_1293,N_696,N_387);
nand U1294 (N_1294,N_738,N_503);
xnor U1295 (N_1295,N_716,N_112);
nand U1296 (N_1296,N_219,N_534);
or U1297 (N_1297,N_219,N_339);
xor U1298 (N_1298,N_266,N_522);
and U1299 (N_1299,N_394,N_162);
or U1300 (N_1300,N_409,N_546);
nor U1301 (N_1301,N_312,N_133);
xnor U1302 (N_1302,N_26,N_102);
or U1303 (N_1303,N_375,N_196);
nand U1304 (N_1304,N_162,N_266);
and U1305 (N_1305,N_702,N_82);
or U1306 (N_1306,N_572,N_151);
or U1307 (N_1307,N_409,N_671);
xnor U1308 (N_1308,N_671,N_504);
xnor U1309 (N_1309,N_216,N_40);
xor U1310 (N_1310,N_685,N_344);
xnor U1311 (N_1311,N_18,N_618);
xor U1312 (N_1312,N_746,N_482);
nand U1313 (N_1313,N_24,N_447);
and U1314 (N_1314,N_435,N_312);
nor U1315 (N_1315,N_318,N_569);
nand U1316 (N_1316,N_40,N_328);
or U1317 (N_1317,N_292,N_665);
nand U1318 (N_1318,N_712,N_226);
nor U1319 (N_1319,N_89,N_690);
and U1320 (N_1320,N_699,N_109);
nand U1321 (N_1321,N_109,N_126);
nand U1322 (N_1322,N_722,N_473);
and U1323 (N_1323,N_17,N_319);
xor U1324 (N_1324,N_283,N_259);
nor U1325 (N_1325,N_324,N_307);
nor U1326 (N_1326,N_338,N_43);
nor U1327 (N_1327,N_477,N_382);
nand U1328 (N_1328,N_524,N_239);
and U1329 (N_1329,N_265,N_110);
nor U1330 (N_1330,N_310,N_42);
or U1331 (N_1331,N_111,N_538);
nor U1332 (N_1332,N_471,N_603);
and U1333 (N_1333,N_369,N_231);
xor U1334 (N_1334,N_532,N_561);
or U1335 (N_1335,N_274,N_723);
nor U1336 (N_1336,N_258,N_442);
nand U1337 (N_1337,N_358,N_377);
nand U1338 (N_1338,N_306,N_353);
and U1339 (N_1339,N_441,N_522);
and U1340 (N_1340,N_286,N_323);
xnor U1341 (N_1341,N_522,N_496);
nand U1342 (N_1342,N_230,N_105);
nand U1343 (N_1343,N_415,N_24);
nor U1344 (N_1344,N_108,N_32);
xor U1345 (N_1345,N_202,N_566);
nor U1346 (N_1346,N_745,N_471);
nand U1347 (N_1347,N_674,N_511);
xor U1348 (N_1348,N_749,N_184);
or U1349 (N_1349,N_623,N_428);
xnor U1350 (N_1350,N_713,N_127);
and U1351 (N_1351,N_471,N_248);
xor U1352 (N_1352,N_48,N_550);
xor U1353 (N_1353,N_580,N_488);
nand U1354 (N_1354,N_164,N_525);
xor U1355 (N_1355,N_732,N_22);
or U1356 (N_1356,N_0,N_488);
or U1357 (N_1357,N_446,N_248);
and U1358 (N_1358,N_223,N_494);
nand U1359 (N_1359,N_33,N_103);
or U1360 (N_1360,N_238,N_623);
xnor U1361 (N_1361,N_263,N_154);
xor U1362 (N_1362,N_302,N_90);
nor U1363 (N_1363,N_8,N_514);
or U1364 (N_1364,N_441,N_393);
xnor U1365 (N_1365,N_42,N_316);
or U1366 (N_1366,N_180,N_505);
nor U1367 (N_1367,N_591,N_301);
nand U1368 (N_1368,N_441,N_114);
nand U1369 (N_1369,N_90,N_489);
or U1370 (N_1370,N_132,N_647);
nand U1371 (N_1371,N_392,N_389);
xor U1372 (N_1372,N_8,N_331);
xnor U1373 (N_1373,N_375,N_50);
xor U1374 (N_1374,N_478,N_8);
nor U1375 (N_1375,N_227,N_434);
and U1376 (N_1376,N_119,N_369);
nor U1377 (N_1377,N_677,N_222);
nand U1378 (N_1378,N_355,N_46);
and U1379 (N_1379,N_516,N_22);
nor U1380 (N_1380,N_683,N_18);
nand U1381 (N_1381,N_170,N_80);
or U1382 (N_1382,N_270,N_233);
and U1383 (N_1383,N_330,N_182);
nor U1384 (N_1384,N_478,N_442);
and U1385 (N_1385,N_446,N_460);
or U1386 (N_1386,N_132,N_481);
nand U1387 (N_1387,N_684,N_301);
xnor U1388 (N_1388,N_106,N_134);
xnor U1389 (N_1389,N_584,N_423);
nor U1390 (N_1390,N_679,N_225);
and U1391 (N_1391,N_96,N_477);
or U1392 (N_1392,N_65,N_85);
and U1393 (N_1393,N_428,N_705);
and U1394 (N_1394,N_674,N_609);
nor U1395 (N_1395,N_50,N_421);
or U1396 (N_1396,N_511,N_147);
nand U1397 (N_1397,N_669,N_663);
nor U1398 (N_1398,N_482,N_476);
xnor U1399 (N_1399,N_678,N_420);
xnor U1400 (N_1400,N_179,N_571);
xnor U1401 (N_1401,N_450,N_651);
or U1402 (N_1402,N_737,N_151);
or U1403 (N_1403,N_721,N_15);
nand U1404 (N_1404,N_690,N_44);
or U1405 (N_1405,N_417,N_641);
nand U1406 (N_1406,N_450,N_736);
nor U1407 (N_1407,N_612,N_140);
or U1408 (N_1408,N_614,N_435);
nand U1409 (N_1409,N_221,N_214);
nor U1410 (N_1410,N_749,N_260);
or U1411 (N_1411,N_174,N_246);
xnor U1412 (N_1412,N_156,N_272);
xnor U1413 (N_1413,N_137,N_749);
nor U1414 (N_1414,N_458,N_426);
and U1415 (N_1415,N_190,N_437);
nand U1416 (N_1416,N_732,N_304);
or U1417 (N_1417,N_627,N_324);
xnor U1418 (N_1418,N_499,N_576);
xor U1419 (N_1419,N_577,N_541);
xor U1420 (N_1420,N_673,N_411);
and U1421 (N_1421,N_540,N_618);
xnor U1422 (N_1422,N_449,N_61);
xor U1423 (N_1423,N_140,N_692);
nand U1424 (N_1424,N_348,N_497);
or U1425 (N_1425,N_746,N_397);
and U1426 (N_1426,N_67,N_337);
nand U1427 (N_1427,N_305,N_552);
or U1428 (N_1428,N_729,N_227);
and U1429 (N_1429,N_36,N_295);
xnor U1430 (N_1430,N_19,N_223);
xnor U1431 (N_1431,N_202,N_503);
nand U1432 (N_1432,N_414,N_51);
nor U1433 (N_1433,N_7,N_243);
or U1434 (N_1434,N_483,N_583);
and U1435 (N_1435,N_415,N_117);
and U1436 (N_1436,N_469,N_517);
and U1437 (N_1437,N_543,N_187);
or U1438 (N_1438,N_429,N_390);
nand U1439 (N_1439,N_190,N_520);
nor U1440 (N_1440,N_110,N_643);
or U1441 (N_1441,N_120,N_322);
nand U1442 (N_1442,N_698,N_58);
and U1443 (N_1443,N_277,N_144);
nor U1444 (N_1444,N_337,N_603);
nor U1445 (N_1445,N_594,N_277);
xnor U1446 (N_1446,N_565,N_250);
nor U1447 (N_1447,N_501,N_305);
xor U1448 (N_1448,N_276,N_384);
or U1449 (N_1449,N_544,N_731);
nand U1450 (N_1450,N_607,N_415);
nor U1451 (N_1451,N_698,N_127);
nor U1452 (N_1452,N_548,N_270);
nor U1453 (N_1453,N_200,N_593);
xnor U1454 (N_1454,N_169,N_538);
or U1455 (N_1455,N_272,N_98);
or U1456 (N_1456,N_233,N_737);
xor U1457 (N_1457,N_524,N_624);
nand U1458 (N_1458,N_747,N_511);
xor U1459 (N_1459,N_459,N_79);
nand U1460 (N_1460,N_385,N_180);
nor U1461 (N_1461,N_307,N_105);
xnor U1462 (N_1462,N_157,N_72);
nand U1463 (N_1463,N_156,N_277);
nand U1464 (N_1464,N_612,N_8);
nor U1465 (N_1465,N_497,N_16);
or U1466 (N_1466,N_691,N_138);
xor U1467 (N_1467,N_341,N_207);
and U1468 (N_1468,N_176,N_520);
and U1469 (N_1469,N_39,N_706);
and U1470 (N_1470,N_77,N_645);
nand U1471 (N_1471,N_43,N_58);
or U1472 (N_1472,N_16,N_356);
and U1473 (N_1473,N_293,N_553);
and U1474 (N_1474,N_677,N_60);
nor U1475 (N_1475,N_484,N_553);
xnor U1476 (N_1476,N_258,N_462);
nor U1477 (N_1477,N_2,N_187);
nor U1478 (N_1478,N_406,N_652);
and U1479 (N_1479,N_403,N_48);
nor U1480 (N_1480,N_25,N_310);
and U1481 (N_1481,N_515,N_360);
nand U1482 (N_1482,N_126,N_297);
nor U1483 (N_1483,N_134,N_622);
and U1484 (N_1484,N_648,N_16);
nor U1485 (N_1485,N_649,N_651);
xor U1486 (N_1486,N_364,N_171);
nand U1487 (N_1487,N_0,N_642);
nor U1488 (N_1488,N_43,N_301);
nor U1489 (N_1489,N_491,N_668);
or U1490 (N_1490,N_680,N_323);
xnor U1491 (N_1491,N_660,N_120);
nand U1492 (N_1492,N_152,N_23);
nor U1493 (N_1493,N_259,N_642);
nor U1494 (N_1494,N_232,N_606);
or U1495 (N_1495,N_389,N_131);
nand U1496 (N_1496,N_201,N_594);
nand U1497 (N_1497,N_581,N_728);
and U1498 (N_1498,N_615,N_481);
nand U1499 (N_1499,N_684,N_379);
or U1500 (N_1500,N_989,N_785);
nand U1501 (N_1501,N_1418,N_1314);
and U1502 (N_1502,N_1378,N_1143);
xor U1503 (N_1503,N_1078,N_1122);
xor U1504 (N_1504,N_1134,N_1458);
nand U1505 (N_1505,N_1157,N_1474);
nor U1506 (N_1506,N_1127,N_775);
nor U1507 (N_1507,N_1285,N_1469);
nor U1508 (N_1508,N_1217,N_1007);
xor U1509 (N_1509,N_814,N_1245);
nand U1510 (N_1510,N_1296,N_920);
xnor U1511 (N_1511,N_1158,N_784);
and U1512 (N_1512,N_1039,N_937);
nor U1513 (N_1513,N_773,N_1046);
nand U1514 (N_1514,N_1499,N_955);
and U1515 (N_1515,N_798,N_1345);
nor U1516 (N_1516,N_1057,N_1491);
and U1517 (N_1517,N_1337,N_1450);
nand U1518 (N_1518,N_908,N_978);
or U1519 (N_1519,N_847,N_1191);
xnor U1520 (N_1520,N_1045,N_918);
or U1521 (N_1521,N_1249,N_849);
nand U1522 (N_1522,N_1291,N_1124);
or U1523 (N_1523,N_923,N_1253);
xor U1524 (N_1524,N_1148,N_1290);
nor U1525 (N_1525,N_1002,N_1420);
and U1526 (N_1526,N_1184,N_1195);
nand U1527 (N_1527,N_1322,N_870);
or U1528 (N_1528,N_1426,N_1170);
or U1529 (N_1529,N_969,N_794);
xnor U1530 (N_1530,N_1415,N_1343);
nor U1531 (N_1531,N_1106,N_1416);
xor U1532 (N_1532,N_890,N_1279);
nor U1533 (N_1533,N_865,N_990);
nor U1534 (N_1534,N_1301,N_1288);
xor U1535 (N_1535,N_985,N_1094);
nor U1536 (N_1536,N_1451,N_910);
and U1537 (N_1537,N_1029,N_1189);
xnor U1538 (N_1538,N_818,N_988);
or U1539 (N_1539,N_1495,N_1394);
nand U1540 (N_1540,N_1215,N_1321);
and U1541 (N_1541,N_1273,N_850);
xor U1542 (N_1542,N_1088,N_926);
and U1543 (N_1543,N_1477,N_1229);
nor U1544 (N_1544,N_957,N_1333);
nand U1545 (N_1545,N_1284,N_1109);
nand U1546 (N_1546,N_1186,N_1142);
nand U1547 (N_1547,N_858,N_1397);
nor U1548 (N_1548,N_1203,N_1380);
nor U1549 (N_1549,N_1221,N_1409);
nand U1550 (N_1550,N_1270,N_1307);
and U1551 (N_1551,N_1147,N_1208);
xnor U1552 (N_1552,N_1269,N_1072);
xnor U1553 (N_1553,N_1341,N_1062);
nor U1554 (N_1554,N_786,N_1053);
or U1555 (N_1555,N_995,N_1110);
and U1556 (N_1556,N_974,N_1498);
nor U1557 (N_1557,N_1067,N_813);
and U1558 (N_1558,N_885,N_901);
xnor U1559 (N_1559,N_1496,N_991);
xor U1560 (N_1560,N_1452,N_904);
nand U1561 (N_1561,N_1016,N_1370);
xor U1562 (N_1562,N_1299,N_1413);
nor U1563 (N_1563,N_977,N_1289);
nand U1564 (N_1564,N_942,N_919);
xor U1565 (N_1565,N_1459,N_1381);
nand U1566 (N_1566,N_832,N_808);
nand U1567 (N_1567,N_1119,N_1080);
xor U1568 (N_1568,N_1026,N_1254);
or U1569 (N_1569,N_1383,N_1441);
nand U1570 (N_1570,N_1064,N_949);
and U1571 (N_1571,N_928,N_1091);
nor U1572 (N_1572,N_1073,N_799);
or U1573 (N_1573,N_1152,N_833);
nand U1574 (N_1574,N_1017,N_1010);
xnor U1575 (N_1575,N_881,N_1228);
nand U1576 (N_1576,N_1311,N_1406);
nand U1577 (N_1577,N_1049,N_987);
and U1578 (N_1578,N_1081,N_1327);
or U1579 (N_1579,N_780,N_778);
xnor U1580 (N_1580,N_823,N_855);
nor U1581 (N_1581,N_1055,N_1154);
or U1582 (N_1582,N_1070,N_1202);
or U1583 (N_1583,N_779,N_965);
and U1584 (N_1584,N_1271,N_788);
nand U1585 (N_1585,N_1466,N_1464);
nor U1586 (N_1586,N_1144,N_1369);
nor U1587 (N_1587,N_857,N_916);
xor U1588 (N_1588,N_997,N_1357);
and U1589 (N_1589,N_1175,N_1431);
xnor U1590 (N_1590,N_826,N_772);
or U1591 (N_1591,N_1075,N_1163);
nor U1592 (N_1592,N_1281,N_1292);
and U1593 (N_1593,N_860,N_1398);
nand U1594 (N_1594,N_842,N_1190);
nand U1595 (N_1595,N_816,N_1306);
nor U1596 (N_1596,N_1463,N_1318);
nand U1597 (N_1597,N_809,N_1328);
or U1598 (N_1598,N_1137,N_750);
and U1599 (N_1599,N_1389,N_1473);
xnor U1600 (N_1600,N_1128,N_1044);
nor U1601 (N_1601,N_1047,N_1433);
nand U1602 (N_1602,N_970,N_1293);
nand U1603 (N_1603,N_878,N_1353);
nand U1604 (N_1604,N_1324,N_887);
nor U1605 (N_1605,N_934,N_999);
nor U1606 (N_1606,N_1411,N_875);
and U1607 (N_1607,N_962,N_1224);
or U1608 (N_1608,N_992,N_1258);
nand U1609 (N_1609,N_1025,N_1410);
and U1610 (N_1610,N_766,N_1248);
and U1611 (N_1611,N_1034,N_1014);
nand U1612 (N_1612,N_1048,N_1156);
or U1613 (N_1613,N_1437,N_753);
nand U1614 (N_1614,N_966,N_1277);
or U1615 (N_1615,N_1280,N_837);
nor U1616 (N_1616,N_1027,N_1113);
xnor U1617 (N_1617,N_1230,N_1219);
and U1618 (N_1618,N_1188,N_1120);
nor U1619 (N_1619,N_1246,N_1460);
nand U1620 (N_1620,N_1478,N_883);
or U1621 (N_1621,N_1403,N_1022);
nor U1622 (N_1622,N_1182,N_1220);
and U1623 (N_1623,N_1309,N_825);
nor U1624 (N_1624,N_1179,N_895);
nand U1625 (N_1625,N_932,N_1093);
nand U1626 (N_1626,N_1232,N_964);
nor U1627 (N_1627,N_1102,N_956);
nand U1628 (N_1628,N_777,N_1140);
nand U1629 (N_1629,N_915,N_1000);
nand U1630 (N_1630,N_1227,N_1244);
or U1631 (N_1631,N_1283,N_841);
and U1632 (N_1632,N_819,N_776);
and U1633 (N_1633,N_1176,N_1023);
nand U1634 (N_1634,N_1213,N_1334);
nor U1635 (N_1635,N_1085,N_1092);
and U1636 (N_1636,N_1241,N_880);
nor U1637 (N_1637,N_1308,N_1349);
and U1638 (N_1638,N_1196,N_1454);
or U1639 (N_1639,N_947,N_1260);
and U1640 (N_1640,N_864,N_874);
xnor U1641 (N_1641,N_824,N_1461);
nand U1642 (N_1642,N_1272,N_1462);
xnor U1643 (N_1643,N_1356,N_853);
xnor U1644 (N_1644,N_1097,N_968);
xor U1645 (N_1645,N_1139,N_972);
nor U1646 (N_1646,N_1238,N_1236);
or U1647 (N_1647,N_1332,N_1061);
xor U1648 (N_1648,N_1172,N_961);
or U1649 (N_1649,N_1316,N_1368);
or U1650 (N_1650,N_863,N_1342);
xnor U1651 (N_1651,N_872,N_1391);
and U1652 (N_1652,N_1218,N_1050);
xor U1653 (N_1653,N_973,N_954);
nor U1654 (N_1654,N_1468,N_951);
nand U1655 (N_1655,N_764,N_1252);
nor U1656 (N_1656,N_1123,N_1274);
xor U1657 (N_1657,N_886,N_1111);
or U1658 (N_1658,N_1435,N_1302);
xnor U1659 (N_1659,N_1058,N_1261);
and U1660 (N_1660,N_1065,N_1011);
xor U1661 (N_1661,N_802,N_1497);
nor U1662 (N_1662,N_1231,N_1024);
nand U1663 (N_1663,N_1432,N_790);
and U1664 (N_1664,N_1362,N_804);
xor U1665 (N_1665,N_1425,N_948);
nand U1666 (N_1666,N_1040,N_1372);
nor U1667 (N_1667,N_845,N_1376);
and U1668 (N_1668,N_1149,N_1367);
nor U1669 (N_1669,N_940,N_1087);
nand U1670 (N_1670,N_1449,N_1226);
xnor U1671 (N_1671,N_1185,N_1256);
and U1672 (N_1672,N_1052,N_754);
and U1673 (N_1673,N_755,N_1197);
or U1674 (N_1674,N_1038,N_1257);
or U1675 (N_1675,N_1255,N_828);
and U1676 (N_1676,N_1103,N_1090);
and U1677 (N_1677,N_938,N_867);
and U1678 (N_1678,N_1446,N_771);
and U1679 (N_1679,N_791,N_1338);
xnor U1680 (N_1680,N_907,N_1076);
nor U1681 (N_1681,N_861,N_1493);
nand U1682 (N_1682,N_1159,N_1247);
or U1683 (N_1683,N_1297,N_1096);
nor U1684 (N_1684,N_797,N_994);
nand U1685 (N_1685,N_1212,N_1239);
xnor U1686 (N_1686,N_758,N_840);
or U1687 (N_1687,N_1487,N_1206);
or U1688 (N_1688,N_1222,N_1108);
and U1689 (N_1689,N_1167,N_1001);
or U1690 (N_1690,N_1069,N_1282);
or U1691 (N_1691,N_1135,N_1201);
or U1692 (N_1692,N_1417,N_1198);
xnor U1693 (N_1693,N_789,N_752);
and U1694 (N_1694,N_1205,N_1374);
and U1695 (N_1695,N_1440,N_1412);
and U1696 (N_1696,N_1099,N_811);
or U1697 (N_1697,N_896,N_1329);
nand U1698 (N_1698,N_927,N_1174);
xnor U1699 (N_1699,N_1265,N_759);
nor U1700 (N_1700,N_1267,N_1118);
nand U1701 (N_1701,N_1481,N_767);
nor U1702 (N_1702,N_1408,N_1177);
or U1703 (N_1703,N_1371,N_1077);
and U1704 (N_1704,N_993,N_1181);
xnor U1705 (N_1705,N_882,N_1428);
nand U1706 (N_1706,N_876,N_1275);
or U1707 (N_1707,N_1008,N_1216);
and U1708 (N_1708,N_1330,N_909);
and U1709 (N_1709,N_821,N_820);
or U1710 (N_1710,N_1107,N_1171);
and U1711 (N_1711,N_1340,N_905);
nand U1712 (N_1712,N_1161,N_1350);
xor U1713 (N_1713,N_1325,N_975);
and U1714 (N_1714,N_751,N_774);
nand U1715 (N_1715,N_1490,N_792);
xnor U1716 (N_1716,N_950,N_1482);
xnor U1717 (N_1717,N_877,N_980);
xor U1718 (N_1718,N_1373,N_1287);
xnor U1719 (N_1719,N_1492,N_998);
nand U1720 (N_1720,N_1488,N_1015);
or U1721 (N_1721,N_1209,N_946);
nor U1722 (N_1722,N_1089,N_859);
nor U1723 (N_1723,N_1095,N_1243);
or U1724 (N_1724,N_1155,N_756);
or U1725 (N_1725,N_930,N_1145);
nand U1726 (N_1726,N_1384,N_1200);
and U1727 (N_1727,N_1033,N_871);
nand U1728 (N_1728,N_1169,N_924);
and U1729 (N_1729,N_1294,N_1315);
nor U1730 (N_1730,N_1347,N_1377);
and U1731 (N_1731,N_1323,N_1268);
nor U1732 (N_1732,N_1125,N_1427);
nor U1733 (N_1733,N_769,N_1443);
xnor U1734 (N_1734,N_1422,N_787);
nor U1735 (N_1735,N_1402,N_1178);
and U1736 (N_1736,N_1051,N_1304);
xor U1737 (N_1737,N_827,N_976);
and U1738 (N_1738,N_931,N_1471);
or U1739 (N_1739,N_761,N_914);
nor U1740 (N_1740,N_1138,N_1259);
or U1741 (N_1741,N_936,N_1153);
or U1742 (N_1742,N_1086,N_1348);
nand U1743 (N_1743,N_1021,N_1194);
xnor U1744 (N_1744,N_1313,N_903);
nand U1745 (N_1745,N_1278,N_971);
and U1746 (N_1746,N_1352,N_1183);
and U1747 (N_1747,N_1424,N_1164);
nand U1748 (N_1748,N_1475,N_1317);
and U1749 (N_1749,N_862,N_803);
xnor U1750 (N_1750,N_783,N_800);
nand U1751 (N_1751,N_838,N_1359);
nand U1752 (N_1752,N_1436,N_1331);
xor U1753 (N_1753,N_917,N_935);
xor U1754 (N_1754,N_815,N_1013);
xor U1755 (N_1755,N_1004,N_793);
nor U1756 (N_1756,N_1121,N_1361);
or U1757 (N_1757,N_806,N_1366);
and U1758 (N_1758,N_1438,N_817);
and U1759 (N_1759,N_944,N_1214);
or U1760 (N_1760,N_967,N_981);
nor U1761 (N_1761,N_1115,N_1430);
and U1762 (N_1762,N_1117,N_1100);
or U1763 (N_1763,N_913,N_760);
or U1764 (N_1764,N_1101,N_835);
nor U1765 (N_1765,N_1160,N_1303);
or U1766 (N_1766,N_1455,N_1305);
or U1767 (N_1767,N_1453,N_1083);
and U1768 (N_1768,N_1396,N_1421);
xnor U1769 (N_1769,N_831,N_1434);
nand U1770 (N_1770,N_1346,N_1358);
nand U1771 (N_1771,N_1063,N_979);
nor U1772 (N_1772,N_1484,N_1030);
and U1773 (N_1773,N_1479,N_952);
nand U1774 (N_1774,N_884,N_1112);
xnor U1775 (N_1775,N_1400,N_854);
xor U1776 (N_1776,N_822,N_851);
and U1777 (N_1777,N_929,N_925);
or U1778 (N_1778,N_1326,N_844);
or U1779 (N_1779,N_1448,N_1079);
xor U1780 (N_1780,N_1365,N_1028);
nor U1781 (N_1781,N_1192,N_1130);
xnor U1782 (N_1782,N_906,N_1439);
or U1783 (N_1783,N_1129,N_830);
and U1784 (N_1784,N_1251,N_1150);
xor U1785 (N_1785,N_1066,N_1233);
xnor U1786 (N_1786,N_1242,N_1060);
or U1787 (N_1787,N_781,N_866);
nand U1788 (N_1788,N_1019,N_1355);
xor U1789 (N_1789,N_1465,N_1003);
nor U1790 (N_1790,N_1489,N_939);
and U1791 (N_1791,N_1467,N_943);
nand U1792 (N_1792,N_1401,N_983);
nor U1793 (N_1793,N_1476,N_899);
or U1794 (N_1794,N_836,N_941);
nor U1795 (N_1795,N_1470,N_1031);
nor U1796 (N_1796,N_891,N_1382);
nor U1797 (N_1797,N_768,N_1210);
and U1798 (N_1798,N_856,N_1390);
nand U1799 (N_1799,N_1483,N_1295);
nor U1800 (N_1800,N_1320,N_1056);
xor U1801 (N_1801,N_1006,N_1054);
nand U1802 (N_1802,N_1180,N_1354);
nand U1803 (N_1803,N_1018,N_1360);
or U1804 (N_1804,N_888,N_1419);
nor U1805 (N_1805,N_1486,N_1041);
nor U1806 (N_1806,N_1235,N_810);
and U1807 (N_1807,N_1131,N_1379);
xor U1808 (N_1808,N_960,N_1363);
nor U1809 (N_1809,N_1351,N_889);
nand U1810 (N_1810,N_958,N_1104);
xnor U1811 (N_1811,N_1312,N_801);
and U1812 (N_1812,N_1036,N_795);
xnor U1813 (N_1813,N_894,N_1429);
xnor U1814 (N_1814,N_1445,N_1074);
xnor U1815 (N_1815,N_1375,N_1114);
nor U1816 (N_1816,N_1263,N_996);
xnor U1817 (N_1817,N_1187,N_911);
xnor U1818 (N_1818,N_1266,N_1395);
xor U1819 (N_1819,N_902,N_765);
nor U1820 (N_1820,N_843,N_1204);
nand U1821 (N_1821,N_1151,N_839);
or U1822 (N_1822,N_897,N_1472);
and U1823 (N_1823,N_1193,N_1240);
or U1824 (N_1824,N_912,N_1298);
and U1825 (N_1825,N_1387,N_1300);
or U1826 (N_1826,N_1494,N_1414);
and U1827 (N_1827,N_1457,N_1032);
xnor U1828 (N_1828,N_1105,N_1250);
nand U1829 (N_1829,N_762,N_1173);
xnor U1830 (N_1830,N_829,N_1082);
and U1831 (N_1831,N_770,N_1335);
and U1832 (N_1832,N_1392,N_1005);
nand U1833 (N_1833,N_1084,N_873);
or U1834 (N_1834,N_986,N_1168);
or U1835 (N_1835,N_922,N_898);
nand U1836 (N_1836,N_1166,N_1407);
and U1837 (N_1837,N_1405,N_1447);
or U1838 (N_1838,N_1264,N_1234);
xnor U1839 (N_1839,N_1225,N_1286);
nor U1840 (N_1840,N_1146,N_1199);
xor U1841 (N_1841,N_1132,N_1037);
and U1842 (N_1842,N_1035,N_1393);
nor U1843 (N_1843,N_1344,N_1068);
xnor U1844 (N_1844,N_848,N_1126);
or U1845 (N_1845,N_812,N_1310);
nand U1846 (N_1846,N_1043,N_1456);
nor U1847 (N_1847,N_1276,N_1020);
nand U1848 (N_1848,N_963,N_1042);
or U1849 (N_1849,N_1399,N_763);
xor U1850 (N_1850,N_805,N_1336);
nor U1851 (N_1851,N_1385,N_868);
xor U1852 (N_1852,N_1136,N_893);
nor U1853 (N_1853,N_959,N_1262);
and U1854 (N_1854,N_796,N_1404);
and U1855 (N_1855,N_1319,N_1386);
and U1856 (N_1856,N_945,N_1223);
or U1857 (N_1857,N_1165,N_1207);
nor U1858 (N_1858,N_1480,N_1009);
nor U1859 (N_1859,N_982,N_933);
nor U1860 (N_1860,N_869,N_1442);
or U1861 (N_1861,N_1012,N_1211);
or U1862 (N_1862,N_984,N_1444);
nor U1863 (N_1863,N_852,N_1388);
or U1864 (N_1864,N_807,N_846);
nand U1865 (N_1865,N_1098,N_1141);
xor U1866 (N_1866,N_1162,N_900);
nand U1867 (N_1867,N_1423,N_1485);
nor U1868 (N_1868,N_953,N_1364);
or U1869 (N_1869,N_892,N_1059);
nand U1870 (N_1870,N_1133,N_1116);
or U1871 (N_1871,N_834,N_1237);
nor U1872 (N_1872,N_1339,N_921);
or U1873 (N_1873,N_757,N_1071);
nand U1874 (N_1874,N_879,N_782);
nand U1875 (N_1875,N_1268,N_986);
or U1876 (N_1876,N_1187,N_814);
or U1877 (N_1877,N_953,N_1043);
nor U1878 (N_1878,N_905,N_1057);
xnor U1879 (N_1879,N_1310,N_1020);
xor U1880 (N_1880,N_776,N_788);
nor U1881 (N_1881,N_993,N_1383);
nor U1882 (N_1882,N_1317,N_1450);
nor U1883 (N_1883,N_882,N_1319);
or U1884 (N_1884,N_1374,N_841);
xor U1885 (N_1885,N_838,N_999);
nand U1886 (N_1886,N_1106,N_1115);
nand U1887 (N_1887,N_1397,N_786);
nand U1888 (N_1888,N_1339,N_1499);
nor U1889 (N_1889,N_978,N_1040);
xor U1890 (N_1890,N_1487,N_1382);
and U1891 (N_1891,N_1199,N_1009);
xor U1892 (N_1892,N_1056,N_1370);
nand U1893 (N_1893,N_917,N_1173);
or U1894 (N_1894,N_1250,N_849);
nand U1895 (N_1895,N_1499,N_1360);
nand U1896 (N_1896,N_1087,N_1013);
or U1897 (N_1897,N_1365,N_965);
nand U1898 (N_1898,N_973,N_1312);
nand U1899 (N_1899,N_837,N_1222);
and U1900 (N_1900,N_1215,N_781);
xnor U1901 (N_1901,N_1039,N_1229);
or U1902 (N_1902,N_888,N_796);
or U1903 (N_1903,N_822,N_1223);
nand U1904 (N_1904,N_1304,N_790);
nand U1905 (N_1905,N_801,N_1397);
nor U1906 (N_1906,N_1394,N_785);
and U1907 (N_1907,N_1476,N_1498);
nor U1908 (N_1908,N_1009,N_955);
nand U1909 (N_1909,N_1125,N_1487);
xnor U1910 (N_1910,N_1125,N_881);
or U1911 (N_1911,N_1019,N_1081);
nand U1912 (N_1912,N_1288,N_1322);
nand U1913 (N_1913,N_1046,N_959);
nor U1914 (N_1914,N_1465,N_1351);
xor U1915 (N_1915,N_1219,N_768);
nor U1916 (N_1916,N_1442,N_1210);
or U1917 (N_1917,N_1308,N_1138);
or U1918 (N_1918,N_780,N_828);
nand U1919 (N_1919,N_1464,N_900);
or U1920 (N_1920,N_867,N_842);
and U1921 (N_1921,N_1449,N_844);
nand U1922 (N_1922,N_1174,N_1459);
xor U1923 (N_1923,N_761,N_1439);
nand U1924 (N_1924,N_795,N_860);
nor U1925 (N_1925,N_1014,N_1101);
or U1926 (N_1926,N_1475,N_1401);
nor U1927 (N_1927,N_863,N_1385);
nand U1928 (N_1928,N_1031,N_1362);
nor U1929 (N_1929,N_958,N_1437);
and U1930 (N_1930,N_877,N_1067);
and U1931 (N_1931,N_1142,N_938);
nor U1932 (N_1932,N_1448,N_1290);
nand U1933 (N_1933,N_1256,N_1322);
or U1934 (N_1934,N_1085,N_1442);
nor U1935 (N_1935,N_989,N_1301);
and U1936 (N_1936,N_1200,N_954);
nor U1937 (N_1937,N_1111,N_1410);
nand U1938 (N_1938,N_1088,N_804);
or U1939 (N_1939,N_1363,N_1075);
or U1940 (N_1940,N_1483,N_1055);
and U1941 (N_1941,N_1214,N_871);
nor U1942 (N_1942,N_1305,N_1428);
nand U1943 (N_1943,N_824,N_1483);
and U1944 (N_1944,N_1272,N_794);
or U1945 (N_1945,N_1409,N_1141);
and U1946 (N_1946,N_1067,N_903);
nand U1947 (N_1947,N_1087,N_1381);
nor U1948 (N_1948,N_985,N_1122);
xnor U1949 (N_1949,N_860,N_1488);
or U1950 (N_1950,N_886,N_1076);
nand U1951 (N_1951,N_1227,N_1406);
nor U1952 (N_1952,N_1054,N_1226);
or U1953 (N_1953,N_1178,N_1351);
nand U1954 (N_1954,N_822,N_1132);
nand U1955 (N_1955,N_1451,N_1422);
nand U1956 (N_1956,N_1085,N_1157);
nor U1957 (N_1957,N_960,N_830);
and U1958 (N_1958,N_1158,N_1484);
nand U1959 (N_1959,N_769,N_1035);
nor U1960 (N_1960,N_1299,N_1175);
nand U1961 (N_1961,N_1050,N_1163);
xnor U1962 (N_1962,N_1392,N_1310);
nor U1963 (N_1963,N_891,N_1040);
or U1964 (N_1964,N_996,N_1473);
or U1965 (N_1965,N_1481,N_1249);
nand U1966 (N_1966,N_752,N_1069);
or U1967 (N_1967,N_886,N_1007);
nand U1968 (N_1968,N_1436,N_1130);
and U1969 (N_1969,N_764,N_1337);
xor U1970 (N_1970,N_1273,N_1240);
and U1971 (N_1971,N_1202,N_877);
xnor U1972 (N_1972,N_1193,N_1110);
nand U1973 (N_1973,N_823,N_1311);
and U1974 (N_1974,N_865,N_1256);
nand U1975 (N_1975,N_982,N_1441);
and U1976 (N_1976,N_941,N_886);
xnor U1977 (N_1977,N_950,N_854);
nor U1978 (N_1978,N_943,N_1140);
nor U1979 (N_1979,N_1499,N_1110);
xnor U1980 (N_1980,N_1135,N_892);
nand U1981 (N_1981,N_1226,N_1295);
nand U1982 (N_1982,N_1414,N_1249);
or U1983 (N_1983,N_1371,N_951);
or U1984 (N_1984,N_1308,N_1171);
nand U1985 (N_1985,N_1385,N_1376);
nor U1986 (N_1986,N_1052,N_859);
nand U1987 (N_1987,N_1014,N_1052);
xnor U1988 (N_1988,N_1290,N_1036);
nand U1989 (N_1989,N_848,N_1234);
nand U1990 (N_1990,N_1283,N_1181);
xor U1991 (N_1991,N_1012,N_1497);
and U1992 (N_1992,N_1491,N_1459);
nand U1993 (N_1993,N_1129,N_1213);
nor U1994 (N_1994,N_1407,N_1000);
nand U1995 (N_1995,N_1332,N_810);
or U1996 (N_1996,N_1481,N_1318);
nor U1997 (N_1997,N_880,N_1310);
nand U1998 (N_1998,N_1085,N_1342);
and U1999 (N_1999,N_1239,N_1469);
and U2000 (N_2000,N_783,N_1125);
and U2001 (N_2001,N_1439,N_1191);
xor U2002 (N_2002,N_866,N_1064);
nand U2003 (N_2003,N_794,N_860);
xnor U2004 (N_2004,N_1403,N_1390);
and U2005 (N_2005,N_1257,N_1108);
xor U2006 (N_2006,N_1036,N_841);
and U2007 (N_2007,N_944,N_1149);
nor U2008 (N_2008,N_1400,N_1213);
and U2009 (N_2009,N_1092,N_1106);
xor U2010 (N_2010,N_1479,N_1404);
xor U2011 (N_2011,N_1457,N_1405);
xor U2012 (N_2012,N_1241,N_785);
or U2013 (N_2013,N_915,N_1357);
nor U2014 (N_2014,N_1141,N_1289);
nor U2015 (N_2015,N_990,N_956);
or U2016 (N_2016,N_1413,N_1082);
nor U2017 (N_2017,N_1150,N_1392);
or U2018 (N_2018,N_1345,N_1423);
nand U2019 (N_2019,N_1437,N_1414);
and U2020 (N_2020,N_1211,N_799);
xor U2021 (N_2021,N_1042,N_838);
nor U2022 (N_2022,N_1325,N_1009);
nor U2023 (N_2023,N_1141,N_1077);
and U2024 (N_2024,N_1250,N_1433);
nor U2025 (N_2025,N_1392,N_972);
nand U2026 (N_2026,N_790,N_965);
nand U2027 (N_2027,N_1407,N_1191);
nand U2028 (N_2028,N_813,N_775);
and U2029 (N_2029,N_1348,N_1304);
nor U2030 (N_2030,N_903,N_1477);
xor U2031 (N_2031,N_1420,N_833);
or U2032 (N_2032,N_1369,N_943);
or U2033 (N_2033,N_1084,N_958);
nor U2034 (N_2034,N_1383,N_886);
or U2035 (N_2035,N_1006,N_1328);
and U2036 (N_2036,N_847,N_1292);
or U2037 (N_2037,N_990,N_1482);
nand U2038 (N_2038,N_1143,N_1152);
nor U2039 (N_2039,N_1190,N_758);
nand U2040 (N_2040,N_1364,N_1335);
nor U2041 (N_2041,N_1159,N_1141);
or U2042 (N_2042,N_1049,N_1394);
or U2043 (N_2043,N_874,N_1299);
and U2044 (N_2044,N_896,N_1169);
nand U2045 (N_2045,N_759,N_1054);
nor U2046 (N_2046,N_993,N_1013);
nor U2047 (N_2047,N_1287,N_1464);
nor U2048 (N_2048,N_1353,N_1455);
and U2049 (N_2049,N_1216,N_957);
nor U2050 (N_2050,N_1488,N_899);
xor U2051 (N_2051,N_842,N_1416);
and U2052 (N_2052,N_1362,N_930);
nand U2053 (N_2053,N_1392,N_965);
nor U2054 (N_2054,N_1249,N_985);
and U2055 (N_2055,N_1060,N_1259);
xnor U2056 (N_2056,N_820,N_1228);
and U2057 (N_2057,N_1043,N_1445);
and U2058 (N_2058,N_1360,N_1449);
xor U2059 (N_2059,N_1202,N_849);
xnor U2060 (N_2060,N_940,N_781);
or U2061 (N_2061,N_922,N_1440);
nor U2062 (N_2062,N_797,N_804);
nor U2063 (N_2063,N_873,N_1055);
or U2064 (N_2064,N_1462,N_1323);
nor U2065 (N_2065,N_987,N_1495);
nor U2066 (N_2066,N_1028,N_1374);
xnor U2067 (N_2067,N_1143,N_923);
nor U2068 (N_2068,N_1402,N_1486);
or U2069 (N_2069,N_1172,N_1187);
and U2070 (N_2070,N_1399,N_989);
or U2071 (N_2071,N_1293,N_1299);
xnor U2072 (N_2072,N_1079,N_864);
and U2073 (N_2073,N_1206,N_759);
and U2074 (N_2074,N_1300,N_951);
xnor U2075 (N_2075,N_1255,N_950);
nand U2076 (N_2076,N_899,N_967);
and U2077 (N_2077,N_958,N_1063);
nand U2078 (N_2078,N_1356,N_886);
or U2079 (N_2079,N_1301,N_1163);
or U2080 (N_2080,N_802,N_1332);
xnor U2081 (N_2081,N_1131,N_1040);
nor U2082 (N_2082,N_1082,N_1150);
nand U2083 (N_2083,N_780,N_874);
nand U2084 (N_2084,N_771,N_1261);
and U2085 (N_2085,N_1342,N_967);
xor U2086 (N_2086,N_1253,N_767);
or U2087 (N_2087,N_1008,N_1143);
and U2088 (N_2088,N_1073,N_755);
xor U2089 (N_2089,N_1224,N_1490);
nand U2090 (N_2090,N_753,N_883);
xnor U2091 (N_2091,N_782,N_1375);
or U2092 (N_2092,N_1499,N_1007);
nor U2093 (N_2093,N_1431,N_914);
or U2094 (N_2094,N_1348,N_1321);
nor U2095 (N_2095,N_934,N_1167);
nand U2096 (N_2096,N_1013,N_851);
or U2097 (N_2097,N_944,N_937);
nor U2098 (N_2098,N_901,N_1362);
or U2099 (N_2099,N_1375,N_908);
or U2100 (N_2100,N_1339,N_1168);
or U2101 (N_2101,N_1344,N_941);
nor U2102 (N_2102,N_1044,N_1468);
and U2103 (N_2103,N_1167,N_1228);
and U2104 (N_2104,N_777,N_1418);
or U2105 (N_2105,N_946,N_1466);
xor U2106 (N_2106,N_949,N_1129);
and U2107 (N_2107,N_1362,N_1407);
and U2108 (N_2108,N_930,N_1168);
or U2109 (N_2109,N_1157,N_1137);
xor U2110 (N_2110,N_821,N_986);
nor U2111 (N_2111,N_1282,N_1257);
nand U2112 (N_2112,N_926,N_877);
and U2113 (N_2113,N_976,N_982);
or U2114 (N_2114,N_887,N_1338);
xor U2115 (N_2115,N_1198,N_1168);
nor U2116 (N_2116,N_978,N_1409);
or U2117 (N_2117,N_953,N_842);
or U2118 (N_2118,N_1002,N_968);
or U2119 (N_2119,N_1101,N_1474);
xor U2120 (N_2120,N_1480,N_936);
and U2121 (N_2121,N_1404,N_944);
xnor U2122 (N_2122,N_1259,N_783);
and U2123 (N_2123,N_1044,N_860);
nor U2124 (N_2124,N_1422,N_1041);
and U2125 (N_2125,N_1415,N_985);
nor U2126 (N_2126,N_1098,N_1491);
or U2127 (N_2127,N_895,N_1013);
and U2128 (N_2128,N_1331,N_1322);
xnor U2129 (N_2129,N_1434,N_1236);
xor U2130 (N_2130,N_1372,N_831);
or U2131 (N_2131,N_1323,N_781);
nor U2132 (N_2132,N_986,N_1242);
xnor U2133 (N_2133,N_757,N_1215);
nand U2134 (N_2134,N_1369,N_1388);
xnor U2135 (N_2135,N_1221,N_790);
nand U2136 (N_2136,N_1444,N_1291);
and U2137 (N_2137,N_904,N_987);
and U2138 (N_2138,N_1420,N_996);
xor U2139 (N_2139,N_1086,N_967);
nor U2140 (N_2140,N_1287,N_1401);
and U2141 (N_2141,N_1391,N_1498);
and U2142 (N_2142,N_1160,N_1027);
and U2143 (N_2143,N_961,N_1232);
nor U2144 (N_2144,N_826,N_1227);
nand U2145 (N_2145,N_1490,N_1457);
or U2146 (N_2146,N_840,N_1499);
nor U2147 (N_2147,N_1219,N_1211);
and U2148 (N_2148,N_930,N_951);
or U2149 (N_2149,N_1365,N_799);
xor U2150 (N_2150,N_1169,N_827);
and U2151 (N_2151,N_1372,N_1338);
and U2152 (N_2152,N_1452,N_1383);
or U2153 (N_2153,N_1479,N_1041);
and U2154 (N_2154,N_1230,N_977);
or U2155 (N_2155,N_1392,N_1213);
nand U2156 (N_2156,N_1265,N_913);
or U2157 (N_2157,N_890,N_1097);
nand U2158 (N_2158,N_1038,N_996);
nor U2159 (N_2159,N_903,N_1328);
or U2160 (N_2160,N_985,N_1464);
and U2161 (N_2161,N_1159,N_1484);
or U2162 (N_2162,N_865,N_855);
nor U2163 (N_2163,N_800,N_1431);
nor U2164 (N_2164,N_1166,N_1471);
nor U2165 (N_2165,N_784,N_758);
and U2166 (N_2166,N_1000,N_799);
nand U2167 (N_2167,N_772,N_999);
nor U2168 (N_2168,N_990,N_1421);
nor U2169 (N_2169,N_782,N_1453);
and U2170 (N_2170,N_1185,N_833);
xor U2171 (N_2171,N_1299,N_1049);
nand U2172 (N_2172,N_1338,N_1047);
and U2173 (N_2173,N_1010,N_1304);
xnor U2174 (N_2174,N_1161,N_1168);
xnor U2175 (N_2175,N_1114,N_967);
xor U2176 (N_2176,N_1415,N_861);
xnor U2177 (N_2177,N_877,N_932);
nand U2178 (N_2178,N_862,N_752);
nand U2179 (N_2179,N_1453,N_1420);
nand U2180 (N_2180,N_1198,N_1125);
or U2181 (N_2181,N_1047,N_1423);
nand U2182 (N_2182,N_1075,N_1347);
or U2183 (N_2183,N_1117,N_1043);
nor U2184 (N_2184,N_971,N_843);
or U2185 (N_2185,N_1000,N_1071);
or U2186 (N_2186,N_912,N_1109);
xnor U2187 (N_2187,N_1483,N_1456);
and U2188 (N_2188,N_1077,N_775);
nand U2189 (N_2189,N_856,N_755);
and U2190 (N_2190,N_1390,N_1072);
xor U2191 (N_2191,N_873,N_1185);
nor U2192 (N_2192,N_1217,N_1130);
nand U2193 (N_2193,N_894,N_1358);
nor U2194 (N_2194,N_1352,N_1460);
or U2195 (N_2195,N_1091,N_1055);
nor U2196 (N_2196,N_1296,N_857);
nor U2197 (N_2197,N_772,N_1001);
xnor U2198 (N_2198,N_1255,N_817);
or U2199 (N_2199,N_1099,N_945);
and U2200 (N_2200,N_845,N_1359);
nor U2201 (N_2201,N_1163,N_1055);
xnor U2202 (N_2202,N_772,N_960);
nand U2203 (N_2203,N_843,N_1465);
nand U2204 (N_2204,N_1125,N_893);
nand U2205 (N_2205,N_1007,N_933);
nand U2206 (N_2206,N_1224,N_1340);
nor U2207 (N_2207,N_1429,N_1268);
xnor U2208 (N_2208,N_979,N_1347);
nand U2209 (N_2209,N_1251,N_919);
nor U2210 (N_2210,N_1367,N_922);
nand U2211 (N_2211,N_1247,N_1465);
and U2212 (N_2212,N_1149,N_1392);
and U2213 (N_2213,N_837,N_1457);
nand U2214 (N_2214,N_1485,N_769);
nor U2215 (N_2215,N_814,N_1031);
or U2216 (N_2216,N_1484,N_906);
and U2217 (N_2217,N_760,N_1098);
or U2218 (N_2218,N_1353,N_932);
xnor U2219 (N_2219,N_838,N_1481);
nor U2220 (N_2220,N_1064,N_1301);
or U2221 (N_2221,N_1449,N_771);
nand U2222 (N_2222,N_1425,N_1291);
and U2223 (N_2223,N_819,N_1111);
xor U2224 (N_2224,N_1483,N_994);
or U2225 (N_2225,N_1238,N_1103);
or U2226 (N_2226,N_1102,N_879);
nor U2227 (N_2227,N_1353,N_1367);
nor U2228 (N_2228,N_1418,N_1444);
nor U2229 (N_2229,N_968,N_1334);
xnor U2230 (N_2230,N_1346,N_1018);
nor U2231 (N_2231,N_1228,N_1421);
and U2232 (N_2232,N_959,N_1386);
nor U2233 (N_2233,N_1018,N_1004);
or U2234 (N_2234,N_1162,N_1151);
and U2235 (N_2235,N_1073,N_913);
xor U2236 (N_2236,N_1356,N_765);
nor U2237 (N_2237,N_1459,N_1145);
nor U2238 (N_2238,N_1315,N_876);
nor U2239 (N_2239,N_1182,N_1468);
nand U2240 (N_2240,N_1217,N_1385);
nor U2241 (N_2241,N_923,N_1380);
nand U2242 (N_2242,N_1022,N_1435);
xor U2243 (N_2243,N_1341,N_1013);
or U2244 (N_2244,N_1257,N_1254);
nor U2245 (N_2245,N_895,N_1479);
or U2246 (N_2246,N_1116,N_1444);
and U2247 (N_2247,N_1193,N_975);
nor U2248 (N_2248,N_810,N_822);
nor U2249 (N_2249,N_951,N_1221);
and U2250 (N_2250,N_1688,N_1707);
or U2251 (N_2251,N_1757,N_1594);
xor U2252 (N_2252,N_1886,N_1817);
and U2253 (N_2253,N_1950,N_2156);
nand U2254 (N_2254,N_1796,N_1839);
nand U2255 (N_2255,N_1939,N_2058);
or U2256 (N_2256,N_2130,N_1765);
nor U2257 (N_2257,N_2001,N_2008);
nor U2258 (N_2258,N_1769,N_2135);
or U2259 (N_2259,N_2121,N_1721);
nor U2260 (N_2260,N_1596,N_1531);
nand U2261 (N_2261,N_1890,N_1872);
nor U2262 (N_2262,N_2122,N_1927);
or U2263 (N_2263,N_1789,N_2101);
or U2264 (N_2264,N_2212,N_1970);
xor U2265 (N_2265,N_2023,N_1589);
xnor U2266 (N_2266,N_1763,N_1510);
and U2267 (N_2267,N_1916,N_2225);
nand U2268 (N_2268,N_1631,N_2091);
nor U2269 (N_2269,N_1928,N_1802);
nor U2270 (N_2270,N_1552,N_1961);
nor U2271 (N_2271,N_1785,N_1737);
or U2272 (N_2272,N_1523,N_2035);
and U2273 (N_2273,N_1585,N_1893);
nor U2274 (N_2274,N_2235,N_1827);
nand U2275 (N_2275,N_1692,N_1912);
nor U2276 (N_2276,N_1726,N_1808);
nand U2277 (N_2277,N_2024,N_1851);
nand U2278 (N_2278,N_2015,N_1674);
xnor U2279 (N_2279,N_1693,N_1551);
or U2280 (N_2280,N_2173,N_1669);
nor U2281 (N_2281,N_1538,N_2188);
xor U2282 (N_2282,N_1843,N_2016);
or U2283 (N_2283,N_1899,N_1641);
xor U2284 (N_2284,N_1925,N_1597);
and U2285 (N_2285,N_2195,N_2017);
nor U2286 (N_2286,N_2103,N_1579);
nand U2287 (N_2287,N_1629,N_2020);
xnor U2288 (N_2288,N_1547,N_1984);
nand U2289 (N_2289,N_1572,N_1553);
or U2290 (N_2290,N_1718,N_1979);
and U2291 (N_2291,N_2033,N_1951);
nand U2292 (N_2292,N_1573,N_1710);
xnor U2293 (N_2293,N_1588,N_1584);
xor U2294 (N_2294,N_1704,N_1617);
xor U2295 (N_2295,N_1744,N_2192);
and U2296 (N_2296,N_2113,N_2233);
or U2297 (N_2297,N_1847,N_1515);
xor U2298 (N_2298,N_1766,N_2232);
and U2299 (N_2299,N_1842,N_1840);
and U2300 (N_2300,N_1870,N_1557);
or U2301 (N_2301,N_1971,N_1920);
nor U2302 (N_2302,N_1603,N_2168);
and U2303 (N_2303,N_2115,N_2175);
and U2304 (N_2304,N_1580,N_1944);
nor U2305 (N_2305,N_2067,N_2132);
nand U2306 (N_2306,N_1694,N_2234);
nand U2307 (N_2307,N_1772,N_1773);
or U2308 (N_2308,N_1712,N_2134);
and U2309 (N_2309,N_1517,N_1781);
and U2310 (N_2310,N_1685,N_1564);
nor U2311 (N_2311,N_1754,N_1706);
or U2312 (N_2312,N_1592,N_2145);
or U2313 (N_2313,N_1982,N_1749);
nand U2314 (N_2314,N_1973,N_1683);
and U2315 (N_2315,N_2153,N_1625);
xnor U2316 (N_2316,N_2095,N_1730);
or U2317 (N_2317,N_2037,N_2018);
nor U2318 (N_2318,N_2204,N_1559);
and U2319 (N_2319,N_2026,N_1977);
xnor U2320 (N_2320,N_2075,N_1638);
nand U2321 (N_2321,N_1963,N_1917);
and U2322 (N_2322,N_1965,N_2106);
nand U2323 (N_2323,N_1775,N_2177);
xnor U2324 (N_2324,N_2073,N_2083);
nor U2325 (N_2325,N_1924,N_2158);
or U2326 (N_2326,N_2150,N_2244);
and U2327 (N_2327,N_1941,N_1569);
nor U2328 (N_2328,N_1501,N_1663);
and U2329 (N_2329,N_1732,N_1864);
nand U2330 (N_2330,N_2201,N_2111);
xnor U2331 (N_2331,N_1975,N_1542);
nor U2332 (N_2332,N_1606,N_1915);
xor U2333 (N_2333,N_1505,N_1703);
and U2334 (N_2334,N_2102,N_2151);
and U2335 (N_2335,N_1891,N_1616);
and U2336 (N_2336,N_2059,N_1659);
xor U2337 (N_2337,N_2193,N_2000);
nor U2338 (N_2338,N_1932,N_1823);
or U2339 (N_2339,N_2057,N_2160);
nor U2340 (N_2340,N_1664,N_2055);
nand U2341 (N_2341,N_1957,N_2239);
xor U2342 (N_2342,N_1904,N_2143);
or U2343 (N_2343,N_1896,N_1881);
xor U2344 (N_2344,N_2074,N_1605);
and U2345 (N_2345,N_1648,N_1562);
or U2346 (N_2346,N_2162,N_1675);
and U2347 (N_2347,N_1846,N_1987);
xor U2348 (N_2348,N_2219,N_1980);
nor U2349 (N_2349,N_1770,N_1554);
nand U2350 (N_2350,N_1504,N_1623);
nor U2351 (N_2351,N_1956,N_1993);
nand U2352 (N_2352,N_1998,N_2155);
and U2353 (N_2353,N_2199,N_1608);
and U2354 (N_2354,N_1621,N_1645);
and U2355 (N_2355,N_2220,N_1709);
xnor U2356 (N_2356,N_1780,N_2187);
nand U2357 (N_2357,N_2003,N_1892);
nor U2358 (N_2358,N_1880,N_2021);
or U2359 (N_2359,N_1844,N_1529);
and U2360 (N_2360,N_1946,N_1978);
or U2361 (N_2361,N_1705,N_2078);
nand U2362 (N_2362,N_1527,N_1815);
or U2363 (N_2363,N_1500,N_1541);
nor U2364 (N_2364,N_1691,N_1952);
nor U2365 (N_2365,N_2041,N_2005);
nand U2366 (N_2366,N_1696,N_1614);
or U2367 (N_2367,N_1649,N_1940);
nand U2368 (N_2368,N_2194,N_1662);
and U2369 (N_2369,N_2131,N_2242);
xor U2370 (N_2370,N_1642,N_2137);
nand U2371 (N_2371,N_1530,N_1988);
nand U2372 (N_2372,N_1755,N_1700);
nand U2373 (N_2373,N_1787,N_1860);
or U2374 (N_2374,N_1561,N_2043);
or U2375 (N_2375,N_1908,N_1752);
nor U2376 (N_2376,N_1832,N_1816);
nand U2377 (N_2377,N_1563,N_2191);
or U2378 (N_2378,N_2246,N_2129);
or U2379 (N_2379,N_1637,N_2149);
and U2380 (N_2380,N_1852,N_1660);
xnor U2381 (N_2381,N_2152,N_1581);
nor U2382 (N_2382,N_1680,N_1673);
xor U2383 (N_2383,N_1636,N_1905);
nand U2384 (N_2384,N_1933,N_1930);
or U2385 (N_2385,N_2185,N_1566);
or U2386 (N_2386,N_2120,N_1871);
or U2387 (N_2387,N_2133,N_1513);
nand U2388 (N_2388,N_1508,N_1604);
xor U2389 (N_2389,N_2228,N_1738);
xor U2390 (N_2390,N_1879,N_2032);
nor U2391 (N_2391,N_2070,N_1830);
xor U2392 (N_2392,N_1742,N_2056);
xor U2393 (N_2393,N_1677,N_1797);
or U2394 (N_2394,N_1514,N_1503);
nor U2395 (N_2395,N_2241,N_2142);
xnor U2396 (N_2396,N_2226,N_2064);
nand U2397 (N_2397,N_1740,N_1964);
and U2398 (N_2398,N_1985,N_1953);
and U2399 (N_2399,N_1714,N_1795);
or U2400 (N_2400,N_1945,N_2011);
nor U2401 (N_2401,N_1593,N_1931);
nand U2402 (N_2402,N_1613,N_2012);
or U2403 (N_2403,N_2161,N_1814);
xnor U2404 (N_2404,N_1518,N_1828);
and U2405 (N_2405,N_2197,N_1615);
or U2406 (N_2406,N_1657,N_1655);
nor U2407 (N_2407,N_1690,N_1969);
nor U2408 (N_2408,N_1929,N_1923);
nor U2409 (N_2409,N_1720,N_1768);
nand U2410 (N_2410,N_1914,N_2092);
nand U2411 (N_2411,N_2097,N_2227);
xnor U2412 (N_2412,N_2109,N_2218);
or U2413 (N_2413,N_2082,N_1751);
xor U2414 (N_2414,N_1767,N_2049);
nor U2415 (N_2415,N_2123,N_1902);
or U2416 (N_2416,N_1997,N_1936);
nor U2417 (N_2417,N_1724,N_1962);
and U2418 (N_2418,N_1822,N_1824);
nor U2419 (N_2419,N_2046,N_1595);
or U2420 (N_2420,N_1736,N_2163);
nor U2421 (N_2421,N_2025,N_2139);
or U2422 (N_2422,N_1974,N_1521);
nand U2423 (N_2423,N_1550,N_1653);
or U2424 (N_2424,N_1507,N_1620);
nor U2425 (N_2425,N_1570,N_1540);
nor U2426 (N_2426,N_1783,N_2215);
nor U2427 (N_2427,N_1511,N_2108);
or U2428 (N_2428,N_2211,N_1715);
nor U2429 (N_2429,N_2209,N_1670);
xor U2430 (N_2430,N_1831,N_2069);
xor U2431 (N_2431,N_1866,N_1804);
nand U2432 (N_2432,N_1644,N_1624);
xnor U2433 (N_2433,N_1897,N_1834);
or U2434 (N_2434,N_1667,N_1539);
nand U2435 (N_2435,N_1520,N_1635);
nor U2436 (N_2436,N_1666,N_1509);
nand U2437 (N_2437,N_1735,N_1528);
xor U2438 (N_2438,N_2042,N_1602);
nor U2439 (N_2439,N_2088,N_1888);
and U2440 (N_2440,N_1838,N_2216);
xnor U2441 (N_2441,N_2182,N_1853);
xor U2442 (N_2442,N_2223,N_1942);
nor U2443 (N_2443,N_1702,N_1898);
nor U2444 (N_2444,N_2240,N_1650);
nor U2445 (N_2445,N_2198,N_1565);
nor U2446 (N_2446,N_1889,N_1793);
and U2447 (N_2447,N_2062,N_1678);
and U2448 (N_2448,N_1723,N_1725);
and U2449 (N_2449,N_2063,N_2022);
xor U2450 (N_2450,N_2052,N_1661);
xor U2451 (N_2451,N_1800,N_1578);
and U2452 (N_2452,N_1991,N_1799);
nor U2453 (N_2453,N_2098,N_1771);
nor U2454 (N_2454,N_1859,N_2159);
or U2455 (N_2455,N_2200,N_2084);
and U2456 (N_2456,N_2141,N_1652);
nor U2457 (N_2457,N_1876,N_1654);
and U2458 (N_2458,N_1922,N_1938);
nand U2459 (N_2459,N_1634,N_1756);
and U2460 (N_2460,N_1676,N_1825);
nor U2461 (N_2461,N_2183,N_1746);
xor U2462 (N_2462,N_1989,N_2090);
or U2463 (N_2463,N_1733,N_1607);
and U2464 (N_2464,N_1829,N_2050);
and U2465 (N_2465,N_1618,N_1525);
nor U2466 (N_2466,N_1656,N_1711);
xnor U2467 (N_2467,N_2004,N_1845);
nand U2468 (N_2468,N_1609,N_2224);
nand U2469 (N_2469,N_2007,N_2019);
and U2470 (N_2470,N_1812,N_2171);
nor U2471 (N_2471,N_1728,N_2061);
nor U2472 (N_2472,N_2030,N_2221);
nor U2473 (N_2473,N_1729,N_2214);
nand U2474 (N_2474,N_1972,N_1826);
nand U2475 (N_2475,N_2047,N_1610);
nor U2476 (N_2476,N_1958,N_2060);
nand U2477 (N_2477,N_1805,N_1907);
xnor U2478 (N_2478,N_1687,N_2071);
xor U2479 (N_2479,N_1906,N_1526);
xnor U2480 (N_2480,N_1764,N_1992);
nand U2481 (N_2481,N_2076,N_1698);
nor U2482 (N_2482,N_1682,N_2144);
xnor U2483 (N_2483,N_1586,N_2100);
and U2484 (N_2484,N_2154,N_2245);
nor U2485 (N_2485,N_1748,N_1679);
nor U2486 (N_2486,N_2045,N_1926);
nand U2487 (N_2487,N_2013,N_2208);
nor U2488 (N_2488,N_2205,N_1809);
or U2489 (N_2489,N_1909,N_1619);
or U2490 (N_2490,N_1807,N_1532);
nand U2491 (N_2491,N_1782,N_1960);
nor U2492 (N_2492,N_2036,N_1937);
nor U2493 (N_2493,N_1821,N_2093);
nand U2494 (N_2494,N_2107,N_1546);
and U2495 (N_2495,N_1760,N_1697);
nand U2496 (N_2496,N_2105,N_1856);
nand U2497 (N_2497,N_1741,N_1713);
nand U2498 (N_2498,N_1622,N_2124);
xnor U2499 (N_2499,N_1684,N_1778);
nor U2500 (N_2500,N_2029,N_1719);
nor U2501 (N_2501,N_1591,N_1801);
nor U2502 (N_2502,N_1739,N_2247);
and U2503 (N_2503,N_1976,N_1516);
and U2504 (N_2504,N_1633,N_2066);
nand U2505 (N_2505,N_2174,N_1502);
or U2506 (N_2506,N_2099,N_1983);
xor U2507 (N_2507,N_2147,N_2014);
xor U2508 (N_2508,N_1813,N_2217);
or U2509 (N_2509,N_1919,N_2010);
or U2510 (N_2510,N_2034,N_1981);
xnor U2511 (N_2511,N_2086,N_1867);
and U2512 (N_2512,N_1632,N_1576);
xor U2513 (N_2513,N_2190,N_2087);
nor U2514 (N_2514,N_2170,N_1626);
and U2515 (N_2515,N_1794,N_1558);
and U2516 (N_2516,N_1996,N_2169);
nand U2517 (N_2517,N_1798,N_1868);
or U2518 (N_2518,N_2202,N_2065);
nor U2519 (N_2519,N_2181,N_1762);
or U2520 (N_2520,N_1668,N_1598);
nor U2521 (N_2521,N_2117,N_1863);
and U2522 (N_2522,N_2028,N_2039);
or U2523 (N_2523,N_1689,N_2126);
nand U2524 (N_2524,N_2027,N_2230);
xor U2525 (N_2525,N_1837,N_1555);
and U2526 (N_2526,N_2140,N_1994);
xnor U2527 (N_2527,N_1861,N_2165);
xor U2528 (N_2528,N_1671,N_2089);
or U2529 (N_2529,N_2196,N_1672);
and U2530 (N_2530,N_1883,N_1921);
nand U2531 (N_2531,N_2094,N_1918);
xnor U2532 (N_2532,N_1885,N_1791);
nand U2533 (N_2533,N_2053,N_2231);
nand U2534 (N_2534,N_1583,N_1776);
and U2535 (N_2535,N_2112,N_1865);
nand U2536 (N_2536,N_2068,N_2157);
nand U2537 (N_2537,N_2167,N_1750);
xnor U2538 (N_2538,N_1699,N_1758);
xnor U2539 (N_2539,N_2031,N_1900);
nand U2540 (N_2540,N_1716,N_2002);
nand U2541 (N_2541,N_1966,N_2236);
and U2542 (N_2542,N_1884,N_2237);
nand U2543 (N_2543,N_1792,N_1786);
nand U2544 (N_2544,N_2243,N_2072);
or U2545 (N_2545,N_1811,N_1955);
nand U2546 (N_2546,N_1887,N_1895);
xor U2547 (N_2547,N_1537,N_2206);
nand U2548 (N_2548,N_1999,N_1545);
or U2549 (N_2549,N_1855,N_1934);
or U2550 (N_2550,N_2009,N_1935);
nand U2551 (N_2551,N_1524,N_2178);
nor U2552 (N_2552,N_1858,N_1878);
nand U2553 (N_2553,N_2127,N_1533);
nor U2554 (N_2554,N_2138,N_1747);
or U2555 (N_2555,N_1522,N_1873);
and U2556 (N_2556,N_2080,N_1877);
nand U2557 (N_2557,N_1968,N_2006);
or U2558 (N_2558,N_1986,N_1777);
nor U2559 (N_2559,N_1544,N_2128);
or U2560 (N_2560,N_1759,N_1820);
nor U2561 (N_2561,N_1568,N_2116);
nor U2562 (N_2562,N_1627,N_1803);
xnor U2563 (N_2563,N_2118,N_2125);
or U2564 (N_2564,N_1506,N_2119);
and U2565 (N_2565,N_1639,N_1841);
and U2566 (N_2566,N_1628,N_1582);
nand U2567 (N_2567,N_1630,N_1665);
xor U2568 (N_2568,N_2210,N_1818);
and U2569 (N_2569,N_1774,N_1727);
nor U2570 (N_2570,N_1788,N_1835);
nand U2571 (N_2571,N_2054,N_1836);
nand U2572 (N_2572,N_1848,N_2048);
or U2573 (N_2573,N_2180,N_2136);
nand U2574 (N_2574,N_1534,N_1536);
nor U2575 (N_2575,N_1784,N_2085);
xnor U2576 (N_2576,N_1910,N_1519);
nand U2577 (N_2577,N_1901,N_1874);
xor U2578 (N_2578,N_1913,N_1753);
nor U2579 (N_2579,N_1743,N_2081);
and U2580 (N_2580,N_1850,N_1535);
or U2581 (N_2581,N_2079,N_1819);
nand U2582 (N_2582,N_1731,N_2146);
xnor U2583 (N_2583,N_2114,N_1745);
and U2584 (N_2584,N_1882,N_2189);
or U2585 (N_2585,N_1990,N_1849);
and U2586 (N_2586,N_1854,N_1911);
nor U2587 (N_2587,N_1701,N_1686);
and U2588 (N_2588,N_2164,N_2096);
and U2589 (N_2589,N_1790,N_2172);
and U2590 (N_2590,N_1571,N_2207);
nor U2591 (N_2591,N_1875,N_2176);
and U2592 (N_2592,N_1548,N_1640);
and U2593 (N_2593,N_1894,N_1959);
nor U2594 (N_2594,N_1611,N_1695);
xnor U2595 (N_2595,N_2044,N_1681);
nor U2596 (N_2596,N_1567,N_2203);
and U2597 (N_2597,N_2110,N_1612);
nand U2598 (N_2598,N_1587,N_1995);
and U2599 (N_2599,N_1708,N_1643);
nor U2600 (N_2600,N_1543,N_1948);
nor U2601 (N_2601,N_1560,N_1949);
nor U2602 (N_2602,N_1600,N_1556);
or U2603 (N_2603,N_1862,N_2213);
or U2604 (N_2604,N_1903,N_2179);
or U2605 (N_2605,N_2148,N_1512);
nand U2606 (N_2606,N_2184,N_1647);
and U2607 (N_2607,N_1599,N_1779);
xnor U2608 (N_2608,N_2040,N_1857);
xor U2609 (N_2609,N_1601,N_1734);
xor U2610 (N_2610,N_2186,N_2222);
and U2611 (N_2611,N_1549,N_2104);
and U2612 (N_2612,N_1717,N_1590);
nand U2613 (N_2613,N_2038,N_1943);
nand U2614 (N_2614,N_1646,N_2166);
nor U2615 (N_2615,N_2238,N_1574);
nor U2616 (N_2616,N_1651,N_1947);
xnor U2617 (N_2617,N_1806,N_1722);
and U2618 (N_2618,N_1575,N_1761);
or U2619 (N_2619,N_2248,N_1658);
nor U2620 (N_2620,N_1869,N_1967);
nor U2621 (N_2621,N_2051,N_1954);
xnor U2622 (N_2622,N_2249,N_2077);
nor U2623 (N_2623,N_2229,N_1833);
nand U2624 (N_2624,N_1577,N_1810);
nor U2625 (N_2625,N_1671,N_2146);
nand U2626 (N_2626,N_2062,N_1775);
nor U2627 (N_2627,N_2169,N_1717);
nor U2628 (N_2628,N_1537,N_1801);
xnor U2629 (N_2629,N_1732,N_1788);
nor U2630 (N_2630,N_1536,N_1592);
nand U2631 (N_2631,N_1524,N_2038);
or U2632 (N_2632,N_1779,N_1653);
nor U2633 (N_2633,N_2020,N_1591);
or U2634 (N_2634,N_2234,N_1658);
xnor U2635 (N_2635,N_1839,N_1638);
nor U2636 (N_2636,N_1707,N_2084);
nand U2637 (N_2637,N_2213,N_1512);
or U2638 (N_2638,N_1700,N_1709);
xor U2639 (N_2639,N_2171,N_1638);
and U2640 (N_2640,N_2079,N_2022);
xor U2641 (N_2641,N_1904,N_2067);
nor U2642 (N_2642,N_2053,N_1547);
or U2643 (N_2643,N_1627,N_1558);
nor U2644 (N_2644,N_1765,N_1896);
xor U2645 (N_2645,N_1635,N_1572);
nor U2646 (N_2646,N_2190,N_1522);
or U2647 (N_2647,N_2065,N_1642);
or U2648 (N_2648,N_1639,N_2058);
xnor U2649 (N_2649,N_1972,N_2151);
nor U2650 (N_2650,N_1773,N_2177);
or U2651 (N_2651,N_1885,N_1731);
or U2652 (N_2652,N_1713,N_2246);
and U2653 (N_2653,N_1780,N_1553);
nor U2654 (N_2654,N_1827,N_1507);
nor U2655 (N_2655,N_2150,N_1609);
nor U2656 (N_2656,N_2073,N_1937);
nand U2657 (N_2657,N_2003,N_2187);
nand U2658 (N_2658,N_1509,N_2019);
xor U2659 (N_2659,N_1731,N_2231);
xor U2660 (N_2660,N_2176,N_1535);
nand U2661 (N_2661,N_1963,N_2193);
nor U2662 (N_2662,N_1848,N_1979);
nand U2663 (N_2663,N_1706,N_2059);
or U2664 (N_2664,N_1557,N_2096);
or U2665 (N_2665,N_2135,N_2066);
nand U2666 (N_2666,N_2132,N_1871);
xor U2667 (N_2667,N_1548,N_2114);
and U2668 (N_2668,N_2221,N_1973);
xor U2669 (N_2669,N_1839,N_1515);
xor U2670 (N_2670,N_1617,N_2156);
nand U2671 (N_2671,N_1656,N_1723);
xor U2672 (N_2672,N_1773,N_2167);
nand U2673 (N_2673,N_1548,N_1729);
and U2674 (N_2674,N_1620,N_2053);
nand U2675 (N_2675,N_1672,N_2038);
nand U2676 (N_2676,N_1699,N_1887);
nor U2677 (N_2677,N_2221,N_1630);
xor U2678 (N_2678,N_1586,N_1661);
or U2679 (N_2679,N_2079,N_1665);
xor U2680 (N_2680,N_1742,N_1748);
and U2681 (N_2681,N_1704,N_1547);
or U2682 (N_2682,N_1980,N_1624);
nor U2683 (N_2683,N_1889,N_1959);
xnor U2684 (N_2684,N_1612,N_1855);
and U2685 (N_2685,N_2191,N_1785);
and U2686 (N_2686,N_2089,N_2147);
nor U2687 (N_2687,N_1705,N_2219);
and U2688 (N_2688,N_1507,N_1524);
or U2689 (N_2689,N_1794,N_1819);
nand U2690 (N_2690,N_1670,N_1879);
or U2691 (N_2691,N_2139,N_2023);
xor U2692 (N_2692,N_2156,N_1837);
and U2693 (N_2693,N_2064,N_1897);
nor U2694 (N_2694,N_1912,N_1509);
or U2695 (N_2695,N_1730,N_2209);
nor U2696 (N_2696,N_1761,N_1865);
nor U2697 (N_2697,N_1702,N_1669);
or U2698 (N_2698,N_2095,N_1548);
xor U2699 (N_2699,N_2092,N_1649);
xnor U2700 (N_2700,N_2038,N_1725);
nor U2701 (N_2701,N_1651,N_1916);
or U2702 (N_2702,N_1871,N_2152);
nand U2703 (N_2703,N_1891,N_2180);
nor U2704 (N_2704,N_1898,N_1523);
nand U2705 (N_2705,N_1735,N_1679);
nor U2706 (N_2706,N_2188,N_1784);
and U2707 (N_2707,N_1500,N_1972);
xnor U2708 (N_2708,N_2116,N_1613);
xor U2709 (N_2709,N_1546,N_2188);
and U2710 (N_2710,N_2177,N_1963);
nand U2711 (N_2711,N_1926,N_2017);
xnor U2712 (N_2712,N_1695,N_2139);
nor U2713 (N_2713,N_1766,N_1648);
nor U2714 (N_2714,N_2121,N_1934);
or U2715 (N_2715,N_2055,N_1903);
nand U2716 (N_2716,N_1571,N_1815);
nor U2717 (N_2717,N_1515,N_1895);
or U2718 (N_2718,N_1694,N_1561);
nor U2719 (N_2719,N_1981,N_1769);
nor U2720 (N_2720,N_1966,N_2201);
nor U2721 (N_2721,N_2049,N_1945);
nor U2722 (N_2722,N_2170,N_1528);
nand U2723 (N_2723,N_2060,N_1742);
or U2724 (N_2724,N_1937,N_2166);
nor U2725 (N_2725,N_2140,N_1572);
or U2726 (N_2726,N_2222,N_1976);
or U2727 (N_2727,N_1814,N_1971);
and U2728 (N_2728,N_1920,N_1522);
or U2729 (N_2729,N_2070,N_1926);
or U2730 (N_2730,N_2014,N_2067);
xor U2731 (N_2731,N_1512,N_1993);
nor U2732 (N_2732,N_2228,N_1995);
nand U2733 (N_2733,N_1700,N_1522);
nor U2734 (N_2734,N_1558,N_1772);
nor U2735 (N_2735,N_2064,N_1894);
nor U2736 (N_2736,N_1655,N_2022);
nand U2737 (N_2737,N_2173,N_1707);
nand U2738 (N_2738,N_2067,N_1712);
nor U2739 (N_2739,N_2144,N_2141);
nand U2740 (N_2740,N_1668,N_1684);
xor U2741 (N_2741,N_1567,N_1600);
and U2742 (N_2742,N_1961,N_1505);
nand U2743 (N_2743,N_1992,N_1927);
xor U2744 (N_2744,N_2235,N_1881);
nor U2745 (N_2745,N_1519,N_1903);
or U2746 (N_2746,N_1557,N_2147);
and U2747 (N_2747,N_1509,N_1880);
xnor U2748 (N_2748,N_2203,N_1600);
nor U2749 (N_2749,N_2064,N_1835);
and U2750 (N_2750,N_1646,N_1962);
nor U2751 (N_2751,N_1535,N_1817);
or U2752 (N_2752,N_1671,N_1659);
nor U2753 (N_2753,N_1562,N_1953);
nor U2754 (N_2754,N_2040,N_1940);
xnor U2755 (N_2755,N_1829,N_1976);
or U2756 (N_2756,N_2165,N_1766);
nand U2757 (N_2757,N_2166,N_1899);
nor U2758 (N_2758,N_1539,N_2023);
and U2759 (N_2759,N_1993,N_2204);
xnor U2760 (N_2760,N_1863,N_2134);
nor U2761 (N_2761,N_2065,N_1903);
nand U2762 (N_2762,N_1994,N_1975);
and U2763 (N_2763,N_1517,N_1767);
or U2764 (N_2764,N_1603,N_2052);
xor U2765 (N_2765,N_2180,N_1904);
nand U2766 (N_2766,N_2052,N_1956);
xor U2767 (N_2767,N_1815,N_1944);
nand U2768 (N_2768,N_1804,N_2016);
and U2769 (N_2769,N_2236,N_1542);
nand U2770 (N_2770,N_2040,N_1643);
xnor U2771 (N_2771,N_1897,N_1682);
nand U2772 (N_2772,N_2228,N_1721);
nor U2773 (N_2773,N_1647,N_2072);
nor U2774 (N_2774,N_1501,N_1778);
or U2775 (N_2775,N_1561,N_1991);
or U2776 (N_2776,N_1897,N_1602);
nor U2777 (N_2777,N_1896,N_1550);
and U2778 (N_2778,N_1932,N_1764);
or U2779 (N_2779,N_1890,N_1553);
and U2780 (N_2780,N_2158,N_1802);
nand U2781 (N_2781,N_1907,N_1639);
and U2782 (N_2782,N_2097,N_2162);
xnor U2783 (N_2783,N_1951,N_2134);
nor U2784 (N_2784,N_2114,N_2083);
nand U2785 (N_2785,N_2019,N_1572);
xor U2786 (N_2786,N_1855,N_2218);
nand U2787 (N_2787,N_1868,N_1959);
nand U2788 (N_2788,N_1740,N_1750);
or U2789 (N_2789,N_1609,N_2242);
nor U2790 (N_2790,N_1624,N_1684);
and U2791 (N_2791,N_2236,N_2011);
or U2792 (N_2792,N_2152,N_2078);
nor U2793 (N_2793,N_2239,N_2133);
nand U2794 (N_2794,N_1722,N_1974);
and U2795 (N_2795,N_2169,N_1827);
nand U2796 (N_2796,N_1684,N_1860);
xor U2797 (N_2797,N_2086,N_2050);
xor U2798 (N_2798,N_1917,N_1895);
and U2799 (N_2799,N_2157,N_2007);
nand U2800 (N_2800,N_2141,N_2119);
nor U2801 (N_2801,N_1644,N_2015);
xor U2802 (N_2802,N_2106,N_2154);
or U2803 (N_2803,N_1986,N_1845);
nand U2804 (N_2804,N_1708,N_1896);
and U2805 (N_2805,N_2018,N_1688);
or U2806 (N_2806,N_1669,N_1572);
and U2807 (N_2807,N_1728,N_1639);
or U2808 (N_2808,N_1575,N_2079);
and U2809 (N_2809,N_1866,N_1977);
nor U2810 (N_2810,N_1798,N_1836);
xor U2811 (N_2811,N_1624,N_1786);
nand U2812 (N_2812,N_1518,N_2000);
nand U2813 (N_2813,N_1635,N_1805);
nand U2814 (N_2814,N_1518,N_1956);
and U2815 (N_2815,N_2124,N_1550);
nand U2816 (N_2816,N_1780,N_1707);
and U2817 (N_2817,N_1670,N_1808);
and U2818 (N_2818,N_1562,N_1613);
xnor U2819 (N_2819,N_1557,N_1579);
nand U2820 (N_2820,N_1871,N_1888);
xnor U2821 (N_2821,N_2128,N_1680);
xnor U2822 (N_2822,N_1830,N_2172);
nor U2823 (N_2823,N_1537,N_1999);
and U2824 (N_2824,N_1848,N_1711);
and U2825 (N_2825,N_1648,N_1688);
nor U2826 (N_2826,N_2199,N_2218);
xnor U2827 (N_2827,N_2102,N_2193);
or U2828 (N_2828,N_2220,N_2173);
nor U2829 (N_2829,N_1902,N_1576);
or U2830 (N_2830,N_2101,N_1906);
nand U2831 (N_2831,N_2069,N_1765);
nand U2832 (N_2832,N_1571,N_1511);
nand U2833 (N_2833,N_2191,N_1872);
and U2834 (N_2834,N_1784,N_1665);
nand U2835 (N_2835,N_2014,N_2164);
nor U2836 (N_2836,N_1769,N_2006);
xor U2837 (N_2837,N_2023,N_2225);
nand U2838 (N_2838,N_2024,N_2181);
nor U2839 (N_2839,N_1958,N_1643);
and U2840 (N_2840,N_1540,N_2172);
or U2841 (N_2841,N_2029,N_1507);
and U2842 (N_2842,N_2068,N_2052);
xor U2843 (N_2843,N_1749,N_1764);
and U2844 (N_2844,N_1630,N_1598);
or U2845 (N_2845,N_2093,N_2051);
nor U2846 (N_2846,N_1639,N_1597);
nand U2847 (N_2847,N_1657,N_2036);
or U2848 (N_2848,N_1616,N_1936);
nor U2849 (N_2849,N_1510,N_1888);
or U2850 (N_2850,N_1766,N_2239);
and U2851 (N_2851,N_1645,N_1926);
xnor U2852 (N_2852,N_1767,N_1733);
nand U2853 (N_2853,N_2203,N_2061);
xnor U2854 (N_2854,N_2047,N_1521);
and U2855 (N_2855,N_2103,N_1512);
and U2856 (N_2856,N_1807,N_1773);
nor U2857 (N_2857,N_2172,N_1959);
nand U2858 (N_2858,N_1955,N_1967);
nand U2859 (N_2859,N_2039,N_1539);
nand U2860 (N_2860,N_1811,N_1934);
or U2861 (N_2861,N_2037,N_2029);
xnor U2862 (N_2862,N_1603,N_1677);
or U2863 (N_2863,N_2100,N_2074);
nand U2864 (N_2864,N_1508,N_1989);
nand U2865 (N_2865,N_2006,N_1750);
xor U2866 (N_2866,N_1865,N_2218);
or U2867 (N_2867,N_2049,N_1891);
nand U2868 (N_2868,N_1618,N_2127);
or U2869 (N_2869,N_1531,N_1586);
nor U2870 (N_2870,N_1697,N_2190);
nand U2871 (N_2871,N_1747,N_1734);
and U2872 (N_2872,N_2082,N_1765);
or U2873 (N_2873,N_2157,N_2190);
xor U2874 (N_2874,N_1599,N_1879);
nor U2875 (N_2875,N_1607,N_2229);
and U2876 (N_2876,N_2169,N_1651);
nand U2877 (N_2877,N_1597,N_1688);
xnor U2878 (N_2878,N_1546,N_2068);
xor U2879 (N_2879,N_1670,N_1909);
xor U2880 (N_2880,N_1688,N_2088);
and U2881 (N_2881,N_2224,N_2248);
nor U2882 (N_2882,N_1817,N_2046);
nand U2883 (N_2883,N_1581,N_2021);
or U2884 (N_2884,N_1596,N_1720);
or U2885 (N_2885,N_1970,N_1957);
and U2886 (N_2886,N_2001,N_1617);
or U2887 (N_2887,N_1831,N_1979);
nor U2888 (N_2888,N_1564,N_1582);
nor U2889 (N_2889,N_2030,N_1509);
and U2890 (N_2890,N_1880,N_1862);
or U2891 (N_2891,N_1976,N_2104);
or U2892 (N_2892,N_1599,N_1826);
xor U2893 (N_2893,N_2229,N_1544);
nand U2894 (N_2894,N_2033,N_1774);
xor U2895 (N_2895,N_1989,N_1770);
xnor U2896 (N_2896,N_2187,N_1913);
nand U2897 (N_2897,N_1722,N_1810);
nor U2898 (N_2898,N_1670,N_1689);
and U2899 (N_2899,N_1609,N_2135);
xnor U2900 (N_2900,N_1761,N_1691);
and U2901 (N_2901,N_1748,N_1572);
and U2902 (N_2902,N_1517,N_1929);
nand U2903 (N_2903,N_2230,N_1904);
xor U2904 (N_2904,N_1848,N_2093);
nand U2905 (N_2905,N_1650,N_1731);
or U2906 (N_2906,N_1939,N_1875);
and U2907 (N_2907,N_2092,N_1582);
xor U2908 (N_2908,N_1678,N_1956);
nand U2909 (N_2909,N_1933,N_2174);
nand U2910 (N_2910,N_2217,N_2105);
xor U2911 (N_2911,N_1527,N_2080);
nor U2912 (N_2912,N_2076,N_1884);
xnor U2913 (N_2913,N_1528,N_2008);
nor U2914 (N_2914,N_1679,N_1523);
xnor U2915 (N_2915,N_1775,N_1840);
nor U2916 (N_2916,N_1993,N_1918);
and U2917 (N_2917,N_1951,N_2013);
and U2918 (N_2918,N_2164,N_2167);
or U2919 (N_2919,N_1656,N_1706);
and U2920 (N_2920,N_1723,N_1557);
nor U2921 (N_2921,N_1521,N_2040);
xor U2922 (N_2922,N_1763,N_1539);
xor U2923 (N_2923,N_1919,N_2082);
xnor U2924 (N_2924,N_1903,N_1673);
nand U2925 (N_2925,N_1652,N_1559);
xor U2926 (N_2926,N_2012,N_1618);
xnor U2927 (N_2927,N_1943,N_1756);
or U2928 (N_2928,N_1537,N_1577);
and U2929 (N_2929,N_2169,N_1674);
or U2930 (N_2930,N_1956,N_1750);
xnor U2931 (N_2931,N_1544,N_2192);
nand U2932 (N_2932,N_1873,N_1763);
xor U2933 (N_2933,N_1520,N_1550);
nor U2934 (N_2934,N_2051,N_1808);
nand U2935 (N_2935,N_1710,N_1926);
nor U2936 (N_2936,N_1618,N_1818);
or U2937 (N_2937,N_2022,N_1648);
or U2938 (N_2938,N_2079,N_2090);
or U2939 (N_2939,N_1914,N_1951);
and U2940 (N_2940,N_1781,N_1633);
nor U2941 (N_2941,N_1636,N_2139);
or U2942 (N_2942,N_1519,N_1960);
nand U2943 (N_2943,N_1929,N_2105);
or U2944 (N_2944,N_1508,N_2138);
xor U2945 (N_2945,N_2046,N_1869);
nand U2946 (N_2946,N_1513,N_2165);
nand U2947 (N_2947,N_1678,N_1505);
xor U2948 (N_2948,N_2127,N_2046);
and U2949 (N_2949,N_1613,N_1716);
or U2950 (N_2950,N_1697,N_1749);
xnor U2951 (N_2951,N_2023,N_1867);
xnor U2952 (N_2952,N_2134,N_1606);
nand U2953 (N_2953,N_2120,N_1600);
and U2954 (N_2954,N_1727,N_1972);
and U2955 (N_2955,N_1600,N_1644);
nand U2956 (N_2956,N_1562,N_1807);
or U2957 (N_2957,N_1575,N_1650);
nand U2958 (N_2958,N_1574,N_2041);
nor U2959 (N_2959,N_1791,N_2214);
xnor U2960 (N_2960,N_2014,N_1811);
or U2961 (N_2961,N_2162,N_2062);
and U2962 (N_2962,N_1973,N_1685);
nand U2963 (N_2963,N_2246,N_2235);
nor U2964 (N_2964,N_2213,N_1899);
xnor U2965 (N_2965,N_1695,N_2217);
nor U2966 (N_2966,N_2190,N_1541);
or U2967 (N_2967,N_1758,N_1842);
and U2968 (N_2968,N_1876,N_2150);
xor U2969 (N_2969,N_1844,N_2048);
or U2970 (N_2970,N_1579,N_1869);
nor U2971 (N_2971,N_1913,N_2005);
nor U2972 (N_2972,N_1749,N_1973);
xor U2973 (N_2973,N_2021,N_2211);
and U2974 (N_2974,N_1586,N_1523);
nor U2975 (N_2975,N_1905,N_1943);
nor U2976 (N_2976,N_1566,N_1692);
xnor U2977 (N_2977,N_2058,N_1828);
nand U2978 (N_2978,N_2206,N_1738);
xor U2979 (N_2979,N_2247,N_1720);
or U2980 (N_2980,N_2198,N_1808);
nor U2981 (N_2981,N_1542,N_2179);
nand U2982 (N_2982,N_2214,N_2134);
and U2983 (N_2983,N_2111,N_1868);
xnor U2984 (N_2984,N_2034,N_2142);
nor U2985 (N_2985,N_1560,N_1691);
xor U2986 (N_2986,N_1983,N_2222);
nand U2987 (N_2987,N_2141,N_1994);
xor U2988 (N_2988,N_1733,N_2133);
nor U2989 (N_2989,N_1620,N_2077);
or U2990 (N_2990,N_1659,N_1608);
nor U2991 (N_2991,N_2061,N_1534);
or U2992 (N_2992,N_1727,N_1931);
nand U2993 (N_2993,N_1823,N_1608);
nand U2994 (N_2994,N_2225,N_1572);
or U2995 (N_2995,N_1629,N_1521);
nor U2996 (N_2996,N_2091,N_2018);
or U2997 (N_2997,N_2232,N_1566);
and U2998 (N_2998,N_1855,N_1768);
and U2999 (N_2999,N_2225,N_1686);
and UO_0 (O_0,N_2330,N_2952);
nand UO_1 (O_1,N_2707,N_2462);
nand UO_2 (O_2,N_2653,N_2279);
or UO_3 (O_3,N_2399,N_2484);
and UO_4 (O_4,N_2455,N_2449);
or UO_5 (O_5,N_2986,N_2789);
nor UO_6 (O_6,N_2460,N_2508);
or UO_7 (O_7,N_2562,N_2610);
and UO_8 (O_8,N_2721,N_2271);
nand UO_9 (O_9,N_2407,N_2543);
nand UO_10 (O_10,N_2253,N_2301);
nor UO_11 (O_11,N_2328,N_2684);
and UO_12 (O_12,N_2414,N_2617);
xor UO_13 (O_13,N_2589,N_2490);
and UO_14 (O_14,N_2578,N_2257);
nand UO_15 (O_15,N_2528,N_2926);
nand UO_16 (O_16,N_2337,N_2322);
xnor UO_17 (O_17,N_2637,N_2560);
nand UO_18 (O_18,N_2519,N_2379);
and UO_19 (O_19,N_2964,N_2458);
or UO_20 (O_20,N_2318,N_2896);
and UO_21 (O_21,N_2385,N_2402);
and UO_22 (O_22,N_2607,N_2970);
nor UO_23 (O_23,N_2639,N_2456);
or UO_24 (O_24,N_2930,N_2281);
xor UO_25 (O_25,N_2856,N_2259);
xor UO_26 (O_26,N_2640,N_2715);
and UO_27 (O_27,N_2650,N_2877);
nor UO_28 (O_28,N_2906,N_2737);
or UO_29 (O_29,N_2424,N_2536);
and UO_30 (O_30,N_2558,N_2552);
nand UO_31 (O_31,N_2500,N_2944);
or UO_32 (O_32,N_2924,N_2418);
and UO_33 (O_33,N_2838,N_2442);
or UO_34 (O_34,N_2570,N_2932);
or UO_35 (O_35,N_2574,N_2692);
or UO_36 (O_36,N_2312,N_2450);
nor UO_37 (O_37,N_2674,N_2808);
xor UO_38 (O_38,N_2995,N_2400);
or UO_39 (O_39,N_2818,N_2396);
or UO_40 (O_40,N_2710,N_2306);
nand UO_41 (O_41,N_2783,N_2367);
nand UO_42 (O_42,N_2439,N_2940);
xor UO_43 (O_43,N_2358,N_2515);
xor UO_44 (O_44,N_2530,N_2647);
nand UO_45 (O_45,N_2605,N_2485);
nor UO_46 (O_46,N_2767,N_2738);
or UO_47 (O_47,N_2711,N_2912);
xor UO_48 (O_48,N_2889,N_2649);
xnor UO_49 (O_49,N_2459,N_2324);
and UO_50 (O_50,N_2730,N_2611);
xor UO_51 (O_51,N_2966,N_2894);
or UO_52 (O_52,N_2983,N_2817);
and UO_53 (O_53,N_2935,N_2825);
nand UO_54 (O_54,N_2526,N_2822);
xor UO_55 (O_55,N_2495,N_2916);
nor UO_56 (O_56,N_2993,N_2643);
nor UO_57 (O_57,N_2941,N_2507);
and UO_58 (O_58,N_2440,N_2394);
and UO_59 (O_59,N_2572,N_2869);
and UO_60 (O_60,N_2800,N_2561);
nor UO_61 (O_61,N_2901,N_2364);
xor UO_62 (O_62,N_2996,N_2777);
nand UO_63 (O_63,N_2757,N_2290);
nand UO_64 (O_64,N_2489,N_2447);
or UO_65 (O_65,N_2261,N_2727);
nand UO_66 (O_66,N_2582,N_2579);
nor UO_67 (O_67,N_2759,N_2251);
nor UO_68 (O_68,N_2585,N_2307);
xnor UO_69 (O_69,N_2383,N_2457);
xor UO_70 (O_70,N_2753,N_2881);
nor UO_71 (O_71,N_2850,N_2310);
xor UO_72 (O_72,N_2883,N_2331);
and UO_73 (O_73,N_2412,N_2566);
xor UO_74 (O_74,N_2670,N_2915);
nor UO_75 (O_75,N_2422,N_2875);
nor UO_76 (O_76,N_2360,N_2491);
nand UO_77 (O_77,N_2280,N_2660);
xor UO_78 (O_78,N_2776,N_2648);
nor UO_79 (O_79,N_2565,N_2588);
or UO_80 (O_80,N_2946,N_2876);
nand UO_81 (O_81,N_2775,N_2746);
or UO_82 (O_82,N_2339,N_2819);
or UO_83 (O_83,N_2343,N_2833);
nand UO_84 (O_84,N_2854,N_2813);
or UO_85 (O_85,N_2677,N_2867);
and UO_86 (O_86,N_2398,N_2803);
and UO_87 (O_87,N_2874,N_2262);
nor UO_88 (O_88,N_2269,N_2370);
nand UO_89 (O_89,N_2614,N_2812);
nor UO_90 (O_90,N_2722,N_2428);
nand UO_91 (O_91,N_2750,N_2371);
xor UO_92 (O_92,N_2796,N_2778);
xor UO_93 (O_93,N_2569,N_2992);
xor UO_94 (O_94,N_2619,N_2938);
xnor UO_95 (O_95,N_2401,N_2288);
xor UO_96 (O_96,N_2705,N_2918);
nand UO_97 (O_97,N_2387,N_2942);
nand UO_98 (O_98,N_2657,N_2327);
nand UO_99 (O_99,N_2836,N_2268);
xor UO_100 (O_100,N_2904,N_2583);
and UO_101 (O_101,N_2505,N_2443);
xor UO_102 (O_102,N_2701,N_2673);
or UO_103 (O_103,N_2446,N_2735);
and UO_104 (O_104,N_2863,N_2454);
xnor UO_105 (O_105,N_2474,N_2999);
xor UO_106 (O_106,N_2294,N_2700);
nand UO_107 (O_107,N_2763,N_2523);
nor UO_108 (O_108,N_2356,N_2962);
nor UO_109 (O_109,N_2405,N_2470);
xor UO_110 (O_110,N_2511,N_2628);
or UO_111 (O_111,N_2250,N_2359);
nand UO_112 (O_112,N_2499,N_2537);
nor UO_113 (O_113,N_2603,N_2622);
or UO_114 (O_114,N_2873,N_2732);
or UO_115 (O_115,N_2802,N_2580);
nand UO_116 (O_116,N_2917,N_2656);
and UO_117 (O_117,N_2606,N_2682);
or UO_118 (O_118,N_2512,N_2974);
nand UO_119 (O_119,N_2849,N_2571);
xnor UO_120 (O_120,N_2404,N_2847);
nor UO_121 (O_121,N_2464,N_2529);
and UO_122 (O_122,N_2340,N_2954);
nor UO_123 (O_123,N_2806,N_2563);
nor UO_124 (O_124,N_2870,N_2544);
nor UO_125 (O_125,N_2934,N_2888);
and UO_126 (O_126,N_2551,N_2785);
and UO_127 (O_127,N_2299,N_2305);
nor UO_128 (O_128,N_2586,N_2821);
nor UO_129 (O_129,N_2958,N_2843);
xnor UO_130 (O_130,N_2754,N_2827);
and UO_131 (O_131,N_2975,N_2885);
nor UO_132 (O_132,N_2406,N_2680);
nand UO_133 (O_133,N_2898,N_2357);
nor UO_134 (O_134,N_2953,N_2300);
or UO_135 (O_135,N_2403,N_2316);
nor UO_136 (O_136,N_2909,N_2659);
nand UO_137 (O_137,N_2591,N_2273);
nand UO_138 (O_138,N_2745,N_2839);
or UO_139 (O_139,N_2483,N_2351);
or UO_140 (O_140,N_2646,N_2516);
xor UO_141 (O_141,N_2641,N_2304);
nand UO_142 (O_142,N_2937,N_2718);
and UO_143 (O_143,N_2807,N_2765);
or UO_144 (O_144,N_2998,N_2335);
nor UO_145 (O_145,N_2429,N_2264);
nor UO_146 (O_146,N_2286,N_2728);
or UO_147 (O_147,N_2960,N_2630);
nor UO_148 (O_148,N_2716,N_2609);
and UO_149 (O_149,N_2501,N_2432);
xor UO_150 (O_150,N_2602,N_2488);
and UO_151 (O_151,N_2797,N_2465);
xnor UO_152 (O_152,N_2830,N_2476);
nor UO_153 (O_153,N_2631,N_2948);
or UO_154 (O_154,N_2900,N_2895);
or UO_155 (O_155,N_2349,N_2726);
and UO_156 (O_156,N_2514,N_2842);
xor UO_157 (O_157,N_2671,N_2840);
nand UO_158 (O_158,N_2503,N_2920);
xor UO_159 (O_159,N_2548,N_2270);
or UO_160 (O_160,N_2595,N_2756);
xor UO_161 (O_161,N_2581,N_2309);
nand UO_162 (O_162,N_2604,N_2487);
nor UO_163 (O_163,N_2568,N_2252);
xor UO_164 (O_164,N_2687,N_2448);
and UO_165 (O_165,N_2265,N_2771);
and UO_166 (O_166,N_2620,N_2471);
and UO_167 (O_167,N_2793,N_2597);
nand UO_168 (O_168,N_2768,N_2892);
or UO_169 (O_169,N_2553,N_2633);
xnor UO_170 (O_170,N_2409,N_2729);
or UO_171 (O_171,N_2661,N_2770);
or UO_172 (O_172,N_2903,N_2890);
nor UO_173 (O_173,N_2764,N_2740);
or UO_174 (O_174,N_2751,N_2527);
nand UO_175 (O_175,N_2391,N_2734);
and UO_176 (O_176,N_2635,N_2593);
nand UO_177 (O_177,N_2928,N_2278);
xnor UO_178 (O_178,N_2472,N_2662);
xnor UO_179 (O_179,N_2366,N_2302);
and UO_180 (O_180,N_2596,N_2277);
nand UO_181 (O_181,N_2625,N_2323);
nand UO_182 (O_182,N_2627,N_2296);
and UO_183 (O_183,N_2547,N_2535);
and UO_184 (O_184,N_2598,N_2961);
and UO_185 (O_185,N_2678,N_2969);
nand UO_186 (O_186,N_2857,N_2858);
and UO_187 (O_187,N_2742,N_2355);
nand UO_188 (O_188,N_2760,N_2498);
and UO_189 (O_189,N_2263,N_2698);
nor UO_190 (O_190,N_2720,N_2434);
nand UO_191 (O_191,N_2976,N_2258);
nand UO_192 (O_192,N_2717,N_2697);
nor UO_193 (O_193,N_2688,N_2786);
nand UO_194 (O_194,N_2815,N_2467);
nand UO_195 (O_195,N_2666,N_2882);
nand UO_196 (O_196,N_2744,N_2291);
or UO_197 (O_197,N_2347,N_2636);
nor UO_198 (O_198,N_2590,N_2524);
xnor UO_199 (O_199,N_2539,N_2787);
or UO_200 (O_200,N_2390,N_2564);
and UO_201 (O_201,N_2397,N_2616);
nor UO_202 (O_202,N_2334,N_2749);
or UO_203 (O_203,N_2353,N_2654);
nand UO_204 (O_204,N_2779,N_2284);
nor UO_205 (O_205,N_2979,N_2899);
or UO_206 (O_206,N_2546,N_2438);
xor UO_207 (O_207,N_2599,N_2411);
or UO_208 (O_208,N_2860,N_2445);
or UO_209 (O_209,N_2274,N_2477);
or UO_210 (O_210,N_2923,N_2984);
xnor UO_211 (O_211,N_2987,N_2897);
nand UO_212 (O_212,N_2626,N_2315);
nand UO_213 (O_213,N_2731,N_2762);
xor UO_214 (O_214,N_2559,N_2834);
nand UO_215 (O_215,N_2473,N_2341);
nor UO_216 (O_216,N_2266,N_2844);
and UO_217 (O_217,N_2913,N_2982);
nor UO_218 (O_218,N_2865,N_2550);
and UO_219 (O_219,N_2420,N_2798);
and UO_220 (O_220,N_2837,N_2933);
or UO_221 (O_221,N_2621,N_2545);
or UO_222 (O_222,N_2283,N_2652);
and UO_223 (O_223,N_2408,N_2413);
or UO_224 (O_224,N_2880,N_2292);
and UO_225 (O_225,N_2493,N_2879);
or UO_226 (O_226,N_2425,N_2829);
or UO_227 (O_227,N_2748,N_2384);
xnor UO_228 (O_228,N_2267,N_2664);
or UO_229 (O_229,N_2855,N_2478);
nand UO_230 (O_230,N_2835,N_2575);
xor UO_231 (O_231,N_2902,N_2790);
nor UO_232 (O_232,N_2372,N_2708);
xnor UO_233 (O_233,N_2520,N_2828);
or UO_234 (O_234,N_2592,N_2336);
xor UO_235 (O_235,N_2668,N_2685);
nor UO_236 (O_236,N_2861,N_2809);
or UO_237 (O_237,N_2496,N_2376);
nor UO_238 (O_238,N_2321,N_2618);
nand UO_239 (O_239,N_2922,N_2971);
nor UO_240 (O_240,N_2441,N_2494);
and UO_241 (O_241,N_2612,N_2949);
or UO_242 (O_242,N_2461,N_2344);
nor UO_243 (O_243,N_2794,N_2363);
xor UO_244 (O_244,N_2816,N_2823);
nand UO_245 (O_245,N_2638,N_2696);
nand UO_246 (O_246,N_2451,N_2644);
and UO_247 (O_247,N_2276,N_2416);
nor UO_248 (O_248,N_2521,N_2846);
nor UO_249 (O_249,N_2377,N_2957);
nor UO_250 (O_250,N_2695,N_2361);
xnor UO_251 (O_251,N_2848,N_2739);
xnor UO_252 (O_252,N_2820,N_2921);
nor UO_253 (O_253,N_2393,N_2792);
xor UO_254 (O_254,N_2805,N_2629);
and UO_255 (O_255,N_2741,N_2725);
xor UO_256 (O_256,N_2706,N_2632);
nor UO_257 (O_257,N_2541,N_2985);
nor UO_258 (O_258,N_2887,N_2557);
and UO_259 (O_259,N_2772,N_2479);
and UO_260 (O_260,N_2513,N_2824);
or UO_261 (O_261,N_2338,N_2782);
nand UO_262 (O_262,N_2943,N_2486);
xnor UO_263 (O_263,N_2348,N_2781);
and UO_264 (O_264,N_2320,N_2905);
nor UO_265 (O_265,N_2645,N_2686);
or UO_266 (O_266,N_2799,N_2410);
nor UO_267 (O_267,N_2255,N_2502);
xor UO_268 (O_268,N_2430,N_2851);
xor UO_269 (O_269,N_2272,N_2852);
nor UO_270 (O_270,N_2368,N_2554);
xnor UO_271 (O_271,N_2421,N_2482);
xnor UO_272 (O_272,N_2965,N_2893);
nor UO_273 (O_273,N_2382,N_2814);
xor UO_274 (O_274,N_2973,N_2919);
and UO_275 (O_275,N_2676,N_2665);
or UO_276 (O_276,N_2466,N_2587);
and UO_277 (O_277,N_2667,N_2936);
or UO_278 (O_278,N_2791,N_2350);
and UO_279 (O_279,N_2378,N_2955);
or UO_280 (O_280,N_2801,N_2314);
nand UO_281 (O_281,N_2702,N_2532);
and UO_282 (O_282,N_2555,N_2872);
and UO_283 (O_283,N_2373,N_2931);
xor UO_284 (O_284,N_2287,N_2947);
nor UO_285 (O_285,N_2342,N_2910);
or UO_286 (O_286,N_2567,N_2504);
and UO_287 (O_287,N_2886,N_2573);
or UO_288 (O_288,N_2709,N_2285);
and UO_289 (O_289,N_2991,N_2594);
nand UO_290 (O_290,N_2699,N_2497);
nand UO_291 (O_291,N_2540,N_2988);
or UO_292 (O_292,N_2380,N_2981);
and UO_293 (O_293,N_2752,N_2615);
xor UO_294 (O_294,N_2841,N_2866);
nor UO_295 (O_295,N_2436,N_2968);
and UO_296 (O_296,N_2989,N_2282);
or UO_297 (O_297,N_2313,N_2788);
and UO_298 (O_298,N_2747,N_2375);
and UO_299 (O_299,N_2864,N_2452);
and UO_300 (O_300,N_2733,N_2345);
nand UO_301 (O_301,N_2419,N_2362);
or UO_302 (O_302,N_2533,N_2365);
or UO_303 (O_303,N_2386,N_2784);
and UO_304 (O_304,N_2859,N_2769);
or UO_305 (O_305,N_2469,N_2427);
and UO_306 (O_306,N_2978,N_2415);
or UO_307 (O_307,N_2518,N_2542);
nand UO_308 (O_308,N_2525,N_2758);
nand UO_309 (O_309,N_2963,N_2795);
nor UO_310 (O_310,N_2690,N_2927);
xor UO_311 (O_311,N_2297,N_2990);
nand UO_312 (O_312,N_2468,N_2845);
xor UO_313 (O_313,N_2997,N_2433);
nor UO_314 (O_314,N_2714,N_2289);
xnor UO_315 (O_315,N_2994,N_2719);
or UO_316 (O_316,N_2319,N_2723);
and UO_317 (O_317,N_2853,N_2939);
and UO_318 (O_318,N_2925,N_2389);
nand UO_319 (O_319,N_2694,N_2914);
xor UO_320 (O_320,N_2743,N_2980);
nand UO_321 (O_321,N_2766,N_2298);
or UO_322 (O_322,N_2826,N_2584);
and UO_323 (O_323,N_2950,N_2908);
or UO_324 (O_324,N_2613,N_2773);
xnor UO_325 (O_325,N_2332,N_2945);
or UO_326 (O_326,N_2506,N_2303);
nor UO_327 (O_327,N_2534,N_2577);
xnor UO_328 (O_328,N_2481,N_2395);
xnor UO_329 (O_329,N_2972,N_2480);
xor UO_330 (O_330,N_2293,N_2260);
xor UO_331 (O_331,N_2703,N_2538);
nor UO_332 (O_332,N_2862,N_2755);
and UO_333 (O_333,N_2967,N_2907);
or UO_334 (O_334,N_2556,N_2669);
nand UO_335 (O_335,N_2724,N_2704);
xor UO_336 (O_336,N_2642,N_2663);
nor UO_337 (O_337,N_2426,N_2463);
nor UO_338 (O_338,N_2325,N_2679);
or UO_339 (O_339,N_2333,N_2522);
and UO_340 (O_340,N_2634,N_2658);
nor UO_341 (O_341,N_2417,N_2517);
nand UO_342 (O_342,N_2374,N_2929);
and UO_343 (O_343,N_2675,N_2655);
or UO_344 (O_344,N_2256,N_2672);
and UO_345 (O_345,N_2811,N_2959);
xor UO_346 (O_346,N_2254,N_2531);
nor UO_347 (O_347,N_2868,N_2681);
xor UO_348 (O_348,N_2691,N_2951);
nor UO_349 (O_349,N_2275,N_2369);
xor UO_350 (O_350,N_2326,N_2329);
xor UO_351 (O_351,N_2392,N_2761);
or UO_352 (O_352,N_2810,N_2693);
or UO_353 (O_353,N_2832,N_2804);
nor UO_354 (O_354,N_2354,N_2977);
nor UO_355 (O_355,N_2601,N_2736);
or UO_356 (O_356,N_2509,N_2689);
nor UO_357 (O_357,N_2431,N_2435);
or UO_358 (O_358,N_2295,N_2651);
nor UO_359 (O_359,N_2311,N_2891);
nand UO_360 (O_360,N_2423,N_2317);
nor UO_361 (O_361,N_2871,N_2624);
xnor UO_362 (O_362,N_2510,N_2608);
nand UO_363 (O_363,N_2437,N_2713);
or UO_364 (O_364,N_2884,N_2346);
nor UO_365 (O_365,N_2831,N_2308);
nand UO_366 (O_366,N_2352,N_2381);
xnor UO_367 (O_367,N_2683,N_2878);
xor UO_368 (O_368,N_2600,N_2623);
or UO_369 (O_369,N_2388,N_2475);
or UO_370 (O_370,N_2774,N_2549);
nand UO_371 (O_371,N_2576,N_2956);
or UO_372 (O_372,N_2911,N_2492);
nand UO_373 (O_373,N_2453,N_2444);
nor UO_374 (O_374,N_2780,N_2712);
and UO_375 (O_375,N_2819,N_2502);
nand UO_376 (O_376,N_2943,N_2647);
xnor UO_377 (O_377,N_2869,N_2516);
xnor UO_378 (O_378,N_2738,N_2649);
nand UO_379 (O_379,N_2325,N_2991);
xnor UO_380 (O_380,N_2456,N_2977);
and UO_381 (O_381,N_2543,N_2353);
nor UO_382 (O_382,N_2366,N_2478);
nand UO_383 (O_383,N_2818,N_2845);
and UO_384 (O_384,N_2499,N_2430);
nand UO_385 (O_385,N_2570,N_2984);
xor UO_386 (O_386,N_2699,N_2489);
and UO_387 (O_387,N_2863,N_2530);
and UO_388 (O_388,N_2987,N_2495);
nor UO_389 (O_389,N_2473,N_2333);
and UO_390 (O_390,N_2509,N_2374);
and UO_391 (O_391,N_2577,N_2811);
xnor UO_392 (O_392,N_2907,N_2404);
and UO_393 (O_393,N_2688,N_2793);
xor UO_394 (O_394,N_2782,N_2936);
nor UO_395 (O_395,N_2850,N_2670);
xor UO_396 (O_396,N_2483,N_2325);
xor UO_397 (O_397,N_2535,N_2807);
nor UO_398 (O_398,N_2801,N_2448);
xor UO_399 (O_399,N_2525,N_2590);
nand UO_400 (O_400,N_2412,N_2292);
and UO_401 (O_401,N_2556,N_2651);
xor UO_402 (O_402,N_2464,N_2833);
xnor UO_403 (O_403,N_2399,N_2737);
xnor UO_404 (O_404,N_2720,N_2867);
xnor UO_405 (O_405,N_2459,N_2796);
xnor UO_406 (O_406,N_2422,N_2948);
or UO_407 (O_407,N_2752,N_2872);
or UO_408 (O_408,N_2356,N_2708);
xnor UO_409 (O_409,N_2951,N_2805);
or UO_410 (O_410,N_2818,N_2253);
nor UO_411 (O_411,N_2972,N_2394);
nor UO_412 (O_412,N_2531,N_2789);
and UO_413 (O_413,N_2333,N_2927);
nand UO_414 (O_414,N_2605,N_2584);
xor UO_415 (O_415,N_2569,N_2923);
or UO_416 (O_416,N_2727,N_2400);
nor UO_417 (O_417,N_2618,N_2979);
nand UO_418 (O_418,N_2364,N_2882);
or UO_419 (O_419,N_2308,N_2747);
xnor UO_420 (O_420,N_2312,N_2781);
nand UO_421 (O_421,N_2517,N_2926);
nor UO_422 (O_422,N_2466,N_2645);
xor UO_423 (O_423,N_2878,N_2432);
nor UO_424 (O_424,N_2970,N_2555);
and UO_425 (O_425,N_2762,N_2865);
nor UO_426 (O_426,N_2657,N_2786);
nand UO_427 (O_427,N_2879,N_2823);
and UO_428 (O_428,N_2581,N_2250);
xnor UO_429 (O_429,N_2793,N_2733);
nor UO_430 (O_430,N_2774,N_2907);
xnor UO_431 (O_431,N_2856,N_2748);
nand UO_432 (O_432,N_2945,N_2928);
xor UO_433 (O_433,N_2621,N_2601);
nand UO_434 (O_434,N_2283,N_2516);
and UO_435 (O_435,N_2441,N_2393);
nor UO_436 (O_436,N_2907,N_2545);
nor UO_437 (O_437,N_2535,N_2679);
nor UO_438 (O_438,N_2488,N_2449);
nor UO_439 (O_439,N_2356,N_2890);
xnor UO_440 (O_440,N_2890,N_2484);
nand UO_441 (O_441,N_2570,N_2545);
nand UO_442 (O_442,N_2390,N_2713);
xor UO_443 (O_443,N_2642,N_2330);
and UO_444 (O_444,N_2400,N_2810);
or UO_445 (O_445,N_2398,N_2323);
nand UO_446 (O_446,N_2820,N_2689);
xnor UO_447 (O_447,N_2392,N_2487);
and UO_448 (O_448,N_2976,N_2904);
and UO_449 (O_449,N_2488,N_2656);
and UO_450 (O_450,N_2581,N_2941);
and UO_451 (O_451,N_2657,N_2357);
nand UO_452 (O_452,N_2801,N_2884);
nor UO_453 (O_453,N_2846,N_2622);
or UO_454 (O_454,N_2350,N_2522);
or UO_455 (O_455,N_2299,N_2880);
nor UO_456 (O_456,N_2995,N_2594);
and UO_457 (O_457,N_2915,N_2742);
nor UO_458 (O_458,N_2669,N_2383);
nand UO_459 (O_459,N_2417,N_2543);
xnor UO_460 (O_460,N_2673,N_2588);
xnor UO_461 (O_461,N_2900,N_2688);
and UO_462 (O_462,N_2775,N_2844);
and UO_463 (O_463,N_2877,N_2889);
and UO_464 (O_464,N_2398,N_2284);
xnor UO_465 (O_465,N_2312,N_2318);
nor UO_466 (O_466,N_2323,N_2394);
and UO_467 (O_467,N_2974,N_2936);
xor UO_468 (O_468,N_2459,N_2437);
nor UO_469 (O_469,N_2549,N_2752);
nand UO_470 (O_470,N_2694,N_2303);
xor UO_471 (O_471,N_2931,N_2925);
or UO_472 (O_472,N_2522,N_2690);
and UO_473 (O_473,N_2572,N_2924);
nor UO_474 (O_474,N_2411,N_2953);
xnor UO_475 (O_475,N_2678,N_2618);
xor UO_476 (O_476,N_2627,N_2609);
nand UO_477 (O_477,N_2541,N_2848);
or UO_478 (O_478,N_2800,N_2792);
nor UO_479 (O_479,N_2358,N_2919);
and UO_480 (O_480,N_2311,N_2303);
nand UO_481 (O_481,N_2649,N_2605);
and UO_482 (O_482,N_2273,N_2313);
nand UO_483 (O_483,N_2479,N_2705);
nor UO_484 (O_484,N_2973,N_2507);
nand UO_485 (O_485,N_2837,N_2974);
nand UO_486 (O_486,N_2698,N_2993);
and UO_487 (O_487,N_2313,N_2371);
or UO_488 (O_488,N_2268,N_2924);
and UO_489 (O_489,N_2988,N_2411);
xnor UO_490 (O_490,N_2866,N_2791);
nor UO_491 (O_491,N_2403,N_2452);
nor UO_492 (O_492,N_2280,N_2508);
nand UO_493 (O_493,N_2917,N_2313);
nand UO_494 (O_494,N_2981,N_2796);
and UO_495 (O_495,N_2293,N_2328);
nor UO_496 (O_496,N_2304,N_2322);
nor UO_497 (O_497,N_2627,N_2703);
and UO_498 (O_498,N_2768,N_2641);
nor UO_499 (O_499,N_2550,N_2412);
endmodule