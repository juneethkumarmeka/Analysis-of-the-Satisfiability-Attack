module basic_2500_25000_3000_50_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nand U0 (N_0,In_2189,In_1207);
and U1 (N_1,In_2121,In_1719);
and U2 (N_2,In_678,In_576);
and U3 (N_3,In_1204,In_964);
nor U4 (N_4,In_1673,In_112);
or U5 (N_5,In_743,In_188);
nor U6 (N_6,In_1159,In_1331);
or U7 (N_7,In_905,In_812);
nand U8 (N_8,In_1452,In_2285);
xor U9 (N_9,In_2295,In_918);
nand U10 (N_10,In_582,In_1200);
xnor U11 (N_11,In_953,In_445);
or U12 (N_12,In_197,In_2237);
or U13 (N_13,In_2430,In_1541);
nand U14 (N_14,In_1524,In_1744);
and U15 (N_15,In_2082,In_2396);
nand U16 (N_16,In_532,In_2427);
xnor U17 (N_17,In_1471,In_1013);
or U18 (N_18,In_1948,In_2131);
nor U19 (N_19,In_1727,In_13);
or U20 (N_20,In_1988,In_2315);
nand U21 (N_21,In_1255,In_585);
and U22 (N_22,In_1298,In_2344);
xnor U23 (N_23,In_1632,In_1151);
or U24 (N_24,In_958,In_876);
xnor U25 (N_25,In_1281,In_1350);
and U26 (N_26,In_2196,In_1691);
or U27 (N_27,In_1770,In_2221);
or U28 (N_28,In_1001,In_1902);
nor U29 (N_29,In_2041,In_895);
nor U30 (N_30,In_1669,In_496);
and U31 (N_31,In_2087,In_1737);
xnor U32 (N_32,In_611,In_2277);
xor U33 (N_33,In_1733,In_1143);
xnor U34 (N_34,In_829,In_1370);
nand U35 (N_35,In_1112,In_1163);
xor U36 (N_36,In_1037,In_815);
nand U37 (N_37,In_1484,In_365);
xor U38 (N_38,In_971,In_38);
or U39 (N_39,In_909,In_708);
nor U40 (N_40,In_1111,In_482);
and U41 (N_41,In_2266,In_2472);
or U42 (N_42,In_1102,In_1138);
and U43 (N_43,In_1392,In_1100);
nand U44 (N_44,In_942,In_465);
xnor U45 (N_45,In_258,In_646);
and U46 (N_46,In_252,In_1650);
nand U47 (N_47,In_650,In_54);
nand U48 (N_48,In_1859,In_64);
xnor U49 (N_49,In_200,In_343);
nand U50 (N_50,In_67,In_270);
xor U51 (N_51,In_2089,In_1269);
and U52 (N_52,In_1630,In_34);
nor U53 (N_53,In_619,In_1713);
and U54 (N_54,In_2370,In_1542);
xnor U55 (N_55,In_658,In_291);
nor U56 (N_56,In_1603,In_1909);
and U57 (N_57,In_442,In_2003);
nand U58 (N_58,In_693,In_689);
nand U59 (N_59,In_840,In_1879);
or U60 (N_60,In_584,In_1206);
and U61 (N_61,In_1870,In_2416);
nor U62 (N_62,In_1181,In_2387);
and U63 (N_63,In_849,In_2167);
and U64 (N_64,In_1208,In_775);
nand U65 (N_65,In_85,In_2479);
or U66 (N_66,In_627,In_2020);
nand U67 (N_67,In_1365,In_901);
nand U68 (N_68,In_1494,In_336);
and U69 (N_69,In_457,In_2239);
nor U70 (N_70,In_1394,In_1134);
nor U71 (N_71,In_912,In_2160);
xor U72 (N_72,In_1294,In_441);
nor U73 (N_73,In_2234,In_1817);
nand U74 (N_74,In_2246,In_158);
or U75 (N_75,In_2108,In_1818);
nor U76 (N_76,In_305,In_667);
nand U77 (N_77,In_104,In_512);
nor U78 (N_78,In_1676,In_822);
or U79 (N_79,In_1738,In_1462);
nand U80 (N_80,In_525,In_1186);
xnor U81 (N_81,In_295,In_558);
and U82 (N_82,In_2325,In_769);
or U83 (N_83,In_2471,In_1055);
nand U84 (N_84,In_599,In_1447);
nand U85 (N_85,In_1606,In_2179);
and U86 (N_86,In_366,In_1108);
xor U87 (N_87,In_488,In_1481);
nand U88 (N_88,In_1495,In_81);
xor U89 (N_89,In_1074,In_1604);
nor U90 (N_90,In_87,In_925);
xnor U91 (N_91,In_641,In_334);
nor U92 (N_92,In_861,In_1157);
xor U93 (N_93,In_987,In_1476);
and U94 (N_94,In_1141,In_1465);
or U95 (N_95,In_2203,In_390);
and U96 (N_96,In_2352,In_1071);
or U97 (N_97,In_2200,In_2092);
xor U98 (N_98,In_317,In_2068);
xnor U99 (N_99,In_1537,In_893);
or U100 (N_100,In_817,In_1075);
nor U101 (N_101,In_344,In_2126);
and U102 (N_102,In_537,In_2429);
xor U103 (N_103,In_202,In_1527);
nand U104 (N_104,In_2379,In_2495);
or U105 (N_105,In_2103,In_1881);
or U106 (N_106,In_836,In_2313);
nor U107 (N_107,In_1964,In_2447);
nand U108 (N_108,In_621,In_312);
nor U109 (N_109,In_320,In_51);
nand U110 (N_110,In_1982,In_1000);
or U111 (N_111,In_345,In_950);
xor U112 (N_112,In_1778,In_740);
and U113 (N_113,In_2097,In_278);
nor U114 (N_114,In_2454,In_164);
or U115 (N_115,In_1219,In_567);
or U116 (N_116,In_2415,In_1608);
nor U117 (N_117,In_123,In_1903);
or U118 (N_118,In_1026,In_1963);
and U119 (N_119,In_91,In_1862);
xnor U120 (N_120,In_1573,In_1979);
nand U121 (N_121,In_1498,In_157);
nand U122 (N_122,In_1786,In_2127);
nand U123 (N_123,In_1863,In_1414);
xnor U124 (N_124,In_1344,In_1795);
nand U125 (N_125,In_721,In_2371);
xnor U126 (N_126,In_1296,In_1554);
and U127 (N_127,In_1101,In_141);
and U128 (N_128,In_1272,In_2268);
or U129 (N_129,In_1671,In_311);
xor U130 (N_130,In_290,In_555);
or U131 (N_131,In_1560,In_1656);
nand U132 (N_132,In_139,In_761);
nor U133 (N_133,In_2073,In_348);
xnor U134 (N_134,In_520,In_1087);
nand U135 (N_135,In_2141,In_423);
and U136 (N_136,In_122,In_435);
nor U137 (N_137,In_2069,In_2044);
nand U138 (N_138,In_1752,In_1999);
or U139 (N_139,In_2485,In_1872);
xnor U140 (N_140,In_1068,In_982);
xnor U141 (N_141,In_31,In_1580);
xor U142 (N_142,In_1215,In_308);
nor U143 (N_143,In_2349,In_1168);
xor U144 (N_144,In_86,In_694);
xor U145 (N_145,In_1287,In_2300);
and U146 (N_146,In_1299,In_208);
or U147 (N_147,In_1592,In_374);
xnor U148 (N_148,In_951,In_923);
and U149 (N_149,In_604,In_709);
nand U150 (N_150,In_484,In_1959);
nand U151 (N_151,In_2148,In_2445);
or U152 (N_152,In_371,In_381);
nor U153 (N_153,In_1658,In_975);
or U154 (N_154,In_945,In_917);
or U155 (N_155,In_786,In_1225);
and U156 (N_156,In_1285,In_767);
or U157 (N_157,In_172,In_2305);
xnor U158 (N_158,In_2362,In_2381);
or U159 (N_159,In_1397,In_1758);
nand U160 (N_160,In_1193,In_1639);
xnor U161 (N_161,In_1239,In_1563);
or U162 (N_162,In_700,In_1077);
or U163 (N_163,In_1472,In_924);
nor U164 (N_164,In_2223,In_2135);
xor U165 (N_165,In_885,In_970);
nor U166 (N_166,In_105,In_1336);
and U167 (N_167,In_1871,In_1289);
and U168 (N_168,In_352,In_1492);
or U169 (N_169,In_2130,In_1785);
or U170 (N_170,In_375,In_102);
or U171 (N_171,In_404,In_1304);
nand U172 (N_172,In_359,In_1939);
or U173 (N_173,In_1437,In_376);
or U174 (N_174,In_1850,In_1990);
xor U175 (N_175,In_427,In_233);
nand U176 (N_176,In_1073,In_1060);
and U177 (N_177,In_960,In_1516);
and U178 (N_178,In_1780,In_2410);
nor U179 (N_179,In_230,In_56);
and U180 (N_180,In_1968,In_115);
xnor U181 (N_181,In_1984,In_1756);
nor U182 (N_182,In_1051,In_1806);
xor U183 (N_183,In_287,In_1805);
nor U184 (N_184,In_1897,In_1257);
or U185 (N_185,In_307,In_811);
and U186 (N_186,In_2122,In_755);
and U187 (N_187,In_262,In_706);
nor U188 (N_188,In_2154,In_2156);
or U189 (N_189,In_2259,In_1403);
nand U190 (N_190,In_741,In_2132);
nand U191 (N_191,In_841,In_1677);
nor U192 (N_192,In_1674,In_2047);
nor U193 (N_193,In_43,In_699);
nor U194 (N_194,In_670,In_96);
xnor U195 (N_195,In_1624,In_957);
or U196 (N_196,In_2348,In_2010);
or U197 (N_197,In_1464,In_2107);
or U198 (N_198,In_28,In_518);
nand U199 (N_199,In_2438,In_421);
nor U200 (N_200,In_1653,In_1904);
and U201 (N_201,In_2399,In_2441);
nand U202 (N_202,In_926,In_2390);
nand U203 (N_203,In_1381,In_2011);
nor U204 (N_204,In_1029,In_797);
nand U205 (N_205,In_826,In_1199);
xnor U206 (N_206,In_1442,In_1547);
nor U207 (N_207,In_1132,In_873);
and U208 (N_208,In_810,In_221);
or U209 (N_209,In_2321,In_1035);
or U210 (N_210,In_2157,In_1006);
nor U211 (N_211,In_1970,In_2473);
or U212 (N_212,In_247,In_527);
nand U213 (N_213,In_63,In_1845);
nor U214 (N_214,In_2317,In_1705);
nand U215 (N_215,In_425,In_595);
xor U216 (N_216,In_1475,In_2493);
xnor U217 (N_217,In_1179,In_408);
xnor U218 (N_218,In_2384,In_827);
nor U219 (N_219,In_219,In_587);
and U220 (N_220,In_48,In_1133);
nand U221 (N_221,In_1218,In_2307);
nor U222 (N_222,In_1998,In_825);
or U223 (N_223,In_1423,In_1076);
nor U224 (N_224,In_322,In_563);
nand U225 (N_225,In_2455,In_2147);
nor U226 (N_226,In_1975,In_1238);
xor U227 (N_227,In_1779,In_1231);
nor U228 (N_228,In_707,In_1341);
and U229 (N_229,In_1877,In_1314);
nor U230 (N_230,In_1406,In_1154);
and U231 (N_231,In_2014,In_673);
xor U232 (N_232,In_1022,In_522);
nor U233 (N_233,In_1918,In_1503);
nor U234 (N_234,In_874,In_1564);
and U235 (N_235,In_996,In_1891);
and U236 (N_236,In_1349,In_939);
nand U237 (N_237,In_1976,In_1091);
and U238 (N_238,In_214,In_898);
nor U239 (N_239,In_931,In_2146);
nand U240 (N_240,In_2161,In_2330);
and U241 (N_241,In_309,In_1109);
xor U242 (N_242,In_758,In_1623);
or U243 (N_243,In_733,In_195);
xor U244 (N_244,In_596,In_380);
and U245 (N_245,In_253,In_1416);
nand U246 (N_246,In_1679,In_422);
xor U247 (N_247,In_517,In_534);
and U248 (N_248,In_903,In_439);
and U249 (N_249,In_2149,In_2474);
and U250 (N_250,In_1966,In_2328);
nor U251 (N_251,In_456,In_2347);
nand U252 (N_252,In_1435,In_326);
nor U253 (N_253,In_1843,In_185);
nor U254 (N_254,In_2091,In_902);
nor U255 (N_255,In_980,In_434);
or U256 (N_256,In_640,In_1633);
nand U257 (N_257,In_1927,In_1142);
nor U258 (N_258,In_2414,In_1252);
nor U259 (N_259,In_437,In_701);
and U260 (N_260,In_1345,In_990);
xnor U261 (N_261,In_1140,In_973);
xnor U262 (N_262,In_1728,In_179);
nand U263 (N_263,In_356,In_1625);
nand U264 (N_264,In_1703,In_1931);
nand U265 (N_265,In_722,In_998);
xnor U266 (N_266,In_377,In_1506);
xnor U267 (N_267,In_2004,In_549);
and U268 (N_268,In_2331,In_175);
nor U269 (N_269,In_572,In_932);
and U270 (N_270,In_1565,In_248);
nor U271 (N_271,In_462,In_93);
nor U272 (N_272,In_1346,In_203);
and U273 (N_273,In_1268,In_145);
and U274 (N_274,In_178,In_1509);
and U275 (N_275,In_686,In_507);
and U276 (N_276,In_2007,In_1613);
and U277 (N_277,In_1059,In_550);
xnor U278 (N_278,In_97,In_2385);
nand U279 (N_279,In_1561,In_1546);
and U280 (N_280,In_1512,In_1764);
or U281 (N_281,In_1690,In_192);
xor U282 (N_282,In_776,In_1688);
or U283 (N_283,In_631,In_639);
nor U284 (N_284,In_273,In_2487);
and U285 (N_285,In_362,In_360);
and U286 (N_286,In_1823,In_400);
and U287 (N_287,In_1522,In_935);
xor U288 (N_288,In_162,In_2282);
nand U289 (N_289,In_2088,In_2120);
nor U290 (N_290,In_1254,In_2338);
or U291 (N_291,In_1905,In_1742);
and U292 (N_292,In_2053,In_744);
nor U293 (N_293,In_796,In_1295);
and U294 (N_294,In_1427,In_1153);
and U295 (N_295,In_2163,In_1274);
nand U296 (N_296,In_1096,In_2065);
nor U297 (N_297,In_1020,In_1167);
and U298 (N_298,In_1648,In_206);
nand U299 (N_299,In_647,In_2383);
nand U300 (N_300,In_994,In_1947);
nand U301 (N_301,In_1267,In_363);
nand U302 (N_302,In_1119,In_1213);
and U303 (N_303,In_341,In_896);
and U304 (N_304,In_1701,In_1558);
and U305 (N_305,In_553,In_1422);
nor U306 (N_306,In_983,In_1064);
and U307 (N_307,In_947,In_2115);
nor U308 (N_308,In_1740,In_2211);
xnor U309 (N_309,In_1513,In_2212);
nand U310 (N_310,In_1155,In_1368);
xor U311 (N_311,In_1960,In_1042);
xor U312 (N_312,In_142,In_2095);
and U313 (N_313,In_430,In_937);
nor U314 (N_314,In_2403,In_2143);
or U315 (N_315,In_2358,In_2378);
or U316 (N_316,In_346,In_78);
and U317 (N_317,In_681,In_1605);
nand U318 (N_318,In_1478,In_1994);
nor U319 (N_319,In_147,In_1681);
xnor U320 (N_320,In_23,In_2094);
and U321 (N_321,In_332,In_20);
nor U322 (N_322,In_2027,In_1875);
xor U323 (N_323,In_2166,In_1115);
xnor U324 (N_324,In_1810,In_2293);
and U325 (N_325,In_862,In_1470);
nand U326 (N_326,In_1293,In_259);
or U327 (N_327,In_494,In_2434);
nor U328 (N_328,In_125,In_715);
nor U329 (N_329,In_1027,In_636);
and U330 (N_330,In_560,In_2116);
or U331 (N_331,In_267,In_2025);
nor U332 (N_332,In_351,In_2210);
nand U333 (N_333,In_547,In_263);
or U334 (N_334,In_729,In_559);
xnor U335 (N_335,In_1644,In_293);
or U336 (N_336,In_2492,In_760);
nor U337 (N_337,In_1849,In_1209);
and U338 (N_338,In_1454,In_1885);
nor U339 (N_339,In_834,In_2476);
or U340 (N_340,In_73,In_1283);
or U341 (N_341,In_154,In_2446);
nand U342 (N_342,In_569,In_807);
nand U343 (N_343,In_1340,In_1820);
and U344 (N_344,In_1233,In_1226);
nor U345 (N_345,In_237,In_1887);
nor U346 (N_346,In_226,In_2428);
xor U347 (N_347,In_2021,In_2102);
xnor U348 (N_348,In_510,In_1259);
and U349 (N_349,In_2288,In_1685);
or U350 (N_350,In_1396,In_1807);
or U351 (N_351,In_402,In_1842);
and U352 (N_352,In_1145,In_2017);
nor U353 (N_353,In_2105,In_1894);
or U354 (N_354,In_418,In_1754);
xnor U355 (N_355,In_2213,In_1388);
and U356 (N_356,In_1695,In_933);
or U357 (N_357,In_657,In_1708);
xnor U358 (N_358,In_2216,In_80);
nor U359 (N_359,In_991,In_2248);
and U360 (N_360,In_2437,In_2114);
xor U361 (N_361,In_1008,In_1874);
nand U362 (N_362,In_571,In_1194);
nand U363 (N_363,In_1348,In_6);
xnor U364 (N_364,In_2228,In_1878);
nor U365 (N_365,In_1171,In_1985);
or U366 (N_366,In_746,In_850);
nor U367 (N_367,In_1487,In_1914);
xor U368 (N_368,In_2261,In_1458);
nand U369 (N_369,In_1360,In_846);
xor U370 (N_370,In_1444,In_2483);
nand U371 (N_371,In_634,In_2458);
or U372 (N_372,In_2243,In_774);
nor U373 (N_373,In_524,In_1665);
nand U374 (N_374,In_1407,In_804);
and U375 (N_375,In_659,In_505);
or U376 (N_376,In_176,In_656);
xnor U377 (N_377,In_2128,In_1347);
xor U378 (N_378,In_1544,In_544);
nand U379 (N_379,In_1932,In_712);
nor U380 (N_380,In_762,In_1356);
nand U381 (N_381,In_1337,In_1821);
nor U382 (N_382,In_1774,In_844);
nand U383 (N_383,In_1655,In_2034);
nand U384 (N_384,In_1363,In_1854);
and U385 (N_385,In_2225,In_1614);
and U386 (N_386,In_1362,In_1330);
or U387 (N_387,In_1236,In_463);
and U388 (N_388,In_2486,In_424);
nand U389 (N_389,In_573,In_1722);
xor U390 (N_390,In_682,In_35);
nor U391 (N_391,In_1716,In_2298);
and U392 (N_392,In_2283,In_899);
xor U393 (N_393,In_606,In_1352);
xnor U394 (N_394,In_82,In_459);
nand U395 (N_395,In_1972,In_454);
nor U396 (N_396,In_99,In_855);
or U397 (N_397,In_1371,In_1057);
and U398 (N_398,In_401,In_564);
xnor U399 (N_399,In_677,In_76);
xnor U400 (N_400,In_1479,In_704);
nand U401 (N_401,In_392,In_1867);
nand U402 (N_402,In_1460,In_2076);
and U403 (N_403,In_1402,In_2245);
nor U404 (N_404,In_1504,In_1989);
or U405 (N_405,In_2098,In_1925);
nand U406 (N_406,In_1196,In_406);
xnor U407 (N_407,In_1583,In_1529);
xnor U408 (N_408,In_1880,In_734);
nand U409 (N_409,In_331,In_1577);
xor U410 (N_410,In_1803,In_2112);
or U411 (N_411,In_808,In_1080);
or U412 (N_412,In_394,In_2155);
and U413 (N_413,In_1014,In_1715);
and U414 (N_414,In_2468,In_1591);
nand U415 (N_415,In_2072,In_2360);
nor U416 (N_416,In_570,In_1528);
or U417 (N_417,In_416,In_283);
nand U418 (N_418,In_372,In_1514);
and U419 (N_419,In_2035,In_1431);
xor U420 (N_420,In_633,In_1599);
and U421 (N_421,In_2327,In_2273);
xnor U422 (N_422,In_913,In_1865);
and U423 (N_423,In_1853,In_2405);
xnor U424 (N_424,In_432,In_329);
and U425 (N_425,In_2319,In_1152);
nor U426 (N_426,In_1343,In_1729);
nand U427 (N_427,In_133,In_2463);
xor U428 (N_428,In_2341,In_218);
or U429 (N_429,In_1316,In_730);
or U430 (N_430,In_1819,In_1212);
nand U431 (N_431,In_2356,In_412);
or U432 (N_432,In_2465,In_1790);
nor U433 (N_433,In_2443,In_720);
nor U434 (N_434,In_791,In_1773);
and U435 (N_435,In_1329,In_100);
xor U436 (N_436,In_961,In_388);
xnor U437 (N_437,In_235,In_18);
and U438 (N_438,In_349,In_49);
nor U439 (N_439,In_1714,In_816);
xnor U440 (N_440,In_954,In_303);
nand U441 (N_441,In_541,In_1611);
and U442 (N_442,In_379,In_2110);
and U443 (N_443,In_2482,In_1019);
and U444 (N_444,In_72,In_2172);
nor U445 (N_445,In_628,In_845);
nor U446 (N_446,In_2113,In_1949);
nand U447 (N_447,In_1572,In_2051);
or U448 (N_448,In_450,In_1389);
xor U449 (N_449,In_1712,In_1243);
and U450 (N_450,In_1686,In_749);
and U451 (N_451,In_735,In_88);
nand U452 (N_452,In_436,In_1463);
xnor U453 (N_453,In_1801,In_1070);
nand U454 (N_454,In_126,In_369);
xor U455 (N_455,In_47,In_1297);
nand U456 (N_456,In_1505,In_491);
or U457 (N_457,In_1868,In_2393);
xor U458 (N_458,In_224,In_2236);
or U459 (N_459,In_2368,In_1266);
and U460 (N_460,In_2395,In_2070);
nor U461 (N_461,In_325,In_1755);
nor U462 (N_462,In_2235,In_2032);
nor U463 (N_463,In_1923,In_33);
nand U464 (N_464,In_2039,In_1228);
or U465 (N_465,In_1775,In_1657);
xor U466 (N_466,In_1830,In_37);
xnor U467 (N_467,In_2409,In_1707);
and U468 (N_468,In_1275,In_2314);
xor U469 (N_469,In_1978,In_1327);
or U470 (N_470,In_429,In_1082);
nand U471 (N_471,In_1488,In_613);
nor U472 (N_472,In_2240,In_66);
nor U473 (N_473,In_1136,In_1223);
and U474 (N_474,In_493,In_62);
nand U475 (N_475,In_231,In_1459);
xor U476 (N_476,In_1915,In_385);
nand U477 (N_477,In_319,In_521);
nand U478 (N_478,In_2180,In_1203);
xor U479 (N_479,In_1493,In_1958);
nor U480 (N_480,In_2013,In_1130);
nand U481 (N_481,In_1626,In_1569);
xor U482 (N_482,In_490,In_552);
or U483 (N_483,In_1496,In_1284);
xor U484 (N_484,In_1873,In_1375);
nor U485 (N_485,In_2018,In_1847);
or U486 (N_486,In_159,In_1602);
nor U487 (N_487,In_1321,In_431);
xor U488 (N_488,In_1137,In_2176);
xnor U489 (N_489,In_2133,In_177);
or U490 (N_490,In_671,In_608);
and U491 (N_491,In_2177,In_1156);
nor U492 (N_492,In_948,In_603);
or U493 (N_493,In_455,In_395);
xnor U494 (N_494,In_1753,In_578);
nor U495 (N_495,In_472,In_819);
or U496 (N_496,In_1763,In_687);
nor U497 (N_497,In_1093,In_1114);
nor U498 (N_498,In_1084,In_1376);
and U499 (N_499,In_892,In_1164);
xor U500 (N_500,In_1081,In_788);
nand U501 (N_501,In_1056,In_1324);
nand U502 (N_502,In_993,In_765);
xnor U503 (N_503,In_2290,In_661);
nand U504 (N_504,In_399,In_275);
or U505 (N_505,In_872,In_1161);
or U506 (N_506,In_2030,N_330);
nand U507 (N_507,In_2144,In_792);
nor U508 (N_508,In_2040,In_668);
nor U509 (N_509,In_1467,In_1067);
and U510 (N_510,In_2253,In_1663);
or U511 (N_511,N_349,In_2181);
and U512 (N_512,In_1757,In_1575);
nand U513 (N_513,In_2392,N_429);
nor U514 (N_514,In_1262,In_2480);
nor U515 (N_515,In_1398,N_71);
or U516 (N_516,N_456,N_482);
and U517 (N_517,In_828,In_272);
nand U518 (N_518,In_1113,N_417);
xnor U519 (N_519,In_1131,In_130);
or U520 (N_520,In_251,In_1800);
nand U521 (N_521,N_77,N_62);
and U522 (N_522,In_852,In_1);
xnor U523 (N_523,N_26,N_361);
xor U524 (N_524,In_1936,In_1216);
nor U525 (N_525,In_70,In_1711);
nor U526 (N_526,In_127,In_1033);
xor U527 (N_527,N_88,N_288);
and U528 (N_528,In_2217,In_2449);
nor U529 (N_529,In_239,In_1117);
or U530 (N_530,In_581,In_2407);
nor U531 (N_531,N_201,In_1767);
xor U532 (N_532,N_310,In_5);
or U533 (N_533,N_411,In_2372);
nor U534 (N_534,N_300,In_41);
and U535 (N_535,In_1310,In_838);
xnor U536 (N_536,N_446,In_2291);
nor U537 (N_537,In_2152,N_332);
and U538 (N_538,In_2165,In_327);
xor U539 (N_539,N_293,In_1973);
xor U540 (N_540,In_2164,In_1997);
and U541 (N_541,In_1974,In_1021);
nor U542 (N_542,In_1461,In_1128);
nor U543 (N_543,In_2323,In_2081);
nor U544 (N_544,In_140,In_2276);
or U545 (N_545,In_1405,In_280);
and U546 (N_546,In_151,N_169);
xnor U547 (N_547,In_95,In_847);
nor U548 (N_548,N_266,In_1002);
or U549 (N_549,In_1610,In_764);
nand U550 (N_550,In_116,In_489);
and U551 (N_551,In_1693,N_74);
or U552 (N_552,N_4,In_717);
xor U553 (N_553,N_408,N_255);
or U554 (N_554,In_1937,In_2150);
and U555 (N_555,In_763,In_995);
xor U556 (N_556,In_568,In_1519);
and U557 (N_557,In_44,In_2101);
and U558 (N_558,In_1832,In_2012);
and U559 (N_559,In_649,In_1649);
nor U560 (N_560,In_1489,In_2138);
nand U561 (N_561,In_1270,In_2294);
or U562 (N_562,In_1121,In_2334);
and U563 (N_563,In_1249,N_51);
nor U564 (N_564,N_412,In_279);
or U565 (N_565,N_393,In_2206);
or U566 (N_566,N_147,In_301);
nor U567 (N_567,In_887,In_1490);
or U568 (N_568,In_1559,In_1172);
nor U569 (N_569,In_156,N_102);
nand U570 (N_570,N_448,N_104);
and U571 (N_571,In_189,In_2475);
nand U572 (N_572,In_1598,N_216);
xor U573 (N_573,In_257,In_1828);
nand U574 (N_574,N_76,In_65);
nand U575 (N_575,N_473,In_1311);
and U576 (N_576,In_1896,In_616);
and U577 (N_577,In_2262,In_234);
and U578 (N_578,In_21,N_33);
nand U579 (N_579,In_675,In_2085);
or U580 (N_580,In_1190,N_59);
and U581 (N_581,N_474,N_127);
nand U582 (N_582,N_25,N_82);
xor U583 (N_583,In_2111,In_1230);
nor U584 (N_584,In_1198,N_381);
or U585 (N_585,In_2380,N_125);
or U586 (N_586,N_441,N_275);
nand U587 (N_587,In_1670,In_39);
nor U588 (N_588,N_222,N_319);
nand U589 (N_589,N_174,In_618);
nor U590 (N_590,In_2366,In_1651);
nor U591 (N_591,In_2028,In_648);
nand U592 (N_592,In_1838,In_2440);
or U593 (N_593,In_652,N_123);
nand U594 (N_594,In_727,In_2351);
xnor U595 (N_595,In_1508,N_164);
xnor U596 (N_596,In_2036,In_1678);
nand U597 (N_597,In_153,In_1248);
nand U598 (N_598,In_1412,In_719);
and U599 (N_599,In_94,In_2345);
and U600 (N_600,N_491,In_963);
nor U601 (N_601,In_1557,In_1421);
nand U602 (N_602,In_389,In_265);
and U603 (N_603,In_1804,In_662);
or U604 (N_604,N_93,In_1095);
nand U605 (N_605,In_1278,In_732);
nand U606 (N_606,In_2241,In_881);
nor U607 (N_607,N_409,In_818);
nor U608 (N_608,N_449,In_1860);
xnor U609 (N_609,In_593,In_1301);
or U610 (N_610,In_543,In_1759);
nand U611 (N_611,In_2208,In_2432);
xnor U612 (N_612,N_471,In_1386);
xor U613 (N_613,In_575,In_1617);
or U614 (N_614,In_222,N_57);
xnor U615 (N_615,In_2099,In_736);
or U616 (N_616,In_897,N_400);
and U617 (N_617,N_132,In_920);
or U618 (N_618,N_252,N_476);
and U619 (N_619,In_118,In_2063);
and U620 (N_620,N_140,In_2139);
nand U621 (N_621,In_1024,In_27);
xor U622 (N_622,In_106,N_463);
nor U623 (N_623,In_138,In_1240);
nand U624 (N_624,N_419,In_1578);
nor U625 (N_625,In_1576,In_413);
or U626 (N_626,In_60,N_53);
or U627 (N_627,In_1680,In_90);
nor U628 (N_628,In_629,In_771);
nand U629 (N_629,In_801,N_168);
and U630 (N_630,In_199,In_986);
or U631 (N_631,In_1277,N_395);
nor U632 (N_632,In_997,In_174);
and U633 (N_633,In_523,In_2287);
or U634 (N_634,In_1784,In_1276);
nand U635 (N_635,In_617,In_979);
or U636 (N_636,In_620,N_486);
nor U637 (N_637,In_426,In_2481);
nor U638 (N_638,N_20,In_2123);
or U639 (N_639,In_877,In_2412);
nor U640 (N_640,In_2006,N_219);
nor U641 (N_641,In_1253,In_446);
or U642 (N_642,In_1652,In_702);
nor U643 (N_643,N_239,In_2364);
nor U644 (N_644,In_2369,In_2142);
and U645 (N_645,In_1306,In_794);
xor U646 (N_646,In_1992,In_1382);
and U647 (N_647,N_402,In_444);
or U648 (N_648,N_439,In_1395);
nand U649 (N_649,In_25,In_2136);
or U650 (N_650,N_133,N_358);
xor U651 (N_651,N_98,N_498);
xnor U652 (N_652,In_2022,In_1353);
xor U653 (N_653,In_168,In_1263);
and U654 (N_654,In_2119,In_2158);
and U655 (N_655,N_28,N_296);
or U656 (N_656,N_321,N_186);
nor U657 (N_657,In_1882,In_398);
xnor U658 (N_658,N_422,In_1919);
and U659 (N_659,In_2340,In_2272);
xnor U660 (N_660,In_1566,In_1025);
nand U661 (N_661,In_2489,N_155);
and U662 (N_662,In_215,N_130);
nand U663 (N_663,In_2312,In_1271);
or U664 (N_664,In_1781,In_802);
nor U665 (N_665,In_1748,N_386);
nor U666 (N_666,N_183,In_2079);
nor U667 (N_667,In_467,In_1718);
or U668 (N_668,N_63,In_1696);
nand U669 (N_669,In_1908,In_1788);
nand U670 (N_670,In_2297,N_470);
nand U671 (N_671,In_1526,In_1468);
nor U672 (N_672,N_279,In_190);
xnor U673 (N_673,In_2219,N_214);
and U674 (N_674,N_259,In_1942);
nor U675 (N_675,N_371,In_989);
nand U676 (N_676,N_475,In_1826);
or U677 (N_677,In_737,In_453);
xnor U678 (N_678,N_284,In_1359);
nand U679 (N_679,In_396,N_243);
nor U680 (N_680,In_1040,N_337);
xor U681 (N_681,In_1050,In_2386);
nor U682 (N_682,In_2151,In_1856);
or U683 (N_683,In_1053,N_205);
nand U684 (N_684,In_1247,N_105);
or U685 (N_685,In_978,In_2491);
or U686 (N_686,N_110,In_1004);
xnor U687 (N_687,In_57,N_148);
xnor U688 (N_688,In_1104,N_285);
nor U689 (N_689,N_397,In_1892);
or U690 (N_690,In_403,N_60);
xor U691 (N_691,In_1265,N_339);
xnor U692 (N_692,In_1917,In_1833);
nand U693 (N_693,N_388,N_220);
xor U694 (N_694,In_2183,In_803);
xnor U695 (N_695,In_2023,In_242);
nor U696 (N_696,In_1393,In_1039);
xor U697 (N_697,N_202,In_2354);
nand U698 (N_698,In_2326,In_298);
nand U699 (N_699,N_128,In_1704);
or U700 (N_700,N_382,In_2118);
xnor U701 (N_701,In_562,In_1258);
nand U702 (N_702,In_1962,N_180);
nor U703 (N_703,N_484,In_124);
and U704 (N_704,In_2000,In_1069);
xnor U705 (N_705,In_1629,In_1010);
nor U706 (N_706,N_12,N_80);
nand U707 (N_707,In_684,In_1579);
xnor U708 (N_708,In_770,N_146);
nor U709 (N_709,In_1661,N_413);
and U710 (N_710,In_2195,In_2400);
nand U711 (N_711,In_651,In_1474);
and U712 (N_712,N_273,In_1308);
xnor U713 (N_713,In_328,In_2460);
xnor U714 (N_714,In_220,In_2140);
nor U715 (N_715,In_2106,In_318);
nor U716 (N_716,In_378,In_672);
xor U717 (N_717,In_193,In_748);
nor U718 (N_718,In_1149,In_725);
xor U719 (N_719,In_1941,In_495);
xor U720 (N_720,N_97,N_217);
or U721 (N_721,In_813,N_256);
xor U722 (N_722,In_1455,N_329);
xor U723 (N_723,In_59,In_1439);
xor U724 (N_724,N_50,N_200);
nand U725 (N_725,In_2071,In_182);
nand U726 (N_726,In_29,In_1411);
xnor U727 (N_727,In_2311,In_83);
or U728 (N_728,N_249,In_713);
nor U729 (N_729,In_1313,In_1366);
nand U730 (N_730,N_410,In_1739);
nor U731 (N_731,In_663,In_831);
nand U732 (N_732,In_692,In_117);
xnor U733 (N_733,In_1169,N_383);
nand U734 (N_734,In_1532,In_1824);
and U735 (N_735,In_1531,In_972);
nand U736 (N_736,In_497,In_1521);
nor U737 (N_737,In_136,N_258);
nand U738 (N_738,N_68,In_475);
xor U739 (N_739,In_256,In_2299);
nand U740 (N_740,In_2420,N_246);
xor U741 (N_741,In_24,In_241);
nor U742 (N_742,In_2230,In_2191);
or U743 (N_743,In_75,In_940);
and U744 (N_744,In_2232,In_1743);
nand U745 (N_745,In_1440,In_1815);
nand U746 (N_746,N_416,N_340);
xnor U747 (N_747,In_289,In_354);
nor U748 (N_748,In_2052,N_276);
xnor U749 (N_749,N_106,In_165);
and U750 (N_750,In_967,In_754);
and U751 (N_751,N_328,In_170);
xor U752 (N_752,In_384,In_1971);
nand U753 (N_753,N_171,In_588);
xnor U754 (N_754,In_806,In_2421);
nor U755 (N_755,In_2361,In_934);
and U756 (N_756,In_2100,N_43);
nor U757 (N_757,In_927,In_2444);
xor U758 (N_758,In_2301,In_451);
nand U759 (N_759,In_2397,N_317);
and U760 (N_760,In_2184,N_23);
and U761 (N_761,In_1288,N_299);
or U762 (N_762,In_137,In_884);
nand U763 (N_763,N_359,N_158);
xor U764 (N_764,In_146,In_46);
nor U765 (N_765,In_889,N_236);
or U766 (N_766,In_1538,N_49);
nand U767 (N_767,N_318,In_784);
nor U768 (N_768,In_1126,N_497);
nor U769 (N_769,In_339,In_42);
xnor U770 (N_770,In_409,In_1787);
xor U771 (N_771,In_1844,In_1646);
xor U772 (N_772,N_418,In_2005);
or U773 (N_773,In_1195,In_601);
nor U774 (N_774,In_1840,N_188);
nor U775 (N_775,N_264,N_465);
xnor U776 (N_776,N_101,N_115);
nand U777 (N_777,In_1058,N_247);
nand U778 (N_778,In_1046,In_1895);
nand U779 (N_779,In_766,In_1229);
or U780 (N_780,In_1952,In_1898);
nand U781 (N_781,In_1745,In_492);
xnor U782 (N_782,In_1099,N_472);
or U783 (N_783,N_179,In_1814);
xnor U784 (N_784,In_2055,In_1072);
or U785 (N_785,In_1436,In_1957);
xnor U786 (N_786,In_1326,N_434);
nor U787 (N_787,In_592,In_1036);
nor U788 (N_788,N_142,In_414);
nand U789 (N_789,N_213,N_89);
and U790 (N_790,N_336,N_477);
nor U791 (N_791,In_2064,N_160);
nor U792 (N_792,In_428,In_411);
xor U793 (N_793,In_502,In_2218);
or U794 (N_794,In_1907,In_1640);
nor U795 (N_795,In_2309,N_163);
nand U796 (N_796,N_490,In_361);
xnor U797 (N_797,N_100,In_1771);
xor U798 (N_798,In_886,In_660);
and U799 (N_799,N_167,N_40);
xnor U800 (N_800,N_399,N_185);
nor U801 (N_801,In_2324,N_39);
nor U802 (N_802,In_1144,In_968);
nand U803 (N_803,In_103,In_2388);
or U804 (N_804,In_1709,N_107);
or U805 (N_805,In_1282,In_1697);
xnor U806 (N_806,In_1802,In_1731);
and U807 (N_807,In_921,In_281);
nor U808 (N_808,N_48,In_625);
xor U809 (N_809,In_2278,In_304);
and U810 (N_810,In_2339,In_53);
nand U811 (N_811,In_1433,In_2424);
nor U812 (N_812,N_153,In_2359);
or U813 (N_813,In_129,In_548);
and U814 (N_814,N_195,In_2350);
nand U815 (N_815,In_1760,In_1593);
xor U816 (N_816,N_257,In_274);
nor U817 (N_817,In_870,In_109);
xor U818 (N_818,In_1609,In_306);
xnor U819 (N_819,N_335,In_1664);
nand U820 (N_820,In_1510,In_1857);
nor U821 (N_821,In_1342,In_2054);
and U822 (N_822,In_2093,N_267);
xor U823 (N_823,In_1995,In_1906);
xor U824 (N_824,In_1858,In_1227);
nor U825 (N_825,In_2043,In_688);
and U826 (N_826,In_26,N_14);
nand U827 (N_827,N_487,In_2185);
xor U828 (N_828,N_352,In_697);
nor U829 (N_829,In_882,In_679);
nand U830 (N_830,In_2357,N_323);
nand U831 (N_831,In_1201,In_2335);
nor U832 (N_832,In_2190,In_878);
xnor U833 (N_833,In_1698,In_500);
nor U834 (N_834,In_1497,In_1237);
nand U835 (N_835,In_928,N_341);
and U836 (N_836,N_280,In_2086);
and U837 (N_837,In_286,In_1920);
xor U838 (N_838,In_1574,In_914);
nand U839 (N_839,In_1762,In_598);
nor U840 (N_840,N_209,N_211);
and U841 (N_841,In_1534,N_390);
xor U842 (N_842,In_1827,In_2037);
and U843 (N_843,In_1234,N_152);
nand U844 (N_844,N_166,In_12);
or U845 (N_845,N_268,In_52);
nand U846 (N_846,In_1041,In_907);
nand U847 (N_847,In_1637,In_1938);
xor U848 (N_848,N_302,N_154);
nand U849 (N_849,N_52,N_141);
nand U850 (N_850,In_966,In_1162);
xor U851 (N_851,In_1515,In_1910);
or U852 (N_852,In_447,In_664);
xor U853 (N_853,In_1482,In_842);
and U854 (N_854,In_1749,In_1486);
xnor U855 (N_855,In_2320,In_1769);
or U856 (N_856,In_1930,In_155);
and U857 (N_857,In_114,N_357);
or U858 (N_858,In_1023,N_99);
or U859 (N_859,In_1636,N_263);
nor U860 (N_860,In_296,In_2247);
nor U861 (N_861,N_415,In_364);
xor U862 (N_862,In_2418,In_15);
or U863 (N_863,N_391,In_477);
or U864 (N_864,N_78,N_234);
nor U865 (N_865,In_217,N_187);
nand U866 (N_866,In_315,N_363);
nand U867 (N_867,In_1499,In_781);
nor U868 (N_868,In_936,N_248);
xor U869 (N_869,In_772,In_2201);
or U870 (N_870,In_1441,In_1783);
or U871 (N_871,In_1940,In_583);
xor U872 (N_872,In_1135,In_1816);
or U873 (N_873,In_941,In_832);
or U874 (N_874,In_2096,N_309);
xor U875 (N_875,In_1191,In_2451);
and U876 (N_876,In_171,In_468);
nor U877 (N_877,In_904,N_13);
xnor U878 (N_878,In_1045,N_121);
and U879 (N_879,In_1015,In_163);
and U880 (N_880,N_29,In_1950);
and U881 (N_881,In_1725,In_1250);
or U882 (N_882,In_1086,In_1720);
or U883 (N_883,In_962,In_160);
xnor U884 (N_884,In_2342,N_66);
or U885 (N_885,In_1672,N_438);
xnor U886 (N_886,In_837,N_269);
and U887 (N_887,In_999,In_2174);
and U888 (N_888,In_2498,In_77);
xnor U889 (N_889,In_2066,In_1016);
nor U890 (N_890,N_372,In_843);
and U891 (N_891,In_922,In_2171);
nand U892 (N_892,In_1700,In_386);
or U893 (N_893,In_250,In_1548);
xnor U894 (N_894,In_2257,N_10);
or U895 (N_895,In_1549,In_1214);
or U896 (N_896,In_871,In_2346);
nor U897 (N_897,N_233,In_1848);
and U898 (N_898,In_1600,In_503);
or U899 (N_899,In_739,N_421);
and U900 (N_900,In_745,N_442);
nand U901 (N_901,In_1846,In_789);
or U902 (N_902,In_1399,N_461);
nor U903 (N_903,N_61,In_1063);
and U904 (N_904,In_910,In_1415);
nor U905 (N_905,In_1721,In_2129);
and U906 (N_906,In_2329,In_2450);
or U907 (N_907,In_1876,In_985);
or U908 (N_908,In_45,N_27);
nand U909 (N_909,In_1595,In_1855);
or U910 (N_910,In_448,In_2457);
or U911 (N_911,In_2436,N_54);
nor U912 (N_912,In_622,In_705);
nand U913 (N_913,In_1540,N_32);
xnor U914 (N_914,In_891,In_1834);
or U915 (N_915,In_915,In_1706);
nor U916 (N_916,In_2205,In_888);
and U917 (N_917,In_919,In_614);
or U918 (N_918,In_976,In_2402);
and U919 (N_919,N_291,In_1668);
and U920 (N_920,In_2249,N_231);
and U921 (N_921,In_1641,N_172);
xnor U922 (N_922,In_529,In_1419);
or U923 (N_923,N_194,In_1980);
nand U924 (N_924,In_1429,N_251);
nor U925 (N_925,N_362,In_2398);
nand U926 (N_926,N_314,In_1635);
nand U927 (N_927,N_122,N_69);
nor U928 (N_928,In_368,N_348);
or U929 (N_929,In_1634,N_199);
nand U930 (N_930,In_201,In_2109);
or U931 (N_931,In_449,In_0);
nor U932 (N_932,In_2153,In_2494);
xnor U933 (N_933,In_186,In_2274);
and U934 (N_934,In_1689,In_410);
xor U935 (N_935,In_580,In_1007);
and U936 (N_936,N_75,In_2296);
nor U937 (N_937,In_198,In_1586);
xor U938 (N_938,In_690,N_450);
and U939 (N_939,In_1502,In_1260);
xor U940 (N_940,N_38,N_385);
nor U941 (N_941,N_150,In_2302);
or U942 (N_942,In_184,N_297);
xnor U943 (N_943,N_120,In_974);
nand U944 (N_944,In_561,N_7);
nand U945 (N_945,In_1734,In_1383);
nor U946 (N_946,In_1951,In_731);
xor U947 (N_947,In_1457,In_1571);
nand U948 (N_948,In_959,In_1332);
xor U949 (N_949,N_143,In_1085);
nor U950 (N_950,In_2422,In_805);
nand U951 (N_951,In_1986,In_2169);
and U952 (N_952,In_1480,In_1182);
nor U953 (N_953,In_790,N_113);
xnor U954 (N_954,N_460,In_1413);
or U955 (N_955,In_1323,In_1615);
or U956 (N_956,In_1552,In_787);
or U957 (N_957,N_261,In_2477);
and U958 (N_958,In_2467,N_157);
nor U959 (N_959,In_440,N_56);
xnor U960 (N_960,In_1987,In_1643);
or U961 (N_961,In_1092,In_297);
and U962 (N_962,In_314,In_2059);
xnor U963 (N_963,In_144,In_355);
and U964 (N_964,In_1122,N_137);
nor U965 (N_965,In_1525,In_9);
xor U966 (N_966,In_485,N_119);
nand U967 (N_967,N_338,In_1003);
and U968 (N_968,N_375,N_206);
xor U969 (N_969,In_1380,N_316);
xnor U970 (N_970,In_2411,In_1235);
and U971 (N_971,In_2038,In_2255);
and U972 (N_972,In_1409,In_1189);
xor U973 (N_973,In_1401,In_1116);
nand U974 (N_974,In_782,In_875);
or U975 (N_975,In_516,In_542);
xnor U976 (N_976,In_2401,In_814);
xor U977 (N_977,In_1694,In_299);
or U978 (N_978,In_277,In_1724);
and U979 (N_979,N_407,In_321);
or U980 (N_980,In_1123,In_1339);
nor U981 (N_981,N_369,In_610);
and U982 (N_982,In_98,In_780);
nor U983 (N_983,N_345,In_626);
or U984 (N_984,In_2029,In_1139);
or U985 (N_985,In_655,N_235);
nand U986 (N_986,In_2074,In_1318);
nor U987 (N_987,N_380,In_1166);
nor U988 (N_988,In_1302,In_1038);
nor U989 (N_989,In_768,N_218);
nor U990 (N_990,In_101,In_865);
and U991 (N_991,N_308,In_1018);
nand U992 (N_992,N_208,In_1926);
nand U993 (N_993,In_1083,In_1286);
or U994 (N_994,In_1094,In_868);
xnor U995 (N_995,In_40,In_1511);
or U996 (N_996,N_16,In_2254);
or U997 (N_997,In_1120,In_1424);
or U998 (N_998,In_1107,In_1264);
xor U999 (N_999,In_1372,In_908);
and U1000 (N_1000,N_37,N_134);
nand U1001 (N_1001,In_131,In_1619);
nor U1002 (N_1002,N_793,N_374);
xor U1003 (N_1003,N_805,In_879);
xnor U1004 (N_1004,In_1921,In_1556);
or U1005 (N_1005,In_2419,N_83);
nor U1006 (N_1006,In_546,In_946);
nor U1007 (N_1007,N_598,In_1106);
or U1008 (N_1008,In_1291,N_801);
nor U1009 (N_1009,N_733,N_396);
or U1010 (N_1010,N_55,N_581);
xor U1011 (N_1011,N_307,N_535);
and U1012 (N_1012,N_58,In_1812);
xnor U1013 (N_1013,In_110,In_438);
and U1014 (N_1014,N_962,N_162);
or U1015 (N_1015,In_350,In_32);
nor U1016 (N_1016,N_283,In_2286);
and U1017 (N_1017,N_654,In_751);
xnor U1018 (N_1018,In_55,N_212);
or U1019 (N_1019,N_84,N_271);
nand U1020 (N_1020,N_627,N_840);
nand U1021 (N_1021,In_820,In_1148);
xnor U1022 (N_1022,N_516,N_468);
nor U1023 (N_1023,In_1777,In_1220);
or U1024 (N_1024,In_1589,In_798);
and U1025 (N_1025,N_617,N_343);
nand U1026 (N_1026,N_350,N_680);
nand U1027 (N_1027,In_795,In_1290);
and U1028 (N_1028,In_209,In_69);
or U1029 (N_1029,In_1682,N_70);
nand U1030 (N_1030,In_1977,N_833);
nor U1031 (N_1031,N_671,N_697);
and U1032 (N_1032,In_108,In_1645);
nor U1033 (N_1033,In_1751,N_718);
or U1034 (N_1034,N_931,In_930);
or U1035 (N_1035,In_238,N_191);
and U1036 (N_1036,In_120,N_679);
and U1037 (N_1037,In_1150,N_333);
nand U1038 (N_1038,N_842,In_1622);
nor U1039 (N_1039,In_1954,In_753);
nor U1040 (N_1040,In_988,N_517);
xnor U1041 (N_1041,In_1945,In_848);
and U1042 (N_1042,In_2242,In_204);
and U1043 (N_1043,N_695,In_1981);
nor U1044 (N_1044,N_737,N_716);
or U1045 (N_1045,In_860,N_272);
or U1046 (N_1046,In_2008,N_994);
nand U1047 (N_1047,N_794,N_898);
nor U1048 (N_1048,In_19,N_609);
xnor U1049 (N_1049,In_2231,In_1187);
nor U1050 (N_1050,In_1723,In_2496);
or U1051 (N_1051,N_230,N_897);
nor U1052 (N_1052,N_519,In_17);
or U1053 (N_1053,N_640,N_736);
and U1054 (N_1054,N_72,In_2453);
nand U1055 (N_1055,N_481,In_1118);
xor U1056 (N_1056,In_107,N_943);
nor U1057 (N_1057,In_2056,In_1809);
and U1058 (N_1058,N_451,In_1408);
and U1059 (N_1059,In_1776,In_2188);
or U1060 (N_1060,In_1692,N_774);
nor U1061 (N_1061,N_564,N_877);
xor U1062 (N_1062,In_612,N_156);
nand U1063 (N_1063,N_687,N_813);
xnor U1064 (N_1064,In_1184,In_1079);
and U1065 (N_1065,In_2367,N_177);
nand U1066 (N_1066,N_605,In_665);
and U1067 (N_1067,N_991,N_867);
or U1068 (N_1068,N_770,In_1924);
and U1069 (N_1069,In_1065,N_538);
nor U1070 (N_1070,In_433,In_324);
nor U1071 (N_1071,N_865,N_221);
nand U1072 (N_1072,In_859,N_301);
or U1073 (N_1073,In_1953,In_243);
xor U1074 (N_1074,N_747,In_58);
and U1075 (N_1075,N_758,N_922);
nor U1076 (N_1076,N_632,N_776);
nor U1077 (N_1077,In_1841,In_1443);
nor U1078 (N_1078,In_2244,N_954);
and U1079 (N_1079,In_696,In_2229);
nand U1080 (N_1080,N_838,N_646);
and U1081 (N_1081,N_528,In_742);
or U1082 (N_1082,In_2117,N_118);
and U1083 (N_1083,In_1702,In_854);
and U1084 (N_1084,N_190,In_1173);
nor U1085 (N_1085,N_822,In_779);
nor U1086 (N_1086,N_554,N_530);
nor U1087 (N_1087,N_295,N_548);
nor U1088 (N_1088,In_1612,In_2049);
and U1089 (N_1089,N_506,N_550);
and U1090 (N_1090,N_739,N_643);
xnor U1091 (N_1091,N_729,N_701);
xnor U1092 (N_1092,N_709,In_2394);
and U1093 (N_1093,In_2222,In_2220);
or U1094 (N_1094,In_1518,N_956);
xnor U1095 (N_1095,In_166,In_1683);
nand U1096 (N_1096,In_1627,N_675);
or U1097 (N_1097,In_2462,In_161);
or U1098 (N_1098,In_1355,N_227);
or U1099 (N_1099,In_1741,In_1146);
or U1100 (N_1100,N_22,N_953);
or U1101 (N_1101,N_126,In_1794);
nor U1102 (N_1102,N_965,In_1420);
and U1103 (N_1103,N_197,In_486);
and U1104 (N_1104,In_1886,In_1835);
nand U1105 (N_1105,In_1533,In_691);
nand U1106 (N_1106,In_1996,In_1450);
nand U1107 (N_1107,N_501,N_974);
nand U1108 (N_1108,In_1660,N_573);
nor U1109 (N_1109,N_580,In_1307);
xor U1110 (N_1110,In_821,N_601);
xor U1111 (N_1111,In_183,N_500);
or U1112 (N_1112,N_287,In_1098);
or U1113 (N_1113,N_880,In_508);
and U1114 (N_1114,In_2333,In_1553);
nor U1115 (N_1115,In_1900,N_902);
xnor U1116 (N_1116,N_870,N_852);
and U1117 (N_1117,In_1967,In_2304);
nand U1118 (N_1118,N_864,N_703);
or U1119 (N_1119,N_746,In_119);
and U1120 (N_1120,In_1048,In_373);
nand U1121 (N_1121,N_967,N_561);
nor U1122 (N_1122,N_558,N_798);
xnor U1123 (N_1123,N_959,N_136);
and U1124 (N_1124,In_2078,N_45);
xnor U1125 (N_1125,In_148,N_346);
or U1126 (N_1126,N_151,In_2275);
or U1127 (N_1127,In_1687,In_1555);
xor U1128 (N_1128,In_2033,N_809);
nor U1129 (N_1129,In_1221,N_569);
or U1130 (N_1130,N_771,In_2186);
or U1131 (N_1131,N_557,In_2058);
and U1132 (N_1132,N_826,N_178);
xor U1133 (N_1133,N_376,N_630);
or U1134 (N_1134,N_963,In_1012);
and U1135 (N_1135,N_281,In_180);
nand U1136 (N_1136,N_367,N_420);
xor U1137 (N_1137,In_1335,In_2145);
nand U1138 (N_1138,In_167,In_1536);
and U1139 (N_1139,In_268,In_1836);
or U1140 (N_1140,In_526,In_212);
xnor U1141 (N_1141,N_821,N_0);
nor U1142 (N_1142,In_1430,N_225);
nand U1143 (N_1143,In_2279,In_1273);
xor U1144 (N_1144,In_835,N_30);
or U1145 (N_1145,In_1034,In_1451);
nand U1146 (N_1146,N_526,N_930);
and U1147 (N_1147,N_176,N_882);
nand U1148 (N_1148,N_876,In_461);
and U1149 (N_1149,In_2124,N_799);
or U1150 (N_1150,In_2391,In_264);
nor U1151 (N_1151,N_676,N_92);
xor U1152 (N_1152,In_383,In_2192);
and U1153 (N_1153,N_551,In_227);
or U1154 (N_1154,N_641,N_610);
nand U1155 (N_1155,In_1666,N_305);
nand U1156 (N_1156,In_2,In_2343);
nor U1157 (N_1157,N_745,In_515);
nor U1158 (N_1158,In_2016,N_433);
nand U1159 (N_1159,In_1261,In_420);
nand U1160 (N_1160,N_444,In_2363);
and U1161 (N_1161,In_680,In_1761);
or U1162 (N_1162,In_1338,In_1570);
or U1163 (N_1163,N_848,N_764);
or U1164 (N_1164,N_529,In_1601);
xnor U1165 (N_1165,In_1387,N_837);
nand U1166 (N_1166,N_752,N_81);
and U1167 (N_1167,In_2046,N_496);
or U1168 (N_1168,In_600,N_634);
or U1169 (N_1169,N_884,N_145);
nand U1170 (N_1170,N_64,N_896);
xor U1171 (N_1171,In_213,N_278);
nand U1172 (N_1172,N_684,In_2435);
or U1173 (N_1173,N_114,In_1588);
nor U1174 (N_1174,In_1078,In_285);
xnor U1175 (N_1175,In_1955,In_271);
or U1176 (N_1176,N_594,N_432);
nand U1177 (N_1177,N_995,In_1768);
xnor U1178 (N_1178,In_540,In_358);
and U1179 (N_1179,In_2233,N_19);
xor U1180 (N_1180,N_91,N_277);
nor U1181 (N_1181,In_1912,In_134);
or U1182 (N_1182,In_2214,In_2303);
or U1183 (N_1183,N_161,N_270);
or U1184 (N_1184,N_648,In_2464);
nor U1185 (N_1185,In_1675,N_403);
nand U1186 (N_1186,In_2448,N_241);
nand U1187 (N_1187,In_783,N_754);
and U1188 (N_1188,In_1300,In_1922);
or U1189 (N_1189,N_389,N_427);
or U1190 (N_1190,In_169,In_952);
or U1191 (N_1191,N_740,In_632);
or U1192 (N_1192,N_883,In_11);
and U1193 (N_1193,In_228,N_812);
nor U1194 (N_1194,N_658,N_699);
nor U1195 (N_1195,N_1,In_1434);
xor U1196 (N_1196,In_1319,N_914);
or U1197 (N_1197,N_131,In_2251);
and U1198 (N_1198,In_1969,In_545);
or U1199 (N_1199,N_588,N_478);
and U1200 (N_1200,In_1049,N_86);
nand U1201 (N_1201,N_559,N_431);
or U1202 (N_1202,N_414,In_747);
or U1203 (N_1203,In_777,N_306);
or U1204 (N_1204,In_2178,In_1943);
nor U1205 (N_1205,In_683,In_1032);
xor U1206 (N_1206,In_1062,N_198);
nand U1207 (N_1207,N_242,N_846);
xor U1208 (N_1208,In_464,In_597);
or U1209 (N_1209,In_1888,In_476);
xnor U1210 (N_1210,In_2137,N_398);
and U1211 (N_1211,N_979,In_1211);
and U1212 (N_1212,N_572,In_643);
or U1213 (N_1213,In_2269,N_921);
or U1214 (N_1214,N_936,In_1210);
nand U1215 (N_1215,In_911,N_523);
or U1216 (N_1216,In_2382,N_629);
or U1217 (N_1217,N_303,In_466);
and U1218 (N_1218,In_1956,In_1232);
nand U1219 (N_1219,N_917,In_302);
nor U1220 (N_1220,In_469,In_246);
or U1221 (N_1221,In_1562,In_869);
nor U1222 (N_1222,N_696,In_1054);
nor U1223 (N_1223,N_724,N_575);
and U1224 (N_1224,In_506,N_534);
nand U1225 (N_1225,N_311,In_2209);
xnor U1226 (N_1226,N_772,In_1839);
and U1227 (N_1227,N_691,In_551);
and U1228 (N_1228,N_570,In_1456);
or U1229 (N_1229,In_1911,In_1616);
xor U1230 (N_1230,N_874,N_459);
nor U1231 (N_1231,In_1364,N_726);
or U1232 (N_1232,N_116,In_1596);
and U1233 (N_1233,In_294,In_8);
or U1234 (N_1234,In_2194,N_379);
or U1235 (N_1235,N_653,In_955);
nand U1236 (N_1236,N_993,N_705);
and U1237 (N_1237,In_726,N_485);
nand U1238 (N_1238,N_964,N_565);
xor U1239 (N_1239,N_250,In_1088);
xor U1240 (N_1240,N_505,In_528);
xnor U1241 (N_1241,In_1245,N_888);
xnor U1242 (N_1242,In_1305,N_469);
or U1243 (N_1243,In_2198,In_759);
xnor U1244 (N_1244,N_304,N_73);
nand U1245 (N_1245,In_225,In_2075);
or U1246 (N_1246,N_757,N_881);
nor U1247 (N_1247,In_718,In_2062);
xnor U1248 (N_1248,In_1446,In_2197);
nor U1249 (N_1249,In_382,N_215);
xor U1250 (N_1250,In_1251,In_417);
or U1251 (N_1251,In_2478,N_857);
and U1252 (N_1252,In_194,In_74);
nand U1253 (N_1253,N_360,N_144);
or U1254 (N_1254,N_606,N_830);
nand U1255 (N_1255,N_457,N_365);
and U1256 (N_1256,N_678,In_2204);
and U1257 (N_1257,N_424,N_274);
and U1258 (N_1258,In_2159,In_1175);
nand U1259 (N_1259,In_2057,N_996);
or U1260 (N_1260,In_624,N_878);
or U1261 (N_1261,In_1747,In_2264);
nand U1262 (N_1262,In_906,N_808);
or U1263 (N_1263,In_2439,N_828);
and U1264 (N_1264,In_2375,N_804);
and U1265 (N_1265,N_437,In_938);
nand U1266 (N_1266,In_405,N_555);
nor U1267 (N_1267,In_1944,In_2026);
or U1268 (N_1268,N_899,N_732);
and U1269 (N_1269,In_1684,N_825);
nand U1270 (N_1270,N_41,N_927);
nand U1271 (N_1271,In_2134,N_613);
nand U1272 (N_1272,In_483,In_1883);
and U1273 (N_1273,In_2316,N_525);
and U1274 (N_1274,N_911,In_1799);
nand U1275 (N_1275,In_471,N_983);
nand U1276 (N_1276,In_2497,N_807);
xor U1277 (N_1277,In_2215,In_1241);
xor U1278 (N_1278,N_326,In_2459);
nand U1279 (N_1279,N_693,In_2090);
xnor U1280 (N_1280,In_1011,N_681);
xnor U1281 (N_1281,N_520,In_2168);
nand U1282 (N_1282,N_912,In_1205);
xor U1283 (N_1283,In_565,N_847);
xnor U1284 (N_1284,In_2289,N_549);
xnor U1285 (N_1285,N_642,N_325);
or U1286 (N_1286,N_334,In_254);
and U1287 (N_1287,N_182,In_1631);
nor U1288 (N_1288,In_479,N_875);
xnor U1289 (N_1289,In_2202,N_90);
nand U1290 (N_1290,In_2355,N_910);
or U1291 (N_1291,N_908,In_1279);
xnor U1292 (N_1292,In_531,N_950);
and U1293 (N_1293,In_187,N_547);
xor U1294 (N_1294,N_493,N_773);
or U1295 (N_1295,In_728,In_714);
nor U1296 (N_1296,N_783,In_1466);
nand U1297 (N_1297,N_511,N_203);
nand U1298 (N_1298,In_2306,In_1197);
xnor U1299 (N_1299,In_316,N_313);
nand U1300 (N_1300,In_2083,N_173);
xor U1301 (N_1301,N_692,N_524);
and U1302 (N_1302,N_720,In_2281);
and U1303 (N_1303,In_2461,N_795);
nand U1304 (N_1304,In_2404,In_1483);
xor U1305 (N_1305,In_1659,In_1961);
nor U1306 (N_1306,N_961,In_1913);
nand U1307 (N_1307,In_1369,N_937);
and U1308 (N_1308,N_894,In_2263);
xor U1309 (N_1309,In_609,N_871);
nor U1310 (N_1310,In_1852,N_971);
or U1311 (N_1311,In_1618,In_809);
nor U1312 (N_1312,In_1322,In_335);
nand U1313 (N_1313,In_2170,In_1765);
and U1314 (N_1314,N_831,N_574);
or U1315 (N_1315,N_290,In_1303);
and U1316 (N_1316,In_605,In_2452);
nand U1317 (N_1317,In_150,In_211);
and U1318 (N_1318,In_2433,N_784);
xnor U1319 (N_1319,In_143,N_893);
nand U1320 (N_1320,N_928,N_563);
nor U1321 (N_1321,In_2256,In_800);
nand U1322 (N_1322,In_1654,In_866);
and U1323 (N_1323,N_464,In_863);
nand U1324 (N_1324,N_226,In_513);
or U1325 (N_1325,In_2009,N_748);
nand U1326 (N_1326,In_1946,N_527);
or U1327 (N_1327,In_2284,N_532);
nand U1328 (N_1328,In_1185,N_94);
and U1329 (N_1329,N_579,N_999);
xor U1330 (N_1330,In_2469,N_834);
nor U1331 (N_1331,In_984,N_44);
nor U1332 (N_1332,N_915,N_356);
or U1333 (N_1333,In_949,N_111);
xnor U1334 (N_1334,In_2250,N_566);
nand U1335 (N_1335,In_2227,In_566);
nand U1336 (N_1336,In_2353,N_392);
nand U1337 (N_1337,In_1103,In_509);
xnor U1338 (N_1338,In_1501,N_95);
and U1339 (N_1339,In_1869,In_793);
nor U1340 (N_1340,N_635,In_2408);
nor U1341 (N_1341,In_1730,N_909);
and U1342 (N_1342,N_932,N_512);
or U1343 (N_1343,In_607,N_761);
nand U1344 (N_1344,N_986,In_284);
nor U1345 (N_1345,In_1568,N_513);
nand U1346 (N_1346,In_1811,N_514);
or U1347 (N_1347,In_2199,In_1993);
and U1348 (N_1348,N_714,In_1043);
and U1349 (N_1349,N_34,In_1097);
nor U1350 (N_1350,In_1315,N_426);
xor U1351 (N_1351,In_773,N_975);
xnor U1352 (N_1352,In_900,N_651);
nand U1353 (N_1353,N_968,In_2260);
nand U1354 (N_1354,N_568,In_2484);
or U1355 (N_1355,N_952,N_700);
nor U1356 (N_1356,In_839,In_1183);
or U1357 (N_1357,In_2373,In_1129);
and U1358 (N_1358,N_753,N_666);
nor U1359 (N_1359,In_943,N_435);
xor U1360 (N_1360,N_312,N_224);
xnor U1361 (N_1361,N_713,N_531);
and U1362 (N_1362,In_2182,N_667);
and U1363 (N_1363,In_676,In_824);
nor U1364 (N_1364,N_31,In_330);
nand U1365 (N_1365,N_750,In_535);
nor U1366 (N_1366,N_907,N_430);
xor U1367 (N_1367,In_1901,In_1933);
xnor U1368 (N_1368,In_113,N_769);
and U1369 (N_1369,N_712,In_1791);
nand U1370 (N_1370,N_751,In_22);
xor U1371 (N_1371,N_546,N_728);
nand U1372 (N_1372,N_87,In_1584);
nand U1373 (N_1373,In_533,In_1935);
nand U1374 (N_1374,In_1292,In_89);
and U1375 (N_1375,In_1217,N_638);
or U1376 (N_1376,N_607,In_1597);
or U1377 (N_1377,In_313,N_521);
or U1378 (N_1378,N_698,In_1662);
xnor U1379 (N_1379,In_260,N_677);
and U1380 (N_1380,In_1192,In_2374);
or U1381 (N_1381,In_135,In_1543);
or U1382 (N_1382,N_567,In_1890);
and U1383 (N_1383,N_802,N_997);
or U1384 (N_1384,N_817,N_518);
xor U1385 (N_1385,In_1317,In_478);
nor U1386 (N_1386,In_615,In_981);
and U1387 (N_1387,N_850,In_68);
nor U1388 (N_1388,N_543,N_672);
nor U1389 (N_1389,In_1545,N_425);
and U1390 (N_1390,N_502,In_1417);
and U1391 (N_1391,In_1165,N_711);
or U1392 (N_1392,N_704,In_695);
nor U1393 (N_1393,N_650,In_890);
xnor U1394 (N_1394,In_1864,In_944);
xor U1395 (N_1395,In_1174,N_644);
nand U1396 (N_1396,N_286,In_1066);
or U1397 (N_1397,In_1517,In_556);
xor U1398 (N_1398,N_855,N_649);
or U1399 (N_1399,In_2442,N_749);
xnor U1400 (N_1400,In_191,N_742);
and U1401 (N_1401,In_310,N_466);
xor U1402 (N_1402,N_342,N_839);
and U1403 (N_1403,N_440,N_576);
xor U1404 (N_1404,N_879,In_685);
and U1405 (N_1405,In_2224,N_603);
or U1406 (N_1406,In_1717,In_249);
nor U1407 (N_1407,N_522,In_1374);
and U1408 (N_1408,N_2,In_1312);
xnor U1409 (N_1409,In_387,N_686);
and U1410 (N_1410,N_320,N_604);
nor U1411 (N_1411,N_15,In_229);
and U1412 (N_1412,N_823,In_916);
or U1413 (N_1413,In_1377,N_428);
nand U1414 (N_1414,N_661,In_1798);
xor U1415 (N_1415,N_782,N_327);
xnor U1416 (N_1416,N_614,In_2019);
xor U1417 (N_1417,N_6,In_1110);
and U1418 (N_1418,In_1124,In_1410);
and U1419 (N_1419,N_384,N_969);
xnor U1420 (N_1420,N_985,In_1750);
nand U1421 (N_1421,N_889,N_988);
and U1422 (N_1422,N_940,In_1017);
or U1423 (N_1423,In_1177,N_887);
xor U1424 (N_1424,N_656,N_719);
or U1425 (N_1425,In_499,N_590);
nand U1426 (N_1426,In_240,N_824);
and U1427 (N_1427,In_1170,In_1280);
or U1428 (N_1428,In_1491,In_1620);
xnor U1429 (N_1429,N_533,In_1789);
and U1430 (N_1430,In_152,In_269);
nand U1431 (N_1431,In_2322,N_394);
and U1432 (N_1432,N_958,N_619);
nand U1433 (N_1433,N_149,N_925);
xor U1434 (N_1434,N_331,In_2377);
nand U1435 (N_1435,N_939,N_289);
or U1436 (N_1436,N_443,In_132);
and U1437 (N_1437,N_404,In_79);
nand U1438 (N_1438,In_14,In_1242);
nor U1439 (N_1439,N_616,In_1507);
xor U1440 (N_1440,N_886,In_1325);
and U1441 (N_1441,N_982,In_965);
nand U1442 (N_1442,N_447,In_391);
nand U1443 (N_1443,In_519,In_823);
nor U1444 (N_1444,In_635,N_835);
xor U1445 (N_1445,In_645,N_597);
and U1446 (N_1446,In_2061,N_595);
nand U1447 (N_1447,In_992,In_536);
nor U1448 (N_1448,N_228,N_621);
nand U1449 (N_1449,In_674,In_255);
nor U1450 (N_1450,N_890,N_647);
and U1451 (N_1451,N_103,In_2175);
xnor U1452 (N_1452,In_778,In_323);
nand U1453 (N_1453,In_669,In_2015);
or U1454 (N_1454,N_976,In_977);
and U1455 (N_1455,In_216,N_866);
and U1456 (N_1456,In_397,In_2490);
nor U1457 (N_1457,In_1367,In_630);
nor U1458 (N_1458,In_2084,In_1582);
nor U1459 (N_1459,N_920,N_625);
and U1460 (N_1460,In_1520,N_344);
nor U1461 (N_1461,N_918,N_636);
nand U1462 (N_1462,In_2389,N_683);
and U1463 (N_1463,N_65,In_2173);
xor U1464 (N_1464,In_121,N_545);
xor U1465 (N_1465,In_2280,N_663);
and U1466 (N_1466,In_149,N_366);
nand U1467 (N_1467,N_322,N_763);
nand U1468 (N_1468,N_377,N_504);
and U1469 (N_1469,In_1477,In_1361);
xnor U1470 (N_1470,In_2456,N_670);
xor U1471 (N_1471,N_387,N_96);
nand U1472 (N_1472,In_799,N_906);
xnor U1473 (N_1473,N_135,In_244);
nand U1474 (N_1474,N_347,N_853);
xnor U1475 (N_1475,In_1188,In_1453);
xnor U1476 (N_1476,In_30,N_765);
or U1477 (N_1477,N_139,In_2413);
or U1478 (N_1478,In_2187,In_1180);
nand U1479 (N_1479,In_2125,N_797);
nor U1480 (N_1480,In_1473,In_1726);
or U1481 (N_1481,N_282,N_129);
xor U1482 (N_1482,In_1432,In_282);
nor U1483 (N_1483,In_1965,N_238);
and U1484 (N_1484,In_128,In_1797);
or U1485 (N_1485,In_1551,N_353);
and U1486 (N_1486,In_1309,N_891);
nand U1487 (N_1487,In_833,In_1550);
nand U1488 (N_1488,N_503,N_189);
nor U1489 (N_1489,In_2332,In_1861);
nand U1490 (N_1490,In_1628,N_36);
or U1491 (N_1491,In_353,N_645);
nand U1492 (N_1492,N_738,In_1469);
nand U1493 (N_1493,N_662,In_2002);
nand U1494 (N_1494,In_393,N_652);
nand U1495 (N_1495,N_951,In_1358);
nor U1496 (N_1496,In_590,In_3);
nand U1497 (N_1497,In_2310,N_17);
xor U1498 (N_1498,In_1127,N_723);
nand U1499 (N_1499,N_990,N_929);
or U1500 (N_1500,N_181,N_364);
xor U1501 (N_1501,In_473,N_1098);
and U1502 (N_1502,N_1142,In_2271);
and U1503 (N_1503,N_972,In_1448);
or U1504 (N_1504,In_2067,In_1746);
or U1505 (N_1505,In_210,N_1389);
xor U1506 (N_1506,N_1318,N_1314);
and U1507 (N_1507,N_935,In_2207);
or U1508 (N_1508,N_1008,N_1072);
nand U1509 (N_1509,N_1446,In_853);
nand U1510 (N_1510,N_1205,N_1157);
xor U1511 (N_1511,In_1449,N_1050);
nand U1512 (N_1512,N_1384,N_1092);
nand U1513 (N_1513,N_780,N_1221);
or U1514 (N_1514,In_340,In_2162);
xor U1515 (N_1515,In_443,N_781);
nor U1516 (N_1516,N_1174,N_1197);
or U1517 (N_1517,N_1159,N_1320);
xor U1518 (N_1518,N_1045,N_845);
nor U1519 (N_1519,N_1278,In_2425);
nor U1520 (N_1520,N_47,N_67);
xor U1521 (N_1521,N_1160,N_1224);
or U1522 (N_1522,N_454,N_1448);
xor U1523 (N_1523,N_1262,In_1428);
nand U1524 (N_1524,In_2470,N_1149);
nor U1525 (N_1525,In_724,N_1071);
xor U1526 (N_1526,N_948,N_892);
and U1527 (N_1527,N_1091,N_1207);
nand U1528 (N_1528,N_1427,N_1288);
and U1529 (N_1529,N_735,N_1196);
or U1530 (N_1530,N_1173,N_210);
nor U1531 (N_1531,N_1139,In_1866);
nor U1532 (N_1532,N_1260,In_530);
xnor U1533 (N_1533,In_577,N_1246);
and U1534 (N_1534,N_1300,N_1078);
nand U1535 (N_1535,N_1307,In_864);
nand U1536 (N_1536,N_1478,N_957);
nor U1537 (N_1537,N_1015,In_4);
and U1538 (N_1538,In_1061,N_1476);
nor U1539 (N_1539,In_716,N_1390);
xnor U1540 (N_1540,N_1394,N_868);
xnor U1541 (N_1541,N_11,N_1352);
xnor U1542 (N_1542,N_843,N_944);
nor U1543 (N_1543,N_1035,In_1426);
nor U1544 (N_1544,In_1390,In_698);
nor U1545 (N_1545,N_1374,In_738);
xor U1546 (N_1546,N_1455,N_1415);
or U1547 (N_1547,N_1214,N_562);
or U1548 (N_1548,N_1003,N_1203);
or U1549 (N_1549,N_1188,In_2337);
or U1550 (N_1550,N_1379,N_820);
nor U1551 (N_1551,N_1162,N_924);
xnor U1552 (N_1552,N_253,N_1313);
nor U1553 (N_1553,In_830,In_579);
or U1554 (N_1554,N_1106,N_1341);
and U1555 (N_1555,N_1178,N_1402);
or U1556 (N_1556,N_1412,N_1466);
nor U1557 (N_1557,In_1642,N_159);
nor U1558 (N_1558,In_1837,N_1047);
xor U1559 (N_1559,N_1470,N_1021);
nand U1560 (N_1560,N_1070,N_1373);
or U1561 (N_1561,N_1344,N_1225);
xor U1562 (N_1562,In_1158,In_1090);
nor U1563 (N_1563,N_1122,N_1444);
nand U1564 (N_1564,N_1428,N_980);
or U1565 (N_1565,N_1425,N_117);
nor U1566 (N_1566,N_1116,N_1193);
or U1567 (N_1567,N_1132,N_707);
nand U1568 (N_1568,N_1356,N_245);
and U1569 (N_1569,N_1258,N_919);
or U1570 (N_1570,N_1283,N_1234);
nand U1571 (N_1571,N_1458,In_61);
nand U1572 (N_1572,In_1916,N_1451);
nand U1573 (N_1573,N_862,N_1292);
nor U1574 (N_1574,N_1083,N_1460);
or U1575 (N_1575,In_785,In_1028);
nand U1576 (N_1576,In_1928,In_2050);
or U1577 (N_1577,N_1365,In_245);
and U1578 (N_1578,N_1269,N_818);
and U1579 (N_1579,N_539,N_509);
nor U1580 (N_1580,N_1492,N_665);
nor U1581 (N_1581,In_1334,In_196);
xnor U1582 (N_1582,N_1311,N_1326);
nor U1583 (N_1583,N_655,N_1378);
nand U1584 (N_1584,N_1324,N_885);
xnor U1585 (N_1585,N_1275,In_557);
xor U1586 (N_1586,N_1038,N_1317);
nor U1587 (N_1587,In_498,In_2077);
nand U1588 (N_1588,N_1184,N_1377);
nand U1589 (N_1589,N_1380,In_1638);
xor U1590 (N_1590,In_367,N_1481);
nor U1591 (N_1591,N_1084,In_1581);
or U1592 (N_1592,N_587,N_1349);
or U1593 (N_1593,In_2292,In_1328);
nand U1594 (N_1594,N_1241,N_1357);
and U1595 (N_1595,N_593,N_775);
or U1596 (N_1596,N_1371,N_1163);
or U1597 (N_1597,In_1438,N_1218);
or U1598 (N_1598,In_2499,N_298);
nor U1599 (N_1599,N_1034,In_1782);
and U1600 (N_1600,N_1299,In_1418);
or U1601 (N_1601,In_1351,N_1302);
nand U1602 (N_1602,N_611,In_586);
nor U1603 (N_1603,N_552,N_624);
nor U1604 (N_1604,N_1490,N_1494);
or U1605 (N_1605,N_1382,N_1175);
xor U1606 (N_1606,In_514,N_1147);
and U1607 (N_1607,N_35,N_1226);
nand U1608 (N_1608,N_1325,N_800);
and U1609 (N_1609,In_1647,N_596);
and U1610 (N_1610,In_851,N_1407);
and U1611 (N_1611,N_1279,N_1102);
or U1612 (N_1612,N_378,N_1245);
and U1613 (N_1613,N_1354,N_196);
nand U1614 (N_1614,N_1426,N_1027);
nor U1615 (N_1615,N_586,N_1040);
nand U1616 (N_1616,N_1408,N_1335);
and U1617 (N_1617,N_592,N_947);
xor U1618 (N_1618,N_1136,N_1169);
xor U1619 (N_1619,N_260,N_861);
xor U1620 (N_1620,In_594,In_181);
nand U1621 (N_1621,N_706,N_1396);
xor U1622 (N_1622,N_1247,N_1222);
nor U1623 (N_1623,N_811,N_1110);
nor U1624 (N_1624,N_819,In_2318);
and U1625 (N_1625,N_1154,N_368);
or U1626 (N_1626,N_109,N_731);
xnor U1627 (N_1627,In_1808,In_2031);
and U1628 (N_1628,In_1825,N_138);
or U1629 (N_1629,N_792,N_734);
nand U1630 (N_1630,N_1430,N_659);
xor U1631 (N_1631,N_1235,N_1489);
nor U1632 (N_1632,In_1621,N_992);
xor U1633 (N_1633,N_1243,N_973);
xor U1634 (N_1634,N_1453,N_1057);
nor U1635 (N_1635,In_1772,In_2308);
and U1636 (N_1636,In_511,N_494);
nand U1637 (N_1637,N_544,In_1587);
xnor U1638 (N_1638,In_1831,N_872);
or U1639 (N_1639,N_405,N_1381);
or U1640 (N_1640,N_1165,N_1310);
or U1641 (N_1641,N_599,N_727);
nand U1642 (N_1642,N_1473,N_863);
and U1643 (N_1643,N_1145,In_2376);
or U1644 (N_1644,In_415,N_262);
nor U1645 (N_1645,N_1082,In_1178);
xnor U1646 (N_1646,N_229,N_1437);
or U1647 (N_1647,N_1210,N_1264);
nand U1648 (N_1648,N_1066,N_1308);
nand U1649 (N_1649,In_333,N_1353);
nand U1650 (N_1650,In_2193,N_756);
nand U1651 (N_1651,N_1261,In_1147);
nand U1652 (N_1652,N_1461,N_1309);
xnor U1653 (N_1653,N_1231,N_1398);
or U1654 (N_1654,N_488,N_1181);
xnor U1655 (N_1655,N_689,In_1244);
nand U1656 (N_1656,N_240,N_791);
xnor U1657 (N_1657,N_1167,In_703);
or U1658 (N_1658,N_1331,N_1158);
and U1659 (N_1659,N_628,N_1445);
xnor U1660 (N_1660,N_1011,In_338);
nand U1661 (N_1661,N_1041,In_487);
nand U1662 (N_1662,N_721,N_223);
nor U1663 (N_1663,In_1667,N_1340);
nand U1664 (N_1664,In_642,N_370);
and U1665 (N_1665,N_1467,N_744);
or U1666 (N_1666,N_1447,N_933);
or U1667 (N_1667,N_1395,N_423);
nand U1668 (N_1668,N_945,N_1002);
or U1669 (N_1669,In_1822,N_540);
or U1670 (N_1670,N_1315,N_1183);
and U1671 (N_1671,N_1401,N_1345);
or U1672 (N_1672,N_1074,N_1417);
xnor U1673 (N_1673,N_1495,N_1272);
and U1674 (N_1674,N_165,N_1252);
xor U1675 (N_1675,N_1423,N_1176);
and U1676 (N_1676,N_1161,N_934);
nand U1677 (N_1677,N_1255,N_1126);
and U1678 (N_1678,N_984,In_750);
nor U1679 (N_1679,In_856,N_1383);
nand U1680 (N_1680,In_10,In_2080);
nand U1681 (N_1681,In_2060,N_1334);
nand U1682 (N_1682,N_743,In_370);
nor U1683 (N_1683,N_1130,N_620);
nand U1684 (N_1684,N_796,N_1124);
nor U1685 (N_1685,N_787,N_688);
xor U1686 (N_1686,N_193,N_1404);
xnor U1687 (N_1687,In_638,In_623);
nor U1688 (N_1688,N_600,N_1268);
and U1689 (N_1689,N_1464,N_1485);
or U1690 (N_1690,In_1333,N_730);
nand U1691 (N_1691,In_2406,N_1433);
nor U1692 (N_1692,In_1176,N_829);
nand U1693 (N_1693,N_1032,N_462);
nand U1694 (N_1694,N_1164,N_942);
nor U1695 (N_1695,N_602,In_1736);
or U1696 (N_1696,N_844,N_9);
and U1697 (N_1697,N_981,N_1118);
nor U1698 (N_1698,N_1025,In_2104);
or U1699 (N_1699,N_1266,N_1399);
xor U1700 (N_1700,N_1179,In_261);
and U1701 (N_1701,N_1097,N_851);
or U1702 (N_1702,In_969,N_1351);
xnor U1703 (N_1703,N_673,N_1350);
and U1704 (N_1704,In_1899,N_1304);
xnor U1705 (N_1705,N_170,N_1217);
nor U1706 (N_1706,In_2045,N_790);
or U1707 (N_1707,N_998,N_1128);
and U1708 (N_1708,N_1244,N_453);
and U1709 (N_1709,N_626,In_1125);
xnor U1710 (N_1710,N_637,N_690);
nand U1711 (N_1711,N_1228,In_538);
or U1712 (N_1712,N_1434,N_1387);
or U1713 (N_1713,In_407,N_1199);
nor U1714 (N_1714,N_1232,N_1085);
xnor U1715 (N_1715,N_1194,N_1290);
nor U1716 (N_1716,N_207,In_574);
nand U1717 (N_1717,N_24,N_1296);
or U1718 (N_1718,N_1479,N_1219);
or U1719 (N_1719,N_1409,N_46);
xnor U1720 (N_1720,N_1029,In_236);
xnor U1721 (N_1721,N_1018,N_479);
xor U1722 (N_1722,N_1172,In_2258);
or U1723 (N_1723,N_1020,In_1160);
nor U1724 (N_1724,N_1348,N_1198);
nor U1725 (N_1725,In_2267,In_1523);
and U1726 (N_1726,In_481,N_622);
xnor U1727 (N_1727,N_741,N_1431);
nor U1728 (N_1728,N_1212,N_1223);
nor U1729 (N_1729,N_1363,N_1462);
or U1730 (N_1730,N_1477,N_495);
or U1731 (N_1731,N_970,N_904);
and U1732 (N_1732,In_1889,In_591);
or U1733 (N_1733,N_542,N_1497);
xnor U1734 (N_1734,N_1282,N_589);
or U1735 (N_1735,N_1090,In_1400);
nand U1736 (N_1736,N_1347,N_1120);
nand U1737 (N_1737,In_752,In_589);
nor U1738 (N_1738,In_1005,In_1792);
and U1739 (N_1739,In_1404,N_1043);
or U1740 (N_1740,N_1364,N_1216);
or U1741 (N_1741,N_1251,N_1010);
or U1742 (N_1742,N_3,In_71);
xnor U1743 (N_1743,N_1143,N_1422);
nor U1744 (N_1744,In_342,In_458);
nor U1745 (N_1745,In_50,N_1405);
nand U1746 (N_1746,N_905,N_841);
and U1747 (N_1747,N_1359,In_1934);
nor U1748 (N_1748,In_232,N_1483);
or U1749 (N_1749,N_1094,N_237);
or U1750 (N_1750,In_84,N_1254);
or U1751 (N_1751,N_1281,N_1285);
and U1752 (N_1752,N_1185,In_1539);
nand U1753 (N_1753,In_1044,N_1328);
or U1754 (N_1754,N_553,N_324);
xnor U1755 (N_1755,N_108,In_2265);
nor U1756 (N_1756,N_1248,N_1019);
xor U1757 (N_1757,In_880,N_955);
nand U1758 (N_1758,N_1026,N_480);
nand U1759 (N_1759,N_1441,N_1330);
nor U1760 (N_1760,In_1009,In_1089);
nor U1761 (N_1761,N_766,N_1442);
xor U1762 (N_1762,N_669,N_42);
nor U1763 (N_1763,In_1445,N_1037);
nor U1764 (N_1764,In_266,N_1095);
or U1765 (N_1765,N_401,N_1491);
xnor U1766 (N_1766,N_1321,N_1493);
and U1767 (N_1767,N_901,N_1187);
nor U1768 (N_1768,N_941,In_1983);
nor U1769 (N_1769,N_265,N_1306);
or U1770 (N_1770,N_768,N_873);
nand U1771 (N_1771,In_474,In_2488);
xor U1772 (N_1772,N_1170,N_633);
or U1773 (N_1773,N_814,N_1171);
nor U1774 (N_1774,N_1312,In_1585);
xnor U1775 (N_1775,N_1443,N_1141);
nand U1776 (N_1776,N_1293,In_1851);
xor U1777 (N_1777,N_1305,N_355);
or U1778 (N_1778,N_507,N_1406);
and U1779 (N_1779,N_1230,N_1099);
nor U1780 (N_1780,N_1146,N_1286);
nor U1781 (N_1781,N_1284,N_1229);
nor U1782 (N_1782,N_1468,N_571);
xor U1783 (N_1783,N_1294,In_2238);
and U1784 (N_1784,N_1209,N_373);
nor U1785 (N_1785,In_1530,N_1061);
xnor U1786 (N_1786,In_2270,In_1766);
and U1787 (N_1787,N_1257,In_602);
or U1788 (N_1788,N_1112,In_207);
and U1789 (N_1789,N_759,N_1182);
nor U1790 (N_1790,N_1004,In_2226);
xor U1791 (N_1791,N_292,N_1088);
nand U1792 (N_1792,N_816,N_1459);
and U1793 (N_1793,N_1432,In_757);
nor U1794 (N_1794,N_827,N_1051);
or U1795 (N_1795,N_1280,N_8);
nor U1796 (N_1796,N_1397,In_2001);
xnor U1797 (N_1797,N_664,In_894);
nor U1798 (N_1798,N_1265,In_1929);
nand U1799 (N_1799,N_1113,N_895);
nor U1800 (N_1800,In_554,N_1463);
nand U1801 (N_1801,N_777,N_1342);
xnor U1802 (N_1802,N_1457,N_1189);
or U1803 (N_1803,In_2466,N_560);
nor U1804 (N_1804,In_92,N_1054);
and U1805 (N_1805,N_1213,N_1336);
xor U1806 (N_1806,N_1093,In_956);
and U1807 (N_1807,In_1813,In_929);
xor U1808 (N_1808,In_1607,N_1469);
nand U1809 (N_1809,N_18,N_1206);
xnor U1810 (N_1810,N_755,In_1732);
or U1811 (N_1811,N_1303,N_618);
xnor U1812 (N_1812,N_1127,N_1067);
xor U1813 (N_1813,In_1031,In_1893);
nor U1814 (N_1814,N_1227,N_1263);
and U1815 (N_1815,N_1023,N_1101);
and U1816 (N_1816,In_654,N_1480);
nand U1817 (N_1817,N_682,In_1991);
or U1818 (N_1818,N_1086,N_708);
or U1819 (N_1819,N_1115,In_644);
xor U1820 (N_1820,N_1100,N_1316);
nor U1821 (N_1821,N_1376,N_112);
nand U1822 (N_1822,N_657,N_1073);
or U1823 (N_1823,N_556,N_1372);
nand U1824 (N_1824,N_1056,N_1276);
xnor U1825 (N_1825,N_585,N_1488);
nand U1826 (N_1826,N_175,In_756);
or U1827 (N_1827,N_1475,In_1796);
xnor U1828 (N_1828,N_1104,N_1028);
nand U1829 (N_1829,N_806,N_1343);
or U1830 (N_1830,N_1007,N_1044);
nor U1831 (N_1831,N_1200,N_79);
and U1832 (N_1832,In_2426,N_1013);
nor U1833 (N_1833,N_1392,In_2042);
or U1834 (N_1834,N_1456,N_1339);
and U1835 (N_1835,N_1062,N_1080);
and U1836 (N_1836,N_1250,N_1220);
and U1837 (N_1837,N_1411,In_1829);
xor U1838 (N_1838,N_1081,N_1117);
and U1839 (N_1839,In_452,N_1273);
nor U1840 (N_1840,In_723,N_1487);
xnor U1841 (N_1841,N_1153,N_923);
nand U1842 (N_1842,N_715,N_1060);
nor U1843 (N_1843,N_1429,N_725);
or U1844 (N_1844,N_1418,N_515);
nor U1845 (N_1845,In_7,In_292);
nand U1846 (N_1846,N_1360,In_1030);
nand U1847 (N_1847,In_1222,N_786);
nand U1848 (N_1848,N_354,In_1246);
or U1849 (N_1849,N_578,N_1063);
or U1850 (N_1850,N_1177,N_1289);
nand U1851 (N_1851,In_2365,N_452);
or U1852 (N_1852,N_1119,N_1096);
or U1853 (N_1853,N_1048,N_1240);
and U1854 (N_1854,N_978,N_1253);
nor U1855 (N_1855,In_1793,In_111);
xor U1856 (N_1856,In_711,N_1486);
nor U1857 (N_1857,N_1059,N_832);
xnor U1858 (N_1858,N_1400,N_1366);
and U1859 (N_1859,In_460,N_762);
xnor U1860 (N_1860,N_966,N_184);
or U1861 (N_1861,N_1482,N_204);
xor U1862 (N_1862,N_1420,N_1068);
and U1863 (N_1863,In_337,N_21);
nand U1864 (N_1864,N_1454,N_1065);
xnor U1865 (N_1865,N_685,N_1271);
nor U1866 (N_1866,N_1155,N_1109);
or U1867 (N_1867,In_1256,N_1256);
nor U1868 (N_1868,N_1075,N_1024);
nor U1869 (N_1869,In_1699,N_1237);
and U1870 (N_1870,N_1036,N_608);
or U1871 (N_1871,N_1180,N_508);
nand U1872 (N_1872,In_173,N_1016);
xnor U1873 (N_1873,N_1355,In_2431);
or U1874 (N_1874,In_867,N_1440);
xnor U1875 (N_1875,N_1295,In_1384);
and U1876 (N_1876,N_859,N_584);
xnor U1877 (N_1877,In_1379,N_1166);
and U1878 (N_1878,N_788,N_1009);
and U1879 (N_1879,N_445,N_1439);
nor U1880 (N_1880,In_16,N_1017);
nor U1881 (N_1881,N_1416,In_2336);
and U1882 (N_1882,N_1137,In_2423);
or U1883 (N_1883,N_1049,N_254);
nand U1884 (N_1884,N_1211,In_1425);
and U1885 (N_1885,N_1208,N_244);
or U1886 (N_1886,N_858,N_1069);
or U1887 (N_1887,N_5,N_1287);
and U1888 (N_1888,N_1393,In_419);
xor U1889 (N_1889,In_276,N_1403);
or U1890 (N_1890,N_717,N_1332);
nand U1891 (N_1891,N_1323,N_1298);
nand U1892 (N_1892,N_674,N_836);
nand U1893 (N_1893,N_1267,N_1001);
and U1894 (N_1894,In_223,N_1484);
xnor U1895 (N_1895,N_1438,N_1386);
nand U1896 (N_1896,N_639,N_1192);
and U1897 (N_1897,N_1076,N_849);
nand U1898 (N_1898,In_1224,N_232);
nor U1899 (N_1899,N_1055,N_1135);
or U1900 (N_1900,In_857,N_1151);
and U1901 (N_1901,N_660,N_1498);
or U1902 (N_1902,N_916,N_1046);
or U1903 (N_1903,N_1125,In_1385);
nor U1904 (N_1904,N_537,N_1152);
nor U1905 (N_1905,N_489,N_1000);
nand U1906 (N_1906,N_1033,N_903);
nor U1907 (N_1907,N_1089,N_1058);
nand U1908 (N_1908,In_1535,N_702);
nand U1909 (N_1909,N_1005,N_1087);
nor U1910 (N_1910,N_949,N_1201);
or U1911 (N_1911,In_1052,N_1413);
nand U1912 (N_1912,N_778,N_860);
nor U1913 (N_1913,In_1378,N_406);
nand U1914 (N_1914,N_615,N_1322);
or U1915 (N_1915,N_1014,N_1238);
and U1916 (N_1916,N_1449,In_357);
xnor U1917 (N_1917,N_1133,N_960);
or U1918 (N_1918,In_347,N_1435);
xor U1919 (N_1919,N_1111,In_504);
nand U1920 (N_1920,N_85,N_612);
nor U1921 (N_1921,N_1259,N_900);
nor U1922 (N_1922,N_1358,N_1421);
nand U1923 (N_1923,N_1236,N_536);
nor U1924 (N_1924,N_192,N_1370);
and U1925 (N_1925,N_492,N_1419);
or U1926 (N_1926,N_294,N_1140);
xor U1927 (N_1927,N_1202,In_858);
nor U1928 (N_1928,N_124,N_1131);
xor U1929 (N_1929,N_1052,N_1436);
or U1930 (N_1930,In_1590,In_883);
xnor U1931 (N_1931,N_1297,N_869);
and U1932 (N_1932,N_1301,N_1114);
and U1933 (N_1933,N_483,N_1150);
or U1934 (N_1934,N_1123,N_1053);
nor U1935 (N_1935,N_499,N_987);
or U1936 (N_1936,In_2252,N_315);
xnor U1937 (N_1937,N_1190,N_455);
and U1938 (N_1938,In_470,N_1242);
nand U1939 (N_1939,N_1148,N_913);
and U1940 (N_1940,N_760,N_1368);
nand U1941 (N_1941,N_1333,N_1144);
nor U1942 (N_1942,N_668,N_1012);
nand U1943 (N_1943,N_1042,In_205);
nor U1944 (N_1944,N_1414,N_1105);
and U1945 (N_1945,N_1362,N_1450);
nand U1946 (N_1946,N_694,N_591);
nand U1947 (N_1947,In_2417,In_480);
xor U1948 (N_1948,N_1274,N_854);
nand U1949 (N_1949,In_1594,N_1103);
nand U1950 (N_1950,N_1107,N_1006);
and U1951 (N_1951,N_785,N_1239);
nand U1952 (N_1952,N_1195,In_1320);
xor U1953 (N_1953,N_577,N_1338);
xor U1954 (N_1954,In_1047,N_1156);
nor U1955 (N_1955,N_1329,N_1121);
and U1956 (N_1956,N_1079,N_938);
nor U1957 (N_1957,In_1357,N_946);
nand U1958 (N_1958,N_1499,N_1367);
or U1959 (N_1959,N_1291,N_1375);
nor U1960 (N_1960,N_1249,In_539);
nor U1961 (N_1961,N_541,N_1391);
nand U1962 (N_1962,In_1202,In_1735);
or U1963 (N_1963,N_1204,In_666);
nand U1964 (N_1964,In_501,In_1567);
and U1965 (N_1965,N_1388,In_710);
nand U1966 (N_1966,N_1031,N_1108);
and U1967 (N_1967,N_351,N_926);
nand U1968 (N_1968,N_1134,N_977);
nand U1969 (N_1969,N_1233,In_637);
nor U1970 (N_1970,N_623,N_710);
and U1971 (N_1971,N_789,N_583);
nor U1972 (N_1972,N_1465,N_1030);
or U1973 (N_1973,N_815,N_1191);
or U1974 (N_1974,N_1337,N_458);
or U1975 (N_1975,In_1884,N_1129);
xnor U1976 (N_1976,In_2024,N_1077);
and U1977 (N_1977,N_803,N_1369);
and U1978 (N_1978,N_1471,N_1361);
or U1979 (N_1979,N_722,N_1410);
xor U1980 (N_1980,N_1385,N_856);
and U1981 (N_1981,N_1277,N_810);
nor U1982 (N_1982,N_1496,N_1424);
nor U1983 (N_1983,In_300,In_1391);
and U1984 (N_1984,N_1472,In_36);
and U1985 (N_1985,N_582,In_1500);
nor U1986 (N_1986,In_653,N_1319);
and U1987 (N_1987,N_767,N_436);
nand U1988 (N_1988,N_1186,In_1373);
nand U1989 (N_1989,In_1105,N_467);
xnor U1990 (N_1990,N_631,N_1022);
or U1991 (N_1991,N_510,N_1346);
nor U1992 (N_1992,N_1474,In_288);
nor U1993 (N_1993,N_1215,In_1710);
xor U1994 (N_1994,In_1485,N_989);
xor U1995 (N_1995,N_1168,N_1138);
and U1996 (N_1996,N_779,N_1452);
or U1997 (N_1997,N_1064,N_1327);
or U1998 (N_1998,N_1039,In_2048);
xor U1999 (N_1999,N_1270,In_1354);
or U2000 (N_2000,N_1629,N_1914);
or U2001 (N_2001,N_1608,N_1678);
and U2002 (N_2002,N_1984,N_1665);
nand U2003 (N_2003,N_1863,N_1601);
or U2004 (N_2004,N_1825,N_1876);
nor U2005 (N_2005,N_1642,N_1945);
nor U2006 (N_2006,N_1892,N_1756);
and U2007 (N_2007,N_1571,N_1508);
and U2008 (N_2008,N_1729,N_1619);
nor U2009 (N_2009,N_1784,N_1819);
nand U2010 (N_2010,N_1765,N_1920);
nor U2011 (N_2011,N_1919,N_1744);
and U2012 (N_2012,N_1823,N_1746);
or U2013 (N_2013,N_1593,N_1523);
nand U2014 (N_2014,N_1858,N_1921);
nor U2015 (N_2015,N_1805,N_1961);
and U2016 (N_2016,N_1649,N_1627);
and U2017 (N_2017,N_1993,N_1607);
nand U2018 (N_2018,N_1834,N_1621);
nor U2019 (N_2019,N_1562,N_1987);
and U2020 (N_2020,N_1950,N_1506);
xnor U2021 (N_2021,N_1997,N_1618);
or U2022 (N_2022,N_1926,N_1934);
nor U2023 (N_2023,N_1998,N_1887);
nand U2024 (N_2024,N_1543,N_1898);
xnor U2025 (N_2025,N_1874,N_1894);
nand U2026 (N_2026,N_1771,N_1534);
nand U2027 (N_2027,N_1776,N_1962);
or U2028 (N_2028,N_1943,N_1766);
or U2029 (N_2029,N_1809,N_1503);
xnor U2030 (N_2030,N_1884,N_1905);
nor U2031 (N_2031,N_1636,N_1970);
or U2032 (N_2032,N_1868,N_1720);
or U2033 (N_2033,N_1605,N_1676);
xor U2034 (N_2034,N_1994,N_1718);
nor U2035 (N_2035,N_1979,N_1925);
nor U2036 (N_2036,N_1846,N_1947);
and U2037 (N_2037,N_1739,N_1515);
and U2038 (N_2038,N_1668,N_1799);
xor U2039 (N_2039,N_1745,N_1963);
and U2040 (N_2040,N_1566,N_1606);
xnor U2041 (N_2041,N_1680,N_1500);
nand U2042 (N_2042,N_1779,N_1587);
or U2043 (N_2043,N_1575,N_1933);
nand U2044 (N_2044,N_1940,N_1581);
and U2045 (N_2045,N_1999,N_1527);
or U2046 (N_2046,N_1883,N_1710);
nand U2047 (N_2047,N_1688,N_1693);
xnor U2048 (N_2048,N_1661,N_1567);
or U2049 (N_2049,N_1888,N_1531);
nand U2050 (N_2050,N_1599,N_1808);
nor U2051 (N_2051,N_1501,N_1760);
or U2052 (N_2052,N_1553,N_1786);
nand U2053 (N_2053,N_1681,N_1773);
xnor U2054 (N_2054,N_1740,N_1836);
nand U2055 (N_2055,N_1737,N_1651);
and U2056 (N_2056,N_1980,N_1707);
xor U2057 (N_2057,N_1936,N_1517);
or U2058 (N_2058,N_1538,N_1570);
and U2059 (N_2059,N_1832,N_1859);
and U2060 (N_2060,N_1758,N_1817);
xnor U2061 (N_2061,N_1948,N_1613);
and U2062 (N_2062,N_1754,N_1939);
nand U2063 (N_2063,N_1528,N_1828);
or U2064 (N_2064,N_1841,N_1896);
and U2065 (N_2065,N_1937,N_1670);
nand U2066 (N_2066,N_1848,N_1816);
nor U2067 (N_2067,N_1644,N_1991);
or U2068 (N_2068,N_1713,N_1731);
or U2069 (N_2069,N_1938,N_1869);
xor U2070 (N_2070,N_1787,N_1639);
or U2071 (N_2071,N_1510,N_1540);
nor U2072 (N_2072,N_1781,N_1549);
or U2073 (N_2073,N_1864,N_1539);
or U2074 (N_2074,N_1647,N_1769);
xnor U2075 (N_2075,N_1958,N_1954);
nor U2076 (N_2076,N_1922,N_1723);
nand U2077 (N_2077,N_1717,N_1721);
xnor U2078 (N_2078,N_1546,N_1525);
nand U2079 (N_2079,N_1986,N_1861);
nand U2080 (N_2080,N_1638,N_1658);
and U2081 (N_2081,N_1985,N_1989);
xor U2082 (N_2082,N_1885,N_1568);
nor U2083 (N_2083,N_1911,N_1694);
or U2084 (N_2084,N_1547,N_1951);
nand U2085 (N_2085,N_1873,N_1632);
nand U2086 (N_2086,N_1650,N_1524);
and U2087 (N_2087,N_1502,N_1901);
nand U2088 (N_2088,N_1519,N_1573);
xnor U2089 (N_2089,N_1886,N_1747);
and U2090 (N_2090,N_1923,N_1611);
nor U2091 (N_2091,N_1663,N_1625);
xnor U2092 (N_2092,N_1586,N_1903);
nor U2093 (N_2093,N_1514,N_1851);
or U2094 (N_2094,N_1821,N_1910);
nor U2095 (N_2095,N_1709,N_1912);
xor U2096 (N_2096,N_1978,N_1685);
xnor U2097 (N_2097,N_1576,N_1704);
xor U2098 (N_2098,N_1700,N_1855);
nand U2099 (N_2099,N_1603,N_1695);
xor U2100 (N_2100,N_1879,N_1957);
nand U2101 (N_2101,N_1965,N_1830);
nand U2102 (N_2102,N_1541,N_1730);
or U2103 (N_2103,N_1862,N_1792);
xor U2104 (N_2104,N_1992,N_1902);
and U2105 (N_2105,N_1907,N_1774);
nand U2106 (N_2106,N_1634,N_1529);
xnor U2107 (N_2107,N_1913,N_1533);
nand U2108 (N_2108,N_1722,N_1866);
xor U2109 (N_2109,N_1666,N_1964);
xor U2110 (N_2110,N_1968,N_1872);
and U2111 (N_2111,N_1631,N_1972);
or U2112 (N_2112,N_1881,N_1827);
nand U2113 (N_2113,N_1520,N_1662);
xnor U2114 (N_2114,N_1609,N_1516);
or U2115 (N_2115,N_1790,N_1509);
or U2116 (N_2116,N_1690,N_1699);
nor U2117 (N_2117,N_1782,N_1837);
or U2118 (N_2118,N_1824,N_1585);
nor U2119 (N_2119,N_1583,N_1918);
nand U2120 (N_2120,N_1840,N_1917);
nor U2121 (N_2121,N_1620,N_1715);
or U2122 (N_2122,N_1791,N_1598);
or U2123 (N_2123,N_1518,N_1574);
xnor U2124 (N_2124,N_1526,N_1692);
xnor U2125 (N_2125,N_1743,N_1882);
nand U2126 (N_2126,N_1798,N_1780);
nor U2127 (N_2127,N_1615,N_1844);
nand U2128 (N_2128,N_1860,N_1749);
and U2129 (N_2129,N_1675,N_1899);
or U2130 (N_2130,N_1640,N_1677);
nand U2131 (N_2131,N_1904,N_1974);
xnor U2132 (N_2132,N_1597,N_1915);
or U2133 (N_2133,N_1889,N_1702);
nor U2134 (N_2134,N_1877,N_1826);
and U2135 (N_2135,N_1708,N_1600);
xor U2136 (N_2136,N_1617,N_1591);
nor U2137 (N_2137,N_1667,N_1612);
and U2138 (N_2138,N_1537,N_1548);
and U2139 (N_2139,N_1838,N_1969);
and U2140 (N_2140,N_1726,N_1772);
nand U2141 (N_2141,N_1513,N_1829);
or U2142 (N_2142,N_1990,N_1810);
xnor U2143 (N_2143,N_1588,N_1724);
nand U2144 (N_2144,N_1697,N_1748);
nand U2145 (N_2145,N_1815,N_1656);
and U2146 (N_2146,N_1622,N_1560);
and U2147 (N_2147,N_1735,N_1545);
and U2148 (N_2148,N_1628,N_1988);
and U2149 (N_2149,N_1897,N_1755);
xnor U2150 (N_2150,N_1953,N_1935);
and U2151 (N_2151,N_1946,N_1927);
or U2152 (N_2152,N_1981,N_1807);
nand U2153 (N_2153,N_1800,N_1626);
xor U2154 (N_2154,N_1818,N_1645);
xor U2155 (N_2155,N_1698,N_1763);
xor U2156 (N_2156,N_1785,N_1561);
nand U2157 (N_2157,N_1512,N_1852);
xnor U2158 (N_2158,N_1504,N_1719);
or U2159 (N_2159,N_1880,N_1891);
or U2160 (N_2160,N_1752,N_1850);
or U2161 (N_2161,N_1975,N_1732);
or U2162 (N_2162,N_1716,N_1687);
nor U2163 (N_2163,N_1594,N_1610);
xor U2164 (N_2164,N_1655,N_1811);
and U2165 (N_2165,N_1857,N_1557);
xnor U2166 (N_2166,N_1564,N_1712);
and U2167 (N_2167,N_1674,N_1983);
nor U2168 (N_2168,N_1856,N_1584);
or U2169 (N_2169,N_1569,N_1982);
or U2170 (N_2170,N_1558,N_1689);
or U2171 (N_2171,N_1582,N_1602);
nor U2172 (N_2172,N_1664,N_1931);
nor U2173 (N_2173,N_1660,N_1854);
and U2174 (N_2174,N_1742,N_1550);
nor U2175 (N_2175,N_1757,N_1806);
nand U2176 (N_2176,N_1579,N_1853);
nand U2177 (N_2177,N_1686,N_1909);
xor U2178 (N_2178,N_1973,N_1795);
nand U2179 (N_2179,N_1893,N_1802);
and U2180 (N_2180,N_1511,N_1959);
or U2181 (N_2181,N_1820,N_1803);
xor U2182 (N_2182,N_1895,N_1554);
nand U2183 (N_2183,N_1589,N_1555);
and U2184 (N_2184,N_1535,N_1793);
nand U2185 (N_2185,N_1867,N_1839);
nor U2186 (N_2186,N_1623,N_1750);
and U2187 (N_2187,N_1653,N_1616);
or U2188 (N_2188,N_1556,N_1849);
nor U2189 (N_2189,N_1734,N_1682);
nor U2190 (N_2190,N_1635,N_1522);
xnor U2191 (N_2191,N_1768,N_1778);
and U2192 (N_2192,N_1835,N_1812);
xnor U2193 (N_2193,N_1565,N_1648);
and U2194 (N_2194,N_1738,N_1604);
or U2195 (N_2195,N_1842,N_1996);
nand U2196 (N_2196,N_1563,N_1696);
xor U2197 (N_2197,N_1507,N_1966);
nor U2198 (N_2198,N_1833,N_1736);
xnor U2199 (N_2199,N_1870,N_1701);
nor U2200 (N_2200,N_1930,N_1843);
nand U2201 (N_2201,N_1952,N_1783);
nor U2202 (N_2202,N_1847,N_1967);
nor U2203 (N_2203,N_1971,N_1762);
nand U2204 (N_2204,N_1572,N_1671);
or U2205 (N_2205,N_1878,N_1542);
and U2206 (N_2206,N_1727,N_1592);
and U2207 (N_2207,N_1669,N_1711);
nor U2208 (N_2208,N_1794,N_1960);
or U2209 (N_2209,N_1916,N_1741);
nor U2210 (N_2210,N_1875,N_1764);
nor U2211 (N_2211,N_1753,N_1552);
nand U2212 (N_2212,N_1759,N_1590);
nor U2213 (N_2213,N_1654,N_1944);
nor U2214 (N_2214,N_1871,N_1643);
or U2215 (N_2215,N_1797,N_1672);
nand U2216 (N_2216,N_1941,N_1614);
or U2217 (N_2217,N_1977,N_1646);
and U2218 (N_2218,N_1932,N_1956);
nor U2219 (N_2219,N_1955,N_1530);
or U2220 (N_2220,N_1641,N_1691);
nand U2221 (N_2221,N_1908,N_1796);
and U2222 (N_2222,N_1706,N_1637);
xnor U2223 (N_2223,N_1942,N_1831);
nand U2224 (N_2224,N_1890,N_1761);
and U2225 (N_2225,N_1900,N_1577);
xor U2226 (N_2226,N_1929,N_1789);
xnor U2227 (N_2227,N_1580,N_1728);
or U2228 (N_2228,N_1976,N_1777);
or U2229 (N_2229,N_1813,N_1801);
nor U2230 (N_2230,N_1775,N_1924);
or U2231 (N_2231,N_1673,N_1657);
or U2232 (N_2232,N_1865,N_1822);
and U2233 (N_2233,N_1845,N_1725);
xor U2234 (N_2234,N_1521,N_1551);
or U2235 (N_2235,N_1714,N_1751);
and U2236 (N_2236,N_1949,N_1559);
xor U2237 (N_2237,N_1532,N_1733);
nand U2238 (N_2238,N_1679,N_1683);
xor U2239 (N_2239,N_1804,N_1596);
xor U2240 (N_2240,N_1995,N_1814);
and U2241 (N_2241,N_1652,N_1630);
nand U2242 (N_2242,N_1505,N_1544);
nor U2243 (N_2243,N_1705,N_1906);
and U2244 (N_2244,N_1770,N_1536);
nor U2245 (N_2245,N_1595,N_1659);
nor U2246 (N_2246,N_1928,N_1578);
and U2247 (N_2247,N_1624,N_1767);
and U2248 (N_2248,N_1788,N_1684);
nand U2249 (N_2249,N_1703,N_1633);
or U2250 (N_2250,N_1579,N_1923);
nor U2251 (N_2251,N_1539,N_1997);
and U2252 (N_2252,N_1752,N_1799);
and U2253 (N_2253,N_1990,N_1716);
xor U2254 (N_2254,N_1952,N_1613);
or U2255 (N_2255,N_1885,N_1932);
nand U2256 (N_2256,N_1799,N_1708);
nand U2257 (N_2257,N_1603,N_1644);
nand U2258 (N_2258,N_1794,N_1693);
nor U2259 (N_2259,N_1778,N_1733);
and U2260 (N_2260,N_1730,N_1753);
xor U2261 (N_2261,N_1645,N_1527);
xnor U2262 (N_2262,N_1542,N_1825);
and U2263 (N_2263,N_1537,N_1927);
xnor U2264 (N_2264,N_1810,N_1534);
and U2265 (N_2265,N_1880,N_1562);
or U2266 (N_2266,N_1677,N_1941);
nand U2267 (N_2267,N_1871,N_1989);
xor U2268 (N_2268,N_1551,N_1507);
or U2269 (N_2269,N_1914,N_1834);
xnor U2270 (N_2270,N_1862,N_1543);
nand U2271 (N_2271,N_1533,N_1810);
and U2272 (N_2272,N_1554,N_1776);
nor U2273 (N_2273,N_1578,N_1955);
or U2274 (N_2274,N_1813,N_1961);
nand U2275 (N_2275,N_1930,N_1868);
xnor U2276 (N_2276,N_1862,N_1925);
nand U2277 (N_2277,N_1769,N_1738);
nor U2278 (N_2278,N_1616,N_1740);
xnor U2279 (N_2279,N_1836,N_1550);
and U2280 (N_2280,N_1622,N_1561);
or U2281 (N_2281,N_1604,N_1826);
nand U2282 (N_2282,N_1735,N_1693);
xor U2283 (N_2283,N_1545,N_1593);
xnor U2284 (N_2284,N_1806,N_1611);
or U2285 (N_2285,N_1914,N_1692);
and U2286 (N_2286,N_1847,N_1854);
nor U2287 (N_2287,N_1718,N_1728);
and U2288 (N_2288,N_1741,N_1828);
and U2289 (N_2289,N_1612,N_1819);
nand U2290 (N_2290,N_1700,N_1878);
nand U2291 (N_2291,N_1719,N_1819);
and U2292 (N_2292,N_1714,N_1899);
nor U2293 (N_2293,N_1670,N_1568);
or U2294 (N_2294,N_1643,N_1774);
xnor U2295 (N_2295,N_1947,N_1887);
xor U2296 (N_2296,N_1574,N_1851);
nand U2297 (N_2297,N_1986,N_1729);
and U2298 (N_2298,N_1883,N_1805);
nor U2299 (N_2299,N_1863,N_1801);
nor U2300 (N_2300,N_1729,N_1801);
xnor U2301 (N_2301,N_1746,N_1861);
nand U2302 (N_2302,N_1825,N_1849);
or U2303 (N_2303,N_1795,N_1749);
or U2304 (N_2304,N_1894,N_1716);
nor U2305 (N_2305,N_1698,N_1527);
xnor U2306 (N_2306,N_1620,N_1806);
nand U2307 (N_2307,N_1552,N_1810);
or U2308 (N_2308,N_1978,N_1726);
xor U2309 (N_2309,N_1500,N_1986);
or U2310 (N_2310,N_1695,N_1931);
and U2311 (N_2311,N_1772,N_1566);
xnor U2312 (N_2312,N_1707,N_1696);
nand U2313 (N_2313,N_1846,N_1741);
nor U2314 (N_2314,N_1508,N_1976);
nand U2315 (N_2315,N_1736,N_1758);
nand U2316 (N_2316,N_1790,N_1609);
nor U2317 (N_2317,N_1956,N_1821);
or U2318 (N_2318,N_1716,N_1865);
nand U2319 (N_2319,N_1950,N_1568);
or U2320 (N_2320,N_1555,N_1889);
xor U2321 (N_2321,N_1537,N_1858);
nand U2322 (N_2322,N_1966,N_1794);
or U2323 (N_2323,N_1790,N_1676);
and U2324 (N_2324,N_1606,N_1524);
or U2325 (N_2325,N_1757,N_1707);
or U2326 (N_2326,N_1589,N_1902);
and U2327 (N_2327,N_1778,N_1806);
and U2328 (N_2328,N_1720,N_1867);
xor U2329 (N_2329,N_1727,N_1738);
or U2330 (N_2330,N_1818,N_1947);
nand U2331 (N_2331,N_1637,N_1607);
nand U2332 (N_2332,N_1561,N_1907);
nor U2333 (N_2333,N_1877,N_1882);
xnor U2334 (N_2334,N_1745,N_1989);
or U2335 (N_2335,N_1751,N_1884);
nor U2336 (N_2336,N_1884,N_1514);
nand U2337 (N_2337,N_1671,N_1834);
nor U2338 (N_2338,N_1562,N_1686);
or U2339 (N_2339,N_1678,N_1535);
or U2340 (N_2340,N_1988,N_1926);
or U2341 (N_2341,N_1665,N_1907);
nor U2342 (N_2342,N_1511,N_1900);
and U2343 (N_2343,N_1735,N_1998);
or U2344 (N_2344,N_1986,N_1523);
xor U2345 (N_2345,N_1607,N_1768);
xnor U2346 (N_2346,N_1728,N_1858);
xnor U2347 (N_2347,N_1542,N_1661);
nor U2348 (N_2348,N_1573,N_1860);
or U2349 (N_2349,N_1740,N_1892);
xor U2350 (N_2350,N_1557,N_1654);
and U2351 (N_2351,N_1667,N_1983);
and U2352 (N_2352,N_1640,N_1983);
xnor U2353 (N_2353,N_1659,N_1832);
nor U2354 (N_2354,N_1830,N_1877);
nor U2355 (N_2355,N_1730,N_1672);
or U2356 (N_2356,N_1591,N_1759);
and U2357 (N_2357,N_1969,N_1514);
nand U2358 (N_2358,N_1775,N_1727);
nor U2359 (N_2359,N_1550,N_1961);
and U2360 (N_2360,N_1716,N_1621);
or U2361 (N_2361,N_1710,N_1969);
or U2362 (N_2362,N_1578,N_1963);
nor U2363 (N_2363,N_1549,N_1678);
or U2364 (N_2364,N_1513,N_1655);
nand U2365 (N_2365,N_1725,N_1594);
and U2366 (N_2366,N_1586,N_1524);
nor U2367 (N_2367,N_1842,N_1737);
and U2368 (N_2368,N_1959,N_1870);
nand U2369 (N_2369,N_1744,N_1674);
nand U2370 (N_2370,N_1985,N_1768);
and U2371 (N_2371,N_1699,N_1924);
xnor U2372 (N_2372,N_1563,N_1586);
nand U2373 (N_2373,N_1765,N_1651);
nand U2374 (N_2374,N_1931,N_1712);
nand U2375 (N_2375,N_1928,N_1740);
or U2376 (N_2376,N_1509,N_1742);
nor U2377 (N_2377,N_1801,N_1566);
nand U2378 (N_2378,N_1780,N_1573);
nand U2379 (N_2379,N_1751,N_1532);
xnor U2380 (N_2380,N_1743,N_1751);
or U2381 (N_2381,N_1711,N_1645);
nor U2382 (N_2382,N_1541,N_1762);
xnor U2383 (N_2383,N_1963,N_1949);
xor U2384 (N_2384,N_1737,N_1934);
and U2385 (N_2385,N_1662,N_1743);
nand U2386 (N_2386,N_1570,N_1722);
nand U2387 (N_2387,N_1898,N_1671);
or U2388 (N_2388,N_1765,N_1986);
xnor U2389 (N_2389,N_1611,N_1685);
nor U2390 (N_2390,N_1937,N_1690);
nor U2391 (N_2391,N_1788,N_1901);
or U2392 (N_2392,N_1594,N_1898);
and U2393 (N_2393,N_1534,N_1841);
nand U2394 (N_2394,N_1844,N_1864);
nor U2395 (N_2395,N_1592,N_1647);
xor U2396 (N_2396,N_1647,N_1928);
nor U2397 (N_2397,N_1709,N_1995);
nand U2398 (N_2398,N_1741,N_1804);
xnor U2399 (N_2399,N_1611,N_1830);
or U2400 (N_2400,N_1783,N_1883);
or U2401 (N_2401,N_1699,N_1910);
and U2402 (N_2402,N_1855,N_1948);
and U2403 (N_2403,N_1962,N_1644);
or U2404 (N_2404,N_1851,N_1670);
nand U2405 (N_2405,N_1962,N_1809);
nor U2406 (N_2406,N_1520,N_1994);
or U2407 (N_2407,N_1502,N_1689);
and U2408 (N_2408,N_1586,N_1654);
xor U2409 (N_2409,N_1631,N_1927);
xnor U2410 (N_2410,N_1696,N_1792);
nor U2411 (N_2411,N_1518,N_1649);
nor U2412 (N_2412,N_1985,N_1845);
or U2413 (N_2413,N_1789,N_1560);
or U2414 (N_2414,N_1982,N_1690);
nor U2415 (N_2415,N_1908,N_1807);
nor U2416 (N_2416,N_1560,N_1655);
and U2417 (N_2417,N_1937,N_1582);
xor U2418 (N_2418,N_1745,N_1500);
nor U2419 (N_2419,N_1686,N_1948);
xor U2420 (N_2420,N_1968,N_1738);
nand U2421 (N_2421,N_1851,N_1988);
or U2422 (N_2422,N_1597,N_1652);
xnor U2423 (N_2423,N_1643,N_1652);
or U2424 (N_2424,N_1517,N_1888);
nand U2425 (N_2425,N_1776,N_1507);
nor U2426 (N_2426,N_1830,N_1944);
xnor U2427 (N_2427,N_1624,N_1565);
and U2428 (N_2428,N_1872,N_1687);
and U2429 (N_2429,N_1902,N_1620);
nand U2430 (N_2430,N_1520,N_1885);
nor U2431 (N_2431,N_1920,N_1951);
and U2432 (N_2432,N_1755,N_1749);
nor U2433 (N_2433,N_1973,N_1971);
nor U2434 (N_2434,N_1669,N_1517);
or U2435 (N_2435,N_1695,N_1722);
or U2436 (N_2436,N_1674,N_1733);
xnor U2437 (N_2437,N_1615,N_1647);
nand U2438 (N_2438,N_1695,N_1645);
or U2439 (N_2439,N_1700,N_1806);
xnor U2440 (N_2440,N_1990,N_1978);
nand U2441 (N_2441,N_1689,N_1893);
nand U2442 (N_2442,N_1752,N_1867);
nand U2443 (N_2443,N_1688,N_1963);
and U2444 (N_2444,N_1839,N_1813);
nand U2445 (N_2445,N_1560,N_1775);
xor U2446 (N_2446,N_1980,N_1958);
or U2447 (N_2447,N_1864,N_1672);
nand U2448 (N_2448,N_1503,N_1929);
or U2449 (N_2449,N_1668,N_1941);
and U2450 (N_2450,N_1749,N_1506);
xor U2451 (N_2451,N_1975,N_1738);
or U2452 (N_2452,N_1678,N_1848);
nand U2453 (N_2453,N_1850,N_1938);
or U2454 (N_2454,N_1591,N_1990);
nand U2455 (N_2455,N_1820,N_1903);
and U2456 (N_2456,N_1948,N_1523);
or U2457 (N_2457,N_1907,N_1992);
nand U2458 (N_2458,N_1861,N_1729);
and U2459 (N_2459,N_1761,N_1854);
nor U2460 (N_2460,N_1945,N_1875);
or U2461 (N_2461,N_1542,N_1962);
and U2462 (N_2462,N_1798,N_1520);
or U2463 (N_2463,N_1816,N_1883);
or U2464 (N_2464,N_1709,N_1522);
and U2465 (N_2465,N_1595,N_1862);
xor U2466 (N_2466,N_1837,N_1769);
nand U2467 (N_2467,N_1998,N_1682);
and U2468 (N_2468,N_1756,N_1750);
and U2469 (N_2469,N_1572,N_1568);
or U2470 (N_2470,N_1568,N_1836);
nor U2471 (N_2471,N_1715,N_1846);
nor U2472 (N_2472,N_1877,N_1704);
or U2473 (N_2473,N_1842,N_1656);
and U2474 (N_2474,N_1894,N_1576);
and U2475 (N_2475,N_1598,N_1896);
and U2476 (N_2476,N_1585,N_1599);
and U2477 (N_2477,N_1868,N_1707);
or U2478 (N_2478,N_1892,N_1606);
or U2479 (N_2479,N_1846,N_1913);
nand U2480 (N_2480,N_1850,N_1952);
nand U2481 (N_2481,N_1942,N_1822);
or U2482 (N_2482,N_1920,N_1833);
nand U2483 (N_2483,N_1592,N_1782);
nand U2484 (N_2484,N_1913,N_1635);
and U2485 (N_2485,N_1548,N_1759);
or U2486 (N_2486,N_1836,N_1751);
nor U2487 (N_2487,N_1534,N_1872);
nand U2488 (N_2488,N_1808,N_1776);
nand U2489 (N_2489,N_1959,N_1559);
nand U2490 (N_2490,N_1875,N_1575);
xor U2491 (N_2491,N_1703,N_1768);
and U2492 (N_2492,N_1656,N_1615);
xor U2493 (N_2493,N_1962,N_1511);
or U2494 (N_2494,N_1888,N_1817);
nand U2495 (N_2495,N_1813,N_1959);
nor U2496 (N_2496,N_1765,N_1512);
xnor U2497 (N_2497,N_1819,N_1838);
or U2498 (N_2498,N_1841,N_1594);
or U2499 (N_2499,N_1690,N_1576);
and U2500 (N_2500,N_2390,N_2000);
and U2501 (N_2501,N_2041,N_2449);
xnor U2502 (N_2502,N_2331,N_2388);
nor U2503 (N_2503,N_2306,N_2012);
and U2504 (N_2504,N_2206,N_2359);
nor U2505 (N_2505,N_2278,N_2383);
xor U2506 (N_2506,N_2344,N_2322);
or U2507 (N_2507,N_2029,N_2290);
nor U2508 (N_2508,N_2349,N_2375);
and U2509 (N_2509,N_2469,N_2251);
and U2510 (N_2510,N_2490,N_2242);
xnor U2511 (N_2511,N_2389,N_2401);
xor U2512 (N_2512,N_2455,N_2396);
nor U2513 (N_2513,N_2124,N_2122);
xnor U2514 (N_2514,N_2131,N_2297);
nor U2515 (N_2515,N_2072,N_2275);
nand U2516 (N_2516,N_2031,N_2445);
nor U2517 (N_2517,N_2234,N_2162);
nand U2518 (N_2518,N_2354,N_2193);
nor U2519 (N_2519,N_2304,N_2332);
and U2520 (N_2520,N_2498,N_2194);
nand U2521 (N_2521,N_2285,N_2456);
nor U2522 (N_2522,N_2220,N_2374);
xor U2523 (N_2523,N_2033,N_2319);
xnor U2524 (N_2524,N_2446,N_2093);
and U2525 (N_2525,N_2026,N_2288);
or U2526 (N_2526,N_2071,N_2148);
nand U2527 (N_2527,N_2164,N_2059);
nor U2528 (N_2528,N_2398,N_2064);
xor U2529 (N_2529,N_2014,N_2001);
nand U2530 (N_2530,N_2257,N_2021);
or U2531 (N_2531,N_2249,N_2461);
xnor U2532 (N_2532,N_2235,N_2168);
and U2533 (N_2533,N_2002,N_2320);
nand U2534 (N_2534,N_2423,N_2066);
and U2535 (N_2535,N_2136,N_2287);
and U2536 (N_2536,N_2296,N_2070);
xnor U2537 (N_2537,N_2318,N_2092);
xor U2538 (N_2538,N_2454,N_2310);
nor U2539 (N_2539,N_2274,N_2419);
nor U2540 (N_2540,N_2203,N_2458);
xnor U2541 (N_2541,N_2459,N_2341);
or U2542 (N_2542,N_2244,N_2317);
and U2543 (N_2543,N_2025,N_2229);
nor U2544 (N_2544,N_2085,N_2163);
nand U2545 (N_2545,N_2049,N_2007);
and U2546 (N_2546,N_2178,N_2345);
nand U2547 (N_2547,N_2057,N_2003);
nand U2548 (N_2548,N_2065,N_2460);
or U2549 (N_2549,N_2335,N_2447);
xnor U2550 (N_2550,N_2422,N_2139);
and U2551 (N_2551,N_2437,N_2201);
and U2552 (N_2552,N_2160,N_2470);
or U2553 (N_2553,N_2183,N_2333);
and U2554 (N_2554,N_2264,N_2156);
and U2555 (N_2555,N_2327,N_2165);
nor U2556 (N_2556,N_2429,N_2247);
nor U2557 (N_2557,N_2427,N_2202);
nor U2558 (N_2558,N_2110,N_2410);
or U2559 (N_2559,N_2425,N_2030);
nor U2560 (N_2560,N_2323,N_2051);
xor U2561 (N_2561,N_2191,N_2276);
nor U2562 (N_2562,N_2100,N_2017);
xor U2563 (N_2563,N_2279,N_2062);
nor U2564 (N_2564,N_2137,N_2240);
or U2565 (N_2565,N_2166,N_2097);
xnor U2566 (N_2566,N_2364,N_2439);
nor U2567 (N_2567,N_2146,N_2260);
xor U2568 (N_2568,N_2102,N_2385);
or U2569 (N_2569,N_2262,N_2495);
xnor U2570 (N_2570,N_2265,N_2267);
nand U2571 (N_2571,N_2207,N_2232);
nand U2572 (N_2572,N_2491,N_2431);
xor U2573 (N_2573,N_2121,N_2176);
or U2574 (N_2574,N_2208,N_2329);
and U2575 (N_2575,N_2263,N_2302);
or U2576 (N_2576,N_2105,N_2330);
nor U2577 (N_2577,N_2067,N_2069);
xor U2578 (N_2578,N_2357,N_2411);
nand U2579 (N_2579,N_2301,N_2312);
and U2580 (N_2580,N_2395,N_2473);
nand U2581 (N_2581,N_2482,N_2409);
nand U2582 (N_2582,N_2205,N_2078);
xor U2583 (N_2583,N_2213,N_2352);
or U2584 (N_2584,N_2119,N_2204);
and U2585 (N_2585,N_2334,N_2032);
nor U2586 (N_2586,N_2252,N_2298);
xnor U2587 (N_2587,N_2315,N_2476);
nand U2588 (N_2588,N_2045,N_2080);
nor U2589 (N_2589,N_2231,N_2196);
or U2590 (N_2590,N_2038,N_2272);
xor U2591 (N_2591,N_2015,N_2358);
xnor U2592 (N_2592,N_2426,N_2488);
or U2593 (N_2593,N_2462,N_2484);
nor U2594 (N_2594,N_2467,N_2087);
nor U2595 (N_2595,N_2496,N_2363);
and U2596 (N_2596,N_2039,N_2442);
and U2597 (N_2597,N_2475,N_2369);
nor U2598 (N_2598,N_2403,N_2351);
or U2599 (N_2599,N_2010,N_2060);
nand U2600 (N_2600,N_2299,N_2083);
or U2601 (N_2601,N_2474,N_2273);
nor U2602 (N_2602,N_2348,N_2372);
or U2603 (N_2603,N_2440,N_2186);
nand U2604 (N_2604,N_2211,N_2424);
xor U2605 (N_2605,N_2173,N_2241);
or U2606 (N_2606,N_2120,N_2394);
nor U2607 (N_2607,N_2271,N_2313);
nand U2608 (N_2608,N_2169,N_2144);
xor U2609 (N_2609,N_2292,N_2406);
or U2610 (N_2610,N_2150,N_2471);
xor U2611 (N_2611,N_2487,N_2103);
nand U2612 (N_2612,N_2174,N_2326);
and U2613 (N_2613,N_2035,N_2384);
xor U2614 (N_2614,N_2068,N_2457);
xor U2615 (N_2615,N_2036,N_2436);
or U2616 (N_2616,N_2195,N_2126);
xor U2617 (N_2617,N_2305,N_2192);
nand U2618 (N_2618,N_2382,N_2481);
and U2619 (N_2619,N_2309,N_2266);
or U2620 (N_2620,N_2238,N_2228);
and U2621 (N_2621,N_2413,N_2073);
xor U2622 (N_2622,N_2289,N_2008);
and U2623 (N_2623,N_2006,N_2020);
nand U2624 (N_2624,N_2114,N_2081);
nor U2625 (N_2625,N_2198,N_2189);
nand U2626 (N_2626,N_2155,N_2356);
nor U2627 (N_2627,N_2259,N_2005);
or U2628 (N_2628,N_2339,N_2056);
and U2629 (N_2629,N_2223,N_2089);
nor U2630 (N_2630,N_2418,N_2337);
or U2631 (N_2631,N_2421,N_2478);
nor U2632 (N_2632,N_2443,N_2101);
and U2633 (N_2633,N_2149,N_2061);
nor U2634 (N_2634,N_2052,N_2404);
xor U2635 (N_2635,N_2245,N_2107);
nor U2636 (N_2636,N_2050,N_2258);
and U2637 (N_2637,N_2493,N_2058);
nor U2638 (N_2638,N_2397,N_2082);
nand U2639 (N_2639,N_2226,N_2172);
nor U2640 (N_2640,N_2353,N_2415);
and U2641 (N_2641,N_2098,N_2291);
and U2642 (N_2642,N_2453,N_2261);
nand U2643 (N_2643,N_2355,N_2044);
nand U2644 (N_2644,N_2116,N_2040);
nor U2645 (N_2645,N_2111,N_2379);
nand U2646 (N_2646,N_2253,N_2376);
nand U2647 (N_2647,N_2308,N_2043);
nand U2648 (N_2648,N_2016,N_2400);
nor U2649 (N_2649,N_2132,N_2371);
and U2650 (N_2650,N_2286,N_2479);
or U2651 (N_2651,N_2294,N_2464);
or U2652 (N_2652,N_2485,N_2167);
nor U2653 (N_2653,N_2325,N_2377);
xor U2654 (N_2654,N_2115,N_2412);
or U2655 (N_2655,N_2281,N_2210);
nand U2656 (N_2656,N_2405,N_2347);
and U2657 (N_2657,N_2343,N_2350);
nor U2658 (N_2658,N_2284,N_2141);
nand U2659 (N_2659,N_2328,N_2336);
nor U2660 (N_2660,N_2316,N_2366);
nor U2661 (N_2661,N_2477,N_2143);
xnor U2662 (N_2662,N_2130,N_2048);
nor U2663 (N_2663,N_2441,N_2187);
nand U2664 (N_2664,N_2361,N_2147);
or U2665 (N_2665,N_2188,N_2280);
nor U2666 (N_2666,N_2074,N_2268);
and U2667 (N_2667,N_2293,N_2159);
and U2668 (N_2668,N_2435,N_2138);
nor U2669 (N_2669,N_2209,N_2179);
xor U2670 (N_2670,N_2387,N_2019);
xor U2671 (N_2671,N_2282,N_2157);
and U2672 (N_2672,N_2434,N_2090);
xor U2673 (N_2673,N_2311,N_2129);
nand U2674 (N_2674,N_2123,N_2135);
or U2675 (N_2675,N_2133,N_2054);
nor U2676 (N_2676,N_2407,N_2218);
nand U2677 (N_2677,N_2451,N_2145);
xor U2678 (N_2678,N_2084,N_2125);
xor U2679 (N_2679,N_2380,N_2248);
nor U2680 (N_2680,N_2024,N_2483);
nor U2681 (N_2681,N_2055,N_2112);
and U2682 (N_2682,N_2200,N_2117);
xor U2683 (N_2683,N_2047,N_2236);
xor U2684 (N_2684,N_2321,N_2381);
nand U2685 (N_2685,N_2037,N_2499);
xnor U2686 (N_2686,N_2221,N_2199);
xnor U2687 (N_2687,N_2324,N_2450);
nor U2688 (N_2688,N_2185,N_2212);
nor U2689 (N_2689,N_2393,N_2079);
and U2690 (N_2690,N_2362,N_2108);
nor U2691 (N_2691,N_2215,N_2127);
or U2692 (N_2692,N_2452,N_2433);
and U2693 (N_2693,N_2161,N_2018);
nor U2694 (N_2694,N_2128,N_2300);
and U2695 (N_2695,N_2307,N_2094);
nand U2696 (N_2696,N_2134,N_2180);
xnor U2697 (N_2697,N_2270,N_2414);
nor U2698 (N_2698,N_2170,N_2346);
xor U2699 (N_2699,N_2239,N_2340);
nor U2700 (N_2700,N_2444,N_2432);
and U2701 (N_2701,N_2486,N_2011);
xnor U2702 (N_2702,N_2184,N_2466);
nor U2703 (N_2703,N_2053,N_2468);
nand U2704 (N_2704,N_2237,N_2338);
nand U2705 (N_2705,N_2225,N_2028);
or U2706 (N_2706,N_2256,N_2182);
xor U2707 (N_2707,N_2255,N_2153);
and U2708 (N_2708,N_2140,N_2408);
xor U2709 (N_2709,N_2095,N_2027);
xor U2710 (N_2710,N_2042,N_2392);
and U2711 (N_2711,N_2013,N_2277);
nor U2712 (N_2712,N_2378,N_2214);
nand U2713 (N_2713,N_2386,N_2365);
nand U2714 (N_2714,N_2086,N_2233);
or U2715 (N_2715,N_2494,N_2216);
xnor U2716 (N_2716,N_2190,N_2106);
nand U2717 (N_2717,N_2076,N_2391);
nand U2718 (N_2718,N_2370,N_2246);
or U2719 (N_2719,N_2472,N_2243);
or U2720 (N_2720,N_2109,N_2152);
or U2721 (N_2721,N_2181,N_2046);
nand U2722 (N_2722,N_2171,N_2283);
nor U2723 (N_2723,N_2099,N_2142);
xnor U2724 (N_2724,N_2254,N_2091);
or U2725 (N_2725,N_2004,N_2492);
and U2726 (N_2726,N_2420,N_2063);
nand U2727 (N_2727,N_2177,N_2022);
xnor U2728 (N_2728,N_2088,N_2230);
and U2729 (N_2729,N_2360,N_2104);
or U2730 (N_2730,N_2428,N_2463);
nand U2731 (N_2731,N_2367,N_2250);
nor U2732 (N_2732,N_2096,N_2314);
nor U2733 (N_2733,N_2113,N_2154);
and U2734 (N_2734,N_2448,N_2465);
or U2735 (N_2735,N_2224,N_2269);
nand U2736 (N_2736,N_2217,N_2023);
or U2737 (N_2737,N_2077,N_2402);
and U2738 (N_2738,N_2118,N_2219);
nor U2739 (N_2739,N_2222,N_2158);
or U2740 (N_2740,N_2489,N_2009);
nor U2741 (N_2741,N_2151,N_2417);
and U2742 (N_2742,N_2430,N_2175);
and U2743 (N_2743,N_2416,N_2497);
and U2744 (N_2744,N_2295,N_2197);
nand U2745 (N_2745,N_2034,N_2342);
and U2746 (N_2746,N_2303,N_2227);
nand U2747 (N_2747,N_2368,N_2438);
and U2748 (N_2748,N_2075,N_2399);
or U2749 (N_2749,N_2373,N_2480);
xor U2750 (N_2750,N_2370,N_2379);
and U2751 (N_2751,N_2152,N_2438);
nand U2752 (N_2752,N_2081,N_2384);
nand U2753 (N_2753,N_2367,N_2134);
nor U2754 (N_2754,N_2025,N_2446);
xor U2755 (N_2755,N_2379,N_2225);
or U2756 (N_2756,N_2239,N_2090);
nand U2757 (N_2757,N_2343,N_2250);
and U2758 (N_2758,N_2484,N_2398);
nor U2759 (N_2759,N_2298,N_2177);
xnor U2760 (N_2760,N_2330,N_2071);
nand U2761 (N_2761,N_2009,N_2379);
xnor U2762 (N_2762,N_2030,N_2407);
nand U2763 (N_2763,N_2294,N_2358);
and U2764 (N_2764,N_2018,N_2070);
nor U2765 (N_2765,N_2325,N_2114);
nor U2766 (N_2766,N_2151,N_2378);
xnor U2767 (N_2767,N_2106,N_2175);
and U2768 (N_2768,N_2266,N_2058);
and U2769 (N_2769,N_2092,N_2211);
or U2770 (N_2770,N_2121,N_2253);
xor U2771 (N_2771,N_2212,N_2491);
nand U2772 (N_2772,N_2383,N_2007);
xnor U2773 (N_2773,N_2258,N_2357);
xor U2774 (N_2774,N_2455,N_2494);
nor U2775 (N_2775,N_2253,N_2411);
and U2776 (N_2776,N_2126,N_2320);
and U2777 (N_2777,N_2046,N_2296);
nor U2778 (N_2778,N_2484,N_2086);
nand U2779 (N_2779,N_2177,N_2236);
and U2780 (N_2780,N_2097,N_2139);
nor U2781 (N_2781,N_2017,N_2012);
nand U2782 (N_2782,N_2068,N_2148);
nor U2783 (N_2783,N_2298,N_2277);
nor U2784 (N_2784,N_2301,N_2014);
or U2785 (N_2785,N_2475,N_2025);
xor U2786 (N_2786,N_2490,N_2029);
nor U2787 (N_2787,N_2454,N_2090);
xnor U2788 (N_2788,N_2413,N_2481);
nor U2789 (N_2789,N_2312,N_2418);
nand U2790 (N_2790,N_2401,N_2241);
xnor U2791 (N_2791,N_2293,N_2147);
or U2792 (N_2792,N_2490,N_2137);
and U2793 (N_2793,N_2428,N_2163);
nor U2794 (N_2794,N_2419,N_2109);
nand U2795 (N_2795,N_2108,N_2106);
xnor U2796 (N_2796,N_2293,N_2485);
or U2797 (N_2797,N_2060,N_2465);
xor U2798 (N_2798,N_2018,N_2278);
and U2799 (N_2799,N_2469,N_2013);
or U2800 (N_2800,N_2451,N_2278);
or U2801 (N_2801,N_2392,N_2405);
xor U2802 (N_2802,N_2172,N_2433);
nor U2803 (N_2803,N_2485,N_2247);
or U2804 (N_2804,N_2018,N_2353);
or U2805 (N_2805,N_2189,N_2383);
and U2806 (N_2806,N_2388,N_2275);
xor U2807 (N_2807,N_2467,N_2138);
and U2808 (N_2808,N_2051,N_2017);
or U2809 (N_2809,N_2033,N_2001);
nor U2810 (N_2810,N_2324,N_2207);
and U2811 (N_2811,N_2337,N_2278);
or U2812 (N_2812,N_2499,N_2194);
xor U2813 (N_2813,N_2111,N_2178);
nor U2814 (N_2814,N_2090,N_2327);
xor U2815 (N_2815,N_2206,N_2128);
and U2816 (N_2816,N_2235,N_2383);
xor U2817 (N_2817,N_2057,N_2158);
nand U2818 (N_2818,N_2335,N_2221);
and U2819 (N_2819,N_2494,N_2142);
and U2820 (N_2820,N_2195,N_2410);
or U2821 (N_2821,N_2348,N_2064);
nor U2822 (N_2822,N_2030,N_2090);
or U2823 (N_2823,N_2285,N_2103);
or U2824 (N_2824,N_2469,N_2054);
or U2825 (N_2825,N_2459,N_2355);
nor U2826 (N_2826,N_2487,N_2498);
nand U2827 (N_2827,N_2417,N_2139);
or U2828 (N_2828,N_2324,N_2234);
xnor U2829 (N_2829,N_2406,N_2452);
nor U2830 (N_2830,N_2364,N_2169);
nor U2831 (N_2831,N_2134,N_2111);
nor U2832 (N_2832,N_2074,N_2077);
nor U2833 (N_2833,N_2220,N_2229);
nand U2834 (N_2834,N_2434,N_2284);
or U2835 (N_2835,N_2304,N_2445);
or U2836 (N_2836,N_2309,N_2140);
xnor U2837 (N_2837,N_2275,N_2479);
xnor U2838 (N_2838,N_2249,N_2175);
nand U2839 (N_2839,N_2442,N_2249);
or U2840 (N_2840,N_2170,N_2008);
nand U2841 (N_2841,N_2147,N_2272);
nor U2842 (N_2842,N_2077,N_2046);
or U2843 (N_2843,N_2344,N_2159);
and U2844 (N_2844,N_2421,N_2230);
xnor U2845 (N_2845,N_2435,N_2012);
or U2846 (N_2846,N_2170,N_2448);
nor U2847 (N_2847,N_2022,N_2043);
and U2848 (N_2848,N_2332,N_2264);
nor U2849 (N_2849,N_2091,N_2258);
xnor U2850 (N_2850,N_2291,N_2143);
nor U2851 (N_2851,N_2058,N_2178);
or U2852 (N_2852,N_2396,N_2476);
and U2853 (N_2853,N_2400,N_2039);
nand U2854 (N_2854,N_2072,N_2238);
nand U2855 (N_2855,N_2057,N_2317);
nand U2856 (N_2856,N_2177,N_2238);
xnor U2857 (N_2857,N_2011,N_2439);
or U2858 (N_2858,N_2469,N_2179);
nor U2859 (N_2859,N_2233,N_2398);
nor U2860 (N_2860,N_2022,N_2198);
nand U2861 (N_2861,N_2366,N_2471);
nor U2862 (N_2862,N_2315,N_2132);
nor U2863 (N_2863,N_2323,N_2261);
nand U2864 (N_2864,N_2025,N_2344);
and U2865 (N_2865,N_2109,N_2463);
xnor U2866 (N_2866,N_2037,N_2278);
nor U2867 (N_2867,N_2309,N_2284);
and U2868 (N_2868,N_2076,N_2316);
nand U2869 (N_2869,N_2147,N_2055);
nand U2870 (N_2870,N_2166,N_2474);
xnor U2871 (N_2871,N_2206,N_2124);
nand U2872 (N_2872,N_2080,N_2250);
and U2873 (N_2873,N_2499,N_2091);
xor U2874 (N_2874,N_2302,N_2025);
or U2875 (N_2875,N_2200,N_2241);
xnor U2876 (N_2876,N_2206,N_2149);
or U2877 (N_2877,N_2134,N_2093);
nor U2878 (N_2878,N_2238,N_2079);
or U2879 (N_2879,N_2446,N_2172);
nor U2880 (N_2880,N_2026,N_2476);
nand U2881 (N_2881,N_2360,N_2114);
or U2882 (N_2882,N_2089,N_2406);
nor U2883 (N_2883,N_2322,N_2149);
xor U2884 (N_2884,N_2142,N_2245);
nor U2885 (N_2885,N_2254,N_2234);
nand U2886 (N_2886,N_2185,N_2315);
nand U2887 (N_2887,N_2317,N_2150);
and U2888 (N_2888,N_2305,N_2043);
nand U2889 (N_2889,N_2493,N_2304);
xnor U2890 (N_2890,N_2207,N_2242);
xor U2891 (N_2891,N_2001,N_2103);
xnor U2892 (N_2892,N_2262,N_2036);
xor U2893 (N_2893,N_2442,N_2303);
nor U2894 (N_2894,N_2391,N_2433);
nor U2895 (N_2895,N_2108,N_2318);
nor U2896 (N_2896,N_2061,N_2041);
nor U2897 (N_2897,N_2154,N_2225);
and U2898 (N_2898,N_2271,N_2145);
nand U2899 (N_2899,N_2083,N_2268);
xor U2900 (N_2900,N_2304,N_2137);
xor U2901 (N_2901,N_2199,N_2341);
or U2902 (N_2902,N_2474,N_2081);
nor U2903 (N_2903,N_2093,N_2367);
and U2904 (N_2904,N_2193,N_2231);
xor U2905 (N_2905,N_2241,N_2003);
nor U2906 (N_2906,N_2071,N_2105);
xor U2907 (N_2907,N_2034,N_2098);
nor U2908 (N_2908,N_2243,N_2352);
xnor U2909 (N_2909,N_2056,N_2227);
nand U2910 (N_2910,N_2493,N_2153);
and U2911 (N_2911,N_2340,N_2113);
nand U2912 (N_2912,N_2198,N_2143);
xnor U2913 (N_2913,N_2287,N_2428);
nand U2914 (N_2914,N_2260,N_2001);
xor U2915 (N_2915,N_2339,N_2230);
or U2916 (N_2916,N_2009,N_2410);
xor U2917 (N_2917,N_2014,N_2121);
or U2918 (N_2918,N_2395,N_2130);
nand U2919 (N_2919,N_2447,N_2169);
xnor U2920 (N_2920,N_2346,N_2071);
and U2921 (N_2921,N_2090,N_2106);
or U2922 (N_2922,N_2375,N_2037);
nand U2923 (N_2923,N_2193,N_2173);
xor U2924 (N_2924,N_2202,N_2269);
nand U2925 (N_2925,N_2151,N_2034);
nor U2926 (N_2926,N_2038,N_2250);
xor U2927 (N_2927,N_2399,N_2361);
or U2928 (N_2928,N_2429,N_2376);
nand U2929 (N_2929,N_2085,N_2454);
or U2930 (N_2930,N_2227,N_2335);
and U2931 (N_2931,N_2052,N_2423);
or U2932 (N_2932,N_2233,N_2237);
nor U2933 (N_2933,N_2190,N_2470);
nor U2934 (N_2934,N_2202,N_2281);
nand U2935 (N_2935,N_2205,N_2004);
nor U2936 (N_2936,N_2347,N_2410);
and U2937 (N_2937,N_2132,N_2267);
nand U2938 (N_2938,N_2281,N_2084);
and U2939 (N_2939,N_2232,N_2345);
nor U2940 (N_2940,N_2457,N_2064);
nand U2941 (N_2941,N_2219,N_2280);
nand U2942 (N_2942,N_2407,N_2041);
and U2943 (N_2943,N_2080,N_2376);
or U2944 (N_2944,N_2278,N_2120);
or U2945 (N_2945,N_2149,N_2250);
nor U2946 (N_2946,N_2247,N_2259);
nor U2947 (N_2947,N_2187,N_2386);
nand U2948 (N_2948,N_2376,N_2489);
nand U2949 (N_2949,N_2372,N_2274);
and U2950 (N_2950,N_2281,N_2002);
nor U2951 (N_2951,N_2112,N_2377);
and U2952 (N_2952,N_2108,N_2168);
nor U2953 (N_2953,N_2430,N_2325);
or U2954 (N_2954,N_2379,N_2308);
xor U2955 (N_2955,N_2362,N_2429);
xnor U2956 (N_2956,N_2039,N_2094);
nor U2957 (N_2957,N_2119,N_2160);
nor U2958 (N_2958,N_2049,N_2064);
or U2959 (N_2959,N_2397,N_2369);
nor U2960 (N_2960,N_2408,N_2103);
or U2961 (N_2961,N_2461,N_2172);
nor U2962 (N_2962,N_2201,N_2396);
and U2963 (N_2963,N_2225,N_2262);
nand U2964 (N_2964,N_2476,N_2447);
nand U2965 (N_2965,N_2496,N_2158);
nand U2966 (N_2966,N_2402,N_2255);
xor U2967 (N_2967,N_2094,N_2372);
nand U2968 (N_2968,N_2173,N_2453);
and U2969 (N_2969,N_2407,N_2275);
or U2970 (N_2970,N_2440,N_2132);
nor U2971 (N_2971,N_2350,N_2306);
nor U2972 (N_2972,N_2270,N_2073);
and U2973 (N_2973,N_2116,N_2263);
nand U2974 (N_2974,N_2069,N_2244);
xor U2975 (N_2975,N_2207,N_2032);
and U2976 (N_2976,N_2328,N_2279);
nand U2977 (N_2977,N_2429,N_2030);
nand U2978 (N_2978,N_2155,N_2335);
nor U2979 (N_2979,N_2273,N_2116);
and U2980 (N_2980,N_2067,N_2406);
xnor U2981 (N_2981,N_2279,N_2046);
nand U2982 (N_2982,N_2419,N_2361);
and U2983 (N_2983,N_2064,N_2219);
or U2984 (N_2984,N_2471,N_2252);
nand U2985 (N_2985,N_2464,N_2148);
or U2986 (N_2986,N_2314,N_2430);
or U2987 (N_2987,N_2027,N_2399);
or U2988 (N_2988,N_2421,N_2090);
nor U2989 (N_2989,N_2286,N_2051);
or U2990 (N_2990,N_2125,N_2094);
xor U2991 (N_2991,N_2173,N_2062);
nor U2992 (N_2992,N_2457,N_2016);
and U2993 (N_2993,N_2006,N_2077);
and U2994 (N_2994,N_2062,N_2300);
or U2995 (N_2995,N_2296,N_2326);
nand U2996 (N_2996,N_2351,N_2419);
xnor U2997 (N_2997,N_2250,N_2191);
xor U2998 (N_2998,N_2427,N_2042);
xnor U2999 (N_2999,N_2243,N_2274);
nor U3000 (N_3000,N_2557,N_2564);
nand U3001 (N_3001,N_2537,N_2719);
nand U3002 (N_3002,N_2690,N_2895);
xor U3003 (N_3003,N_2643,N_2806);
nand U3004 (N_3004,N_2613,N_2575);
or U3005 (N_3005,N_2525,N_2515);
or U3006 (N_3006,N_2593,N_2636);
and U3007 (N_3007,N_2620,N_2845);
xor U3008 (N_3008,N_2664,N_2574);
nand U3009 (N_3009,N_2999,N_2792);
xnor U3010 (N_3010,N_2622,N_2508);
nor U3011 (N_3011,N_2814,N_2832);
xor U3012 (N_3012,N_2710,N_2542);
nor U3013 (N_3013,N_2762,N_2990);
or U3014 (N_3014,N_2998,N_2939);
or U3015 (N_3015,N_2700,N_2766);
and U3016 (N_3016,N_2619,N_2791);
and U3017 (N_3017,N_2790,N_2695);
nand U3018 (N_3018,N_2947,N_2943);
and U3019 (N_3019,N_2618,N_2549);
nor U3020 (N_3020,N_2875,N_2603);
nor U3021 (N_3021,N_2873,N_2740);
nor U3022 (N_3022,N_2698,N_2989);
or U3023 (N_3023,N_2800,N_2708);
nor U3024 (N_3024,N_2978,N_2993);
and U3025 (N_3025,N_2848,N_2819);
xnor U3026 (N_3026,N_2759,N_2547);
or U3027 (N_3027,N_2885,N_2551);
nor U3028 (N_3028,N_2519,N_2945);
or U3029 (N_3029,N_2808,N_2706);
xnor U3030 (N_3030,N_2920,N_2765);
nor U3031 (N_3031,N_2805,N_2602);
and U3032 (N_3032,N_2696,N_2611);
nand U3033 (N_3033,N_2995,N_2916);
or U3034 (N_3034,N_2768,N_2763);
xor U3035 (N_3035,N_2915,N_2859);
nor U3036 (N_3036,N_2975,N_2633);
nand U3037 (N_3037,N_2576,N_2968);
or U3038 (N_3038,N_2905,N_2862);
xnor U3039 (N_3039,N_2906,N_2579);
nor U3040 (N_3040,N_2642,N_2799);
xor U3041 (N_3041,N_2510,N_2834);
nand U3042 (N_3042,N_2926,N_2691);
xor U3043 (N_3043,N_2594,N_2645);
or U3044 (N_3044,N_2886,N_2986);
nand U3045 (N_3045,N_2894,N_2704);
and U3046 (N_3046,N_2849,N_2554);
nand U3047 (N_3047,N_2658,N_2528);
nor U3048 (N_3048,N_2601,N_2561);
nand U3049 (N_3049,N_2656,N_2617);
and U3050 (N_3050,N_2935,N_2948);
nand U3051 (N_3051,N_2648,N_2818);
xnor U3052 (N_3052,N_2566,N_2941);
or U3053 (N_3053,N_2864,N_2628);
or U3054 (N_3054,N_2683,N_2828);
and U3055 (N_3055,N_2898,N_2942);
and U3056 (N_3056,N_2946,N_2893);
nor U3057 (N_3057,N_2912,N_2932);
or U3058 (N_3058,N_2521,N_2785);
xor U3059 (N_3059,N_2727,N_2503);
or U3060 (N_3060,N_2937,N_2569);
or U3061 (N_3061,N_2964,N_2539);
xnor U3062 (N_3062,N_2773,N_2546);
and U3063 (N_3063,N_2797,N_2753);
nand U3064 (N_3064,N_2796,N_2505);
nor U3065 (N_3065,N_2694,N_2903);
and U3066 (N_3066,N_2841,N_2925);
nand U3067 (N_3067,N_2982,N_2723);
nor U3068 (N_3068,N_2588,N_2860);
xnor U3069 (N_3069,N_2803,N_2668);
and U3070 (N_3070,N_2777,N_2981);
nand U3071 (N_3071,N_2686,N_2702);
nand U3072 (N_3072,N_2843,N_2587);
xnor U3073 (N_3073,N_2517,N_2991);
or U3074 (N_3074,N_2746,N_2679);
nand U3075 (N_3075,N_2829,N_2764);
xnor U3076 (N_3076,N_2646,N_2928);
nor U3077 (N_3077,N_2623,N_2854);
and U3078 (N_3078,N_2688,N_2853);
xor U3079 (N_3079,N_2703,N_2598);
nor U3080 (N_3080,N_2751,N_2910);
nor U3081 (N_3081,N_2966,N_2626);
or U3082 (N_3082,N_2861,N_2568);
nand U3083 (N_3083,N_2541,N_2634);
xor U3084 (N_3084,N_2596,N_2522);
nand U3085 (N_3085,N_2584,N_2654);
and U3086 (N_3086,N_2835,N_2527);
nand U3087 (N_3087,N_2930,N_2996);
xor U3088 (N_3088,N_2863,N_2612);
nor U3089 (N_3089,N_2722,N_2673);
or U3090 (N_3090,N_2726,N_2555);
xnor U3091 (N_3091,N_2907,N_2504);
or U3092 (N_3092,N_2692,N_2846);
nand U3093 (N_3093,N_2507,N_2571);
or U3094 (N_3094,N_2578,N_2660);
nor U3095 (N_3095,N_2896,N_2544);
nor U3096 (N_3096,N_2630,N_2640);
nand U3097 (N_3097,N_2878,N_2724);
xor U3098 (N_3098,N_2540,N_2994);
and U3099 (N_3099,N_2889,N_2743);
or U3100 (N_3100,N_2592,N_2866);
or U3101 (N_3101,N_2731,N_2631);
xor U3102 (N_3102,N_2933,N_2810);
or U3103 (N_3103,N_2877,N_2625);
nand U3104 (N_3104,N_2938,N_2950);
nor U3105 (N_3105,N_2824,N_2872);
nand U3106 (N_3106,N_2816,N_2855);
or U3107 (N_3107,N_2830,N_2958);
or U3108 (N_3108,N_2616,N_2954);
nor U3109 (N_3109,N_2661,N_2513);
nand U3110 (N_3110,N_2684,N_2899);
xnor U3111 (N_3111,N_2957,N_2931);
nor U3112 (N_3112,N_2530,N_2599);
or U3113 (N_3113,N_2936,N_2783);
nor U3114 (N_3114,N_2586,N_2716);
nor U3115 (N_3115,N_2553,N_2718);
or U3116 (N_3116,N_2581,N_2880);
nor U3117 (N_3117,N_2883,N_2501);
or U3118 (N_3118,N_2637,N_2605);
nand U3119 (N_3119,N_2559,N_2770);
or U3120 (N_3120,N_2742,N_2614);
nand U3121 (N_3121,N_2961,N_2641);
and U3122 (N_3122,N_2715,N_2607);
nand U3123 (N_3123,N_2737,N_2729);
or U3124 (N_3124,N_2739,N_2621);
xor U3125 (N_3125,N_2988,N_2552);
or U3126 (N_3126,N_2831,N_2728);
xor U3127 (N_3127,N_2929,N_2717);
or U3128 (N_3128,N_2881,N_2562);
or U3129 (N_3129,N_2685,N_2672);
nand U3130 (N_3130,N_2965,N_2667);
nor U3131 (N_3131,N_2967,N_2744);
xnor U3132 (N_3132,N_2820,N_2591);
and U3133 (N_3133,N_2887,N_2655);
xnor U3134 (N_3134,N_2771,N_2865);
xnor U3135 (N_3135,N_2526,N_2992);
and U3136 (N_3136,N_2892,N_2535);
nor U3137 (N_3137,N_2748,N_2570);
or U3138 (N_3138,N_2651,N_2977);
and U3139 (N_3139,N_2709,N_2608);
nor U3140 (N_3140,N_2682,N_2548);
nand U3141 (N_3141,N_2678,N_2567);
and U3142 (N_3142,N_2844,N_2750);
xor U3143 (N_3143,N_2629,N_2523);
nor U3144 (N_3144,N_2639,N_2550);
nor U3145 (N_3145,N_2500,N_2680);
or U3146 (N_3146,N_2786,N_2997);
and U3147 (N_3147,N_2676,N_2725);
nor U3148 (N_3148,N_2879,N_2758);
xor U3149 (N_3149,N_2874,N_2852);
or U3150 (N_3150,N_2769,N_2867);
and U3151 (N_3151,N_2884,N_2840);
nor U3152 (N_3152,N_2781,N_2701);
or U3153 (N_3153,N_2520,N_2597);
nor U3154 (N_3154,N_2813,N_2595);
and U3155 (N_3155,N_2825,N_2534);
and U3156 (N_3156,N_2665,N_2610);
or U3157 (N_3157,N_2674,N_2775);
nand U3158 (N_3158,N_2924,N_2827);
or U3159 (N_3159,N_2757,N_2754);
and U3160 (N_3160,N_2801,N_2851);
and U3161 (N_3161,N_2952,N_2543);
nor U3162 (N_3162,N_2518,N_2669);
or U3163 (N_3163,N_2983,N_2802);
xor U3164 (N_3164,N_2735,N_2919);
nand U3165 (N_3165,N_2904,N_2921);
xnor U3166 (N_3166,N_2809,N_2798);
nor U3167 (N_3167,N_2767,N_2951);
nor U3168 (N_3168,N_2755,N_2511);
or U3169 (N_3169,N_2734,N_2638);
nor U3170 (N_3170,N_2745,N_2720);
nand U3171 (N_3171,N_2532,N_2782);
and U3172 (N_3172,N_2502,N_2940);
or U3173 (N_3173,N_2632,N_2826);
nand U3174 (N_3174,N_2652,N_2774);
nor U3175 (N_3175,N_2650,N_2589);
nor U3176 (N_3176,N_2838,N_2772);
xor U3177 (N_3177,N_2934,N_2707);
and U3178 (N_3178,N_2909,N_2624);
nor U3179 (N_3179,N_2897,N_2711);
nor U3180 (N_3180,N_2644,N_2822);
and U3181 (N_3181,N_2963,N_2856);
xnor U3182 (N_3182,N_2752,N_2516);
or U3183 (N_3183,N_2833,N_2927);
nand U3184 (N_3184,N_2647,N_2962);
xnor U3185 (N_3185,N_2615,N_2749);
and U3186 (N_3186,N_2657,N_2980);
or U3187 (N_3187,N_2563,N_2869);
and U3188 (N_3188,N_2776,N_2953);
nor U3189 (N_3189,N_2653,N_2914);
xnor U3190 (N_3190,N_2606,N_2839);
and U3191 (N_3191,N_2812,N_2736);
xnor U3192 (N_3192,N_2697,N_2705);
xor U3193 (N_3193,N_2713,N_2795);
or U3194 (N_3194,N_2604,N_2741);
and U3195 (N_3195,N_2891,N_2949);
nand U3196 (N_3196,N_2918,N_2807);
nand U3197 (N_3197,N_2693,N_2960);
nand U3198 (N_3198,N_2969,N_2956);
xor U3199 (N_3199,N_2804,N_2789);
and U3200 (N_3200,N_2794,N_2649);
nor U3201 (N_3201,N_2842,N_2738);
or U3202 (N_3202,N_2509,N_2681);
nand U3203 (N_3203,N_2900,N_2582);
nand U3204 (N_3204,N_2779,N_2712);
nor U3205 (N_3205,N_2821,N_2970);
and U3206 (N_3206,N_2868,N_2545);
nand U3207 (N_3207,N_2788,N_2922);
and U3208 (N_3208,N_2850,N_2882);
xnor U3209 (N_3209,N_2662,N_2780);
xnor U3210 (N_3210,N_2913,N_2627);
nor U3211 (N_3211,N_2565,N_2512);
xnor U3212 (N_3212,N_2815,N_2760);
nor U3213 (N_3213,N_2979,N_2955);
nand U3214 (N_3214,N_2529,N_2536);
nor U3215 (N_3215,N_2972,N_2663);
nor U3216 (N_3216,N_2971,N_2699);
nand U3217 (N_3217,N_2671,N_2747);
and U3218 (N_3218,N_2901,N_2847);
and U3219 (N_3219,N_2784,N_2659);
and U3220 (N_3220,N_2902,N_2556);
and U3221 (N_3221,N_2721,N_2560);
xnor U3222 (N_3222,N_2538,N_2666);
nand U3223 (N_3223,N_2573,N_2976);
and U3224 (N_3224,N_2572,N_2870);
xor U3225 (N_3225,N_2577,N_2590);
nor U3226 (N_3226,N_2635,N_2944);
xor U3227 (N_3227,N_2675,N_2973);
xnor U3228 (N_3228,N_2580,N_2778);
nor U3229 (N_3229,N_2817,N_2687);
xor U3230 (N_3230,N_2959,N_2524);
or U3231 (N_3231,N_2514,N_2670);
nor U3232 (N_3232,N_2793,N_2506);
nand U3233 (N_3233,N_2585,N_2890);
xnor U3234 (N_3234,N_2600,N_2689);
or U3235 (N_3235,N_2823,N_2531);
xnor U3236 (N_3236,N_2730,N_2677);
nand U3237 (N_3237,N_2609,N_2908);
and U3238 (N_3238,N_2917,N_2911);
xor U3239 (N_3239,N_2984,N_2533);
and U3240 (N_3240,N_2558,N_2923);
or U3241 (N_3241,N_2761,N_2811);
and U3242 (N_3242,N_2714,N_2837);
xor U3243 (N_3243,N_2888,N_2858);
xor U3244 (N_3244,N_2987,N_2857);
xor U3245 (N_3245,N_2732,N_2733);
nand U3246 (N_3246,N_2583,N_2974);
xnor U3247 (N_3247,N_2756,N_2836);
xnor U3248 (N_3248,N_2985,N_2876);
xnor U3249 (N_3249,N_2787,N_2871);
nor U3250 (N_3250,N_2888,N_2715);
nand U3251 (N_3251,N_2869,N_2612);
xor U3252 (N_3252,N_2868,N_2842);
nand U3253 (N_3253,N_2739,N_2721);
nand U3254 (N_3254,N_2882,N_2846);
nor U3255 (N_3255,N_2992,N_2523);
xnor U3256 (N_3256,N_2724,N_2624);
nor U3257 (N_3257,N_2951,N_2948);
or U3258 (N_3258,N_2566,N_2628);
or U3259 (N_3259,N_2671,N_2735);
and U3260 (N_3260,N_2982,N_2915);
nand U3261 (N_3261,N_2764,N_2577);
and U3262 (N_3262,N_2576,N_2794);
xor U3263 (N_3263,N_2905,N_2728);
xnor U3264 (N_3264,N_2580,N_2551);
or U3265 (N_3265,N_2835,N_2556);
or U3266 (N_3266,N_2706,N_2910);
nor U3267 (N_3267,N_2744,N_2809);
and U3268 (N_3268,N_2813,N_2882);
nor U3269 (N_3269,N_2992,N_2537);
and U3270 (N_3270,N_2670,N_2710);
xnor U3271 (N_3271,N_2518,N_2734);
or U3272 (N_3272,N_2676,N_2957);
xor U3273 (N_3273,N_2897,N_2720);
nor U3274 (N_3274,N_2800,N_2882);
xnor U3275 (N_3275,N_2788,N_2550);
nand U3276 (N_3276,N_2948,N_2812);
or U3277 (N_3277,N_2988,N_2779);
and U3278 (N_3278,N_2882,N_2638);
nor U3279 (N_3279,N_2897,N_2783);
xnor U3280 (N_3280,N_2918,N_2820);
and U3281 (N_3281,N_2904,N_2719);
xor U3282 (N_3282,N_2658,N_2674);
nand U3283 (N_3283,N_2756,N_2531);
or U3284 (N_3284,N_2968,N_2797);
and U3285 (N_3285,N_2556,N_2910);
or U3286 (N_3286,N_2774,N_2873);
xor U3287 (N_3287,N_2743,N_2649);
nor U3288 (N_3288,N_2809,N_2986);
xnor U3289 (N_3289,N_2532,N_2858);
nand U3290 (N_3290,N_2829,N_2760);
xor U3291 (N_3291,N_2981,N_2619);
nand U3292 (N_3292,N_2980,N_2843);
nand U3293 (N_3293,N_2884,N_2647);
and U3294 (N_3294,N_2526,N_2936);
and U3295 (N_3295,N_2540,N_2538);
nand U3296 (N_3296,N_2811,N_2710);
and U3297 (N_3297,N_2939,N_2802);
and U3298 (N_3298,N_2764,N_2732);
nand U3299 (N_3299,N_2770,N_2946);
nor U3300 (N_3300,N_2576,N_2809);
and U3301 (N_3301,N_2714,N_2925);
xnor U3302 (N_3302,N_2941,N_2617);
nand U3303 (N_3303,N_2803,N_2532);
xor U3304 (N_3304,N_2536,N_2624);
or U3305 (N_3305,N_2921,N_2872);
nor U3306 (N_3306,N_2588,N_2805);
nor U3307 (N_3307,N_2662,N_2989);
and U3308 (N_3308,N_2702,N_2730);
or U3309 (N_3309,N_2701,N_2657);
and U3310 (N_3310,N_2809,N_2690);
nand U3311 (N_3311,N_2846,N_2784);
nand U3312 (N_3312,N_2705,N_2741);
or U3313 (N_3313,N_2767,N_2781);
xnor U3314 (N_3314,N_2618,N_2676);
and U3315 (N_3315,N_2675,N_2828);
nand U3316 (N_3316,N_2721,N_2965);
or U3317 (N_3317,N_2677,N_2830);
or U3318 (N_3318,N_2712,N_2792);
xor U3319 (N_3319,N_2534,N_2514);
or U3320 (N_3320,N_2702,N_2583);
or U3321 (N_3321,N_2885,N_2685);
and U3322 (N_3322,N_2978,N_2595);
and U3323 (N_3323,N_2508,N_2962);
xor U3324 (N_3324,N_2991,N_2555);
nor U3325 (N_3325,N_2981,N_2552);
nand U3326 (N_3326,N_2875,N_2731);
nand U3327 (N_3327,N_2893,N_2591);
nand U3328 (N_3328,N_2651,N_2554);
xnor U3329 (N_3329,N_2758,N_2732);
xor U3330 (N_3330,N_2895,N_2510);
nand U3331 (N_3331,N_2790,N_2950);
nand U3332 (N_3332,N_2871,N_2975);
and U3333 (N_3333,N_2988,N_2810);
or U3334 (N_3334,N_2834,N_2748);
nand U3335 (N_3335,N_2790,N_2975);
and U3336 (N_3336,N_2513,N_2858);
nor U3337 (N_3337,N_2666,N_2584);
or U3338 (N_3338,N_2610,N_2584);
nand U3339 (N_3339,N_2877,N_2977);
nor U3340 (N_3340,N_2682,N_2516);
and U3341 (N_3341,N_2706,N_2919);
xor U3342 (N_3342,N_2932,N_2867);
xor U3343 (N_3343,N_2919,N_2957);
nor U3344 (N_3344,N_2530,N_2990);
nor U3345 (N_3345,N_2966,N_2552);
xor U3346 (N_3346,N_2530,N_2709);
or U3347 (N_3347,N_2581,N_2507);
nor U3348 (N_3348,N_2520,N_2910);
or U3349 (N_3349,N_2833,N_2809);
or U3350 (N_3350,N_2681,N_2666);
xor U3351 (N_3351,N_2979,N_2670);
and U3352 (N_3352,N_2762,N_2712);
and U3353 (N_3353,N_2502,N_2919);
and U3354 (N_3354,N_2795,N_2941);
nor U3355 (N_3355,N_2686,N_2953);
nand U3356 (N_3356,N_2836,N_2935);
or U3357 (N_3357,N_2778,N_2898);
nor U3358 (N_3358,N_2794,N_2614);
nor U3359 (N_3359,N_2992,N_2572);
xor U3360 (N_3360,N_2561,N_2576);
xor U3361 (N_3361,N_2611,N_2844);
and U3362 (N_3362,N_2945,N_2918);
or U3363 (N_3363,N_2662,N_2733);
and U3364 (N_3364,N_2934,N_2684);
or U3365 (N_3365,N_2941,N_2903);
nand U3366 (N_3366,N_2905,N_2626);
xor U3367 (N_3367,N_2855,N_2515);
and U3368 (N_3368,N_2503,N_2785);
and U3369 (N_3369,N_2556,N_2904);
nand U3370 (N_3370,N_2562,N_2611);
and U3371 (N_3371,N_2840,N_2999);
and U3372 (N_3372,N_2760,N_2677);
nand U3373 (N_3373,N_2626,N_2784);
and U3374 (N_3374,N_2593,N_2612);
nor U3375 (N_3375,N_2511,N_2817);
or U3376 (N_3376,N_2754,N_2665);
nor U3377 (N_3377,N_2907,N_2916);
xnor U3378 (N_3378,N_2870,N_2737);
or U3379 (N_3379,N_2744,N_2826);
and U3380 (N_3380,N_2502,N_2908);
and U3381 (N_3381,N_2802,N_2532);
nor U3382 (N_3382,N_2938,N_2886);
nor U3383 (N_3383,N_2562,N_2742);
and U3384 (N_3384,N_2815,N_2507);
or U3385 (N_3385,N_2602,N_2758);
or U3386 (N_3386,N_2557,N_2762);
nand U3387 (N_3387,N_2702,N_2817);
xor U3388 (N_3388,N_2877,N_2663);
nor U3389 (N_3389,N_2754,N_2740);
xor U3390 (N_3390,N_2736,N_2543);
or U3391 (N_3391,N_2924,N_2616);
xor U3392 (N_3392,N_2940,N_2676);
xnor U3393 (N_3393,N_2528,N_2569);
nand U3394 (N_3394,N_2836,N_2830);
nand U3395 (N_3395,N_2759,N_2751);
nand U3396 (N_3396,N_2593,N_2519);
nand U3397 (N_3397,N_2971,N_2945);
and U3398 (N_3398,N_2855,N_2912);
or U3399 (N_3399,N_2928,N_2774);
or U3400 (N_3400,N_2743,N_2664);
nor U3401 (N_3401,N_2827,N_2642);
or U3402 (N_3402,N_2661,N_2949);
and U3403 (N_3403,N_2786,N_2907);
nand U3404 (N_3404,N_2502,N_2619);
nor U3405 (N_3405,N_2587,N_2854);
and U3406 (N_3406,N_2864,N_2949);
xor U3407 (N_3407,N_2634,N_2747);
xnor U3408 (N_3408,N_2721,N_2613);
or U3409 (N_3409,N_2873,N_2962);
and U3410 (N_3410,N_2647,N_2934);
nor U3411 (N_3411,N_2702,N_2774);
nand U3412 (N_3412,N_2834,N_2932);
or U3413 (N_3413,N_2653,N_2810);
nand U3414 (N_3414,N_2526,N_2721);
or U3415 (N_3415,N_2767,N_2731);
nor U3416 (N_3416,N_2997,N_2504);
nand U3417 (N_3417,N_2807,N_2714);
and U3418 (N_3418,N_2939,N_2923);
or U3419 (N_3419,N_2977,N_2676);
and U3420 (N_3420,N_2704,N_2904);
nand U3421 (N_3421,N_2607,N_2842);
xor U3422 (N_3422,N_2944,N_2710);
and U3423 (N_3423,N_2878,N_2564);
or U3424 (N_3424,N_2790,N_2559);
nand U3425 (N_3425,N_2681,N_2665);
nand U3426 (N_3426,N_2726,N_2874);
xor U3427 (N_3427,N_2667,N_2889);
or U3428 (N_3428,N_2938,N_2519);
nand U3429 (N_3429,N_2995,N_2521);
xnor U3430 (N_3430,N_2597,N_2796);
or U3431 (N_3431,N_2957,N_2529);
and U3432 (N_3432,N_2971,N_2969);
xnor U3433 (N_3433,N_2853,N_2896);
and U3434 (N_3434,N_2653,N_2589);
and U3435 (N_3435,N_2953,N_2813);
and U3436 (N_3436,N_2577,N_2805);
xnor U3437 (N_3437,N_2723,N_2913);
nand U3438 (N_3438,N_2725,N_2520);
and U3439 (N_3439,N_2818,N_2641);
or U3440 (N_3440,N_2997,N_2946);
and U3441 (N_3441,N_2923,N_2815);
nand U3442 (N_3442,N_2896,N_2760);
or U3443 (N_3443,N_2726,N_2714);
or U3444 (N_3444,N_2538,N_2787);
nand U3445 (N_3445,N_2867,N_2911);
xor U3446 (N_3446,N_2871,N_2563);
nand U3447 (N_3447,N_2519,N_2892);
and U3448 (N_3448,N_2841,N_2647);
nor U3449 (N_3449,N_2778,N_2653);
and U3450 (N_3450,N_2997,N_2867);
and U3451 (N_3451,N_2914,N_2779);
nor U3452 (N_3452,N_2999,N_2516);
and U3453 (N_3453,N_2517,N_2527);
nand U3454 (N_3454,N_2766,N_2921);
xor U3455 (N_3455,N_2767,N_2904);
and U3456 (N_3456,N_2961,N_2648);
nand U3457 (N_3457,N_2523,N_2564);
nand U3458 (N_3458,N_2970,N_2938);
xnor U3459 (N_3459,N_2928,N_2923);
and U3460 (N_3460,N_2689,N_2948);
or U3461 (N_3461,N_2741,N_2998);
nand U3462 (N_3462,N_2639,N_2807);
xor U3463 (N_3463,N_2871,N_2795);
nand U3464 (N_3464,N_2521,N_2741);
xor U3465 (N_3465,N_2848,N_2993);
and U3466 (N_3466,N_2861,N_2560);
nand U3467 (N_3467,N_2595,N_2880);
or U3468 (N_3468,N_2642,N_2793);
or U3469 (N_3469,N_2643,N_2815);
xor U3470 (N_3470,N_2812,N_2708);
nor U3471 (N_3471,N_2783,N_2618);
nor U3472 (N_3472,N_2641,N_2957);
or U3473 (N_3473,N_2696,N_2783);
nand U3474 (N_3474,N_2972,N_2616);
nand U3475 (N_3475,N_2916,N_2621);
and U3476 (N_3476,N_2871,N_2799);
xor U3477 (N_3477,N_2508,N_2902);
or U3478 (N_3478,N_2666,N_2754);
nand U3479 (N_3479,N_2880,N_2767);
nor U3480 (N_3480,N_2723,N_2726);
nand U3481 (N_3481,N_2656,N_2644);
and U3482 (N_3482,N_2548,N_2571);
nor U3483 (N_3483,N_2638,N_2676);
or U3484 (N_3484,N_2554,N_2858);
xnor U3485 (N_3485,N_2848,N_2932);
or U3486 (N_3486,N_2776,N_2565);
and U3487 (N_3487,N_2708,N_2518);
xnor U3488 (N_3488,N_2914,N_2648);
nand U3489 (N_3489,N_2532,N_2655);
nand U3490 (N_3490,N_2831,N_2993);
or U3491 (N_3491,N_2661,N_2583);
or U3492 (N_3492,N_2525,N_2734);
and U3493 (N_3493,N_2771,N_2855);
and U3494 (N_3494,N_2531,N_2726);
and U3495 (N_3495,N_2924,N_2629);
nand U3496 (N_3496,N_2884,N_2598);
nand U3497 (N_3497,N_2564,N_2875);
xnor U3498 (N_3498,N_2991,N_2795);
and U3499 (N_3499,N_2806,N_2768);
and U3500 (N_3500,N_3137,N_3274);
nand U3501 (N_3501,N_3125,N_3399);
and U3502 (N_3502,N_3447,N_3465);
nor U3503 (N_3503,N_3169,N_3355);
and U3504 (N_3504,N_3103,N_3064);
and U3505 (N_3505,N_3461,N_3278);
nor U3506 (N_3506,N_3413,N_3194);
and U3507 (N_3507,N_3146,N_3388);
xor U3508 (N_3508,N_3037,N_3150);
or U3509 (N_3509,N_3183,N_3069);
nor U3510 (N_3510,N_3006,N_3121);
xor U3511 (N_3511,N_3029,N_3260);
and U3512 (N_3512,N_3406,N_3055);
xnor U3513 (N_3513,N_3206,N_3249);
nor U3514 (N_3514,N_3191,N_3483);
or U3515 (N_3515,N_3400,N_3306);
nor U3516 (N_3516,N_3396,N_3273);
nor U3517 (N_3517,N_3107,N_3085);
and U3518 (N_3518,N_3386,N_3299);
and U3519 (N_3519,N_3240,N_3032);
and U3520 (N_3520,N_3181,N_3209);
and U3521 (N_3521,N_3226,N_3297);
xor U3522 (N_3522,N_3171,N_3197);
nand U3523 (N_3523,N_3432,N_3418);
nand U3524 (N_3524,N_3268,N_3324);
or U3525 (N_3525,N_3140,N_3459);
or U3526 (N_3526,N_3011,N_3120);
nor U3527 (N_3527,N_3389,N_3426);
xnor U3528 (N_3528,N_3397,N_3127);
nand U3529 (N_3529,N_3437,N_3008);
and U3530 (N_3530,N_3002,N_3091);
nor U3531 (N_3531,N_3155,N_3039);
xor U3532 (N_3532,N_3026,N_3354);
xnor U3533 (N_3533,N_3205,N_3452);
nor U3534 (N_3534,N_3336,N_3250);
or U3535 (N_3535,N_3367,N_3499);
and U3536 (N_3536,N_3112,N_3025);
xnor U3537 (N_3537,N_3496,N_3410);
nor U3538 (N_3538,N_3438,N_3267);
xnor U3539 (N_3539,N_3325,N_3263);
and U3540 (N_3540,N_3247,N_3233);
or U3541 (N_3541,N_3288,N_3356);
and U3542 (N_3542,N_3391,N_3086);
and U3543 (N_3543,N_3427,N_3214);
nand U3544 (N_3544,N_3070,N_3001);
xnor U3545 (N_3545,N_3184,N_3244);
xnor U3546 (N_3546,N_3476,N_3318);
nand U3547 (N_3547,N_3423,N_3298);
nor U3548 (N_3548,N_3380,N_3445);
nand U3549 (N_3549,N_3163,N_3373);
nor U3550 (N_3550,N_3450,N_3072);
and U3551 (N_3551,N_3262,N_3043);
nand U3552 (N_3552,N_3036,N_3007);
nor U3553 (N_3553,N_3302,N_3379);
nand U3554 (N_3554,N_3145,N_3421);
xnor U3555 (N_3555,N_3222,N_3093);
or U3556 (N_3556,N_3168,N_3265);
nor U3557 (N_3557,N_3467,N_3353);
and U3558 (N_3558,N_3454,N_3416);
nand U3559 (N_3559,N_3123,N_3016);
nor U3560 (N_3560,N_3409,N_3160);
or U3561 (N_3561,N_3051,N_3023);
nand U3562 (N_3562,N_3075,N_3176);
and U3563 (N_3563,N_3328,N_3308);
and U3564 (N_3564,N_3449,N_3287);
or U3565 (N_3565,N_3330,N_3204);
and U3566 (N_3566,N_3471,N_3381);
xor U3567 (N_3567,N_3084,N_3082);
or U3568 (N_3568,N_3132,N_3193);
or U3569 (N_3569,N_3407,N_3434);
nand U3570 (N_3570,N_3243,N_3117);
and U3571 (N_3571,N_3192,N_3462);
xnor U3572 (N_3572,N_3048,N_3314);
nand U3573 (N_3573,N_3404,N_3178);
xor U3574 (N_3574,N_3362,N_3215);
xor U3575 (N_3575,N_3478,N_3100);
xor U3576 (N_3576,N_3188,N_3309);
or U3577 (N_3577,N_3174,N_3014);
nor U3578 (N_3578,N_3022,N_3147);
nor U3579 (N_3579,N_3165,N_3073);
nor U3580 (N_3580,N_3216,N_3245);
nand U3581 (N_3581,N_3316,N_3019);
or U3582 (N_3582,N_3370,N_3482);
or U3583 (N_3583,N_3124,N_3097);
nand U3584 (N_3584,N_3119,N_3235);
and U3585 (N_3585,N_3207,N_3469);
nor U3586 (N_3586,N_3394,N_3149);
and U3587 (N_3587,N_3345,N_3106);
nor U3588 (N_3588,N_3387,N_3063);
xnor U3589 (N_3589,N_3311,N_3393);
or U3590 (N_3590,N_3295,N_3315);
nor U3591 (N_3591,N_3472,N_3201);
nand U3592 (N_3592,N_3138,N_3257);
nor U3593 (N_3593,N_3228,N_3313);
nand U3594 (N_3594,N_3027,N_3322);
xor U3595 (N_3595,N_3161,N_3219);
or U3596 (N_3596,N_3275,N_3232);
nor U3597 (N_3597,N_3195,N_3470);
xnor U3598 (N_3598,N_3096,N_3111);
nor U3599 (N_3599,N_3346,N_3211);
or U3600 (N_3600,N_3101,N_3429);
or U3601 (N_3601,N_3110,N_3420);
and U3602 (N_3602,N_3196,N_3083);
xor U3603 (N_3603,N_3365,N_3301);
nor U3604 (N_3604,N_3357,N_3241);
nor U3605 (N_3605,N_3276,N_3337);
or U3606 (N_3606,N_3326,N_3053);
and U3607 (N_3607,N_3464,N_3280);
and U3608 (N_3608,N_3237,N_3102);
nor U3609 (N_3609,N_3347,N_3170);
or U3610 (N_3610,N_3332,N_3348);
nand U3611 (N_3611,N_3341,N_3208);
nand U3612 (N_3612,N_3139,N_3225);
or U3613 (N_3613,N_3492,N_3238);
nand U3614 (N_3614,N_3485,N_3480);
or U3615 (N_3615,N_3272,N_3058);
nand U3616 (N_3616,N_3408,N_3142);
or U3617 (N_3617,N_3143,N_3003);
and U3618 (N_3618,N_3252,N_3259);
xor U3619 (N_3619,N_3078,N_3378);
nand U3620 (N_3620,N_3024,N_3136);
and U3621 (N_3621,N_3497,N_3079);
or U3622 (N_3622,N_3246,N_3071);
nor U3623 (N_3623,N_3342,N_3200);
and U3624 (N_3624,N_3494,N_3360);
and U3625 (N_3625,N_3431,N_3256);
nor U3626 (N_3626,N_3258,N_3368);
nand U3627 (N_3627,N_3475,N_3220);
and U3628 (N_3628,N_3335,N_3374);
and U3629 (N_3629,N_3261,N_3359);
xor U3630 (N_3630,N_3457,N_3131);
and U3631 (N_3631,N_3430,N_3021);
and U3632 (N_3632,N_3187,N_3004);
nand U3633 (N_3633,N_3364,N_3126);
or U3634 (N_3634,N_3153,N_3118);
or U3635 (N_3635,N_3080,N_3433);
and U3636 (N_3636,N_3327,N_3044);
and U3637 (N_3637,N_3415,N_3034);
nor U3638 (N_3638,N_3444,N_3040);
xnor U3639 (N_3639,N_3304,N_3264);
nand U3640 (N_3640,N_3210,N_3054);
nor U3641 (N_3641,N_3479,N_3334);
and U3642 (N_3642,N_3285,N_3015);
or U3643 (N_3643,N_3329,N_3066);
nor U3644 (N_3644,N_3164,N_3283);
nand U3645 (N_3645,N_3375,N_3369);
or U3646 (N_3646,N_3092,N_3134);
nor U3647 (N_3647,N_3213,N_3493);
nand U3648 (N_3648,N_3189,N_3062);
or U3649 (N_3649,N_3251,N_3130);
nor U3650 (N_3650,N_3277,N_3223);
or U3651 (N_3651,N_3012,N_3435);
xor U3652 (N_3652,N_3151,N_3221);
xor U3653 (N_3653,N_3489,N_3144);
or U3654 (N_3654,N_3202,N_3371);
xnor U3655 (N_3655,N_3377,N_3010);
or U3656 (N_3656,N_3116,N_3095);
and U3657 (N_3657,N_3333,N_3060);
nor U3658 (N_3658,N_3088,N_3390);
nor U3659 (N_3659,N_3033,N_3089);
nor U3660 (N_3660,N_3401,N_3271);
nand U3661 (N_3661,N_3372,N_3236);
nor U3662 (N_3662,N_3028,N_3230);
or U3663 (N_3663,N_3425,N_3321);
and U3664 (N_3664,N_3167,N_3081);
nand U3665 (N_3665,N_3133,N_3339);
nor U3666 (N_3666,N_3382,N_3490);
or U3667 (N_3667,N_3203,N_3292);
and U3668 (N_3668,N_3185,N_3474);
or U3669 (N_3669,N_3477,N_3175);
or U3670 (N_3670,N_3254,N_3281);
xnor U3671 (N_3671,N_3229,N_3045);
and U3672 (N_3672,N_3255,N_3152);
nor U3673 (N_3673,N_3279,N_3487);
or U3674 (N_3674,N_3242,N_3340);
or U3675 (N_3675,N_3224,N_3128);
nor U3676 (N_3676,N_3158,N_3439);
nor U3677 (N_3677,N_3234,N_3041);
and U3678 (N_3678,N_3031,N_3108);
nand U3679 (N_3679,N_3186,N_3156);
nor U3680 (N_3680,N_3046,N_3488);
nand U3681 (N_3681,N_3239,N_3392);
xnor U3682 (N_3682,N_3384,N_3269);
nand U3683 (N_3683,N_3344,N_3105);
and U3684 (N_3684,N_3293,N_3148);
nor U3685 (N_3685,N_3227,N_3052);
xor U3686 (N_3686,N_3351,N_3061);
or U3687 (N_3687,N_3486,N_3198);
nor U3688 (N_3688,N_3320,N_3312);
xnor U3689 (N_3689,N_3173,N_3441);
nor U3690 (N_3690,N_3451,N_3074);
or U3691 (N_3691,N_3113,N_3436);
nand U3692 (N_3692,N_3468,N_3350);
nand U3693 (N_3693,N_3484,N_3177);
or U3694 (N_3694,N_3253,N_3352);
xnor U3695 (N_3695,N_3453,N_3491);
nor U3696 (N_3696,N_3319,N_3296);
or U3697 (N_3697,N_3422,N_3018);
nor U3698 (N_3698,N_3218,N_3017);
xnor U3699 (N_3699,N_3307,N_3403);
xnor U3700 (N_3700,N_3109,N_3419);
xnor U3701 (N_3701,N_3428,N_3122);
nand U3702 (N_3702,N_3424,N_3310);
nand U3703 (N_3703,N_3248,N_3231);
or U3704 (N_3704,N_3294,N_3005);
and U3705 (N_3705,N_3172,N_3035);
and U3706 (N_3706,N_3440,N_3498);
nor U3707 (N_3707,N_3456,N_3038);
nor U3708 (N_3708,N_3159,N_3115);
and U3709 (N_3709,N_3135,N_3000);
xor U3710 (N_3710,N_3349,N_3129);
xnor U3711 (N_3711,N_3300,N_3443);
nor U3712 (N_3712,N_3303,N_3442);
nand U3713 (N_3713,N_3455,N_3282);
xnor U3714 (N_3714,N_3317,N_3463);
nor U3715 (N_3715,N_3460,N_3065);
or U3716 (N_3716,N_3289,N_3057);
or U3717 (N_3717,N_3473,N_3290);
nand U3718 (N_3718,N_3090,N_3182);
or U3719 (N_3719,N_3376,N_3411);
or U3720 (N_3720,N_3098,N_3266);
nor U3721 (N_3721,N_3076,N_3059);
or U3722 (N_3722,N_3323,N_3395);
or U3723 (N_3723,N_3009,N_3466);
or U3724 (N_3724,N_3067,N_3481);
and U3725 (N_3725,N_3270,N_3154);
and U3726 (N_3726,N_3361,N_3331);
xnor U3727 (N_3727,N_3383,N_3343);
xnor U3728 (N_3728,N_3042,N_3286);
and U3729 (N_3729,N_3385,N_3077);
nand U3730 (N_3730,N_3458,N_3166);
nor U3731 (N_3731,N_3448,N_3414);
nor U3732 (N_3732,N_3020,N_3114);
xor U3733 (N_3733,N_3087,N_3217);
or U3734 (N_3734,N_3358,N_3446);
xnor U3735 (N_3735,N_3099,N_3284);
nor U3736 (N_3736,N_3398,N_3363);
and U3737 (N_3737,N_3050,N_3180);
and U3738 (N_3738,N_3013,N_3405);
and U3739 (N_3739,N_3104,N_3291);
nand U3740 (N_3740,N_3495,N_3049);
and U3741 (N_3741,N_3199,N_3212);
xor U3742 (N_3742,N_3162,N_3305);
xor U3743 (N_3743,N_3338,N_3190);
nor U3744 (N_3744,N_3157,N_3047);
nor U3745 (N_3745,N_3366,N_3056);
or U3746 (N_3746,N_3141,N_3412);
nor U3747 (N_3747,N_3179,N_3402);
or U3748 (N_3748,N_3417,N_3094);
or U3749 (N_3749,N_3030,N_3068);
xnor U3750 (N_3750,N_3310,N_3355);
nand U3751 (N_3751,N_3008,N_3095);
or U3752 (N_3752,N_3453,N_3219);
nor U3753 (N_3753,N_3467,N_3465);
xor U3754 (N_3754,N_3286,N_3429);
or U3755 (N_3755,N_3479,N_3267);
or U3756 (N_3756,N_3332,N_3032);
or U3757 (N_3757,N_3077,N_3043);
nand U3758 (N_3758,N_3411,N_3436);
nor U3759 (N_3759,N_3451,N_3003);
nand U3760 (N_3760,N_3110,N_3318);
or U3761 (N_3761,N_3124,N_3164);
nand U3762 (N_3762,N_3089,N_3248);
and U3763 (N_3763,N_3337,N_3202);
nor U3764 (N_3764,N_3072,N_3336);
nand U3765 (N_3765,N_3172,N_3124);
or U3766 (N_3766,N_3485,N_3137);
and U3767 (N_3767,N_3037,N_3342);
nor U3768 (N_3768,N_3290,N_3394);
xnor U3769 (N_3769,N_3063,N_3374);
or U3770 (N_3770,N_3496,N_3414);
or U3771 (N_3771,N_3014,N_3039);
or U3772 (N_3772,N_3416,N_3055);
xor U3773 (N_3773,N_3401,N_3446);
nand U3774 (N_3774,N_3142,N_3394);
nand U3775 (N_3775,N_3299,N_3484);
nand U3776 (N_3776,N_3073,N_3351);
or U3777 (N_3777,N_3408,N_3187);
or U3778 (N_3778,N_3446,N_3444);
xnor U3779 (N_3779,N_3310,N_3136);
nand U3780 (N_3780,N_3074,N_3137);
xnor U3781 (N_3781,N_3405,N_3275);
nand U3782 (N_3782,N_3213,N_3210);
nor U3783 (N_3783,N_3145,N_3428);
xor U3784 (N_3784,N_3204,N_3034);
and U3785 (N_3785,N_3233,N_3256);
nand U3786 (N_3786,N_3221,N_3028);
and U3787 (N_3787,N_3319,N_3487);
nor U3788 (N_3788,N_3134,N_3169);
and U3789 (N_3789,N_3191,N_3195);
xnor U3790 (N_3790,N_3229,N_3278);
nor U3791 (N_3791,N_3419,N_3269);
xnor U3792 (N_3792,N_3081,N_3242);
nor U3793 (N_3793,N_3287,N_3091);
and U3794 (N_3794,N_3042,N_3490);
or U3795 (N_3795,N_3204,N_3108);
and U3796 (N_3796,N_3411,N_3090);
xor U3797 (N_3797,N_3482,N_3456);
and U3798 (N_3798,N_3419,N_3237);
nand U3799 (N_3799,N_3314,N_3253);
xor U3800 (N_3800,N_3069,N_3196);
and U3801 (N_3801,N_3074,N_3054);
nor U3802 (N_3802,N_3411,N_3276);
nand U3803 (N_3803,N_3363,N_3383);
and U3804 (N_3804,N_3258,N_3290);
nand U3805 (N_3805,N_3188,N_3073);
nand U3806 (N_3806,N_3357,N_3403);
and U3807 (N_3807,N_3201,N_3272);
xor U3808 (N_3808,N_3077,N_3490);
xor U3809 (N_3809,N_3129,N_3161);
xor U3810 (N_3810,N_3082,N_3031);
nor U3811 (N_3811,N_3211,N_3246);
xor U3812 (N_3812,N_3220,N_3049);
xor U3813 (N_3813,N_3319,N_3403);
xor U3814 (N_3814,N_3381,N_3087);
or U3815 (N_3815,N_3279,N_3108);
and U3816 (N_3816,N_3167,N_3216);
nor U3817 (N_3817,N_3034,N_3390);
and U3818 (N_3818,N_3321,N_3455);
and U3819 (N_3819,N_3108,N_3366);
nand U3820 (N_3820,N_3056,N_3169);
nand U3821 (N_3821,N_3225,N_3020);
nand U3822 (N_3822,N_3162,N_3303);
and U3823 (N_3823,N_3291,N_3449);
nand U3824 (N_3824,N_3037,N_3343);
nor U3825 (N_3825,N_3435,N_3282);
nor U3826 (N_3826,N_3410,N_3257);
nor U3827 (N_3827,N_3177,N_3000);
or U3828 (N_3828,N_3086,N_3311);
xor U3829 (N_3829,N_3226,N_3368);
xnor U3830 (N_3830,N_3125,N_3474);
and U3831 (N_3831,N_3337,N_3169);
xor U3832 (N_3832,N_3031,N_3042);
and U3833 (N_3833,N_3190,N_3375);
and U3834 (N_3834,N_3479,N_3109);
xor U3835 (N_3835,N_3103,N_3248);
or U3836 (N_3836,N_3418,N_3008);
nor U3837 (N_3837,N_3086,N_3255);
nor U3838 (N_3838,N_3306,N_3115);
and U3839 (N_3839,N_3441,N_3445);
xnor U3840 (N_3840,N_3176,N_3047);
nand U3841 (N_3841,N_3057,N_3243);
nand U3842 (N_3842,N_3312,N_3122);
nand U3843 (N_3843,N_3460,N_3351);
xor U3844 (N_3844,N_3093,N_3464);
or U3845 (N_3845,N_3217,N_3213);
or U3846 (N_3846,N_3110,N_3050);
nor U3847 (N_3847,N_3349,N_3451);
and U3848 (N_3848,N_3439,N_3232);
nor U3849 (N_3849,N_3156,N_3437);
xor U3850 (N_3850,N_3034,N_3490);
nand U3851 (N_3851,N_3238,N_3212);
nand U3852 (N_3852,N_3453,N_3086);
nor U3853 (N_3853,N_3424,N_3491);
or U3854 (N_3854,N_3123,N_3084);
xor U3855 (N_3855,N_3400,N_3282);
and U3856 (N_3856,N_3029,N_3182);
nand U3857 (N_3857,N_3160,N_3256);
xnor U3858 (N_3858,N_3104,N_3432);
nand U3859 (N_3859,N_3100,N_3132);
xor U3860 (N_3860,N_3314,N_3206);
nor U3861 (N_3861,N_3092,N_3198);
and U3862 (N_3862,N_3257,N_3277);
and U3863 (N_3863,N_3222,N_3278);
xor U3864 (N_3864,N_3177,N_3019);
or U3865 (N_3865,N_3371,N_3446);
and U3866 (N_3866,N_3332,N_3008);
nand U3867 (N_3867,N_3494,N_3353);
nor U3868 (N_3868,N_3393,N_3046);
or U3869 (N_3869,N_3454,N_3071);
nand U3870 (N_3870,N_3211,N_3204);
and U3871 (N_3871,N_3003,N_3063);
and U3872 (N_3872,N_3103,N_3304);
nand U3873 (N_3873,N_3234,N_3276);
xnor U3874 (N_3874,N_3304,N_3038);
and U3875 (N_3875,N_3107,N_3295);
nor U3876 (N_3876,N_3453,N_3445);
nand U3877 (N_3877,N_3428,N_3079);
nand U3878 (N_3878,N_3303,N_3489);
nand U3879 (N_3879,N_3222,N_3014);
or U3880 (N_3880,N_3106,N_3396);
and U3881 (N_3881,N_3199,N_3237);
and U3882 (N_3882,N_3044,N_3496);
or U3883 (N_3883,N_3310,N_3043);
xnor U3884 (N_3884,N_3111,N_3066);
nor U3885 (N_3885,N_3456,N_3275);
nand U3886 (N_3886,N_3337,N_3458);
or U3887 (N_3887,N_3134,N_3085);
and U3888 (N_3888,N_3183,N_3405);
or U3889 (N_3889,N_3053,N_3152);
nand U3890 (N_3890,N_3256,N_3011);
xnor U3891 (N_3891,N_3272,N_3468);
nor U3892 (N_3892,N_3221,N_3139);
or U3893 (N_3893,N_3378,N_3254);
and U3894 (N_3894,N_3268,N_3113);
nor U3895 (N_3895,N_3086,N_3010);
nand U3896 (N_3896,N_3445,N_3432);
and U3897 (N_3897,N_3214,N_3228);
or U3898 (N_3898,N_3041,N_3186);
nand U3899 (N_3899,N_3116,N_3225);
and U3900 (N_3900,N_3273,N_3421);
nor U3901 (N_3901,N_3324,N_3149);
nand U3902 (N_3902,N_3076,N_3239);
or U3903 (N_3903,N_3363,N_3082);
xnor U3904 (N_3904,N_3035,N_3138);
and U3905 (N_3905,N_3089,N_3439);
nor U3906 (N_3906,N_3040,N_3352);
nor U3907 (N_3907,N_3138,N_3156);
xor U3908 (N_3908,N_3388,N_3227);
nand U3909 (N_3909,N_3049,N_3318);
nand U3910 (N_3910,N_3063,N_3144);
xor U3911 (N_3911,N_3493,N_3347);
nor U3912 (N_3912,N_3477,N_3118);
nand U3913 (N_3913,N_3144,N_3201);
xnor U3914 (N_3914,N_3102,N_3427);
and U3915 (N_3915,N_3016,N_3414);
nand U3916 (N_3916,N_3357,N_3339);
nand U3917 (N_3917,N_3300,N_3048);
and U3918 (N_3918,N_3303,N_3041);
nand U3919 (N_3919,N_3230,N_3093);
and U3920 (N_3920,N_3486,N_3153);
nor U3921 (N_3921,N_3273,N_3409);
or U3922 (N_3922,N_3329,N_3044);
and U3923 (N_3923,N_3267,N_3292);
or U3924 (N_3924,N_3088,N_3471);
nand U3925 (N_3925,N_3031,N_3133);
xnor U3926 (N_3926,N_3093,N_3308);
nor U3927 (N_3927,N_3323,N_3320);
or U3928 (N_3928,N_3405,N_3000);
nand U3929 (N_3929,N_3163,N_3093);
or U3930 (N_3930,N_3042,N_3096);
and U3931 (N_3931,N_3058,N_3200);
nand U3932 (N_3932,N_3075,N_3135);
and U3933 (N_3933,N_3045,N_3075);
or U3934 (N_3934,N_3141,N_3231);
nor U3935 (N_3935,N_3058,N_3275);
or U3936 (N_3936,N_3131,N_3222);
nor U3937 (N_3937,N_3221,N_3170);
nand U3938 (N_3938,N_3170,N_3027);
or U3939 (N_3939,N_3301,N_3013);
nand U3940 (N_3940,N_3327,N_3112);
and U3941 (N_3941,N_3078,N_3413);
nand U3942 (N_3942,N_3376,N_3096);
or U3943 (N_3943,N_3489,N_3296);
nor U3944 (N_3944,N_3160,N_3203);
nand U3945 (N_3945,N_3475,N_3251);
xor U3946 (N_3946,N_3048,N_3369);
or U3947 (N_3947,N_3367,N_3232);
nand U3948 (N_3948,N_3014,N_3010);
xor U3949 (N_3949,N_3345,N_3448);
or U3950 (N_3950,N_3492,N_3170);
or U3951 (N_3951,N_3340,N_3373);
xnor U3952 (N_3952,N_3089,N_3440);
nor U3953 (N_3953,N_3063,N_3018);
and U3954 (N_3954,N_3125,N_3163);
and U3955 (N_3955,N_3090,N_3231);
nand U3956 (N_3956,N_3289,N_3427);
nor U3957 (N_3957,N_3024,N_3303);
xor U3958 (N_3958,N_3313,N_3037);
and U3959 (N_3959,N_3320,N_3246);
or U3960 (N_3960,N_3163,N_3489);
xnor U3961 (N_3961,N_3055,N_3178);
nand U3962 (N_3962,N_3363,N_3454);
nand U3963 (N_3963,N_3120,N_3405);
or U3964 (N_3964,N_3138,N_3215);
xor U3965 (N_3965,N_3081,N_3031);
and U3966 (N_3966,N_3148,N_3030);
xor U3967 (N_3967,N_3228,N_3310);
nand U3968 (N_3968,N_3184,N_3111);
and U3969 (N_3969,N_3163,N_3371);
and U3970 (N_3970,N_3396,N_3138);
and U3971 (N_3971,N_3339,N_3027);
nand U3972 (N_3972,N_3083,N_3145);
nor U3973 (N_3973,N_3194,N_3375);
xnor U3974 (N_3974,N_3264,N_3285);
nor U3975 (N_3975,N_3188,N_3064);
xor U3976 (N_3976,N_3026,N_3113);
nor U3977 (N_3977,N_3077,N_3436);
nor U3978 (N_3978,N_3456,N_3303);
nand U3979 (N_3979,N_3452,N_3289);
nand U3980 (N_3980,N_3365,N_3351);
nand U3981 (N_3981,N_3363,N_3484);
nor U3982 (N_3982,N_3063,N_3078);
nand U3983 (N_3983,N_3484,N_3023);
xor U3984 (N_3984,N_3227,N_3430);
xor U3985 (N_3985,N_3307,N_3297);
or U3986 (N_3986,N_3399,N_3436);
xor U3987 (N_3987,N_3499,N_3011);
nand U3988 (N_3988,N_3334,N_3277);
and U3989 (N_3989,N_3136,N_3210);
nand U3990 (N_3990,N_3058,N_3296);
or U3991 (N_3991,N_3177,N_3356);
nor U3992 (N_3992,N_3156,N_3220);
nor U3993 (N_3993,N_3281,N_3230);
or U3994 (N_3994,N_3152,N_3262);
xnor U3995 (N_3995,N_3451,N_3255);
xnor U3996 (N_3996,N_3289,N_3311);
nor U3997 (N_3997,N_3383,N_3247);
nand U3998 (N_3998,N_3235,N_3011);
nor U3999 (N_3999,N_3133,N_3044);
nand U4000 (N_4000,N_3973,N_3913);
and U4001 (N_4001,N_3996,N_3804);
and U4002 (N_4002,N_3650,N_3991);
or U4003 (N_4003,N_3549,N_3563);
nor U4004 (N_4004,N_3929,N_3942);
nor U4005 (N_4005,N_3888,N_3718);
nand U4006 (N_4006,N_3957,N_3949);
nor U4007 (N_4007,N_3544,N_3510);
nor U4008 (N_4008,N_3986,N_3708);
nor U4009 (N_4009,N_3610,N_3784);
nand U4010 (N_4010,N_3717,N_3691);
xor U4011 (N_4011,N_3770,N_3514);
nand U4012 (N_4012,N_3780,N_3935);
nor U4013 (N_4013,N_3604,N_3899);
xnor U4014 (N_4014,N_3698,N_3798);
nor U4015 (N_4015,N_3795,N_3632);
nor U4016 (N_4016,N_3915,N_3838);
and U4017 (N_4017,N_3832,N_3922);
nor U4018 (N_4018,N_3959,N_3559);
nor U4019 (N_4019,N_3778,N_3883);
and U4020 (N_4020,N_3535,N_3966);
and U4021 (N_4021,N_3672,N_3603);
or U4022 (N_4022,N_3782,N_3794);
or U4023 (N_4023,N_3799,N_3602);
nor U4024 (N_4024,N_3532,N_3618);
nand U4025 (N_4025,N_3684,N_3533);
or U4026 (N_4026,N_3926,N_3677);
or U4027 (N_4027,N_3508,N_3692);
or U4028 (N_4028,N_3852,N_3696);
or U4029 (N_4029,N_3856,N_3867);
nor U4030 (N_4030,N_3593,N_3721);
and U4031 (N_4031,N_3729,N_3983);
or U4032 (N_4032,N_3699,N_3556);
xor U4033 (N_4033,N_3657,N_3979);
nand U4034 (N_4034,N_3938,N_3607);
and U4035 (N_4035,N_3900,N_3790);
or U4036 (N_4036,N_3858,N_3519);
nand U4037 (N_4037,N_3786,N_3526);
nand U4038 (N_4038,N_3665,N_3803);
xor U4039 (N_4039,N_3625,N_3555);
xor U4040 (N_4040,N_3725,N_3847);
xor U4041 (N_4041,N_3741,N_3836);
xnor U4042 (N_4042,N_3507,N_3752);
xor U4043 (N_4043,N_3667,N_3728);
nand U4044 (N_4044,N_3932,N_3686);
xor U4045 (N_4045,N_3828,N_3568);
nand U4046 (N_4046,N_3807,N_3878);
xor U4047 (N_4047,N_3678,N_3873);
or U4048 (N_4048,N_3558,N_3592);
nand U4049 (N_4049,N_3525,N_3636);
xnor U4050 (N_4050,N_3992,N_3641);
or U4051 (N_4051,N_3749,N_3887);
xor U4052 (N_4052,N_3703,N_3953);
or U4053 (N_4053,N_3564,N_3802);
and U4054 (N_4054,N_3861,N_3619);
nor U4055 (N_4055,N_3688,N_3785);
and U4056 (N_4056,N_3761,N_3951);
nand U4057 (N_4057,N_3727,N_3612);
xnor U4058 (N_4058,N_3990,N_3750);
and U4059 (N_4059,N_3809,N_3746);
and U4060 (N_4060,N_3527,N_3542);
or U4061 (N_4061,N_3704,N_3710);
nor U4062 (N_4062,N_3787,N_3895);
nor U4063 (N_4063,N_3766,N_3528);
nand U4064 (N_4064,N_3854,N_3849);
or U4065 (N_4065,N_3781,N_3543);
nor U4066 (N_4066,N_3891,N_3754);
nand U4067 (N_4067,N_3585,N_3606);
and U4068 (N_4068,N_3805,N_3723);
xor U4069 (N_4069,N_3868,N_3818);
xnor U4070 (N_4070,N_3806,N_3826);
nand U4071 (N_4071,N_3904,N_3962);
and U4072 (N_4072,N_3881,N_3715);
nand U4073 (N_4073,N_3976,N_3548);
nor U4074 (N_4074,N_3631,N_3815);
or U4075 (N_4075,N_3652,N_3655);
nand U4076 (N_4076,N_3522,N_3911);
xnor U4077 (N_4077,N_3893,N_3981);
and U4078 (N_4078,N_3898,N_3722);
nor U4079 (N_4079,N_3679,N_3892);
or U4080 (N_4080,N_3582,N_3876);
or U4081 (N_4081,N_3874,N_3946);
or U4082 (N_4082,N_3997,N_3651);
xor U4083 (N_4083,N_3999,N_3751);
nor U4084 (N_4084,N_3767,N_3660);
nor U4085 (N_4085,N_3747,N_3853);
and U4086 (N_4086,N_3768,N_3756);
xor U4087 (N_4087,N_3822,N_3531);
nand U4088 (N_4088,N_3940,N_3748);
xor U4089 (N_4089,N_3624,N_3952);
and U4090 (N_4090,N_3529,N_3726);
xor U4091 (N_4091,N_3877,N_3580);
nand U4092 (N_4092,N_3575,N_3759);
nand U4093 (N_4093,N_3812,N_3740);
xnor U4094 (N_4094,N_3909,N_3709);
and U4095 (N_4095,N_3864,N_3960);
nand U4096 (N_4096,N_3705,N_3646);
or U4097 (N_4097,N_3536,N_3865);
nor U4098 (N_4098,N_3565,N_3605);
xnor U4099 (N_4099,N_3987,N_3956);
and U4100 (N_4100,N_3616,N_3863);
and U4101 (N_4101,N_3623,N_3884);
nand U4102 (N_4102,N_3843,N_3654);
nand U4103 (N_4103,N_3994,N_3872);
and U4104 (N_4104,N_3681,N_3998);
nand U4105 (N_4105,N_3560,N_3742);
or U4106 (N_4106,N_3842,N_3554);
xor U4107 (N_4107,N_3967,N_3524);
and U4108 (N_4108,N_3907,N_3534);
xor U4109 (N_4109,N_3820,N_3923);
nand U4110 (N_4110,N_3896,N_3955);
and U4111 (N_4111,N_3816,N_3775);
or U4112 (N_4112,N_3644,N_3914);
and U4113 (N_4113,N_3680,N_3903);
nand U4114 (N_4114,N_3889,N_3902);
nor U4115 (N_4115,N_3628,N_3642);
nand U4116 (N_4116,N_3682,N_3813);
nand U4117 (N_4117,N_3882,N_3954);
or U4118 (N_4118,N_3941,N_3588);
nand U4119 (N_4119,N_3640,N_3615);
nand U4120 (N_4120,N_3894,N_3755);
nand U4121 (N_4121,N_3701,N_3885);
xor U4122 (N_4122,N_3591,N_3505);
xor U4123 (N_4123,N_3738,N_3662);
xor U4124 (N_4124,N_3792,N_3827);
or U4125 (N_4125,N_3779,N_3706);
or U4126 (N_4126,N_3598,N_3875);
nand U4127 (N_4127,N_3601,N_3594);
and U4128 (N_4128,N_3783,N_3919);
and U4129 (N_4129,N_3869,N_3659);
nand U4130 (N_4130,N_3918,N_3924);
nor U4131 (N_4131,N_3859,N_3578);
or U4132 (N_4132,N_3694,N_3714);
xnor U4133 (N_4133,N_3944,N_3579);
nand U4134 (N_4134,N_3673,N_3653);
and U4135 (N_4135,N_3521,N_3974);
xnor U4136 (N_4136,N_3661,N_3576);
xor U4137 (N_4137,N_3656,N_3734);
nor U4138 (N_4138,N_3921,N_3958);
nand U4139 (N_4139,N_3733,N_3939);
and U4140 (N_4140,N_3945,N_3511);
nand U4141 (N_4141,N_3985,N_3622);
and U4142 (N_4142,N_3933,N_3897);
and U4143 (N_4143,N_3712,N_3515);
nor U4144 (N_4144,N_3562,N_3608);
nand U4145 (N_4145,N_3927,N_3648);
xor U4146 (N_4146,N_3948,N_3629);
nor U4147 (N_4147,N_3971,N_3936);
xnor U4148 (N_4148,N_3545,N_3504);
xor U4149 (N_4149,N_3988,N_3512);
and U4150 (N_4150,N_3553,N_3664);
nand U4151 (N_4151,N_3689,N_3586);
or U4152 (N_4152,N_3931,N_3745);
xnor U4153 (N_4153,N_3937,N_3724);
nand U4154 (N_4154,N_3764,N_3583);
or U4155 (N_4155,N_3774,N_3848);
and U4156 (N_4156,N_3736,N_3716);
and U4157 (N_4157,N_3757,N_3829);
xnor U4158 (N_4158,N_3551,N_3972);
and U4159 (N_4159,N_3697,N_3530);
or U4160 (N_4160,N_3500,N_3866);
nor U4161 (N_4161,N_3666,N_3516);
nand U4162 (N_4162,N_3573,N_3763);
nand U4163 (N_4163,N_3860,N_3925);
or U4164 (N_4164,N_3762,N_3934);
xnor U4165 (N_4165,N_3683,N_3796);
xnor U4166 (N_4166,N_3817,N_3808);
or U4167 (N_4167,N_3633,N_3513);
xor U4168 (N_4168,N_3916,N_3503);
and U4169 (N_4169,N_3871,N_3744);
nand U4170 (N_4170,N_3658,N_3502);
nor U4171 (N_4171,N_3737,N_3581);
and U4172 (N_4172,N_3571,N_3574);
nand U4173 (N_4173,N_3595,N_3520);
and U4174 (N_4174,N_3577,N_3980);
nor U4175 (N_4175,N_3765,N_3614);
or U4176 (N_4176,N_3584,N_3850);
xor U4177 (N_4177,N_3674,N_3791);
or U4178 (N_4178,N_3643,N_3518);
xnor U4179 (N_4179,N_3824,N_3645);
nor U4180 (N_4180,N_3590,N_3982);
nand U4181 (N_4181,N_3634,N_3541);
and U4182 (N_4182,N_3839,N_3995);
and U4183 (N_4183,N_3840,N_3908);
nor U4184 (N_4184,N_3506,N_3993);
and U4185 (N_4185,N_3621,N_3823);
and U4186 (N_4186,N_3685,N_3901);
and U4187 (N_4187,N_3857,N_3639);
or U4188 (N_4188,N_3731,N_3713);
and U4189 (N_4189,N_3797,N_3509);
nor U4190 (N_4190,N_3695,N_3669);
xnor U4191 (N_4191,N_3810,N_3928);
or U4192 (N_4192,N_3647,N_3819);
xnor U4193 (N_4193,N_3841,N_3676);
and U4194 (N_4194,N_3950,N_3830);
nor U4195 (N_4195,N_3735,N_3572);
nand U4196 (N_4196,N_3912,N_3964);
xor U4197 (N_4197,N_3930,N_3620);
nor U4198 (N_4198,N_3635,N_3567);
nor U4199 (N_4199,N_3837,N_3977);
xor U4200 (N_4200,N_3814,N_3501);
or U4201 (N_4201,N_3550,N_3788);
and U4202 (N_4202,N_3637,N_3920);
nor U4203 (N_4203,N_3879,N_3906);
or U4204 (N_4204,N_3587,N_3569);
xnor U4205 (N_4205,N_3566,N_3719);
xor U4206 (N_4206,N_3552,N_3589);
nand U4207 (N_4207,N_3561,N_3917);
nor U4208 (N_4208,N_3675,N_3880);
nand U4209 (N_4209,N_3570,N_3711);
or U4210 (N_4210,N_3538,N_3975);
or U4211 (N_4211,N_3771,N_3546);
xnor U4212 (N_4212,N_3831,N_3961);
xor U4213 (N_4213,N_3969,N_3947);
nor U4214 (N_4214,N_3630,N_3821);
xor U4215 (N_4215,N_3539,N_3968);
xor U4216 (N_4216,N_3905,N_3776);
nand U4217 (N_4217,N_3720,N_3965);
nand U4218 (N_4218,N_3537,N_3943);
nor U4219 (N_4219,N_3978,N_3600);
xor U4220 (N_4220,N_3626,N_3963);
xor U4221 (N_4221,N_3772,N_3687);
xnor U4222 (N_4222,N_3769,N_3835);
or U4223 (N_4223,N_3851,N_3760);
and U4224 (N_4224,N_3855,N_3970);
nand U4225 (N_4225,N_3693,N_3890);
nand U4226 (N_4226,N_3557,N_3649);
nor U4227 (N_4227,N_3663,N_3886);
or U4228 (N_4228,N_3989,N_3668);
or U4229 (N_4229,N_3743,N_3671);
nand U4230 (N_4230,N_3789,N_3777);
nor U4231 (N_4231,N_3910,N_3547);
and U4232 (N_4232,N_3540,N_3844);
or U4233 (N_4233,N_3825,N_3670);
or U4234 (N_4234,N_3599,N_3758);
nand U4235 (N_4235,N_3739,N_3793);
nand U4236 (N_4236,N_3597,N_3611);
and U4237 (N_4237,N_3984,N_3523);
nand U4238 (N_4238,N_3627,N_3834);
or U4239 (N_4239,N_3801,N_3845);
and U4240 (N_4240,N_3773,N_3862);
xor U4241 (N_4241,N_3811,N_3707);
nor U4242 (N_4242,N_3753,N_3833);
nand U4243 (N_4243,N_3613,N_3517);
nor U4244 (N_4244,N_3609,N_3702);
nor U4245 (N_4245,N_3846,N_3800);
nor U4246 (N_4246,N_3638,N_3690);
nor U4247 (N_4247,N_3730,N_3732);
xnor U4248 (N_4248,N_3870,N_3700);
xor U4249 (N_4249,N_3596,N_3617);
xnor U4250 (N_4250,N_3597,N_3775);
or U4251 (N_4251,N_3779,N_3753);
nor U4252 (N_4252,N_3839,N_3714);
xor U4253 (N_4253,N_3834,N_3846);
xnor U4254 (N_4254,N_3644,N_3632);
or U4255 (N_4255,N_3734,N_3679);
xor U4256 (N_4256,N_3979,N_3894);
or U4257 (N_4257,N_3533,N_3692);
nand U4258 (N_4258,N_3994,N_3810);
xnor U4259 (N_4259,N_3863,N_3935);
xnor U4260 (N_4260,N_3919,N_3561);
and U4261 (N_4261,N_3717,N_3911);
nand U4262 (N_4262,N_3937,N_3846);
nor U4263 (N_4263,N_3500,N_3809);
nor U4264 (N_4264,N_3636,N_3841);
or U4265 (N_4265,N_3828,N_3933);
and U4266 (N_4266,N_3611,N_3951);
nand U4267 (N_4267,N_3622,N_3735);
and U4268 (N_4268,N_3524,N_3826);
or U4269 (N_4269,N_3753,N_3853);
nor U4270 (N_4270,N_3704,N_3513);
or U4271 (N_4271,N_3875,N_3695);
or U4272 (N_4272,N_3768,N_3957);
nand U4273 (N_4273,N_3636,N_3608);
or U4274 (N_4274,N_3772,N_3969);
and U4275 (N_4275,N_3632,N_3528);
xor U4276 (N_4276,N_3816,N_3709);
nand U4277 (N_4277,N_3645,N_3796);
or U4278 (N_4278,N_3922,N_3958);
or U4279 (N_4279,N_3897,N_3579);
xor U4280 (N_4280,N_3509,N_3537);
nor U4281 (N_4281,N_3806,N_3815);
nor U4282 (N_4282,N_3847,N_3951);
xnor U4283 (N_4283,N_3780,N_3906);
nand U4284 (N_4284,N_3670,N_3921);
xnor U4285 (N_4285,N_3693,N_3656);
and U4286 (N_4286,N_3913,N_3779);
xor U4287 (N_4287,N_3941,N_3758);
nand U4288 (N_4288,N_3682,N_3767);
nor U4289 (N_4289,N_3889,N_3855);
and U4290 (N_4290,N_3868,N_3866);
or U4291 (N_4291,N_3685,N_3804);
nor U4292 (N_4292,N_3793,N_3551);
and U4293 (N_4293,N_3762,N_3825);
and U4294 (N_4294,N_3828,N_3814);
nand U4295 (N_4295,N_3794,N_3875);
and U4296 (N_4296,N_3507,N_3854);
nand U4297 (N_4297,N_3615,N_3751);
nor U4298 (N_4298,N_3640,N_3749);
or U4299 (N_4299,N_3721,N_3983);
nand U4300 (N_4300,N_3634,N_3864);
xor U4301 (N_4301,N_3761,N_3880);
or U4302 (N_4302,N_3760,N_3504);
and U4303 (N_4303,N_3978,N_3597);
nand U4304 (N_4304,N_3802,N_3679);
xor U4305 (N_4305,N_3534,N_3915);
and U4306 (N_4306,N_3662,N_3607);
xor U4307 (N_4307,N_3809,N_3946);
xor U4308 (N_4308,N_3632,N_3604);
nand U4309 (N_4309,N_3906,N_3844);
or U4310 (N_4310,N_3988,N_3655);
and U4311 (N_4311,N_3812,N_3766);
nor U4312 (N_4312,N_3668,N_3809);
nor U4313 (N_4313,N_3679,N_3643);
xnor U4314 (N_4314,N_3887,N_3903);
nand U4315 (N_4315,N_3775,N_3871);
and U4316 (N_4316,N_3729,N_3879);
xnor U4317 (N_4317,N_3641,N_3921);
xor U4318 (N_4318,N_3792,N_3955);
or U4319 (N_4319,N_3703,N_3841);
xnor U4320 (N_4320,N_3774,N_3511);
nand U4321 (N_4321,N_3670,N_3715);
or U4322 (N_4322,N_3790,N_3983);
or U4323 (N_4323,N_3753,N_3848);
nor U4324 (N_4324,N_3818,N_3819);
nand U4325 (N_4325,N_3520,N_3642);
or U4326 (N_4326,N_3916,N_3629);
nor U4327 (N_4327,N_3629,N_3739);
and U4328 (N_4328,N_3669,N_3719);
xnor U4329 (N_4329,N_3603,N_3544);
and U4330 (N_4330,N_3697,N_3815);
and U4331 (N_4331,N_3746,N_3917);
or U4332 (N_4332,N_3633,N_3906);
nand U4333 (N_4333,N_3530,N_3836);
or U4334 (N_4334,N_3842,N_3521);
nand U4335 (N_4335,N_3797,N_3697);
xor U4336 (N_4336,N_3585,N_3521);
nor U4337 (N_4337,N_3749,N_3743);
nor U4338 (N_4338,N_3561,N_3915);
and U4339 (N_4339,N_3981,N_3674);
and U4340 (N_4340,N_3579,N_3707);
xnor U4341 (N_4341,N_3883,N_3627);
nand U4342 (N_4342,N_3998,N_3938);
xnor U4343 (N_4343,N_3720,N_3977);
nand U4344 (N_4344,N_3544,N_3966);
nor U4345 (N_4345,N_3822,N_3764);
nor U4346 (N_4346,N_3592,N_3942);
or U4347 (N_4347,N_3973,N_3669);
nor U4348 (N_4348,N_3653,N_3877);
nor U4349 (N_4349,N_3818,N_3984);
nor U4350 (N_4350,N_3622,N_3872);
xor U4351 (N_4351,N_3940,N_3785);
nand U4352 (N_4352,N_3742,N_3656);
xnor U4353 (N_4353,N_3990,N_3916);
nor U4354 (N_4354,N_3861,N_3533);
nand U4355 (N_4355,N_3814,N_3992);
xnor U4356 (N_4356,N_3795,N_3833);
or U4357 (N_4357,N_3754,N_3739);
and U4358 (N_4358,N_3836,N_3897);
nor U4359 (N_4359,N_3814,N_3700);
or U4360 (N_4360,N_3516,N_3871);
and U4361 (N_4361,N_3796,N_3627);
nand U4362 (N_4362,N_3844,N_3617);
and U4363 (N_4363,N_3615,N_3955);
nor U4364 (N_4364,N_3587,N_3849);
xnor U4365 (N_4365,N_3952,N_3555);
and U4366 (N_4366,N_3985,N_3675);
nor U4367 (N_4367,N_3736,N_3562);
nand U4368 (N_4368,N_3566,N_3675);
and U4369 (N_4369,N_3761,N_3503);
xor U4370 (N_4370,N_3538,N_3995);
nor U4371 (N_4371,N_3922,N_3622);
and U4372 (N_4372,N_3691,N_3863);
nor U4373 (N_4373,N_3774,N_3510);
nand U4374 (N_4374,N_3528,N_3676);
nand U4375 (N_4375,N_3910,N_3791);
nor U4376 (N_4376,N_3989,N_3903);
or U4377 (N_4377,N_3778,N_3953);
or U4378 (N_4378,N_3540,N_3845);
and U4379 (N_4379,N_3506,N_3835);
nor U4380 (N_4380,N_3724,N_3675);
and U4381 (N_4381,N_3805,N_3819);
and U4382 (N_4382,N_3739,N_3959);
xnor U4383 (N_4383,N_3973,N_3774);
xnor U4384 (N_4384,N_3602,N_3650);
nand U4385 (N_4385,N_3698,N_3764);
nand U4386 (N_4386,N_3673,N_3548);
or U4387 (N_4387,N_3710,N_3636);
or U4388 (N_4388,N_3686,N_3927);
or U4389 (N_4389,N_3674,N_3564);
xnor U4390 (N_4390,N_3571,N_3679);
nor U4391 (N_4391,N_3981,N_3524);
and U4392 (N_4392,N_3588,N_3780);
or U4393 (N_4393,N_3869,N_3523);
nor U4394 (N_4394,N_3963,N_3518);
or U4395 (N_4395,N_3692,N_3558);
xor U4396 (N_4396,N_3874,N_3763);
nor U4397 (N_4397,N_3656,N_3858);
xnor U4398 (N_4398,N_3872,N_3884);
or U4399 (N_4399,N_3700,N_3640);
and U4400 (N_4400,N_3870,N_3853);
and U4401 (N_4401,N_3798,N_3782);
nor U4402 (N_4402,N_3907,N_3512);
xor U4403 (N_4403,N_3597,N_3668);
or U4404 (N_4404,N_3500,N_3727);
nand U4405 (N_4405,N_3689,N_3775);
or U4406 (N_4406,N_3501,N_3884);
nor U4407 (N_4407,N_3847,N_3591);
xor U4408 (N_4408,N_3833,N_3813);
and U4409 (N_4409,N_3834,N_3787);
and U4410 (N_4410,N_3960,N_3756);
or U4411 (N_4411,N_3953,N_3609);
and U4412 (N_4412,N_3917,N_3609);
or U4413 (N_4413,N_3863,N_3824);
and U4414 (N_4414,N_3584,N_3597);
nand U4415 (N_4415,N_3571,N_3729);
or U4416 (N_4416,N_3799,N_3883);
nor U4417 (N_4417,N_3660,N_3863);
or U4418 (N_4418,N_3592,N_3573);
xnor U4419 (N_4419,N_3822,N_3891);
and U4420 (N_4420,N_3671,N_3505);
nor U4421 (N_4421,N_3638,N_3547);
nand U4422 (N_4422,N_3982,N_3605);
xor U4423 (N_4423,N_3940,N_3623);
nand U4424 (N_4424,N_3627,N_3672);
and U4425 (N_4425,N_3876,N_3780);
xnor U4426 (N_4426,N_3558,N_3910);
nor U4427 (N_4427,N_3785,N_3948);
and U4428 (N_4428,N_3755,N_3816);
nor U4429 (N_4429,N_3563,N_3804);
nor U4430 (N_4430,N_3977,N_3518);
xnor U4431 (N_4431,N_3592,N_3693);
or U4432 (N_4432,N_3505,N_3810);
or U4433 (N_4433,N_3861,N_3655);
or U4434 (N_4434,N_3929,N_3524);
xor U4435 (N_4435,N_3636,N_3781);
xnor U4436 (N_4436,N_3721,N_3548);
nand U4437 (N_4437,N_3865,N_3873);
or U4438 (N_4438,N_3682,N_3774);
or U4439 (N_4439,N_3660,N_3799);
or U4440 (N_4440,N_3613,N_3750);
xnor U4441 (N_4441,N_3753,N_3545);
nand U4442 (N_4442,N_3979,N_3692);
nand U4443 (N_4443,N_3772,N_3848);
and U4444 (N_4444,N_3942,N_3519);
xor U4445 (N_4445,N_3581,N_3709);
nand U4446 (N_4446,N_3656,N_3839);
xnor U4447 (N_4447,N_3552,N_3977);
or U4448 (N_4448,N_3940,N_3853);
or U4449 (N_4449,N_3854,N_3967);
nor U4450 (N_4450,N_3715,N_3814);
or U4451 (N_4451,N_3976,N_3862);
nor U4452 (N_4452,N_3553,N_3518);
and U4453 (N_4453,N_3844,N_3960);
xnor U4454 (N_4454,N_3553,N_3776);
and U4455 (N_4455,N_3544,N_3652);
xnor U4456 (N_4456,N_3937,N_3609);
nand U4457 (N_4457,N_3739,N_3682);
nand U4458 (N_4458,N_3635,N_3628);
nand U4459 (N_4459,N_3561,N_3690);
nor U4460 (N_4460,N_3841,N_3873);
xor U4461 (N_4461,N_3992,N_3986);
or U4462 (N_4462,N_3999,N_3588);
or U4463 (N_4463,N_3624,N_3884);
and U4464 (N_4464,N_3928,N_3688);
xor U4465 (N_4465,N_3942,N_3833);
or U4466 (N_4466,N_3884,N_3999);
xor U4467 (N_4467,N_3707,N_3552);
xnor U4468 (N_4468,N_3863,N_3868);
nor U4469 (N_4469,N_3577,N_3907);
or U4470 (N_4470,N_3565,N_3923);
nor U4471 (N_4471,N_3600,N_3982);
nand U4472 (N_4472,N_3844,N_3934);
and U4473 (N_4473,N_3528,N_3648);
nor U4474 (N_4474,N_3617,N_3882);
nor U4475 (N_4475,N_3867,N_3704);
and U4476 (N_4476,N_3513,N_3951);
nand U4477 (N_4477,N_3539,N_3824);
or U4478 (N_4478,N_3616,N_3858);
xnor U4479 (N_4479,N_3543,N_3689);
nor U4480 (N_4480,N_3904,N_3716);
nand U4481 (N_4481,N_3671,N_3543);
nor U4482 (N_4482,N_3749,N_3606);
or U4483 (N_4483,N_3607,N_3703);
nor U4484 (N_4484,N_3637,N_3768);
nand U4485 (N_4485,N_3952,N_3804);
nand U4486 (N_4486,N_3611,N_3998);
or U4487 (N_4487,N_3566,N_3838);
xnor U4488 (N_4488,N_3828,N_3629);
or U4489 (N_4489,N_3826,N_3841);
xnor U4490 (N_4490,N_3717,N_3851);
and U4491 (N_4491,N_3973,N_3595);
or U4492 (N_4492,N_3998,N_3901);
nor U4493 (N_4493,N_3687,N_3531);
xnor U4494 (N_4494,N_3962,N_3871);
or U4495 (N_4495,N_3614,N_3701);
or U4496 (N_4496,N_3992,N_3600);
xor U4497 (N_4497,N_3703,N_3632);
nor U4498 (N_4498,N_3619,N_3568);
or U4499 (N_4499,N_3935,N_3926);
xnor U4500 (N_4500,N_4110,N_4396);
xor U4501 (N_4501,N_4099,N_4214);
nand U4502 (N_4502,N_4415,N_4182);
nor U4503 (N_4503,N_4123,N_4255);
or U4504 (N_4504,N_4398,N_4282);
nor U4505 (N_4505,N_4472,N_4073);
and U4506 (N_4506,N_4471,N_4039);
nor U4507 (N_4507,N_4476,N_4117);
or U4508 (N_4508,N_4306,N_4355);
xnor U4509 (N_4509,N_4218,N_4288);
nand U4510 (N_4510,N_4145,N_4058);
and U4511 (N_4511,N_4079,N_4393);
or U4512 (N_4512,N_4247,N_4050);
and U4513 (N_4513,N_4049,N_4443);
nor U4514 (N_4514,N_4234,N_4114);
or U4515 (N_4515,N_4430,N_4297);
xnor U4516 (N_4516,N_4485,N_4186);
or U4517 (N_4517,N_4104,N_4468);
nand U4518 (N_4518,N_4394,N_4409);
xor U4519 (N_4519,N_4286,N_4047);
xor U4520 (N_4520,N_4364,N_4169);
nor U4521 (N_4521,N_4360,N_4298);
nor U4522 (N_4522,N_4413,N_4420);
nand U4523 (N_4523,N_4438,N_4236);
or U4524 (N_4524,N_4264,N_4275);
nor U4525 (N_4525,N_4347,N_4412);
nand U4526 (N_4526,N_4313,N_4192);
xor U4527 (N_4527,N_4008,N_4051);
nand U4528 (N_4528,N_4144,N_4404);
xnor U4529 (N_4529,N_4097,N_4400);
nand U4530 (N_4530,N_4034,N_4055);
or U4531 (N_4531,N_4054,N_4273);
nor U4532 (N_4532,N_4450,N_4482);
nor U4533 (N_4533,N_4249,N_4378);
and U4534 (N_4534,N_4451,N_4124);
nand U4535 (N_4535,N_4066,N_4277);
nor U4536 (N_4536,N_4194,N_4291);
xor U4537 (N_4537,N_4109,N_4102);
nor U4538 (N_4538,N_4159,N_4258);
nand U4539 (N_4539,N_4287,N_4311);
or U4540 (N_4540,N_4452,N_4025);
and U4541 (N_4541,N_4022,N_4209);
nor U4542 (N_4542,N_4361,N_4017);
or U4543 (N_4543,N_4294,N_4065);
nand U4544 (N_4544,N_4279,N_4268);
or U4545 (N_4545,N_4310,N_4441);
or U4546 (N_4546,N_4187,N_4377);
nand U4547 (N_4547,N_4375,N_4293);
nand U4548 (N_4548,N_4416,N_4316);
and U4549 (N_4549,N_4067,N_4333);
nand U4550 (N_4550,N_4308,N_4334);
nand U4551 (N_4551,N_4053,N_4350);
nor U4552 (N_4552,N_4447,N_4344);
or U4553 (N_4553,N_4033,N_4204);
and U4554 (N_4554,N_4084,N_4388);
nand U4555 (N_4555,N_4399,N_4405);
nor U4556 (N_4556,N_4354,N_4425);
or U4557 (N_4557,N_4418,N_4189);
and U4558 (N_4558,N_4238,N_4351);
or U4559 (N_4559,N_4335,N_4184);
xor U4560 (N_4560,N_4095,N_4357);
nor U4561 (N_4561,N_4496,N_4081);
nor U4562 (N_4562,N_4410,N_4202);
nand U4563 (N_4563,N_4101,N_4001);
or U4564 (N_4564,N_4337,N_4385);
and U4565 (N_4565,N_4487,N_4307);
nand U4566 (N_4566,N_4417,N_4370);
nand U4567 (N_4567,N_4453,N_4040);
or U4568 (N_4568,N_4078,N_4281);
nand U4569 (N_4569,N_4088,N_4480);
nor U4570 (N_4570,N_4036,N_4115);
or U4571 (N_4571,N_4455,N_4086);
xnor U4572 (N_4572,N_4367,N_4029);
xnor U4573 (N_4573,N_4188,N_4440);
and U4574 (N_4574,N_4203,N_4449);
or U4575 (N_4575,N_4241,N_4434);
nor U4576 (N_4576,N_4406,N_4057);
nand U4577 (N_4577,N_4469,N_4111);
nand U4578 (N_4578,N_4063,N_4250);
or U4579 (N_4579,N_4136,N_4295);
and U4580 (N_4580,N_4387,N_4183);
and U4581 (N_4581,N_4106,N_4301);
xor U4582 (N_4582,N_4037,N_4220);
xnor U4583 (N_4583,N_4042,N_4374);
or U4584 (N_4584,N_4402,N_4401);
or U4585 (N_4585,N_4479,N_4386);
and U4586 (N_4586,N_4325,N_4197);
xnor U4587 (N_4587,N_4225,N_4201);
xnor U4588 (N_4588,N_4475,N_4363);
and U4589 (N_4589,N_4177,N_4075);
nor U4590 (N_4590,N_4271,N_4213);
or U4591 (N_4591,N_4092,N_4024);
and U4592 (N_4592,N_4390,N_4373);
nand U4593 (N_4593,N_4215,N_4445);
xnor U4594 (N_4594,N_4164,N_4314);
or U4595 (N_4595,N_4312,N_4219);
or U4596 (N_4596,N_4148,N_4135);
and U4597 (N_4597,N_4019,N_4478);
or U4598 (N_4598,N_4224,N_4243);
nor U4599 (N_4599,N_4369,N_4368);
and U4600 (N_4600,N_4221,N_4062);
nor U4601 (N_4601,N_4226,N_4199);
or U4602 (N_4602,N_4459,N_4230);
or U4603 (N_4603,N_4392,N_4423);
xnor U4604 (N_4604,N_4432,N_4484);
nand U4605 (N_4605,N_4082,N_4163);
nor U4606 (N_4606,N_4191,N_4069);
nor U4607 (N_4607,N_4331,N_4171);
nand U4608 (N_4608,N_4437,N_4251);
nor U4609 (N_4609,N_4030,N_4353);
nor U4610 (N_4610,N_4495,N_4462);
and U4611 (N_4611,N_4113,N_4041);
xnor U4612 (N_4612,N_4210,N_4276);
xor U4613 (N_4613,N_4460,N_4151);
nand U4614 (N_4614,N_4003,N_4132);
and U4615 (N_4615,N_4465,N_4242);
nand U4616 (N_4616,N_4427,N_4232);
and U4617 (N_4617,N_4077,N_4231);
xnor U4618 (N_4618,N_4456,N_4160);
nor U4619 (N_4619,N_4379,N_4179);
nand U4620 (N_4620,N_4365,N_4384);
and U4621 (N_4621,N_4020,N_4309);
or U4622 (N_4622,N_4269,N_4157);
or U4623 (N_4623,N_4146,N_4481);
or U4624 (N_4624,N_4349,N_4428);
nor U4625 (N_4625,N_4080,N_4004);
nand U4626 (N_4626,N_4228,N_4499);
nor U4627 (N_4627,N_4137,N_4270);
xor U4628 (N_4628,N_4116,N_4190);
nand U4629 (N_4629,N_4457,N_4252);
and U4630 (N_4630,N_4407,N_4257);
xnor U4631 (N_4631,N_4071,N_4149);
nor U4632 (N_4632,N_4380,N_4015);
nor U4633 (N_4633,N_4152,N_4166);
and U4634 (N_4634,N_4035,N_4346);
nand U4635 (N_4635,N_4296,N_4429);
and U4636 (N_4636,N_4319,N_4324);
nor U4637 (N_4637,N_4139,N_4473);
nand U4638 (N_4638,N_4285,N_4359);
or U4639 (N_4639,N_4222,N_4383);
and U4640 (N_4640,N_4498,N_4074);
or U4641 (N_4641,N_4076,N_4208);
xor U4642 (N_4642,N_4422,N_4127);
and U4643 (N_4643,N_4094,N_4060);
nor U4644 (N_4644,N_4336,N_4464);
nand U4645 (N_4645,N_4403,N_4138);
or U4646 (N_4646,N_4267,N_4463);
nand U4647 (N_4647,N_4283,N_4332);
xnor U4648 (N_4648,N_4320,N_4175);
nand U4649 (N_4649,N_4007,N_4227);
nor U4650 (N_4650,N_4072,N_4431);
and U4651 (N_4651,N_4474,N_4489);
xnor U4652 (N_4652,N_4343,N_4289);
or U4653 (N_4653,N_4193,N_4292);
or U4654 (N_4654,N_4180,N_4435);
nand U4655 (N_4655,N_4005,N_4326);
and U4656 (N_4656,N_4170,N_4128);
xnor U4657 (N_4657,N_4059,N_4248);
or U4658 (N_4658,N_4090,N_4112);
nor U4659 (N_4659,N_4263,N_4056);
and U4660 (N_4660,N_4064,N_4176);
nand U4661 (N_4661,N_4358,N_4200);
nand U4662 (N_4662,N_4131,N_4046);
and U4663 (N_4663,N_4439,N_4356);
or U4664 (N_4664,N_4143,N_4173);
nand U4665 (N_4665,N_4240,N_4305);
nand U4666 (N_4666,N_4391,N_4016);
or U4667 (N_4667,N_4198,N_4129);
nand U4668 (N_4668,N_4419,N_4010);
and U4669 (N_4669,N_4239,N_4206);
or U4670 (N_4670,N_4245,N_4329);
nand U4671 (N_4671,N_4362,N_4491);
and U4672 (N_4672,N_4207,N_4235);
nor U4673 (N_4673,N_4253,N_4426);
xnor U4674 (N_4674,N_4376,N_4290);
xor U4675 (N_4675,N_4038,N_4013);
nand U4676 (N_4676,N_4299,N_4096);
or U4677 (N_4677,N_4266,N_4223);
and U4678 (N_4678,N_4317,N_4321);
nor U4679 (N_4679,N_4216,N_4408);
nor U4680 (N_4680,N_4284,N_4421);
nand U4681 (N_4681,N_4083,N_4167);
nor U4682 (N_4682,N_4246,N_4488);
nor U4683 (N_4683,N_4028,N_4107);
and U4684 (N_4684,N_4023,N_4260);
xor U4685 (N_4685,N_4211,N_4304);
or U4686 (N_4686,N_4126,N_4256);
and U4687 (N_4687,N_4133,N_4070);
and U4688 (N_4688,N_4342,N_4161);
xnor U4689 (N_4689,N_4461,N_4483);
nand U4690 (N_4690,N_4091,N_4068);
nor U4691 (N_4691,N_4093,N_4382);
nand U4692 (N_4692,N_4486,N_4061);
and U4693 (N_4693,N_4466,N_4205);
or U4694 (N_4694,N_4442,N_4140);
or U4695 (N_4695,N_4155,N_4278);
or U4696 (N_4696,N_4244,N_4233);
xnor U4697 (N_4697,N_4045,N_4009);
or U4698 (N_4698,N_4444,N_4318);
nand U4699 (N_4699,N_4103,N_4181);
nand U4700 (N_4700,N_4323,N_4454);
and U4701 (N_4701,N_4156,N_4446);
nand U4702 (N_4702,N_4389,N_4031);
nor U4703 (N_4703,N_4172,N_4217);
or U4704 (N_4704,N_4492,N_4340);
and U4705 (N_4705,N_4153,N_4302);
nand U4706 (N_4706,N_4327,N_4012);
nor U4707 (N_4707,N_4021,N_4371);
and U4708 (N_4708,N_4490,N_4470);
nand U4709 (N_4709,N_4006,N_4158);
nor U4710 (N_4710,N_4119,N_4026);
nor U4711 (N_4711,N_4014,N_4147);
xnor U4712 (N_4712,N_4120,N_4048);
nor U4713 (N_4713,N_4458,N_4162);
nand U4714 (N_4714,N_4280,N_4044);
xor U4715 (N_4715,N_4467,N_4168);
xnor U4716 (N_4716,N_4000,N_4237);
nor U4717 (N_4717,N_4027,N_4142);
and U4718 (N_4718,N_4043,N_4352);
nand U4719 (N_4719,N_4125,N_4322);
nor U4720 (N_4720,N_4141,N_4032);
or U4721 (N_4721,N_4178,N_4348);
and U4722 (N_4722,N_4098,N_4262);
nand U4723 (N_4723,N_4018,N_4341);
xor U4724 (N_4724,N_4011,N_4345);
or U4725 (N_4725,N_4254,N_4195);
nand U4726 (N_4726,N_4196,N_4300);
nor U4727 (N_4727,N_4424,N_4411);
nor U4728 (N_4728,N_4315,N_4395);
or U4729 (N_4729,N_4397,N_4002);
nor U4730 (N_4730,N_4150,N_4089);
nand U4731 (N_4731,N_4414,N_4052);
xnor U4732 (N_4732,N_4108,N_4185);
nand U4733 (N_4733,N_4436,N_4212);
nand U4734 (N_4734,N_4174,N_4303);
or U4735 (N_4735,N_4497,N_4118);
nor U4736 (N_4736,N_4477,N_4122);
nor U4737 (N_4737,N_4366,N_4339);
or U4738 (N_4738,N_4372,N_4494);
nand U4739 (N_4739,N_4165,N_4261);
nor U4740 (N_4740,N_4265,N_4328);
and U4741 (N_4741,N_4100,N_4433);
xor U4742 (N_4742,N_4154,N_4229);
or U4743 (N_4743,N_4381,N_4274);
nand U4744 (N_4744,N_4134,N_4259);
xor U4745 (N_4745,N_4272,N_4130);
or U4746 (N_4746,N_4121,N_4338);
and U4747 (N_4747,N_4330,N_4493);
nand U4748 (N_4748,N_4448,N_4105);
or U4749 (N_4749,N_4085,N_4087);
xnor U4750 (N_4750,N_4242,N_4289);
xnor U4751 (N_4751,N_4202,N_4167);
nand U4752 (N_4752,N_4257,N_4037);
and U4753 (N_4753,N_4489,N_4339);
nand U4754 (N_4754,N_4092,N_4408);
nand U4755 (N_4755,N_4333,N_4215);
nor U4756 (N_4756,N_4167,N_4229);
or U4757 (N_4757,N_4413,N_4263);
and U4758 (N_4758,N_4479,N_4390);
xnor U4759 (N_4759,N_4430,N_4346);
xnor U4760 (N_4760,N_4383,N_4273);
nor U4761 (N_4761,N_4437,N_4300);
nand U4762 (N_4762,N_4370,N_4386);
and U4763 (N_4763,N_4059,N_4153);
and U4764 (N_4764,N_4190,N_4201);
and U4765 (N_4765,N_4186,N_4160);
nand U4766 (N_4766,N_4415,N_4372);
and U4767 (N_4767,N_4189,N_4118);
nand U4768 (N_4768,N_4406,N_4476);
nor U4769 (N_4769,N_4422,N_4431);
or U4770 (N_4770,N_4098,N_4166);
nor U4771 (N_4771,N_4279,N_4490);
nand U4772 (N_4772,N_4427,N_4033);
or U4773 (N_4773,N_4141,N_4187);
nor U4774 (N_4774,N_4405,N_4182);
xnor U4775 (N_4775,N_4119,N_4313);
xnor U4776 (N_4776,N_4466,N_4467);
or U4777 (N_4777,N_4293,N_4018);
and U4778 (N_4778,N_4113,N_4279);
and U4779 (N_4779,N_4385,N_4236);
or U4780 (N_4780,N_4343,N_4328);
xor U4781 (N_4781,N_4145,N_4082);
and U4782 (N_4782,N_4283,N_4109);
nor U4783 (N_4783,N_4185,N_4230);
and U4784 (N_4784,N_4479,N_4017);
xnor U4785 (N_4785,N_4022,N_4027);
nand U4786 (N_4786,N_4001,N_4332);
or U4787 (N_4787,N_4492,N_4174);
xnor U4788 (N_4788,N_4281,N_4054);
nor U4789 (N_4789,N_4194,N_4496);
and U4790 (N_4790,N_4255,N_4160);
nor U4791 (N_4791,N_4374,N_4161);
xnor U4792 (N_4792,N_4028,N_4459);
or U4793 (N_4793,N_4206,N_4244);
nand U4794 (N_4794,N_4039,N_4286);
or U4795 (N_4795,N_4152,N_4129);
or U4796 (N_4796,N_4145,N_4287);
and U4797 (N_4797,N_4469,N_4346);
nand U4798 (N_4798,N_4441,N_4453);
and U4799 (N_4799,N_4257,N_4042);
or U4800 (N_4800,N_4059,N_4470);
nand U4801 (N_4801,N_4286,N_4117);
or U4802 (N_4802,N_4201,N_4207);
nor U4803 (N_4803,N_4003,N_4078);
or U4804 (N_4804,N_4132,N_4395);
or U4805 (N_4805,N_4318,N_4237);
xnor U4806 (N_4806,N_4161,N_4019);
nand U4807 (N_4807,N_4370,N_4059);
xnor U4808 (N_4808,N_4307,N_4019);
nand U4809 (N_4809,N_4194,N_4126);
nand U4810 (N_4810,N_4484,N_4141);
nand U4811 (N_4811,N_4335,N_4091);
and U4812 (N_4812,N_4079,N_4319);
nor U4813 (N_4813,N_4008,N_4081);
nand U4814 (N_4814,N_4101,N_4239);
nand U4815 (N_4815,N_4342,N_4469);
nand U4816 (N_4816,N_4290,N_4272);
xor U4817 (N_4817,N_4423,N_4069);
and U4818 (N_4818,N_4227,N_4068);
or U4819 (N_4819,N_4271,N_4499);
xor U4820 (N_4820,N_4187,N_4331);
nor U4821 (N_4821,N_4308,N_4454);
nand U4822 (N_4822,N_4422,N_4201);
nand U4823 (N_4823,N_4426,N_4403);
nor U4824 (N_4824,N_4234,N_4218);
and U4825 (N_4825,N_4499,N_4004);
or U4826 (N_4826,N_4131,N_4496);
nand U4827 (N_4827,N_4245,N_4175);
nand U4828 (N_4828,N_4455,N_4254);
and U4829 (N_4829,N_4306,N_4061);
xor U4830 (N_4830,N_4237,N_4320);
nor U4831 (N_4831,N_4114,N_4482);
and U4832 (N_4832,N_4286,N_4176);
xor U4833 (N_4833,N_4426,N_4069);
and U4834 (N_4834,N_4192,N_4262);
nand U4835 (N_4835,N_4311,N_4018);
or U4836 (N_4836,N_4288,N_4148);
and U4837 (N_4837,N_4243,N_4015);
xor U4838 (N_4838,N_4400,N_4374);
nor U4839 (N_4839,N_4163,N_4125);
nor U4840 (N_4840,N_4468,N_4350);
and U4841 (N_4841,N_4340,N_4205);
nand U4842 (N_4842,N_4104,N_4001);
nand U4843 (N_4843,N_4401,N_4456);
nand U4844 (N_4844,N_4005,N_4087);
xor U4845 (N_4845,N_4341,N_4330);
or U4846 (N_4846,N_4453,N_4297);
and U4847 (N_4847,N_4372,N_4113);
or U4848 (N_4848,N_4301,N_4194);
xnor U4849 (N_4849,N_4091,N_4128);
xor U4850 (N_4850,N_4225,N_4203);
and U4851 (N_4851,N_4049,N_4213);
and U4852 (N_4852,N_4341,N_4270);
or U4853 (N_4853,N_4363,N_4261);
xnor U4854 (N_4854,N_4397,N_4340);
nand U4855 (N_4855,N_4164,N_4056);
nor U4856 (N_4856,N_4318,N_4145);
xor U4857 (N_4857,N_4389,N_4441);
nand U4858 (N_4858,N_4093,N_4461);
nand U4859 (N_4859,N_4047,N_4080);
xor U4860 (N_4860,N_4016,N_4338);
nor U4861 (N_4861,N_4125,N_4052);
nand U4862 (N_4862,N_4334,N_4330);
nand U4863 (N_4863,N_4313,N_4238);
or U4864 (N_4864,N_4495,N_4006);
nor U4865 (N_4865,N_4319,N_4254);
xor U4866 (N_4866,N_4079,N_4363);
xor U4867 (N_4867,N_4152,N_4067);
and U4868 (N_4868,N_4450,N_4441);
or U4869 (N_4869,N_4446,N_4323);
or U4870 (N_4870,N_4129,N_4205);
xor U4871 (N_4871,N_4292,N_4134);
xnor U4872 (N_4872,N_4354,N_4028);
and U4873 (N_4873,N_4244,N_4016);
nor U4874 (N_4874,N_4358,N_4296);
and U4875 (N_4875,N_4062,N_4311);
nand U4876 (N_4876,N_4055,N_4467);
xnor U4877 (N_4877,N_4331,N_4053);
or U4878 (N_4878,N_4107,N_4318);
nor U4879 (N_4879,N_4095,N_4155);
nor U4880 (N_4880,N_4323,N_4259);
xor U4881 (N_4881,N_4399,N_4129);
nand U4882 (N_4882,N_4437,N_4139);
xnor U4883 (N_4883,N_4453,N_4088);
or U4884 (N_4884,N_4394,N_4200);
nor U4885 (N_4885,N_4499,N_4395);
xnor U4886 (N_4886,N_4443,N_4051);
and U4887 (N_4887,N_4350,N_4115);
nor U4888 (N_4888,N_4398,N_4464);
and U4889 (N_4889,N_4041,N_4173);
xnor U4890 (N_4890,N_4163,N_4398);
nand U4891 (N_4891,N_4084,N_4493);
or U4892 (N_4892,N_4378,N_4325);
or U4893 (N_4893,N_4444,N_4421);
or U4894 (N_4894,N_4077,N_4009);
and U4895 (N_4895,N_4235,N_4480);
nor U4896 (N_4896,N_4366,N_4217);
or U4897 (N_4897,N_4150,N_4475);
nand U4898 (N_4898,N_4294,N_4072);
nor U4899 (N_4899,N_4005,N_4295);
nand U4900 (N_4900,N_4187,N_4378);
xnor U4901 (N_4901,N_4335,N_4486);
and U4902 (N_4902,N_4394,N_4389);
and U4903 (N_4903,N_4455,N_4167);
and U4904 (N_4904,N_4050,N_4323);
and U4905 (N_4905,N_4350,N_4110);
and U4906 (N_4906,N_4281,N_4349);
and U4907 (N_4907,N_4200,N_4447);
and U4908 (N_4908,N_4113,N_4194);
nand U4909 (N_4909,N_4136,N_4486);
nand U4910 (N_4910,N_4040,N_4134);
and U4911 (N_4911,N_4149,N_4439);
nor U4912 (N_4912,N_4264,N_4303);
xnor U4913 (N_4913,N_4358,N_4210);
nor U4914 (N_4914,N_4091,N_4080);
xnor U4915 (N_4915,N_4482,N_4340);
nand U4916 (N_4916,N_4138,N_4125);
xor U4917 (N_4917,N_4153,N_4475);
nor U4918 (N_4918,N_4475,N_4303);
nor U4919 (N_4919,N_4355,N_4101);
xor U4920 (N_4920,N_4301,N_4244);
xor U4921 (N_4921,N_4236,N_4489);
xor U4922 (N_4922,N_4054,N_4268);
xor U4923 (N_4923,N_4344,N_4437);
nand U4924 (N_4924,N_4041,N_4279);
and U4925 (N_4925,N_4365,N_4150);
nor U4926 (N_4926,N_4308,N_4012);
nand U4927 (N_4927,N_4191,N_4000);
nor U4928 (N_4928,N_4125,N_4297);
and U4929 (N_4929,N_4379,N_4390);
nor U4930 (N_4930,N_4396,N_4268);
nor U4931 (N_4931,N_4318,N_4441);
and U4932 (N_4932,N_4131,N_4339);
nand U4933 (N_4933,N_4220,N_4046);
or U4934 (N_4934,N_4217,N_4136);
nor U4935 (N_4935,N_4181,N_4460);
nor U4936 (N_4936,N_4447,N_4434);
nand U4937 (N_4937,N_4435,N_4244);
and U4938 (N_4938,N_4142,N_4446);
or U4939 (N_4939,N_4311,N_4110);
or U4940 (N_4940,N_4297,N_4370);
and U4941 (N_4941,N_4301,N_4087);
nand U4942 (N_4942,N_4379,N_4461);
nor U4943 (N_4943,N_4213,N_4348);
xnor U4944 (N_4944,N_4423,N_4168);
nand U4945 (N_4945,N_4291,N_4131);
xnor U4946 (N_4946,N_4454,N_4301);
nor U4947 (N_4947,N_4179,N_4234);
or U4948 (N_4948,N_4359,N_4338);
and U4949 (N_4949,N_4391,N_4224);
nand U4950 (N_4950,N_4388,N_4096);
and U4951 (N_4951,N_4325,N_4320);
nor U4952 (N_4952,N_4333,N_4048);
nor U4953 (N_4953,N_4361,N_4357);
nand U4954 (N_4954,N_4197,N_4144);
xor U4955 (N_4955,N_4464,N_4341);
xor U4956 (N_4956,N_4416,N_4064);
and U4957 (N_4957,N_4199,N_4227);
nor U4958 (N_4958,N_4204,N_4175);
nand U4959 (N_4959,N_4022,N_4460);
nor U4960 (N_4960,N_4409,N_4309);
nand U4961 (N_4961,N_4302,N_4174);
nor U4962 (N_4962,N_4129,N_4468);
nand U4963 (N_4963,N_4320,N_4221);
nand U4964 (N_4964,N_4260,N_4488);
and U4965 (N_4965,N_4008,N_4392);
nor U4966 (N_4966,N_4133,N_4190);
xnor U4967 (N_4967,N_4293,N_4334);
nor U4968 (N_4968,N_4105,N_4142);
nand U4969 (N_4969,N_4461,N_4068);
xnor U4970 (N_4970,N_4008,N_4328);
nand U4971 (N_4971,N_4233,N_4093);
nor U4972 (N_4972,N_4100,N_4215);
or U4973 (N_4973,N_4114,N_4238);
and U4974 (N_4974,N_4023,N_4146);
nor U4975 (N_4975,N_4225,N_4434);
nand U4976 (N_4976,N_4093,N_4011);
and U4977 (N_4977,N_4053,N_4220);
nor U4978 (N_4978,N_4471,N_4180);
or U4979 (N_4979,N_4351,N_4473);
nand U4980 (N_4980,N_4447,N_4247);
xor U4981 (N_4981,N_4243,N_4013);
nand U4982 (N_4982,N_4283,N_4417);
or U4983 (N_4983,N_4486,N_4443);
nand U4984 (N_4984,N_4443,N_4139);
nand U4985 (N_4985,N_4428,N_4490);
nor U4986 (N_4986,N_4483,N_4331);
nand U4987 (N_4987,N_4234,N_4070);
or U4988 (N_4988,N_4179,N_4062);
or U4989 (N_4989,N_4131,N_4292);
nand U4990 (N_4990,N_4449,N_4061);
nor U4991 (N_4991,N_4412,N_4156);
and U4992 (N_4992,N_4317,N_4000);
or U4993 (N_4993,N_4328,N_4150);
or U4994 (N_4994,N_4074,N_4426);
nor U4995 (N_4995,N_4318,N_4369);
and U4996 (N_4996,N_4082,N_4310);
nor U4997 (N_4997,N_4393,N_4217);
or U4998 (N_4998,N_4209,N_4138);
xnor U4999 (N_4999,N_4346,N_4476);
and U5000 (N_5000,N_4707,N_4511);
xnor U5001 (N_5001,N_4634,N_4543);
or U5002 (N_5002,N_4930,N_4858);
or U5003 (N_5003,N_4598,N_4842);
nand U5004 (N_5004,N_4507,N_4925);
and U5005 (N_5005,N_4603,N_4540);
nand U5006 (N_5006,N_4750,N_4653);
nor U5007 (N_5007,N_4831,N_4773);
nor U5008 (N_5008,N_4965,N_4664);
or U5009 (N_5009,N_4835,N_4997);
nand U5010 (N_5010,N_4865,N_4607);
or U5011 (N_5011,N_4912,N_4524);
nor U5012 (N_5012,N_4646,N_4798);
and U5013 (N_5013,N_4875,N_4864);
or U5014 (N_5014,N_4545,N_4849);
or U5015 (N_5015,N_4819,N_4719);
nor U5016 (N_5016,N_4906,N_4928);
and U5017 (N_5017,N_4574,N_4728);
nor U5018 (N_5018,N_4971,N_4960);
nand U5019 (N_5019,N_4886,N_4887);
nor U5020 (N_5020,N_4983,N_4876);
and U5021 (N_5021,N_4624,N_4878);
xnor U5022 (N_5022,N_4921,N_4527);
nand U5023 (N_5023,N_4844,N_4872);
xnor U5024 (N_5024,N_4643,N_4622);
nand U5025 (N_5025,N_4775,N_4947);
and U5026 (N_5026,N_4706,N_4771);
xnor U5027 (N_5027,N_4594,N_4924);
nand U5028 (N_5028,N_4525,N_4929);
and U5029 (N_5029,N_4609,N_4592);
and U5030 (N_5030,N_4587,N_4569);
and U5031 (N_5031,N_4568,N_4591);
nor U5032 (N_5032,N_4923,N_4563);
nor U5033 (N_5033,N_4825,N_4927);
or U5034 (N_5034,N_4789,N_4623);
xnor U5035 (N_5035,N_4804,N_4920);
xor U5036 (N_5036,N_4790,N_4754);
nor U5037 (N_5037,N_4704,N_4839);
and U5038 (N_5038,N_4767,N_4584);
and U5039 (N_5039,N_4846,N_4548);
xnor U5040 (N_5040,N_4717,N_4940);
xnor U5041 (N_5041,N_4630,N_4772);
and U5042 (N_5042,N_4820,N_4816);
or U5043 (N_5043,N_4894,N_4691);
nor U5044 (N_5044,N_4583,N_4784);
xor U5045 (N_5045,N_4963,N_4892);
nor U5046 (N_5046,N_4575,N_4870);
xor U5047 (N_5047,N_4905,N_4654);
and U5048 (N_5048,N_4559,N_4700);
and U5049 (N_5049,N_4671,N_4600);
xnor U5050 (N_5050,N_4838,N_4703);
or U5051 (N_5051,N_4514,N_4791);
or U5052 (N_5052,N_4991,N_4686);
or U5053 (N_5053,N_4557,N_4948);
nand U5054 (N_5054,N_4943,N_4737);
or U5055 (N_5055,N_4663,N_4582);
and U5056 (N_5056,N_4796,N_4736);
and U5057 (N_5057,N_4677,N_4951);
or U5058 (N_5058,N_4797,N_4627);
and U5059 (N_5059,N_4861,N_4828);
nor U5060 (N_5060,N_4708,N_4946);
nand U5061 (N_5061,N_4644,N_4682);
and U5062 (N_5062,N_4958,N_4765);
xnor U5063 (N_5063,N_4778,N_4652);
nor U5064 (N_5064,N_4513,N_4818);
nor U5065 (N_5065,N_4919,N_4730);
and U5066 (N_5066,N_4724,N_4942);
nor U5067 (N_5067,N_4638,N_4933);
xor U5068 (N_5068,N_4841,N_4670);
nand U5069 (N_5069,N_4764,N_4648);
nand U5070 (N_5070,N_4815,N_4571);
and U5071 (N_5071,N_4610,N_4823);
xor U5072 (N_5072,N_4679,N_4562);
nand U5073 (N_5073,N_4649,N_4783);
nor U5074 (N_5074,N_4745,N_4873);
or U5075 (N_5075,N_4890,N_4877);
nand U5076 (N_5076,N_4751,N_4732);
nor U5077 (N_5077,N_4689,N_4697);
nor U5078 (N_5078,N_4599,N_4589);
nor U5079 (N_5079,N_4911,N_4544);
or U5080 (N_5080,N_4945,N_4860);
xor U5081 (N_5081,N_4547,N_4981);
or U5082 (N_5082,N_4519,N_4803);
nor U5083 (N_5083,N_4554,N_4931);
nor U5084 (N_5084,N_4883,N_4917);
xnor U5085 (N_5085,N_4802,N_4982);
nand U5086 (N_5086,N_4807,N_4901);
or U5087 (N_5087,N_4505,N_4684);
xor U5088 (N_5088,N_4725,N_4535);
nand U5089 (N_5089,N_4998,N_4749);
nand U5090 (N_5090,N_4673,N_4961);
nor U5091 (N_5091,N_4659,N_4521);
nor U5092 (N_5092,N_4884,N_4969);
nand U5093 (N_5093,N_4989,N_4687);
and U5094 (N_5094,N_4962,N_4821);
nand U5095 (N_5095,N_4692,N_4693);
xnor U5096 (N_5096,N_4613,N_4944);
nand U5097 (N_5097,N_4848,N_4702);
nor U5098 (N_5098,N_4777,N_4629);
nor U5099 (N_5099,N_4738,N_4851);
xnor U5100 (N_5100,N_4561,N_4635);
and U5101 (N_5101,N_4832,N_4556);
nand U5102 (N_5102,N_4529,N_4874);
nand U5103 (N_5103,N_4502,N_4531);
xor U5104 (N_5104,N_4770,N_4900);
nand U5105 (N_5105,N_4827,N_4722);
nand U5106 (N_5106,N_4840,N_4782);
and U5107 (N_5107,N_4723,N_4896);
nand U5108 (N_5108,N_4898,N_4938);
or U5109 (N_5109,N_4551,N_4579);
nor U5110 (N_5110,N_4585,N_4760);
nor U5111 (N_5111,N_4808,N_4862);
nor U5112 (N_5112,N_4987,N_4726);
nor U5113 (N_5113,N_4537,N_4633);
and U5114 (N_5114,N_4941,N_4731);
xnor U5115 (N_5115,N_4979,N_4956);
or U5116 (N_5116,N_4993,N_4758);
or U5117 (N_5117,N_4665,N_4578);
and U5118 (N_5118,N_4647,N_4867);
nand U5119 (N_5119,N_4833,N_4939);
or U5120 (N_5120,N_4739,N_4996);
xnor U5121 (N_5121,N_4553,N_4666);
and U5122 (N_5122,N_4757,N_4805);
nand U5123 (N_5123,N_4716,N_4893);
and U5124 (N_5124,N_4918,N_4904);
xnor U5125 (N_5125,N_4588,N_4786);
nor U5126 (N_5126,N_4955,N_4645);
nor U5127 (N_5127,N_4552,N_4964);
nor U5128 (N_5128,N_4605,N_4581);
xor U5129 (N_5129,N_4992,N_4512);
nor U5130 (N_5130,N_4658,N_4970);
and U5131 (N_5131,N_4680,N_4573);
and U5132 (N_5132,N_4856,N_4576);
nand U5133 (N_5133,N_4761,N_4834);
nand U5134 (N_5134,N_4566,N_4994);
or U5135 (N_5135,N_4766,N_4972);
xnor U5136 (N_5136,N_4657,N_4735);
nand U5137 (N_5137,N_4685,N_4888);
xnor U5138 (N_5138,N_4558,N_4715);
nor U5139 (N_5139,N_4678,N_4601);
xor U5140 (N_5140,N_4866,N_4619);
and U5141 (N_5141,N_4616,N_4967);
and U5142 (N_5142,N_4595,N_4880);
xor U5143 (N_5143,N_4549,N_4759);
and U5144 (N_5144,N_4564,N_4500);
nor U5145 (N_5145,N_4534,N_4694);
xnor U5146 (N_5146,N_4885,N_4640);
nand U5147 (N_5147,N_4533,N_4953);
nand U5148 (N_5148,N_4668,N_4968);
nor U5149 (N_5149,N_4596,N_4800);
nor U5150 (N_5150,N_4632,N_4621);
or U5151 (N_5151,N_4546,N_4625);
nor U5152 (N_5152,N_4871,N_4597);
or U5153 (N_5153,N_4516,N_4812);
xor U5154 (N_5154,N_4853,N_4515);
or U5155 (N_5155,N_4781,N_4614);
xor U5156 (N_5156,N_4949,N_4727);
or U5157 (N_5157,N_4857,N_4980);
xor U5158 (N_5158,N_4879,N_4526);
nor U5159 (N_5159,N_4520,N_4889);
xnor U5160 (N_5160,N_4631,N_4608);
nand U5161 (N_5161,N_4711,N_4538);
xnor U5162 (N_5162,N_4822,N_4916);
nor U5163 (N_5163,N_4617,N_4744);
nand U5164 (N_5164,N_4743,N_4674);
and U5165 (N_5165,N_4714,N_4701);
or U5166 (N_5166,N_4984,N_4952);
xor U5167 (N_5167,N_4934,N_4746);
nor U5168 (N_5168,N_4586,N_4620);
or U5169 (N_5169,N_4713,N_4530);
nor U5170 (N_5170,N_4604,N_4902);
or U5171 (N_5171,N_4779,N_4672);
nand U5172 (N_5172,N_4854,N_4935);
nand U5173 (N_5173,N_4976,N_4895);
or U5174 (N_5174,N_4999,N_4626);
and U5175 (N_5175,N_4826,N_4830);
xor U5176 (N_5176,N_4705,N_4903);
nand U5177 (N_5177,N_4528,N_4813);
nand U5178 (N_5178,N_4618,N_4748);
xnor U5179 (N_5179,N_4932,N_4506);
nor U5180 (N_5180,N_4504,N_4541);
xnor U5181 (N_5181,N_4661,N_4909);
or U5182 (N_5182,N_4740,N_4690);
nor U5183 (N_5183,N_4995,N_4795);
and U5184 (N_5184,N_4660,N_4676);
xor U5185 (N_5185,N_4794,N_4628);
and U5186 (N_5186,N_4733,N_4852);
or U5187 (N_5187,N_4710,N_4780);
xnor U5188 (N_5188,N_4642,N_4509);
or U5189 (N_5189,N_4988,N_4845);
xnor U5190 (N_5190,N_4712,N_4926);
xnor U5191 (N_5191,N_4606,N_4639);
nor U5192 (N_5192,N_4763,N_4667);
nand U5193 (N_5193,N_4824,N_4572);
and U5194 (N_5194,N_4651,N_4914);
or U5195 (N_5195,N_4899,N_4774);
nand U5196 (N_5196,N_4729,N_4847);
and U5197 (N_5197,N_4580,N_4570);
nand U5198 (N_5198,N_4501,N_4954);
nand U5199 (N_5199,N_4810,N_4806);
nand U5200 (N_5200,N_4734,N_4709);
and U5201 (N_5201,N_4937,N_4721);
xor U5202 (N_5202,N_4836,N_4550);
or U5203 (N_5203,N_4699,N_4542);
and U5204 (N_5204,N_4532,N_4762);
xnor U5205 (N_5205,N_4590,N_4656);
nor U5206 (N_5206,N_4641,N_4753);
nand U5207 (N_5207,N_4650,N_4897);
nor U5208 (N_5208,N_4882,N_4755);
nor U5209 (N_5209,N_4913,N_4907);
and U5210 (N_5210,N_4817,N_4869);
nand U5211 (N_5211,N_4611,N_4522);
or U5212 (N_5212,N_4776,N_4855);
or U5213 (N_5213,N_4742,N_4688);
nand U5214 (N_5214,N_4787,N_4747);
and U5215 (N_5215,N_4503,N_4799);
and U5216 (N_5216,N_4850,N_4669);
or U5217 (N_5217,N_4966,N_4752);
xnor U5218 (N_5218,N_4959,N_4577);
nor U5219 (N_5219,N_4510,N_4859);
nor U5220 (N_5220,N_4560,N_4977);
and U5221 (N_5221,N_4974,N_4837);
nor U5222 (N_5222,N_4565,N_4636);
or U5223 (N_5223,N_4695,N_4655);
and U5224 (N_5224,N_4922,N_4718);
xnor U5225 (N_5225,N_4868,N_4788);
xnor U5226 (N_5226,N_4518,N_4891);
nand U5227 (N_5227,N_4612,N_4792);
xnor U5228 (N_5228,N_4769,N_4881);
and U5229 (N_5229,N_4950,N_4829);
nand U5230 (N_5230,N_4536,N_4508);
nor U5231 (N_5231,N_4978,N_4681);
nor U5232 (N_5232,N_4908,N_4602);
nor U5233 (N_5233,N_4985,N_4675);
and U5234 (N_5234,N_4801,N_4975);
and U5235 (N_5235,N_4523,N_4915);
or U5236 (N_5236,N_4986,N_4863);
xor U5237 (N_5237,N_4637,N_4615);
nand U5238 (N_5238,N_4683,N_4698);
xor U5239 (N_5239,N_4957,N_4555);
and U5240 (N_5240,N_4696,N_4936);
xor U5241 (N_5241,N_4990,N_4814);
and U5242 (N_5242,N_4785,N_4811);
or U5243 (N_5243,N_4809,N_4843);
nor U5244 (N_5244,N_4567,N_4662);
xnor U5245 (N_5245,N_4741,N_4973);
and U5246 (N_5246,N_4768,N_4539);
xor U5247 (N_5247,N_4517,N_4720);
xor U5248 (N_5248,N_4793,N_4910);
nor U5249 (N_5249,N_4593,N_4756);
or U5250 (N_5250,N_4529,N_4857);
xor U5251 (N_5251,N_4631,N_4709);
xor U5252 (N_5252,N_4558,N_4828);
xnor U5253 (N_5253,N_4503,N_4690);
and U5254 (N_5254,N_4841,N_4886);
or U5255 (N_5255,N_4661,N_4621);
xnor U5256 (N_5256,N_4983,N_4840);
xor U5257 (N_5257,N_4630,N_4959);
nand U5258 (N_5258,N_4827,N_4795);
nand U5259 (N_5259,N_4996,N_4582);
nor U5260 (N_5260,N_4822,N_4772);
nor U5261 (N_5261,N_4980,N_4554);
nor U5262 (N_5262,N_4739,N_4586);
nor U5263 (N_5263,N_4842,N_4902);
and U5264 (N_5264,N_4749,N_4853);
and U5265 (N_5265,N_4571,N_4814);
nor U5266 (N_5266,N_4581,N_4652);
or U5267 (N_5267,N_4924,N_4527);
and U5268 (N_5268,N_4606,N_4988);
xnor U5269 (N_5269,N_4655,N_4850);
and U5270 (N_5270,N_4545,N_4831);
and U5271 (N_5271,N_4822,N_4919);
or U5272 (N_5272,N_4563,N_4759);
nor U5273 (N_5273,N_4680,N_4907);
and U5274 (N_5274,N_4600,N_4978);
nand U5275 (N_5275,N_4750,N_4787);
and U5276 (N_5276,N_4620,N_4780);
and U5277 (N_5277,N_4933,N_4775);
and U5278 (N_5278,N_4629,N_4618);
and U5279 (N_5279,N_4558,N_4726);
or U5280 (N_5280,N_4930,N_4548);
or U5281 (N_5281,N_4844,N_4623);
xor U5282 (N_5282,N_4913,N_4533);
and U5283 (N_5283,N_4516,N_4756);
xor U5284 (N_5284,N_4825,N_4881);
nor U5285 (N_5285,N_4692,N_4522);
or U5286 (N_5286,N_4673,N_4680);
xnor U5287 (N_5287,N_4572,N_4775);
and U5288 (N_5288,N_4988,N_4930);
nor U5289 (N_5289,N_4931,N_4922);
nand U5290 (N_5290,N_4965,N_4514);
and U5291 (N_5291,N_4766,N_4700);
and U5292 (N_5292,N_4659,N_4730);
nand U5293 (N_5293,N_4618,N_4669);
xor U5294 (N_5294,N_4719,N_4868);
xor U5295 (N_5295,N_4892,N_4693);
xor U5296 (N_5296,N_4648,N_4623);
xor U5297 (N_5297,N_4644,N_4904);
or U5298 (N_5298,N_4843,N_4962);
or U5299 (N_5299,N_4828,N_4680);
xor U5300 (N_5300,N_4645,N_4710);
xnor U5301 (N_5301,N_4964,N_4594);
xor U5302 (N_5302,N_4765,N_4666);
xnor U5303 (N_5303,N_4543,N_4630);
nor U5304 (N_5304,N_4543,N_4566);
xnor U5305 (N_5305,N_4540,N_4902);
xnor U5306 (N_5306,N_4926,N_4693);
nand U5307 (N_5307,N_4789,N_4669);
xor U5308 (N_5308,N_4929,N_4589);
and U5309 (N_5309,N_4991,N_4511);
nand U5310 (N_5310,N_4856,N_4665);
or U5311 (N_5311,N_4755,N_4974);
nor U5312 (N_5312,N_4749,N_4985);
nor U5313 (N_5313,N_4887,N_4743);
and U5314 (N_5314,N_4864,N_4843);
xor U5315 (N_5315,N_4687,N_4652);
or U5316 (N_5316,N_4637,N_4547);
nor U5317 (N_5317,N_4527,N_4707);
xnor U5318 (N_5318,N_4751,N_4552);
xor U5319 (N_5319,N_4735,N_4881);
nand U5320 (N_5320,N_4925,N_4622);
nor U5321 (N_5321,N_4895,N_4527);
and U5322 (N_5322,N_4956,N_4968);
xnor U5323 (N_5323,N_4534,N_4758);
xor U5324 (N_5324,N_4557,N_4598);
xor U5325 (N_5325,N_4660,N_4704);
or U5326 (N_5326,N_4733,N_4700);
xnor U5327 (N_5327,N_4769,N_4997);
xor U5328 (N_5328,N_4763,N_4844);
nor U5329 (N_5329,N_4830,N_4557);
and U5330 (N_5330,N_4696,N_4900);
nand U5331 (N_5331,N_4582,N_4965);
and U5332 (N_5332,N_4924,N_4566);
and U5333 (N_5333,N_4705,N_4652);
xor U5334 (N_5334,N_4820,N_4718);
or U5335 (N_5335,N_4617,N_4971);
and U5336 (N_5336,N_4835,N_4918);
nand U5337 (N_5337,N_4548,N_4808);
xor U5338 (N_5338,N_4624,N_4906);
xnor U5339 (N_5339,N_4659,N_4545);
or U5340 (N_5340,N_4685,N_4945);
and U5341 (N_5341,N_4622,N_4905);
nand U5342 (N_5342,N_4934,N_4785);
or U5343 (N_5343,N_4821,N_4690);
xnor U5344 (N_5344,N_4745,N_4879);
and U5345 (N_5345,N_4536,N_4741);
or U5346 (N_5346,N_4710,N_4945);
nor U5347 (N_5347,N_4580,N_4662);
xnor U5348 (N_5348,N_4921,N_4891);
xnor U5349 (N_5349,N_4891,N_4893);
nor U5350 (N_5350,N_4676,N_4722);
nand U5351 (N_5351,N_4684,N_4695);
and U5352 (N_5352,N_4666,N_4677);
or U5353 (N_5353,N_4747,N_4943);
and U5354 (N_5354,N_4759,N_4949);
and U5355 (N_5355,N_4784,N_4530);
xor U5356 (N_5356,N_4851,N_4528);
nand U5357 (N_5357,N_4681,N_4523);
or U5358 (N_5358,N_4776,N_4758);
nor U5359 (N_5359,N_4521,N_4625);
xnor U5360 (N_5360,N_4871,N_4648);
or U5361 (N_5361,N_4561,N_4804);
nor U5362 (N_5362,N_4614,N_4664);
nor U5363 (N_5363,N_4746,N_4794);
and U5364 (N_5364,N_4730,N_4666);
xnor U5365 (N_5365,N_4976,N_4512);
xnor U5366 (N_5366,N_4507,N_4853);
nor U5367 (N_5367,N_4984,N_4545);
xor U5368 (N_5368,N_4978,N_4856);
nor U5369 (N_5369,N_4645,N_4521);
nor U5370 (N_5370,N_4541,N_4994);
nor U5371 (N_5371,N_4806,N_4876);
nand U5372 (N_5372,N_4742,N_4689);
or U5373 (N_5373,N_4657,N_4768);
nand U5374 (N_5374,N_4756,N_4500);
xnor U5375 (N_5375,N_4614,N_4915);
xor U5376 (N_5376,N_4726,N_4644);
nor U5377 (N_5377,N_4584,N_4799);
or U5378 (N_5378,N_4603,N_4552);
xnor U5379 (N_5379,N_4714,N_4568);
nand U5380 (N_5380,N_4899,N_4896);
xnor U5381 (N_5381,N_4632,N_4879);
or U5382 (N_5382,N_4580,N_4504);
xor U5383 (N_5383,N_4657,N_4501);
or U5384 (N_5384,N_4802,N_4986);
nor U5385 (N_5385,N_4621,N_4708);
nand U5386 (N_5386,N_4719,N_4610);
xnor U5387 (N_5387,N_4704,N_4576);
or U5388 (N_5388,N_4581,N_4941);
xnor U5389 (N_5389,N_4950,N_4567);
xnor U5390 (N_5390,N_4514,N_4970);
nand U5391 (N_5391,N_4642,N_4750);
xnor U5392 (N_5392,N_4888,N_4919);
nor U5393 (N_5393,N_4754,N_4930);
or U5394 (N_5394,N_4860,N_4528);
and U5395 (N_5395,N_4951,N_4997);
nand U5396 (N_5396,N_4968,N_4678);
xor U5397 (N_5397,N_4702,N_4589);
nand U5398 (N_5398,N_4745,N_4730);
nand U5399 (N_5399,N_4528,N_4726);
and U5400 (N_5400,N_4665,N_4684);
nand U5401 (N_5401,N_4982,N_4563);
xor U5402 (N_5402,N_4857,N_4633);
nor U5403 (N_5403,N_4984,N_4692);
or U5404 (N_5404,N_4619,N_4825);
or U5405 (N_5405,N_4874,N_4559);
or U5406 (N_5406,N_4946,N_4997);
xnor U5407 (N_5407,N_4714,N_4954);
xor U5408 (N_5408,N_4969,N_4525);
nor U5409 (N_5409,N_4736,N_4873);
or U5410 (N_5410,N_4915,N_4694);
nor U5411 (N_5411,N_4981,N_4649);
and U5412 (N_5412,N_4705,N_4860);
or U5413 (N_5413,N_4741,N_4818);
xnor U5414 (N_5414,N_4705,N_4516);
or U5415 (N_5415,N_4764,N_4743);
nand U5416 (N_5416,N_4683,N_4807);
nand U5417 (N_5417,N_4683,N_4905);
nor U5418 (N_5418,N_4612,N_4659);
xnor U5419 (N_5419,N_4721,N_4986);
nor U5420 (N_5420,N_4761,N_4757);
or U5421 (N_5421,N_4942,N_4763);
nor U5422 (N_5422,N_4942,N_4506);
and U5423 (N_5423,N_4736,N_4916);
nand U5424 (N_5424,N_4590,N_4692);
nor U5425 (N_5425,N_4849,N_4881);
xnor U5426 (N_5426,N_4772,N_4985);
nor U5427 (N_5427,N_4892,N_4937);
or U5428 (N_5428,N_4528,N_4550);
nand U5429 (N_5429,N_4585,N_4785);
xnor U5430 (N_5430,N_4694,N_4850);
or U5431 (N_5431,N_4796,N_4764);
and U5432 (N_5432,N_4948,N_4806);
nand U5433 (N_5433,N_4913,N_4938);
nor U5434 (N_5434,N_4659,N_4917);
nand U5435 (N_5435,N_4597,N_4823);
nor U5436 (N_5436,N_4593,N_4674);
or U5437 (N_5437,N_4543,N_4999);
nand U5438 (N_5438,N_4536,N_4930);
nand U5439 (N_5439,N_4896,N_4533);
nor U5440 (N_5440,N_4566,N_4685);
and U5441 (N_5441,N_4796,N_4929);
xnor U5442 (N_5442,N_4999,N_4996);
and U5443 (N_5443,N_4595,N_4665);
nor U5444 (N_5444,N_4608,N_4521);
or U5445 (N_5445,N_4907,N_4876);
nand U5446 (N_5446,N_4981,N_4821);
nand U5447 (N_5447,N_4583,N_4518);
and U5448 (N_5448,N_4553,N_4531);
nand U5449 (N_5449,N_4647,N_4859);
xor U5450 (N_5450,N_4555,N_4855);
nand U5451 (N_5451,N_4598,N_4682);
nor U5452 (N_5452,N_4564,N_4740);
nand U5453 (N_5453,N_4777,N_4752);
and U5454 (N_5454,N_4623,N_4781);
nor U5455 (N_5455,N_4636,N_4969);
nor U5456 (N_5456,N_4889,N_4663);
nor U5457 (N_5457,N_4977,N_4631);
and U5458 (N_5458,N_4517,N_4850);
nand U5459 (N_5459,N_4801,N_4967);
nor U5460 (N_5460,N_4630,N_4906);
xor U5461 (N_5461,N_4625,N_4866);
nand U5462 (N_5462,N_4516,N_4807);
or U5463 (N_5463,N_4955,N_4517);
nand U5464 (N_5464,N_4735,N_4829);
and U5465 (N_5465,N_4631,N_4841);
nand U5466 (N_5466,N_4897,N_4766);
xnor U5467 (N_5467,N_4560,N_4621);
and U5468 (N_5468,N_4724,N_4659);
nand U5469 (N_5469,N_4820,N_4570);
or U5470 (N_5470,N_4721,N_4839);
and U5471 (N_5471,N_4744,N_4756);
nor U5472 (N_5472,N_4695,N_4585);
and U5473 (N_5473,N_4902,N_4769);
or U5474 (N_5474,N_4772,N_4698);
xnor U5475 (N_5475,N_4857,N_4527);
xor U5476 (N_5476,N_4972,N_4669);
and U5477 (N_5477,N_4893,N_4578);
or U5478 (N_5478,N_4514,N_4657);
nor U5479 (N_5479,N_4854,N_4645);
nor U5480 (N_5480,N_4892,N_4817);
nor U5481 (N_5481,N_4934,N_4878);
nor U5482 (N_5482,N_4510,N_4990);
or U5483 (N_5483,N_4876,N_4909);
nor U5484 (N_5484,N_4874,N_4761);
nor U5485 (N_5485,N_4667,N_4969);
and U5486 (N_5486,N_4772,N_4914);
and U5487 (N_5487,N_4696,N_4848);
or U5488 (N_5488,N_4954,N_4711);
or U5489 (N_5489,N_4950,N_4655);
nand U5490 (N_5490,N_4608,N_4731);
xor U5491 (N_5491,N_4521,N_4813);
or U5492 (N_5492,N_4915,N_4998);
xnor U5493 (N_5493,N_4626,N_4699);
or U5494 (N_5494,N_4582,N_4706);
nand U5495 (N_5495,N_4950,N_4642);
nor U5496 (N_5496,N_4615,N_4995);
nor U5497 (N_5497,N_4508,N_4991);
or U5498 (N_5498,N_4862,N_4638);
nor U5499 (N_5499,N_4881,N_4917);
nor U5500 (N_5500,N_5435,N_5393);
or U5501 (N_5501,N_5185,N_5402);
or U5502 (N_5502,N_5007,N_5036);
or U5503 (N_5503,N_5060,N_5113);
nor U5504 (N_5504,N_5129,N_5433);
and U5505 (N_5505,N_5035,N_5451);
and U5506 (N_5506,N_5398,N_5331);
nor U5507 (N_5507,N_5055,N_5464);
nand U5508 (N_5508,N_5071,N_5133);
and U5509 (N_5509,N_5267,N_5021);
nor U5510 (N_5510,N_5265,N_5008);
or U5511 (N_5511,N_5458,N_5088);
or U5512 (N_5512,N_5198,N_5170);
xnor U5513 (N_5513,N_5274,N_5015);
or U5514 (N_5514,N_5406,N_5281);
and U5515 (N_5515,N_5394,N_5273);
nor U5516 (N_5516,N_5243,N_5352);
xor U5517 (N_5517,N_5335,N_5030);
and U5518 (N_5518,N_5364,N_5200);
or U5519 (N_5519,N_5090,N_5130);
nor U5520 (N_5520,N_5147,N_5315);
and U5521 (N_5521,N_5428,N_5468);
nor U5522 (N_5522,N_5410,N_5320);
xor U5523 (N_5523,N_5403,N_5239);
and U5524 (N_5524,N_5095,N_5100);
xor U5525 (N_5525,N_5348,N_5152);
nand U5526 (N_5526,N_5268,N_5411);
and U5527 (N_5527,N_5231,N_5233);
nor U5528 (N_5528,N_5103,N_5077);
xor U5529 (N_5529,N_5079,N_5010);
and U5530 (N_5530,N_5087,N_5238);
and U5531 (N_5531,N_5374,N_5346);
nand U5532 (N_5532,N_5380,N_5080);
xnor U5533 (N_5533,N_5298,N_5156);
xor U5534 (N_5534,N_5167,N_5391);
nor U5535 (N_5535,N_5277,N_5019);
xnor U5536 (N_5536,N_5182,N_5025);
nand U5537 (N_5537,N_5323,N_5251);
nand U5538 (N_5538,N_5086,N_5122);
nand U5539 (N_5539,N_5199,N_5023);
and U5540 (N_5540,N_5221,N_5295);
or U5541 (N_5541,N_5218,N_5442);
and U5542 (N_5542,N_5191,N_5165);
or U5543 (N_5543,N_5017,N_5214);
nor U5544 (N_5544,N_5001,N_5487);
and U5545 (N_5545,N_5121,N_5118);
and U5546 (N_5546,N_5284,N_5498);
and U5547 (N_5547,N_5259,N_5094);
or U5548 (N_5548,N_5353,N_5407);
nand U5549 (N_5549,N_5369,N_5461);
nor U5550 (N_5550,N_5249,N_5057);
xnor U5551 (N_5551,N_5151,N_5232);
xor U5552 (N_5552,N_5494,N_5479);
nor U5553 (N_5553,N_5042,N_5341);
nand U5554 (N_5554,N_5116,N_5083);
or U5555 (N_5555,N_5271,N_5179);
nor U5556 (N_5556,N_5467,N_5423);
xor U5557 (N_5557,N_5029,N_5386);
xnor U5558 (N_5558,N_5171,N_5050);
nand U5559 (N_5559,N_5127,N_5375);
or U5560 (N_5560,N_5154,N_5046);
xor U5561 (N_5561,N_5356,N_5110);
nand U5562 (N_5562,N_5054,N_5104);
nand U5563 (N_5563,N_5308,N_5430);
nand U5564 (N_5564,N_5157,N_5400);
or U5565 (N_5565,N_5260,N_5324);
and U5566 (N_5566,N_5220,N_5318);
nor U5567 (N_5567,N_5416,N_5262);
nand U5568 (N_5568,N_5219,N_5016);
nor U5569 (N_5569,N_5026,N_5443);
nor U5570 (N_5570,N_5244,N_5293);
xor U5571 (N_5571,N_5449,N_5068);
nand U5572 (N_5572,N_5377,N_5186);
xnor U5573 (N_5573,N_5414,N_5033);
xor U5574 (N_5574,N_5076,N_5074);
and U5575 (N_5575,N_5256,N_5045);
and U5576 (N_5576,N_5304,N_5114);
and U5577 (N_5577,N_5063,N_5477);
or U5578 (N_5578,N_5497,N_5344);
and U5579 (N_5579,N_5067,N_5302);
or U5580 (N_5580,N_5062,N_5491);
or U5581 (N_5581,N_5069,N_5206);
nand U5582 (N_5582,N_5290,N_5164);
or U5583 (N_5583,N_5405,N_5031);
xnor U5584 (N_5584,N_5078,N_5203);
or U5585 (N_5585,N_5455,N_5395);
xor U5586 (N_5586,N_5229,N_5466);
and U5587 (N_5587,N_5120,N_5371);
xor U5588 (N_5588,N_5447,N_5043);
and U5589 (N_5589,N_5176,N_5081);
and U5590 (N_5590,N_5034,N_5059);
xnor U5591 (N_5591,N_5246,N_5459);
nor U5592 (N_5592,N_5044,N_5223);
and U5593 (N_5593,N_5299,N_5276);
nor U5594 (N_5594,N_5099,N_5119);
or U5595 (N_5595,N_5453,N_5158);
xnor U5596 (N_5596,N_5205,N_5480);
nor U5597 (N_5597,N_5495,N_5193);
nand U5598 (N_5598,N_5338,N_5061);
or U5599 (N_5599,N_5000,N_5485);
or U5600 (N_5600,N_5162,N_5013);
xor U5601 (N_5601,N_5316,N_5149);
or U5602 (N_5602,N_5161,N_5066);
nand U5603 (N_5603,N_5228,N_5250);
nand U5604 (N_5604,N_5038,N_5195);
and U5605 (N_5605,N_5384,N_5392);
and U5606 (N_5606,N_5311,N_5349);
and U5607 (N_5607,N_5388,N_5148);
or U5608 (N_5608,N_5201,N_5168);
nor U5609 (N_5609,N_5396,N_5093);
xor U5610 (N_5610,N_5385,N_5009);
nand U5611 (N_5611,N_5240,N_5286);
nand U5612 (N_5612,N_5270,N_5209);
nor U5613 (N_5613,N_5360,N_5145);
xor U5614 (N_5614,N_5269,N_5471);
and U5615 (N_5615,N_5436,N_5051);
xor U5616 (N_5616,N_5247,N_5415);
nand U5617 (N_5617,N_5465,N_5470);
xnor U5618 (N_5618,N_5215,N_5355);
xor U5619 (N_5619,N_5106,N_5330);
and U5620 (N_5620,N_5279,N_5175);
nand U5621 (N_5621,N_5383,N_5413);
or U5622 (N_5622,N_5289,N_5022);
or U5623 (N_5623,N_5091,N_5417);
xnor U5624 (N_5624,N_5217,N_5139);
xor U5625 (N_5625,N_5359,N_5301);
nor U5626 (N_5626,N_5048,N_5202);
xor U5627 (N_5627,N_5303,N_5213);
xnor U5628 (N_5628,N_5150,N_5365);
xor U5629 (N_5629,N_5125,N_5446);
xor U5630 (N_5630,N_5160,N_5112);
nand U5631 (N_5631,N_5257,N_5437);
nand U5632 (N_5632,N_5474,N_5463);
xor U5633 (N_5633,N_5389,N_5155);
xnor U5634 (N_5634,N_5387,N_5362);
xor U5635 (N_5635,N_5325,N_5439);
or U5636 (N_5636,N_5272,N_5336);
xor U5637 (N_5637,N_5137,N_5313);
and U5638 (N_5638,N_5163,N_5254);
nor U5639 (N_5639,N_5107,N_5224);
nor U5640 (N_5640,N_5169,N_5288);
and U5641 (N_5641,N_5138,N_5089);
and U5642 (N_5642,N_5366,N_5492);
or U5643 (N_5643,N_5018,N_5342);
nor U5644 (N_5644,N_5327,N_5136);
nand U5645 (N_5645,N_5431,N_5404);
nand U5646 (N_5646,N_5053,N_5172);
and U5647 (N_5647,N_5073,N_5141);
and U5648 (N_5648,N_5332,N_5230);
nor U5649 (N_5649,N_5222,N_5280);
nor U5650 (N_5650,N_5351,N_5420);
and U5651 (N_5651,N_5204,N_5032);
nor U5652 (N_5652,N_5134,N_5027);
or U5653 (N_5653,N_5159,N_5181);
and U5654 (N_5654,N_5419,N_5135);
or U5655 (N_5655,N_5367,N_5292);
nand U5656 (N_5656,N_5006,N_5020);
nand U5657 (N_5657,N_5226,N_5343);
or U5658 (N_5658,N_5372,N_5421);
nor U5659 (N_5659,N_5258,N_5399);
nand U5660 (N_5660,N_5197,N_5475);
nor U5661 (N_5661,N_5339,N_5300);
nor U5662 (N_5662,N_5340,N_5337);
nand U5663 (N_5663,N_5212,N_5049);
and U5664 (N_5664,N_5422,N_5306);
nor U5665 (N_5665,N_5357,N_5275);
or U5666 (N_5666,N_5363,N_5287);
xnor U5667 (N_5667,N_5153,N_5005);
nand U5668 (N_5668,N_5473,N_5345);
xor U5669 (N_5669,N_5216,N_5333);
xnor U5670 (N_5670,N_5028,N_5483);
or U5671 (N_5671,N_5143,N_5187);
and U5672 (N_5672,N_5312,N_5040);
xor U5673 (N_5673,N_5462,N_5314);
nor U5674 (N_5674,N_5370,N_5450);
xor U5675 (N_5675,N_5285,N_5457);
and U5676 (N_5676,N_5438,N_5358);
nand U5677 (N_5677,N_5291,N_5058);
xor U5678 (N_5678,N_5004,N_5310);
or U5679 (N_5679,N_5052,N_5378);
or U5680 (N_5680,N_5486,N_5101);
xor U5681 (N_5681,N_5178,N_5041);
nand U5682 (N_5682,N_5166,N_5441);
nand U5683 (N_5683,N_5490,N_5070);
or U5684 (N_5684,N_5266,N_5064);
nor U5685 (N_5685,N_5444,N_5253);
or U5686 (N_5686,N_5242,N_5211);
or U5687 (N_5687,N_5011,N_5472);
or U5688 (N_5688,N_5173,N_5123);
and U5689 (N_5689,N_5207,N_5322);
nor U5690 (N_5690,N_5452,N_5499);
xor U5691 (N_5691,N_5189,N_5037);
nand U5692 (N_5692,N_5194,N_5482);
nor U5693 (N_5693,N_5192,N_5084);
nand U5694 (N_5694,N_5361,N_5108);
xor U5695 (N_5695,N_5196,N_5177);
xor U5696 (N_5696,N_5460,N_5319);
or U5697 (N_5697,N_5075,N_5124);
nor U5698 (N_5698,N_5117,N_5003);
nand U5699 (N_5699,N_5245,N_5131);
nor U5700 (N_5700,N_5328,N_5132);
nand U5701 (N_5701,N_5115,N_5329);
nand U5702 (N_5702,N_5282,N_5376);
and U5703 (N_5703,N_5448,N_5190);
xnor U5704 (N_5704,N_5085,N_5255);
and U5705 (N_5705,N_5082,N_5373);
nand U5706 (N_5706,N_5401,N_5296);
and U5707 (N_5707,N_5309,N_5305);
xor U5708 (N_5708,N_5484,N_5261);
xnor U5709 (N_5709,N_5334,N_5183);
nand U5710 (N_5710,N_5140,N_5409);
nand U5711 (N_5711,N_5412,N_5263);
xnor U5712 (N_5712,N_5469,N_5111);
xnor U5713 (N_5713,N_5126,N_5012);
nor U5714 (N_5714,N_5368,N_5208);
or U5715 (N_5715,N_5264,N_5321);
or U5716 (N_5716,N_5235,N_5184);
nand U5717 (N_5717,N_5489,N_5252);
nand U5718 (N_5718,N_5476,N_5426);
and U5719 (N_5719,N_5237,N_5096);
xor U5720 (N_5720,N_5379,N_5105);
nand U5721 (N_5721,N_5072,N_5481);
nand U5722 (N_5722,N_5180,N_5174);
nor U5723 (N_5723,N_5496,N_5456);
nand U5724 (N_5724,N_5109,N_5418);
nor U5725 (N_5725,N_5424,N_5024);
xor U5726 (N_5726,N_5397,N_5432);
and U5727 (N_5727,N_5065,N_5098);
xnor U5728 (N_5728,N_5047,N_5248);
nand U5729 (N_5729,N_5002,N_5381);
nand U5730 (N_5730,N_5014,N_5146);
xor U5731 (N_5731,N_5454,N_5294);
or U5732 (N_5732,N_5354,N_5056);
and U5733 (N_5733,N_5429,N_5210);
or U5734 (N_5734,N_5317,N_5102);
xor U5735 (N_5735,N_5408,N_5493);
or U5736 (N_5736,N_5382,N_5144);
and U5737 (N_5737,N_5434,N_5097);
xnor U5738 (N_5738,N_5227,N_5283);
nand U5739 (N_5739,N_5039,N_5236);
nor U5740 (N_5740,N_5440,N_5478);
xnor U5741 (N_5741,N_5347,N_5425);
nand U5742 (N_5742,N_5092,N_5278);
xor U5743 (N_5743,N_5445,N_5427);
nor U5744 (N_5744,N_5307,N_5241);
and U5745 (N_5745,N_5225,N_5297);
nand U5746 (N_5746,N_5326,N_5234);
or U5747 (N_5747,N_5188,N_5142);
and U5748 (N_5748,N_5488,N_5390);
or U5749 (N_5749,N_5128,N_5350);
or U5750 (N_5750,N_5195,N_5177);
xor U5751 (N_5751,N_5039,N_5174);
and U5752 (N_5752,N_5498,N_5008);
or U5753 (N_5753,N_5003,N_5129);
and U5754 (N_5754,N_5024,N_5020);
and U5755 (N_5755,N_5186,N_5023);
or U5756 (N_5756,N_5421,N_5023);
xor U5757 (N_5757,N_5448,N_5094);
nand U5758 (N_5758,N_5481,N_5200);
nor U5759 (N_5759,N_5253,N_5466);
nand U5760 (N_5760,N_5428,N_5396);
xnor U5761 (N_5761,N_5430,N_5006);
and U5762 (N_5762,N_5436,N_5347);
xnor U5763 (N_5763,N_5299,N_5055);
nor U5764 (N_5764,N_5139,N_5359);
xnor U5765 (N_5765,N_5466,N_5060);
nand U5766 (N_5766,N_5106,N_5430);
and U5767 (N_5767,N_5039,N_5485);
or U5768 (N_5768,N_5079,N_5025);
xnor U5769 (N_5769,N_5469,N_5139);
nor U5770 (N_5770,N_5300,N_5001);
or U5771 (N_5771,N_5403,N_5387);
and U5772 (N_5772,N_5000,N_5036);
and U5773 (N_5773,N_5188,N_5483);
xor U5774 (N_5774,N_5057,N_5380);
xor U5775 (N_5775,N_5466,N_5142);
nor U5776 (N_5776,N_5191,N_5463);
or U5777 (N_5777,N_5210,N_5482);
nand U5778 (N_5778,N_5085,N_5342);
nor U5779 (N_5779,N_5073,N_5129);
xnor U5780 (N_5780,N_5329,N_5356);
xnor U5781 (N_5781,N_5154,N_5232);
xnor U5782 (N_5782,N_5082,N_5400);
or U5783 (N_5783,N_5203,N_5028);
nor U5784 (N_5784,N_5128,N_5237);
or U5785 (N_5785,N_5490,N_5018);
or U5786 (N_5786,N_5053,N_5408);
xnor U5787 (N_5787,N_5030,N_5161);
nor U5788 (N_5788,N_5152,N_5366);
nand U5789 (N_5789,N_5144,N_5095);
nor U5790 (N_5790,N_5419,N_5477);
and U5791 (N_5791,N_5462,N_5187);
nand U5792 (N_5792,N_5498,N_5170);
and U5793 (N_5793,N_5067,N_5365);
and U5794 (N_5794,N_5158,N_5065);
xor U5795 (N_5795,N_5302,N_5460);
or U5796 (N_5796,N_5228,N_5465);
or U5797 (N_5797,N_5082,N_5351);
nand U5798 (N_5798,N_5141,N_5414);
and U5799 (N_5799,N_5429,N_5168);
and U5800 (N_5800,N_5113,N_5457);
or U5801 (N_5801,N_5437,N_5214);
nand U5802 (N_5802,N_5136,N_5236);
and U5803 (N_5803,N_5043,N_5179);
and U5804 (N_5804,N_5456,N_5293);
nor U5805 (N_5805,N_5488,N_5427);
and U5806 (N_5806,N_5072,N_5283);
nor U5807 (N_5807,N_5097,N_5225);
xnor U5808 (N_5808,N_5229,N_5289);
nand U5809 (N_5809,N_5401,N_5229);
xor U5810 (N_5810,N_5249,N_5024);
xor U5811 (N_5811,N_5215,N_5116);
nand U5812 (N_5812,N_5101,N_5082);
and U5813 (N_5813,N_5177,N_5031);
and U5814 (N_5814,N_5235,N_5283);
nor U5815 (N_5815,N_5445,N_5093);
nor U5816 (N_5816,N_5021,N_5427);
nor U5817 (N_5817,N_5266,N_5371);
nor U5818 (N_5818,N_5154,N_5110);
nor U5819 (N_5819,N_5125,N_5315);
and U5820 (N_5820,N_5117,N_5012);
or U5821 (N_5821,N_5270,N_5006);
nand U5822 (N_5822,N_5425,N_5000);
or U5823 (N_5823,N_5148,N_5314);
xor U5824 (N_5824,N_5128,N_5014);
nand U5825 (N_5825,N_5134,N_5037);
and U5826 (N_5826,N_5096,N_5350);
xor U5827 (N_5827,N_5448,N_5015);
xor U5828 (N_5828,N_5221,N_5077);
or U5829 (N_5829,N_5033,N_5431);
nand U5830 (N_5830,N_5294,N_5471);
nand U5831 (N_5831,N_5030,N_5048);
nor U5832 (N_5832,N_5039,N_5372);
nand U5833 (N_5833,N_5365,N_5373);
nand U5834 (N_5834,N_5150,N_5007);
and U5835 (N_5835,N_5048,N_5332);
xor U5836 (N_5836,N_5159,N_5474);
or U5837 (N_5837,N_5153,N_5454);
nor U5838 (N_5838,N_5082,N_5348);
and U5839 (N_5839,N_5428,N_5269);
nor U5840 (N_5840,N_5064,N_5039);
nor U5841 (N_5841,N_5114,N_5306);
xnor U5842 (N_5842,N_5199,N_5493);
nor U5843 (N_5843,N_5457,N_5355);
nand U5844 (N_5844,N_5331,N_5270);
or U5845 (N_5845,N_5214,N_5198);
nand U5846 (N_5846,N_5241,N_5230);
or U5847 (N_5847,N_5380,N_5282);
xor U5848 (N_5848,N_5073,N_5257);
xor U5849 (N_5849,N_5369,N_5455);
and U5850 (N_5850,N_5227,N_5198);
and U5851 (N_5851,N_5490,N_5123);
xnor U5852 (N_5852,N_5229,N_5165);
xnor U5853 (N_5853,N_5255,N_5073);
and U5854 (N_5854,N_5090,N_5278);
nor U5855 (N_5855,N_5294,N_5371);
or U5856 (N_5856,N_5377,N_5028);
and U5857 (N_5857,N_5350,N_5144);
xor U5858 (N_5858,N_5141,N_5361);
nor U5859 (N_5859,N_5200,N_5374);
nand U5860 (N_5860,N_5150,N_5298);
nor U5861 (N_5861,N_5321,N_5485);
xnor U5862 (N_5862,N_5443,N_5164);
xnor U5863 (N_5863,N_5109,N_5415);
nand U5864 (N_5864,N_5267,N_5414);
nand U5865 (N_5865,N_5063,N_5403);
or U5866 (N_5866,N_5126,N_5157);
and U5867 (N_5867,N_5372,N_5069);
nor U5868 (N_5868,N_5429,N_5294);
or U5869 (N_5869,N_5404,N_5367);
and U5870 (N_5870,N_5357,N_5369);
nand U5871 (N_5871,N_5283,N_5429);
nor U5872 (N_5872,N_5165,N_5313);
nor U5873 (N_5873,N_5007,N_5258);
xor U5874 (N_5874,N_5246,N_5142);
nand U5875 (N_5875,N_5482,N_5077);
nor U5876 (N_5876,N_5067,N_5478);
xnor U5877 (N_5877,N_5351,N_5046);
and U5878 (N_5878,N_5259,N_5156);
or U5879 (N_5879,N_5037,N_5277);
xor U5880 (N_5880,N_5050,N_5446);
xor U5881 (N_5881,N_5214,N_5193);
xor U5882 (N_5882,N_5319,N_5029);
nand U5883 (N_5883,N_5177,N_5485);
nand U5884 (N_5884,N_5177,N_5005);
xor U5885 (N_5885,N_5179,N_5398);
or U5886 (N_5886,N_5430,N_5287);
nor U5887 (N_5887,N_5027,N_5315);
xnor U5888 (N_5888,N_5135,N_5042);
nand U5889 (N_5889,N_5332,N_5306);
xnor U5890 (N_5890,N_5046,N_5035);
or U5891 (N_5891,N_5157,N_5379);
nand U5892 (N_5892,N_5050,N_5243);
nor U5893 (N_5893,N_5448,N_5006);
nand U5894 (N_5894,N_5093,N_5142);
or U5895 (N_5895,N_5343,N_5183);
nor U5896 (N_5896,N_5380,N_5284);
xnor U5897 (N_5897,N_5348,N_5298);
and U5898 (N_5898,N_5028,N_5366);
xnor U5899 (N_5899,N_5472,N_5268);
and U5900 (N_5900,N_5474,N_5332);
xor U5901 (N_5901,N_5424,N_5420);
or U5902 (N_5902,N_5166,N_5373);
or U5903 (N_5903,N_5365,N_5186);
nand U5904 (N_5904,N_5234,N_5095);
nand U5905 (N_5905,N_5085,N_5419);
or U5906 (N_5906,N_5225,N_5237);
xor U5907 (N_5907,N_5079,N_5147);
or U5908 (N_5908,N_5375,N_5030);
xnor U5909 (N_5909,N_5299,N_5103);
or U5910 (N_5910,N_5276,N_5311);
and U5911 (N_5911,N_5318,N_5145);
or U5912 (N_5912,N_5179,N_5468);
nand U5913 (N_5913,N_5409,N_5406);
or U5914 (N_5914,N_5190,N_5345);
nor U5915 (N_5915,N_5043,N_5018);
xor U5916 (N_5916,N_5080,N_5337);
nor U5917 (N_5917,N_5081,N_5211);
and U5918 (N_5918,N_5166,N_5160);
xor U5919 (N_5919,N_5318,N_5250);
nor U5920 (N_5920,N_5128,N_5090);
nor U5921 (N_5921,N_5491,N_5295);
and U5922 (N_5922,N_5087,N_5421);
nor U5923 (N_5923,N_5104,N_5458);
nor U5924 (N_5924,N_5231,N_5361);
xor U5925 (N_5925,N_5445,N_5213);
or U5926 (N_5926,N_5161,N_5122);
or U5927 (N_5927,N_5081,N_5470);
or U5928 (N_5928,N_5287,N_5265);
and U5929 (N_5929,N_5075,N_5372);
nor U5930 (N_5930,N_5324,N_5382);
and U5931 (N_5931,N_5211,N_5262);
nor U5932 (N_5932,N_5287,N_5234);
nand U5933 (N_5933,N_5356,N_5370);
or U5934 (N_5934,N_5018,N_5045);
nand U5935 (N_5935,N_5029,N_5307);
xor U5936 (N_5936,N_5037,N_5396);
xor U5937 (N_5937,N_5140,N_5084);
and U5938 (N_5938,N_5178,N_5255);
and U5939 (N_5939,N_5152,N_5398);
xnor U5940 (N_5940,N_5355,N_5109);
or U5941 (N_5941,N_5179,N_5452);
xnor U5942 (N_5942,N_5024,N_5367);
or U5943 (N_5943,N_5059,N_5319);
and U5944 (N_5944,N_5187,N_5454);
or U5945 (N_5945,N_5388,N_5315);
nand U5946 (N_5946,N_5082,N_5496);
nand U5947 (N_5947,N_5184,N_5228);
xnor U5948 (N_5948,N_5265,N_5338);
or U5949 (N_5949,N_5149,N_5494);
nor U5950 (N_5950,N_5144,N_5449);
xnor U5951 (N_5951,N_5406,N_5326);
or U5952 (N_5952,N_5249,N_5316);
xor U5953 (N_5953,N_5085,N_5471);
and U5954 (N_5954,N_5128,N_5137);
xor U5955 (N_5955,N_5412,N_5469);
and U5956 (N_5956,N_5196,N_5466);
nand U5957 (N_5957,N_5166,N_5209);
or U5958 (N_5958,N_5433,N_5042);
xor U5959 (N_5959,N_5380,N_5242);
xnor U5960 (N_5960,N_5111,N_5173);
xnor U5961 (N_5961,N_5199,N_5478);
nand U5962 (N_5962,N_5186,N_5024);
or U5963 (N_5963,N_5029,N_5449);
or U5964 (N_5964,N_5134,N_5458);
or U5965 (N_5965,N_5237,N_5449);
nand U5966 (N_5966,N_5034,N_5262);
nor U5967 (N_5967,N_5282,N_5123);
nor U5968 (N_5968,N_5214,N_5293);
or U5969 (N_5969,N_5127,N_5402);
or U5970 (N_5970,N_5074,N_5296);
nand U5971 (N_5971,N_5315,N_5142);
nand U5972 (N_5972,N_5481,N_5091);
or U5973 (N_5973,N_5463,N_5049);
nor U5974 (N_5974,N_5060,N_5340);
nor U5975 (N_5975,N_5495,N_5258);
or U5976 (N_5976,N_5109,N_5177);
and U5977 (N_5977,N_5396,N_5097);
nand U5978 (N_5978,N_5000,N_5214);
nand U5979 (N_5979,N_5296,N_5190);
and U5980 (N_5980,N_5074,N_5336);
or U5981 (N_5981,N_5201,N_5105);
nand U5982 (N_5982,N_5434,N_5030);
nand U5983 (N_5983,N_5269,N_5498);
and U5984 (N_5984,N_5438,N_5190);
nor U5985 (N_5985,N_5439,N_5270);
nor U5986 (N_5986,N_5036,N_5015);
and U5987 (N_5987,N_5368,N_5095);
xor U5988 (N_5988,N_5265,N_5384);
and U5989 (N_5989,N_5031,N_5339);
nor U5990 (N_5990,N_5042,N_5170);
nand U5991 (N_5991,N_5445,N_5129);
and U5992 (N_5992,N_5426,N_5041);
and U5993 (N_5993,N_5124,N_5015);
xnor U5994 (N_5994,N_5115,N_5174);
and U5995 (N_5995,N_5444,N_5280);
nor U5996 (N_5996,N_5095,N_5158);
nor U5997 (N_5997,N_5134,N_5046);
nand U5998 (N_5998,N_5245,N_5065);
and U5999 (N_5999,N_5323,N_5449);
nor U6000 (N_6000,N_5867,N_5586);
and U6001 (N_6001,N_5729,N_5687);
and U6002 (N_6002,N_5797,N_5569);
nor U6003 (N_6003,N_5741,N_5823);
nor U6004 (N_6004,N_5572,N_5834);
xnor U6005 (N_6005,N_5896,N_5664);
and U6006 (N_6006,N_5578,N_5519);
nor U6007 (N_6007,N_5606,N_5788);
or U6008 (N_6008,N_5699,N_5818);
or U6009 (N_6009,N_5610,N_5798);
and U6010 (N_6010,N_5608,N_5879);
nand U6011 (N_6011,N_5785,N_5645);
and U6012 (N_6012,N_5558,N_5705);
and U6013 (N_6013,N_5767,N_5667);
nor U6014 (N_6014,N_5912,N_5794);
and U6015 (N_6015,N_5778,N_5697);
nand U6016 (N_6016,N_5943,N_5702);
and U6017 (N_6017,N_5573,N_5542);
and U6018 (N_6018,N_5829,N_5890);
or U6019 (N_6019,N_5724,N_5791);
or U6020 (N_6020,N_5539,N_5700);
xnor U6021 (N_6021,N_5979,N_5977);
nand U6022 (N_6022,N_5605,N_5948);
xnor U6023 (N_6023,N_5596,N_5865);
xnor U6024 (N_6024,N_5760,N_5905);
xnor U6025 (N_6025,N_5955,N_5826);
xor U6026 (N_6026,N_5956,N_5528);
xor U6027 (N_6027,N_5627,N_5968);
or U6028 (N_6028,N_5692,N_5560);
nand U6029 (N_6029,N_5711,N_5551);
or U6030 (N_6030,N_5727,N_5655);
and U6031 (N_6031,N_5874,N_5999);
nor U6032 (N_6032,N_5568,N_5515);
xor U6033 (N_6033,N_5684,N_5671);
and U6034 (N_6034,N_5967,N_5775);
and U6035 (N_6035,N_5747,N_5925);
and U6036 (N_6036,N_5696,N_5830);
nand U6037 (N_6037,N_5628,N_5982);
xor U6038 (N_6038,N_5839,N_5926);
or U6039 (N_6039,N_5854,N_5712);
nor U6040 (N_6040,N_5765,N_5891);
and U6041 (N_6041,N_5786,N_5562);
nand U6042 (N_6042,N_5672,N_5929);
or U6043 (N_6043,N_5603,N_5601);
nand U6044 (N_6044,N_5810,N_5595);
and U6045 (N_6045,N_5587,N_5592);
xnor U6046 (N_6046,N_5793,N_5716);
and U6047 (N_6047,N_5679,N_5766);
or U6048 (N_6048,N_5589,N_5670);
nand U6049 (N_6049,N_5548,N_5907);
xnor U6050 (N_6050,N_5772,N_5517);
or U6051 (N_6051,N_5880,N_5876);
and U6052 (N_6052,N_5915,N_5647);
nand U6053 (N_6053,N_5535,N_5631);
nand U6054 (N_6054,N_5918,N_5644);
xnor U6055 (N_6055,N_5878,N_5707);
and U6056 (N_6056,N_5846,N_5753);
and U6057 (N_6057,N_5782,N_5506);
nand U6058 (N_6058,N_5933,N_5504);
nand U6059 (N_6059,N_5825,N_5739);
and U6060 (N_6060,N_5989,N_5502);
nand U6061 (N_6061,N_5768,N_5897);
nand U6062 (N_6062,N_5734,N_5582);
nor U6063 (N_6063,N_5527,N_5799);
xnor U6064 (N_6064,N_5969,N_5660);
or U6065 (N_6065,N_5930,N_5756);
nor U6066 (N_6066,N_5708,N_5629);
nor U6067 (N_6067,N_5526,N_5927);
xnor U6068 (N_6068,N_5632,N_5530);
nor U6069 (N_6069,N_5850,N_5722);
nand U6070 (N_6070,N_5698,N_5646);
and U6071 (N_6071,N_5590,N_5959);
and U6072 (N_6072,N_5966,N_5514);
xor U6073 (N_6073,N_5892,N_5773);
or U6074 (N_6074,N_5614,N_5621);
or U6075 (N_6075,N_5884,N_5990);
nor U6076 (N_6076,N_5972,N_5923);
xnor U6077 (N_6077,N_5599,N_5790);
and U6078 (N_6078,N_5809,N_5703);
and U6079 (N_6079,N_5963,N_5721);
xnor U6080 (N_6080,N_5777,N_5507);
or U6081 (N_6081,N_5988,N_5758);
nand U6082 (N_6082,N_5849,N_5748);
xnor U6083 (N_6083,N_5900,N_5857);
and U6084 (N_6084,N_5730,N_5998);
nand U6085 (N_6085,N_5709,N_5640);
or U6086 (N_6086,N_5661,N_5508);
or U6087 (N_6087,N_5691,N_5561);
or U6088 (N_6088,N_5870,N_5577);
and U6089 (N_6089,N_5780,N_5863);
xor U6090 (N_6090,N_5885,N_5565);
nand U6091 (N_6091,N_5913,N_5648);
nor U6092 (N_6092,N_5754,N_5733);
and U6093 (N_6093,N_5581,N_5649);
nand U6094 (N_6094,N_5804,N_5835);
xnor U6095 (N_6095,N_5750,N_5550);
and U6096 (N_6096,N_5624,N_5801);
nand U6097 (N_6097,N_5690,N_5841);
nand U6098 (N_6098,N_5936,N_5620);
nor U6099 (N_6099,N_5570,N_5940);
nor U6100 (N_6100,N_5718,N_5685);
nor U6101 (N_6101,N_5832,N_5513);
and U6102 (N_6102,N_5787,N_5749);
nor U6103 (N_6103,N_5735,N_5752);
nor U6104 (N_6104,N_5639,N_5942);
xnor U6105 (N_6105,N_5531,N_5657);
xnor U6106 (N_6106,N_5806,N_5673);
or U6107 (N_6107,N_5976,N_5680);
xor U6108 (N_6108,N_5899,N_5505);
nand U6109 (N_6109,N_5662,N_5833);
xnor U6110 (N_6110,N_5824,N_5789);
xnor U6111 (N_6111,N_5686,N_5813);
xnor U6112 (N_6112,N_5992,N_5537);
nor U6113 (N_6113,N_5638,N_5622);
nor U6114 (N_6114,N_5553,N_5529);
nand U6115 (N_6115,N_5975,N_5591);
or U6116 (N_6116,N_5625,N_5973);
nor U6117 (N_6117,N_5952,N_5802);
xor U6118 (N_6118,N_5575,N_5909);
nand U6119 (N_6119,N_5889,N_5873);
xor U6120 (N_6120,N_5808,N_5994);
nor U6121 (N_6121,N_5944,N_5883);
or U6122 (N_6122,N_5745,N_5946);
nand U6123 (N_6123,N_5731,N_5904);
or U6124 (N_6124,N_5866,N_5842);
xor U6125 (N_6125,N_5524,N_5509);
nand U6126 (N_6126,N_5759,N_5616);
xnor U6127 (N_6127,N_5755,N_5911);
nand U6128 (N_6128,N_5997,N_5888);
nand U6129 (N_6129,N_5953,N_5853);
nor U6130 (N_6130,N_5985,N_5633);
or U6131 (N_6131,N_5996,N_5770);
and U6132 (N_6132,N_5961,N_5983);
nand U6133 (N_6133,N_5774,N_5844);
or U6134 (N_6134,N_5934,N_5795);
nand U6135 (N_6135,N_5970,N_5688);
nand U6136 (N_6136,N_5919,N_5761);
xnor U6137 (N_6137,N_5917,N_5643);
and U6138 (N_6138,N_5964,N_5831);
or U6139 (N_6139,N_5984,N_5860);
or U6140 (N_6140,N_5500,N_5594);
and U6141 (N_6141,N_5869,N_5555);
nand U6142 (N_6142,N_5609,N_5847);
nand U6143 (N_6143,N_5630,N_5965);
and U6144 (N_6144,N_5838,N_5675);
or U6145 (N_6145,N_5652,N_5681);
and U6146 (N_6146,N_5819,N_5937);
xnor U6147 (N_6147,N_5674,N_5738);
or U6148 (N_6148,N_5861,N_5552);
and U6149 (N_6149,N_5534,N_5784);
nor U6150 (N_6150,N_5613,N_5597);
nand U6151 (N_6151,N_5820,N_5931);
and U6152 (N_6152,N_5836,N_5993);
nor U6153 (N_6153,N_5541,N_5903);
and U6154 (N_6154,N_5611,N_5837);
xor U6155 (N_6155,N_5776,N_5714);
xnor U6156 (N_6156,N_5864,N_5945);
nor U6157 (N_6157,N_5805,N_5882);
xnor U6158 (N_6158,N_5615,N_5579);
and U6159 (N_6159,N_5618,N_5957);
nand U6160 (N_6160,N_5843,N_5779);
nand U6161 (N_6161,N_5726,N_5576);
and U6162 (N_6162,N_5821,N_5580);
xor U6163 (N_6163,N_5949,N_5512);
or U6164 (N_6164,N_5991,N_5901);
xnor U6165 (N_6165,N_5704,N_5851);
nand U6166 (N_6166,N_5962,N_5895);
nor U6167 (N_6167,N_5523,N_5852);
and U6168 (N_6168,N_5746,N_5653);
xnor U6169 (N_6169,N_5763,N_5725);
and U6170 (N_6170,N_5737,N_5668);
xor U6171 (N_6171,N_5563,N_5859);
and U6172 (N_6172,N_5736,N_5938);
nor U6173 (N_6173,N_5566,N_5939);
and U6174 (N_6174,N_5769,N_5980);
nand U6175 (N_6175,N_5886,N_5981);
nor U6176 (N_6176,N_5812,N_5567);
nor U6177 (N_6177,N_5525,N_5619);
nor U6178 (N_6178,N_5532,N_5855);
and U6179 (N_6179,N_5845,N_5574);
or U6180 (N_6180,N_5792,N_5920);
or U6181 (N_6181,N_5593,N_5706);
and U6182 (N_6182,N_5862,N_5693);
nand U6183 (N_6183,N_5585,N_5715);
nor U6184 (N_6184,N_5583,N_5695);
nand U6185 (N_6185,N_5800,N_5807);
and U6186 (N_6186,N_5742,N_5908);
or U6187 (N_6187,N_5954,N_5713);
or U6188 (N_6188,N_5636,N_5612);
nor U6189 (N_6189,N_5602,N_5871);
xnor U6190 (N_6190,N_5543,N_5683);
nand U6191 (N_6191,N_5922,N_5719);
xnor U6192 (N_6192,N_5520,N_5656);
nand U6193 (N_6193,N_5554,N_5564);
nand U6194 (N_6194,N_5898,N_5947);
xnor U6195 (N_6195,N_5971,N_5893);
and U6196 (N_6196,N_5941,N_5856);
or U6197 (N_6197,N_5663,N_5764);
nor U6198 (N_6198,N_5701,N_5666);
and U6199 (N_6199,N_5635,N_5815);
nand U6200 (N_6200,N_5522,N_5626);
and U6201 (N_6201,N_5651,N_5676);
and U6202 (N_6202,N_5974,N_5511);
and U6203 (N_6203,N_5694,N_5678);
nor U6204 (N_6204,N_5516,N_5559);
nor U6205 (N_6205,N_5728,N_5538);
nand U6206 (N_6206,N_5814,N_5545);
and U6207 (N_6207,N_5783,N_5995);
nor U6208 (N_6208,N_5598,N_5877);
nand U6209 (N_6209,N_5669,N_5811);
xnor U6210 (N_6210,N_5924,N_5935);
and U6211 (N_6211,N_5536,N_5617);
nand U6212 (N_6212,N_5960,N_5875);
and U6213 (N_6213,N_5796,N_5677);
or U6214 (N_6214,N_5958,N_5501);
nor U6215 (N_6215,N_5910,N_5637);
nor U6216 (N_6216,N_5906,N_5518);
and U6217 (N_6217,N_5744,N_5928);
nand U6218 (N_6218,N_5723,N_5510);
nor U6219 (N_6219,N_5521,N_5503);
and U6220 (N_6220,N_5932,N_5547);
nor U6221 (N_6221,N_5827,N_5914);
nand U6222 (N_6222,N_5549,N_5887);
xor U6223 (N_6223,N_5781,N_5740);
nor U6224 (N_6224,N_5816,N_5751);
xnor U6225 (N_6225,N_5916,N_5604);
nor U6226 (N_6226,N_5717,N_5817);
nand U6227 (N_6227,N_5642,N_5641);
and U6228 (N_6228,N_5600,N_5757);
nor U6229 (N_6229,N_5533,N_5828);
or U6230 (N_6230,N_5544,N_5732);
nand U6231 (N_6231,N_5654,N_5634);
or U6232 (N_6232,N_5822,N_5557);
nor U6233 (N_6233,N_5894,N_5868);
nand U6234 (N_6234,N_5540,N_5872);
nand U6235 (N_6235,N_5987,N_5921);
nand U6236 (N_6236,N_5978,N_5710);
nor U6237 (N_6237,N_5571,N_5720);
xor U6238 (N_6238,N_5682,N_5689);
nand U6239 (N_6239,N_5659,N_5762);
and U6240 (N_6240,N_5588,N_5623);
nor U6241 (N_6241,N_5650,N_5840);
or U6242 (N_6242,N_5902,N_5607);
xnor U6243 (N_6243,N_5584,N_5771);
nor U6244 (N_6244,N_5950,N_5858);
nand U6245 (N_6245,N_5986,N_5881);
nor U6246 (N_6246,N_5743,N_5803);
and U6247 (N_6247,N_5951,N_5658);
nand U6248 (N_6248,N_5546,N_5556);
and U6249 (N_6249,N_5848,N_5665);
or U6250 (N_6250,N_5524,N_5985);
and U6251 (N_6251,N_5900,N_5573);
xor U6252 (N_6252,N_5501,N_5667);
xor U6253 (N_6253,N_5826,N_5740);
xnor U6254 (N_6254,N_5917,N_5609);
and U6255 (N_6255,N_5960,N_5668);
nor U6256 (N_6256,N_5576,N_5958);
and U6257 (N_6257,N_5652,N_5640);
xor U6258 (N_6258,N_5637,N_5549);
and U6259 (N_6259,N_5645,N_5557);
nand U6260 (N_6260,N_5642,N_5761);
nor U6261 (N_6261,N_5611,N_5760);
or U6262 (N_6262,N_5518,N_5689);
xor U6263 (N_6263,N_5831,N_5862);
nor U6264 (N_6264,N_5932,N_5657);
nand U6265 (N_6265,N_5980,N_5931);
nand U6266 (N_6266,N_5785,N_5694);
or U6267 (N_6267,N_5551,N_5504);
nand U6268 (N_6268,N_5559,N_5673);
xor U6269 (N_6269,N_5761,N_5862);
nor U6270 (N_6270,N_5854,N_5578);
nand U6271 (N_6271,N_5749,N_5637);
nand U6272 (N_6272,N_5919,N_5768);
and U6273 (N_6273,N_5778,N_5571);
nor U6274 (N_6274,N_5516,N_5724);
nor U6275 (N_6275,N_5885,N_5869);
and U6276 (N_6276,N_5695,N_5500);
nor U6277 (N_6277,N_5554,N_5504);
xnor U6278 (N_6278,N_5656,N_5990);
nand U6279 (N_6279,N_5807,N_5810);
nor U6280 (N_6280,N_5834,N_5620);
nand U6281 (N_6281,N_5885,N_5744);
nor U6282 (N_6282,N_5767,N_5653);
xnor U6283 (N_6283,N_5579,N_5957);
and U6284 (N_6284,N_5592,N_5666);
and U6285 (N_6285,N_5844,N_5576);
nor U6286 (N_6286,N_5849,N_5752);
nand U6287 (N_6287,N_5895,N_5654);
xnor U6288 (N_6288,N_5776,N_5638);
or U6289 (N_6289,N_5815,N_5915);
and U6290 (N_6290,N_5854,N_5610);
nand U6291 (N_6291,N_5807,N_5910);
and U6292 (N_6292,N_5552,N_5701);
nand U6293 (N_6293,N_5594,N_5679);
and U6294 (N_6294,N_5585,N_5760);
or U6295 (N_6295,N_5893,N_5888);
xor U6296 (N_6296,N_5933,N_5539);
or U6297 (N_6297,N_5939,N_5519);
xnor U6298 (N_6298,N_5635,N_5924);
nor U6299 (N_6299,N_5978,N_5899);
xnor U6300 (N_6300,N_5618,N_5982);
or U6301 (N_6301,N_5930,N_5886);
or U6302 (N_6302,N_5998,N_5857);
and U6303 (N_6303,N_5703,N_5887);
nand U6304 (N_6304,N_5981,N_5946);
or U6305 (N_6305,N_5928,N_5717);
nor U6306 (N_6306,N_5722,N_5911);
xor U6307 (N_6307,N_5923,N_5623);
nor U6308 (N_6308,N_5700,N_5871);
and U6309 (N_6309,N_5722,N_5711);
or U6310 (N_6310,N_5865,N_5723);
nor U6311 (N_6311,N_5621,N_5580);
nand U6312 (N_6312,N_5701,N_5867);
nor U6313 (N_6313,N_5675,N_5804);
xor U6314 (N_6314,N_5728,N_5799);
and U6315 (N_6315,N_5623,N_5746);
or U6316 (N_6316,N_5597,N_5662);
nand U6317 (N_6317,N_5905,N_5823);
nor U6318 (N_6318,N_5618,N_5683);
nand U6319 (N_6319,N_5836,N_5524);
and U6320 (N_6320,N_5992,N_5726);
or U6321 (N_6321,N_5733,N_5724);
nor U6322 (N_6322,N_5614,N_5587);
xnor U6323 (N_6323,N_5593,N_5628);
nand U6324 (N_6324,N_5539,N_5890);
or U6325 (N_6325,N_5895,N_5921);
nand U6326 (N_6326,N_5901,N_5764);
xnor U6327 (N_6327,N_5545,N_5580);
nor U6328 (N_6328,N_5525,N_5652);
nor U6329 (N_6329,N_5571,N_5963);
and U6330 (N_6330,N_5907,N_5895);
nor U6331 (N_6331,N_5523,N_5940);
xnor U6332 (N_6332,N_5999,N_5648);
nand U6333 (N_6333,N_5957,N_5829);
nand U6334 (N_6334,N_5529,N_5717);
xnor U6335 (N_6335,N_5567,N_5906);
or U6336 (N_6336,N_5645,N_5940);
nand U6337 (N_6337,N_5902,N_5575);
and U6338 (N_6338,N_5736,N_5724);
or U6339 (N_6339,N_5728,N_5782);
nor U6340 (N_6340,N_5903,N_5939);
nor U6341 (N_6341,N_5722,N_5532);
or U6342 (N_6342,N_5964,N_5937);
nand U6343 (N_6343,N_5595,N_5837);
or U6344 (N_6344,N_5810,N_5667);
nor U6345 (N_6345,N_5881,N_5594);
xnor U6346 (N_6346,N_5732,N_5886);
and U6347 (N_6347,N_5954,N_5757);
nor U6348 (N_6348,N_5506,N_5635);
xor U6349 (N_6349,N_5860,N_5677);
and U6350 (N_6350,N_5758,N_5601);
and U6351 (N_6351,N_5572,N_5561);
xor U6352 (N_6352,N_5703,N_5764);
and U6353 (N_6353,N_5646,N_5602);
xnor U6354 (N_6354,N_5902,N_5623);
or U6355 (N_6355,N_5704,N_5934);
nand U6356 (N_6356,N_5689,N_5731);
xnor U6357 (N_6357,N_5511,N_5708);
or U6358 (N_6358,N_5729,N_5673);
nor U6359 (N_6359,N_5806,N_5810);
or U6360 (N_6360,N_5785,N_5566);
xor U6361 (N_6361,N_5504,N_5938);
nand U6362 (N_6362,N_5696,N_5513);
nand U6363 (N_6363,N_5608,N_5932);
nand U6364 (N_6364,N_5647,N_5774);
and U6365 (N_6365,N_5602,N_5917);
or U6366 (N_6366,N_5702,N_5866);
nor U6367 (N_6367,N_5766,N_5760);
nor U6368 (N_6368,N_5951,N_5711);
nand U6369 (N_6369,N_5520,N_5793);
and U6370 (N_6370,N_5992,N_5738);
xnor U6371 (N_6371,N_5745,N_5904);
nor U6372 (N_6372,N_5630,N_5779);
and U6373 (N_6373,N_5819,N_5973);
nor U6374 (N_6374,N_5689,N_5654);
xor U6375 (N_6375,N_5571,N_5916);
and U6376 (N_6376,N_5777,N_5927);
nand U6377 (N_6377,N_5994,N_5890);
xor U6378 (N_6378,N_5632,N_5590);
xnor U6379 (N_6379,N_5813,N_5661);
nand U6380 (N_6380,N_5873,N_5602);
nor U6381 (N_6381,N_5909,N_5994);
xnor U6382 (N_6382,N_5874,N_5636);
and U6383 (N_6383,N_5870,N_5731);
and U6384 (N_6384,N_5860,N_5558);
nand U6385 (N_6385,N_5746,N_5904);
and U6386 (N_6386,N_5670,N_5692);
or U6387 (N_6387,N_5802,N_5923);
or U6388 (N_6388,N_5980,N_5636);
xnor U6389 (N_6389,N_5504,N_5937);
nand U6390 (N_6390,N_5735,N_5996);
nand U6391 (N_6391,N_5739,N_5890);
xnor U6392 (N_6392,N_5955,N_5695);
or U6393 (N_6393,N_5702,N_5629);
xnor U6394 (N_6394,N_5785,N_5788);
xnor U6395 (N_6395,N_5711,N_5921);
xor U6396 (N_6396,N_5750,N_5583);
or U6397 (N_6397,N_5548,N_5924);
or U6398 (N_6398,N_5637,N_5500);
and U6399 (N_6399,N_5541,N_5618);
nand U6400 (N_6400,N_5551,N_5769);
and U6401 (N_6401,N_5737,N_5674);
or U6402 (N_6402,N_5991,N_5785);
nand U6403 (N_6403,N_5972,N_5862);
nand U6404 (N_6404,N_5643,N_5579);
or U6405 (N_6405,N_5718,N_5524);
nor U6406 (N_6406,N_5870,N_5530);
nand U6407 (N_6407,N_5904,N_5574);
or U6408 (N_6408,N_5925,N_5825);
and U6409 (N_6409,N_5974,N_5996);
xor U6410 (N_6410,N_5751,N_5747);
nand U6411 (N_6411,N_5669,N_5997);
nor U6412 (N_6412,N_5660,N_5822);
and U6413 (N_6413,N_5941,N_5925);
and U6414 (N_6414,N_5919,N_5784);
nand U6415 (N_6415,N_5856,N_5690);
xnor U6416 (N_6416,N_5909,N_5950);
xnor U6417 (N_6417,N_5942,N_5843);
nor U6418 (N_6418,N_5862,N_5665);
nor U6419 (N_6419,N_5946,N_5610);
nor U6420 (N_6420,N_5930,N_5616);
or U6421 (N_6421,N_5763,N_5591);
or U6422 (N_6422,N_5711,N_5545);
nand U6423 (N_6423,N_5992,N_5694);
nor U6424 (N_6424,N_5571,N_5739);
or U6425 (N_6425,N_5853,N_5883);
or U6426 (N_6426,N_5858,N_5642);
or U6427 (N_6427,N_5720,N_5958);
nand U6428 (N_6428,N_5785,N_5758);
xor U6429 (N_6429,N_5803,N_5980);
and U6430 (N_6430,N_5839,N_5907);
nand U6431 (N_6431,N_5950,N_5659);
nor U6432 (N_6432,N_5905,N_5606);
nand U6433 (N_6433,N_5629,N_5760);
nor U6434 (N_6434,N_5929,N_5822);
nor U6435 (N_6435,N_5568,N_5519);
and U6436 (N_6436,N_5642,N_5608);
xnor U6437 (N_6437,N_5603,N_5880);
and U6438 (N_6438,N_5738,N_5911);
nor U6439 (N_6439,N_5556,N_5889);
and U6440 (N_6440,N_5972,N_5728);
and U6441 (N_6441,N_5844,N_5838);
or U6442 (N_6442,N_5775,N_5640);
nor U6443 (N_6443,N_5778,N_5655);
xor U6444 (N_6444,N_5970,N_5920);
nand U6445 (N_6445,N_5725,N_5736);
nand U6446 (N_6446,N_5633,N_5574);
nand U6447 (N_6447,N_5528,N_5546);
xnor U6448 (N_6448,N_5639,N_5822);
nand U6449 (N_6449,N_5755,N_5645);
nand U6450 (N_6450,N_5665,N_5785);
or U6451 (N_6451,N_5949,N_5600);
xor U6452 (N_6452,N_5931,N_5793);
or U6453 (N_6453,N_5734,N_5592);
or U6454 (N_6454,N_5919,N_5970);
or U6455 (N_6455,N_5558,N_5986);
nand U6456 (N_6456,N_5738,N_5788);
xor U6457 (N_6457,N_5607,N_5892);
nor U6458 (N_6458,N_5623,N_5749);
nor U6459 (N_6459,N_5561,N_5542);
nor U6460 (N_6460,N_5978,N_5747);
xor U6461 (N_6461,N_5791,N_5526);
nand U6462 (N_6462,N_5621,N_5547);
and U6463 (N_6463,N_5955,N_5723);
nand U6464 (N_6464,N_5713,N_5571);
nor U6465 (N_6465,N_5958,N_5694);
nand U6466 (N_6466,N_5653,N_5696);
xor U6467 (N_6467,N_5646,N_5620);
nor U6468 (N_6468,N_5696,N_5688);
xor U6469 (N_6469,N_5969,N_5869);
and U6470 (N_6470,N_5735,N_5592);
nor U6471 (N_6471,N_5738,N_5832);
nor U6472 (N_6472,N_5763,N_5680);
nand U6473 (N_6473,N_5603,N_5876);
nor U6474 (N_6474,N_5965,N_5703);
or U6475 (N_6475,N_5676,N_5898);
nor U6476 (N_6476,N_5766,N_5682);
xor U6477 (N_6477,N_5759,N_5826);
and U6478 (N_6478,N_5679,N_5967);
xor U6479 (N_6479,N_5844,N_5877);
or U6480 (N_6480,N_5625,N_5868);
or U6481 (N_6481,N_5915,N_5909);
nand U6482 (N_6482,N_5896,N_5635);
nor U6483 (N_6483,N_5703,N_5945);
nand U6484 (N_6484,N_5610,N_5834);
and U6485 (N_6485,N_5760,N_5709);
or U6486 (N_6486,N_5835,N_5766);
or U6487 (N_6487,N_5771,N_5529);
and U6488 (N_6488,N_5833,N_5549);
xor U6489 (N_6489,N_5827,N_5854);
nand U6490 (N_6490,N_5588,N_5995);
nand U6491 (N_6491,N_5531,N_5688);
nor U6492 (N_6492,N_5816,N_5598);
nand U6493 (N_6493,N_5742,N_5629);
xnor U6494 (N_6494,N_5858,N_5806);
xnor U6495 (N_6495,N_5931,N_5746);
nor U6496 (N_6496,N_5962,N_5721);
nand U6497 (N_6497,N_5558,N_5993);
xnor U6498 (N_6498,N_5514,N_5591);
nand U6499 (N_6499,N_5797,N_5633);
xor U6500 (N_6500,N_6100,N_6411);
nor U6501 (N_6501,N_6143,N_6373);
or U6502 (N_6502,N_6159,N_6339);
xor U6503 (N_6503,N_6184,N_6241);
and U6504 (N_6504,N_6356,N_6341);
or U6505 (N_6505,N_6235,N_6165);
or U6506 (N_6506,N_6126,N_6125);
nor U6507 (N_6507,N_6409,N_6270);
nor U6508 (N_6508,N_6224,N_6458);
nand U6509 (N_6509,N_6368,N_6249);
or U6510 (N_6510,N_6042,N_6251);
nand U6511 (N_6511,N_6280,N_6268);
and U6512 (N_6512,N_6275,N_6226);
and U6513 (N_6513,N_6222,N_6155);
nand U6514 (N_6514,N_6490,N_6331);
xnor U6515 (N_6515,N_6117,N_6323);
nand U6516 (N_6516,N_6414,N_6383);
or U6517 (N_6517,N_6421,N_6273);
nor U6518 (N_6518,N_6336,N_6276);
and U6519 (N_6519,N_6021,N_6320);
and U6520 (N_6520,N_6462,N_6020);
nand U6521 (N_6521,N_6046,N_6427);
or U6522 (N_6522,N_6007,N_6037);
nand U6523 (N_6523,N_6419,N_6253);
and U6524 (N_6524,N_6113,N_6044);
xnor U6525 (N_6525,N_6154,N_6285);
or U6526 (N_6526,N_6358,N_6343);
nor U6527 (N_6527,N_6310,N_6340);
or U6528 (N_6528,N_6298,N_6203);
and U6529 (N_6529,N_6284,N_6095);
or U6530 (N_6530,N_6363,N_6434);
nand U6531 (N_6531,N_6277,N_6269);
nand U6532 (N_6532,N_6430,N_6231);
or U6533 (N_6533,N_6170,N_6319);
and U6534 (N_6534,N_6148,N_6166);
nand U6535 (N_6535,N_6473,N_6426);
xnor U6536 (N_6536,N_6064,N_6408);
nor U6537 (N_6537,N_6294,N_6288);
and U6538 (N_6538,N_6167,N_6147);
and U6539 (N_6539,N_6352,N_6066);
nand U6540 (N_6540,N_6296,N_6024);
or U6541 (N_6541,N_6232,N_6134);
and U6542 (N_6542,N_6479,N_6460);
or U6543 (N_6543,N_6333,N_6332);
nand U6544 (N_6544,N_6428,N_6257);
or U6545 (N_6545,N_6412,N_6264);
and U6546 (N_6546,N_6443,N_6461);
and U6547 (N_6547,N_6015,N_6201);
nor U6548 (N_6548,N_6348,N_6200);
xor U6549 (N_6549,N_6176,N_6417);
nand U6550 (N_6550,N_6039,N_6048);
nor U6551 (N_6551,N_6008,N_6199);
or U6552 (N_6552,N_6440,N_6403);
nand U6553 (N_6553,N_6110,N_6193);
nand U6554 (N_6554,N_6173,N_6013);
or U6555 (N_6555,N_6367,N_6136);
nor U6556 (N_6556,N_6171,N_6211);
or U6557 (N_6557,N_6228,N_6314);
nor U6558 (N_6558,N_6009,N_6289);
and U6559 (N_6559,N_6279,N_6056);
and U6560 (N_6560,N_6189,N_6150);
or U6561 (N_6561,N_6355,N_6149);
nor U6562 (N_6562,N_6471,N_6469);
or U6563 (N_6563,N_6478,N_6106);
nand U6564 (N_6564,N_6040,N_6192);
or U6565 (N_6565,N_6115,N_6220);
xnor U6566 (N_6566,N_6213,N_6243);
nor U6567 (N_6567,N_6422,N_6001);
or U6568 (N_6568,N_6286,N_6190);
nor U6569 (N_6569,N_6030,N_6255);
and U6570 (N_6570,N_6000,N_6181);
nor U6571 (N_6571,N_6011,N_6062);
nor U6572 (N_6572,N_6396,N_6194);
or U6573 (N_6573,N_6087,N_6272);
and U6574 (N_6574,N_6137,N_6499);
xor U6575 (N_6575,N_6395,N_6182);
or U6576 (N_6576,N_6006,N_6082);
nand U6577 (N_6577,N_6245,N_6472);
xor U6578 (N_6578,N_6326,N_6078);
nor U6579 (N_6579,N_6389,N_6405);
nand U6580 (N_6580,N_6233,N_6315);
nor U6581 (N_6581,N_6236,N_6488);
nor U6582 (N_6582,N_6088,N_6342);
and U6583 (N_6583,N_6256,N_6386);
or U6584 (N_6584,N_6299,N_6109);
or U6585 (N_6585,N_6244,N_6129);
or U6586 (N_6586,N_6209,N_6071);
and U6587 (N_6587,N_6198,N_6357);
and U6588 (N_6588,N_6442,N_6085);
or U6589 (N_6589,N_6486,N_6450);
xor U6590 (N_6590,N_6305,N_6123);
nor U6591 (N_6591,N_6187,N_6105);
xor U6592 (N_6592,N_6210,N_6097);
and U6593 (N_6593,N_6350,N_6025);
nor U6594 (N_6594,N_6494,N_6438);
nor U6595 (N_6595,N_6262,N_6445);
or U6596 (N_6596,N_6041,N_6379);
xnor U6597 (N_6597,N_6197,N_6308);
or U6598 (N_6598,N_6242,N_6174);
nor U6599 (N_6599,N_6391,N_6346);
nand U6600 (N_6600,N_6101,N_6112);
xnor U6601 (N_6601,N_6365,N_6334);
and U6602 (N_6602,N_6207,N_6160);
and U6603 (N_6603,N_6072,N_6073);
and U6604 (N_6604,N_6397,N_6327);
nor U6605 (N_6605,N_6047,N_6292);
nand U6606 (N_6606,N_6309,N_6484);
and U6607 (N_6607,N_6477,N_6359);
nor U6608 (N_6608,N_6075,N_6446);
nor U6609 (N_6609,N_6274,N_6407);
nand U6610 (N_6610,N_6475,N_6023);
nand U6611 (N_6611,N_6212,N_6059);
xor U6612 (N_6612,N_6079,N_6108);
nor U6613 (N_6613,N_6423,N_6138);
nor U6614 (N_6614,N_6033,N_6385);
nand U6615 (N_6615,N_6074,N_6283);
nand U6616 (N_6616,N_6361,N_6467);
or U6617 (N_6617,N_6287,N_6083);
nor U6618 (N_6618,N_6103,N_6002);
and U6619 (N_6619,N_6317,N_6145);
or U6620 (N_6620,N_6351,N_6151);
and U6621 (N_6621,N_6297,N_6218);
nor U6622 (N_6622,N_6400,N_6436);
xor U6623 (N_6623,N_6324,N_6225);
nand U6624 (N_6624,N_6238,N_6043);
nor U6625 (N_6625,N_6202,N_6457);
xnor U6626 (N_6626,N_6240,N_6335);
xor U6627 (N_6627,N_6448,N_6399);
or U6628 (N_6628,N_6487,N_6433);
nor U6629 (N_6629,N_6254,N_6261);
nand U6630 (N_6630,N_6168,N_6402);
nand U6631 (N_6631,N_6077,N_6474);
or U6632 (N_6632,N_6019,N_6360);
xor U6633 (N_6633,N_6153,N_6258);
and U6634 (N_6634,N_6466,N_6052);
nor U6635 (N_6635,N_6259,N_6034);
and U6636 (N_6636,N_6304,N_6293);
or U6637 (N_6637,N_6420,N_6035);
xnor U6638 (N_6638,N_6012,N_6191);
xor U6639 (N_6639,N_6177,N_6322);
nor U6640 (N_6640,N_6164,N_6321);
or U6641 (N_6641,N_6424,N_6004);
xnor U6642 (N_6642,N_6169,N_6162);
xor U6643 (N_6643,N_6435,N_6265);
and U6644 (N_6644,N_6133,N_6328);
or U6645 (N_6645,N_6057,N_6493);
or U6646 (N_6646,N_6470,N_6084);
or U6647 (N_6647,N_6416,N_6406);
or U6648 (N_6648,N_6055,N_6489);
xor U6649 (N_6649,N_6371,N_6152);
nand U6650 (N_6650,N_6377,N_6463);
nand U6651 (N_6651,N_6104,N_6076);
and U6652 (N_6652,N_6263,N_6054);
and U6653 (N_6653,N_6067,N_6390);
nand U6654 (N_6654,N_6441,N_6131);
nor U6655 (N_6655,N_6130,N_6161);
nand U6656 (N_6656,N_6338,N_6080);
nand U6657 (N_6657,N_6157,N_6345);
nand U6658 (N_6658,N_6185,N_6344);
nor U6659 (N_6659,N_6158,N_6318);
nor U6660 (N_6660,N_6480,N_6204);
and U6661 (N_6661,N_6329,N_6455);
nor U6662 (N_6662,N_6290,N_6482);
or U6663 (N_6663,N_6398,N_6234);
xor U6664 (N_6664,N_6163,N_6432);
and U6665 (N_6665,N_6229,N_6447);
or U6666 (N_6666,N_6401,N_6239);
nand U6667 (N_6667,N_6032,N_6219);
nand U6668 (N_6668,N_6495,N_6127);
xor U6669 (N_6669,N_6491,N_6038);
and U6670 (N_6670,N_6096,N_6387);
nor U6671 (N_6671,N_6028,N_6465);
xnor U6672 (N_6672,N_6139,N_6050);
nand U6673 (N_6673,N_6223,N_6121);
nor U6674 (N_6674,N_6388,N_6092);
and U6675 (N_6675,N_6295,N_6330);
xor U6676 (N_6676,N_6300,N_6017);
and U6677 (N_6677,N_6156,N_6459);
nor U6678 (N_6678,N_6188,N_6058);
xor U6679 (N_6679,N_6124,N_6354);
xnor U6680 (N_6680,N_6206,N_6370);
nand U6681 (N_6681,N_6311,N_6146);
nor U6682 (N_6682,N_6049,N_6347);
nor U6683 (N_6683,N_6195,N_6237);
nand U6684 (N_6684,N_6378,N_6413);
xor U6685 (N_6685,N_6483,N_6302);
and U6686 (N_6686,N_6005,N_6141);
nor U6687 (N_6687,N_6144,N_6393);
nor U6688 (N_6688,N_6102,N_6392);
and U6689 (N_6689,N_6364,N_6306);
nor U6690 (N_6690,N_6282,N_6183);
and U6691 (N_6691,N_6464,N_6230);
and U6692 (N_6692,N_6116,N_6031);
and U6693 (N_6693,N_6090,N_6415);
and U6694 (N_6694,N_6452,N_6120);
nor U6695 (N_6695,N_6429,N_6369);
and U6696 (N_6696,N_6376,N_6142);
or U6697 (N_6697,N_6266,N_6439);
or U6698 (N_6698,N_6215,N_6221);
nand U6699 (N_6699,N_6036,N_6481);
xor U6700 (N_6700,N_6068,N_6312);
xnor U6701 (N_6701,N_6119,N_6260);
nor U6702 (N_6702,N_6451,N_6026);
and U6703 (N_6703,N_6325,N_6065);
xnor U6704 (N_6704,N_6349,N_6404);
xor U6705 (N_6705,N_6196,N_6093);
nand U6706 (N_6706,N_6111,N_6476);
or U6707 (N_6707,N_6453,N_6029);
nor U6708 (N_6708,N_6316,N_6069);
and U6709 (N_6709,N_6375,N_6186);
or U6710 (N_6710,N_6362,N_6063);
and U6711 (N_6711,N_6410,N_6018);
nor U6712 (N_6712,N_6172,N_6122);
nor U6713 (N_6713,N_6394,N_6492);
nand U6714 (N_6714,N_6061,N_6227);
nor U6715 (N_6715,N_6291,N_6010);
and U6716 (N_6716,N_6246,N_6281);
and U6717 (N_6717,N_6303,N_6384);
nor U6718 (N_6718,N_6248,N_6070);
xnor U6719 (N_6719,N_6250,N_6114);
nor U6720 (N_6720,N_6178,N_6278);
or U6721 (N_6721,N_6016,N_6485);
nand U6722 (N_6722,N_6252,N_6498);
nand U6723 (N_6723,N_6179,N_6267);
nor U6724 (N_6724,N_6060,N_6214);
nand U6725 (N_6725,N_6132,N_6045);
or U6726 (N_6726,N_6468,N_6027);
xnor U6727 (N_6727,N_6217,N_6098);
or U6728 (N_6728,N_6128,N_6208);
xor U6729 (N_6729,N_6081,N_6135);
nand U6730 (N_6730,N_6118,N_6051);
nand U6731 (N_6731,N_6456,N_6337);
nand U6732 (N_6732,N_6089,N_6372);
and U6733 (N_6733,N_6366,N_6107);
xnor U6734 (N_6734,N_6301,N_6091);
or U6735 (N_6735,N_6425,N_6003);
xnor U6736 (N_6736,N_6180,N_6271);
and U6737 (N_6737,N_6094,N_6497);
nor U6738 (N_6738,N_6381,N_6449);
xnor U6739 (N_6739,N_6307,N_6014);
nor U6740 (N_6740,N_6418,N_6437);
nand U6741 (N_6741,N_6382,N_6216);
or U6742 (N_6742,N_6022,N_6313);
nand U6743 (N_6743,N_6140,N_6496);
or U6744 (N_6744,N_6086,N_6053);
nor U6745 (N_6745,N_6431,N_6444);
or U6746 (N_6746,N_6099,N_6454);
nor U6747 (N_6747,N_6247,N_6175);
nor U6748 (N_6748,N_6353,N_6380);
nor U6749 (N_6749,N_6205,N_6374);
and U6750 (N_6750,N_6494,N_6120);
nand U6751 (N_6751,N_6102,N_6357);
and U6752 (N_6752,N_6043,N_6445);
xor U6753 (N_6753,N_6240,N_6205);
nand U6754 (N_6754,N_6357,N_6320);
nor U6755 (N_6755,N_6341,N_6209);
and U6756 (N_6756,N_6062,N_6146);
or U6757 (N_6757,N_6247,N_6231);
nand U6758 (N_6758,N_6156,N_6403);
and U6759 (N_6759,N_6017,N_6175);
or U6760 (N_6760,N_6285,N_6298);
xnor U6761 (N_6761,N_6499,N_6041);
nor U6762 (N_6762,N_6201,N_6164);
and U6763 (N_6763,N_6201,N_6170);
nand U6764 (N_6764,N_6186,N_6208);
or U6765 (N_6765,N_6074,N_6148);
and U6766 (N_6766,N_6296,N_6318);
and U6767 (N_6767,N_6032,N_6156);
nand U6768 (N_6768,N_6439,N_6453);
nand U6769 (N_6769,N_6060,N_6485);
or U6770 (N_6770,N_6311,N_6233);
and U6771 (N_6771,N_6360,N_6207);
and U6772 (N_6772,N_6384,N_6301);
xor U6773 (N_6773,N_6239,N_6461);
and U6774 (N_6774,N_6404,N_6147);
xor U6775 (N_6775,N_6157,N_6232);
xnor U6776 (N_6776,N_6211,N_6196);
nand U6777 (N_6777,N_6164,N_6404);
and U6778 (N_6778,N_6349,N_6156);
nand U6779 (N_6779,N_6215,N_6365);
and U6780 (N_6780,N_6126,N_6438);
xor U6781 (N_6781,N_6045,N_6118);
nand U6782 (N_6782,N_6079,N_6008);
nor U6783 (N_6783,N_6415,N_6330);
nand U6784 (N_6784,N_6133,N_6052);
or U6785 (N_6785,N_6195,N_6022);
nor U6786 (N_6786,N_6221,N_6444);
nor U6787 (N_6787,N_6328,N_6487);
nor U6788 (N_6788,N_6285,N_6225);
nand U6789 (N_6789,N_6000,N_6289);
or U6790 (N_6790,N_6234,N_6211);
xor U6791 (N_6791,N_6245,N_6295);
xnor U6792 (N_6792,N_6132,N_6214);
or U6793 (N_6793,N_6339,N_6239);
or U6794 (N_6794,N_6322,N_6393);
nand U6795 (N_6795,N_6186,N_6393);
nor U6796 (N_6796,N_6241,N_6273);
and U6797 (N_6797,N_6311,N_6230);
nand U6798 (N_6798,N_6167,N_6239);
xor U6799 (N_6799,N_6183,N_6015);
nand U6800 (N_6800,N_6374,N_6116);
xor U6801 (N_6801,N_6089,N_6155);
or U6802 (N_6802,N_6190,N_6442);
nor U6803 (N_6803,N_6466,N_6338);
xnor U6804 (N_6804,N_6171,N_6227);
xnor U6805 (N_6805,N_6297,N_6446);
nor U6806 (N_6806,N_6063,N_6100);
or U6807 (N_6807,N_6040,N_6132);
nor U6808 (N_6808,N_6428,N_6446);
or U6809 (N_6809,N_6386,N_6321);
nor U6810 (N_6810,N_6175,N_6457);
and U6811 (N_6811,N_6041,N_6151);
nor U6812 (N_6812,N_6444,N_6142);
xor U6813 (N_6813,N_6407,N_6002);
nor U6814 (N_6814,N_6176,N_6299);
and U6815 (N_6815,N_6103,N_6268);
or U6816 (N_6816,N_6436,N_6339);
nor U6817 (N_6817,N_6074,N_6140);
and U6818 (N_6818,N_6334,N_6061);
nand U6819 (N_6819,N_6355,N_6210);
nand U6820 (N_6820,N_6244,N_6374);
nand U6821 (N_6821,N_6204,N_6341);
xor U6822 (N_6822,N_6356,N_6463);
nor U6823 (N_6823,N_6144,N_6436);
xor U6824 (N_6824,N_6052,N_6039);
nand U6825 (N_6825,N_6050,N_6378);
xnor U6826 (N_6826,N_6167,N_6150);
or U6827 (N_6827,N_6258,N_6099);
nand U6828 (N_6828,N_6212,N_6441);
nor U6829 (N_6829,N_6233,N_6045);
or U6830 (N_6830,N_6154,N_6483);
xnor U6831 (N_6831,N_6145,N_6394);
or U6832 (N_6832,N_6116,N_6383);
or U6833 (N_6833,N_6000,N_6034);
nand U6834 (N_6834,N_6481,N_6237);
or U6835 (N_6835,N_6006,N_6190);
and U6836 (N_6836,N_6221,N_6487);
xnor U6837 (N_6837,N_6161,N_6221);
and U6838 (N_6838,N_6083,N_6043);
xnor U6839 (N_6839,N_6035,N_6468);
and U6840 (N_6840,N_6494,N_6144);
nor U6841 (N_6841,N_6416,N_6227);
and U6842 (N_6842,N_6132,N_6320);
nand U6843 (N_6843,N_6258,N_6366);
and U6844 (N_6844,N_6037,N_6267);
and U6845 (N_6845,N_6348,N_6434);
or U6846 (N_6846,N_6136,N_6371);
xnor U6847 (N_6847,N_6037,N_6134);
or U6848 (N_6848,N_6016,N_6185);
xor U6849 (N_6849,N_6186,N_6081);
nor U6850 (N_6850,N_6268,N_6236);
nand U6851 (N_6851,N_6220,N_6174);
nor U6852 (N_6852,N_6362,N_6192);
or U6853 (N_6853,N_6366,N_6103);
and U6854 (N_6854,N_6332,N_6326);
xnor U6855 (N_6855,N_6260,N_6107);
and U6856 (N_6856,N_6043,N_6373);
xor U6857 (N_6857,N_6164,N_6053);
xnor U6858 (N_6858,N_6093,N_6137);
or U6859 (N_6859,N_6499,N_6055);
or U6860 (N_6860,N_6086,N_6407);
xnor U6861 (N_6861,N_6043,N_6150);
or U6862 (N_6862,N_6010,N_6278);
or U6863 (N_6863,N_6432,N_6344);
and U6864 (N_6864,N_6062,N_6387);
xor U6865 (N_6865,N_6004,N_6320);
xor U6866 (N_6866,N_6459,N_6191);
xnor U6867 (N_6867,N_6077,N_6498);
and U6868 (N_6868,N_6132,N_6270);
and U6869 (N_6869,N_6001,N_6112);
and U6870 (N_6870,N_6366,N_6244);
and U6871 (N_6871,N_6027,N_6068);
or U6872 (N_6872,N_6068,N_6017);
xnor U6873 (N_6873,N_6031,N_6010);
nor U6874 (N_6874,N_6004,N_6347);
nand U6875 (N_6875,N_6149,N_6078);
nor U6876 (N_6876,N_6141,N_6343);
nor U6877 (N_6877,N_6111,N_6107);
xnor U6878 (N_6878,N_6392,N_6069);
xnor U6879 (N_6879,N_6419,N_6119);
nand U6880 (N_6880,N_6470,N_6198);
xnor U6881 (N_6881,N_6072,N_6457);
nor U6882 (N_6882,N_6332,N_6122);
xor U6883 (N_6883,N_6400,N_6185);
nand U6884 (N_6884,N_6241,N_6461);
and U6885 (N_6885,N_6208,N_6184);
xnor U6886 (N_6886,N_6333,N_6062);
or U6887 (N_6887,N_6260,N_6393);
or U6888 (N_6888,N_6440,N_6406);
xnor U6889 (N_6889,N_6003,N_6027);
nor U6890 (N_6890,N_6424,N_6405);
or U6891 (N_6891,N_6216,N_6344);
or U6892 (N_6892,N_6382,N_6320);
xnor U6893 (N_6893,N_6222,N_6230);
nand U6894 (N_6894,N_6091,N_6259);
xnor U6895 (N_6895,N_6053,N_6315);
nor U6896 (N_6896,N_6080,N_6178);
or U6897 (N_6897,N_6256,N_6387);
nor U6898 (N_6898,N_6117,N_6341);
xnor U6899 (N_6899,N_6324,N_6336);
nor U6900 (N_6900,N_6030,N_6421);
nor U6901 (N_6901,N_6018,N_6342);
nand U6902 (N_6902,N_6348,N_6257);
nand U6903 (N_6903,N_6090,N_6141);
xnor U6904 (N_6904,N_6010,N_6276);
or U6905 (N_6905,N_6289,N_6157);
or U6906 (N_6906,N_6308,N_6108);
nor U6907 (N_6907,N_6487,N_6359);
nand U6908 (N_6908,N_6281,N_6152);
nor U6909 (N_6909,N_6212,N_6484);
nand U6910 (N_6910,N_6166,N_6437);
nor U6911 (N_6911,N_6141,N_6121);
nor U6912 (N_6912,N_6139,N_6385);
nand U6913 (N_6913,N_6107,N_6212);
nand U6914 (N_6914,N_6263,N_6041);
xnor U6915 (N_6915,N_6152,N_6065);
nand U6916 (N_6916,N_6376,N_6392);
or U6917 (N_6917,N_6177,N_6462);
nand U6918 (N_6918,N_6449,N_6405);
nor U6919 (N_6919,N_6023,N_6292);
nand U6920 (N_6920,N_6336,N_6008);
xnor U6921 (N_6921,N_6054,N_6448);
xor U6922 (N_6922,N_6207,N_6356);
or U6923 (N_6923,N_6162,N_6204);
and U6924 (N_6924,N_6295,N_6426);
or U6925 (N_6925,N_6227,N_6477);
xnor U6926 (N_6926,N_6292,N_6449);
and U6927 (N_6927,N_6068,N_6493);
xor U6928 (N_6928,N_6352,N_6372);
or U6929 (N_6929,N_6340,N_6235);
and U6930 (N_6930,N_6215,N_6357);
and U6931 (N_6931,N_6024,N_6489);
and U6932 (N_6932,N_6471,N_6012);
or U6933 (N_6933,N_6455,N_6341);
or U6934 (N_6934,N_6025,N_6409);
or U6935 (N_6935,N_6497,N_6035);
and U6936 (N_6936,N_6486,N_6149);
nor U6937 (N_6937,N_6356,N_6329);
nor U6938 (N_6938,N_6013,N_6316);
or U6939 (N_6939,N_6185,N_6284);
xor U6940 (N_6940,N_6057,N_6209);
nand U6941 (N_6941,N_6314,N_6447);
nand U6942 (N_6942,N_6471,N_6177);
and U6943 (N_6943,N_6210,N_6326);
nor U6944 (N_6944,N_6442,N_6039);
nand U6945 (N_6945,N_6009,N_6145);
xnor U6946 (N_6946,N_6089,N_6092);
xnor U6947 (N_6947,N_6313,N_6467);
nand U6948 (N_6948,N_6231,N_6239);
or U6949 (N_6949,N_6246,N_6176);
xor U6950 (N_6950,N_6458,N_6284);
nor U6951 (N_6951,N_6311,N_6025);
nand U6952 (N_6952,N_6150,N_6211);
nand U6953 (N_6953,N_6339,N_6495);
and U6954 (N_6954,N_6006,N_6264);
xnor U6955 (N_6955,N_6058,N_6222);
nand U6956 (N_6956,N_6475,N_6478);
or U6957 (N_6957,N_6431,N_6357);
nand U6958 (N_6958,N_6497,N_6335);
xnor U6959 (N_6959,N_6062,N_6329);
and U6960 (N_6960,N_6407,N_6487);
nor U6961 (N_6961,N_6063,N_6243);
and U6962 (N_6962,N_6211,N_6305);
or U6963 (N_6963,N_6111,N_6292);
or U6964 (N_6964,N_6064,N_6063);
nand U6965 (N_6965,N_6416,N_6480);
nand U6966 (N_6966,N_6418,N_6086);
or U6967 (N_6967,N_6318,N_6094);
nand U6968 (N_6968,N_6008,N_6375);
and U6969 (N_6969,N_6153,N_6100);
nor U6970 (N_6970,N_6433,N_6038);
and U6971 (N_6971,N_6488,N_6275);
nand U6972 (N_6972,N_6252,N_6117);
and U6973 (N_6973,N_6427,N_6430);
xnor U6974 (N_6974,N_6432,N_6332);
nor U6975 (N_6975,N_6019,N_6005);
nand U6976 (N_6976,N_6164,N_6068);
or U6977 (N_6977,N_6425,N_6053);
nand U6978 (N_6978,N_6461,N_6124);
and U6979 (N_6979,N_6394,N_6300);
or U6980 (N_6980,N_6200,N_6308);
and U6981 (N_6981,N_6122,N_6234);
and U6982 (N_6982,N_6423,N_6266);
xnor U6983 (N_6983,N_6383,N_6231);
nand U6984 (N_6984,N_6386,N_6151);
nor U6985 (N_6985,N_6204,N_6192);
or U6986 (N_6986,N_6325,N_6438);
nand U6987 (N_6987,N_6024,N_6463);
nand U6988 (N_6988,N_6094,N_6412);
nor U6989 (N_6989,N_6456,N_6464);
nor U6990 (N_6990,N_6332,N_6465);
or U6991 (N_6991,N_6343,N_6120);
nand U6992 (N_6992,N_6405,N_6207);
nand U6993 (N_6993,N_6338,N_6481);
nor U6994 (N_6994,N_6327,N_6186);
and U6995 (N_6995,N_6059,N_6458);
xnor U6996 (N_6996,N_6035,N_6265);
or U6997 (N_6997,N_6114,N_6073);
or U6998 (N_6998,N_6399,N_6243);
xnor U6999 (N_6999,N_6298,N_6202);
xnor U7000 (N_7000,N_6873,N_6718);
and U7001 (N_7001,N_6854,N_6796);
xor U7002 (N_7002,N_6871,N_6610);
and U7003 (N_7003,N_6935,N_6754);
and U7004 (N_7004,N_6661,N_6911);
and U7005 (N_7005,N_6868,N_6933);
nand U7006 (N_7006,N_6500,N_6716);
nand U7007 (N_7007,N_6581,N_6749);
and U7008 (N_7008,N_6930,N_6870);
nand U7009 (N_7009,N_6968,N_6626);
and U7010 (N_7010,N_6770,N_6580);
and U7011 (N_7011,N_6502,N_6606);
or U7012 (N_7012,N_6746,N_6638);
and U7013 (N_7013,N_6909,N_6812);
or U7014 (N_7014,N_6691,N_6984);
and U7015 (N_7015,N_6627,N_6841);
or U7016 (N_7016,N_6510,N_6522);
and U7017 (N_7017,N_6687,N_6684);
or U7018 (N_7018,N_6863,N_6820);
nand U7019 (N_7019,N_6623,N_6750);
and U7020 (N_7020,N_6711,N_6817);
or U7021 (N_7021,N_6619,N_6617);
or U7022 (N_7022,N_6975,N_6766);
and U7023 (N_7023,N_6967,N_6989);
or U7024 (N_7024,N_6587,N_6938);
nor U7025 (N_7025,N_6825,N_6640);
xor U7026 (N_7026,N_6705,N_6700);
and U7027 (N_7027,N_6655,N_6912);
or U7028 (N_7028,N_6709,N_6887);
nand U7029 (N_7029,N_6722,N_6795);
or U7030 (N_7030,N_6620,N_6904);
xor U7031 (N_7031,N_6641,N_6890);
and U7032 (N_7032,N_6879,N_6557);
nor U7033 (N_7033,N_6925,N_6513);
and U7034 (N_7034,N_6940,N_6618);
xor U7035 (N_7035,N_6827,N_6560);
or U7036 (N_7036,N_6979,N_6877);
and U7037 (N_7037,N_6998,N_6567);
xnor U7038 (N_7038,N_6678,N_6565);
or U7039 (N_7039,N_6633,N_6538);
and U7040 (N_7040,N_6537,N_6974);
and U7041 (N_7041,N_6931,N_6927);
and U7042 (N_7042,N_6835,N_6582);
or U7043 (N_7043,N_6818,N_6710);
nor U7044 (N_7044,N_6695,N_6521);
or U7045 (N_7045,N_6954,N_6839);
and U7046 (N_7046,N_6816,N_6544);
and U7047 (N_7047,N_6571,N_6900);
or U7048 (N_7048,N_6908,N_6913);
nor U7049 (N_7049,N_6558,N_6578);
nand U7050 (N_7050,N_6759,N_6785);
nor U7051 (N_7051,N_6834,N_6692);
xnor U7052 (N_7052,N_6531,N_6595);
or U7053 (N_7053,N_6788,N_6862);
xor U7054 (N_7054,N_6650,N_6708);
xor U7055 (N_7055,N_6971,N_6823);
nand U7056 (N_7056,N_6961,N_6965);
and U7057 (N_7057,N_6952,N_6992);
or U7058 (N_7058,N_6664,N_6613);
and U7059 (N_7059,N_6985,N_6679);
and U7060 (N_7060,N_6555,N_6859);
or U7061 (N_7061,N_6955,N_6597);
xor U7062 (N_7062,N_6784,N_6808);
and U7063 (N_7063,N_6585,N_6760);
nand U7064 (N_7064,N_6986,N_6739);
nand U7065 (N_7065,N_6778,N_6880);
nor U7066 (N_7066,N_6712,N_6583);
xor U7067 (N_7067,N_6704,N_6507);
or U7068 (N_7068,N_6901,N_6864);
nand U7069 (N_7069,N_6720,N_6694);
nor U7070 (N_7070,N_6689,N_6806);
xor U7071 (N_7071,N_6781,N_6858);
nand U7072 (N_7072,N_6721,N_6636);
or U7073 (N_7073,N_6794,N_6762);
and U7074 (N_7074,N_6990,N_6801);
or U7075 (N_7075,N_6844,N_6942);
xnor U7076 (N_7076,N_6520,N_6508);
xor U7077 (N_7077,N_6574,N_6719);
or U7078 (N_7078,N_6934,N_6543);
or U7079 (N_7079,N_6630,N_6556);
and U7080 (N_7080,N_6736,N_6889);
or U7081 (N_7081,N_6973,N_6653);
and U7082 (N_7082,N_6607,N_6742);
and U7083 (N_7083,N_6811,N_6635);
or U7084 (N_7084,N_6535,N_6732);
nand U7085 (N_7085,N_6789,N_6672);
or U7086 (N_7086,N_6683,N_6956);
xnor U7087 (N_7087,N_6509,N_6591);
nor U7088 (N_7088,N_6928,N_6576);
nand U7089 (N_7089,N_6857,N_6637);
nand U7090 (N_7090,N_6939,N_6550);
and U7091 (N_7091,N_6698,N_6849);
xor U7092 (N_7092,N_6686,N_6603);
and U7093 (N_7093,N_6612,N_6920);
nand U7094 (N_7094,N_6696,N_6907);
nor U7095 (N_7095,N_6621,N_6561);
nor U7096 (N_7096,N_6847,N_6822);
or U7097 (N_7097,N_6552,N_6614);
xor U7098 (N_7098,N_6564,N_6598);
or U7099 (N_7099,N_6648,N_6645);
and U7100 (N_7100,N_6805,N_6815);
xor U7101 (N_7101,N_6504,N_6548);
nor U7102 (N_7102,N_6670,N_6734);
nand U7103 (N_7103,N_6511,N_6518);
or U7104 (N_7104,N_6562,N_6758);
nor U7105 (N_7105,N_6966,N_6671);
or U7106 (N_7106,N_6586,N_6951);
nand U7107 (N_7107,N_6833,N_6733);
or U7108 (N_7108,N_6804,N_6763);
and U7109 (N_7109,N_6897,N_6947);
nor U7110 (N_7110,N_6668,N_6830);
nand U7111 (N_7111,N_6895,N_6505);
nor U7112 (N_7112,N_6501,N_6802);
and U7113 (N_7113,N_6723,N_6737);
and U7114 (N_7114,N_6579,N_6832);
nor U7115 (N_7115,N_6950,N_6738);
nand U7116 (N_7116,N_6642,N_6919);
nand U7117 (N_7117,N_6793,N_6838);
xnor U7118 (N_7118,N_6988,N_6547);
nor U7119 (N_7119,N_6608,N_6707);
and U7120 (N_7120,N_6682,N_6876);
nand U7121 (N_7121,N_6918,N_6549);
nor U7122 (N_7122,N_6601,N_6681);
and U7123 (N_7123,N_6665,N_6765);
nor U7124 (N_7124,N_6916,N_6821);
and U7125 (N_7125,N_6546,N_6977);
xnor U7126 (N_7126,N_6753,N_6615);
nand U7127 (N_7127,N_6554,N_6569);
xor U7128 (N_7128,N_6885,N_6748);
and U7129 (N_7129,N_6660,N_6878);
xnor U7130 (N_7130,N_6590,N_6893);
or U7131 (N_7131,N_6768,N_6663);
or U7132 (N_7132,N_6755,N_6667);
nand U7133 (N_7133,N_6514,N_6829);
or U7134 (N_7134,N_6570,N_6563);
nor U7135 (N_7135,N_6775,N_6525);
or U7136 (N_7136,N_6851,N_6976);
or U7137 (N_7137,N_6905,N_6730);
or U7138 (N_7138,N_6631,N_6756);
or U7139 (N_7139,N_6814,N_6970);
xor U7140 (N_7140,N_6943,N_6809);
nand U7141 (N_7141,N_6677,N_6790);
or U7142 (N_7142,N_6972,N_6588);
or U7143 (N_7143,N_6899,N_6803);
nand U7144 (N_7144,N_6884,N_6517);
and U7145 (N_7145,N_6741,N_6902);
xnor U7146 (N_7146,N_6852,N_6875);
or U7147 (N_7147,N_6800,N_6532);
and U7148 (N_7148,N_6503,N_6666);
and U7149 (N_7149,N_6725,N_6969);
nand U7150 (N_7150,N_6945,N_6850);
nor U7151 (N_7151,N_6837,N_6728);
or U7152 (N_7152,N_6602,N_6553);
xnor U7153 (N_7153,N_6680,N_6632);
xor U7154 (N_7154,N_6639,N_6515);
and U7155 (N_7155,N_6924,N_6752);
nor U7156 (N_7156,N_6991,N_6669);
nor U7157 (N_7157,N_6528,N_6605);
or U7158 (N_7158,N_6964,N_6724);
and U7159 (N_7159,N_6519,N_6926);
xnor U7160 (N_7160,N_6516,N_6600);
xnor U7161 (N_7161,N_6656,N_6810);
and U7162 (N_7162,N_6922,N_6845);
and U7163 (N_7163,N_6995,N_6886);
and U7164 (N_7164,N_6596,N_6717);
xnor U7165 (N_7165,N_6616,N_6727);
and U7166 (N_7166,N_6949,N_6512);
nor U7167 (N_7167,N_6767,N_6959);
xor U7168 (N_7168,N_6757,N_6575);
or U7169 (N_7169,N_6994,N_6828);
xnor U7170 (N_7170,N_6624,N_6798);
xor U7171 (N_7171,N_6688,N_6882);
or U7172 (N_7172,N_6604,N_6651);
nor U7173 (N_7173,N_6978,N_6731);
nor U7174 (N_7174,N_6853,N_6874);
nor U7175 (N_7175,N_6568,N_6894);
nor U7176 (N_7176,N_6764,N_6846);
and U7177 (N_7177,N_6848,N_6921);
and U7178 (N_7178,N_6843,N_6892);
nand U7179 (N_7179,N_6527,N_6799);
xor U7180 (N_7180,N_6948,N_6826);
nor U7181 (N_7181,N_6609,N_6960);
nand U7182 (N_7182,N_6644,N_6628);
or U7183 (N_7183,N_6963,N_6714);
nor U7184 (N_7184,N_6540,N_6903);
xor U7185 (N_7185,N_6593,N_6906);
xnor U7186 (N_7186,N_6744,N_6780);
and U7187 (N_7187,N_6701,N_6779);
nor U7188 (N_7188,N_6888,N_6654);
nor U7189 (N_7189,N_6713,N_6923);
or U7190 (N_7190,N_6962,N_6634);
xor U7191 (N_7191,N_6577,N_6611);
xor U7192 (N_7192,N_6566,N_6869);
xor U7193 (N_7193,N_6898,N_6840);
and U7194 (N_7194,N_6944,N_6813);
xor U7195 (N_7195,N_6551,N_6958);
nand U7196 (N_7196,N_6774,N_6524);
and U7197 (N_7197,N_6771,N_6526);
or U7198 (N_7198,N_6915,N_6659);
xor U7199 (N_7199,N_6860,N_6594);
and U7200 (N_7200,N_6941,N_6536);
xor U7201 (N_7201,N_6745,N_6523);
nor U7202 (N_7202,N_6676,N_6539);
nor U7203 (N_7203,N_6541,N_6861);
and U7204 (N_7204,N_6751,N_6831);
nand U7205 (N_7205,N_6572,N_6592);
nor U7206 (N_7206,N_6983,N_6530);
and U7207 (N_7207,N_6652,N_6647);
and U7208 (N_7208,N_6629,N_6693);
and U7209 (N_7209,N_6910,N_6792);
nand U7210 (N_7210,N_6881,N_6929);
nand U7211 (N_7211,N_6896,N_6545);
nor U7212 (N_7212,N_6706,N_6534);
and U7213 (N_7213,N_6891,N_6957);
nor U7214 (N_7214,N_6740,N_6743);
nand U7215 (N_7215,N_6883,N_6726);
nor U7216 (N_7216,N_6715,N_6787);
and U7217 (N_7217,N_6993,N_6622);
and U7218 (N_7218,N_6932,N_6657);
nand U7219 (N_7219,N_6842,N_6865);
nand U7220 (N_7220,N_6953,N_6776);
xor U7221 (N_7221,N_6782,N_6777);
and U7222 (N_7222,N_6773,N_6855);
nor U7223 (N_7223,N_6769,N_6836);
or U7224 (N_7224,N_6542,N_6658);
or U7225 (N_7225,N_6673,N_6791);
nor U7226 (N_7226,N_6702,N_6761);
xor U7227 (N_7227,N_6735,N_6690);
nor U7228 (N_7228,N_6573,N_6999);
nor U7229 (N_7229,N_6982,N_6786);
and U7230 (N_7230,N_6936,N_6866);
nor U7231 (N_7231,N_6937,N_6649);
nand U7232 (N_7232,N_6703,N_6643);
nand U7233 (N_7233,N_6867,N_6917);
nand U7234 (N_7234,N_6981,N_6872);
nor U7235 (N_7235,N_6697,N_6699);
nor U7236 (N_7236,N_6819,N_6807);
xor U7237 (N_7237,N_6625,N_6589);
nor U7238 (N_7238,N_6674,N_6856);
nand U7239 (N_7239,N_6747,N_6824);
nand U7240 (N_7240,N_6946,N_6783);
or U7241 (N_7241,N_6675,N_6662);
xor U7242 (N_7242,N_6599,N_6914);
and U7243 (N_7243,N_6529,N_6729);
xor U7244 (N_7244,N_6996,N_6559);
nand U7245 (N_7245,N_6685,N_6506);
nor U7246 (N_7246,N_6797,N_6646);
or U7247 (N_7247,N_6533,N_6584);
nand U7248 (N_7248,N_6772,N_6987);
xnor U7249 (N_7249,N_6980,N_6997);
or U7250 (N_7250,N_6998,N_6601);
or U7251 (N_7251,N_6779,N_6633);
nand U7252 (N_7252,N_6955,N_6654);
or U7253 (N_7253,N_6626,N_6505);
nand U7254 (N_7254,N_6546,N_6562);
and U7255 (N_7255,N_6678,N_6681);
and U7256 (N_7256,N_6721,N_6634);
nand U7257 (N_7257,N_6583,N_6510);
and U7258 (N_7258,N_6500,N_6819);
nand U7259 (N_7259,N_6562,N_6665);
and U7260 (N_7260,N_6615,N_6839);
xor U7261 (N_7261,N_6527,N_6850);
or U7262 (N_7262,N_6615,N_6680);
nor U7263 (N_7263,N_6610,N_6608);
xnor U7264 (N_7264,N_6716,N_6753);
nand U7265 (N_7265,N_6930,N_6828);
or U7266 (N_7266,N_6578,N_6858);
nand U7267 (N_7267,N_6819,N_6920);
nand U7268 (N_7268,N_6781,N_6822);
and U7269 (N_7269,N_6514,N_6649);
xor U7270 (N_7270,N_6703,N_6750);
nor U7271 (N_7271,N_6651,N_6566);
and U7272 (N_7272,N_6763,N_6787);
or U7273 (N_7273,N_6773,N_6924);
nand U7274 (N_7274,N_6528,N_6926);
and U7275 (N_7275,N_6987,N_6642);
nand U7276 (N_7276,N_6649,N_6681);
nor U7277 (N_7277,N_6988,N_6930);
and U7278 (N_7278,N_6873,N_6665);
or U7279 (N_7279,N_6812,N_6927);
xor U7280 (N_7280,N_6517,N_6792);
xnor U7281 (N_7281,N_6537,N_6550);
or U7282 (N_7282,N_6762,N_6791);
or U7283 (N_7283,N_6981,N_6858);
nand U7284 (N_7284,N_6677,N_6596);
nand U7285 (N_7285,N_6838,N_6842);
nor U7286 (N_7286,N_6986,N_6814);
and U7287 (N_7287,N_6889,N_6668);
or U7288 (N_7288,N_6715,N_6692);
nand U7289 (N_7289,N_6581,N_6735);
and U7290 (N_7290,N_6688,N_6773);
xor U7291 (N_7291,N_6856,N_6890);
and U7292 (N_7292,N_6817,N_6992);
or U7293 (N_7293,N_6741,N_6730);
xnor U7294 (N_7294,N_6859,N_6933);
nand U7295 (N_7295,N_6529,N_6846);
nand U7296 (N_7296,N_6866,N_6768);
xor U7297 (N_7297,N_6846,N_6669);
and U7298 (N_7298,N_6788,N_6879);
nand U7299 (N_7299,N_6990,N_6543);
nand U7300 (N_7300,N_6684,N_6928);
or U7301 (N_7301,N_6642,N_6571);
nand U7302 (N_7302,N_6504,N_6716);
nor U7303 (N_7303,N_6540,N_6926);
and U7304 (N_7304,N_6650,N_6533);
nand U7305 (N_7305,N_6538,N_6722);
nand U7306 (N_7306,N_6528,N_6919);
nand U7307 (N_7307,N_6941,N_6749);
xnor U7308 (N_7308,N_6992,N_6968);
nor U7309 (N_7309,N_6831,N_6923);
or U7310 (N_7310,N_6634,N_6867);
or U7311 (N_7311,N_6766,N_6882);
nor U7312 (N_7312,N_6914,N_6698);
xor U7313 (N_7313,N_6852,N_6773);
or U7314 (N_7314,N_6851,N_6637);
nor U7315 (N_7315,N_6719,N_6890);
or U7316 (N_7316,N_6803,N_6630);
nor U7317 (N_7317,N_6591,N_6665);
nand U7318 (N_7318,N_6854,N_6932);
nor U7319 (N_7319,N_6626,N_6762);
xnor U7320 (N_7320,N_6500,N_6671);
xor U7321 (N_7321,N_6650,N_6866);
nand U7322 (N_7322,N_6791,N_6953);
nand U7323 (N_7323,N_6911,N_6654);
nand U7324 (N_7324,N_6909,N_6766);
nand U7325 (N_7325,N_6876,N_6561);
xor U7326 (N_7326,N_6572,N_6820);
nand U7327 (N_7327,N_6543,N_6643);
or U7328 (N_7328,N_6559,N_6600);
xor U7329 (N_7329,N_6507,N_6642);
nor U7330 (N_7330,N_6693,N_6843);
or U7331 (N_7331,N_6589,N_6691);
xor U7332 (N_7332,N_6827,N_6743);
nor U7333 (N_7333,N_6682,N_6980);
xor U7334 (N_7334,N_6687,N_6559);
nor U7335 (N_7335,N_6932,N_6997);
nor U7336 (N_7336,N_6801,N_6566);
nand U7337 (N_7337,N_6508,N_6649);
or U7338 (N_7338,N_6612,N_6780);
nand U7339 (N_7339,N_6831,N_6856);
xor U7340 (N_7340,N_6736,N_6609);
nand U7341 (N_7341,N_6944,N_6523);
xnor U7342 (N_7342,N_6704,N_6674);
nor U7343 (N_7343,N_6871,N_6896);
or U7344 (N_7344,N_6663,N_6660);
or U7345 (N_7345,N_6970,N_6652);
and U7346 (N_7346,N_6560,N_6505);
nor U7347 (N_7347,N_6581,N_6671);
xor U7348 (N_7348,N_6592,N_6617);
and U7349 (N_7349,N_6552,N_6889);
nand U7350 (N_7350,N_6631,N_6971);
or U7351 (N_7351,N_6577,N_6990);
nand U7352 (N_7352,N_6995,N_6989);
nand U7353 (N_7353,N_6629,N_6957);
xor U7354 (N_7354,N_6560,N_6502);
nor U7355 (N_7355,N_6879,N_6653);
or U7356 (N_7356,N_6888,N_6866);
xnor U7357 (N_7357,N_6804,N_6718);
nor U7358 (N_7358,N_6538,N_6892);
nand U7359 (N_7359,N_6986,N_6754);
or U7360 (N_7360,N_6703,N_6655);
nand U7361 (N_7361,N_6719,N_6958);
or U7362 (N_7362,N_6947,N_6835);
nand U7363 (N_7363,N_6801,N_6805);
and U7364 (N_7364,N_6645,N_6840);
or U7365 (N_7365,N_6896,N_6945);
xor U7366 (N_7366,N_6978,N_6542);
nand U7367 (N_7367,N_6654,N_6765);
and U7368 (N_7368,N_6543,N_6827);
nor U7369 (N_7369,N_6957,N_6633);
or U7370 (N_7370,N_6540,N_6805);
nor U7371 (N_7371,N_6699,N_6843);
nor U7372 (N_7372,N_6519,N_6618);
xor U7373 (N_7373,N_6750,N_6933);
and U7374 (N_7374,N_6855,N_6615);
xor U7375 (N_7375,N_6738,N_6821);
xnor U7376 (N_7376,N_6619,N_6938);
xnor U7377 (N_7377,N_6553,N_6616);
nand U7378 (N_7378,N_6852,N_6531);
nor U7379 (N_7379,N_6891,N_6584);
and U7380 (N_7380,N_6529,N_6536);
xnor U7381 (N_7381,N_6946,N_6952);
nand U7382 (N_7382,N_6818,N_6892);
or U7383 (N_7383,N_6760,N_6658);
or U7384 (N_7384,N_6863,N_6650);
and U7385 (N_7385,N_6614,N_6626);
nand U7386 (N_7386,N_6677,N_6688);
or U7387 (N_7387,N_6639,N_6948);
or U7388 (N_7388,N_6888,N_6933);
nand U7389 (N_7389,N_6982,N_6619);
nand U7390 (N_7390,N_6786,N_6922);
xnor U7391 (N_7391,N_6862,N_6952);
nand U7392 (N_7392,N_6638,N_6839);
or U7393 (N_7393,N_6776,N_6807);
nand U7394 (N_7394,N_6727,N_6536);
and U7395 (N_7395,N_6707,N_6592);
nand U7396 (N_7396,N_6590,N_6610);
nor U7397 (N_7397,N_6952,N_6718);
nor U7398 (N_7398,N_6829,N_6782);
nor U7399 (N_7399,N_6994,N_6796);
and U7400 (N_7400,N_6508,N_6660);
xor U7401 (N_7401,N_6542,N_6846);
and U7402 (N_7402,N_6567,N_6574);
and U7403 (N_7403,N_6955,N_6556);
or U7404 (N_7404,N_6791,N_6664);
nor U7405 (N_7405,N_6667,N_6996);
and U7406 (N_7406,N_6801,N_6770);
xor U7407 (N_7407,N_6712,N_6528);
or U7408 (N_7408,N_6629,N_6624);
or U7409 (N_7409,N_6754,N_6689);
xnor U7410 (N_7410,N_6883,N_6812);
nor U7411 (N_7411,N_6769,N_6851);
or U7412 (N_7412,N_6643,N_6939);
xor U7413 (N_7413,N_6781,N_6849);
xnor U7414 (N_7414,N_6833,N_6981);
and U7415 (N_7415,N_6988,N_6910);
xor U7416 (N_7416,N_6530,N_6575);
nand U7417 (N_7417,N_6920,N_6893);
and U7418 (N_7418,N_6629,N_6673);
nor U7419 (N_7419,N_6616,N_6519);
nor U7420 (N_7420,N_6583,N_6752);
nor U7421 (N_7421,N_6558,N_6562);
nor U7422 (N_7422,N_6926,N_6760);
nand U7423 (N_7423,N_6707,N_6858);
and U7424 (N_7424,N_6922,N_6732);
and U7425 (N_7425,N_6987,N_6907);
and U7426 (N_7426,N_6634,N_6756);
or U7427 (N_7427,N_6799,N_6768);
and U7428 (N_7428,N_6747,N_6812);
nand U7429 (N_7429,N_6512,N_6944);
nor U7430 (N_7430,N_6978,N_6700);
or U7431 (N_7431,N_6780,N_6719);
nand U7432 (N_7432,N_6698,N_6717);
and U7433 (N_7433,N_6758,N_6720);
or U7434 (N_7434,N_6774,N_6554);
nand U7435 (N_7435,N_6775,N_6599);
nor U7436 (N_7436,N_6810,N_6919);
and U7437 (N_7437,N_6649,N_6803);
nor U7438 (N_7438,N_6642,N_6745);
nor U7439 (N_7439,N_6554,N_6990);
or U7440 (N_7440,N_6653,N_6928);
nor U7441 (N_7441,N_6917,N_6557);
or U7442 (N_7442,N_6594,N_6704);
nor U7443 (N_7443,N_6759,N_6692);
or U7444 (N_7444,N_6582,N_6671);
xnor U7445 (N_7445,N_6689,N_6549);
nand U7446 (N_7446,N_6728,N_6813);
nor U7447 (N_7447,N_6619,N_6725);
or U7448 (N_7448,N_6908,N_6759);
xor U7449 (N_7449,N_6794,N_6756);
nand U7450 (N_7450,N_6743,N_6759);
nand U7451 (N_7451,N_6651,N_6574);
and U7452 (N_7452,N_6827,N_6898);
xor U7453 (N_7453,N_6501,N_6807);
or U7454 (N_7454,N_6937,N_6722);
nor U7455 (N_7455,N_6913,N_6866);
or U7456 (N_7456,N_6640,N_6608);
nor U7457 (N_7457,N_6575,N_6956);
and U7458 (N_7458,N_6867,N_6696);
or U7459 (N_7459,N_6675,N_6915);
nor U7460 (N_7460,N_6910,N_6843);
xnor U7461 (N_7461,N_6712,N_6593);
nor U7462 (N_7462,N_6971,N_6959);
or U7463 (N_7463,N_6972,N_6605);
or U7464 (N_7464,N_6775,N_6579);
or U7465 (N_7465,N_6549,N_6873);
xor U7466 (N_7466,N_6884,N_6970);
xor U7467 (N_7467,N_6811,N_6530);
nor U7468 (N_7468,N_6780,N_6724);
and U7469 (N_7469,N_6664,N_6580);
nor U7470 (N_7470,N_6962,N_6505);
xor U7471 (N_7471,N_6828,N_6810);
xor U7472 (N_7472,N_6752,N_6563);
nor U7473 (N_7473,N_6855,N_6529);
nand U7474 (N_7474,N_6675,N_6838);
and U7475 (N_7475,N_6987,N_6524);
and U7476 (N_7476,N_6961,N_6511);
or U7477 (N_7477,N_6559,N_6577);
nand U7478 (N_7478,N_6905,N_6702);
xor U7479 (N_7479,N_6739,N_6742);
or U7480 (N_7480,N_6656,N_6909);
nor U7481 (N_7481,N_6891,N_6509);
and U7482 (N_7482,N_6890,N_6525);
and U7483 (N_7483,N_6542,N_6502);
nand U7484 (N_7484,N_6693,N_6895);
and U7485 (N_7485,N_6933,N_6819);
xnor U7486 (N_7486,N_6950,N_6881);
and U7487 (N_7487,N_6947,N_6860);
or U7488 (N_7488,N_6986,N_6985);
nand U7489 (N_7489,N_6504,N_6551);
nand U7490 (N_7490,N_6955,N_6603);
nand U7491 (N_7491,N_6919,N_6838);
nor U7492 (N_7492,N_6543,N_6583);
and U7493 (N_7493,N_6900,N_6666);
xor U7494 (N_7494,N_6784,N_6511);
xor U7495 (N_7495,N_6887,N_6906);
and U7496 (N_7496,N_6923,N_6755);
nand U7497 (N_7497,N_6957,N_6871);
nor U7498 (N_7498,N_6920,N_6991);
and U7499 (N_7499,N_6857,N_6679);
nor U7500 (N_7500,N_7498,N_7146);
or U7501 (N_7501,N_7260,N_7081);
nor U7502 (N_7502,N_7021,N_7065);
xor U7503 (N_7503,N_7332,N_7376);
and U7504 (N_7504,N_7040,N_7417);
nand U7505 (N_7505,N_7177,N_7261);
xor U7506 (N_7506,N_7351,N_7272);
or U7507 (N_7507,N_7025,N_7475);
xnor U7508 (N_7508,N_7124,N_7147);
nor U7509 (N_7509,N_7467,N_7002);
nand U7510 (N_7510,N_7200,N_7201);
nor U7511 (N_7511,N_7275,N_7449);
xor U7512 (N_7512,N_7185,N_7056);
or U7513 (N_7513,N_7127,N_7446);
nor U7514 (N_7514,N_7120,N_7335);
nor U7515 (N_7515,N_7368,N_7122);
nor U7516 (N_7516,N_7451,N_7284);
and U7517 (N_7517,N_7315,N_7270);
or U7518 (N_7518,N_7219,N_7349);
and U7519 (N_7519,N_7393,N_7344);
nand U7520 (N_7520,N_7019,N_7080);
xnor U7521 (N_7521,N_7194,N_7346);
nor U7522 (N_7522,N_7366,N_7231);
nand U7523 (N_7523,N_7391,N_7059);
nor U7524 (N_7524,N_7278,N_7265);
nor U7525 (N_7525,N_7064,N_7497);
nor U7526 (N_7526,N_7115,N_7015);
nand U7527 (N_7527,N_7092,N_7212);
nand U7528 (N_7528,N_7420,N_7104);
or U7529 (N_7529,N_7189,N_7378);
nor U7530 (N_7530,N_7471,N_7214);
nand U7531 (N_7531,N_7439,N_7491);
nand U7532 (N_7532,N_7241,N_7360);
or U7533 (N_7533,N_7448,N_7145);
or U7534 (N_7534,N_7271,N_7313);
or U7535 (N_7535,N_7269,N_7342);
and U7536 (N_7536,N_7428,N_7061);
nand U7537 (N_7537,N_7049,N_7459);
nand U7538 (N_7538,N_7257,N_7247);
and U7539 (N_7539,N_7401,N_7184);
xor U7540 (N_7540,N_7440,N_7091);
nand U7541 (N_7541,N_7418,N_7388);
and U7542 (N_7542,N_7217,N_7097);
nor U7543 (N_7543,N_7340,N_7051);
nand U7544 (N_7544,N_7263,N_7044);
xor U7545 (N_7545,N_7370,N_7159);
and U7546 (N_7546,N_7469,N_7282);
and U7547 (N_7547,N_7211,N_7453);
nor U7548 (N_7548,N_7011,N_7334);
nand U7549 (N_7549,N_7310,N_7208);
nor U7550 (N_7550,N_7010,N_7390);
nor U7551 (N_7551,N_7224,N_7238);
xnor U7552 (N_7552,N_7033,N_7389);
xnor U7553 (N_7553,N_7307,N_7109);
or U7554 (N_7554,N_7431,N_7038);
xor U7555 (N_7555,N_7444,N_7112);
nand U7556 (N_7556,N_7007,N_7287);
nor U7557 (N_7557,N_7487,N_7377);
or U7558 (N_7558,N_7463,N_7317);
nor U7559 (N_7559,N_7402,N_7465);
and U7560 (N_7560,N_7365,N_7165);
nand U7561 (N_7561,N_7062,N_7020);
and U7562 (N_7562,N_7077,N_7476);
nand U7563 (N_7563,N_7470,N_7462);
nand U7564 (N_7564,N_7041,N_7464);
and U7565 (N_7565,N_7216,N_7111);
xor U7566 (N_7566,N_7244,N_7142);
nand U7567 (N_7567,N_7379,N_7399);
nor U7568 (N_7568,N_7255,N_7037);
or U7569 (N_7569,N_7005,N_7302);
or U7570 (N_7570,N_7098,N_7067);
xnor U7571 (N_7571,N_7437,N_7006);
and U7572 (N_7572,N_7234,N_7358);
and U7573 (N_7573,N_7477,N_7450);
nor U7574 (N_7574,N_7248,N_7350);
xnor U7575 (N_7575,N_7172,N_7353);
and U7576 (N_7576,N_7071,N_7482);
and U7577 (N_7577,N_7429,N_7423);
nor U7578 (N_7578,N_7249,N_7032);
and U7579 (N_7579,N_7012,N_7093);
nand U7580 (N_7580,N_7452,N_7341);
nor U7581 (N_7581,N_7321,N_7083);
or U7582 (N_7582,N_7144,N_7156);
nand U7583 (N_7583,N_7347,N_7001);
and U7584 (N_7584,N_7055,N_7298);
or U7585 (N_7585,N_7186,N_7179);
nor U7586 (N_7586,N_7096,N_7014);
xor U7587 (N_7587,N_7094,N_7395);
xnor U7588 (N_7588,N_7430,N_7258);
and U7589 (N_7589,N_7008,N_7246);
or U7590 (N_7590,N_7057,N_7494);
nor U7591 (N_7591,N_7447,N_7100);
nor U7592 (N_7592,N_7264,N_7461);
nand U7593 (N_7593,N_7496,N_7023);
nor U7594 (N_7594,N_7394,N_7387);
or U7595 (N_7595,N_7196,N_7419);
and U7596 (N_7596,N_7410,N_7408);
or U7597 (N_7597,N_7213,N_7054);
nor U7598 (N_7598,N_7103,N_7045);
nand U7599 (N_7599,N_7132,N_7352);
nor U7600 (N_7600,N_7336,N_7000);
and U7601 (N_7601,N_7082,N_7375);
and U7602 (N_7602,N_7004,N_7076);
nor U7603 (N_7603,N_7027,N_7286);
and U7604 (N_7604,N_7479,N_7130);
xnor U7605 (N_7605,N_7079,N_7193);
nor U7606 (N_7606,N_7424,N_7039);
nand U7607 (N_7607,N_7236,N_7293);
nor U7608 (N_7608,N_7297,N_7288);
or U7609 (N_7609,N_7114,N_7279);
and U7610 (N_7610,N_7119,N_7035);
nand U7611 (N_7611,N_7228,N_7308);
nor U7612 (N_7612,N_7421,N_7170);
and U7613 (N_7613,N_7309,N_7210);
nor U7614 (N_7614,N_7303,N_7171);
and U7615 (N_7615,N_7267,N_7441);
or U7616 (N_7616,N_7187,N_7473);
and U7617 (N_7617,N_7233,N_7197);
and U7618 (N_7618,N_7486,N_7483);
xor U7619 (N_7619,N_7253,N_7403);
and U7620 (N_7620,N_7128,N_7058);
nand U7621 (N_7621,N_7405,N_7325);
xor U7622 (N_7622,N_7031,N_7140);
or U7623 (N_7623,N_7169,N_7204);
xor U7624 (N_7624,N_7474,N_7126);
xnor U7625 (N_7625,N_7074,N_7289);
and U7626 (N_7626,N_7359,N_7443);
or U7627 (N_7627,N_7392,N_7131);
xnor U7628 (N_7628,N_7036,N_7090);
nor U7629 (N_7629,N_7356,N_7283);
and U7630 (N_7630,N_7151,N_7101);
xor U7631 (N_7631,N_7239,N_7295);
nor U7632 (N_7632,N_7107,N_7316);
nor U7633 (N_7633,N_7409,N_7488);
nor U7634 (N_7634,N_7043,N_7285);
nand U7635 (N_7635,N_7398,N_7337);
nand U7636 (N_7636,N_7268,N_7277);
and U7637 (N_7637,N_7426,N_7125);
and U7638 (N_7638,N_7415,N_7445);
or U7639 (N_7639,N_7078,N_7118);
xnor U7640 (N_7640,N_7180,N_7138);
or U7641 (N_7641,N_7085,N_7427);
nor U7642 (N_7642,N_7134,N_7361);
or U7643 (N_7643,N_7195,N_7385);
xnor U7644 (N_7644,N_7484,N_7243);
nor U7645 (N_7645,N_7068,N_7318);
nand U7646 (N_7646,N_7167,N_7312);
or U7647 (N_7647,N_7164,N_7442);
or U7648 (N_7648,N_7306,N_7183);
or U7649 (N_7649,N_7137,N_7129);
nor U7650 (N_7650,N_7225,N_7468);
nand U7651 (N_7651,N_7148,N_7320);
xnor U7652 (N_7652,N_7017,N_7075);
nor U7653 (N_7653,N_7139,N_7034);
xor U7654 (N_7654,N_7113,N_7291);
xnor U7655 (N_7655,N_7086,N_7173);
and U7656 (N_7656,N_7181,N_7105);
and U7657 (N_7657,N_7456,N_7163);
or U7658 (N_7658,N_7435,N_7072);
or U7659 (N_7659,N_7157,N_7324);
nand U7660 (N_7660,N_7220,N_7262);
nor U7661 (N_7661,N_7161,N_7191);
xnor U7662 (N_7662,N_7481,N_7136);
nand U7663 (N_7663,N_7357,N_7089);
xor U7664 (N_7664,N_7158,N_7251);
and U7665 (N_7665,N_7434,N_7371);
nand U7666 (N_7666,N_7455,N_7460);
or U7667 (N_7667,N_7386,N_7382);
or U7668 (N_7668,N_7182,N_7166);
xor U7669 (N_7669,N_7489,N_7478);
xor U7670 (N_7670,N_7102,N_7454);
and U7671 (N_7671,N_7205,N_7466);
nor U7672 (N_7672,N_7168,N_7354);
or U7673 (N_7673,N_7432,N_7070);
and U7674 (N_7674,N_7372,N_7229);
nand U7675 (N_7675,N_7150,N_7493);
xnor U7676 (N_7676,N_7333,N_7304);
and U7677 (N_7677,N_7433,N_7227);
or U7678 (N_7678,N_7422,N_7198);
or U7679 (N_7679,N_7235,N_7190);
nor U7680 (N_7680,N_7322,N_7222);
xnor U7681 (N_7681,N_7328,N_7117);
or U7682 (N_7682,N_7296,N_7259);
nor U7683 (N_7683,N_7053,N_7276);
nand U7684 (N_7684,N_7013,N_7381);
and U7685 (N_7685,N_7123,N_7343);
nand U7686 (N_7686,N_7492,N_7206);
or U7687 (N_7687,N_7363,N_7273);
xor U7688 (N_7688,N_7022,N_7254);
xnor U7689 (N_7689,N_7106,N_7030);
nand U7690 (N_7690,N_7345,N_7348);
nor U7691 (N_7691,N_7485,N_7199);
or U7692 (N_7692,N_7373,N_7202);
or U7693 (N_7693,N_7162,N_7028);
nand U7694 (N_7694,N_7406,N_7226);
nand U7695 (N_7695,N_7384,N_7438);
or U7696 (N_7696,N_7047,N_7149);
and U7697 (N_7697,N_7160,N_7069);
nor U7698 (N_7698,N_7153,N_7018);
or U7699 (N_7699,N_7141,N_7073);
or U7700 (N_7700,N_7188,N_7436);
nor U7701 (N_7701,N_7084,N_7330);
xor U7702 (N_7702,N_7060,N_7294);
nor U7703 (N_7703,N_7338,N_7411);
and U7704 (N_7704,N_7135,N_7397);
nand U7705 (N_7705,N_7274,N_7300);
nor U7706 (N_7706,N_7009,N_7480);
and U7707 (N_7707,N_7490,N_7108);
or U7708 (N_7708,N_7245,N_7425);
xor U7709 (N_7709,N_7024,N_7412);
nor U7710 (N_7710,N_7016,N_7063);
or U7711 (N_7711,N_7046,N_7299);
nor U7712 (N_7712,N_7116,N_7499);
xnor U7713 (N_7713,N_7230,N_7369);
xor U7714 (N_7714,N_7301,N_7305);
or U7715 (N_7715,N_7280,N_7052);
xor U7716 (N_7716,N_7413,N_7133);
nand U7717 (N_7717,N_7457,N_7250);
xor U7718 (N_7718,N_7292,N_7314);
nand U7719 (N_7719,N_7174,N_7311);
nor U7720 (N_7720,N_7209,N_7290);
xor U7721 (N_7721,N_7240,N_7042);
nor U7722 (N_7722,N_7331,N_7203);
nand U7723 (N_7723,N_7026,N_7364);
nor U7724 (N_7724,N_7003,N_7066);
nand U7725 (N_7725,N_7266,N_7327);
or U7726 (N_7726,N_7383,N_7192);
nor U7727 (N_7727,N_7029,N_7458);
nor U7728 (N_7728,N_7110,N_7099);
nand U7729 (N_7729,N_7326,N_7256);
or U7730 (N_7730,N_7319,N_7088);
xnor U7731 (N_7731,N_7242,N_7218);
or U7732 (N_7732,N_7367,N_7281);
xnor U7733 (N_7733,N_7472,N_7237);
and U7734 (N_7734,N_7329,N_7155);
nand U7735 (N_7735,N_7121,N_7339);
or U7736 (N_7736,N_7176,N_7223);
and U7737 (N_7737,N_7095,N_7048);
nor U7738 (N_7738,N_7416,N_7396);
and U7739 (N_7739,N_7221,N_7087);
nor U7740 (N_7740,N_7175,N_7143);
nor U7741 (N_7741,N_7404,N_7400);
or U7742 (N_7742,N_7380,N_7252);
or U7743 (N_7743,N_7178,N_7154);
and U7744 (N_7744,N_7407,N_7362);
or U7745 (N_7745,N_7050,N_7152);
nor U7746 (N_7746,N_7232,N_7215);
and U7747 (N_7747,N_7355,N_7495);
nor U7748 (N_7748,N_7323,N_7207);
nand U7749 (N_7749,N_7374,N_7414);
or U7750 (N_7750,N_7031,N_7042);
and U7751 (N_7751,N_7380,N_7183);
nor U7752 (N_7752,N_7305,N_7275);
nand U7753 (N_7753,N_7497,N_7468);
or U7754 (N_7754,N_7179,N_7386);
nor U7755 (N_7755,N_7222,N_7078);
or U7756 (N_7756,N_7046,N_7068);
nor U7757 (N_7757,N_7322,N_7000);
xor U7758 (N_7758,N_7036,N_7264);
nand U7759 (N_7759,N_7279,N_7428);
xnor U7760 (N_7760,N_7263,N_7075);
nor U7761 (N_7761,N_7468,N_7411);
xnor U7762 (N_7762,N_7400,N_7361);
or U7763 (N_7763,N_7489,N_7440);
and U7764 (N_7764,N_7145,N_7116);
nor U7765 (N_7765,N_7483,N_7337);
or U7766 (N_7766,N_7368,N_7343);
nand U7767 (N_7767,N_7467,N_7489);
and U7768 (N_7768,N_7201,N_7082);
xnor U7769 (N_7769,N_7045,N_7382);
nand U7770 (N_7770,N_7457,N_7291);
xor U7771 (N_7771,N_7074,N_7212);
nor U7772 (N_7772,N_7125,N_7174);
and U7773 (N_7773,N_7100,N_7449);
nand U7774 (N_7774,N_7143,N_7255);
nor U7775 (N_7775,N_7114,N_7122);
or U7776 (N_7776,N_7426,N_7480);
nor U7777 (N_7777,N_7188,N_7447);
nand U7778 (N_7778,N_7467,N_7147);
nand U7779 (N_7779,N_7226,N_7212);
or U7780 (N_7780,N_7440,N_7083);
xnor U7781 (N_7781,N_7333,N_7103);
or U7782 (N_7782,N_7339,N_7418);
nand U7783 (N_7783,N_7239,N_7487);
nand U7784 (N_7784,N_7304,N_7150);
nor U7785 (N_7785,N_7163,N_7476);
nand U7786 (N_7786,N_7351,N_7192);
xor U7787 (N_7787,N_7440,N_7185);
or U7788 (N_7788,N_7369,N_7004);
nand U7789 (N_7789,N_7347,N_7358);
or U7790 (N_7790,N_7060,N_7075);
nand U7791 (N_7791,N_7499,N_7295);
xor U7792 (N_7792,N_7326,N_7038);
or U7793 (N_7793,N_7171,N_7202);
and U7794 (N_7794,N_7276,N_7295);
nand U7795 (N_7795,N_7068,N_7012);
xor U7796 (N_7796,N_7148,N_7491);
nand U7797 (N_7797,N_7115,N_7091);
and U7798 (N_7798,N_7303,N_7086);
or U7799 (N_7799,N_7323,N_7498);
nor U7800 (N_7800,N_7442,N_7061);
nor U7801 (N_7801,N_7405,N_7463);
or U7802 (N_7802,N_7109,N_7350);
nor U7803 (N_7803,N_7173,N_7091);
xnor U7804 (N_7804,N_7414,N_7058);
nor U7805 (N_7805,N_7493,N_7081);
or U7806 (N_7806,N_7334,N_7467);
or U7807 (N_7807,N_7442,N_7294);
or U7808 (N_7808,N_7441,N_7002);
xor U7809 (N_7809,N_7459,N_7271);
and U7810 (N_7810,N_7408,N_7234);
and U7811 (N_7811,N_7316,N_7401);
nand U7812 (N_7812,N_7011,N_7049);
nor U7813 (N_7813,N_7337,N_7306);
nor U7814 (N_7814,N_7028,N_7103);
nor U7815 (N_7815,N_7159,N_7298);
nand U7816 (N_7816,N_7009,N_7189);
or U7817 (N_7817,N_7197,N_7300);
xnor U7818 (N_7818,N_7106,N_7082);
nand U7819 (N_7819,N_7106,N_7028);
xnor U7820 (N_7820,N_7137,N_7301);
and U7821 (N_7821,N_7107,N_7113);
or U7822 (N_7822,N_7390,N_7488);
xor U7823 (N_7823,N_7231,N_7336);
and U7824 (N_7824,N_7065,N_7387);
nand U7825 (N_7825,N_7065,N_7111);
and U7826 (N_7826,N_7059,N_7304);
nand U7827 (N_7827,N_7197,N_7199);
and U7828 (N_7828,N_7115,N_7151);
or U7829 (N_7829,N_7380,N_7385);
or U7830 (N_7830,N_7428,N_7085);
nor U7831 (N_7831,N_7427,N_7324);
xnor U7832 (N_7832,N_7001,N_7497);
xor U7833 (N_7833,N_7187,N_7060);
and U7834 (N_7834,N_7070,N_7221);
nand U7835 (N_7835,N_7474,N_7448);
and U7836 (N_7836,N_7382,N_7372);
nand U7837 (N_7837,N_7494,N_7194);
and U7838 (N_7838,N_7185,N_7100);
nand U7839 (N_7839,N_7036,N_7174);
nor U7840 (N_7840,N_7014,N_7385);
xor U7841 (N_7841,N_7030,N_7298);
nand U7842 (N_7842,N_7278,N_7440);
or U7843 (N_7843,N_7084,N_7425);
and U7844 (N_7844,N_7412,N_7026);
nor U7845 (N_7845,N_7277,N_7153);
xor U7846 (N_7846,N_7499,N_7062);
or U7847 (N_7847,N_7052,N_7389);
nor U7848 (N_7848,N_7122,N_7322);
nor U7849 (N_7849,N_7303,N_7212);
nand U7850 (N_7850,N_7494,N_7155);
nor U7851 (N_7851,N_7342,N_7155);
xnor U7852 (N_7852,N_7011,N_7305);
or U7853 (N_7853,N_7063,N_7138);
and U7854 (N_7854,N_7169,N_7323);
or U7855 (N_7855,N_7116,N_7240);
xor U7856 (N_7856,N_7325,N_7134);
and U7857 (N_7857,N_7351,N_7371);
xnor U7858 (N_7858,N_7277,N_7310);
nand U7859 (N_7859,N_7078,N_7150);
or U7860 (N_7860,N_7300,N_7284);
or U7861 (N_7861,N_7317,N_7232);
xor U7862 (N_7862,N_7284,N_7478);
xor U7863 (N_7863,N_7455,N_7350);
nor U7864 (N_7864,N_7290,N_7064);
nand U7865 (N_7865,N_7315,N_7311);
and U7866 (N_7866,N_7499,N_7355);
nand U7867 (N_7867,N_7471,N_7088);
and U7868 (N_7868,N_7043,N_7476);
and U7869 (N_7869,N_7162,N_7199);
xor U7870 (N_7870,N_7203,N_7330);
nand U7871 (N_7871,N_7012,N_7381);
and U7872 (N_7872,N_7102,N_7251);
and U7873 (N_7873,N_7488,N_7475);
nand U7874 (N_7874,N_7310,N_7289);
and U7875 (N_7875,N_7301,N_7276);
and U7876 (N_7876,N_7365,N_7423);
or U7877 (N_7877,N_7263,N_7004);
nor U7878 (N_7878,N_7356,N_7456);
or U7879 (N_7879,N_7238,N_7432);
nand U7880 (N_7880,N_7189,N_7098);
nand U7881 (N_7881,N_7353,N_7368);
and U7882 (N_7882,N_7343,N_7469);
and U7883 (N_7883,N_7144,N_7075);
nand U7884 (N_7884,N_7378,N_7406);
nand U7885 (N_7885,N_7143,N_7492);
or U7886 (N_7886,N_7369,N_7452);
and U7887 (N_7887,N_7451,N_7283);
nor U7888 (N_7888,N_7249,N_7108);
nand U7889 (N_7889,N_7337,N_7418);
and U7890 (N_7890,N_7096,N_7332);
nor U7891 (N_7891,N_7337,N_7150);
nand U7892 (N_7892,N_7498,N_7043);
nor U7893 (N_7893,N_7262,N_7016);
nor U7894 (N_7894,N_7432,N_7438);
or U7895 (N_7895,N_7416,N_7105);
xor U7896 (N_7896,N_7075,N_7247);
nor U7897 (N_7897,N_7492,N_7332);
xor U7898 (N_7898,N_7353,N_7163);
nand U7899 (N_7899,N_7279,N_7290);
or U7900 (N_7900,N_7108,N_7224);
or U7901 (N_7901,N_7231,N_7068);
and U7902 (N_7902,N_7220,N_7397);
or U7903 (N_7903,N_7199,N_7366);
xnor U7904 (N_7904,N_7077,N_7232);
or U7905 (N_7905,N_7449,N_7060);
and U7906 (N_7906,N_7192,N_7126);
xor U7907 (N_7907,N_7276,N_7131);
xor U7908 (N_7908,N_7224,N_7093);
xor U7909 (N_7909,N_7052,N_7340);
or U7910 (N_7910,N_7200,N_7309);
nor U7911 (N_7911,N_7008,N_7173);
or U7912 (N_7912,N_7113,N_7236);
nor U7913 (N_7913,N_7462,N_7362);
nand U7914 (N_7914,N_7410,N_7423);
xnor U7915 (N_7915,N_7044,N_7051);
and U7916 (N_7916,N_7243,N_7289);
or U7917 (N_7917,N_7333,N_7408);
xnor U7918 (N_7918,N_7429,N_7489);
or U7919 (N_7919,N_7012,N_7190);
and U7920 (N_7920,N_7256,N_7300);
and U7921 (N_7921,N_7471,N_7436);
or U7922 (N_7922,N_7068,N_7466);
nor U7923 (N_7923,N_7470,N_7377);
xnor U7924 (N_7924,N_7312,N_7484);
or U7925 (N_7925,N_7337,N_7048);
xnor U7926 (N_7926,N_7321,N_7294);
xnor U7927 (N_7927,N_7105,N_7089);
or U7928 (N_7928,N_7268,N_7457);
and U7929 (N_7929,N_7346,N_7221);
nor U7930 (N_7930,N_7188,N_7205);
nand U7931 (N_7931,N_7028,N_7499);
xnor U7932 (N_7932,N_7246,N_7302);
or U7933 (N_7933,N_7080,N_7070);
nand U7934 (N_7934,N_7356,N_7369);
or U7935 (N_7935,N_7451,N_7447);
nor U7936 (N_7936,N_7016,N_7395);
nand U7937 (N_7937,N_7174,N_7265);
nor U7938 (N_7938,N_7223,N_7101);
or U7939 (N_7939,N_7265,N_7040);
nor U7940 (N_7940,N_7459,N_7342);
nand U7941 (N_7941,N_7485,N_7055);
nand U7942 (N_7942,N_7228,N_7272);
nand U7943 (N_7943,N_7043,N_7218);
nand U7944 (N_7944,N_7099,N_7158);
nand U7945 (N_7945,N_7258,N_7386);
or U7946 (N_7946,N_7021,N_7300);
nor U7947 (N_7947,N_7456,N_7294);
or U7948 (N_7948,N_7363,N_7338);
or U7949 (N_7949,N_7034,N_7165);
nand U7950 (N_7950,N_7287,N_7443);
or U7951 (N_7951,N_7423,N_7173);
nor U7952 (N_7952,N_7188,N_7304);
nand U7953 (N_7953,N_7183,N_7243);
nand U7954 (N_7954,N_7057,N_7225);
and U7955 (N_7955,N_7018,N_7197);
nand U7956 (N_7956,N_7102,N_7071);
or U7957 (N_7957,N_7126,N_7396);
and U7958 (N_7958,N_7406,N_7131);
xor U7959 (N_7959,N_7045,N_7061);
nand U7960 (N_7960,N_7212,N_7298);
xnor U7961 (N_7961,N_7267,N_7369);
or U7962 (N_7962,N_7023,N_7017);
nor U7963 (N_7963,N_7366,N_7171);
and U7964 (N_7964,N_7031,N_7451);
and U7965 (N_7965,N_7201,N_7297);
xor U7966 (N_7966,N_7161,N_7190);
nor U7967 (N_7967,N_7226,N_7235);
or U7968 (N_7968,N_7393,N_7164);
xnor U7969 (N_7969,N_7276,N_7260);
nand U7970 (N_7970,N_7087,N_7491);
xor U7971 (N_7971,N_7185,N_7373);
and U7972 (N_7972,N_7363,N_7328);
and U7973 (N_7973,N_7242,N_7114);
nor U7974 (N_7974,N_7391,N_7137);
nand U7975 (N_7975,N_7222,N_7327);
nor U7976 (N_7976,N_7212,N_7281);
and U7977 (N_7977,N_7073,N_7231);
or U7978 (N_7978,N_7106,N_7314);
xor U7979 (N_7979,N_7270,N_7127);
and U7980 (N_7980,N_7352,N_7036);
nand U7981 (N_7981,N_7361,N_7163);
nand U7982 (N_7982,N_7416,N_7461);
xor U7983 (N_7983,N_7144,N_7225);
xor U7984 (N_7984,N_7368,N_7262);
nand U7985 (N_7985,N_7051,N_7169);
nand U7986 (N_7986,N_7200,N_7370);
nand U7987 (N_7987,N_7463,N_7196);
and U7988 (N_7988,N_7342,N_7053);
or U7989 (N_7989,N_7104,N_7054);
xor U7990 (N_7990,N_7175,N_7385);
nand U7991 (N_7991,N_7322,N_7463);
xnor U7992 (N_7992,N_7095,N_7088);
nor U7993 (N_7993,N_7488,N_7358);
xnor U7994 (N_7994,N_7149,N_7291);
xor U7995 (N_7995,N_7004,N_7108);
xor U7996 (N_7996,N_7008,N_7496);
and U7997 (N_7997,N_7490,N_7208);
xor U7998 (N_7998,N_7306,N_7054);
or U7999 (N_7999,N_7287,N_7010);
xor U8000 (N_8000,N_7583,N_7576);
and U8001 (N_8001,N_7694,N_7663);
nand U8002 (N_8002,N_7742,N_7879);
nor U8003 (N_8003,N_7633,N_7771);
nor U8004 (N_8004,N_7676,N_7626);
or U8005 (N_8005,N_7957,N_7632);
and U8006 (N_8006,N_7927,N_7672);
or U8007 (N_8007,N_7665,N_7873);
xnor U8008 (N_8008,N_7553,N_7974);
and U8009 (N_8009,N_7648,N_7819);
or U8010 (N_8010,N_7785,N_7714);
xnor U8011 (N_8011,N_7662,N_7745);
xor U8012 (N_8012,N_7791,N_7966);
nor U8013 (N_8013,N_7808,N_7530);
nand U8014 (N_8014,N_7956,N_7853);
nor U8015 (N_8015,N_7989,N_7994);
nor U8016 (N_8016,N_7949,N_7826);
or U8017 (N_8017,N_7992,N_7552);
nand U8018 (N_8018,N_7522,N_7589);
or U8019 (N_8019,N_7737,N_7881);
nand U8020 (N_8020,N_7611,N_7809);
xor U8021 (N_8021,N_7963,N_7794);
nor U8022 (N_8022,N_7834,N_7656);
nand U8023 (N_8023,N_7536,N_7871);
and U8024 (N_8024,N_7897,N_7658);
xnor U8025 (N_8025,N_7977,N_7807);
nor U8026 (N_8026,N_7914,N_7947);
nor U8027 (N_8027,N_7607,N_7603);
xnor U8028 (N_8028,N_7810,N_7524);
nand U8029 (N_8029,N_7752,N_7503);
or U8030 (N_8030,N_7890,N_7911);
nand U8031 (N_8031,N_7624,N_7910);
nand U8032 (N_8032,N_7684,N_7731);
or U8033 (N_8033,N_7972,N_7670);
nand U8034 (N_8034,N_7998,N_7969);
nor U8035 (N_8035,N_7551,N_7644);
xnor U8036 (N_8036,N_7891,N_7582);
xor U8037 (N_8037,N_7820,N_7738);
nand U8038 (N_8038,N_7701,N_7800);
nor U8039 (N_8039,N_7909,N_7850);
nand U8040 (N_8040,N_7874,N_7702);
nand U8041 (N_8041,N_7606,N_7599);
nand U8042 (N_8042,N_7541,N_7840);
xnor U8043 (N_8043,N_7926,N_7619);
and U8044 (N_8044,N_7796,N_7842);
and U8045 (N_8045,N_7801,N_7955);
and U8046 (N_8046,N_7993,N_7678);
or U8047 (N_8047,N_7939,N_7844);
or U8048 (N_8048,N_7691,N_7726);
and U8049 (N_8049,N_7637,N_7650);
nand U8050 (N_8050,N_7841,N_7778);
nand U8051 (N_8051,N_7675,N_7723);
nand U8052 (N_8052,N_7770,N_7520);
and U8053 (N_8053,N_7903,N_7860);
and U8054 (N_8054,N_7715,N_7882);
xor U8055 (N_8055,N_7877,N_7880);
or U8056 (N_8056,N_7932,N_7667);
or U8057 (N_8057,N_7560,N_7629);
xor U8058 (N_8058,N_7788,N_7900);
or U8059 (N_8059,N_7968,N_7704);
nor U8060 (N_8060,N_7557,N_7627);
nor U8061 (N_8061,N_7542,N_7734);
nand U8062 (N_8062,N_7651,N_7588);
xnor U8063 (N_8063,N_7609,N_7511);
and U8064 (N_8064,N_7941,N_7790);
xor U8065 (N_8065,N_7995,N_7744);
or U8066 (N_8066,N_7519,N_7740);
and U8067 (N_8067,N_7793,N_7575);
xnor U8068 (N_8068,N_7766,N_7616);
nor U8069 (N_8069,N_7931,N_7570);
and U8070 (N_8070,N_7686,N_7539);
or U8071 (N_8071,N_7846,N_7677);
xnor U8072 (N_8072,N_7918,N_7933);
nand U8073 (N_8073,N_7913,N_7830);
xnor U8074 (N_8074,N_7755,N_7516);
nand U8075 (N_8075,N_7535,N_7525);
nor U8076 (N_8076,N_7783,N_7905);
xor U8077 (N_8077,N_7655,N_7602);
nor U8078 (N_8078,N_7780,N_7502);
or U8079 (N_8079,N_7849,N_7598);
nor U8080 (N_8080,N_7869,N_7805);
and U8081 (N_8081,N_7513,N_7761);
nor U8082 (N_8082,N_7549,N_7540);
xnor U8083 (N_8083,N_7855,N_7950);
xnor U8084 (N_8084,N_7716,N_7875);
xor U8085 (N_8085,N_7943,N_7856);
nand U8086 (N_8086,N_7827,N_7951);
nor U8087 (N_8087,N_7645,N_7917);
nor U8088 (N_8088,N_7703,N_7854);
and U8089 (N_8089,N_7828,N_7825);
or U8090 (N_8090,N_7837,N_7823);
nor U8091 (N_8091,N_7741,N_7868);
nor U8092 (N_8092,N_7514,N_7639);
and U8093 (N_8093,N_7728,N_7527);
and U8094 (N_8094,N_7548,N_7501);
nor U8095 (N_8095,N_7685,N_7774);
xnor U8096 (N_8096,N_7721,N_7781);
and U8097 (N_8097,N_7625,N_7547);
nor U8098 (N_8098,N_7517,N_7628);
nor U8099 (N_8099,N_7669,N_7690);
and U8100 (N_8100,N_7990,N_7699);
nor U8101 (N_8101,N_7979,N_7858);
nand U8102 (N_8102,N_7554,N_7521);
nor U8103 (N_8103,N_7889,N_7649);
nand U8104 (N_8104,N_7732,N_7848);
or U8105 (N_8105,N_7776,N_7787);
and U8106 (N_8106,N_7505,N_7657);
nand U8107 (N_8107,N_7526,N_7775);
and U8108 (N_8108,N_7580,N_7967);
nand U8109 (N_8109,N_7811,N_7550);
or U8110 (N_8110,N_7509,N_7660);
nand U8111 (N_8111,N_7982,N_7757);
xnor U8112 (N_8112,N_7803,N_7661);
and U8113 (N_8113,N_7824,N_7762);
nor U8114 (N_8114,N_7812,N_7773);
and U8115 (N_8115,N_7946,N_7700);
and U8116 (N_8116,N_7708,N_7935);
nand U8117 (N_8117,N_7952,N_7936);
xor U8118 (N_8118,N_7743,N_7821);
xnor U8119 (N_8119,N_7727,N_7833);
and U8120 (N_8120,N_7971,N_7679);
xnor U8121 (N_8121,N_7797,N_7806);
nand U8122 (N_8122,N_7861,N_7862);
nor U8123 (N_8123,N_7634,N_7887);
or U8124 (N_8124,N_7733,N_7985);
nand U8125 (N_8125,N_7852,N_7707);
nor U8126 (N_8126,N_7567,N_7577);
nand U8127 (N_8127,N_7578,N_7713);
and U8128 (N_8128,N_7872,N_7585);
and U8129 (N_8129,N_7729,N_7747);
nor U8130 (N_8130,N_7748,N_7789);
nor U8131 (N_8131,N_7635,N_7885);
and U8132 (N_8132,N_7753,N_7558);
nand U8133 (N_8133,N_7565,N_7865);
or U8134 (N_8134,N_7839,N_7822);
nand U8135 (N_8135,N_7590,N_7904);
or U8136 (N_8136,N_7813,N_7640);
xor U8137 (N_8137,N_7620,N_7934);
and U8138 (N_8138,N_7984,N_7930);
nor U8139 (N_8139,N_7673,N_7912);
nor U8140 (N_8140,N_7768,N_7646);
and U8141 (N_8141,N_7654,N_7940);
or U8142 (N_8142,N_7643,N_7712);
nand U8143 (N_8143,N_7980,N_7674);
xor U8144 (N_8144,N_7614,N_7717);
or U8145 (N_8145,N_7978,N_7636);
or U8146 (N_8146,N_7693,N_7593);
and U8147 (N_8147,N_7546,N_7622);
nand U8148 (N_8148,N_7581,N_7817);
nor U8149 (N_8149,N_7937,N_7739);
nand U8150 (N_8150,N_7705,N_7597);
nor U8151 (N_8151,N_7604,N_7991);
nor U8152 (N_8152,N_7845,N_7605);
xnor U8153 (N_8153,N_7601,N_7559);
nand U8154 (N_8154,N_7786,N_7760);
nor U8155 (N_8155,N_7749,N_7534);
and U8156 (N_8156,N_7659,N_7544);
nand U8157 (N_8157,N_7682,N_7591);
or U8158 (N_8158,N_7523,N_7864);
nor U8159 (N_8159,N_7894,N_7981);
or U8160 (N_8160,N_7531,N_7960);
nor U8161 (N_8161,N_7987,N_7746);
nand U8162 (N_8162,N_7866,N_7863);
nor U8163 (N_8163,N_7569,N_7698);
nand U8164 (N_8164,N_7916,N_7587);
nor U8165 (N_8165,N_7689,N_7942);
nor U8166 (N_8166,N_7876,N_7504);
nor U8167 (N_8167,N_7986,N_7764);
xor U8168 (N_8168,N_7617,N_7666);
nor U8169 (N_8169,N_7896,N_7512);
nand U8170 (N_8170,N_7621,N_7851);
or U8171 (N_8171,N_7832,N_7722);
nor U8172 (N_8172,N_7901,N_7999);
or U8173 (N_8173,N_7958,N_7928);
xnor U8174 (N_8174,N_7573,N_7938);
or U8175 (N_8175,N_7754,N_7718);
nand U8176 (N_8176,N_7596,N_7532);
nand U8177 (N_8177,N_7953,N_7692);
or U8178 (N_8178,N_7618,N_7906);
and U8179 (N_8179,N_7816,N_7996);
xor U8180 (N_8180,N_7735,N_7507);
and U8181 (N_8181,N_7561,N_7528);
nor U8182 (N_8182,N_7795,N_7829);
or U8183 (N_8183,N_7594,N_7668);
nand U8184 (N_8184,N_7562,N_7867);
or U8185 (N_8185,N_7518,N_7962);
or U8186 (N_8186,N_7959,N_7921);
nand U8187 (N_8187,N_7997,N_7572);
nand U8188 (N_8188,N_7556,N_7653);
xnor U8189 (N_8189,N_7506,N_7870);
nand U8190 (N_8190,N_7647,N_7719);
and U8191 (N_8191,N_7683,N_7652);
xnor U8192 (N_8192,N_7922,N_7608);
xor U8193 (N_8193,N_7584,N_7763);
xnor U8194 (N_8194,N_7835,N_7759);
and U8195 (N_8195,N_7695,N_7564);
nor U8196 (N_8196,N_7681,N_7884);
and U8197 (N_8197,N_7769,N_7784);
and U8198 (N_8198,N_7767,N_7765);
nand U8199 (N_8199,N_7574,N_7924);
nor U8200 (N_8200,N_7595,N_7907);
and U8201 (N_8201,N_7592,N_7915);
nor U8202 (N_8202,N_7892,N_7612);
nor U8203 (N_8203,N_7965,N_7543);
or U8204 (N_8204,N_7970,N_7988);
xor U8205 (N_8205,N_7838,N_7983);
nand U8206 (N_8206,N_7908,N_7706);
or U8207 (N_8207,N_7725,N_7571);
nand U8208 (N_8208,N_7730,N_7533);
xor U8209 (N_8209,N_7680,N_7893);
or U8210 (N_8210,N_7898,N_7586);
nand U8211 (N_8211,N_7782,N_7802);
and U8212 (N_8212,N_7510,N_7919);
and U8213 (N_8213,N_7814,N_7973);
xor U8214 (N_8214,N_7920,N_7724);
xor U8215 (N_8215,N_7709,N_7883);
and U8216 (N_8216,N_7500,N_7756);
xnor U8217 (N_8217,N_7847,N_7697);
xor U8218 (N_8218,N_7751,N_7515);
nand U8219 (N_8219,N_7687,N_7710);
and U8220 (N_8220,N_7537,N_7804);
nand U8221 (N_8221,N_7857,N_7615);
and U8222 (N_8222,N_7799,N_7641);
and U8223 (N_8223,N_7818,N_7579);
nor U8224 (N_8224,N_7945,N_7631);
xor U8225 (N_8225,N_7642,N_7711);
nand U8226 (N_8226,N_7671,N_7613);
and U8227 (N_8227,N_7798,N_7836);
nor U8228 (N_8228,N_7777,N_7944);
nor U8229 (N_8229,N_7568,N_7630);
nor U8230 (N_8230,N_7792,N_7566);
nand U8231 (N_8231,N_7720,N_7664);
and U8232 (N_8232,N_7976,N_7750);
nand U8233 (N_8233,N_7895,N_7954);
or U8234 (N_8234,N_7610,N_7929);
or U8235 (N_8235,N_7888,N_7538);
and U8236 (N_8236,N_7815,N_7925);
nor U8237 (N_8237,N_7555,N_7696);
and U8238 (N_8238,N_7902,N_7878);
or U8239 (N_8239,N_7688,N_7508);
and U8240 (N_8240,N_7623,N_7886);
and U8241 (N_8241,N_7545,N_7758);
xor U8242 (N_8242,N_7923,N_7899);
and U8243 (N_8243,N_7563,N_7948);
nand U8244 (N_8244,N_7600,N_7529);
xor U8245 (N_8245,N_7831,N_7779);
xnor U8246 (N_8246,N_7843,N_7736);
xnor U8247 (N_8247,N_7859,N_7964);
nor U8248 (N_8248,N_7772,N_7638);
nor U8249 (N_8249,N_7975,N_7961);
or U8250 (N_8250,N_7503,N_7865);
nor U8251 (N_8251,N_7580,N_7547);
xnor U8252 (N_8252,N_7761,N_7941);
xnor U8253 (N_8253,N_7857,N_7752);
and U8254 (N_8254,N_7676,N_7999);
or U8255 (N_8255,N_7508,N_7812);
xor U8256 (N_8256,N_7815,N_7678);
and U8257 (N_8257,N_7637,N_7922);
or U8258 (N_8258,N_7602,N_7547);
nand U8259 (N_8259,N_7566,N_7551);
nand U8260 (N_8260,N_7815,N_7539);
or U8261 (N_8261,N_7681,N_7973);
xnor U8262 (N_8262,N_7686,N_7872);
nor U8263 (N_8263,N_7995,N_7646);
xor U8264 (N_8264,N_7790,N_7858);
xnor U8265 (N_8265,N_7869,N_7662);
xor U8266 (N_8266,N_7671,N_7567);
or U8267 (N_8267,N_7560,N_7759);
xnor U8268 (N_8268,N_7643,N_7978);
and U8269 (N_8269,N_7589,N_7621);
xnor U8270 (N_8270,N_7504,N_7794);
xor U8271 (N_8271,N_7538,N_7521);
xnor U8272 (N_8272,N_7801,N_7743);
and U8273 (N_8273,N_7626,N_7872);
and U8274 (N_8274,N_7721,N_7841);
or U8275 (N_8275,N_7605,N_7789);
or U8276 (N_8276,N_7848,N_7987);
or U8277 (N_8277,N_7642,N_7968);
or U8278 (N_8278,N_7691,N_7857);
nand U8279 (N_8279,N_7656,N_7626);
nor U8280 (N_8280,N_7745,N_7800);
nand U8281 (N_8281,N_7570,N_7862);
nand U8282 (N_8282,N_7718,N_7833);
or U8283 (N_8283,N_7839,N_7798);
nor U8284 (N_8284,N_7960,N_7924);
nor U8285 (N_8285,N_7729,N_7727);
or U8286 (N_8286,N_7764,N_7659);
and U8287 (N_8287,N_7818,N_7663);
nand U8288 (N_8288,N_7581,N_7708);
and U8289 (N_8289,N_7905,N_7613);
xnor U8290 (N_8290,N_7624,N_7563);
nand U8291 (N_8291,N_7955,N_7854);
nand U8292 (N_8292,N_7639,N_7951);
nand U8293 (N_8293,N_7985,N_7990);
nand U8294 (N_8294,N_7873,N_7837);
or U8295 (N_8295,N_7646,N_7913);
or U8296 (N_8296,N_7713,N_7570);
and U8297 (N_8297,N_7614,N_7775);
nor U8298 (N_8298,N_7741,N_7748);
nor U8299 (N_8299,N_7632,N_7585);
nor U8300 (N_8300,N_7612,N_7602);
and U8301 (N_8301,N_7833,N_7946);
nor U8302 (N_8302,N_7965,N_7780);
nand U8303 (N_8303,N_7635,N_7848);
xor U8304 (N_8304,N_7698,N_7780);
or U8305 (N_8305,N_7635,N_7750);
nor U8306 (N_8306,N_7951,N_7862);
and U8307 (N_8307,N_7744,N_7689);
and U8308 (N_8308,N_7724,N_7545);
nor U8309 (N_8309,N_7809,N_7749);
and U8310 (N_8310,N_7778,N_7620);
nand U8311 (N_8311,N_7601,N_7981);
and U8312 (N_8312,N_7598,N_7773);
or U8313 (N_8313,N_7641,N_7687);
nand U8314 (N_8314,N_7599,N_7744);
nand U8315 (N_8315,N_7822,N_7523);
or U8316 (N_8316,N_7552,N_7912);
xnor U8317 (N_8317,N_7651,N_7895);
nand U8318 (N_8318,N_7736,N_7859);
and U8319 (N_8319,N_7926,N_7728);
nand U8320 (N_8320,N_7946,N_7777);
or U8321 (N_8321,N_7883,N_7767);
nand U8322 (N_8322,N_7744,N_7985);
or U8323 (N_8323,N_7754,N_7699);
nor U8324 (N_8324,N_7520,N_7884);
or U8325 (N_8325,N_7640,N_7644);
xor U8326 (N_8326,N_7660,N_7724);
nor U8327 (N_8327,N_7735,N_7824);
or U8328 (N_8328,N_7513,N_7928);
or U8329 (N_8329,N_7835,N_7859);
and U8330 (N_8330,N_7510,N_7506);
nor U8331 (N_8331,N_7545,N_7933);
or U8332 (N_8332,N_7744,N_7733);
nor U8333 (N_8333,N_7557,N_7675);
nor U8334 (N_8334,N_7907,N_7622);
nand U8335 (N_8335,N_7744,N_7817);
and U8336 (N_8336,N_7574,N_7701);
nand U8337 (N_8337,N_7970,N_7578);
nor U8338 (N_8338,N_7619,N_7673);
xor U8339 (N_8339,N_7943,N_7642);
nand U8340 (N_8340,N_7738,N_7850);
xnor U8341 (N_8341,N_7747,N_7702);
nor U8342 (N_8342,N_7508,N_7964);
and U8343 (N_8343,N_7607,N_7543);
or U8344 (N_8344,N_7800,N_7620);
xor U8345 (N_8345,N_7612,N_7501);
and U8346 (N_8346,N_7695,N_7556);
and U8347 (N_8347,N_7719,N_7633);
nor U8348 (N_8348,N_7619,N_7694);
nor U8349 (N_8349,N_7988,N_7903);
or U8350 (N_8350,N_7925,N_7890);
or U8351 (N_8351,N_7522,N_7682);
or U8352 (N_8352,N_7916,N_7764);
and U8353 (N_8353,N_7933,N_7800);
nor U8354 (N_8354,N_7801,N_7990);
nand U8355 (N_8355,N_7543,N_7862);
nand U8356 (N_8356,N_7944,N_7823);
or U8357 (N_8357,N_7524,N_7870);
nor U8358 (N_8358,N_7618,N_7627);
and U8359 (N_8359,N_7967,N_7724);
and U8360 (N_8360,N_7826,N_7842);
xor U8361 (N_8361,N_7720,N_7542);
or U8362 (N_8362,N_7524,N_7747);
nand U8363 (N_8363,N_7971,N_7784);
and U8364 (N_8364,N_7840,N_7911);
or U8365 (N_8365,N_7937,N_7985);
or U8366 (N_8366,N_7758,N_7930);
nand U8367 (N_8367,N_7814,N_7812);
and U8368 (N_8368,N_7867,N_7927);
nand U8369 (N_8369,N_7798,N_7604);
nand U8370 (N_8370,N_7703,N_7770);
and U8371 (N_8371,N_7710,N_7822);
xnor U8372 (N_8372,N_7970,N_7915);
nand U8373 (N_8373,N_7688,N_7977);
nand U8374 (N_8374,N_7648,N_7940);
or U8375 (N_8375,N_7946,N_7977);
nor U8376 (N_8376,N_7959,N_7591);
nand U8377 (N_8377,N_7843,N_7764);
or U8378 (N_8378,N_7733,N_7528);
nand U8379 (N_8379,N_7601,N_7752);
nand U8380 (N_8380,N_7639,N_7988);
nand U8381 (N_8381,N_7594,N_7578);
nor U8382 (N_8382,N_7732,N_7871);
nor U8383 (N_8383,N_7993,N_7792);
and U8384 (N_8384,N_7980,N_7943);
nand U8385 (N_8385,N_7685,N_7969);
xor U8386 (N_8386,N_7587,N_7897);
or U8387 (N_8387,N_7559,N_7823);
and U8388 (N_8388,N_7944,N_7746);
nor U8389 (N_8389,N_7994,N_7856);
nand U8390 (N_8390,N_7802,N_7592);
or U8391 (N_8391,N_7836,N_7588);
or U8392 (N_8392,N_7964,N_7691);
xor U8393 (N_8393,N_7757,N_7556);
xnor U8394 (N_8394,N_7871,N_7917);
and U8395 (N_8395,N_7959,N_7517);
nand U8396 (N_8396,N_7718,N_7934);
nand U8397 (N_8397,N_7907,N_7617);
or U8398 (N_8398,N_7942,N_7548);
nor U8399 (N_8399,N_7940,N_7677);
xnor U8400 (N_8400,N_7546,N_7965);
xnor U8401 (N_8401,N_7558,N_7859);
or U8402 (N_8402,N_7680,N_7733);
nor U8403 (N_8403,N_7880,N_7579);
nand U8404 (N_8404,N_7574,N_7664);
or U8405 (N_8405,N_7742,N_7831);
xor U8406 (N_8406,N_7820,N_7687);
nor U8407 (N_8407,N_7701,N_7554);
or U8408 (N_8408,N_7553,N_7826);
and U8409 (N_8409,N_7932,N_7970);
xnor U8410 (N_8410,N_7880,N_7693);
nor U8411 (N_8411,N_7822,N_7583);
and U8412 (N_8412,N_7992,N_7724);
xor U8413 (N_8413,N_7601,N_7646);
nand U8414 (N_8414,N_7918,N_7810);
or U8415 (N_8415,N_7780,N_7804);
nand U8416 (N_8416,N_7993,N_7872);
and U8417 (N_8417,N_7560,N_7795);
nand U8418 (N_8418,N_7632,N_7975);
and U8419 (N_8419,N_7601,N_7633);
or U8420 (N_8420,N_7866,N_7623);
nand U8421 (N_8421,N_7773,N_7635);
and U8422 (N_8422,N_7889,N_7940);
nand U8423 (N_8423,N_7553,N_7919);
and U8424 (N_8424,N_7876,N_7869);
and U8425 (N_8425,N_7749,N_7849);
xnor U8426 (N_8426,N_7613,N_7912);
nand U8427 (N_8427,N_7764,N_7913);
or U8428 (N_8428,N_7785,N_7806);
xor U8429 (N_8429,N_7829,N_7817);
nand U8430 (N_8430,N_7834,N_7846);
or U8431 (N_8431,N_7502,N_7652);
nand U8432 (N_8432,N_7629,N_7769);
xor U8433 (N_8433,N_7654,N_7767);
nor U8434 (N_8434,N_7634,N_7521);
xor U8435 (N_8435,N_7874,N_7955);
nand U8436 (N_8436,N_7945,N_7510);
xnor U8437 (N_8437,N_7783,N_7891);
nand U8438 (N_8438,N_7543,N_7790);
nor U8439 (N_8439,N_7847,N_7796);
or U8440 (N_8440,N_7855,N_7755);
nand U8441 (N_8441,N_7540,N_7505);
nand U8442 (N_8442,N_7548,N_7812);
nor U8443 (N_8443,N_7902,N_7901);
nor U8444 (N_8444,N_7923,N_7904);
or U8445 (N_8445,N_7789,N_7617);
nand U8446 (N_8446,N_7640,N_7591);
and U8447 (N_8447,N_7607,N_7963);
and U8448 (N_8448,N_7777,N_7988);
and U8449 (N_8449,N_7890,N_7927);
nand U8450 (N_8450,N_7612,N_7874);
xnor U8451 (N_8451,N_7635,N_7735);
or U8452 (N_8452,N_7595,N_7603);
xnor U8453 (N_8453,N_7920,N_7698);
nand U8454 (N_8454,N_7966,N_7682);
xnor U8455 (N_8455,N_7600,N_7743);
or U8456 (N_8456,N_7899,N_7760);
and U8457 (N_8457,N_7874,N_7748);
and U8458 (N_8458,N_7763,N_7554);
nand U8459 (N_8459,N_7704,N_7824);
nand U8460 (N_8460,N_7571,N_7791);
xor U8461 (N_8461,N_7869,N_7864);
xnor U8462 (N_8462,N_7884,N_7993);
nand U8463 (N_8463,N_7922,N_7744);
nor U8464 (N_8464,N_7992,N_7921);
nor U8465 (N_8465,N_7569,N_7748);
nor U8466 (N_8466,N_7669,N_7649);
nor U8467 (N_8467,N_7666,N_7857);
nor U8468 (N_8468,N_7817,N_7995);
or U8469 (N_8469,N_7878,N_7749);
nand U8470 (N_8470,N_7769,N_7910);
and U8471 (N_8471,N_7905,N_7994);
nand U8472 (N_8472,N_7694,N_7606);
nand U8473 (N_8473,N_7795,N_7604);
nand U8474 (N_8474,N_7796,N_7617);
nor U8475 (N_8475,N_7921,N_7859);
or U8476 (N_8476,N_7983,N_7848);
nand U8477 (N_8477,N_7754,N_7577);
xor U8478 (N_8478,N_7739,N_7684);
nor U8479 (N_8479,N_7800,N_7959);
or U8480 (N_8480,N_7550,N_7733);
or U8481 (N_8481,N_7542,N_7678);
xnor U8482 (N_8482,N_7676,N_7732);
nand U8483 (N_8483,N_7568,N_7697);
xor U8484 (N_8484,N_7636,N_7761);
and U8485 (N_8485,N_7973,N_7981);
xor U8486 (N_8486,N_7835,N_7973);
or U8487 (N_8487,N_7875,N_7516);
xor U8488 (N_8488,N_7530,N_7952);
xnor U8489 (N_8489,N_7622,N_7592);
nor U8490 (N_8490,N_7779,N_7663);
or U8491 (N_8491,N_7669,N_7548);
nand U8492 (N_8492,N_7979,N_7876);
or U8493 (N_8493,N_7776,N_7889);
nand U8494 (N_8494,N_7515,N_7626);
or U8495 (N_8495,N_7983,N_7893);
xnor U8496 (N_8496,N_7541,N_7876);
or U8497 (N_8497,N_7985,N_7940);
xnor U8498 (N_8498,N_7711,N_7752);
xnor U8499 (N_8499,N_7750,N_7736);
nor U8500 (N_8500,N_8105,N_8153);
or U8501 (N_8501,N_8234,N_8026);
nand U8502 (N_8502,N_8368,N_8027);
and U8503 (N_8503,N_8076,N_8282);
xor U8504 (N_8504,N_8428,N_8132);
or U8505 (N_8505,N_8213,N_8187);
or U8506 (N_8506,N_8041,N_8062);
or U8507 (N_8507,N_8165,N_8366);
xnor U8508 (N_8508,N_8006,N_8379);
nor U8509 (N_8509,N_8162,N_8468);
nand U8510 (N_8510,N_8161,N_8400);
and U8511 (N_8511,N_8416,N_8499);
xnor U8512 (N_8512,N_8114,N_8023);
xor U8513 (N_8513,N_8044,N_8123);
or U8514 (N_8514,N_8049,N_8286);
and U8515 (N_8515,N_8295,N_8382);
nor U8516 (N_8516,N_8140,N_8448);
nor U8517 (N_8517,N_8211,N_8119);
and U8518 (N_8518,N_8219,N_8135);
nor U8519 (N_8519,N_8024,N_8125);
nand U8520 (N_8520,N_8152,N_8306);
or U8521 (N_8521,N_8070,N_8052);
nor U8522 (N_8522,N_8178,N_8430);
xnor U8523 (N_8523,N_8055,N_8293);
xnor U8524 (N_8524,N_8142,N_8484);
nand U8525 (N_8525,N_8439,N_8216);
and U8526 (N_8526,N_8494,N_8012);
nor U8527 (N_8527,N_8248,N_8465);
xnor U8528 (N_8528,N_8003,N_8245);
xnor U8529 (N_8529,N_8361,N_8157);
nand U8530 (N_8530,N_8181,N_8159);
nand U8531 (N_8531,N_8313,N_8230);
nor U8532 (N_8532,N_8015,N_8010);
and U8533 (N_8533,N_8089,N_8004);
nor U8534 (N_8534,N_8288,N_8253);
and U8535 (N_8535,N_8087,N_8461);
or U8536 (N_8536,N_8482,N_8127);
or U8537 (N_8537,N_8281,N_8111);
or U8538 (N_8538,N_8000,N_8297);
xor U8539 (N_8539,N_8378,N_8200);
or U8540 (N_8540,N_8365,N_8303);
nand U8541 (N_8541,N_8183,N_8016);
nand U8542 (N_8542,N_8201,N_8294);
nand U8543 (N_8543,N_8207,N_8324);
nand U8544 (N_8544,N_8374,N_8071);
xnor U8545 (N_8545,N_8490,N_8155);
or U8546 (N_8546,N_8498,N_8054);
xor U8547 (N_8547,N_8192,N_8443);
and U8548 (N_8548,N_8092,N_8255);
and U8549 (N_8549,N_8491,N_8014);
nand U8550 (N_8550,N_8455,N_8040);
xor U8551 (N_8551,N_8496,N_8098);
or U8552 (N_8552,N_8221,N_8462);
and U8553 (N_8553,N_8080,N_8241);
or U8554 (N_8554,N_8097,N_8031);
and U8555 (N_8555,N_8053,N_8384);
xnor U8556 (N_8556,N_8032,N_8130);
nor U8557 (N_8557,N_8316,N_8436);
xnor U8558 (N_8558,N_8321,N_8141);
and U8559 (N_8559,N_8019,N_8225);
xnor U8560 (N_8560,N_8488,N_8419);
and U8561 (N_8561,N_8423,N_8007);
nand U8562 (N_8562,N_8486,N_8243);
and U8563 (N_8563,N_8239,N_8085);
xnor U8564 (N_8564,N_8069,N_8391);
and U8565 (N_8565,N_8137,N_8059);
nand U8566 (N_8566,N_8339,N_8353);
xnor U8567 (N_8567,N_8256,N_8247);
xor U8568 (N_8568,N_8445,N_8300);
nor U8569 (N_8569,N_8199,N_8249);
and U8570 (N_8570,N_8326,N_8463);
nor U8571 (N_8571,N_8106,N_8263);
and U8572 (N_8572,N_8226,N_8264);
nand U8573 (N_8573,N_8072,N_8325);
and U8574 (N_8574,N_8220,N_8291);
or U8575 (N_8575,N_8240,N_8095);
nand U8576 (N_8576,N_8056,N_8341);
or U8577 (N_8577,N_8269,N_8454);
nor U8578 (N_8578,N_8037,N_8437);
or U8579 (N_8579,N_8184,N_8317);
nand U8580 (N_8580,N_8381,N_8146);
and U8581 (N_8581,N_8047,N_8377);
and U8582 (N_8582,N_8458,N_8474);
xor U8583 (N_8583,N_8021,N_8398);
xor U8584 (N_8584,N_8126,N_8081);
xor U8585 (N_8585,N_8174,N_8101);
nand U8586 (N_8586,N_8198,N_8261);
xnor U8587 (N_8587,N_8168,N_8327);
and U8588 (N_8588,N_8193,N_8279);
or U8589 (N_8589,N_8438,N_8479);
nand U8590 (N_8590,N_8328,N_8215);
nand U8591 (N_8591,N_8338,N_8158);
and U8592 (N_8592,N_8359,N_8143);
and U8593 (N_8593,N_8495,N_8138);
and U8594 (N_8594,N_8418,N_8196);
nor U8595 (N_8595,N_8068,N_8077);
nand U8596 (N_8596,N_8229,N_8402);
nand U8597 (N_8597,N_8380,N_8383);
or U8598 (N_8598,N_8011,N_8470);
and U8599 (N_8599,N_8453,N_8287);
xnor U8600 (N_8600,N_8354,N_8242);
nor U8601 (N_8601,N_8449,N_8270);
or U8602 (N_8602,N_8360,N_8265);
nor U8603 (N_8603,N_8170,N_8289);
and U8604 (N_8604,N_8434,N_8322);
or U8605 (N_8605,N_8075,N_8404);
nand U8606 (N_8606,N_8120,N_8441);
nand U8607 (N_8607,N_8048,N_8148);
xor U8608 (N_8608,N_8493,N_8109);
xnor U8609 (N_8609,N_8456,N_8371);
nor U8610 (N_8610,N_8259,N_8393);
xor U8611 (N_8611,N_8426,N_8409);
or U8612 (N_8612,N_8078,N_8172);
nor U8613 (N_8613,N_8442,N_8236);
or U8614 (N_8614,N_8290,N_8369);
nor U8615 (N_8615,N_8411,N_8103);
nand U8616 (N_8616,N_8145,N_8179);
and U8617 (N_8617,N_8376,N_8335);
or U8618 (N_8618,N_8396,N_8357);
and U8619 (N_8619,N_8232,N_8260);
nor U8620 (N_8620,N_8464,N_8009);
nor U8621 (N_8621,N_8312,N_8315);
or U8622 (N_8622,N_8314,N_8110);
xnor U8623 (N_8623,N_8460,N_8233);
xnor U8624 (N_8624,N_8262,N_8244);
xor U8625 (N_8625,N_8214,N_8476);
nor U8626 (N_8626,N_8133,N_8331);
or U8627 (N_8627,N_8005,N_8018);
xnor U8628 (N_8628,N_8086,N_8417);
xnor U8629 (N_8629,N_8307,N_8008);
xnor U8630 (N_8630,N_8188,N_8082);
or U8631 (N_8631,N_8227,N_8191);
or U8632 (N_8632,N_8083,N_8292);
nor U8633 (N_8633,N_8190,N_8115);
or U8634 (N_8634,N_8189,N_8452);
nand U8635 (N_8635,N_8348,N_8283);
xnor U8636 (N_8636,N_8030,N_8074);
or U8637 (N_8637,N_8296,N_8171);
or U8638 (N_8638,N_8131,N_8169);
xor U8639 (N_8639,N_8446,N_8001);
nor U8640 (N_8640,N_8246,N_8223);
xor U8641 (N_8641,N_8309,N_8431);
nor U8642 (N_8642,N_8013,N_8136);
nand U8643 (N_8643,N_8222,N_8299);
nand U8644 (N_8644,N_8096,N_8375);
nor U8645 (N_8645,N_8336,N_8166);
nand U8646 (N_8646,N_8403,N_8094);
and U8647 (N_8647,N_8285,N_8235);
and U8648 (N_8648,N_8002,N_8258);
xor U8649 (N_8649,N_8407,N_8421);
nand U8650 (N_8650,N_8203,N_8124);
xnor U8651 (N_8651,N_8257,N_8319);
or U8652 (N_8652,N_8043,N_8405);
xnor U8653 (N_8653,N_8277,N_8356);
and U8654 (N_8654,N_8301,N_8406);
nand U8655 (N_8655,N_8061,N_8401);
nor U8656 (N_8656,N_8150,N_8063);
nand U8657 (N_8657,N_8035,N_8390);
or U8658 (N_8658,N_8266,N_8029);
and U8659 (N_8659,N_8414,N_8351);
xnor U8660 (N_8660,N_8420,N_8099);
nor U8661 (N_8661,N_8173,N_8058);
and U8662 (N_8662,N_8066,N_8206);
nor U8663 (N_8663,N_8067,N_8149);
nor U8664 (N_8664,N_8394,N_8268);
or U8665 (N_8665,N_8091,N_8182);
nor U8666 (N_8666,N_8251,N_8250);
nor U8667 (N_8667,N_8466,N_8333);
nand U8668 (N_8668,N_8349,N_8386);
nand U8669 (N_8669,N_8489,N_8334);
nand U8670 (N_8670,N_8363,N_8284);
nor U8671 (N_8671,N_8228,N_8433);
or U8672 (N_8672,N_8163,N_8485);
nor U8673 (N_8673,N_8471,N_8042);
xnor U8674 (N_8674,N_8274,N_8395);
and U8675 (N_8675,N_8050,N_8129);
nand U8676 (N_8676,N_8330,N_8435);
or U8677 (N_8677,N_8345,N_8342);
nor U8678 (N_8678,N_8372,N_8039);
and U8679 (N_8679,N_8046,N_8164);
nor U8680 (N_8680,N_8298,N_8065);
nand U8681 (N_8681,N_8057,N_8432);
and U8682 (N_8682,N_8090,N_8202);
or U8683 (N_8683,N_8478,N_8025);
and U8684 (N_8684,N_8177,N_8311);
xor U8685 (N_8685,N_8045,N_8212);
nor U8686 (N_8686,N_8147,N_8459);
and U8687 (N_8687,N_8128,N_8079);
nor U8688 (N_8688,N_8273,N_8424);
or U8689 (N_8689,N_8195,N_8318);
nor U8690 (N_8690,N_8408,N_8472);
nand U8691 (N_8691,N_8477,N_8362);
nor U8692 (N_8692,N_8038,N_8118);
nand U8693 (N_8693,N_8180,N_8276);
nor U8694 (N_8694,N_8122,N_8473);
nand U8695 (N_8695,N_8167,N_8440);
nor U8696 (N_8696,N_8340,N_8160);
xor U8697 (N_8697,N_8217,N_8389);
nor U8698 (N_8698,N_8280,N_8370);
nor U8699 (N_8699,N_8112,N_8194);
and U8700 (N_8700,N_8104,N_8084);
and U8701 (N_8701,N_8469,N_8238);
and U8702 (N_8702,N_8415,N_8352);
nand U8703 (N_8703,N_8305,N_8310);
nand U8704 (N_8704,N_8186,N_8224);
or U8705 (N_8705,N_8254,N_8410);
nand U8706 (N_8706,N_8205,N_8175);
xnor U8707 (N_8707,N_8060,N_8154);
nand U8708 (N_8708,N_8102,N_8185);
xnor U8709 (N_8709,N_8051,N_8427);
xor U8710 (N_8710,N_8036,N_8064);
nand U8711 (N_8711,N_8323,N_8457);
and U8712 (N_8712,N_8022,N_8467);
or U8713 (N_8713,N_8451,N_8108);
nand U8714 (N_8714,N_8367,N_8358);
nor U8715 (N_8715,N_8073,N_8373);
nor U8716 (N_8716,N_8151,N_8208);
and U8717 (N_8717,N_8392,N_8332);
or U8718 (N_8718,N_8344,N_8425);
and U8719 (N_8719,N_8278,N_8034);
and U8720 (N_8720,N_8218,N_8483);
nor U8721 (N_8721,N_8388,N_8204);
and U8722 (N_8722,N_8480,N_8267);
or U8723 (N_8723,N_8346,N_8475);
or U8724 (N_8724,N_8107,N_8093);
and U8725 (N_8725,N_8134,N_8100);
xnor U8726 (N_8726,N_8028,N_8385);
xor U8727 (N_8727,N_8343,N_8116);
or U8728 (N_8728,N_8320,N_8350);
and U8729 (N_8729,N_8329,N_8113);
nand U8730 (N_8730,N_8156,N_8272);
xnor U8731 (N_8731,N_8347,N_8497);
nand U8732 (N_8732,N_8399,N_8231);
and U8733 (N_8733,N_8209,N_8412);
nor U8734 (N_8734,N_8302,N_8088);
xor U8735 (N_8735,N_8117,N_8275);
nand U8736 (N_8736,N_8308,N_8429);
or U8737 (N_8737,N_8355,N_8364);
nor U8738 (N_8738,N_8237,N_8492);
and U8739 (N_8739,N_8033,N_8450);
xnor U8740 (N_8740,N_8176,N_8387);
xor U8741 (N_8741,N_8271,N_8413);
and U8742 (N_8742,N_8121,N_8487);
or U8743 (N_8743,N_8197,N_8252);
nand U8744 (N_8744,N_8422,N_8481);
and U8745 (N_8745,N_8397,N_8020);
nand U8746 (N_8746,N_8017,N_8447);
or U8747 (N_8747,N_8139,N_8144);
nand U8748 (N_8748,N_8444,N_8304);
nor U8749 (N_8749,N_8210,N_8337);
or U8750 (N_8750,N_8380,N_8189);
and U8751 (N_8751,N_8228,N_8410);
or U8752 (N_8752,N_8303,N_8457);
nor U8753 (N_8753,N_8222,N_8302);
nand U8754 (N_8754,N_8059,N_8148);
nand U8755 (N_8755,N_8239,N_8068);
and U8756 (N_8756,N_8256,N_8474);
or U8757 (N_8757,N_8075,N_8178);
or U8758 (N_8758,N_8474,N_8046);
xor U8759 (N_8759,N_8138,N_8365);
nand U8760 (N_8760,N_8194,N_8417);
nor U8761 (N_8761,N_8293,N_8174);
or U8762 (N_8762,N_8351,N_8362);
xnor U8763 (N_8763,N_8189,N_8430);
nand U8764 (N_8764,N_8300,N_8023);
nor U8765 (N_8765,N_8068,N_8292);
nand U8766 (N_8766,N_8198,N_8099);
or U8767 (N_8767,N_8359,N_8091);
xor U8768 (N_8768,N_8195,N_8361);
nand U8769 (N_8769,N_8169,N_8242);
xor U8770 (N_8770,N_8322,N_8185);
nor U8771 (N_8771,N_8424,N_8466);
xor U8772 (N_8772,N_8237,N_8434);
xor U8773 (N_8773,N_8117,N_8066);
nand U8774 (N_8774,N_8252,N_8207);
and U8775 (N_8775,N_8497,N_8250);
nor U8776 (N_8776,N_8317,N_8279);
nand U8777 (N_8777,N_8167,N_8371);
and U8778 (N_8778,N_8079,N_8326);
or U8779 (N_8779,N_8489,N_8010);
nor U8780 (N_8780,N_8111,N_8161);
xor U8781 (N_8781,N_8278,N_8468);
or U8782 (N_8782,N_8041,N_8258);
nor U8783 (N_8783,N_8097,N_8309);
xor U8784 (N_8784,N_8069,N_8194);
nand U8785 (N_8785,N_8184,N_8101);
nor U8786 (N_8786,N_8102,N_8168);
nor U8787 (N_8787,N_8087,N_8476);
nand U8788 (N_8788,N_8386,N_8261);
or U8789 (N_8789,N_8495,N_8128);
nor U8790 (N_8790,N_8444,N_8084);
and U8791 (N_8791,N_8382,N_8004);
or U8792 (N_8792,N_8081,N_8073);
or U8793 (N_8793,N_8441,N_8370);
nor U8794 (N_8794,N_8172,N_8348);
xnor U8795 (N_8795,N_8075,N_8429);
or U8796 (N_8796,N_8307,N_8364);
and U8797 (N_8797,N_8101,N_8485);
and U8798 (N_8798,N_8463,N_8325);
xor U8799 (N_8799,N_8209,N_8139);
nand U8800 (N_8800,N_8154,N_8347);
nand U8801 (N_8801,N_8290,N_8396);
xnor U8802 (N_8802,N_8472,N_8433);
or U8803 (N_8803,N_8280,N_8111);
or U8804 (N_8804,N_8032,N_8111);
nand U8805 (N_8805,N_8038,N_8035);
nor U8806 (N_8806,N_8022,N_8235);
and U8807 (N_8807,N_8306,N_8160);
nand U8808 (N_8808,N_8409,N_8349);
xnor U8809 (N_8809,N_8259,N_8205);
or U8810 (N_8810,N_8463,N_8408);
nand U8811 (N_8811,N_8130,N_8331);
or U8812 (N_8812,N_8098,N_8066);
xor U8813 (N_8813,N_8323,N_8224);
nand U8814 (N_8814,N_8456,N_8271);
nand U8815 (N_8815,N_8189,N_8132);
xor U8816 (N_8816,N_8343,N_8418);
and U8817 (N_8817,N_8055,N_8330);
or U8818 (N_8818,N_8071,N_8009);
xnor U8819 (N_8819,N_8017,N_8081);
nand U8820 (N_8820,N_8014,N_8228);
and U8821 (N_8821,N_8056,N_8064);
and U8822 (N_8822,N_8263,N_8309);
nor U8823 (N_8823,N_8332,N_8350);
nand U8824 (N_8824,N_8471,N_8084);
xor U8825 (N_8825,N_8137,N_8072);
and U8826 (N_8826,N_8332,N_8462);
and U8827 (N_8827,N_8247,N_8248);
nor U8828 (N_8828,N_8254,N_8219);
xnor U8829 (N_8829,N_8170,N_8345);
xnor U8830 (N_8830,N_8076,N_8046);
or U8831 (N_8831,N_8424,N_8461);
nor U8832 (N_8832,N_8105,N_8218);
nand U8833 (N_8833,N_8399,N_8321);
or U8834 (N_8834,N_8035,N_8094);
and U8835 (N_8835,N_8101,N_8206);
or U8836 (N_8836,N_8148,N_8296);
nor U8837 (N_8837,N_8448,N_8337);
xor U8838 (N_8838,N_8240,N_8455);
nand U8839 (N_8839,N_8229,N_8453);
or U8840 (N_8840,N_8094,N_8354);
nor U8841 (N_8841,N_8394,N_8302);
nand U8842 (N_8842,N_8425,N_8491);
nand U8843 (N_8843,N_8372,N_8466);
xor U8844 (N_8844,N_8176,N_8059);
and U8845 (N_8845,N_8114,N_8318);
or U8846 (N_8846,N_8289,N_8100);
and U8847 (N_8847,N_8415,N_8384);
and U8848 (N_8848,N_8299,N_8262);
xnor U8849 (N_8849,N_8174,N_8114);
nand U8850 (N_8850,N_8484,N_8174);
xor U8851 (N_8851,N_8167,N_8419);
nor U8852 (N_8852,N_8466,N_8327);
xor U8853 (N_8853,N_8102,N_8144);
nor U8854 (N_8854,N_8264,N_8187);
nor U8855 (N_8855,N_8256,N_8461);
and U8856 (N_8856,N_8442,N_8133);
and U8857 (N_8857,N_8396,N_8439);
or U8858 (N_8858,N_8268,N_8300);
and U8859 (N_8859,N_8398,N_8337);
and U8860 (N_8860,N_8209,N_8181);
nand U8861 (N_8861,N_8386,N_8437);
and U8862 (N_8862,N_8095,N_8348);
or U8863 (N_8863,N_8149,N_8233);
nor U8864 (N_8864,N_8453,N_8167);
or U8865 (N_8865,N_8074,N_8129);
and U8866 (N_8866,N_8340,N_8408);
and U8867 (N_8867,N_8320,N_8307);
or U8868 (N_8868,N_8449,N_8317);
xor U8869 (N_8869,N_8474,N_8204);
xnor U8870 (N_8870,N_8079,N_8441);
xor U8871 (N_8871,N_8344,N_8177);
nand U8872 (N_8872,N_8195,N_8461);
nand U8873 (N_8873,N_8457,N_8130);
nor U8874 (N_8874,N_8337,N_8088);
nand U8875 (N_8875,N_8029,N_8449);
nand U8876 (N_8876,N_8025,N_8376);
and U8877 (N_8877,N_8213,N_8100);
or U8878 (N_8878,N_8243,N_8459);
or U8879 (N_8879,N_8427,N_8183);
or U8880 (N_8880,N_8226,N_8038);
xnor U8881 (N_8881,N_8099,N_8167);
nand U8882 (N_8882,N_8102,N_8405);
nor U8883 (N_8883,N_8074,N_8149);
xnor U8884 (N_8884,N_8379,N_8317);
and U8885 (N_8885,N_8026,N_8322);
or U8886 (N_8886,N_8300,N_8470);
nand U8887 (N_8887,N_8006,N_8120);
and U8888 (N_8888,N_8478,N_8172);
or U8889 (N_8889,N_8258,N_8470);
or U8890 (N_8890,N_8258,N_8379);
or U8891 (N_8891,N_8445,N_8025);
xnor U8892 (N_8892,N_8039,N_8095);
or U8893 (N_8893,N_8344,N_8097);
nor U8894 (N_8894,N_8127,N_8028);
or U8895 (N_8895,N_8050,N_8094);
nor U8896 (N_8896,N_8013,N_8018);
nor U8897 (N_8897,N_8071,N_8237);
nor U8898 (N_8898,N_8470,N_8093);
or U8899 (N_8899,N_8300,N_8441);
xnor U8900 (N_8900,N_8022,N_8051);
xnor U8901 (N_8901,N_8475,N_8079);
nand U8902 (N_8902,N_8228,N_8486);
nor U8903 (N_8903,N_8383,N_8492);
xnor U8904 (N_8904,N_8002,N_8134);
and U8905 (N_8905,N_8333,N_8199);
nand U8906 (N_8906,N_8398,N_8284);
xor U8907 (N_8907,N_8399,N_8039);
nor U8908 (N_8908,N_8242,N_8257);
and U8909 (N_8909,N_8023,N_8069);
xnor U8910 (N_8910,N_8079,N_8435);
or U8911 (N_8911,N_8210,N_8471);
nor U8912 (N_8912,N_8160,N_8122);
nand U8913 (N_8913,N_8367,N_8487);
and U8914 (N_8914,N_8272,N_8294);
nor U8915 (N_8915,N_8239,N_8379);
nor U8916 (N_8916,N_8042,N_8393);
and U8917 (N_8917,N_8101,N_8294);
xor U8918 (N_8918,N_8280,N_8387);
or U8919 (N_8919,N_8037,N_8179);
xor U8920 (N_8920,N_8444,N_8425);
and U8921 (N_8921,N_8199,N_8019);
xor U8922 (N_8922,N_8324,N_8268);
nand U8923 (N_8923,N_8130,N_8263);
nand U8924 (N_8924,N_8435,N_8201);
and U8925 (N_8925,N_8290,N_8193);
or U8926 (N_8926,N_8280,N_8134);
and U8927 (N_8927,N_8330,N_8472);
nand U8928 (N_8928,N_8343,N_8480);
and U8929 (N_8929,N_8322,N_8337);
or U8930 (N_8930,N_8142,N_8144);
xor U8931 (N_8931,N_8399,N_8487);
or U8932 (N_8932,N_8071,N_8423);
xnor U8933 (N_8933,N_8028,N_8012);
nor U8934 (N_8934,N_8240,N_8044);
and U8935 (N_8935,N_8132,N_8328);
xnor U8936 (N_8936,N_8298,N_8393);
nand U8937 (N_8937,N_8489,N_8416);
xor U8938 (N_8938,N_8104,N_8329);
nor U8939 (N_8939,N_8257,N_8326);
nand U8940 (N_8940,N_8417,N_8483);
and U8941 (N_8941,N_8167,N_8484);
xor U8942 (N_8942,N_8293,N_8208);
or U8943 (N_8943,N_8024,N_8101);
xor U8944 (N_8944,N_8288,N_8424);
or U8945 (N_8945,N_8353,N_8395);
and U8946 (N_8946,N_8187,N_8163);
or U8947 (N_8947,N_8052,N_8102);
xnor U8948 (N_8948,N_8274,N_8087);
xor U8949 (N_8949,N_8358,N_8122);
nor U8950 (N_8950,N_8410,N_8156);
and U8951 (N_8951,N_8224,N_8412);
or U8952 (N_8952,N_8012,N_8423);
or U8953 (N_8953,N_8246,N_8310);
or U8954 (N_8954,N_8168,N_8045);
nand U8955 (N_8955,N_8254,N_8275);
nand U8956 (N_8956,N_8081,N_8067);
nand U8957 (N_8957,N_8358,N_8267);
and U8958 (N_8958,N_8156,N_8159);
or U8959 (N_8959,N_8488,N_8271);
or U8960 (N_8960,N_8183,N_8279);
nor U8961 (N_8961,N_8147,N_8439);
nand U8962 (N_8962,N_8401,N_8251);
nor U8963 (N_8963,N_8141,N_8412);
or U8964 (N_8964,N_8476,N_8452);
nand U8965 (N_8965,N_8014,N_8470);
xor U8966 (N_8966,N_8018,N_8490);
nand U8967 (N_8967,N_8078,N_8349);
nand U8968 (N_8968,N_8181,N_8352);
nor U8969 (N_8969,N_8058,N_8305);
nor U8970 (N_8970,N_8380,N_8384);
nand U8971 (N_8971,N_8420,N_8211);
nand U8972 (N_8972,N_8143,N_8032);
xor U8973 (N_8973,N_8365,N_8387);
nor U8974 (N_8974,N_8190,N_8475);
and U8975 (N_8975,N_8304,N_8293);
or U8976 (N_8976,N_8478,N_8369);
nor U8977 (N_8977,N_8328,N_8038);
nand U8978 (N_8978,N_8452,N_8195);
nor U8979 (N_8979,N_8062,N_8032);
nand U8980 (N_8980,N_8297,N_8046);
or U8981 (N_8981,N_8302,N_8165);
or U8982 (N_8982,N_8285,N_8269);
or U8983 (N_8983,N_8441,N_8065);
nor U8984 (N_8984,N_8046,N_8053);
nand U8985 (N_8985,N_8377,N_8255);
nand U8986 (N_8986,N_8382,N_8261);
nor U8987 (N_8987,N_8291,N_8354);
xor U8988 (N_8988,N_8213,N_8323);
nor U8989 (N_8989,N_8205,N_8264);
or U8990 (N_8990,N_8105,N_8247);
and U8991 (N_8991,N_8071,N_8263);
nor U8992 (N_8992,N_8022,N_8307);
and U8993 (N_8993,N_8418,N_8358);
and U8994 (N_8994,N_8399,N_8377);
nor U8995 (N_8995,N_8494,N_8401);
nand U8996 (N_8996,N_8138,N_8369);
xor U8997 (N_8997,N_8228,N_8425);
or U8998 (N_8998,N_8200,N_8239);
or U8999 (N_8999,N_8001,N_8044);
xnor U9000 (N_9000,N_8583,N_8733);
nand U9001 (N_9001,N_8831,N_8557);
nor U9002 (N_9002,N_8775,N_8757);
nor U9003 (N_9003,N_8967,N_8734);
or U9004 (N_9004,N_8839,N_8944);
nor U9005 (N_9005,N_8568,N_8903);
nand U9006 (N_9006,N_8842,N_8600);
or U9007 (N_9007,N_8559,N_8803);
xnor U9008 (N_9008,N_8740,N_8615);
and U9009 (N_9009,N_8784,N_8597);
nand U9010 (N_9010,N_8828,N_8850);
or U9011 (N_9011,N_8922,N_8991);
or U9012 (N_9012,N_8694,N_8960);
xnor U9013 (N_9013,N_8943,N_8780);
or U9014 (N_9014,N_8779,N_8676);
or U9015 (N_9015,N_8560,N_8681);
nand U9016 (N_9016,N_8946,N_8720);
and U9017 (N_9017,N_8987,N_8719);
or U9018 (N_9018,N_8692,N_8723);
nand U9019 (N_9019,N_8999,N_8730);
or U9020 (N_9020,N_8728,N_8710);
nor U9021 (N_9021,N_8675,N_8966);
nand U9022 (N_9022,N_8797,N_8558);
nand U9023 (N_9023,N_8622,N_8766);
xor U9024 (N_9024,N_8737,N_8501);
or U9025 (N_9025,N_8826,N_8636);
nor U9026 (N_9026,N_8616,N_8974);
nor U9027 (N_9027,N_8591,N_8990);
xnor U9028 (N_9028,N_8652,N_8918);
and U9029 (N_9029,N_8908,N_8588);
xor U9030 (N_9030,N_8644,N_8874);
nor U9031 (N_9031,N_8919,N_8716);
and U9032 (N_9032,N_8537,N_8892);
nor U9033 (N_9033,N_8662,N_8672);
xnor U9034 (N_9034,N_8935,N_8660);
and U9035 (N_9035,N_8785,N_8579);
nor U9036 (N_9036,N_8576,N_8542);
and U9037 (N_9037,N_8637,N_8880);
nor U9038 (N_9038,N_8679,N_8882);
and U9039 (N_9039,N_8952,N_8947);
xor U9040 (N_9040,N_8760,N_8798);
nor U9041 (N_9041,N_8848,N_8836);
xor U9042 (N_9042,N_8879,N_8586);
xnor U9043 (N_9043,N_8742,N_8701);
and U9044 (N_9044,N_8659,N_8735);
xor U9045 (N_9045,N_8691,N_8685);
nand U9046 (N_9046,N_8608,N_8902);
nand U9047 (N_9047,N_8645,N_8631);
xnor U9048 (N_9048,N_8771,N_8623);
or U9049 (N_9049,N_8863,N_8657);
or U9050 (N_9050,N_8578,N_8746);
and U9051 (N_9051,N_8988,N_8704);
or U9052 (N_9052,N_8849,N_8641);
or U9053 (N_9053,N_8890,N_8577);
nand U9054 (N_9054,N_8605,N_8614);
and U9055 (N_9055,N_8612,N_8810);
nor U9056 (N_9056,N_8706,N_8787);
and U9057 (N_9057,N_8975,N_8599);
nor U9058 (N_9058,N_8811,N_8971);
xnor U9059 (N_9059,N_8711,N_8629);
xor U9060 (N_9060,N_8653,N_8920);
xor U9061 (N_9061,N_8620,N_8671);
or U9062 (N_9062,N_8980,N_8756);
nor U9063 (N_9063,N_8518,N_8893);
nand U9064 (N_9064,N_8511,N_8926);
and U9065 (N_9065,N_8650,N_8862);
nor U9066 (N_9066,N_8630,N_8950);
and U9067 (N_9067,N_8869,N_8546);
or U9068 (N_9068,N_8707,N_8833);
and U9069 (N_9069,N_8914,N_8989);
xnor U9070 (N_9070,N_8555,N_8921);
xnor U9071 (N_9071,N_8635,N_8886);
and U9072 (N_9072,N_8697,N_8736);
and U9073 (N_9073,N_8743,N_8674);
nand U9074 (N_9074,N_8695,N_8817);
nor U9075 (N_9075,N_8522,N_8993);
xor U9076 (N_9076,N_8529,N_8617);
or U9077 (N_9077,N_8729,N_8801);
nand U9078 (N_9078,N_8953,N_8643);
and U9079 (N_9079,N_8673,N_8596);
nand U9080 (N_9080,N_8891,N_8503);
nor U9081 (N_9081,N_8783,N_8954);
or U9082 (N_9082,N_8561,N_8544);
or U9083 (N_9083,N_8940,N_8851);
xor U9084 (N_9084,N_8872,N_8603);
xnor U9085 (N_9085,N_8765,N_8881);
nor U9086 (N_9086,N_8773,N_8747);
and U9087 (N_9087,N_8654,N_8913);
and U9088 (N_9088,N_8687,N_8633);
nand U9089 (N_9089,N_8651,N_8992);
nor U9090 (N_9090,N_8776,N_8648);
or U9091 (N_9091,N_8661,N_8900);
nor U9092 (N_9092,N_8843,N_8649);
xnor U9093 (N_9093,N_8984,N_8572);
xor U9094 (N_9094,N_8976,N_8517);
and U9095 (N_9095,N_8889,N_8748);
or U9096 (N_9096,N_8625,N_8689);
or U9097 (N_9097,N_8684,N_8670);
xnor U9098 (N_9098,N_8875,N_8794);
nand U9099 (N_9099,N_8937,N_8871);
or U9100 (N_9100,N_8806,N_8959);
nand U9101 (N_9101,N_8864,N_8721);
or U9102 (N_9102,N_8915,N_8807);
xor U9103 (N_9103,N_8996,N_8972);
nand U9104 (N_9104,N_8702,N_8824);
nand U9105 (N_9105,N_8956,N_8854);
nor U9106 (N_9106,N_8613,N_8516);
nand U9107 (N_9107,N_8865,N_8580);
nand U9108 (N_9108,N_8796,N_8745);
or U9109 (N_9109,N_8678,N_8752);
xnor U9110 (N_9110,N_8994,N_8667);
nand U9111 (N_9111,N_8538,N_8853);
or U9112 (N_9112,N_8632,N_8741);
nand U9113 (N_9113,N_8858,N_8677);
nor U9114 (N_9114,N_8938,N_8834);
xnor U9115 (N_9115,N_8977,N_8963);
xnor U9116 (N_9116,N_8770,N_8878);
nand U9117 (N_9117,N_8604,N_8852);
or U9118 (N_9118,N_8714,N_8540);
nand U9119 (N_9119,N_8820,N_8951);
nand U9120 (N_9120,N_8793,N_8762);
nand U9121 (N_9121,N_8751,N_8717);
or U9122 (N_9122,N_8981,N_8593);
nor U9123 (N_9123,N_8936,N_8524);
or U9124 (N_9124,N_8727,N_8982);
and U9125 (N_9125,N_8825,N_8961);
nand U9126 (N_9126,N_8957,N_8822);
xnor U9127 (N_9127,N_8777,N_8931);
or U9128 (N_9128,N_8545,N_8722);
xor U9129 (N_9129,N_8724,N_8680);
and U9130 (N_9130,N_8927,N_8782);
or U9131 (N_9131,N_8590,N_8581);
xnor U9132 (N_9132,N_8816,N_8911);
xnor U9133 (N_9133,N_8898,N_8536);
or U9134 (N_9134,N_8505,N_8642);
and U9135 (N_9135,N_8844,N_8640);
xnor U9136 (N_9136,N_8838,N_8543);
nor U9137 (N_9137,N_8755,N_8929);
nand U9138 (N_9138,N_8827,N_8781);
and U9139 (N_9139,N_8768,N_8532);
nand U9140 (N_9140,N_8666,N_8986);
xnor U9141 (N_9141,N_8949,N_8815);
and U9142 (N_9142,N_8514,N_8837);
or U9143 (N_9143,N_8708,N_8574);
nand U9144 (N_9144,N_8792,N_8703);
nor U9145 (N_9145,N_8700,N_8983);
nor U9146 (N_9146,N_8932,N_8563);
or U9147 (N_9147,N_8821,N_8928);
nor U9148 (N_9148,N_8606,N_8690);
nand U9149 (N_9149,N_8513,N_8609);
and U9150 (N_9150,N_8669,N_8763);
or U9151 (N_9151,N_8634,N_8598);
xnor U9152 (N_9152,N_8530,N_8772);
xnor U9153 (N_9153,N_8589,N_8948);
or U9154 (N_9154,N_8571,N_8539);
nor U9155 (N_9155,N_8904,N_8958);
nand U9156 (N_9156,N_8533,N_8830);
nand U9157 (N_9157,N_8841,N_8705);
or U9158 (N_9158,N_8916,N_8582);
xor U9159 (N_9159,N_8658,N_8739);
xor U9160 (N_9160,N_8925,N_8767);
or U9161 (N_9161,N_8769,N_8726);
or U9162 (N_9162,N_8738,N_8550);
xor U9163 (N_9163,N_8970,N_8535);
and U9164 (N_9164,N_8715,N_8646);
nor U9165 (N_9165,N_8698,N_8638);
xor U9166 (N_9166,N_8786,N_8894);
or U9167 (N_9167,N_8527,N_8512);
and U9168 (N_9168,N_8528,N_8713);
nand U9169 (N_9169,N_8761,N_8699);
and U9170 (N_9170,N_8800,N_8541);
xor U9171 (N_9171,N_8523,N_8978);
or U9172 (N_9172,N_8507,N_8997);
and U9173 (N_9173,N_8602,N_8812);
and U9174 (N_9174,N_8998,N_8778);
nand U9175 (N_9175,N_8930,N_8664);
xor U9176 (N_9176,N_8718,N_8709);
or U9177 (N_9177,N_8870,N_8732);
nand U9178 (N_9178,N_8868,N_8791);
or U9179 (N_9179,N_8744,N_8508);
or U9180 (N_9180,N_8519,N_8554);
xor U9181 (N_9181,N_8509,N_8683);
xor U9182 (N_9182,N_8968,N_8909);
or U9183 (N_9183,N_8570,N_8587);
nand U9184 (N_9184,N_8855,N_8573);
nor U9185 (N_9185,N_8985,N_8548);
xor U9186 (N_9186,N_8515,N_8655);
xor U9187 (N_9187,N_8877,N_8525);
nor U9188 (N_9188,N_8910,N_8534);
nand U9189 (N_9189,N_8823,N_8567);
nand U9190 (N_9190,N_8790,N_8885);
nor U9191 (N_9191,N_8696,N_8663);
nor U9192 (N_9192,N_8813,N_8955);
nand U9193 (N_9193,N_8564,N_8887);
and U9194 (N_9194,N_8725,N_8753);
or U9195 (N_9195,N_8934,N_8814);
and U9196 (N_9196,N_8500,N_8627);
or U9197 (N_9197,N_8788,N_8750);
or U9198 (N_9198,N_8686,N_8607);
xnor U9199 (N_9199,N_8795,N_8502);
nand U9200 (N_9200,N_8585,N_8553);
and U9201 (N_9201,N_8912,N_8688);
xnor U9202 (N_9202,N_8504,N_8565);
xor U9203 (N_9203,N_8626,N_8526);
or U9204 (N_9204,N_8506,N_8595);
nand U9205 (N_9205,N_8876,N_8924);
or U9206 (N_9206,N_8835,N_8712);
nor U9207 (N_9207,N_8860,N_8556);
and U9208 (N_9208,N_8846,N_8520);
nor U9209 (N_9209,N_8758,N_8531);
and U9210 (N_9210,N_8799,N_8939);
nand U9211 (N_9211,N_8867,N_8547);
and U9212 (N_9212,N_8866,N_8805);
nor U9213 (N_9213,N_8624,N_8668);
or U9214 (N_9214,N_8964,N_8857);
and U9215 (N_9215,N_8521,N_8619);
nor U9216 (N_9216,N_8618,N_8552);
xor U9217 (N_9217,N_8639,N_8941);
xnor U9218 (N_9218,N_8884,N_8789);
and U9219 (N_9219,N_8933,N_8901);
xnor U9220 (N_9220,N_8979,N_8856);
nor U9221 (N_9221,N_8883,N_8923);
nor U9222 (N_9222,N_8895,N_8549);
nand U9223 (N_9223,N_8621,N_8899);
or U9224 (N_9224,N_8601,N_8917);
or U9225 (N_9225,N_8962,N_8973);
nand U9226 (N_9226,N_8682,N_8819);
nand U9227 (N_9227,N_8861,N_8965);
nor U9228 (N_9228,N_8610,N_8905);
nor U9229 (N_9229,N_8566,N_8628);
xor U9230 (N_9230,N_8551,N_8592);
nor U9231 (N_9231,N_8859,N_8907);
nor U9232 (N_9232,N_8845,N_8665);
and U9233 (N_9233,N_8840,N_8594);
or U9234 (N_9234,N_8829,N_8764);
nand U9235 (N_9235,N_8569,N_8818);
or U9236 (N_9236,N_8693,N_8969);
xnor U9237 (N_9237,N_8774,N_8802);
and U9238 (N_9238,N_8945,N_8896);
and U9239 (N_9239,N_8584,N_8656);
xnor U9240 (N_9240,N_8611,N_8759);
and U9241 (N_9241,N_8575,N_8562);
or U9242 (N_9242,N_8804,N_8809);
nand U9243 (N_9243,N_8510,N_8873);
and U9244 (N_9244,N_8754,N_8995);
xor U9245 (N_9245,N_8808,N_8647);
or U9246 (N_9246,N_8906,N_8749);
or U9247 (N_9247,N_8888,N_8832);
or U9248 (N_9248,N_8897,N_8731);
xnor U9249 (N_9249,N_8942,N_8847);
and U9250 (N_9250,N_8833,N_8554);
xor U9251 (N_9251,N_8531,N_8761);
or U9252 (N_9252,N_8630,N_8617);
or U9253 (N_9253,N_8916,N_8940);
nor U9254 (N_9254,N_8903,N_8961);
and U9255 (N_9255,N_8768,N_8727);
nor U9256 (N_9256,N_8515,N_8567);
xor U9257 (N_9257,N_8664,N_8825);
xnor U9258 (N_9258,N_8768,N_8746);
or U9259 (N_9259,N_8902,N_8758);
nand U9260 (N_9260,N_8931,N_8885);
nand U9261 (N_9261,N_8782,N_8630);
xnor U9262 (N_9262,N_8943,N_8787);
or U9263 (N_9263,N_8923,N_8796);
and U9264 (N_9264,N_8560,N_8580);
or U9265 (N_9265,N_8952,N_8638);
xnor U9266 (N_9266,N_8784,N_8904);
nand U9267 (N_9267,N_8954,N_8771);
nor U9268 (N_9268,N_8593,N_8708);
nor U9269 (N_9269,N_8708,N_8553);
nor U9270 (N_9270,N_8794,N_8726);
and U9271 (N_9271,N_8557,N_8998);
nand U9272 (N_9272,N_8550,N_8675);
nor U9273 (N_9273,N_8892,N_8741);
or U9274 (N_9274,N_8734,N_8864);
xnor U9275 (N_9275,N_8800,N_8850);
nand U9276 (N_9276,N_8931,N_8784);
nand U9277 (N_9277,N_8582,N_8896);
or U9278 (N_9278,N_8592,N_8680);
nor U9279 (N_9279,N_8983,N_8812);
nand U9280 (N_9280,N_8824,N_8568);
nand U9281 (N_9281,N_8839,N_8840);
nor U9282 (N_9282,N_8713,N_8562);
nor U9283 (N_9283,N_8556,N_8695);
xor U9284 (N_9284,N_8886,N_8916);
and U9285 (N_9285,N_8789,N_8708);
and U9286 (N_9286,N_8602,N_8912);
or U9287 (N_9287,N_8576,N_8636);
and U9288 (N_9288,N_8891,N_8920);
or U9289 (N_9289,N_8740,N_8634);
nor U9290 (N_9290,N_8699,N_8720);
xor U9291 (N_9291,N_8810,N_8761);
or U9292 (N_9292,N_8760,N_8776);
xor U9293 (N_9293,N_8934,N_8893);
nor U9294 (N_9294,N_8941,N_8816);
or U9295 (N_9295,N_8571,N_8973);
or U9296 (N_9296,N_8554,N_8569);
nand U9297 (N_9297,N_8663,N_8523);
and U9298 (N_9298,N_8772,N_8613);
or U9299 (N_9299,N_8960,N_8863);
xnor U9300 (N_9300,N_8684,N_8699);
and U9301 (N_9301,N_8661,N_8906);
nor U9302 (N_9302,N_8799,N_8738);
or U9303 (N_9303,N_8879,N_8551);
nor U9304 (N_9304,N_8662,N_8737);
or U9305 (N_9305,N_8661,N_8665);
and U9306 (N_9306,N_8959,N_8977);
or U9307 (N_9307,N_8619,N_8867);
or U9308 (N_9308,N_8758,N_8567);
nand U9309 (N_9309,N_8723,N_8725);
or U9310 (N_9310,N_8562,N_8832);
xor U9311 (N_9311,N_8606,N_8862);
or U9312 (N_9312,N_8875,N_8649);
and U9313 (N_9313,N_8985,N_8783);
nor U9314 (N_9314,N_8572,N_8548);
nand U9315 (N_9315,N_8814,N_8921);
or U9316 (N_9316,N_8603,N_8660);
or U9317 (N_9317,N_8708,N_8814);
nand U9318 (N_9318,N_8590,N_8741);
nand U9319 (N_9319,N_8763,N_8921);
nor U9320 (N_9320,N_8820,N_8878);
or U9321 (N_9321,N_8539,N_8725);
nor U9322 (N_9322,N_8574,N_8846);
and U9323 (N_9323,N_8978,N_8858);
xor U9324 (N_9324,N_8641,N_8996);
xor U9325 (N_9325,N_8688,N_8606);
xor U9326 (N_9326,N_8821,N_8743);
xor U9327 (N_9327,N_8631,N_8828);
and U9328 (N_9328,N_8555,N_8536);
nor U9329 (N_9329,N_8540,N_8657);
xor U9330 (N_9330,N_8592,N_8772);
nand U9331 (N_9331,N_8798,N_8842);
xor U9332 (N_9332,N_8781,N_8968);
nor U9333 (N_9333,N_8674,N_8834);
nand U9334 (N_9334,N_8736,N_8677);
nor U9335 (N_9335,N_8516,N_8509);
nor U9336 (N_9336,N_8735,N_8740);
and U9337 (N_9337,N_8894,N_8762);
nor U9338 (N_9338,N_8725,N_8834);
and U9339 (N_9339,N_8860,N_8767);
nand U9340 (N_9340,N_8984,N_8793);
xnor U9341 (N_9341,N_8986,N_8931);
nand U9342 (N_9342,N_8516,N_8756);
or U9343 (N_9343,N_8938,N_8795);
xnor U9344 (N_9344,N_8861,N_8529);
and U9345 (N_9345,N_8574,N_8679);
nand U9346 (N_9346,N_8847,N_8966);
nand U9347 (N_9347,N_8960,N_8670);
and U9348 (N_9348,N_8821,N_8882);
and U9349 (N_9349,N_8753,N_8647);
nor U9350 (N_9350,N_8772,N_8926);
and U9351 (N_9351,N_8753,N_8576);
and U9352 (N_9352,N_8515,N_8966);
or U9353 (N_9353,N_8915,N_8545);
nand U9354 (N_9354,N_8773,N_8825);
xnor U9355 (N_9355,N_8698,N_8711);
xor U9356 (N_9356,N_8647,N_8939);
nor U9357 (N_9357,N_8838,N_8756);
xnor U9358 (N_9358,N_8781,N_8852);
xnor U9359 (N_9359,N_8627,N_8711);
and U9360 (N_9360,N_8745,N_8600);
nor U9361 (N_9361,N_8784,N_8712);
and U9362 (N_9362,N_8810,N_8584);
nand U9363 (N_9363,N_8628,N_8991);
nor U9364 (N_9364,N_8888,N_8790);
nand U9365 (N_9365,N_8916,N_8806);
or U9366 (N_9366,N_8730,N_8684);
or U9367 (N_9367,N_8742,N_8757);
nand U9368 (N_9368,N_8619,N_8952);
nor U9369 (N_9369,N_8567,N_8775);
xor U9370 (N_9370,N_8729,N_8677);
xor U9371 (N_9371,N_8929,N_8705);
nand U9372 (N_9372,N_8893,N_8694);
or U9373 (N_9373,N_8878,N_8881);
or U9374 (N_9374,N_8738,N_8542);
nor U9375 (N_9375,N_8848,N_8837);
and U9376 (N_9376,N_8927,N_8759);
xnor U9377 (N_9377,N_8921,N_8502);
nand U9378 (N_9378,N_8912,N_8603);
nor U9379 (N_9379,N_8763,N_8751);
nor U9380 (N_9380,N_8914,N_8739);
xor U9381 (N_9381,N_8671,N_8673);
or U9382 (N_9382,N_8716,N_8915);
or U9383 (N_9383,N_8602,N_8584);
nor U9384 (N_9384,N_8888,N_8723);
and U9385 (N_9385,N_8953,N_8522);
xor U9386 (N_9386,N_8670,N_8823);
or U9387 (N_9387,N_8848,N_8656);
nand U9388 (N_9388,N_8514,N_8892);
or U9389 (N_9389,N_8629,N_8521);
xnor U9390 (N_9390,N_8520,N_8818);
and U9391 (N_9391,N_8802,N_8792);
or U9392 (N_9392,N_8650,N_8703);
nand U9393 (N_9393,N_8569,N_8587);
nand U9394 (N_9394,N_8954,N_8647);
or U9395 (N_9395,N_8594,N_8552);
or U9396 (N_9396,N_8611,N_8528);
xnor U9397 (N_9397,N_8922,N_8502);
nor U9398 (N_9398,N_8763,N_8526);
or U9399 (N_9399,N_8658,N_8902);
nand U9400 (N_9400,N_8878,N_8969);
or U9401 (N_9401,N_8559,N_8853);
xor U9402 (N_9402,N_8961,N_8863);
nor U9403 (N_9403,N_8646,N_8711);
nor U9404 (N_9404,N_8717,N_8814);
and U9405 (N_9405,N_8580,N_8783);
or U9406 (N_9406,N_8776,N_8990);
nand U9407 (N_9407,N_8679,N_8855);
nor U9408 (N_9408,N_8712,N_8606);
and U9409 (N_9409,N_8570,N_8512);
and U9410 (N_9410,N_8860,N_8836);
or U9411 (N_9411,N_8548,N_8797);
xnor U9412 (N_9412,N_8733,N_8943);
xnor U9413 (N_9413,N_8629,N_8736);
nor U9414 (N_9414,N_8854,N_8744);
xor U9415 (N_9415,N_8862,N_8574);
and U9416 (N_9416,N_8594,N_8660);
nand U9417 (N_9417,N_8670,N_8884);
nor U9418 (N_9418,N_8912,N_8906);
nor U9419 (N_9419,N_8665,N_8801);
nand U9420 (N_9420,N_8581,N_8567);
xnor U9421 (N_9421,N_8771,N_8608);
or U9422 (N_9422,N_8914,N_8527);
nand U9423 (N_9423,N_8707,N_8509);
and U9424 (N_9424,N_8887,N_8869);
nor U9425 (N_9425,N_8828,N_8992);
or U9426 (N_9426,N_8644,N_8789);
and U9427 (N_9427,N_8714,N_8932);
and U9428 (N_9428,N_8608,N_8581);
and U9429 (N_9429,N_8799,N_8844);
and U9430 (N_9430,N_8909,N_8938);
and U9431 (N_9431,N_8831,N_8755);
xnor U9432 (N_9432,N_8733,N_8763);
or U9433 (N_9433,N_8882,N_8571);
or U9434 (N_9434,N_8549,N_8952);
or U9435 (N_9435,N_8617,N_8891);
and U9436 (N_9436,N_8789,N_8662);
xnor U9437 (N_9437,N_8682,N_8964);
nor U9438 (N_9438,N_8993,N_8650);
xor U9439 (N_9439,N_8776,N_8974);
xor U9440 (N_9440,N_8546,N_8525);
xor U9441 (N_9441,N_8984,N_8671);
xor U9442 (N_9442,N_8679,N_8990);
xor U9443 (N_9443,N_8940,N_8711);
or U9444 (N_9444,N_8709,N_8513);
nor U9445 (N_9445,N_8902,N_8807);
nand U9446 (N_9446,N_8510,N_8663);
and U9447 (N_9447,N_8635,N_8841);
xor U9448 (N_9448,N_8712,N_8767);
xor U9449 (N_9449,N_8631,N_8661);
xnor U9450 (N_9450,N_8525,N_8792);
nor U9451 (N_9451,N_8928,N_8578);
and U9452 (N_9452,N_8912,N_8792);
nand U9453 (N_9453,N_8533,N_8699);
or U9454 (N_9454,N_8988,N_8653);
nor U9455 (N_9455,N_8869,N_8957);
xnor U9456 (N_9456,N_8925,N_8748);
nand U9457 (N_9457,N_8614,N_8679);
and U9458 (N_9458,N_8588,N_8839);
and U9459 (N_9459,N_8630,N_8568);
nand U9460 (N_9460,N_8714,N_8706);
or U9461 (N_9461,N_8538,N_8753);
or U9462 (N_9462,N_8544,N_8722);
and U9463 (N_9463,N_8522,N_8536);
and U9464 (N_9464,N_8625,N_8928);
and U9465 (N_9465,N_8914,N_8628);
or U9466 (N_9466,N_8970,N_8745);
nand U9467 (N_9467,N_8715,N_8591);
nand U9468 (N_9468,N_8904,N_8642);
nor U9469 (N_9469,N_8514,N_8894);
and U9470 (N_9470,N_8846,N_8744);
nor U9471 (N_9471,N_8859,N_8740);
xor U9472 (N_9472,N_8946,N_8825);
nor U9473 (N_9473,N_8594,N_8839);
xnor U9474 (N_9474,N_8946,N_8919);
or U9475 (N_9475,N_8722,N_8698);
or U9476 (N_9476,N_8992,N_8553);
or U9477 (N_9477,N_8644,N_8554);
xnor U9478 (N_9478,N_8848,N_8628);
or U9479 (N_9479,N_8858,N_8889);
or U9480 (N_9480,N_8536,N_8631);
or U9481 (N_9481,N_8589,N_8791);
and U9482 (N_9482,N_8521,N_8553);
nor U9483 (N_9483,N_8548,N_8526);
or U9484 (N_9484,N_8658,N_8765);
and U9485 (N_9485,N_8853,N_8627);
nand U9486 (N_9486,N_8970,N_8779);
or U9487 (N_9487,N_8504,N_8791);
nor U9488 (N_9488,N_8811,N_8587);
xor U9489 (N_9489,N_8939,N_8571);
nand U9490 (N_9490,N_8855,N_8569);
xnor U9491 (N_9491,N_8922,N_8861);
or U9492 (N_9492,N_8677,N_8794);
and U9493 (N_9493,N_8920,N_8687);
nor U9494 (N_9494,N_8586,N_8978);
and U9495 (N_9495,N_8783,N_8633);
nand U9496 (N_9496,N_8755,N_8744);
nand U9497 (N_9497,N_8887,N_8667);
xor U9498 (N_9498,N_8802,N_8595);
and U9499 (N_9499,N_8796,N_8568);
and U9500 (N_9500,N_9019,N_9397);
and U9501 (N_9501,N_9240,N_9303);
or U9502 (N_9502,N_9471,N_9372);
xnor U9503 (N_9503,N_9400,N_9042);
nand U9504 (N_9504,N_9158,N_9237);
nand U9505 (N_9505,N_9252,N_9073);
and U9506 (N_9506,N_9496,N_9263);
xnor U9507 (N_9507,N_9467,N_9379);
xor U9508 (N_9508,N_9211,N_9103);
or U9509 (N_9509,N_9183,N_9302);
nand U9510 (N_9510,N_9316,N_9175);
nor U9511 (N_9511,N_9254,N_9480);
nand U9512 (N_9512,N_9454,N_9179);
nor U9513 (N_9513,N_9007,N_9222);
or U9514 (N_9514,N_9061,N_9398);
xor U9515 (N_9515,N_9258,N_9220);
nand U9516 (N_9516,N_9416,N_9203);
or U9517 (N_9517,N_9050,N_9020);
nand U9518 (N_9518,N_9361,N_9148);
nor U9519 (N_9519,N_9250,N_9439);
nor U9520 (N_9520,N_9321,N_9425);
xnor U9521 (N_9521,N_9466,N_9077);
nand U9522 (N_9522,N_9185,N_9189);
nor U9523 (N_9523,N_9325,N_9352);
and U9524 (N_9524,N_9359,N_9125);
nor U9525 (N_9525,N_9449,N_9229);
xnor U9526 (N_9526,N_9230,N_9349);
and U9527 (N_9527,N_9193,N_9478);
nor U9528 (N_9528,N_9241,N_9364);
nand U9529 (N_9529,N_9371,N_9065);
nand U9530 (N_9530,N_9119,N_9226);
xor U9531 (N_9531,N_9054,N_9469);
or U9532 (N_9532,N_9289,N_9084);
or U9533 (N_9533,N_9433,N_9274);
nand U9534 (N_9534,N_9214,N_9368);
or U9535 (N_9535,N_9122,N_9011);
xnor U9536 (N_9536,N_9030,N_9370);
xor U9537 (N_9537,N_9451,N_9408);
nand U9538 (N_9538,N_9221,N_9188);
nand U9539 (N_9539,N_9184,N_9337);
nand U9540 (N_9540,N_9018,N_9431);
nand U9541 (N_9541,N_9197,N_9006);
or U9542 (N_9542,N_9163,N_9135);
nand U9543 (N_9543,N_9487,N_9051);
nor U9544 (N_9544,N_9315,N_9069);
xnor U9545 (N_9545,N_9311,N_9322);
nor U9546 (N_9546,N_9409,N_9426);
xor U9547 (N_9547,N_9173,N_9000);
nor U9548 (N_9548,N_9076,N_9096);
or U9549 (N_9549,N_9473,N_9150);
or U9550 (N_9550,N_9420,N_9381);
and U9551 (N_9551,N_9210,N_9208);
or U9552 (N_9552,N_9396,N_9055);
and U9553 (N_9553,N_9489,N_9291);
nor U9554 (N_9554,N_9190,N_9312);
xnor U9555 (N_9555,N_9114,N_9388);
or U9556 (N_9556,N_9213,N_9198);
xnor U9557 (N_9557,N_9204,N_9376);
and U9558 (N_9558,N_9491,N_9009);
and U9559 (N_9559,N_9106,N_9472);
or U9560 (N_9560,N_9477,N_9402);
nor U9561 (N_9561,N_9110,N_9029);
or U9562 (N_9562,N_9279,N_9448);
or U9563 (N_9563,N_9045,N_9025);
and U9564 (N_9564,N_9165,N_9206);
nand U9565 (N_9565,N_9378,N_9116);
and U9566 (N_9566,N_9046,N_9413);
nand U9567 (N_9567,N_9090,N_9068);
nor U9568 (N_9568,N_9357,N_9374);
nand U9569 (N_9569,N_9299,N_9201);
nand U9570 (N_9570,N_9373,N_9458);
or U9571 (N_9571,N_9281,N_9455);
or U9572 (N_9572,N_9486,N_9212);
or U9573 (N_9573,N_9465,N_9089);
nor U9574 (N_9574,N_9403,N_9334);
and U9575 (N_9575,N_9008,N_9301);
or U9576 (N_9576,N_9350,N_9387);
and U9577 (N_9577,N_9085,N_9259);
nand U9578 (N_9578,N_9355,N_9205);
xor U9579 (N_9579,N_9162,N_9117);
and U9580 (N_9580,N_9479,N_9139);
nor U9581 (N_9581,N_9293,N_9144);
xnor U9582 (N_9582,N_9039,N_9156);
and U9583 (N_9583,N_9481,N_9167);
nand U9584 (N_9584,N_9149,N_9394);
or U9585 (N_9585,N_9186,N_9271);
nor U9586 (N_9586,N_9384,N_9457);
xnor U9587 (N_9587,N_9490,N_9333);
and U9588 (N_9588,N_9497,N_9078);
xor U9589 (N_9589,N_9127,N_9238);
nor U9590 (N_9590,N_9245,N_9236);
or U9591 (N_9591,N_9306,N_9336);
or U9592 (N_9592,N_9243,N_9330);
xor U9593 (N_9593,N_9285,N_9356);
and U9594 (N_9594,N_9354,N_9035);
nand U9595 (N_9595,N_9423,N_9172);
or U9596 (N_9596,N_9217,N_9151);
and U9597 (N_9597,N_9468,N_9421);
nand U9598 (N_9598,N_9120,N_9001);
or U9599 (N_9599,N_9305,N_9192);
and U9600 (N_9600,N_9292,N_9200);
nor U9601 (N_9601,N_9121,N_9326);
and U9602 (N_9602,N_9032,N_9267);
or U9603 (N_9603,N_9016,N_9021);
and U9604 (N_9604,N_9256,N_9328);
and U9605 (N_9605,N_9154,N_9239);
or U9606 (N_9606,N_9434,N_9375);
or U9607 (N_9607,N_9363,N_9176);
xnor U9608 (N_9608,N_9273,N_9242);
and U9609 (N_9609,N_9335,N_9485);
xnor U9610 (N_9610,N_9099,N_9447);
or U9611 (N_9611,N_9474,N_9168);
or U9612 (N_9612,N_9499,N_9475);
or U9613 (N_9613,N_9010,N_9339);
xor U9614 (N_9614,N_9126,N_9304);
and U9615 (N_9615,N_9091,N_9385);
nor U9616 (N_9616,N_9268,N_9191);
and U9617 (N_9617,N_9164,N_9062);
xnor U9618 (N_9618,N_9283,N_9460);
or U9619 (N_9619,N_9253,N_9093);
xor U9620 (N_9620,N_9234,N_9058);
xnor U9621 (N_9621,N_9347,N_9174);
nand U9622 (N_9622,N_9298,N_9445);
nor U9623 (N_9623,N_9227,N_9442);
nand U9624 (N_9624,N_9128,N_9377);
nand U9625 (N_9625,N_9412,N_9170);
or U9626 (N_9626,N_9072,N_9310);
or U9627 (N_9627,N_9071,N_9307);
nor U9628 (N_9628,N_9075,N_9137);
nor U9629 (N_9629,N_9332,N_9041);
xor U9630 (N_9630,N_9470,N_9476);
or U9631 (N_9631,N_9047,N_9160);
and U9632 (N_9632,N_9023,N_9070);
and U9633 (N_9633,N_9251,N_9329);
nand U9634 (N_9634,N_9159,N_9209);
nand U9635 (N_9635,N_9092,N_9284);
and U9636 (N_9636,N_9414,N_9367);
nand U9637 (N_9637,N_9052,N_9436);
nor U9638 (N_9638,N_9083,N_9444);
nand U9639 (N_9639,N_9056,N_9429);
xnor U9640 (N_9640,N_9049,N_9112);
or U9641 (N_9641,N_9202,N_9287);
nand U9642 (N_9642,N_9063,N_9207);
and U9643 (N_9643,N_9080,N_9145);
nand U9644 (N_9644,N_9225,N_9262);
xnor U9645 (N_9645,N_9129,N_9405);
xnor U9646 (N_9646,N_9147,N_9105);
nand U9647 (N_9647,N_9157,N_9133);
nor U9648 (N_9648,N_9319,N_9053);
and U9649 (N_9649,N_9482,N_9483);
and U9650 (N_9650,N_9270,N_9134);
nor U9651 (N_9651,N_9410,N_9022);
and U9652 (N_9652,N_9484,N_9109);
xor U9653 (N_9653,N_9169,N_9180);
nor U9654 (N_9654,N_9343,N_9153);
nand U9655 (N_9655,N_9100,N_9277);
nand U9656 (N_9656,N_9098,N_9309);
xnor U9657 (N_9657,N_9456,N_9235);
or U9658 (N_9658,N_9044,N_9300);
nor U9659 (N_9659,N_9224,N_9358);
xnor U9660 (N_9660,N_9318,N_9081);
or U9661 (N_9661,N_9194,N_9104);
xor U9662 (N_9662,N_9146,N_9288);
and U9663 (N_9663,N_9248,N_9386);
or U9664 (N_9664,N_9215,N_9246);
nor U9665 (N_9665,N_9177,N_9255);
or U9666 (N_9666,N_9432,N_9113);
nor U9667 (N_9667,N_9247,N_9219);
nor U9668 (N_9668,N_9440,N_9462);
xnor U9669 (N_9669,N_9464,N_9026);
or U9670 (N_9670,N_9101,N_9024);
xnor U9671 (N_9671,N_9107,N_9115);
or U9672 (N_9672,N_9048,N_9232);
nor U9673 (N_9673,N_9348,N_9132);
or U9674 (N_9674,N_9111,N_9094);
nand U9675 (N_9675,N_9418,N_9441);
xnor U9676 (N_9676,N_9086,N_9494);
xor U9677 (N_9677,N_9435,N_9278);
nor U9678 (N_9678,N_9131,N_9317);
or U9679 (N_9679,N_9138,N_9040);
nand U9680 (N_9680,N_9275,N_9079);
and U9681 (N_9681,N_9261,N_9417);
and U9682 (N_9682,N_9463,N_9142);
xor U9683 (N_9683,N_9141,N_9216);
nand U9684 (N_9684,N_9282,N_9017);
and U9685 (N_9685,N_9295,N_9401);
or U9686 (N_9686,N_9004,N_9340);
nand U9687 (N_9687,N_9067,N_9108);
xor U9688 (N_9688,N_9257,N_9059);
nand U9689 (N_9689,N_9031,N_9492);
nor U9690 (N_9690,N_9264,N_9323);
xor U9691 (N_9691,N_9231,N_9057);
and U9692 (N_9692,N_9290,N_9269);
and U9693 (N_9693,N_9249,N_9028);
nand U9694 (N_9694,N_9074,N_9344);
and U9695 (N_9695,N_9296,N_9155);
nand U9696 (N_9696,N_9272,N_9260);
xnor U9697 (N_9697,N_9286,N_9452);
and U9698 (N_9698,N_9187,N_9060);
or U9699 (N_9699,N_9390,N_9082);
or U9700 (N_9700,N_9182,N_9228);
xor U9701 (N_9701,N_9351,N_9404);
nor U9702 (N_9702,N_9034,N_9218);
xor U9703 (N_9703,N_9037,N_9199);
nand U9704 (N_9704,N_9036,N_9196);
and U9705 (N_9705,N_9488,N_9143);
nand U9706 (N_9706,N_9012,N_9043);
and U9707 (N_9707,N_9331,N_9123);
nand U9708 (N_9708,N_9320,N_9038);
nor U9709 (N_9709,N_9498,N_9003);
nand U9710 (N_9710,N_9002,N_9389);
and U9711 (N_9711,N_9014,N_9424);
nor U9712 (N_9712,N_9195,N_9118);
and U9713 (N_9713,N_9136,N_9308);
and U9714 (N_9714,N_9391,N_9178);
xnor U9715 (N_9715,N_9280,N_9266);
nor U9716 (N_9716,N_9446,N_9276);
nor U9717 (N_9717,N_9015,N_9265);
and U9718 (N_9718,N_9140,N_9459);
or U9719 (N_9719,N_9066,N_9353);
nand U9720 (N_9720,N_9362,N_9161);
or U9721 (N_9721,N_9411,N_9422);
or U9722 (N_9722,N_9233,N_9097);
nand U9723 (N_9723,N_9366,N_9223);
xnor U9724 (N_9724,N_9453,N_9392);
or U9725 (N_9725,N_9027,N_9171);
nand U9726 (N_9726,N_9181,N_9102);
nand U9727 (N_9727,N_9346,N_9443);
and U9728 (N_9728,N_9380,N_9495);
or U9729 (N_9729,N_9345,N_9415);
or U9730 (N_9730,N_9393,N_9033);
nand U9731 (N_9731,N_9383,N_9088);
xor U9732 (N_9732,N_9395,N_9005);
and U9733 (N_9733,N_9152,N_9437);
xor U9734 (N_9734,N_9365,N_9341);
nor U9735 (N_9735,N_9166,N_9297);
or U9736 (N_9736,N_9294,N_9244);
nand U9737 (N_9737,N_9064,N_9087);
and U9738 (N_9738,N_9124,N_9406);
xnor U9739 (N_9739,N_9327,N_9324);
nand U9740 (N_9740,N_9130,N_9382);
xor U9741 (N_9741,N_9450,N_9493);
xnor U9742 (N_9742,N_9360,N_9399);
or U9743 (N_9743,N_9013,N_9430);
and U9744 (N_9744,N_9342,N_9314);
nand U9745 (N_9745,N_9369,N_9419);
xor U9746 (N_9746,N_9461,N_9427);
and U9747 (N_9747,N_9438,N_9407);
nor U9748 (N_9748,N_9338,N_9428);
and U9749 (N_9749,N_9313,N_9095);
and U9750 (N_9750,N_9118,N_9233);
nor U9751 (N_9751,N_9444,N_9403);
nor U9752 (N_9752,N_9235,N_9411);
and U9753 (N_9753,N_9288,N_9080);
or U9754 (N_9754,N_9306,N_9050);
nand U9755 (N_9755,N_9114,N_9160);
or U9756 (N_9756,N_9106,N_9376);
or U9757 (N_9757,N_9335,N_9321);
xnor U9758 (N_9758,N_9108,N_9418);
and U9759 (N_9759,N_9124,N_9280);
nor U9760 (N_9760,N_9088,N_9232);
and U9761 (N_9761,N_9446,N_9112);
nor U9762 (N_9762,N_9484,N_9040);
nor U9763 (N_9763,N_9035,N_9063);
nor U9764 (N_9764,N_9016,N_9327);
nand U9765 (N_9765,N_9121,N_9466);
and U9766 (N_9766,N_9248,N_9121);
or U9767 (N_9767,N_9156,N_9494);
nor U9768 (N_9768,N_9439,N_9220);
or U9769 (N_9769,N_9412,N_9019);
nand U9770 (N_9770,N_9055,N_9410);
xnor U9771 (N_9771,N_9455,N_9135);
or U9772 (N_9772,N_9138,N_9235);
nor U9773 (N_9773,N_9378,N_9194);
or U9774 (N_9774,N_9325,N_9099);
and U9775 (N_9775,N_9049,N_9181);
or U9776 (N_9776,N_9365,N_9075);
and U9777 (N_9777,N_9008,N_9053);
nand U9778 (N_9778,N_9465,N_9364);
nand U9779 (N_9779,N_9046,N_9469);
nor U9780 (N_9780,N_9271,N_9498);
or U9781 (N_9781,N_9330,N_9107);
and U9782 (N_9782,N_9163,N_9041);
xnor U9783 (N_9783,N_9430,N_9177);
or U9784 (N_9784,N_9047,N_9037);
or U9785 (N_9785,N_9448,N_9265);
nand U9786 (N_9786,N_9390,N_9153);
xnor U9787 (N_9787,N_9187,N_9201);
or U9788 (N_9788,N_9490,N_9439);
and U9789 (N_9789,N_9091,N_9296);
nand U9790 (N_9790,N_9378,N_9060);
nor U9791 (N_9791,N_9328,N_9316);
or U9792 (N_9792,N_9130,N_9468);
nor U9793 (N_9793,N_9308,N_9200);
and U9794 (N_9794,N_9287,N_9201);
or U9795 (N_9795,N_9445,N_9180);
nand U9796 (N_9796,N_9398,N_9068);
nor U9797 (N_9797,N_9226,N_9121);
and U9798 (N_9798,N_9173,N_9262);
xnor U9799 (N_9799,N_9191,N_9414);
nand U9800 (N_9800,N_9248,N_9442);
and U9801 (N_9801,N_9056,N_9029);
nand U9802 (N_9802,N_9060,N_9058);
nor U9803 (N_9803,N_9237,N_9332);
or U9804 (N_9804,N_9236,N_9284);
and U9805 (N_9805,N_9417,N_9223);
xor U9806 (N_9806,N_9449,N_9318);
xnor U9807 (N_9807,N_9152,N_9266);
xor U9808 (N_9808,N_9427,N_9494);
nand U9809 (N_9809,N_9461,N_9437);
nand U9810 (N_9810,N_9269,N_9455);
nand U9811 (N_9811,N_9370,N_9212);
or U9812 (N_9812,N_9263,N_9457);
nand U9813 (N_9813,N_9170,N_9372);
nand U9814 (N_9814,N_9185,N_9254);
xnor U9815 (N_9815,N_9139,N_9205);
xnor U9816 (N_9816,N_9446,N_9057);
or U9817 (N_9817,N_9366,N_9387);
nand U9818 (N_9818,N_9331,N_9132);
xnor U9819 (N_9819,N_9336,N_9207);
or U9820 (N_9820,N_9343,N_9259);
nor U9821 (N_9821,N_9438,N_9465);
nand U9822 (N_9822,N_9382,N_9078);
xor U9823 (N_9823,N_9199,N_9024);
xor U9824 (N_9824,N_9016,N_9129);
xnor U9825 (N_9825,N_9159,N_9483);
and U9826 (N_9826,N_9271,N_9441);
xor U9827 (N_9827,N_9280,N_9259);
nand U9828 (N_9828,N_9210,N_9146);
nor U9829 (N_9829,N_9010,N_9365);
and U9830 (N_9830,N_9405,N_9027);
nor U9831 (N_9831,N_9109,N_9313);
and U9832 (N_9832,N_9231,N_9145);
nand U9833 (N_9833,N_9395,N_9273);
xnor U9834 (N_9834,N_9249,N_9466);
and U9835 (N_9835,N_9409,N_9468);
nor U9836 (N_9836,N_9231,N_9025);
and U9837 (N_9837,N_9417,N_9036);
nand U9838 (N_9838,N_9453,N_9053);
nand U9839 (N_9839,N_9355,N_9337);
xor U9840 (N_9840,N_9343,N_9459);
or U9841 (N_9841,N_9490,N_9313);
or U9842 (N_9842,N_9477,N_9480);
nor U9843 (N_9843,N_9209,N_9219);
nand U9844 (N_9844,N_9372,N_9371);
and U9845 (N_9845,N_9498,N_9328);
nor U9846 (N_9846,N_9337,N_9300);
nor U9847 (N_9847,N_9222,N_9302);
nand U9848 (N_9848,N_9438,N_9208);
and U9849 (N_9849,N_9204,N_9273);
nand U9850 (N_9850,N_9399,N_9345);
nor U9851 (N_9851,N_9179,N_9465);
and U9852 (N_9852,N_9173,N_9454);
or U9853 (N_9853,N_9075,N_9344);
or U9854 (N_9854,N_9257,N_9343);
or U9855 (N_9855,N_9144,N_9495);
nand U9856 (N_9856,N_9406,N_9288);
or U9857 (N_9857,N_9273,N_9289);
or U9858 (N_9858,N_9319,N_9213);
xnor U9859 (N_9859,N_9328,N_9261);
nor U9860 (N_9860,N_9243,N_9392);
or U9861 (N_9861,N_9372,N_9490);
xnor U9862 (N_9862,N_9292,N_9164);
nand U9863 (N_9863,N_9430,N_9115);
nand U9864 (N_9864,N_9200,N_9288);
or U9865 (N_9865,N_9439,N_9107);
nand U9866 (N_9866,N_9179,N_9216);
nor U9867 (N_9867,N_9284,N_9330);
nor U9868 (N_9868,N_9391,N_9432);
and U9869 (N_9869,N_9076,N_9270);
nand U9870 (N_9870,N_9283,N_9121);
or U9871 (N_9871,N_9178,N_9113);
xnor U9872 (N_9872,N_9039,N_9314);
xor U9873 (N_9873,N_9429,N_9053);
nand U9874 (N_9874,N_9294,N_9436);
and U9875 (N_9875,N_9051,N_9248);
nor U9876 (N_9876,N_9390,N_9168);
and U9877 (N_9877,N_9476,N_9235);
and U9878 (N_9878,N_9041,N_9014);
or U9879 (N_9879,N_9341,N_9348);
and U9880 (N_9880,N_9088,N_9341);
nand U9881 (N_9881,N_9144,N_9054);
nand U9882 (N_9882,N_9457,N_9300);
nor U9883 (N_9883,N_9475,N_9220);
xnor U9884 (N_9884,N_9183,N_9389);
xor U9885 (N_9885,N_9178,N_9010);
and U9886 (N_9886,N_9080,N_9106);
nor U9887 (N_9887,N_9400,N_9388);
and U9888 (N_9888,N_9490,N_9078);
or U9889 (N_9889,N_9114,N_9493);
or U9890 (N_9890,N_9011,N_9124);
nor U9891 (N_9891,N_9086,N_9207);
xnor U9892 (N_9892,N_9073,N_9462);
and U9893 (N_9893,N_9378,N_9111);
nand U9894 (N_9894,N_9088,N_9097);
or U9895 (N_9895,N_9314,N_9293);
and U9896 (N_9896,N_9096,N_9056);
nor U9897 (N_9897,N_9163,N_9028);
nor U9898 (N_9898,N_9425,N_9005);
nor U9899 (N_9899,N_9368,N_9159);
and U9900 (N_9900,N_9212,N_9188);
xnor U9901 (N_9901,N_9139,N_9036);
and U9902 (N_9902,N_9464,N_9158);
xor U9903 (N_9903,N_9057,N_9274);
xnor U9904 (N_9904,N_9458,N_9161);
or U9905 (N_9905,N_9082,N_9114);
or U9906 (N_9906,N_9285,N_9069);
xor U9907 (N_9907,N_9365,N_9155);
or U9908 (N_9908,N_9047,N_9006);
nor U9909 (N_9909,N_9434,N_9251);
or U9910 (N_9910,N_9020,N_9255);
nand U9911 (N_9911,N_9311,N_9355);
or U9912 (N_9912,N_9018,N_9353);
or U9913 (N_9913,N_9148,N_9374);
xor U9914 (N_9914,N_9302,N_9364);
nand U9915 (N_9915,N_9278,N_9231);
and U9916 (N_9916,N_9304,N_9169);
nand U9917 (N_9917,N_9163,N_9481);
and U9918 (N_9918,N_9499,N_9147);
or U9919 (N_9919,N_9022,N_9171);
nand U9920 (N_9920,N_9344,N_9055);
or U9921 (N_9921,N_9253,N_9213);
nor U9922 (N_9922,N_9233,N_9136);
nor U9923 (N_9923,N_9216,N_9370);
or U9924 (N_9924,N_9245,N_9093);
and U9925 (N_9925,N_9251,N_9422);
and U9926 (N_9926,N_9337,N_9225);
xor U9927 (N_9927,N_9072,N_9416);
or U9928 (N_9928,N_9188,N_9247);
nand U9929 (N_9929,N_9137,N_9006);
and U9930 (N_9930,N_9019,N_9476);
and U9931 (N_9931,N_9475,N_9400);
nor U9932 (N_9932,N_9391,N_9418);
and U9933 (N_9933,N_9184,N_9158);
nand U9934 (N_9934,N_9135,N_9467);
and U9935 (N_9935,N_9298,N_9197);
nor U9936 (N_9936,N_9307,N_9344);
nand U9937 (N_9937,N_9073,N_9069);
nand U9938 (N_9938,N_9430,N_9436);
nor U9939 (N_9939,N_9119,N_9050);
and U9940 (N_9940,N_9086,N_9336);
and U9941 (N_9941,N_9487,N_9400);
nor U9942 (N_9942,N_9204,N_9379);
nor U9943 (N_9943,N_9047,N_9339);
nand U9944 (N_9944,N_9296,N_9191);
xor U9945 (N_9945,N_9293,N_9033);
or U9946 (N_9946,N_9280,N_9208);
nor U9947 (N_9947,N_9066,N_9041);
and U9948 (N_9948,N_9126,N_9397);
or U9949 (N_9949,N_9157,N_9254);
nor U9950 (N_9950,N_9169,N_9262);
xor U9951 (N_9951,N_9396,N_9178);
xor U9952 (N_9952,N_9170,N_9124);
nand U9953 (N_9953,N_9296,N_9194);
xnor U9954 (N_9954,N_9365,N_9141);
or U9955 (N_9955,N_9471,N_9222);
or U9956 (N_9956,N_9342,N_9344);
and U9957 (N_9957,N_9136,N_9166);
nor U9958 (N_9958,N_9028,N_9168);
and U9959 (N_9959,N_9419,N_9029);
and U9960 (N_9960,N_9142,N_9156);
xor U9961 (N_9961,N_9383,N_9478);
xor U9962 (N_9962,N_9071,N_9496);
xnor U9963 (N_9963,N_9071,N_9289);
or U9964 (N_9964,N_9201,N_9240);
or U9965 (N_9965,N_9494,N_9230);
and U9966 (N_9966,N_9119,N_9259);
xnor U9967 (N_9967,N_9175,N_9475);
nand U9968 (N_9968,N_9043,N_9047);
nand U9969 (N_9969,N_9412,N_9079);
and U9970 (N_9970,N_9019,N_9251);
or U9971 (N_9971,N_9016,N_9061);
or U9972 (N_9972,N_9469,N_9141);
or U9973 (N_9973,N_9269,N_9367);
nand U9974 (N_9974,N_9112,N_9247);
and U9975 (N_9975,N_9450,N_9050);
and U9976 (N_9976,N_9464,N_9004);
nor U9977 (N_9977,N_9024,N_9196);
nand U9978 (N_9978,N_9384,N_9003);
nand U9979 (N_9979,N_9421,N_9324);
xnor U9980 (N_9980,N_9490,N_9183);
nand U9981 (N_9981,N_9209,N_9324);
or U9982 (N_9982,N_9153,N_9114);
and U9983 (N_9983,N_9141,N_9059);
nor U9984 (N_9984,N_9193,N_9167);
nor U9985 (N_9985,N_9410,N_9264);
and U9986 (N_9986,N_9149,N_9366);
nor U9987 (N_9987,N_9017,N_9043);
xnor U9988 (N_9988,N_9198,N_9066);
xnor U9989 (N_9989,N_9285,N_9232);
and U9990 (N_9990,N_9163,N_9019);
nand U9991 (N_9991,N_9008,N_9229);
nor U9992 (N_9992,N_9139,N_9311);
xor U9993 (N_9993,N_9066,N_9383);
xnor U9994 (N_9994,N_9312,N_9428);
nand U9995 (N_9995,N_9400,N_9499);
nor U9996 (N_9996,N_9267,N_9138);
nor U9997 (N_9997,N_9401,N_9166);
nand U9998 (N_9998,N_9358,N_9112);
or U9999 (N_9999,N_9091,N_9372);
or U10000 (N_10000,N_9834,N_9958);
and U10001 (N_10001,N_9757,N_9631);
nor U10002 (N_10002,N_9963,N_9644);
nand U10003 (N_10003,N_9758,N_9756);
and U10004 (N_10004,N_9954,N_9895);
xnor U10005 (N_10005,N_9634,N_9830);
xor U10006 (N_10006,N_9686,N_9725);
xnor U10007 (N_10007,N_9549,N_9682);
or U10008 (N_10008,N_9743,N_9641);
or U10009 (N_10009,N_9558,N_9715);
nand U10010 (N_10010,N_9663,N_9560);
nor U10011 (N_10011,N_9734,N_9987);
or U10012 (N_10012,N_9646,N_9538);
or U10013 (N_10013,N_9600,N_9948);
or U10014 (N_10014,N_9654,N_9852);
nand U10015 (N_10015,N_9739,N_9590);
xnor U10016 (N_10016,N_9796,N_9992);
or U10017 (N_10017,N_9621,N_9694);
nor U10018 (N_10018,N_9604,N_9657);
and U10019 (N_10019,N_9862,N_9705);
or U10020 (N_10020,N_9993,N_9509);
nand U10021 (N_10021,N_9596,N_9607);
or U10022 (N_10022,N_9865,N_9848);
nor U10023 (N_10023,N_9773,N_9662);
xor U10024 (N_10024,N_9615,N_9584);
xor U10025 (N_10025,N_9971,N_9622);
and U10026 (N_10026,N_9599,N_9501);
or U10027 (N_10027,N_9626,N_9577);
nand U10028 (N_10028,N_9548,N_9966);
nand U10029 (N_10029,N_9831,N_9502);
xnor U10030 (N_10030,N_9611,N_9640);
nand U10031 (N_10031,N_9825,N_9962);
and U10032 (N_10032,N_9707,N_9866);
xnor U10033 (N_10033,N_9829,N_9949);
nand U10034 (N_10034,N_9534,N_9979);
nor U10035 (N_10035,N_9961,N_9935);
or U10036 (N_10036,N_9950,N_9770);
nand U10037 (N_10037,N_9585,N_9527);
or U10038 (N_10038,N_9827,N_9781);
nor U10039 (N_10039,N_9785,N_9598);
xor U10040 (N_10040,N_9513,N_9984);
or U10041 (N_10041,N_9815,N_9982);
or U10042 (N_10042,N_9760,N_9991);
nand U10043 (N_10043,N_9813,N_9505);
nor U10044 (N_10044,N_9768,N_9648);
nor U10045 (N_10045,N_9605,N_9575);
xnor U10046 (N_10046,N_9955,N_9944);
or U10047 (N_10047,N_9520,N_9582);
or U10048 (N_10048,N_9701,N_9591);
and U10049 (N_10049,N_9857,N_9587);
or U10050 (N_10050,N_9922,N_9891);
nand U10051 (N_10051,N_9983,N_9824);
or U10052 (N_10052,N_9702,N_9893);
nand U10053 (N_10053,N_9666,N_9875);
xnor U10054 (N_10054,N_9718,N_9897);
or U10055 (N_10055,N_9511,N_9800);
nor U10056 (N_10056,N_9579,N_9717);
nand U10057 (N_10057,N_9706,N_9907);
nand U10058 (N_10058,N_9833,N_9909);
nor U10059 (N_10059,N_9583,N_9592);
xnor U10060 (N_10060,N_9878,N_9661);
or U10061 (N_10061,N_9708,N_9931);
xor U10062 (N_10062,N_9550,N_9767);
xor U10063 (N_10063,N_9793,N_9943);
and U10064 (N_10064,N_9936,N_9782);
and U10065 (N_10065,N_9724,N_9610);
and U10066 (N_10066,N_9603,N_9716);
xor U10067 (N_10067,N_9990,N_9876);
nor U10068 (N_10068,N_9806,N_9899);
and U10069 (N_10069,N_9647,N_9761);
nor U10070 (N_10070,N_9925,N_9742);
or U10071 (N_10071,N_9981,N_9535);
and U10072 (N_10072,N_9602,N_9516);
nand U10073 (N_10073,N_9504,N_9567);
nor U10074 (N_10074,N_9589,N_9776);
nand U10075 (N_10075,N_9749,N_9561);
nand U10076 (N_10076,N_9960,N_9947);
or U10077 (N_10077,N_9506,N_9778);
xnor U10078 (N_10078,N_9737,N_9658);
or U10079 (N_10079,N_9816,N_9789);
or U10080 (N_10080,N_9747,N_9999);
nor U10081 (N_10081,N_9930,N_9555);
nand U10082 (N_10082,N_9517,N_9996);
or U10083 (N_10083,N_9787,N_9855);
or U10084 (N_10084,N_9727,N_9911);
nand U10085 (N_10085,N_9900,N_9945);
xnor U10086 (N_10086,N_9921,N_9632);
nor U10087 (N_10087,N_9653,N_9731);
and U10088 (N_10088,N_9522,N_9942);
xor U10089 (N_10089,N_9914,N_9854);
nand U10090 (N_10090,N_9552,N_9721);
nor U10091 (N_10091,N_9918,N_9571);
and U10092 (N_10092,N_9894,N_9869);
nand U10093 (N_10093,N_9643,N_9569);
xor U10094 (N_10094,N_9978,N_9856);
and U10095 (N_10095,N_9551,N_9629);
nand U10096 (N_10096,N_9753,N_9623);
nand U10097 (N_10097,N_9872,N_9566);
nor U10098 (N_10098,N_9843,N_9881);
nor U10099 (N_10099,N_9529,N_9597);
or U10100 (N_10100,N_9951,N_9545);
or U10101 (N_10101,N_9885,N_9637);
xor U10102 (N_10102,N_9710,N_9847);
nor U10103 (N_10103,N_9559,N_9692);
nand U10104 (N_10104,N_9563,N_9515);
and U10105 (N_10105,N_9803,N_9941);
nand U10106 (N_10106,N_9849,N_9639);
nand U10107 (N_10107,N_9959,N_9606);
nand U10108 (N_10108,N_9539,N_9635);
nand U10109 (N_10109,N_9788,N_9860);
xnor U10110 (N_10110,N_9898,N_9861);
nor U10111 (N_10111,N_9526,N_9953);
nand U10112 (N_10112,N_9904,N_9617);
nor U10113 (N_10113,N_9593,N_9542);
nand U10114 (N_10114,N_9884,N_9573);
nor U10115 (N_10115,N_9874,N_9828);
or U10116 (N_10116,N_9636,N_9888);
and U10117 (N_10117,N_9883,N_9985);
nor U10118 (N_10118,N_9811,N_9687);
xnor U10119 (N_10119,N_9609,N_9798);
xor U10120 (N_10120,N_9524,N_9614);
nor U10121 (N_10121,N_9998,N_9882);
or U10122 (N_10122,N_9932,N_9937);
and U10123 (N_10123,N_9752,N_9871);
nand U10124 (N_10124,N_9576,N_9741);
nor U10125 (N_10125,N_9938,N_9695);
and U10126 (N_10126,N_9858,N_9667);
or U10127 (N_10127,N_9842,N_9809);
or U10128 (N_10128,N_9863,N_9870);
and U10129 (N_10129,N_9818,N_9650);
or U10130 (N_10130,N_9508,N_9656);
nand U10131 (N_10131,N_9927,N_9759);
xor U10132 (N_10132,N_9722,N_9946);
xor U10133 (N_10133,N_9698,N_9988);
and U10134 (N_10134,N_9807,N_9673);
nor U10135 (N_10135,N_9703,N_9832);
xor U10136 (N_10136,N_9810,N_9572);
nand U10137 (N_10137,N_9709,N_9671);
nand U10138 (N_10138,N_9915,N_9926);
and U10139 (N_10139,N_9664,N_9746);
xor U10140 (N_10140,N_9578,N_9821);
or U10141 (N_10141,N_9730,N_9919);
xor U10142 (N_10142,N_9503,N_9714);
nand U10143 (N_10143,N_9887,N_9823);
or U10144 (N_10144,N_9543,N_9586);
nor U10145 (N_10145,N_9917,N_9952);
nand U10146 (N_10146,N_9697,N_9772);
and U10147 (N_10147,N_9525,N_9696);
and U10148 (N_10148,N_9726,N_9808);
and U10149 (N_10149,N_9774,N_9906);
xnor U10150 (N_10150,N_9612,N_9537);
nor U10151 (N_10151,N_9514,N_9700);
nand U10152 (N_10152,N_9512,N_9536);
and U10153 (N_10153,N_9685,N_9690);
nand U10154 (N_10154,N_9674,N_9812);
nand U10155 (N_10155,N_9751,N_9997);
nand U10156 (N_10156,N_9970,N_9836);
xor U10157 (N_10157,N_9994,N_9704);
or U10158 (N_10158,N_9595,N_9713);
or U10159 (N_10159,N_9556,N_9564);
or U10160 (N_10160,N_9972,N_9826);
nand U10161 (N_10161,N_9557,N_9608);
or U10162 (N_10162,N_9581,N_9755);
nor U10163 (N_10163,N_9528,N_9819);
and U10164 (N_10164,N_9839,N_9873);
nor U10165 (N_10165,N_9754,N_9676);
or U10166 (N_10166,N_9628,N_9968);
or U10167 (N_10167,N_9799,N_9570);
nor U10168 (N_10168,N_9840,N_9923);
and U10169 (N_10169,N_9765,N_9892);
xnor U10170 (N_10170,N_9740,N_9678);
nand U10171 (N_10171,N_9601,N_9651);
nand U10172 (N_10172,N_9735,N_9633);
nand U10173 (N_10173,N_9684,N_9780);
or U10174 (N_10174,N_9835,N_9928);
or U10175 (N_10175,N_9507,N_9691);
and U10176 (N_10176,N_9912,N_9521);
nand U10177 (N_10177,N_9896,N_9940);
xor U10178 (N_10178,N_9680,N_9784);
and U10179 (N_10179,N_9613,N_9973);
nor U10180 (N_10180,N_9820,N_9764);
xnor U10181 (N_10181,N_9531,N_9733);
or U10182 (N_10182,N_9804,N_9544);
or U10183 (N_10183,N_9574,N_9546);
and U10184 (N_10184,N_9792,N_9649);
or U10185 (N_10185,N_9879,N_9689);
and U10186 (N_10186,N_9795,N_9630);
and U10187 (N_10187,N_9890,N_9967);
xnor U10188 (N_10188,N_9777,N_9995);
or U10189 (N_10189,N_9619,N_9642);
and U10190 (N_10190,N_9801,N_9976);
nor U10191 (N_10191,N_9791,N_9748);
or U10192 (N_10192,N_9594,N_9977);
and U10193 (N_10193,N_9660,N_9625);
nor U10194 (N_10194,N_9822,N_9723);
nand U10195 (N_10195,N_9920,N_9986);
xnor U10196 (N_10196,N_9889,N_9500);
xnor U10197 (N_10197,N_9845,N_9568);
nor U10198 (N_10198,N_9779,N_9580);
and U10199 (N_10199,N_9533,N_9699);
and U10200 (N_10200,N_9547,N_9837);
nor U10201 (N_10201,N_9519,N_9553);
nand U10202 (N_10202,N_9974,N_9901);
xor U10203 (N_10203,N_9817,N_9880);
nor U10204 (N_10204,N_9775,N_9965);
and U10205 (N_10205,N_9763,N_9956);
xnor U10206 (N_10206,N_9910,N_9797);
nor U10207 (N_10207,N_9805,N_9744);
and U10208 (N_10208,N_9729,N_9638);
and U10209 (N_10209,N_9850,N_9957);
xnor U10210 (N_10210,N_9720,N_9980);
or U10211 (N_10211,N_9939,N_9877);
and U10212 (N_10212,N_9908,N_9924);
xnor U10213 (N_10213,N_9802,N_9745);
nor U10214 (N_10214,N_9933,N_9719);
xnor U10215 (N_10215,N_9620,N_9868);
or U10216 (N_10216,N_9645,N_9736);
or U10217 (N_10217,N_9652,N_9732);
nor U10218 (N_10218,N_9853,N_9670);
and U10219 (N_10219,N_9934,N_9964);
nor U10220 (N_10220,N_9711,N_9624);
nor U10221 (N_10221,N_9588,N_9905);
nor U10222 (N_10222,N_9675,N_9541);
nor U10223 (N_10223,N_9668,N_9864);
xnor U10224 (N_10224,N_9532,N_9783);
nand U10225 (N_10225,N_9867,N_9814);
nor U10226 (N_10226,N_9540,N_9728);
or U10227 (N_10227,N_9616,N_9669);
nand U10228 (N_10228,N_9851,N_9738);
and U10229 (N_10229,N_9530,N_9846);
nor U10230 (N_10230,N_9762,N_9750);
xor U10231 (N_10231,N_9655,N_9929);
nand U10232 (N_10232,N_9677,N_9902);
nand U10233 (N_10233,N_9565,N_9518);
nand U10234 (N_10234,N_9665,N_9989);
and U10235 (N_10235,N_9903,N_9771);
and U10236 (N_10236,N_9618,N_9859);
and U10237 (N_10237,N_9681,N_9627);
and U10238 (N_10238,N_9523,N_9554);
or U10239 (N_10239,N_9886,N_9786);
or U10240 (N_10240,N_9838,N_9969);
nand U10241 (N_10241,N_9913,N_9683);
or U10242 (N_10242,N_9790,N_9712);
nand U10243 (N_10243,N_9672,N_9841);
xnor U10244 (N_10244,N_9679,N_9510);
nand U10245 (N_10245,N_9844,N_9688);
nor U10246 (N_10246,N_9794,N_9693);
nand U10247 (N_10247,N_9659,N_9766);
or U10248 (N_10248,N_9916,N_9562);
and U10249 (N_10249,N_9769,N_9975);
and U10250 (N_10250,N_9684,N_9635);
or U10251 (N_10251,N_9511,N_9958);
and U10252 (N_10252,N_9614,N_9928);
nand U10253 (N_10253,N_9510,N_9976);
nor U10254 (N_10254,N_9547,N_9790);
xor U10255 (N_10255,N_9986,N_9957);
nor U10256 (N_10256,N_9958,N_9692);
xor U10257 (N_10257,N_9938,N_9834);
or U10258 (N_10258,N_9526,N_9666);
nand U10259 (N_10259,N_9559,N_9636);
or U10260 (N_10260,N_9810,N_9936);
and U10261 (N_10261,N_9824,N_9793);
xnor U10262 (N_10262,N_9766,N_9649);
nor U10263 (N_10263,N_9901,N_9667);
and U10264 (N_10264,N_9968,N_9693);
or U10265 (N_10265,N_9661,N_9853);
nor U10266 (N_10266,N_9865,N_9661);
and U10267 (N_10267,N_9868,N_9824);
or U10268 (N_10268,N_9864,N_9674);
nand U10269 (N_10269,N_9642,N_9620);
nand U10270 (N_10270,N_9738,N_9987);
and U10271 (N_10271,N_9782,N_9634);
and U10272 (N_10272,N_9915,N_9996);
nand U10273 (N_10273,N_9703,N_9601);
and U10274 (N_10274,N_9635,N_9967);
nor U10275 (N_10275,N_9517,N_9869);
nand U10276 (N_10276,N_9775,N_9999);
nor U10277 (N_10277,N_9899,N_9556);
xnor U10278 (N_10278,N_9822,N_9826);
or U10279 (N_10279,N_9530,N_9977);
xnor U10280 (N_10280,N_9510,N_9571);
and U10281 (N_10281,N_9512,N_9825);
xor U10282 (N_10282,N_9634,N_9793);
nand U10283 (N_10283,N_9591,N_9809);
nand U10284 (N_10284,N_9565,N_9925);
and U10285 (N_10285,N_9811,N_9879);
nor U10286 (N_10286,N_9967,N_9566);
or U10287 (N_10287,N_9946,N_9675);
nand U10288 (N_10288,N_9661,N_9881);
nand U10289 (N_10289,N_9646,N_9932);
nand U10290 (N_10290,N_9610,N_9687);
nand U10291 (N_10291,N_9603,N_9687);
and U10292 (N_10292,N_9538,N_9768);
xnor U10293 (N_10293,N_9919,N_9567);
nor U10294 (N_10294,N_9510,N_9733);
or U10295 (N_10295,N_9730,N_9863);
nand U10296 (N_10296,N_9723,N_9504);
and U10297 (N_10297,N_9928,N_9776);
and U10298 (N_10298,N_9577,N_9721);
nor U10299 (N_10299,N_9753,N_9875);
or U10300 (N_10300,N_9725,N_9517);
xor U10301 (N_10301,N_9951,N_9583);
xor U10302 (N_10302,N_9726,N_9707);
and U10303 (N_10303,N_9757,N_9682);
and U10304 (N_10304,N_9519,N_9790);
or U10305 (N_10305,N_9733,N_9858);
nand U10306 (N_10306,N_9654,N_9890);
nor U10307 (N_10307,N_9601,N_9976);
and U10308 (N_10308,N_9668,N_9822);
and U10309 (N_10309,N_9963,N_9609);
xor U10310 (N_10310,N_9759,N_9790);
xnor U10311 (N_10311,N_9969,N_9653);
nor U10312 (N_10312,N_9503,N_9720);
nor U10313 (N_10313,N_9500,N_9868);
or U10314 (N_10314,N_9831,N_9559);
nand U10315 (N_10315,N_9518,N_9921);
xnor U10316 (N_10316,N_9642,N_9793);
or U10317 (N_10317,N_9797,N_9764);
xor U10318 (N_10318,N_9576,N_9662);
or U10319 (N_10319,N_9824,N_9680);
nand U10320 (N_10320,N_9527,N_9744);
and U10321 (N_10321,N_9545,N_9768);
nand U10322 (N_10322,N_9887,N_9694);
nor U10323 (N_10323,N_9711,N_9634);
or U10324 (N_10324,N_9535,N_9600);
and U10325 (N_10325,N_9689,N_9655);
nand U10326 (N_10326,N_9651,N_9882);
or U10327 (N_10327,N_9753,N_9563);
and U10328 (N_10328,N_9544,N_9896);
xor U10329 (N_10329,N_9573,N_9571);
xnor U10330 (N_10330,N_9540,N_9860);
and U10331 (N_10331,N_9966,N_9973);
nor U10332 (N_10332,N_9763,N_9693);
nor U10333 (N_10333,N_9506,N_9731);
or U10334 (N_10334,N_9713,N_9738);
xnor U10335 (N_10335,N_9987,N_9826);
and U10336 (N_10336,N_9679,N_9605);
and U10337 (N_10337,N_9812,N_9547);
or U10338 (N_10338,N_9895,N_9557);
nand U10339 (N_10339,N_9939,N_9657);
xnor U10340 (N_10340,N_9985,N_9998);
xor U10341 (N_10341,N_9520,N_9581);
or U10342 (N_10342,N_9571,N_9543);
nand U10343 (N_10343,N_9531,N_9684);
and U10344 (N_10344,N_9610,N_9634);
or U10345 (N_10345,N_9639,N_9916);
or U10346 (N_10346,N_9905,N_9608);
nor U10347 (N_10347,N_9694,N_9644);
nor U10348 (N_10348,N_9907,N_9579);
and U10349 (N_10349,N_9913,N_9550);
or U10350 (N_10350,N_9850,N_9508);
or U10351 (N_10351,N_9509,N_9971);
or U10352 (N_10352,N_9660,N_9892);
or U10353 (N_10353,N_9741,N_9712);
nand U10354 (N_10354,N_9879,N_9528);
nand U10355 (N_10355,N_9924,N_9692);
nor U10356 (N_10356,N_9546,N_9836);
nand U10357 (N_10357,N_9509,N_9764);
nand U10358 (N_10358,N_9551,N_9883);
nor U10359 (N_10359,N_9751,N_9564);
nor U10360 (N_10360,N_9733,N_9633);
and U10361 (N_10361,N_9736,N_9829);
nand U10362 (N_10362,N_9724,N_9567);
or U10363 (N_10363,N_9788,N_9987);
xor U10364 (N_10364,N_9594,N_9606);
nor U10365 (N_10365,N_9655,N_9686);
nand U10366 (N_10366,N_9717,N_9669);
or U10367 (N_10367,N_9722,N_9548);
nor U10368 (N_10368,N_9871,N_9523);
or U10369 (N_10369,N_9912,N_9600);
or U10370 (N_10370,N_9835,N_9796);
nand U10371 (N_10371,N_9819,N_9709);
nand U10372 (N_10372,N_9584,N_9535);
or U10373 (N_10373,N_9648,N_9646);
nor U10374 (N_10374,N_9769,N_9817);
xnor U10375 (N_10375,N_9760,N_9618);
xnor U10376 (N_10376,N_9825,N_9716);
nand U10377 (N_10377,N_9922,N_9627);
xnor U10378 (N_10378,N_9526,N_9644);
or U10379 (N_10379,N_9765,N_9941);
xnor U10380 (N_10380,N_9997,N_9588);
and U10381 (N_10381,N_9683,N_9732);
nor U10382 (N_10382,N_9962,N_9742);
nor U10383 (N_10383,N_9630,N_9773);
nor U10384 (N_10384,N_9903,N_9607);
and U10385 (N_10385,N_9639,N_9783);
xor U10386 (N_10386,N_9673,N_9918);
or U10387 (N_10387,N_9924,N_9902);
and U10388 (N_10388,N_9607,N_9962);
nand U10389 (N_10389,N_9525,N_9788);
or U10390 (N_10390,N_9547,N_9612);
nor U10391 (N_10391,N_9975,N_9594);
or U10392 (N_10392,N_9830,N_9668);
nor U10393 (N_10393,N_9880,N_9546);
nor U10394 (N_10394,N_9514,N_9500);
or U10395 (N_10395,N_9563,N_9778);
nor U10396 (N_10396,N_9716,N_9985);
and U10397 (N_10397,N_9654,N_9988);
and U10398 (N_10398,N_9875,N_9665);
and U10399 (N_10399,N_9586,N_9989);
xor U10400 (N_10400,N_9972,N_9723);
xor U10401 (N_10401,N_9602,N_9975);
nand U10402 (N_10402,N_9969,N_9786);
xor U10403 (N_10403,N_9949,N_9709);
nor U10404 (N_10404,N_9797,N_9694);
nand U10405 (N_10405,N_9969,N_9949);
nand U10406 (N_10406,N_9606,N_9914);
nor U10407 (N_10407,N_9864,N_9787);
or U10408 (N_10408,N_9534,N_9671);
nor U10409 (N_10409,N_9514,N_9776);
nor U10410 (N_10410,N_9833,N_9964);
xor U10411 (N_10411,N_9660,N_9912);
xor U10412 (N_10412,N_9962,N_9757);
or U10413 (N_10413,N_9705,N_9951);
xnor U10414 (N_10414,N_9899,N_9779);
xor U10415 (N_10415,N_9818,N_9903);
nand U10416 (N_10416,N_9782,N_9642);
and U10417 (N_10417,N_9516,N_9802);
xor U10418 (N_10418,N_9848,N_9934);
xor U10419 (N_10419,N_9519,N_9758);
and U10420 (N_10420,N_9784,N_9800);
nor U10421 (N_10421,N_9748,N_9823);
or U10422 (N_10422,N_9954,N_9782);
nor U10423 (N_10423,N_9967,N_9786);
or U10424 (N_10424,N_9606,N_9915);
nand U10425 (N_10425,N_9872,N_9985);
nor U10426 (N_10426,N_9927,N_9526);
or U10427 (N_10427,N_9912,N_9631);
nand U10428 (N_10428,N_9670,N_9858);
nand U10429 (N_10429,N_9519,N_9576);
or U10430 (N_10430,N_9629,N_9873);
nor U10431 (N_10431,N_9543,N_9506);
nor U10432 (N_10432,N_9968,N_9909);
nor U10433 (N_10433,N_9601,N_9655);
nand U10434 (N_10434,N_9526,N_9878);
or U10435 (N_10435,N_9999,N_9754);
or U10436 (N_10436,N_9957,N_9739);
or U10437 (N_10437,N_9787,N_9528);
xor U10438 (N_10438,N_9530,N_9622);
xnor U10439 (N_10439,N_9505,N_9610);
and U10440 (N_10440,N_9864,N_9608);
nor U10441 (N_10441,N_9585,N_9967);
and U10442 (N_10442,N_9591,N_9811);
xnor U10443 (N_10443,N_9753,N_9959);
nor U10444 (N_10444,N_9920,N_9736);
xor U10445 (N_10445,N_9851,N_9776);
and U10446 (N_10446,N_9552,N_9906);
xor U10447 (N_10447,N_9925,N_9718);
xnor U10448 (N_10448,N_9847,N_9599);
nor U10449 (N_10449,N_9696,N_9839);
nand U10450 (N_10450,N_9835,N_9780);
or U10451 (N_10451,N_9699,N_9819);
nand U10452 (N_10452,N_9556,N_9661);
xor U10453 (N_10453,N_9501,N_9945);
xnor U10454 (N_10454,N_9912,N_9630);
nor U10455 (N_10455,N_9658,N_9888);
and U10456 (N_10456,N_9927,N_9793);
nand U10457 (N_10457,N_9864,N_9769);
and U10458 (N_10458,N_9593,N_9946);
and U10459 (N_10459,N_9939,N_9896);
nor U10460 (N_10460,N_9625,N_9794);
nand U10461 (N_10461,N_9645,N_9587);
and U10462 (N_10462,N_9888,N_9688);
or U10463 (N_10463,N_9799,N_9644);
xor U10464 (N_10464,N_9957,N_9807);
and U10465 (N_10465,N_9635,N_9538);
nor U10466 (N_10466,N_9730,N_9530);
nor U10467 (N_10467,N_9758,N_9912);
nand U10468 (N_10468,N_9552,N_9814);
nand U10469 (N_10469,N_9985,N_9681);
and U10470 (N_10470,N_9808,N_9559);
nor U10471 (N_10471,N_9545,N_9904);
xor U10472 (N_10472,N_9911,N_9520);
and U10473 (N_10473,N_9508,N_9613);
xor U10474 (N_10474,N_9762,N_9732);
or U10475 (N_10475,N_9856,N_9961);
and U10476 (N_10476,N_9842,N_9901);
xnor U10477 (N_10477,N_9818,N_9562);
xnor U10478 (N_10478,N_9751,N_9738);
or U10479 (N_10479,N_9917,N_9804);
and U10480 (N_10480,N_9819,N_9669);
xor U10481 (N_10481,N_9504,N_9830);
and U10482 (N_10482,N_9636,N_9611);
nor U10483 (N_10483,N_9533,N_9866);
xor U10484 (N_10484,N_9650,N_9813);
xor U10485 (N_10485,N_9994,N_9767);
xnor U10486 (N_10486,N_9716,N_9519);
and U10487 (N_10487,N_9942,N_9940);
nand U10488 (N_10488,N_9743,N_9683);
and U10489 (N_10489,N_9656,N_9689);
or U10490 (N_10490,N_9708,N_9817);
nand U10491 (N_10491,N_9595,N_9936);
xnor U10492 (N_10492,N_9778,N_9933);
xnor U10493 (N_10493,N_9601,N_9504);
and U10494 (N_10494,N_9963,N_9732);
or U10495 (N_10495,N_9971,N_9916);
or U10496 (N_10496,N_9731,N_9705);
nor U10497 (N_10497,N_9676,N_9951);
or U10498 (N_10498,N_9902,N_9949);
nor U10499 (N_10499,N_9684,N_9790);
nand U10500 (N_10500,N_10386,N_10241);
nand U10501 (N_10501,N_10072,N_10158);
and U10502 (N_10502,N_10467,N_10017);
or U10503 (N_10503,N_10197,N_10019);
or U10504 (N_10504,N_10012,N_10227);
or U10505 (N_10505,N_10151,N_10496);
nand U10506 (N_10506,N_10368,N_10491);
xor U10507 (N_10507,N_10402,N_10294);
nand U10508 (N_10508,N_10417,N_10150);
xor U10509 (N_10509,N_10461,N_10361);
nor U10510 (N_10510,N_10222,N_10442);
xnor U10511 (N_10511,N_10114,N_10199);
and U10512 (N_10512,N_10468,N_10046);
nand U10513 (N_10513,N_10438,N_10425);
nand U10514 (N_10514,N_10000,N_10236);
nand U10515 (N_10515,N_10443,N_10297);
or U10516 (N_10516,N_10245,N_10489);
nor U10517 (N_10517,N_10117,N_10176);
xor U10518 (N_10518,N_10095,N_10166);
xor U10519 (N_10519,N_10265,N_10193);
nor U10520 (N_10520,N_10357,N_10015);
or U10521 (N_10521,N_10484,N_10131);
nand U10522 (N_10522,N_10080,N_10266);
and U10523 (N_10523,N_10454,N_10208);
xnor U10524 (N_10524,N_10397,N_10141);
nand U10525 (N_10525,N_10343,N_10204);
xnor U10526 (N_10526,N_10380,N_10440);
nor U10527 (N_10527,N_10198,N_10211);
or U10528 (N_10528,N_10153,N_10200);
or U10529 (N_10529,N_10486,N_10143);
and U10530 (N_10530,N_10243,N_10161);
nand U10531 (N_10531,N_10326,N_10292);
and U10532 (N_10532,N_10270,N_10394);
and U10533 (N_10533,N_10447,N_10410);
nor U10534 (N_10534,N_10455,N_10273);
and U10535 (N_10535,N_10363,N_10385);
xnor U10536 (N_10536,N_10278,N_10427);
nand U10537 (N_10537,N_10445,N_10331);
or U10538 (N_10538,N_10157,N_10418);
nand U10539 (N_10539,N_10185,N_10182);
nand U10540 (N_10540,N_10372,N_10456);
and U10541 (N_10541,N_10421,N_10003);
xor U10542 (N_10542,N_10162,N_10248);
and U10543 (N_10543,N_10275,N_10173);
nand U10544 (N_10544,N_10287,N_10190);
xnor U10545 (N_10545,N_10170,N_10481);
nor U10546 (N_10546,N_10281,N_10063);
and U10547 (N_10547,N_10459,N_10233);
nor U10548 (N_10548,N_10450,N_10276);
and U10549 (N_10549,N_10487,N_10422);
and U10550 (N_10550,N_10296,N_10317);
or U10551 (N_10551,N_10283,N_10097);
or U10552 (N_10552,N_10498,N_10123);
xnor U10553 (N_10553,N_10262,N_10137);
nor U10554 (N_10554,N_10068,N_10257);
xor U10555 (N_10555,N_10469,N_10007);
nand U10556 (N_10556,N_10269,N_10446);
and U10557 (N_10557,N_10395,N_10099);
and U10558 (N_10558,N_10285,N_10255);
and U10559 (N_10559,N_10074,N_10249);
xnor U10560 (N_10560,N_10356,N_10010);
or U10561 (N_10561,N_10430,N_10240);
and U10562 (N_10562,N_10105,N_10493);
and U10563 (N_10563,N_10164,N_10055);
nand U10564 (N_10564,N_10186,N_10061);
nor U10565 (N_10565,N_10154,N_10100);
xnor U10566 (N_10566,N_10339,N_10094);
and U10567 (N_10567,N_10050,N_10411);
nor U10568 (N_10568,N_10047,N_10079);
nor U10569 (N_10569,N_10439,N_10478);
xnor U10570 (N_10570,N_10124,N_10412);
or U10571 (N_10571,N_10212,N_10414);
or U10572 (N_10572,N_10234,N_10349);
nor U10573 (N_10573,N_10036,N_10284);
or U10574 (N_10574,N_10174,N_10470);
nor U10575 (N_10575,N_10021,N_10256);
or U10576 (N_10576,N_10024,N_10353);
and U10577 (N_10577,N_10136,N_10220);
or U10578 (N_10578,N_10328,N_10319);
or U10579 (N_10579,N_10464,N_10434);
or U10580 (N_10580,N_10277,N_10147);
and U10581 (N_10581,N_10293,N_10355);
nor U10582 (N_10582,N_10235,N_10376);
nand U10583 (N_10583,N_10033,N_10078);
nand U10584 (N_10584,N_10318,N_10300);
or U10585 (N_10585,N_10302,N_10130);
or U10586 (N_10586,N_10098,N_10336);
or U10587 (N_10587,N_10121,N_10022);
nand U10588 (N_10588,N_10112,N_10457);
xor U10589 (N_10589,N_10289,N_10404);
or U10590 (N_10590,N_10118,N_10366);
xor U10591 (N_10591,N_10159,N_10320);
or U10592 (N_10592,N_10031,N_10035);
and U10593 (N_10593,N_10334,N_10303);
and U10594 (N_10594,N_10299,N_10428);
or U10595 (N_10595,N_10217,N_10373);
and U10596 (N_10596,N_10310,N_10383);
and U10597 (N_10597,N_10314,N_10305);
xor U10598 (N_10598,N_10056,N_10044);
xnor U10599 (N_10599,N_10030,N_10230);
nor U10600 (N_10600,N_10347,N_10466);
and U10601 (N_10601,N_10040,N_10145);
and U10602 (N_10602,N_10316,N_10206);
xor U10603 (N_10603,N_10312,N_10436);
nor U10604 (N_10604,N_10238,N_10499);
xnor U10605 (N_10605,N_10377,N_10067);
xor U10606 (N_10606,N_10229,N_10407);
nand U10607 (N_10607,N_10142,N_10110);
nand U10608 (N_10608,N_10350,N_10179);
nor U10609 (N_10609,N_10225,N_10191);
nor U10610 (N_10610,N_10183,N_10156);
and U10611 (N_10611,N_10474,N_10382);
xnor U10612 (N_10612,N_10471,N_10215);
nand U10613 (N_10613,N_10398,N_10420);
xnor U10614 (N_10614,N_10133,N_10253);
or U10615 (N_10615,N_10060,N_10144);
nand U10616 (N_10616,N_10419,N_10274);
xor U10617 (N_10617,N_10004,N_10002);
and U10618 (N_10618,N_10093,N_10125);
and U10619 (N_10619,N_10059,N_10013);
nand U10620 (N_10620,N_10309,N_10090);
or U10621 (N_10621,N_10213,N_10492);
xor U10622 (N_10622,N_10338,N_10387);
nand U10623 (N_10623,N_10108,N_10160);
or U10624 (N_10624,N_10135,N_10237);
nor U10625 (N_10625,N_10052,N_10006);
nor U10626 (N_10626,N_10483,N_10329);
nand U10627 (N_10627,N_10401,N_10202);
xor U10628 (N_10628,N_10152,N_10113);
and U10629 (N_10629,N_10038,N_10458);
nand U10630 (N_10630,N_10034,N_10122);
nand U10631 (N_10631,N_10083,N_10087);
nor U10632 (N_10632,N_10167,N_10494);
nor U10633 (N_10633,N_10129,N_10128);
or U10634 (N_10634,N_10088,N_10239);
and U10635 (N_10635,N_10340,N_10023);
xnor U10636 (N_10636,N_10084,N_10077);
nand U10637 (N_10637,N_10140,N_10037);
nand U10638 (N_10638,N_10379,N_10330);
nor U10639 (N_10639,N_10058,N_10026);
nand U10640 (N_10640,N_10244,N_10221);
nor U10641 (N_10641,N_10096,N_10403);
nor U10642 (N_10642,N_10231,N_10441);
or U10643 (N_10643,N_10264,N_10406);
and U10644 (N_10644,N_10437,N_10168);
nand U10645 (N_10645,N_10399,N_10218);
and U10646 (N_10646,N_10370,N_10335);
and U10647 (N_10647,N_10477,N_10286);
and U10648 (N_10648,N_10452,N_10360);
or U10649 (N_10649,N_10488,N_10272);
nand U10650 (N_10650,N_10261,N_10189);
or U10651 (N_10651,N_10085,N_10195);
or U10652 (N_10652,N_10246,N_10280);
xnor U10653 (N_10653,N_10165,N_10479);
nand U10654 (N_10654,N_10415,N_10432);
xnor U10655 (N_10655,N_10345,N_10252);
or U10656 (N_10656,N_10075,N_10187);
xnor U10657 (N_10657,N_10057,N_10180);
or U10658 (N_10658,N_10313,N_10172);
or U10659 (N_10659,N_10337,N_10460);
or U10660 (N_10660,N_10073,N_10062);
nand U10661 (N_10661,N_10005,N_10371);
and U10662 (N_10662,N_10495,N_10201);
nor U10663 (N_10663,N_10049,N_10444);
and U10664 (N_10664,N_10194,N_10393);
xnor U10665 (N_10665,N_10251,N_10250);
nand U10666 (N_10666,N_10325,N_10396);
nor U10667 (N_10667,N_10175,N_10311);
and U10668 (N_10668,N_10163,N_10341);
or U10669 (N_10669,N_10188,N_10120);
or U10670 (N_10670,N_10223,N_10205);
xor U10671 (N_10671,N_10482,N_10210);
nand U10672 (N_10672,N_10290,N_10381);
nor U10673 (N_10673,N_10463,N_10226);
nor U10674 (N_10674,N_10032,N_10332);
or U10675 (N_10675,N_10138,N_10082);
and U10676 (N_10676,N_10020,N_10025);
or U10677 (N_10677,N_10359,N_10042);
nor U10678 (N_10678,N_10065,N_10134);
nand U10679 (N_10679,N_10041,N_10184);
and U10680 (N_10680,N_10308,N_10092);
nand U10681 (N_10681,N_10267,N_10091);
or U10682 (N_10682,N_10192,N_10354);
or U10683 (N_10683,N_10298,N_10342);
xor U10684 (N_10684,N_10064,N_10008);
xor U10685 (N_10685,N_10258,N_10291);
nand U10686 (N_10686,N_10451,N_10254);
or U10687 (N_10687,N_10365,N_10409);
nand U10688 (N_10688,N_10177,N_10066);
or U10689 (N_10689,N_10224,N_10416);
or U10690 (N_10690,N_10480,N_10155);
and U10691 (N_10691,N_10070,N_10039);
nand U10692 (N_10692,N_10169,N_10369);
and U10693 (N_10693,N_10306,N_10429);
nand U10694 (N_10694,N_10408,N_10358);
and U10695 (N_10695,N_10216,N_10001);
and U10696 (N_10696,N_10423,N_10268);
and U10697 (N_10697,N_10378,N_10146);
and U10698 (N_10698,N_10324,N_10178);
nor U10699 (N_10699,N_10433,N_10214);
nand U10700 (N_10700,N_10126,N_10473);
xor U10701 (N_10701,N_10139,N_10388);
and U10702 (N_10702,N_10111,N_10288);
or U10703 (N_10703,N_10107,N_10400);
xor U10704 (N_10704,N_10203,N_10282);
and U10705 (N_10705,N_10196,N_10242);
or U10706 (N_10706,N_10322,N_10016);
and U10707 (N_10707,N_10069,N_10051);
xnor U10708 (N_10708,N_10271,N_10476);
xnor U10709 (N_10709,N_10048,N_10106);
nor U10710 (N_10710,N_10247,N_10367);
nand U10711 (N_10711,N_10449,N_10104);
nor U10712 (N_10712,N_10391,N_10348);
and U10713 (N_10713,N_10295,N_10323);
or U10714 (N_10714,N_10390,N_10109);
nor U10715 (N_10715,N_10405,N_10315);
and U10716 (N_10716,N_10260,N_10431);
xnor U10717 (N_10717,N_10362,N_10043);
nand U10718 (N_10718,N_10071,N_10148);
nor U10719 (N_10719,N_10011,N_10089);
or U10720 (N_10720,N_10375,N_10475);
or U10721 (N_10721,N_10472,N_10327);
or U10722 (N_10722,N_10102,N_10344);
nor U10723 (N_10723,N_10448,N_10086);
or U10724 (N_10724,N_10490,N_10364);
and U10725 (N_10725,N_10045,N_10384);
xor U10726 (N_10726,N_10219,N_10462);
nand U10727 (N_10727,N_10301,N_10115);
or U10728 (N_10728,N_10279,N_10119);
nand U10729 (N_10729,N_10465,N_10453);
and U10730 (N_10730,N_10232,N_10209);
or U10731 (N_10731,N_10392,N_10307);
or U10732 (N_10732,N_10018,N_10333);
or U10733 (N_10733,N_10081,N_10103);
or U10734 (N_10734,N_10424,N_10076);
nand U10735 (N_10735,N_10027,N_10054);
and U10736 (N_10736,N_10171,N_10181);
and U10737 (N_10737,N_10485,N_10426);
xnor U10738 (N_10738,N_10497,N_10321);
nand U10739 (N_10739,N_10009,N_10028);
or U10740 (N_10740,N_10346,N_10228);
or U10741 (N_10741,N_10053,N_10116);
and U10742 (N_10742,N_10149,N_10413);
and U10743 (N_10743,N_10029,N_10132);
nand U10744 (N_10744,N_10351,N_10374);
nand U10745 (N_10745,N_10127,N_10014);
or U10746 (N_10746,N_10352,N_10101);
or U10747 (N_10747,N_10304,N_10259);
and U10748 (N_10748,N_10207,N_10389);
nand U10749 (N_10749,N_10435,N_10263);
and U10750 (N_10750,N_10072,N_10492);
or U10751 (N_10751,N_10432,N_10276);
nand U10752 (N_10752,N_10450,N_10288);
or U10753 (N_10753,N_10492,N_10001);
xor U10754 (N_10754,N_10032,N_10487);
nand U10755 (N_10755,N_10317,N_10259);
nor U10756 (N_10756,N_10445,N_10282);
nand U10757 (N_10757,N_10200,N_10304);
or U10758 (N_10758,N_10016,N_10190);
nand U10759 (N_10759,N_10169,N_10244);
nor U10760 (N_10760,N_10058,N_10257);
and U10761 (N_10761,N_10351,N_10199);
nor U10762 (N_10762,N_10301,N_10493);
xor U10763 (N_10763,N_10454,N_10365);
nor U10764 (N_10764,N_10045,N_10309);
nand U10765 (N_10765,N_10038,N_10147);
or U10766 (N_10766,N_10194,N_10239);
nor U10767 (N_10767,N_10094,N_10491);
xnor U10768 (N_10768,N_10388,N_10186);
nand U10769 (N_10769,N_10227,N_10010);
or U10770 (N_10770,N_10487,N_10274);
nand U10771 (N_10771,N_10141,N_10123);
xor U10772 (N_10772,N_10379,N_10420);
xor U10773 (N_10773,N_10262,N_10039);
and U10774 (N_10774,N_10267,N_10467);
xnor U10775 (N_10775,N_10421,N_10313);
xnor U10776 (N_10776,N_10479,N_10393);
nor U10777 (N_10777,N_10235,N_10130);
xor U10778 (N_10778,N_10315,N_10158);
nor U10779 (N_10779,N_10136,N_10426);
nor U10780 (N_10780,N_10086,N_10355);
or U10781 (N_10781,N_10198,N_10010);
nor U10782 (N_10782,N_10201,N_10400);
nor U10783 (N_10783,N_10114,N_10239);
nand U10784 (N_10784,N_10129,N_10235);
nand U10785 (N_10785,N_10269,N_10411);
nand U10786 (N_10786,N_10030,N_10000);
and U10787 (N_10787,N_10114,N_10147);
or U10788 (N_10788,N_10164,N_10497);
nand U10789 (N_10789,N_10474,N_10019);
xnor U10790 (N_10790,N_10193,N_10468);
nand U10791 (N_10791,N_10394,N_10489);
xor U10792 (N_10792,N_10281,N_10016);
or U10793 (N_10793,N_10034,N_10499);
and U10794 (N_10794,N_10415,N_10345);
and U10795 (N_10795,N_10188,N_10117);
nand U10796 (N_10796,N_10363,N_10153);
nor U10797 (N_10797,N_10197,N_10307);
or U10798 (N_10798,N_10000,N_10130);
nand U10799 (N_10799,N_10106,N_10488);
xnor U10800 (N_10800,N_10034,N_10367);
or U10801 (N_10801,N_10352,N_10052);
nand U10802 (N_10802,N_10489,N_10411);
or U10803 (N_10803,N_10103,N_10147);
or U10804 (N_10804,N_10185,N_10116);
nor U10805 (N_10805,N_10476,N_10075);
xnor U10806 (N_10806,N_10343,N_10203);
nor U10807 (N_10807,N_10431,N_10038);
nand U10808 (N_10808,N_10227,N_10192);
xor U10809 (N_10809,N_10001,N_10390);
nand U10810 (N_10810,N_10073,N_10435);
or U10811 (N_10811,N_10288,N_10164);
xnor U10812 (N_10812,N_10377,N_10006);
or U10813 (N_10813,N_10493,N_10026);
or U10814 (N_10814,N_10124,N_10129);
nor U10815 (N_10815,N_10338,N_10224);
nor U10816 (N_10816,N_10020,N_10466);
and U10817 (N_10817,N_10056,N_10494);
nor U10818 (N_10818,N_10444,N_10342);
xnor U10819 (N_10819,N_10427,N_10054);
nand U10820 (N_10820,N_10263,N_10277);
nand U10821 (N_10821,N_10007,N_10022);
or U10822 (N_10822,N_10243,N_10129);
or U10823 (N_10823,N_10027,N_10312);
and U10824 (N_10824,N_10270,N_10228);
or U10825 (N_10825,N_10332,N_10091);
nor U10826 (N_10826,N_10009,N_10296);
or U10827 (N_10827,N_10089,N_10139);
xor U10828 (N_10828,N_10238,N_10345);
nand U10829 (N_10829,N_10065,N_10061);
or U10830 (N_10830,N_10483,N_10487);
nand U10831 (N_10831,N_10459,N_10020);
and U10832 (N_10832,N_10178,N_10261);
and U10833 (N_10833,N_10101,N_10481);
nor U10834 (N_10834,N_10208,N_10000);
or U10835 (N_10835,N_10118,N_10362);
xor U10836 (N_10836,N_10284,N_10291);
or U10837 (N_10837,N_10434,N_10053);
and U10838 (N_10838,N_10443,N_10424);
xor U10839 (N_10839,N_10244,N_10075);
and U10840 (N_10840,N_10069,N_10295);
and U10841 (N_10841,N_10069,N_10173);
and U10842 (N_10842,N_10165,N_10173);
or U10843 (N_10843,N_10173,N_10265);
and U10844 (N_10844,N_10390,N_10446);
nand U10845 (N_10845,N_10231,N_10114);
or U10846 (N_10846,N_10475,N_10261);
nand U10847 (N_10847,N_10197,N_10257);
xnor U10848 (N_10848,N_10260,N_10453);
xnor U10849 (N_10849,N_10156,N_10043);
xor U10850 (N_10850,N_10341,N_10401);
nand U10851 (N_10851,N_10024,N_10030);
or U10852 (N_10852,N_10406,N_10472);
and U10853 (N_10853,N_10222,N_10322);
and U10854 (N_10854,N_10007,N_10080);
and U10855 (N_10855,N_10280,N_10419);
nor U10856 (N_10856,N_10269,N_10396);
nor U10857 (N_10857,N_10336,N_10129);
and U10858 (N_10858,N_10276,N_10314);
xnor U10859 (N_10859,N_10306,N_10080);
nand U10860 (N_10860,N_10163,N_10385);
nand U10861 (N_10861,N_10169,N_10255);
nor U10862 (N_10862,N_10119,N_10185);
xor U10863 (N_10863,N_10144,N_10093);
or U10864 (N_10864,N_10160,N_10484);
or U10865 (N_10865,N_10462,N_10378);
nand U10866 (N_10866,N_10106,N_10204);
or U10867 (N_10867,N_10153,N_10471);
or U10868 (N_10868,N_10039,N_10112);
or U10869 (N_10869,N_10479,N_10024);
and U10870 (N_10870,N_10344,N_10425);
or U10871 (N_10871,N_10399,N_10385);
nand U10872 (N_10872,N_10494,N_10034);
or U10873 (N_10873,N_10284,N_10278);
and U10874 (N_10874,N_10052,N_10382);
xor U10875 (N_10875,N_10036,N_10285);
and U10876 (N_10876,N_10284,N_10346);
nand U10877 (N_10877,N_10358,N_10468);
and U10878 (N_10878,N_10285,N_10167);
xor U10879 (N_10879,N_10095,N_10011);
nand U10880 (N_10880,N_10168,N_10352);
and U10881 (N_10881,N_10140,N_10311);
or U10882 (N_10882,N_10104,N_10382);
nand U10883 (N_10883,N_10398,N_10086);
and U10884 (N_10884,N_10175,N_10085);
or U10885 (N_10885,N_10289,N_10186);
nand U10886 (N_10886,N_10452,N_10376);
nand U10887 (N_10887,N_10110,N_10045);
xor U10888 (N_10888,N_10208,N_10487);
or U10889 (N_10889,N_10041,N_10325);
and U10890 (N_10890,N_10195,N_10083);
nor U10891 (N_10891,N_10332,N_10100);
nor U10892 (N_10892,N_10308,N_10190);
nand U10893 (N_10893,N_10390,N_10197);
or U10894 (N_10894,N_10201,N_10259);
xnor U10895 (N_10895,N_10395,N_10090);
or U10896 (N_10896,N_10380,N_10102);
xor U10897 (N_10897,N_10056,N_10100);
nand U10898 (N_10898,N_10421,N_10090);
or U10899 (N_10899,N_10282,N_10433);
nor U10900 (N_10900,N_10266,N_10018);
nand U10901 (N_10901,N_10322,N_10023);
nor U10902 (N_10902,N_10069,N_10235);
or U10903 (N_10903,N_10264,N_10380);
nor U10904 (N_10904,N_10101,N_10232);
or U10905 (N_10905,N_10459,N_10336);
nor U10906 (N_10906,N_10287,N_10357);
and U10907 (N_10907,N_10154,N_10125);
xnor U10908 (N_10908,N_10184,N_10474);
nand U10909 (N_10909,N_10203,N_10046);
nor U10910 (N_10910,N_10067,N_10122);
xnor U10911 (N_10911,N_10199,N_10379);
xor U10912 (N_10912,N_10432,N_10042);
or U10913 (N_10913,N_10313,N_10053);
or U10914 (N_10914,N_10110,N_10090);
or U10915 (N_10915,N_10212,N_10096);
and U10916 (N_10916,N_10497,N_10328);
nor U10917 (N_10917,N_10304,N_10185);
xnor U10918 (N_10918,N_10244,N_10199);
nor U10919 (N_10919,N_10242,N_10282);
nand U10920 (N_10920,N_10387,N_10326);
nor U10921 (N_10921,N_10393,N_10219);
xor U10922 (N_10922,N_10415,N_10493);
and U10923 (N_10923,N_10465,N_10474);
nand U10924 (N_10924,N_10481,N_10200);
xnor U10925 (N_10925,N_10355,N_10128);
xnor U10926 (N_10926,N_10253,N_10230);
nor U10927 (N_10927,N_10215,N_10193);
or U10928 (N_10928,N_10288,N_10077);
or U10929 (N_10929,N_10247,N_10295);
xor U10930 (N_10930,N_10148,N_10467);
and U10931 (N_10931,N_10320,N_10470);
nand U10932 (N_10932,N_10483,N_10247);
nand U10933 (N_10933,N_10373,N_10221);
xor U10934 (N_10934,N_10407,N_10305);
or U10935 (N_10935,N_10493,N_10048);
xnor U10936 (N_10936,N_10461,N_10415);
and U10937 (N_10937,N_10398,N_10046);
nand U10938 (N_10938,N_10011,N_10179);
xor U10939 (N_10939,N_10204,N_10079);
nand U10940 (N_10940,N_10210,N_10199);
nor U10941 (N_10941,N_10068,N_10485);
or U10942 (N_10942,N_10362,N_10429);
nand U10943 (N_10943,N_10335,N_10012);
or U10944 (N_10944,N_10487,N_10198);
xor U10945 (N_10945,N_10028,N_10134);
and U10946 (N_10946,N_10342,N_10108);
and U10947 (N_10947,N_10181,N_10199);
nor U10948 (N_10948,N_10192,N_10240);
and U10949 (N_10949,N_10225,N_10440);
xnor U10950 (N_10950,N_10163,N_10049);
and U10951 (N_10951,N_10257,N_10386);
or U10952 (N_10952,N_10465,N_10482);
or U10953 (N_10953,N_10404,N_10015);
and U10954 (N_10954,N_10282,N_10133);
nor U10955 (N_10955,N_10038,N_10127);
and U10956 (N_10956,N_10103,N_10314);
xor U10957 (N_10957,N_10144,N_10155);
nor U10958 (N_10958,N_10206,N_10066);
nand U10959 (N_10959,N_10013,N_10260);
nor U10960 (N_10960,N_10152,N_10119);
xor U10961 (N_10961,N_10463,N_10364);
nor U10962 (N_10962,N_10173,N_10241);
nand U10963 (N_10963,N_10010,N_10011);
and U10964 (N_10964,N_10200,N_10323);
nand U10965 (N_10965,N_10273,N_10204);
nor U10966 (N_10966,N_10474,N_10352);
nor U10967 (N_10967,N_10496,N_10057);
and U10968 (N_10968,N_10334,N_10037);
nand U10969 (N_10969,N_10143,N_10316);
xnor U10970 (N_10970,N_10401,N_10022);
or U10971 (N_10971,N_10437,N_10435);
xor U10972 (N_10972,N_10464,N_10117);
and U10973 (N_10973,N_10012,N_10236);
and U10974 (N_10974,N_10083,N_10245);
xor U10975 (N_10975,N_10282,N_10221);
xnor U10976 (N_10976,N_10390,N_10408);
or U10977 (N_10977,N_10031,N_10088);
nand U10978 (N_10978,N_10170,N_10110);
xor U10979 (N_10979,N_10392,N_10263);
nand U10980 (N_10980,N_10176,N_10265);
or U10981 (N_10981,N_10067,N_10118);
or U10982 (N_10982,N_10280,N_10424);
xnor U10983 (N_10983,N_10269,N_10294);
xor U10984 (N_10984,N_10400,N_10237);
nand U10985 (N_10985,N_10253,N_10474);
nor U10986 (N_10986,N_10428,N_10317);
or U10987 (N_10987,N_10416,N_10321);
nand U10988 (N_10988,N_10171,N_10285);
nand U10989 (N_10989,N_10252,N_10407);
or U10990 (N_10990,N_10237,N_10362);
xor U10991 (N_10991,N_10255,N_10117);
nand U10992 (N_10992,N_10171,N_10084);
nor U10993 (N_10993,N_10289,N_10071);
or U10994 (N_10994,N_10424,N_10390);
and U10995 (N_10995,N_10152,N_10134);
xnor U10996 (N_10996,N_10497,N_10282);
nor U10997 (N_10997,N_10463,N_10294);
xnor U10998 (N_10998,N_10092,N_10020);
xnor U10999 (N_10999,N_10048,N_10007);
or U11000 (N_11000,N_10544,N_10518);
nor U11001 (N_11001,N_10675,N_10534);
xnor U11002 (N_11002,N_10709,N_10783);
xor U11003 (N_11003,N_10526,N_10761);
or U11004 (N_11004,N_10788,N_10991);
nand U11005 (N_11005,N_10842,N_10716);
nand U11006 (N_11006,N_10656,N_10921);
nand U11007 (N_11007,N_10803,N_10559);
and U11008 (N_11008,N_10732,N_10537);
xnor U11009 (N_11009,N_10851,N_10844);
nor U11010 (N_11010,N_10845,N_10624);
nand U11011 (N_11011,N_10952,N_10999);
and U11012 (N_11012,N_10976,N_10590);
or U11013 (N_11013,N_10517,N_10820);
and U11014 (N_11014,N_10830,N_10577);
and U11015 (N_11015,N_10507,N_10602);
or U11016 (N_11016,N_10661,N_10703);
nand U11017 (N_11017,N_10958,N_10752);
nand U11018 (N_11018,N_10785,N_10668);
nor U11019 (N_11019,N_10913,N_10635);
nor U11020 (N_11020,N_10569,N_10561);
xnor U11021 (N_11021,N_10598,N_10767);
and U11022 (N_11022,N_10794,N_10749);
or U11023 (N_11023,N_10897,N_10814);
nor U11024 (N_11024,N_10560,N_10657);
nand U11025 (N_11025,N_10941,N_10545);
nand U11026 (N_11026,N_10522,N_10562);
nand U11027 (N_11027,N_10521,N_10688);
and U11028 (N_11028,N_10935,N_10950);
or U11029 (N_11029,N_10692,N_10622);
nor U11030 (N_11030,N_10715,N_10736);
and U11031 (N_11031,N_10601,N_10887);
xor U11032 (N_11032,N_10748,N_10707);
nor U11033 (N_11033,N_10972,N_10503);
and U11034 (N_11034,N_10813,N_10939);
or U11035 (N_11035,N_10835,N_10850);
xnor U11036 (N_11036,N_10588,N_10604);
or U11037 (N_11037,N_10556,N_10875);
nor U11038 (N_11038,N_10666,N_10697);
or U11039 (N_11039,N_10658,N_10874);
or U11040 (N_11040,N_10962,N_10937);
and U11041 (N_11041,N_10711,N_10961);
xnor U11042 (N_11042,N_10797,N_10878);
xor U11043 (N_11043,N_10691,N_10873);
and U11044 (N_11044,N_10880,N_10584);
or U11045 (N_11045,N_10804,N_10547);
nor U11046 (N_11046,N_10502,N_10809);
nand U11047 (N_11047,N_10669,N_10791);
or U11048 (N_11048,N_10912,N_10772);
nor U11049 (N_11049,N_10571,N_10539);
or U11050 (N_11050,N_10860,N_10753);
nand U11051 (N_11051,N_10506,N_10895);
nand U11052 (N_11052,N_10701,N_10846);
nand U11053 (N_11053,N_10828,N_10726);
and U11054 (N_11054,N_10898,N_10513);
nor U11055 (N_11055,N_10725,N_10595);
or U11056 (N_11056,N_10970,N_10805);
nor U11057 (N_11057,N_10699,N_10867);
xor U11058 (N_11058,N_10642,N_10731);
and U11059 (N_11059,N_10535,N_10740);
and U11060 (N_11060,N_10869,N_10672);
or U11061 (N_11061,N_10865,N_10536);
or U11062 (N_11062,N_10923,N_10645);
and U11063 (N_11063,N_10784,N_10552);
nor U11064 (N_11064,N_10501,N_10766);
xnor U11065 (N_11065,N_10824,N_10712);
and U11066 (N_11066,N_10574,N_10826);
xor U11067 (N_11067,N_10829,N_10891);
nand U11068 (N_11068,N_10841,N_10614);
or U11069 (N_11069,N_10583,N_10723);
xor U11070 (N_11070,N_10557,N_10930);
xor U11071 (N_11071,N_10558,N_10581);
and U11072 (N_11072,N_10925,N_10837);
nor U11073 (N_11073,N_10884,N_10667);
xnor U11074 (N_11074,N_10644,N_10985);
nand U11075 (N_11075,N_10965,N_10633);
nor U11076 (N_11076,N_10670,N_10983);
nand U11077 (N_11077,N_10717,N_10782);
nand U11078 (N_11078,N_10881,N_10730);
xor U11079 (N_11079,N_10765,N_10567);
or U11080 (N_11080,N_10529,N_10954);
and U11081 (N_11081,N_10647,N_10918);
or U11082 (N_11082,N_10949,N_10959);
nand U11083 (N_11083,N_10682,N_10568);
or U11084 (N_11084,N_10612,N_10678);
xor U11085 (N_11085,N_10754,N_10515);
nor U11086 (N_11086,N_10902,N_10987);
xor U11087 (N_11087,N_10589,N_10505);
xnor U11088 (N_11088,N_10889,N_10508);
or U11089 (N_11089,N_10609,N_10825);
nand U11090 (N_11090,N_10755,N_10735);
nand U11091 (N_11091,N_10836,N_10997);
xor U11092 (N_11092,N_10945,N_10566);
and U11093 (N_11093,N_10579,N_10606);
nand U11094 (N_11094,N_10907,N_10621);
or U11095 (N_11095,N_10582,N_10947);
nand U11096 (N_11096,N_10808,N_10676);
and U11097 (N_11097,N_10674,N_10759);
xor U11098 (N_11098,N_10839,N_10751);
nor U11099 (N_11099,N_10951,N_10871);
nor U11100 (N_11100,N_10520,N_10911);
and U11101 (N_11101,N_10655,N_10650);
nand U11102 (N_11102,N_10696,N_10741);
nor U11103 (N_11103,N_10756,N_10704);
and U11104 (N_11104,N_10768,N_10802);
or U11105 (N_11105,N_10969,N_10861);
nand U11106 (N_11106,N_10806,N_10597);
nor U11107 (N_11107,N_10946,N_10989);
nor U11108 (N_11108,N_10774,N_10868);
nor U11109 (N_11109,N_10863,N_10700);
nand U11110 (N_11110,N_10553,N_10827);
and U11111 (N_11111,N_10527,N_10948);
or U11112 (N_11112,N_10617,N_10660);
or U11113 (N_11113,N_10819,N_10587);
nand U11114 (N_11114,N_10710,N_10936);
nand U11115 (N_11115,N_10996,N_10663);
xnor U11116 (N_11116,N_10719,N_10885);
xnor U11117 (N_11117,N_10616,N_10928);
nor U11118 (N_11118,N_10888,N_10720);
xnor U11119 (N_11119,N_10575,N_10580);
and U11120 (N_11120,N_10840,N_10714);
xnor U11121 (N_11121,N_10778,N_10528);
nor U11122 (N_11122,N_10649,N_10510);
nor U11123 (N_11123,N_10570,N_10611);
nand U11124 (N_11124,N_10833,N_10738);
xor U11125 (N_11125,N_10630,N_10746);
and U11126 (N_11126,N_10857,N_10931);
nand U11127 (N_11127,N_10817,N_10743);
or U11128 (N_11128,N_10648,N_10876);
nor U11129 (N_11129,N_10866,N_10920);
xor U11130 (N_11130,N_10773,N_10727);
and U11131 (N_11131,N_10932,N_10903);
nand U11132 (N_11132,N_10653,N_10810);
and U11133 (N_11133,N_10685,N_10705);
xnor U11134 (N_11134,N_10733,N_10563);
nand U11135 (N_11135,N_10593,N_10693);
xnor U11136 (N_11136,N_10780,N_10679);
nor U11137 (N_11137,N_10728,N_10943);
nand U11138 (N_11138,N_10821,N_10713);
or U11139 (N_11139,N_10524,N_10540);
or U11140 (N_11140,N_10793,N_10525);
and U11141 (N_11141,N_10734,N_10615);
nand U11142 (N_11142,N_10718,N_10516);
and U11143 (N_11143,N_10629,N_10893);
xor U11144 (N_11144,N_10838,N_10599);
nand U11145 (N_11145,N_10512,N_10573);
nand U11146 (N_11146,N_10769,N_10900);
and U11147 (N_11147,N_10790,N_10994);
xnor U11148 (N_11148,N_10671,N_10906);
xnor U11149 (N_11149,N_10933,N_10905);
xor U11150 (N_11150,N_10823,N_10998);
nor U11151 (N_11151,N_10538,N_10681);
nor U11152 (N_11152,N_10684,N_10600);
and U11153 (N_11153,N_10654,N_10729);
xor U11154 (N_11154,N_10781,N_10631);
xnor U11155 (N_11155,N_10957,N_10555);
or U11156 (N_11156,N_10690,N_10694);
or U11157 (N_11157,N_10807,N_10974);
nor U11158 (N_11158,N_10523,N_10564);
nand U11159 (N_11159,N_10585,N_10548);
and U11160 (N_11160,N_10944,N_10971);
nor U11161 (N_11161,N_10576,N_10980);
and U11162 (N_11162,N_10942,N_10739);
or U11163 (N_11163,N_10984,N_10855);
xor U11164 (N_11164,N_10742,N_10618);
xnor U11165 (N_11165,N_10779,N_10924);
nor U11166 (N_11166,N_10532,N_10908);
xnor U11167 (N_11167,N_10993,N_10812);
nand U11168 (N_11168,N_10721,N_10637);
xnor U11169 (N_11169,N_10990,N_10964);
and U11170 (N_11170,N_10687,N_10610);
or U11171 (N_11171,N_10886,N_10916);
or U11172 (N_11172,N_10745,N_10665);
and U11173 (N_11173,N_10787,N_10776);
and U11174 (N_11174,N_10982,N_10892);
nor U11175 (N_11175,N_10822,N_10632);
and U11176 (N_11176,N_10973,N_10659);
xnor U11177 (N_11177,N_10695,N_10914);
and U11178 (N_11178,N_10750,N_10757);
xnor U11179 (N_11179,N_10771,N_10511);
or U11180 (N_11180,N_10634,N_10963);
nor U11181 (N_11181,N_10799,N_10883);
or U11182 (N_11182,N_10966,N_10834);
or U11183 (N_11183,N_10641,N_10901);
and U11184 (N_11184,N_10550,N_10977);
or U11185 (N_11185,N_10968,N_10549);
or U11186 (N_11186,N_10981,N_10764);
xnor U11187 (N_11187,N_10992,N_10796);
and U11188 (N_11188,N_10636,N_10722);
and U11189 (N_11189,N_10986,N_10724);
or U11190 (N_11190,N_10546,N_10879);
nor U11191 (N_11191,N_10603,N_10504);
or U11192 (N_11192,N_10975,N_10514);
or U11193 (N_11193,N_10698,N_10619);
or U11194 (N_11194,N_10929,N_10533);
nand U11195 (N_11195,N_10843,N_10763);
or U11196 (N_11196,N_10858,N_10909);
xor U11197 (N_11197,N_10651,N_10708);
and U11198 (N_11198,N_10770,N_10862);
nand U11199 (N_11199,N_10530,N_10775);
or U11200 (N_11200,N_10628,N_10565);
or U11201 (N_11201,N_10852,N_10683);
and U11202 (N_11202,N_10554,N_10816);
and U11203 (N_11203,N_10919,N_10953);
or U11204 (N_11204,N_10859,N_10531);
or U11205 (N_11205,N_10847,N_10922);
nand U11206 (N_11206,N_10686,N_10811);
xnor U11207 (N_11207,N_10967,N_10872);
nand U11208 (N_11208,N_10896,N_10940);
nor U11209 (N_11209,N_10758,N_10664);
nand U11210 (N_11210,N_10652,N_10543);
nor U11211 (N_11211,N_10762,N_10917);
nor U11212 (N_11212,N_10638,N_10934);
or U11213 (N_11213,N_10623,N_10572);
nor U11214 (N_11214,N_10801,N_10702);
nand U11215 (N_11215,N_10927,N_10578);
and U11216 (N_11216,N_10643,N_10586);
nand U11217 (N_11217,N_10856,N_10795);
xnor U11218 (N_11218,N_10747,N_10864);
and U11219 (N_11219,N_10870,N_10995);
nand U11220 (N_11220,N_10910,N_10853);
nand U11221 (N_11221,N_10798,N_10894);
and U11222 (N_11222,N_10689,N_10815);
or U11223 (N_11223,N_10646,N_10832);
and U11224 (N_11224,N_10960,N_10542);
nor U11225 (N_11225,N_10744,N_10737);
and U11226 (N_11226,N_10662,N_10509);
xnor U11227 (N_11227,N_10608,N_10613);
xnor U11228 (N_11228,N_10988,N_10789);
nor U11229 (N_11229,N_10890,N_10673);
or U11230 (N_11230,N_10607,N_10500);
nand U11231 (N_11231,N_10854,N_10541);
or U11232 (N_11232,N_10979,N_10760);
or U11233 (N_11233,N_10605,N_10620);
nand U11234 (N_11234,N_10904,N_10849);
or U11235 (N_11235,N_10792,N_10831);
nor U11236 (N_11236,N_10818,N_10938);
or U11237 (N_11237,N_10955,N_10596);
nand U11238 (N_11238,N_10956,N_10680);
or U11239 (N_11239,N_10625,N_10677);
nand U11240 (N_11240,N_10626,N_10640);
nand U11241 (N_11241,N_10706,N_10592);
xor U11242 (N_11242,N_10519,N_10848);
and U11243 (N_11243,N_10551,N_10915);
nand U11244 (N_11244,N_10627,N_10899);
nand U11245 (N_11245,N_10877,N_10594);
or U11246 (N_11246,N_10882,N_10786);
and U11247 (N_11247,N_10591,N_10978);
and U11248 (N_11248,N_10639,N_10926);
nand U11249 (N_11249,N_10777,N_10800);
nor U11250 (N_11250,N_10581,N_10915);
xnor U11251 (N_11251,N_10575,N_10593);
nand U11252 (N_11252,N_10803,N_10910);
nor U11253 (N_11253,N_10535,N_10738);
nor U11254 (N_11254,N_10706,N_10579);
and U11255 (N_11255,N_10891,N_10828);
nor U11256 (N_11256,N_10558,N_10670);
xnor U11257 (N_11257,N_10810,N_10899);
and U11258 (N_11258,N_10808,N_10627);
nor U11259 (N_11259,N_10824,N_10897);
nand U11260 (N_11260,N_10840,N_10823);
xor U11261 (N_11261,N_10717,N_10549);
nand U11262 (N_11262,N_10832,N_10882);
nor U11263 (N_11263,N_10589,N_10607);
nor U11264 (N_11264,N_10723,N_10828);
nor U11265 (N_11265,N_10614,N_10929);
nand U11266 (N_11266,N_10513,N_10781);
and U11267 (N_11267,N_10590,N_10513);
or U11268 (N_11268,N_10661,N_10774);
nor U11269 (N_11269,N_10778,N_10800);
or U11270 (N_11270,N_10715,N_10917);
and U11271 (N_11271,N_10895,N_10715);
or U11272 (N_11272,N_10641,N_10745);
nand U11273 (N_11273,N_10745,N_10602);
nor U11274 (N_11274,N_10550,N_10790);
xnor U11275 (N_11275,N_10706,N_10728);
and U11276 (N_11276,N_10812,N_10841);
nor U11277 (N_11277,N_10797,N_10583);
nor U11278 (N_11278,N_10525,N_10775);
xnor U11279 (N_11279,N_10933,N_10554);
nor U11280 (N_11280,N_10614,N_10504);
nor U11281 (N_11281,N_10950,N_10836);
nand U11282 (N_11282,N_10809,N_10579);
nor U11283 (N_11283,N_10942,N_10784);
nand U11284 (N_11284,N_10886,N_10642);
xor U11285 (N_11285,N_10944,N_10697);
and U11286 (N_11286,N_10836,N_10899);
nand U11287 (N_11287,N_10766,N_10772);
or U11288 (N_11288,N_10734,N_10908);
nand U11289 (N_11289,N_10991,N_10736);
and U11290 (N_11290,N_10718,N_10944);
nor U11291 (N_11291,N_10644,N_10665);
nand U11292 (N_11292,N_10725,N_10795);
nor U11293 (N_11293,N_10900,N_10766);
or U11294 (N_11294,N_10902,N_10919);
and U11295 (N_11295,N_10500,N_10758);
nand U11296 (N_11296,N_10518,N_10711);
nand U11297 (N_11297,N_10725,N_10690);
and U11298 (N_11298,N_10568,N_10869);
xor U11299 (N_11299,N_10654,N_10500);
nor U11300 (N_11300,N_10513,N_10593);
nand U11301 (N_11301,N_10878,N_10712);
nor U11302 (N_11302,N_10915,N_10821);
or U11303 (N_11303,N_10611,N_10741);
and U11304 (N_11304,N_10756,N_10923);
nor U11305 (N_11305,N_10994,N_10857);
or U11306 (N_11306,N_10534,N_10799);
xor U11307 (N_11307,N_10677,N_10590);
nor U11308 (N_11308,N_10627,N_10584);
xnor U11309 (N_11309,N_10539,N_10894);
nand U11310 (N_11310,N_10802,N_10838);
and U11311 (N_11311,N_10907,N_10709);
nand U11312 (N_11312,N_10771,N_10663);
xnor U11313 (N_11313,N_10615,N_10533);
nand U11314 (N_11314,N_10905,N_10966);
nand U11315 (N_11315,N_10905,N_10522);
or U11316 (N_11316,N_10609,N_10897);
and U11317 (N_11317,N_10868,N_10788);
nor U11318 (N_11318,N_10797,N_10858);
nor U11319 (N_11319,N_10920,N_10773);
xor U11320 (N_11320,N_10988,N_10636);
nand U11321 (N_11321,N_10613,N_10862);
or U11322 (N_11322,N_10965,N_10658);
or U11323 (N_11323,N_10683,N_10689);
xnor U11324 (N_11324,N_10700,N_10593);
nor U11325 (N_11325,N_10814,N_10504);
nand U11326 (N_11326,N_10853,N_10850);
or U11327 (N_11327,N_10726,N_10770);
nor U11328 (N_11328,N_10623,N_10560);
or U11329 (N_11329,N_10802,N_10732);
nor U11330 (N_11330,N_10882,N_10558);
or U11331 (N_11331,N_10643,N_10951);
and U11332 (N_11332,N_10789,N_10745);
xor U11333 (N_11333,N_10762,N_10603);
nand U11334 (N_11334,N_10798,N_10928);
or U11335 (N_11335,N_10927,N_10852);
xor U11336 (N_11336,N_10973,N_10641);
nand U11337 (N_11337,N_10932,N_10502);
nand U11338 (N_11338,N_10683,N_10890);
xor U11339 (N_11339,N_10741,N_10634);
or U11340 (N_11340,N_10714,N_10943);
or U11341 (N_11341,N_10926,N_10787);
and U11342 (N_11342,N_10919,N_10778);
or U11343 (N_11343,N_10625,N_10988);
or U11344 (N_11344,N_10594,N_10507);
nor U11345 (N_11345,N_10579,N_10593);
nand U11346 (N_11346,N_10742,N_10872);
and U11347 (N_11347,N_10698,N_10733);
xnor U11348 (N_11348,N_10720,N_10764);
nor U11349 (N_11349,N_10779,N_10851);
nor U11350 (N_11350,N_10988,N_10814);
xor U11351 (N_11351,N_10781,N_10878);
or U11352 (N_11352,N_10973,N_10554);
xnor U11353 (N_11353,N_10728,N_10631);
or U11354 (N_11354,N_10616,N_10784);
nor U11355 (N_11355,N_10897,N_10575);
nor U11356 (N_11356,N_10686,N_10860);
nor U11357 (N_11357,N_10828,N_10832);
nor U11358 (N_11358,N_10987,N_10523);
xnor U11359 (N_11359,N_10602,N_10730);
nand U11360 (N_11360,N_10771,N_10626);
nand U11361 (N_11361,N_10953,N_10546);
xor U11362 (N_11362,N_10753,N_10743);
nor U11363 (N_11363,N_10806,N_10858);
nand U11364 (N_11364,N_10792,N_10639);
nand U11365 (N_11365,N_10624,N_10731);
nand U11366 (N_11366,N_10669,N_10516);
nand U11367 (N_11367,N_10993,N_10906);
nand U11368 (N_11368,N_10799,N_10824);
xor U11369 (N_11369,N_10611,N_10703);
nor U11370 (N_11370,N_10672,N_10692);
nor U11371 (N_11371,N_10902,N_10837);
nand U11372 (N_11372,N_10989,N_10938);
or U11373 (N_11373,N_10565,N_10752);
xnor U11374 (N_11374,N_10581,N_10838);
xor U11375 (N_11375,N_10786,N_10753);
or U11376 (N_11376,N_10691,N_10733);
or U11377 (N_11377,N_10926,N_10930);
nor U11378 (N_11378,N_10882,N_10518);
or U11379 (N_11379,N_10700,N_10661);
nand U11380 (N_11380,N_10509,N_10872);
xnor U11381 (N_11381,N_10685,N_10510);
xor U11382 (N_11382,N_10872,N_10558);
and U11383 (N_11383,N_10610,N_10516);
and U11384 (N_11384,N_10567,N_10934);
xor U11385 (N_11385,N_10621,N_10873);
nor U11386 (N_11386,N_10680,N_10775);
nand U11387 (N_11387,N_10981,N_10902);
or U11388 (N_11388,N_10560,N_10690);
xnor U11389 (N_11389,N_10689,N_10552);
or U11390 (N_11390,N_10624,N_10923);
nand U11391 (N_11391,N_10727,N_10565);
xnor U11392 (N_11392,N_10877,N_10854);
nand U11393 (N_11393,N_10767,N_10939);
nor U11394 (N_11394,N_10998,N_10856);
or U11395 (N_11395,N_10771,N_10904);
or U11396 (N_11396,N_10945,N_10932);
nand U11397 (N_11397,N_10570,N_10988);
and U11398 (N_11398,N_10920,N_10593);
and U11399 (N_11399,N_10622,N_10893);
nand U11400 (N_11400,N_10521,N_10587);
or U11401 (N_11401,N_10757,N_10892);
nand U11402 (N_11402,N_10772,N_10858);
nand U11403 (N_11403,N_10725,N_10502);
nor U11404 (N_11404,N_10501,N_10614);
nor U11405 (N_11405,N_10545,N_10971);
nand U11406 (N_11406,N_10657,N_10645);
and U11407 (N_11407,N_10646,N_10771);
nand U11408 (N_11408,N_10881,N_10726);
nand U11409 (N_11409,N_10622,N_10882);
and U11410 (N_11410,N_10557,N_10704);
xnor U11411 (N_11411,N_10576,N_10687);
xnor U11412 (N_11412,N_10594,N_10772);
xor U11413 (N_11413,N_10631,N_10588);
or U11414 (N_11414,N_10749,N_10985);
and U11415 (N_11415,N_10855,N_10779);
and U11416 (N_11416,N_10603,N_10911);
nand U11417 (N_11417,N_10755,N_10977);
xnor U11418 (N_11418,N_10973,N_10752);
xor U11419 (N_11419,N_10532,N_10698);
and U11420 (N_11420,N_10729,N_10710);
or U11421 (N_11421,N_10519,N_10615);
xnor U11422 (N_11422,N_10991,N_10787);
and U11423 (N_11423,N_10997,N_10826);
xnor U11424 (N_11424,N_10779,N_10743);
nand U11425 (N_11425,N_10702,N_10984);
or U11426 (N_11426,N_10980,N_10716);
nor U11427 (N_11427,N_10848,N_10534);
or U11428 (N_11428,N_10553,N_10823);
nor U11429 (N_11429,N_10918,N_10868);
nor U11430 (N_11430,N_10846,N_10811);
or U11431 (N_11431,N_10626,N_10842);
nor U11432 (N_11432,N_10679,N_10531);
or U11433 (N_11433,N_10819,N_10605);
nand U11434 (N_11434,N_10879,N_10542);
xor U11435 (N_11435,N_10740,N_10622);
nand U11436 (N_11436,N_10884,N_10866);
and U11437 (N_11437,N_10651,N_10600);
and U11438 (N_11438,N_10830,N_10928);
nand U11439 (N_11439,N_10791,N_10859);
xnor U11440 (N_11440,N_10690,N_10740);
xor U11441 (N_11441,N_10705,N_10958);
nand U11442 (N_11442,N_10898,N_10966);
nor U11443 (N_11443,N_10577,N_10723);
xnor U11444 (N_11444,N_10705,N_10807);
nand U11445 (N_11445,N_10732,N_10592);
or U11446 (N_11446,N_10631,N_10953);
nand U11447 (N_11447,N_10720,N_10794);
or U11448 (N_11448,N_10769,N_10723);
or U11449 (N_11449,N_10552,N_10644);
nor U11450 (N_11450,N_10912,N_10765);
xor U11451 (N_11451,N_10861,N_10848);
and U11452 (N_11452,N_10658,N_10720);
nand U11453 (N_11453,N_10885,N_10516);
and U11454 (N_11454,N_10811,N_10871);
or U11455 (N_11455,N_10521,N_10669);
nor U11456 (N_11456,N_10760,N_10627);
xor U11457 (N_11457,N_10977,N_10743);
or U11458 (N_11458,N_10829,N_10509);
nor U11459 (N_11459,N_10725,N_10927);
xor U11460 (N_11460,N_10757,N_10734);
nor U11461 (N_11461,N_10564,N_10578);
nand U11462 (N_11462,N_10536,N_10609);
nor U11463 (N_11463,N_10804,N_10918);
nor U11464 (N_11464,N_10568,N_10603);
nor U11465 (N_11465,N_10630,N_10525);
and U11466 (N_11466,N_10573,N_10880);
xor U11467 (N_11467,N_10811,N_10972);
nor U11468 (N_11468,N_10597,N_10980);
and U11469 (N_11469,N_10654,N_10962);
and U11470 (N_11470,N_10942,N_10793);
nor U11471 (N_11471,N_10687,N_10996);
xnor U11472 (N_11472,N_10973,N_10975);
or U11473 (N_11473,N_10655,N_10851);
and U11474 (N_11474,N_10734,N_10564);
xor U11475 (N_11475,N_10945,N_10549);
nor U11476 (N_11476,N_10604,N_10809);
or U11477 (N_11477,N_10550,N_10676);
xnor U11478 (N_11478,N_10837,N_10728);
nor U11479 (N_11479,N_10750,N_10692);
or U11480 (N_11480,N_10777,N_10968);
xor U11481 (N_11481,N_10752,N_10630);
or U11482 (N_11482,N_10512,N_10706);
and U11483 (N_11483,N_10984,N_10691);
and U11484 (N_11484,N_10701,N_10774);
and U11485 (N_11485,N_10820,N_10584);
nand U11486 (N_11486,N_10941,N_10994);
or U11487 (N_11487,N_10577,N_10814);
nor U11488 (N_11488,N_10671,N_10635);
nand U11489 (N_11489,N_10509,N_10975);
or U11490 (N_11490,N_10631,N_10876);
xnor U11491 (N_11491,N_10559,N_10628);
or U11492 (N_11492,N_10588,N_10688);
xnor U11493 (N_11493,N_10580,N_10659);
xnor U11494 (N_11494,N_10833,N_10506);
or U11495 (N_11495,N_10645,N_10511);
and U11496 (N_11496,N_10750,N_10888);
or U11497 (N_11497,N_10606,N_10855);
or U11498 (N_11498,N_10595,N_10734);
nand U11499 (N_11499,N_10941,N_10895);
or U11500 (N_11500,N_11444,N_11399);
or U11501 (N_11501,N_11376,N_11092);
xnor U11502 (N_11502,N_11179,N_11169);
nand U11503 (N_11503,N_11039,N_11289);
and U11504 (N_11504,N_11372,N_11042);
nor U11505 (N_11505,N_11309,N_11240);
xor U11506 (N_11506,N_11493,N_11356);
and U11507 (N_11507,N_11362,N_11364);
or U11508 (N_11508,N_11074,N_11225);
nor U11509 (N_11509,N_11375,N_11165);
or U11510 (N_11510,N_11427,N_11438);
nor U11511 (N_11511,N_11084,N_11020);
xor U11512 (N_11512,N_11062,N_11175);
xor U11513 (N_11513,N_11473,N_11210);
or U11514 (N_11514,N_11170,N_11101);
or U11515 (N_11515,N_11048,N_11023);
nand U11516 (N_11516,N_11047,N_11344);
or U11517 (N_11517,N_11031,N_11328);
and U11518 (N_11518,N_11373,N_11318);
xor U11519 (N_11519,N_11100,N_11035);
or U11520 (N_11520,N_11283,N_11102);
xor U11521 (N_11521,N_11195,N_11063);
or U11522 (N_11522,N_11041,N_11491);
nand U11523 (N_11523,N_11198,N_11208);
nor U11524 (N_11524,N_11423,N_11296);
nor U11525 (N_11525,N_11260,N_11116);
or U11526 (N_11526,N_11290,N_11490);
and U11527 (N_11527,N_11275,N_11222);
or U11528 (N_11528,N_11486,N_11217);
xor U11529 (N_11529,N_11235,N_11163);
nand U11530 (N_11530,N_11361,N_11046);
or U11531 (N_11531,N_11032,N_11040);
nor U11532 (N_11532,N_11252,N_11440);
nand U11533 (N_11533,N_11176,N_11081);
xor U11534 (N_11534,N_11057,N_11347);
nand U11535 (N_11535,N_11434,N_11173);
or U11536 (N_11536,N_11371,N_11406);
nor U11537 (N_11537,N_11421,N_11410);
or U11538 (N_11538,N_11012,N_11397);
xor U11539 (N_11539,N_11124,N_11193);
xor U11540 (N_11540,N_11251,N_11369);
xor U11541 (N_11541,N_11295,N_11329);
nand U11542 (N_11542,N_11317,N_11201);
or U11543 (N_11543,N_11025,N_11182);
xor U11544 (N_11544,N_11013,N_11231);
xnor U11545 (N_11545,N_11332,N_11131);
nor U11546 (N_11546,N_11269,N_11481);
and U11547 (N_11547,N_11273,N_11326);
or U11548 (N_11548,N_11281,N_11130);
nor U11549 (N_11549,N_11096,N_11359);
nand U11550 (N_11550,N_11058,N_11321);
or U11551 (N_11551,N_11036,N_11226);
nand U11552 (N_11552,N_11072,N_11172);
nor U11553 (N_11553,N_11292,N_11327);
nor U11554 (N_11554,N_11016,N_11207);
nand U11555 (N_11555,N_11320,N_11188);
nor U11556 (N_11556,N_11097,N_11052);
nor U11557 (N_11557,N_11075,N_11301);
nand U11558 (N_11558,N_11064,N_11389);
xnor U11559 (N_11559,N_11370,N_11154);
nor U11560 (N_11560,N_11408,N_11133);
xnor U11561 (N_11561,N_11109,N_11139);
nand U11562 (N_11562,N_11211,N_11120);
xor U11563 (N_11563,N_11400,N_11028);
nor U11564 (N_11564,N_11108,N_11196);
xnor U11565 (N_11565,N_11387,N_11117);
or U11566 (N_11566,N_11460,N_11024);
xnor U11567 (N_11567,N_11349,N_11194);
nor U11568 (N_11568,N_11068,N_11443);
nor U11569 (N_11569,N_11302,N_11089);
nor U11570 (N_11570,N_11448,N_11246);
nor U11571 (N_11571,N_11299,N_11128);
or U11572 (N_11572,N_11396,N_11363);
and U11573 (N_11573,N_11294,N_11022);
and U11574 (N_11574,N_11417,N_11187);
xor U11575 (N_11575,N_11428,N_11266);
xor U11576 (N_11576,N_11069,N_11155);
xor U11577 (N_11577,N_11357,N_11243);
or U11578 (N_11578,N_11331,N_11355);
and U11579 (N_11579,N_11245,N_11232);
xor U11580 (N_11580,N_11303,N_11011);
nand U11581 (N_11581,N_11002,N_11216);
or U11582 (N_11582,N_11404,N_11488);
nor U11583 (N_11583,N_11077,N_11464);
xor U11584 (N_11584,N_11457,N_11336);
nor U11585 (N_11585,N_11287,N_11461);
or U11586 (N_11586,N_11066,N_11223);
and U11587 (N_11587,N_11190,N_11413);
or U11588 (N_11588,N_11038,N_11118);
xnor U11589 (N_11589,N_11265,N_11126);
xor U11590 (N_11590,N_11348,N_11095);
or U11591 (N_11591,N_11335,N_11484);
or U11592 (N_11592,N_11454,N_11242);
nor U11593 (N_11593,N_11153,N_11480);
or U11594 (N_11594,N_11307,N_11080);
or U11595 (N_11595,N_11119,N_11450);
or U11596 (N_11596,N_11430,N_11053);
nor U11597 (N_11597,N_11202,N_11380);
xnor U11598 (N_11598,N_11136,N_11293);
nand U11599 (N_11599,N_11026,N_11437);
nand U11600 (N_11600,N_11078,N_11090);
nand U11601 (N_11601,N_11112,N_11033);
nand U11602 (N_11602,N_11455,N_11414);
xor U11603 (N_11603,N_11221,N_11494);
nor U11604 (N_11604,N_11167,N_11435);
or U11605 (N_11605,N_11479,N_11489);
or U11606 (N_11606,N_11358,N_11142);
xnor U11607 (N_11607,N_11407,N_11487);
xor U11608 (N_11608,N_11073,N_11365);
and U11609 (N_11609,N_11360,N_11354);
xnor U11610 (N_11610,N_11151,N_11300);
and U11611 (N_11611,N_11247,N_11145);
or U11612 (N_11612,N_11498,N_11076);
nand U11613 (N_11613,N_11184,N_11227);
xor U11614 (N_11614,N_11267,N_11280);
nor U11615 (N_11615,N_11463,N_11168);
and U11616 (N_11616,N_11157,N_11459);
xor U11617 (N_11617,N_11254,N_11264);
nand U11618 (N_11618,N_11186,N_11496);
xor U11619 (N_11619,N_11277,N_11429);
and U11620 (N_11620,N_11271,N_11161);
xor U11621 (N_11621,N_11219,N_11099);
and U11622 (N_11622,N_11171,N_11367);
nor U11623 (N_11623,N_11409,N_11446);
or U11624 (N_11624,N_11432,N_11050);
and U11625 (N_11625,N_11156,N_11274);
nand U11626 (N_11626,N_11061,N_11451);
or U11627 (N_11627,N_11324,N_11418);
xnor U11628 (N_11628,N_11403,N_11341);
xor U11629 (N_11629,N_11000,N_11310);
xor U11630 (N_11630,N_11143,N_11453);
nand U11631 (N_11631,N_11149,N_11346);
nand U11632 (N_11632,N_11134,N_11070);
xnor U11633 (N_11633,N_11458,N_11044);
and U11634 (N_11634,N_11339,N_11060);
nor U11635 (N_11635,N_11441,N_11366);
xor U11636 (N_11636,N_11475,N_11088);
nor U11637 (N_11637,N_11113,N_11192);
nor U11638 (N_11638,N_11416,N_11314);
and U11639 (N_11639,N_11248,N_11056);
nand U11640 (N_11640,N_11268,N_11306);
nor U11641 (N_11641,N_11467,N_11010);
and U11642 (N_11642,N_11353,N_11449);
and U11643 (N_11643,N_11471,N_11278);
xnor U11644 (N_11644,N_11137,N_11148);
nor U11645 (N_11645,N_11497,N_11104);
and U11646 (N_11646,N_11021,N_11276);
nand U11647 (N_11647,N_11164,N_11203);
and U11648 (N_11648,N_11152,N_11158);
or U11649 (N_11649,N_11395,N_11350);
xor U11650 (N_11650,N_11378,N_11159);
and U11651 (N_11651,N_11174,N_11316);
or U11652 (N_11652,N_11470,N_11442);
or U11653 (N_11653,N_11334,N_11319);
nor U11654 (N_11654,N_11433,N_11018);
or U11655 (N_11655,N_11141,N_11495);
and U11656 (N_11656,N_11422,N_11272);
xnor U11657 (N_11657,N_11140,N_11083);
xnor U11658 (N_11658,N_11178,N_11049);
or U11659 (N_11659,N_11424,N_11313);
nand U11660 (N_11660,N_11391,N_11241);
nor U11661 (N_11661,N_11043,N_11055);
nor U11662 (N_11662,N_11412,N_11127);
nor U11663 (N_11663,N_11094,N_11146);
and U11664 (N_11664,N_11330,N_11037);
xor U11665 (N_11665,N_11233,N_11029);
or U11666 (N_11666,N_11425,N_11286);
and U11667 (N_11667,N_11087,N_11106);
nor U11668 (N_11668,N_11014,N_11114);
xor U11669 (N_11669,N_11253,N_11377);
xor U11670 (N_11670,N_11059,N_11415);
nor U11671 (N_11671,N_11462,N_11067);
nand U11672 (N_11672,N_11098,N_11311);
nor U11673 (N_11673,N_11345,N_11138);
xnor U11674 (N_11674,N_11304,N_11237);
or U11675 (N_11675,N_11282,N_11291);
nor U11676 (N_11676,N_11181,N_11250);
nor U11677 (N_11677,N_11436,N_11374);
nor U11678 (N_11678,N_11085,N_11122);
or U11679 (N_11679,N_11103,N_11419);
or U11680 (N_11680,N_11214,N_11107);
xor U11681 (N_11681,N_11015,N_11177);
and U11682 (N_11682,N_11238,N_11115);
nand U11683 (N_11683,N_11093,N_11006);
nor U11684 (N_11684,N_11343,N_11337);
and U11685 (N_11685,N_11185,N_11492);
or U11686 (N_11686,N_11401,N_11392);
and U11687 (N_11687,N_11009,N_11007);
nand U11688 (N_11688,N_11384,N_11477);
nand U11689 (N_11689,N_11259,N_11288);
or U11690 (N_11690,N_11166,N_11465);
nand U11691 (N_11691,N_11411,N_11205);
nor U11692 (N_11692,N_11447,N_11162);
nor U11693 (N_11693,N_11001,N_11228);
nor U11694 (N_11694,N_11382,N_11499);
or U11695 (N_11695,N_11466,N_11206);
xor U11696 (N_11696,N_11110,N_11004);
nand U11697 (N_11697,N_11308,N_11034);
nor U11698 (N_11698,N_11483,N_11255);
nand U11699 (N_11699,N_11398,N_11452);
and U11700 (N_11700,N_11394,N_11197);
nand U11701 (N_11701,N_11125,N_11469);
nand U11702 (N_11702,N_11215,N_11439);
or U11703 (N_11703,N_11017,N_11123);
nor U11704 (N_11704,N_11183,N_11297);
and U11705 (N_11705,N_11236,N_11209);
xor U11706 (N_11706,N_11144,N_11351);
xnor U11707 (N_11707,N_11474,N_11385);
or U11708 (N_11708,N_11390,N_11135);
or U11709 (N_11709,N_11426,N_11263);
nor U11710 (N_11710,N_11315,N_11132);
xor U11711 (N_11711,N_11340,N_11051);
and U11712 (N_11712,N_11325,N_11333);
nor U11713 (N_11713,N_11472,N_11019);
nand U11714 (N_11714,N_11005,N_11468);
nor U11715 (N_11715,N_11258,N_11147);
and U11716 (N_11716,N_11191,N_11342);
nor U11717 (N_11717,N_11244,N_11379);
nor U11718 (N_11718,N_11381,N_11402);
nor U11719 (N_11719,N_11082,N_11284);
or U11720 (N_11720,N_11305,N_11368);
nor U11721 (N_11721,N_11257,N_11388);
and U11722 (N_11722,N_11256,N_11249);
nand U11723 (N_11723,N_11003,N_11086);
xnor U11724 (N_11724,N_11199,N_11204);
nand U11725 (N_11725,N_11338,N_11230);
nor U11726 (N_11726,N_11111,N_11431);
and U11727 (N_11727,N_11445,N_11224);
and U11728 (N_11728,N_11352,N_11079);
or U11729 (N_11729,N_11129,N_11456);
nor U11730 (N_11730,N_11071,N_11234);
and U11731 (N_11731,N_11160,N_11189);
nor U11732 (N_11732,N_11239,N_11065);
or U11733 (N_11733,N_11279,N_11220);
or U11734 (N_11734,N_11405,N_11285);
nand U11735 (N_11735,N_11229,N_11323);
nand U11736 (N_11736,N_11180,N_11218);
or U11737 (N_11737,N_11478,N_11008);
nand U11738 (N_11738,N_11105,N_11485);
or U11739 (N_11739,N_11393,N_11045);
or U11740 (N_11740,N_11262,N_11261);
nor U11741 (N_11741,N_11150,N_11322);
xor U11742 (N_11742,N_11091,N_11420);
nand U11743 (N_11743,N_11200,N_11213);
xnor U11744 (N_11744,N_11386,N_11030);
and U11745 (N_11745,N_11312,N_11476);
or U11746 (N_11746,N_11298,N_11270);
nor U11747 (N_11747,N_11027,N_11482);
nor U11748 (N_11748,N_11383,N_11121);
nor U11749 (N_11749,N_11054,N_11212);
or U11750 (N_11750,N_11224,N_11074);
or U11751 (N_11751,N_11459,N_11100);
nor U11752 (N_11752,N_11300,N_11401);
and U11753 (N_11753,N_11353,N_11114);
nor U11754 (N_11754,N_11227,N_11448);
nand U11755 (N_11755,N_11309,N_11017);
nor U11756 (N_11756,N_11291,N_11014);
and U11757 (N_11757,N_11448,N_11241);
xor U11758 (N_11758,N_11465,N_11474);
nor U11759 (N_11759,N_11302,N_11248);
or U11760 (N_11760,N_11318,N_11251);
xnor U11761 (N_11761,N_11102,N_11153);
nor U11762 (N_11762,N_11288,N_11334);
or U11763 (N_11763,N_11086,N_11367);
or U11764 (N_11764,N_11261,N_11097);
and U11765 (N_11765,N_11314,N_11290);
and U11766 (N_11766,N_11125,N_11334);
and U11767 (N_11767,N_11008,N_11368);
and U11768 (N_11768,N_11040,N_11471);
xnor U11769 (N_11769,N_11110,N_11035);
nor U11770 (N_11770,N_11308,N_11275);
or U11771 (N_11771,N_11042,N_11420);
xnor U11772 (N_11772,N_11317,N_11179);
nand U11773 (N_11773,N_11415,N_11461);
and U11774 (N_11774,N_11308,N_11095);
xnor U11775 (N_11775,N_11437,N_11451);
xor U11776 (N_11776,N_11330,N_11434);
or U11777 (N_11777,N_11169,N_11494);
nor U11778 (N_11778,N_11358,N_11271);
or U11779 (N_11779,N_11104,N_11265);
xor U11780 (N_11780,N_11164,N_11287);
nand U11781 (N_11781,N_11194,N_11471);
nor U11782 (N_11782,N_11377,N_11301);
nand U11783 (N_11783,N_11318,N_11397);
xor U11784 (N_11784,N_11317,N_11134);
nand U11785 (N_11785,N_11256,N_11248);
nand U11786 (N_11786,N_11153,N_11203);
or U11787 (N_11787,N_11062,N_11401);
or U11788 (N_11788,N_11489,N_11336);
nor U11789 (N_11789,N_11285,N_11429);
nand U11790 (N_11790,N_11263,N_11058);
xor U11791 (N_11791,N_11374,N_11439);
nand U11792 (N_11792,N_11300,N_11176);
nor U11793 (N_11793,N_11071,N_11355);
or U11794 (N_11794,N_11102,N_11419);
nand U11795 (N_11795,N_11284,N_11150);
xor U11796 (N_11796,N_11066,N_11430);
xnor U11797 (N_11797,N_11187,N_11396);
xor U11798 (N_11798,N_11266,N_11425);
xnor U11799 (N_11799,N_11139,N_11310);
nor U11800 (N_11800,N_11320,N_11190);
nor U11801 (N_11801,N_11013,N_11342);
or U11802 (N_11802,N_11363,N_11149);
xor U11803 (N_11803,N_11397,N_11157);
nand U11804 (N_11804,N_11164,N_11350);
and U11805 (N_11805,N_11457,N_11275);
or U11806 (N_11806,N_11484,N_11277);
nor U11807 (N_11807,N_11077,N_11102);
nand U11808 (N_11808,N_11213,N_11334);
or U11809 (N_11809,N_11294,N_11305);
or U11810 (N_11810,N_11409,N_11113);
nor U11811 (N_11811,N_11422,N_11429);
and U11812 (N_11812,N_11056,N_11443);
xor U11813 (N_11813,N_11411,N_11437);
nor U11814 (N_11814,N_11067,N_11143);
nand U11815 (N_11815,N_11455,N_11163);
or U11816 (N_11816,N_11045,N_11376);
or U11817 (N_11817,N_11467,N_11090);
nand U11818 (N_11818,N_11351,N_11429);
nor U11819 (N_11819,N_11216,N_11414);
and U11820 (N_11820,N_11165,N_11188);
nor U11821 (N_11821,N_11104,N_11238);
nor U11822 (N_11822,N_11329,N_11029);
and U11823 (N_11823,N_11018,N_11012);
nand U11824 (N_11824,N_11001,N_11499);
nor U11825 (N_11825,N_11351,N_11357);
nor U11826 (N_11826,N_11208,N_11172);
xnor U11827 (N_11827,N_11492,N_11089);
nor U11828 (N_11828,N_11331,N_11202);
and U11829 (N_11829,N_11036,N_11165);
and U11830 (N_11830,N_11079,N_11282);
xor U11831 (N_11831,N_11051,N_11220);
xnor U11832 (N_11832,N_11008,N_11297);
xnor U11833 (N_11833,N_11071,N_11375);
xnor U11834 (N_11834,N_11083,N_11019);
nor U11835 (N_11835,N_11435,N_11284);
nand U11836 (N_11836,N_11259,N_11225);
nor U11837 (N_11837,N_11020,N_11148);
nand U11838 (N_11838,N_11023,N_11041);
nor U11839 (N_11839,N_11053,N_11027);
and U11840 (N_11840,N_11162,N_11021);
and U11841 (N_11841,N_11007,N_11415);
nor U11842 (N_11842,N_11335,N_11405);
or U11843 (N_11843,N_11136,N_11055);
nor U11844 (N_11844,N_11040,N_11248);
or U11845 (N_11845,N_11478,N_11456);
nand U11846 (N_11846,N_11362,N_11448);
nand U11847 (N_11847,N_11054,N_11137);
xor U11848 (N_11848,N_11366,N_11059);
and U11849 (N_11849,N_11185,N_11238);
and U11850 (N_11850,N_11427,N_11097);
and U11851 (N_11851,N_11172,N_11329);
and U11852 (N_11852,N_11071,N_11102);
or U11853 (N_11853,N_11316,N_11439);
nor U11854 (N_11854,N_11207,N_11171);
and U11855 (N_11855,N_11348,N_11210);
nand U11856 (N_11856,N_11442,N_11212);
xnor U11857 (N_11857,N_11446,N_11180);
nand U11858 (N_11858,N_11118,N_11206);
nor U11859 (N_11859,N_11143,N_11332);
nor U11860 (N_11860,N_11481,N_11056);
xor U11861 (N_11861,N_11270,N_11326);
xor U11862 (N_11862,N_11106,N_11234);
nor U11863 (N_11863,N_11442,N_11372);
xnor U11864 (N_11864,N_11302,N_11341);
xnor U11865 (N_11865,N_11063,N_11458);
nor U11866 (N_11866,N_11351,N_11440);
xor U11867 (N_11867,N_11009,N_11110);
xor U11868 (N_11868,N_11170,N_11113);
xnor U11869 (N_11869,N_11131,N_11275);
or U11870 (N_11870,N_11294,N_11465);
and U11871 (N_11871,N_11074,N_11024);
and U11872 (N_11872,N_11113,N_11252);
nand U11873 (N_11873,N_11453,N_11478);
nor U11874 (N_11874,N_11444,N_11307);
or U11875 (N_11875,N_11251,N_11435);
or U11876 (N_11876,N_11055,N_11433);
xor U11877 (N_11877,N_11320,N_11094);
xnor U11878 (N_11878,N_11145,N_11325);
nand U11879 (N_11879,N_11300,N_11345);
and U11880 (N_11880,N_11423,N_11411);
nor U11881 (N_11881,N_11054,N_11418);
or U11882 (N_11882,N_11017,N_11210);
nand U11883 (N_11883,N_11386,N_11181);
nand U11884 (N_11884,N_11044,N_11342);
xor U11885 (N_11885,N_11394,N_11363);
xnor U11886 (N_11886,N_11076,N_11337);
nand U11887 (N_11887,N_11254,N_11085);
and U11888 (N_11888,N_11115,N_11170);
xor U11889 (N_11889,N_11286,N_11494);
nor U11890 (N_11890,N_11333,N_11468);
nand U11891 (N_11891,N_11371,N_11179);
nand U11892 (N_11892,N_11144,N_11367);
nor U11893 (N_11893,N_11487,N_11484);
nor U11894 (N_11894,N_11236,N_11447);
xor U11895 (N_11895,N_11123,N_11301);
or U11896 (N_11896,N_11343,N_11294);
nor U11897 (N_11897,N_11096,N_11487);
nand U11898 (N_11898,N_11442,N_11181);
nand U11899 (N_11899,N_11282,N_11023);
or U11900 (N_11900,N_11351,N_11225);
or U11901 (N_11901,N_11475,N_11165);
nand U11902 (N_11902,N_11199,N_11430);
xor U11903 (N_11903,N_11356,N_11401);
nand U11904 (N_11904,N_11261,N_11212);
nand U11905 (N_11905,N_11341,N_11251);
nor U11906 (N_11906,N_11423,N_11361);
nor U11907 (N_11907,N_11043,N_11275);
or U11908 (N_11908,N_11318,N_11228);
or U11909 (N_11909,N_11038,N_11493);
and U11910 (N_11910,N_11113,N_11461);
and U11911 (N_11911,N_11170,N_11322);
nor U11912 (N_11912,N_11234,N_11264);
and U11913 (N_11913,N_11057,N_11351);
nand U11914 (N_11914,N_11317,N_11403);
and U11915 (N_11915,N_11255,N_11379);
xor U11916 (N_11916,N_11404,N_11436);
nor U11917 (N_11917,N_11474,N_11486);
and U11918 (N_11918,N_11350,N_11382);
or U11919 (N_11919,N_11005,N_11027);
or U11920 (N_11920,N_11449,N_11016);
or U11921 (N_11921,N_11386,N_11295);
nand U11922 (N_11922,N_11232,N_11027);
nor U11923 (N_11923,N_11474,N_11402);
nand U11924 (N_11924,N_11286,N_11337);
nand U11925 (N_11925,N_11293,N_11200);
or U11926 (N_11926,N_11095,N_11407);
xor U11927 (N_11927,N_11273,N_11176);
xnor U11928 (N_11928,N_11411,N_11323);
nand U11929 (N_11929,N_11351,N_11019);
and U11930 (N_11930,N_11099,N_11468);
or U11931 (N_11931,N_11419,N_11392);
nor U11932 (N_11932,N_11151,N_11083);
nor U11933 (N_11933,N_11141,N_11104);
nand U11934 (N_11934,N_11005,N_11163);
and U11935 (N_11935,N_11474,N_11322);
xor U11936 (N_11936,N_11250,N_11178);
or U11937 (N_11937,N_11073,N_11300);
and U11938 (N_11938,N_11142,N_11357);
nor U11939 (N_11939,N_11387,N_11271);
xor U11940 (N_11940,N_11466,N_11183);
nor U11941 (N_11941,N_11439,N_11491);
xnor U11942 (N_11942,N_11141,N_11044);
nor U11943 (N_11943,N_11025,N_11130);
xor U11944 (N_11944,N_11297,N_11113);
and U11945 (N_11945,N_11140,N_11269);
or U11946 (N_11946,N_11328,N_11493);
xnor U11947 (N_11947,N_11229,N_11215);
nor U11948 (N_11948,N_11112,N_11011);
or U11949 (N_11949,N_11211,N_11279);
or U11950 (N_11950,N_11256,N_11111);
and U11951 (N_11951,N_11452,N_11419);
nor U11952 (N_11952,N_11216,N_11019);
nor U11953 (N_11953,N_11150,N_11179);
or U11954 (N_11954,N_11438,N_11199);
nor U11955 (N_11955,N_11181,N_11404);
nor U11956 (N_11956,N_11191,N_11336);
nand U11957 (N_11957,N_11123,N_11243);
xor U11958 (N_11958,N_11230,N_11085);
xnor U11959 (N_11959,N_11080,N_11003);
nor U11960 (N_11960,N_11210,N_11009);
nand U11961 (N_11961,N_11155,N_11237);
xnor U11962 (N_11962,N_11310,N_11238);
and U11963 (N_11963,N_11344,N_11181);
nand U11964 (N_11964,N_11395,N_11225);
xnor U11965 (N_11965,N_11301,N_11260);
nand U11966 (N_11966,N_11347,N_11203);
xnor U11967 (N_11967,N_11350,N_11402);
or U11968 (N_11968,N_11083,N_11050);
xnor U11969 (N_11969,N_11456,N_11347);
nand U11970 (N_11970,N_11448,N_11335);
xor U11971 (N_11971,N_11413,N_11102);
or U11972 (N_11972,N_11202,N_11089);
xnor U11973 (N_11973,N_11343,N_11243);
and U11974 (N_11974,N_11350,N_11235);
xnor U11975 (N_11975,N_11245,N_11490);
or U11976 (N_11976,N_11071,N_11419);
and U11977 (N_11977,N_11430,N_11331);
xor U11978 (N_11978,N_11178,N_11100);
nand U11979 (N_11979,N_11042,N_11429);
nor U11980 (N_11980,N_11218,N_11234);
xnor U11981 (N_11981,N_11353,N_11137);
nand U11982 (N_11982,N_11146,N_11312);
or U11983 (N_11983,N_11198,N_11187);
nor U11984 (N_11984,N_11310,N_11017);
and U11985 (N_11985,N_11036,N_11345);
nand U11986 (N_11986,N_11092,N_11461);
and U11987 (N_11987,N_11302,N_11357);
xor U11988 (N_11988,N_11235,N_11482);
nand U11989 (N_11989,N_11479,N_11029);
nor U11990 (N_11990,N_11457,N_11422);
nor U11991 (N_11991,N_11255,N_11131);
and U11992 (N_11992,N_11122,N_11340);
and U11993 (N_11993,N_11424,N_11432);
xnor U11994 (N_11994,N_11362,N_11334);
and U11995 (N_11995,N_11400,N_11252);
xnor U11996 (N_11996,N_11099,N_11425);
xnor U11997 (N_11997,N_11408,N_11404);
xor U11998 (N_11998,N_11054,N_11241);
or U11999 (N_11999,N_11058,N_11245);
nand U12000 (N_12000,N_11846,N_11693);
or U12001 (N_12001,N_11764,N_11875);
xnor U12002 (N_12002,N_11997,N_11522);
nand U12003 (N_12003,N_11796,N_11829);
nor U12004 (N_12004,N_11832,N_11763);
nor U12005 (N_12005,N_11971,N_11586);
nand U12006 (N_12006,N_11789,N_11896);
or U12007 (N_12007,N_11739,N_11811);
nand U12008 (N_12008,N_11568,N_11767);
nor U12009 (N_12009,N_11514,N_11743);
and U12010 (N_12010,N_11857,N_11898);
or U12011 (N_12011,N_11707,N_11714);
and U12012 (N_12012,N_11918,N_11863);
and U12013 (N_12013,N_11631,N_11770);
nor U12014 (N_12014,N_11932,N_11625);
or U12015 (N_12015,N_11917,N_11603);
and U12016 (N_12016,N_11654,N_11798);
nand U12017 (N_12017,N_11604,N_11985);
xnor U12018 (N_12018,N_11843,N_11628);
nor U12019 (N_12019,N_11837,N_11675);
and U12020 (N_12020,N_11862,N_11884);
nand U12021 (N_12021,N_11508,N_11699);
nor U12022 (N_12022,N_11683,N_11825);
xnor U12023 (N_12023,N_11511,N_11548);
or U12024 (N_12024,N_11611,N_11874);
nand U12025 (N_12025,N_11519,N_11909);
nand U12026 (N_12026,N_11790,N_11733);
or U12027 (N_12027,N_11804,N_11830);
nor U12028 (N_12028,N_11742,N_11704);
nand U12029 (N_12029,N_11794,N_11945);
or U12030 (N_12030,N_11688,N_11622);
or U12031 (N_12031,N_11881,N_11694);
or U12032 (N_12032,N_11944,N_11686);
nand U12033 (N_12033,N_11878,N_11649);
nor U12034 (N_12034,N_11937,N_11600);
xor U12035 (N_12035,N_11934,N_11859);
nand U12036 (N_12036,N_11984,N_11954);
nor U12037 (N_12037,N_11561,N_11677);
and U12038 (N_12038,N_11847,N_11719);
nor U12039 (N_12039,N_11836,N_11721);
nand U12040 (N_12040,N_11953,N_11822);
xor U12041 (N_12041,N_11947,N_11506);
xnor U12042 (N_12042,N_11637,N_11941);
xnor U12043 (N_12043,N_11550,N_11692);
nand U12044 (N_12044,N_11834,N_11723);
nand U12045 (N_12045,N_11598,N_11988);
nand U12046 (N_12046,N_11907,N_11576);
or U12047 (N_12047,N_11538,N_11690);
xor U12048 (N_12048,N_11575,N_11865);
or U12049 (N_12049,N_11509,N_11980);
nand U12050 (N_12050,N_11957,N_11706);
nor U12051 (N_12051,N_11527,N_11933);
and U12052 (N_12052,N_11962,N_11546);
and U12053 (N_12053,N_11741,N_11620);
nor U12054 (N_12054,N_11793,N_11964);
nor U12055 (N_12055,N_11759,N_11726);
nand U12056 (N_12056,N_11608,N_11810);
nand U12057 (N_12057,N_11840,N_11579);
nor U12058 (N_12058,N_11752,N_11589);
nand U12059 (N_12059,N_11717,N_11872);
nand U12060 (N_12060,N_11922,N_11529);
or U12061 (N_12061,N_11670,N_11593);
and U12062 (N_12062,N_11766,N_11950);
xnor U12063 (N_12063,N_11588,N_11972);
nand U12064 (N_12064,N_11805,N_11607);
or U12065 (N_12065,N_11753,N_11657);
nand U12066 (N_12066,N_11663,N_11740);
nor U12067 (N_12067,N_11816,N_11510);
xnor U12068 (N_12068,N_11525,N_11563);
xnor U12069 (N_12069,N_11856,N_11578);
and U12070 (N_12070,N_11844,N_11999);
xnor U12071 (N_12071,N_11974,N_11720);
xnor U12072 (N_12072,N_11778,N_11786);
or U12073 (N_12073,N_11520,N_11700);
or U12074 (N_12074,N_11737,N_11574);
and U12075 (N_12075,N_11852,N_11919);
nor U12076 (N_12076,N_11921,N_11507);
or U12077 (N_12077,N_11813,N_11923);
xnor U12078 (N_12078,N_11940,N_11814);
or U12079 (N_12079,N_11512,N_11673);
and U12080 (N_12080,N_11781,N_11966);
nor U12081 (N_12081,N_11661,N_11774);
xor U12082 (N_12082,N_11685,N_11653);
xnor U12083 (N_12083,N_11768,N_11993);
nand U12084 (N_12084,N_11695,N_11827);
nand U12085 (N_12085,N_11587,N_11824);
or U12086 (N_12086,N_11869,N_11584);
nand U12087 (N_12087,N_11581,N_11687);
or U12088 (N_12088,N_11571,N_11927);
and U12089 (N_12089,N_11777,N_11833);
nand U12090 (N_12090,N_11744,N_11900);
nand U12091 (N_12091,N_11689,N_11523);
and U12092 (N_12092,N_11965,N_11889);
or U12093 (N_12093,N_11899,N_11638);
and U12094 (N_12094,N_11855,N_11864);
or U12095 (N_12095,N_11678,N_11986);
or U12096 (N_12096,N_11989,N_11903);
and U12097 (N_12097,N_11536,N_11783);
nand U12098 (N_12098,N_11926,N_11682);
and U12099 (N_12099,N_11949,N_11990);
nor U12100 (N_12100,N_11551,N_11658);
and U12101 (N_12101,N_11681,N_11967);
or U12102 (N_12102,N_11842,N_11738);
nor U12103 (N_12103,N_11644,N_11535);
and U12104 (N_12104,N_11925,N_11995);
xnor U12105 (N_12105,N_11596,N_11791);
xnor U12106 (N_12106,N_11616,N_11838);
nor U12107 (N_12107,N_11592,N_11652);
xnor U12108 (N_12108,N_11562,N_11861);
nor U12109 (N_12109,N_11614,N_11975);
nor U12110 (N_12110,N_11930,N_11991);
xor U12111 (N_12111,N_11951,N_11505);
or U12112 (N_12112,N_11660,N_11715);
nand U12113 (N_12113,N_11552,N_11787);
and U12114 (N_12114,N_11886,N_11959);
xor U12115 (N_12115,N_11711,N_11928);
xnor U12116 (N_12116,N_11817,N_11887);
xnor U12117 (N_12117,N_11569,N_11702);
xnor U12118 (N_12118,N_11913,N_11860);
xnor U12119 (N_12119,N_11888,N_11998);
or U12120 (N_12120,N_11877,N_11956);
xor U12121 (N_12121,N_11853,N_11710);
xor U12122 (N_12122,N_11976,N_11808);
or U12123 (N_12123,N_11803,N_11908);
xor U12124 (N_12124,N_11725,N_11996);
or U12125 (N_12125,N_11526,N_11590);
or U12126 (N_12126,N_11772,N_11606);
or U12127 (N_12127,N_11580,N_11601);
and U12128 (N_12128,N_11849,N_11758);
and U12129 (N_12129,N_11671,N_11797);
or U12130 (N_12130,N_11820,N_11792);
and U12131 (N_12131,N_11582,N_11724);
and U12132 (N_12132,N_11558,N_11835);
nor U12133 (N_12133,N_11553,N_11782);
and U12134 (N_12134,N_11655,N_11904);
xnor U12135 (N_12135,N_11615,N_11731);
nor U12136 (N_12136,N_11943,N_11573);
or U12137 (N_12137,N_11595,N_11503);
xor U12138 (N_12138,N_11528,N_11970);
nor U12139 (N_12139,N_11775,N_11848);
nand U12140 (N_12140,N_11708,N_11809);
or U12141 (N_12141,N_11754,N_11876);
or U12142 (N_12142,N_11916,N_11961);
and U12143 (N_12143,N_11597,N_11765);
nor U12144 (N_12144,N_11892,N_11769);
or U12145 (N_12145,N_11564,N_11987);
nor U12146 (N_12146,N_11531,N_11982);
nand U12147 (N_12147,N_11709,N_11559);
xnor U12148 (N_12148,N_11883,N_11659);
nand U12149 (N_12149,N_11524,N_11639);
and U12150 (N_12150,N_11749,N_11555);
or U12151 (N_12151,N_11539,N_11672);
or U12152 (N_12152,N_11910,N_11696);
and U12153 (N_12153,N_11968,N_11501);
xor U12154 (N_12154,N_11697,N_11946);
nand U12155 (N_12155,N_11599,N_11748);
xnor U12156 (N_12156,N_11679,N_11935);
and U12157 (N_12157,N_11634,N_11891);
nand U12158 (N_12158,N_11942,N_11823);
nand U12159 (N_12159,N_11839,N_11880);
nor U12160 (N_12160,N_11806,N_11668);
nand U12161 (N_12161,N_11978,N_11577);
and U12162 (N_12162,N_11969,N_11728);
nand U12163 (N_12163,N_11605,N_11610);
xnor U12164 (N_12164,N_11854,N_11554);
xnor U12165 (N_12165,N_11534,N_11669);
and U12166 (N_12166,N_11831,N_11648);
nor U12167 (N_12167,N_11958,N_11929);
xnor U12168 (N_12168,N_11801,N_11543);
nor U12169 (N_12169,N_11905,N_11756);
xor U12170 (N_12170,N_11641,N_11994);
xor U12171 (N_12171,N_11948,N_11650);
xor U12172 (N_12172,N_11585,N_11556);
and U12173 (N_12173,N_11627,N_11850);
xnor U12174 (N_12174,N_11931,N_11746);
nor U12175 (N_12175,N_11736,N_11936);
xnor U12176 (N_12176,N_11802,N_11828);
xnor U12177 (N_12177,N_11785,N_11979);
nand U12178 (N_12178,N_11537,N_11747);
nand U12179 (N_12179,N_11691,N_11541);
xnor U12180 (N_12180,N_11868,N_11807);
nand U12181 (N_12181,N_11504,N_11521);
or U12182 (N_12182,N_11845,N_11533);
nor U12183 (N_12183,N_11780,N_11776);
nand U12184 (N_12184,N_11915,N_11665);
xnor U12185 (N_12185,N_11762,N_11788);
or U12186 (N_12186,N_11549,N_11799);
and U12187 (N_12187,N_11647,N_11515);
xor U12188 (N_12188,N_11684,N_11635);
nand U12189 (N_12189,N_11906,N_11981);
xor U12190 (N_12190,N_11819,N_11732);
nor U12191 (N_12191,N_11664,N_11730);
nand U12192 (N_12192,N_11713,N_11895);
nor U12193 (N_12193,N_11680,N_11705);
xor U12194 (N_12194,N_11897,N_11722);
nand U12195 (N_12195,N_11885,N_11609);
nand U12196 (N_12196,N_11977,N_11729);
xnor U12197 (N_12197,N_11745,N_11646);
nor U12198 (N_12198,N_11674,N_11757);
or U12199 (N_12199,N_11866,N_11911);
or U12200 (N_12200,N_11651,N_11602);
xnor U12201 (N_12201,N_11901,N_11626);
nand U12202 (N_12202,N_11619,N_11914);
or U12203 (N_12203,N_11902,N_11858);
xnor U12204 (N_12204,N_11516,N_11502);
and U12205 (N_12205,N_11773,N_11924);
and U12206 (N_12206,N_11662,N_11718);
nor U12207 (N_12207,N_11643,N_11667);
or U12208 (N_12208,N_11735,N_11795);
nand U12209 (N_12209,N_11612,N_11629);
nand U12210 (N_12210,N_11530,N_11815);
nand U12211 (N_12211,N_11821,N_11955);
or U12212 (N_12212,N_11560,N_11545);
nor U12213 (N_12213,N_11751,N_11779);
and U12214 (N_12214,N_11500,N_11542);
xor U12215 (N_12215,N_11618,N_11939);
nor U12216 (N_12216,N_11557,N_11621);
and U12217 (N_12217,N_11882,N_11565);
or U12218 (N_12218,N_11952,N_11879);
nand U12219 (N_12219,N_11963,N_11624);
xnor U12220 (N_12220,N_11890,N_11812);
or U12221 (N_12221,N_11656,N_11912);
nor U12222 (N_12222,N_11760,N_11666);
or U12223 (N_12223,N_11701,N_11566);
and U12224 (N_12224,N_11517,N_11960);
nand U12225 (N_12225,N_11518,N_11703);
nor U12226 (N_12226,N_11867,N_11645);
nand U12227 (N_12227,N_11642,N_11633);
or U12228 (N_12228,N_11870,N_11873);
and U12229 (N_12229,N_11544,N_11617);
xnor U12230 (N_12230,N_11636,N_11894);
nor U12231 (N_12231,N_11920,N_11513);
xnor U12232 (N_12232,N_11570,N_11567);
or U12233 (N_12233,N_11784,N_11632);
nor U12234 (N_12234,N_11630,N_11540);
nor U12235 (N_12235,N_11826,N_11992);
and U12236 (N_12236,N_11698,N_11532);
nor U12237 (N_12237,N_11591,N_11727);
xnor U12238 (N_12238,N_11583,N_11771);
nor U12239 (N_12239,N_11613,N_11983);
nand U12240 (N_12240,N_11800,N_11938);
nand U12241 (N_12241,N_11640,N_11712);
nand U12242 (N_12242,N_11755,N_11676);
and U12243 (N_12243,N_11716,N_11893);
xor U12244 (N_12244,N_11761,N_11594);
nor U12245 (N_12245,N_11734,N_11841);
and U12246 (N_12246,N_11623,N_11851);
or U12247 (N_12247,N_11572,N_11818);
and U12248 (N_12248,N_11973,N_11750);
nor U12249 (N_12249,N_11871,N_11547);
xnor U12250 (N_12250,N_11532,N_11953);
nor U12251 (N_12251,N_11812,N_11888);
xor U12252 (N_12252,N_11873,N_11618);
nand U12253 (N_12253,N_11618,N_11570);
and U12254 (N_12254,N_11734,N_11896);
and U12255 (N_12255,N_11834,N_11854);
nand U12256 (N_12256,N_11674,N_11850);
nand U12257 (N_12257,N_11609,N_11707);
xor U12258 (N_12258,N_11696,N_11771);
nor U12259 (N_12259,N_11507,N_11736);
or U12260 (N_12260,N_11714,N_11841);
or U12261 (N_12261,N_11764,N_11758);
and U12262 (N_12262,N_11989,N_11842);
nand U12263 (N_12263,N_11592,N_11801);
nor U12264 (N_12264,N_11717,N_11879);
nor U12265 (N_12265,N_11733,N_11554);
and U12266 (N_12266,N_11554,N_11950);
and U12267 (N_12267,N_11636,N_11580);
and U12268 (N_12268,N_11899,N_11885);
nand U12269 (N_12269,N_11737,N_11563);
and U12270 (N_12270,N_11550,N_11770);
nor U12271 (N_12271,N_11902,N_11663);
or U12272 (N_12272,N_11674,N_11886);
nand U12273 (N_12273,N_11731,N_11568);
xor U12274 (N_12274,N_11597,N_11838);
xnor U12275 (N_12275,N_11776,N_11735);
or U12276 (N_12276,N_11985,N_11653);
and U12277 (N_12277,N_11841,N_11529);
and U12278 (N_12278,N_11930,N_11797);
xnor U12279 (N_12279,N_11625,N_11872);
and U12280 (N_12280,N_11806,N_11820);
or U12281 (N_12281,N_11790,N_11691);
and U12282 (N_12282,N_11838,N_11945);
nor U12283 (N_12283,N_11733,N_11670);
nor U12284 (N_12284,N_11992,N_11711);
or U12285 (N_12285,N_11964,N_11720);
xnor U12286 (N_12286,N_11894,N_11525);
or U12287 (N_12287,N_11612,N_11778);
or U12288 (N_12288,N_11721,N_11807);
xnor U12289 (N_12289,N_11794,N_11690);
nor U12290 (N_12290,N_11938,N_11522);
or U12291 (N_12291,N_11856,N_11977);
xnor U12292 (N_12292,N_11593,N_11969);
and U12293 (N_12293,N_11977,N_11722);
nand U12294 (N_12294,N_11553,N_11932);
and U12295 (N_12295,N_11962,N_11912);
and U12296 (N_12296,N_11673,N_11925);
nor U12297 (N_12297,N_11617,N_11633);
nor U12298 (N_12298,N_11789,N_11758);
nand U12299 (N_12299,N_11798,N_11736);
nand U12300 (N_12300,N_11852,N_11765);
nand U12301 (N_12301,N_11773,N_11509);
xor U12302 (N_12302,N_11689,N_11870);
xnor U12303 (N_12303,N_11868,N_11570);
xor U12304 (N_12304,N_11714,N_11747);
or U12305 (N_12305,N_11772,N_11762);
nor U12306 (N_12306,N_11961,N_11860);
xnor U12307 (N_12307,N_11520,N_11781);
xor U12308 (N_12308,N_11599,N_11780);
and U12309 (N_12309,N_11757,N_11776);
nand U12310 (N_12310,N_11551,N_11994);
nand U12311 (N_12311,N_11608,N_11835);
and U12312 (N_12312,N_11951,N_11929);
xnor U12313 (N_12313,N_11910,N_11625);
nor U12314 (N_12314,N_11504,N_11523);
nor U12315 (N_12315,N_11567,N_11841);
or U12316 (N_12316,N_11997,N_11666);
nor U12317 (N_12317,N_11854,N_11890);
nand U12318 (N_12318,N_11913,N_11639);
xnor U12319 (N_12319,N_11888,N_11561);
and U12320 (N_12320,N_11914,N_11966);
nor U12321 (N_12321,N_11941,N_11922);
xor U12322 (N_12322,N_11605,N_11757);
and U12323 (N_12323,N_11902,N_11571);
and U12324 (N_12324,N_11821,N_11902);
nor U12325 (N_12325,N_11941,N_11965);
nand U12326 (N_12326,N_11703,N_11576);
and U12327 (N_12327,N_11531,N_11934);
xor U12328 (N_12328,N_11518,N_11878);
or U12329 (N_12329,N_11678,N_11864);
nor U12330 (N_12330,N_11617,N_11913);
nor U12331 (N_12331,N_11835,N_11774);
and U12332 (N_12332,N_11977,N_11701);
xor U12333 (N_12333,N_11739,N_11665);
or U12334 (N_12334,N_11615,N_11717);
or U12335 (N_12335,N_11786,N_11628);
nand U12336 (N_12336,N_11717,N_11748);
xnor U12337 (N_12337,N_11849,N_11581);
nand U12338 (N_12338,N_11621,N_11748);
nand U12339 (N_12339,N_11542,N_11778);
nand U12340 (N_12340,N_11544,N_11857);
nor U12341 (N_12341,N_11591,N_11569);
xnor U12342 (N_12342,N_11504,N_11536);
and U12343 (N_12343,N_11795,N_11859);
nand U12344 (N_12344,N_11839,N_11888);
or U12345 (N_12345,N_11800,N_11915);
and U12346 (N_12346,N_11859,N_11831);
or U12347 (N_12347,N_11700,N_11769);
and U12348 (N_12348,N_11600,N_11574);
or U12349 (N_12349,N_11540,N_11568);
xnor U12350 (N_12350,N_11619,N_11507);
nor U12351 (N_12351,N_11628,N_11803);
nand U12352 (N_12352,N_11817,N_11633);
and U12353 (N_12353,N_11650,N_11873);
nor U12354 (N_12354,N_11521,N_11707);
nor U12355 (N_12355,N_11633,N_11747);
nand U12356 (N_12356,N_11657,N_11917);
nand U12357 (N_12357,N_11738,N_11628);
nor U12358 (N_12358,N_11576,N_11585);
xor U12359 (N_12359,N_11983,N_11651);
xnor U12360 (N_12360,N_11927,N_11762);
nand U12361 (N_12361,N_11957,N_11566);
or U12362 (N_12362,N_11873,N_11765);
nand U12363 (N_12363,N_11517,N_11728);
nand U12364 (N_12364,N_11626,N_11596);
nand U12365 (N_12365,N_11776,N_11726);
and U12366 (N_12366,N_11889,N_11700);
nand U12367 (N_12367,N_11796,N_11979);
or U12368 (N_12368,N_11670,N_11838);
xnor U12369 (N_12369,N_11959,N_11710);
nor U12370 (N_12370,N_11652,N_11786);
xnor U12371 (N_12371,N_11988,N_11797);
and U12372 (N_12372,N_11697,N_11937);
nand U12373 (N_12373,N_11600,N_11837);
or U12374 (N_12374,N_11663,N_11767);
nand U12375 (N_12375,N_11824,N_11584);
or U12376 (N_12376,N_11560,N_11988);
or U12377 (N_12377,N_11600,N_11769);
nand U12378 (N_12378,N_11909,N_11726);
and U12379 (N_12379,N_11738,N_11715);
nor U12380 (N_12380,N_11846,N_11902);
nor U12381 (N_12381,N_11786,N_11513);
nand U12382 (N_12382,N_11776,N_11848);
nor U12383 (N_12383,N_11871,N_11797);
and U12384 (N_12384,N_11644,N_11551);
nand U12385 (N_12385,N_11772,N_11999);
or U12386 (N_12386,N_11793,N_11568);
nand U12387 (N_12387,N_11696,N_11895);
xor U12388 (N_12388,N_11967,N_11759);
xnor U12389 (N_12389,N_11841,N_11740);
xor U12390 (N_12390,N_11595,N_11692);
and U12391 (N_12391,N_11751,N_11776);
xnor U12392 (N_12392,N_11506,N_11819);
nand U12393 (N_12393,N_11594,N_11886);
or U12394 (N_12394,N_11704,N_11632);
xnor U12395 (N_12395,N_11783,N_11825);
or U12396 (N_12396,N_11567,N_11921);
or U12397 (N_12397,N_11581,N_11668);
or U12398 (N_12398,N_11712,N_11600);
or U12399 (N_12399,N_11853,N_11511);
or U12400 (N_12400,N_11712,N_11978);
xor U12401 (N_12401,N_11810,N_11706);
or U12402 (N_12402,N_11569,N_11718);
xnor U12403 (N_12403,N_11554,N_11614);
nand U12404 (N_12404,N_11858,N_11912);
or U12405 (N_12405,N_11749,N_11501);
nand U12406 (N_12406,N_11677,N_11863);
xnor U12407 (N_12407,N_11670,N_11653);
nand U12408 (N_12408,N_11521,N_11784);
and U12409 (N_12409,N_11688,N_11963);
or U12410 (N_12410,N_11796,N_11900);
or U12411 (N_12411,N_11629,N_11518);
xnor U12412 (N_12412,N_11986,N_11639);
nand U12413 (N_12413,N_11559,N_11957);
and U12414 (N_12414,N_11957,N_11613);
and U12415 (N_12415,N_11789,N_11548);
nand U12416 (N_12416,N_11730,N_11606);
or U12417 (N_12417,N_11648,N_11992);
xor U12418 (N_12418,N_11938,N_11802);
and U12419 (N_12419,N_11863,N_11704);
xnor U12420 (N_12420,N_11664,N_11634);
or U12421 (N_12421,N_11828,N_11944);
or U12422 (N_12422,N_11924,N_11634);
or U12423 (N_12423,N_11716,N_11610);
and U12424 (N_12424,N_11714,N_11872);
or U12425 (N_12425,N_11554,N_11573);
xor U12426 (N_12426,N_11976,N_11528);
xnor U12427 (N_12427,N_11670,N_11801);
and U12428 (N_12428,N_11837,N_11744);
or U12429 (N_12429,N_11649,N_11973);
nand U12430 (N_12430,N_11648,N_11604);
or U12431 (N_12431,N_11587,N_11620);
nor U12432 (N_12432,N_11682,N_11863);
nor U12433 (N_12433,N_11817,N_11874);
nor U12434 (N_12434,N_11555,N_11757);
or U12435 (N_12435,N_11662,N_11621);
nand U12436 (N_12436,N_11637,N_11634);
and U12437 (N_12437,N_11769,N_11928);
and U12438 (N_12438,N_11536,N_11653);
xor U12439 (N_12439,N_11682,N_11578);
xnor U12440 (N_12440,N_11710,N_11771);
and U12441 (N_12441,N_11932,N_11828);
xor U12442 (N_12442,N_11956,N_11840);
or U12443 (N_12443,N_11850,N_11971);
xnor U12444 (N_12444,N_11659,N_11672);
xnor U12445 (N_12445,N_11636,N_11587);
nand U12446 (N_12446,N_11582,N_11719);
and U12447 (N_12447,N_11833,N_11598);
and U12448 (N_12448,N_11828,N_11927);
or U12449 (N_12449,N_11743,N_11679);
or U12450 (N_12450,N_11830,N_11743);
and U12451 (N_12451,N_11783,N_11653);
nand U12452 (N_12452,N_11908,N_11535);
nand U12453 (N_12453,N_11516,N_11744);
and U12454 (N_12454,N_11505,N_11949);
and U12455 (N_12455,N_11775,N_11803);
xnor U12456 (N_12456,N_11607,N_11789);
or U12457 (N_12457,N_11698,N_11736);
nor U12458 (N_12458,N_11649,N_11531);
nand U12459 (N_12459,N_11601,N_11951);
nand U12460 (N_12460,N_11813,N_11854);
xnor U12461 (N_12461,N_11772,N_11511);
nor U12462 (N_12462,N_11910,N_11689);
nor U12463 (N_12463,N_11905,N_11803);
nand U12464 (N_12464,N_11583,N_11691);
xnor U12465 (N_12465,N_11553,N_11558);
and U12466 (N_12466,N_11953,N_11810);
xor U12467 (N_12467,N_11621,N_11962);
or U12468 (N_12468,N_11569,N_11884);
and U12469 (N_12469,N_11658,N_11674);
nand U12470 (N_12470,N_11888,N_11827);
xnor U12471 (N_12471,N_11656,N_11602);
xor U12472 (N_12472,N_11644,N_11733);
xnor U12473 (N_12473,N_11788,N_11839);
or U12474 (N_12474,N_11807,N_11580);
nor U12475 (N_12475,N_11804,N_11974);
and U12476 (N_12476,N_11960,N_11905);
nand U12477 (N_12477,N_11933,N_11552);
xor U12478 (N_12478,N_11838,N_11612);
xnor U12479 (N_12479,N_11515,N_11959);
and U12480 (N_12480,N_11733,N_11669);
or U12481 (N_12481,N_11984,N_11872);
xor U12482 (N_12482,N_11983,N_11677);
nor U12483 (N_12483,N_11692,N_11526);
nor U12484 (N_12484,N_11891,N_11851);
nor U12485 (N_12485,N_11663,N_11905);
nand U12486 (N_12486,N_11808,N_11946);
xor U12487 (N_12487,N_11635,N_11673);
and U12488 (N_12488,N_11971,N_11627);
and U12489 (N_12489,N_11528,N_11811);
and U12490 (N_12490,N_11760,N_11855);
and U12491 (N_12491,N_11666,N_11635);
or U12492 (N_12492,N_11926,N_11832);
nand U12493 (N_12493,N_11831,N_11653);
and U12494 (N_12494,N_11639,N_11604);
nand U12495 (N_12495,N_11516,N_11698);
nor U12496 (N_12496,N_11867,N_11649);
or U12497 (N_12497,N_11659,N_11774);
or U12498 (N_12498,N_11875,N_11656);
nand U12499 (N_12499,N_11708,N_11558);
nor U12500 (N_12500,N_12289,N_12121);
and U12501 (N_12501,N_12272,N_12404);
xor U12502 (N_12502,N_12168,N_12380);
nor U12503 (N_12503,N_12324,N_12328);
nor U12504 (N_12504,N_12428,N_12152);
or U12505 (N_12505,N_12149,N_12155);
nor U12506 (N_12506,N_12119,N_12217);
nand U12507 (N_12507,N_12263,N_12062);
nand U12508 (N_12508,N_12116,N_12470);
xnor U12509 (N_12509,N_12225,N_12012);
or U12510 (N_12510,N_12177,N_12020);
nor U12511 (N_12511,N_12036,N_12109);
xor U12512 (N_12512,N_12166,N_12189);
nand U12513 (N_12513,N_12201,N_12486);
or U12514 (N_12514,N_12124,N_12133);
and U12515 (N_12515,N_12390,N_12460);
or U12516 (N_12516,N_12331,N_12004);
xnor U12517 (N_12517,N_12264,N_12452);
xor U12518 (N_12518,N_12314,N_12363);
and U12519 (N_12519,N_12374,N_12006);
nor U12520 (N_12520,N_12430,N_12472);
or U12521 (N_12521,N_12199,N_12031);
and U12522 (N_12522,N_12317,N_12110);
nor U12523 (N_12523,N_12340,N_12093);
nand U12524 (N_12524,N_12053,N_12043);
nor U12525 (N_12525,N_12481,N_12044);
xor U12526 (N_12526,N_12196,N_12490);
xnor U12527 (N_12527,N_12250,N_12388);
or U12528 (N_12528,N_12073,N_12045);
or U12529 (N_12529,N_12334,N_12033);
and U12530 (N_12530,N_12478,N_12300);
nand U12531 (N_12531,N_12425,N_12030);
or U12532 (N_12532,N_12157,N_12418);
xor U12533 (N_12533,N_12247,N_12160);
nor U12534 (N_12534,N_12174,N_12091);
or U12535 (N_12535,N_12444,N_12140);
nand U12536 (N_12536,N_12249,N_12156);
xor U12537 (N_12537,N_12268,N_12187);
nor U12538 (N_12538,N_12009,N_12241);
nor U12539 (N_12539,N_12219,N_12059);
and U12540 (N_12540,N_12105,N_12055);
and U12541 (N_12541,N_12106,N_12354);
nand U12542 (N_12542,N_12150,N_12101);
or U12543 (N_12543,N_12415,N_12279);
nand U12544 (N_12544,N_12227,N_12092);
nor U12545 (N_12545,N_12173,N_12099);
nor U12546 (N_12546,N_12089,N_12135);
nor U12547 (N_12547,N_12002,N_12299);
xnor U12548 (N_12548,N_12032,N_12207);
nand U12549 (N_12549,N_12370,N_12497);
xnor U12550 (N_12550,N_12190,N_12286);
nand U12551 (N_12551,N_12401,N_12067);
and U12552 (N_12552,N_12240,N_12474);
or U12553 (N_12553,N_12145,N_12079);
nor U12554 (N_12554,N_12069,N_12327);
and U12555 (N_12555,N_12206,N_12255);
and U12556 (N_12556,N_12267,N_12407);
or U12557 (N_12557,N_12080,N_12096);
or U12558 (N_12558,N_12371,N_12115);
and U12559 (N_12559,N_12086,N_12386);
xnor U12560 (N_12560,N_12066,N_12085);
nor U12561 (N_12561,N_12170,N_12186);
or U12562 (N_12562,N_12381,N_12113);
or U12563 (N_12563,N_12226,N_12471);
xor U12564 (N_12564,N_12253,N_12224);
nand U12565 (N_12565,N_12362,N_12432);
or U12566 (N_12566,N_12266,N_12214);
xor U12567 (N_12567,N_12010,N_12018);
nor U12568 (N_12568,N_12039,N_12368);
xor U12569 (N_12569,N_12395,N_12344);
nand U12570 (N_12570,N_12313,N_12408);
nor U12571 (N_12571,N_12038,N_12146);
xnor U12572 (N_12572,N_12489,N_12469);
nand U12573 (N_12573,N_12366,N_12373);
nor U12574 (N_12574,N_12341,N_12178);
nor U12575 (N_12575,N_12333,N_12284);
and U12576 (N_12576,N_12283,N_12348);
and U12577 (N_12577,N_12143,N_12398);
or U12578 (N_12578,N_12394,N_12194);
and U12579 (N_12579,N_12367,N_12385);
nor U12580 (N_12580,N_12412,N_12054);
nand U12581 (N_12581,N_12052,N_12378);
nand U12582 (N_12582,N_12482,N_12296);
and U12583 (N_12583,N_12280,N_12181);
or U12584 (N_12584,N_12431,N_12137);
nor U12585 (N_12585,N_12082,N_12212);
or U12586 (N_12586,N_12446,N_12271);
xor U12587 (N_12587,N_12223,N_12165);
nand U12588 (N_12588,N_12361,N_12159);
nand U12589 (N_12589,N_12111,N_12123);
or U12590 (N_12590,N_12320,N_12245);
or U12591 (N_12591,N_12007,N_12161);
or U12592 (N_12592,N_12433,N_12304);
nor U12593 (N_12593,N_12202,N_12203);
and U12594 (N_12594,N_12282,N_12466);
nor U12595 (N_12595,N_12318,N_12162);
and U12596 (N_12596,N_12246,N_12274);
nand U12597 (N_12597,N_12376,N_12236);
nand U12598 (N_12598,N_12238,N_12352);
xor U12599 (N_12599,N_12211,N_12322);
and U12600 (N_12600,N_12434,N_12134);
xnor U12601 (N_12601,N_12290,N_12473);
or U12602 (N_12602,N_12426,N_12131);
xor U12603 (N_12603,N_12005,N_12229);
or U12604 (N_12604,N_12015,N_12248);
and U12605 (N_12605,N_12406,N_12335);
xnor U12606 (N_12606,N_12112,N_12493);
xor U12607 (N_12607,N_12025,N_12468);
or U12608 (N_12608,N_12127,N_12485);
and U12609 (N_12609,N_12356,N_12323);
or U12610 (N_12610,N_12421,N_12338);
and U12611 (N_12611,N_12251,N_12442);
nand U12612 (N_12612,N_12281,N_12041);
and U12613 (N_12613,N_12026,N_12278);
nor U12614 (N_12614,N_12494,N_12014);
nand U12615 (N_12615,N_12477,N_12070);
xor U12616 (N_12616,N_12488,N_12037);
and U12617 (N_12617,N_12402,N_12372);
nor U12618 (N_12618,N_12332,N_12013);
and U12619 (N_12619,N_12273,N_12128);
nand U12620 (N_12620,N_12265,N_12213);
and U12621 (N_12621,N_12000,N_12429);
and U12622 (N_12622,N_12384,N_12355);
or U12623 (N_12623,N_12192,N_12021);
or U12624 (N_12624,N_12019,N_12308);
and U12625 (N_12625,N_12369,N_12056);
nor U12626 (N_12626,N_12098,N_12419);
nor U12627 (N_12627,N_12463,N_12063);
nor U12628 (N_12628,N_12158,N_12144);
and U12629 (N_12629,N_12126,N_12254);
nand U12630 (N_12630,N_12405,N_12450);
nand U12631 (N_12631,N_12197,N_12205);
nand U12632 (N_12632,N_12297,N_12357);
xnor U12633 (N_12633,N_12310,N_12084);
and U12634 (N_12634,N_12058,N_12151);
and U12635 (N_12635,N_12411,N_12258);
and U12636 (N_12636,N_12330,N_12464);
xor U12637 (N_12637,N_12076,N_12336);
or U12638 (N_12638,N_12233,N_12060);
xor U12639 (N_12639,N_12094,N_12017);
and U12640 (N_12640,N_12035,N_12292);
xor U12641 (N_12641,N_12321,N_12285);
or U12642 (N_12642,N_12343,N_12438);
nand U12643 (N_12643,N_12024,N_12257);
or U12644 (N_12644,N_12183,N_12100);
nand U12645 (N_12645,N_12209,N_12391);
nor U12646 (N_12646,N_12184,N_12191);
nor U12647 (N_12647,N_12360,N_12277);
nor U12648 (N_12648,N_12455,N_12298);
nor U12649 (N_12649,N_12185,N_12312);
or U12650 (N_12650,N_12410,N_12057);
nand U12651 (N_12651,N_12164,N_12011);
and U12652 (N_12652,N_12072,N_12034);
or U12653 (N_12653,N_12325,N_12364);
and U12654 (N_12654,N_12230,N_12351);
or U12655 (N_12655,N_12074,N_12347);
and U12656 (N_12656,N_12228,N_12068);
xor U12657 (N_12657,N_12262,N_12326);
xor U12658 (N_12658,N_12200,N_12046);
or U12659 (N_12659,N_12008,N_12182);
nor U12660 (N_12660,N_12171,N_12252);
nor U12661 (N_12661,N_12449,N_12193);
or U12662 (N_12662,N_12475,N_12132);
xor U12663 (N_12663,N_12359,N_12003);
or U12664 (N_12664,N_12403,N_12393);
nor U12665 (N_12665,N_12294,N_12422);
nor U12666 (N_12666,N_12275,N_12427);
and U12667 (N_12667,N_12016,N_12048);
nor U12668 (N_12668,N_12118,N_12172);
and U12669 (N_12669,N_12476,N_12028);
and U12670 (N_12670,N_12456,N_12130);
xor U12671 (N_12671,N_12496,N_12022);
or U12672 (N_12672,N_12437,N_12188);
or U12673 (N_12673,N_12392,N_12107);
or U12674 (N_12674,N_12491,N_12396);
nand U12675 (N_12675,N_12305,N_12220);
and U12676 (N_12676,N_12256,N_12029);
nand U12677 (N_12677,N_12163,N_12088);
and U12678 (N_12678,N_12498,N_12218);
and U12679 (N_12679,N_12315,N_12081);
or U12680 (N_12680,N_12458,N_12234);
nand U12681 (N_12681,N_12465,N_12027);
and U12682 (N_12682,N_12120,N_12291);
xor U12683 (N_12683,N_12139,N_12288);
xnor U12684 (N_12684,N_12342,N_12413);
nand U12685 (N_12685,N_12479,N_12269);
xor U12686 (N_12686,N_12484,N_12409);
or U12687 (N_12687,N_12397,N_12353);
nand U12688 (N_12688,N_12339,N_12365);
and U12689 (N_12689,N_12459,N_12179);
xor U12690 (N_12690,N_12232,N_12221);
nor U12691 (N_12691,N_12210,N_12461);
and U12692 (N_12692,N_12329,N_12492);
xnor U12693 (N_12693,N_12042,N_12122);
nor U12694 (N_12694,N_12083,N_12167);
nand U12695 (N_12695,N_12138,N_12379);
or U12696 (N_12696,N_12375,N_12261);
nand U12697 (N_12697,N_12345,N_12441);
nand U12698 (N_12698,N_12195,N_12423);
and U12699 (N_12699,N_12102,N_12142);
nand U12700 (N_12700,N_12420,N_12141);
nand U12701 (N_12701,N_12198,N_12148);
and U12702 (N_12702,N_12001,N_12061);
and U12703 (N_12703,N_12176,N_12451);
and U12704 (N_12704,N_12071,N_12350);
xnor U12705 (N_12705,N_12244,N_12243);
xnor U12706 (N_12706,N_12399,N_12064);
and U12707 (N_12707,N_12337,N_12097);
nor U12708 (N_12708,N_12239,N_12154);
xnor U12709 (N_12709,N_12259,N_12270);
and U12710 (N_12710,N_12114,N_12180);
and U12711 (N_12711,N_12153,N_12454);
nor U12712 (N_12712,N_12075,N_12316);
or U12713 (N_12713,N_12440,N_12104);
nand U12714 (N_12714,N_12295,N_12443);
nand U12715 (N_12715,N_12204,N_12215);
xor U12716 (N_12716,N_12023,N_12208);
or U12717 (N_12717,N_12237,N_12095);
nand U12718 (N_12718,N_12319,N_12483);
nand U12719 (N_12719,N_12103,N_12051);
and U12720 (N_12720,N_12242,N_12435);
nor U12721 (N_12721,N_12276,N_12065);
or U12722 (N_12722,N_12480,N_12387);
xor U12723 (N_12723,N_12175,N_12448);
xnor U12724 (N_12724,N_12377,N_12108);
or U12725 (N_12725,N_12417,N_12077);
nor U12726 (N_12726,N_12389,N_12495);
xnor U12727 (N_12727,N_12047,N_12222);
nor U12728 (N_12728,N_12307,N_12302);
or U12729 (N_12729,N_12382,N_12260);
xor U12730 (N_12730,N_12049,N_12293);
xor U12731 (N_12731,N_12303,N_12040);
nand U12732 (N_12732,N_12346,N_12436);
or U12733 (N_12733,N_12358,N_12447);
and U12734 (N_12734,N_12439,N_12078);
nand U12735 (N_12735,N_12311,N_12416);
or U12736 (N_12736,N_12383,N_12467);
nor U12737 (N_12737,N_12050,N_12125);
xor U12738 (N_12738,N_12400,N_12231);
nand U12739 (N_12739,N_12301,N_12306);
and U12740 (N_12740,N_12216,N_12445);
nor U12741 (N_12741,N_12462,N_12453);
nand U12742 (N_12742,N_12349,N_12090);
nor U12743 (N_12743,N_12487,N_12129);
nor U12744 (N_12744,N_12169,N_12235);
nand U12745 (N_12745,N_12499,N_12414);
nor U12746 (N_12746,N_12424,N_12087);
or U12747 (N_12747,N_12136,N_12309);
xor U12748 (N_12748,N_12457,N_12287);
and U12749 (N_12749,N_12117,N_12147);
nor U12750 (N_12750,N_12338,N_12314);
nor U12751 (N_12751,N_12297,N_12473);
nand U12752 (N_12752,N_12018,N_12491);
and U12753 (N_12753,N_12385,N_12479);
nor U12754 (N_12754,N_12034,N_12164);
and U12755 (N_12755,N_12012,N_12295);
or U12756 (N_12756,N_12338,N_12304);
xnor U12757 (N_12757,N_12275,N_12301);
nand U12758 (N_12758,N_12391,N_12177);
and U12759 (N_12759,N_12314,N_12079);
nor U12760 (N_12760,N_12442,N_12074);
nand U12761 (N_12761,N_12161,N_12303);
xor U12762 (N_12762,N_12032,N_12202);
nor U12763 (N_12763,N_12162,N_12428);
nor U12764 (N_12764,N_12098,N_12244);
nand U12765 (N_12765,N_12195,N_12299);
nand U12766 (N_12766,N_12111,N_12051);
nand U12767 (N_12767,N_12411,N_12471);
xor U12768 (N_12768,N_12057,N_12325);
and U12769 (N_12769,N_12260,N_12071);
nor U12770 (N_12770,N_12388,N_12155);
and U12771 (N_12771,N_12221,N_12041);
nor U12772 (N_12772,N_12075,N_12359);
xnor U12773 (N_12773,N_12336,N_12081);
nand U12774 (N_12774,N_12200,N_12223);
nor U12775 (N_12775,N_12498,N_12008);
nor U12776 (N_12776,N_12170,N_12000);
nand U12777 (N_12777,N_12012,N_12335);
xor U12778 (N_12778,N_12390,N_12020);
and U12779 (N_12779,N_12185,N_12104);
nand U12780 (N_12780,N_12481,N_12229);
xnor U12781 (N_12781,N_12021,N_12465);
and U12782 (N_12782,N_12378,N_12291);
xor U12783 (N_12783,N_12111,N_12133);
or U12784 (N_12784,N_12349,N_12189);
or U12785 (N_12785,N_12029,N_12041);
xor U12786 (N_12786,N_12072,N_12236);
or U12787 (N_12787,N_12182,N_12051);
and U12788 (N_12788,N_12164,N_12202);
nor U12789 (N_12789,N_12061,N_12129);
nor U12790 (N_12790,N_12189,N_12011);
nand U12791 (N_12791,N_12397,N_12096);
or U12792 (N_12792,N_12484,N_12420);
or U12793 (N_12793,N_12099,N_12077);
nor U12794 (N_12794,N_12348,N_12454);
or U12795 (N_12795,N_12258,N_12453);
xor U12796 (N_12796,N_12155,N_12180);
and U12797 (N_12797,N_12475,N_12151);
or U12798 (N_12798,N_12093,N_12151);
or U12799 (N_12799,N_12385,N_12040);
and U12800 (N_12800,N_12323,N_12074);
or U12801 (N_12801,N_12376,N_12012);
or U12802 (N_12802,N_12071,N_12196);
nand U12803 (N_12803,N_12312,N_12376);
nor U12804 (N_12804,N_12186,N_12086);
or U12805 (N_12805,N_12214,N_12092);
or U12806 (N_12806,N_12021,N_12230);
xnor U12807 (N_12807,N_12211,N_12139);
nor U12808 (N_12808,N_12208,N_12263);
nand U12809 (N_12809,N_12233,N_12426);
xor U12810 (N_12810,N_12186,N_12286);
nand U12811 (N_12811,N_12319,N_12055);
or U12812 (N_12812,N_12283,N_12035);
or U12813 (N_12813,N_12280,N_12211);
xor U12814 (N_12814,N_12259,N_12177);
nand U12815 (N_12815,N_12481,N_12465);
and U12816 (N_12816,N_12253,N_12369);
xor U12817 (N_12817,N_12402,N_12135);
and U12818 (N_12818,N_12057,N_12216);
and U12819 (N_12819,N_12199,N_12198);
and U12820 (N_12820,N_12373,N_12156);
xnor U12821 (N_12821,N_12390,N_12129);
nor U12822 (N_12822,N_12139,N_12309);
xnor U12823 (N_12823,N_12349,N_12214);
nor U12824 (N_12824,N_12096,N_12230);
nor U12825 (N_12825,N_12069,N_12415);
nand U12826 (N_12826,N_12244,N_12012);
nand U12827 (N_12827,N_12344,N_12196);
or U12828 (N_12828,N_12464,N_12393);
or U12829 (N_12829,N_12223,N_12190);
nand U12830 (N_12830,N_12400,N_12333);
nor U12831 (N_12831,N_12342,N_12307);
nand U12832 (N_12832,N_12419,N_12210);
xnor U12833 (N_12833,N_12344,N_12128);
nand U12834 (N_12834,N_12076,N_12429);
nor U12835 (N_12835,N_12084,N_12240);
and U12836 (N_12836,N_12381,N_12474);
and U12837 (N_12837,N_12284,N_12477);
or U12838 (N_12838,N_12276,N_12239);
nor U12839 (N_12839,N_12029,N_12328);
nand U12840 (N_12840,N_12200,N_12337);
and U12841 (N_12841,N_12394,N_12259);
nor U12842 (N_12842,N_12386,N_12125);
and U12843 (N_12843,N_12058,N_12006);
and U12844 (N_12844,N_12007,N_12159);
or U12845 (N_12845,N_12063,N_12432);
and U12846 (N_12846,N_12434,N_12374);
nand U12847 (N_12847,N_12229,N_12475);
xnor U12848 (N_12848,N_12478,N_12001);
nor U12849 (N_12849,N_12025,N_12137);
xor U12850 (N_12850,N_12410,N_12286);
xor U12851 (N_12851,N_12300,N_12260);
and U12852 (N_12852,N_12162,N_12346);
nor U12853 (N_12853,N_12306,N_12251);
xnor U12854 (N_12854,N_12346,N_12352);
and U12855 (N_12855,N_12012,N_12489);
xnor U12856 (N_12856,N_12338,N_12311);
or U12857 (N_12857,N_12399,N_12140);
or U12858 (N_12858,N_12363,N_12222);
xnor U12859 (N_12859,N_12431,N_12104);
and U12860 (N_12860,N_12361,N_12450);
nor U12861 (N_12861,N_12382,N_12321);
nand U12862 (N_12862,N_12111,N_12347);
or U12863 (N_12863,N_12258,N_12037);
nand U12864 (N_12864,N_12003,N_12378);
or U12865 (N_12865,N_12051,N_12470);
nor U12866 (N_12866,N_12434,N_12175);
or U12867 (N_12867,N_12133,N_12076);
and U12868 (N_12868,N_12407,N_12436);
xor U12869 (N_12869,N_12304,N_12101);
nor U12870 (N_12870,N_12376,N_12087);
nand U12871 (N_12871,N_12194,N_12456);
and U12872 (N_12872,N_12198,N_12026);
xnor U12873 (N_12873,N_12009,N_12492);
xnor U12874 (N_12874,N_12157,N_12233);
nand U12875 (N_12875,N_12443,N_12071);
or U12876 (N_12876,N_12196,N_12357);
nor U12877 (N_12877,N_12052,N_12332);
nand U12878 (N_12878,N_12315,N_12328);
xor U12879 (N_12879,N_12037,N_12456);
or U12880 (N_12880,N_12117,N_12376);
nor U12881 (N_12881,N_12449,N_12216);
nand U12882 (N_12882,N_12476,N_12440);
nor U12883 (N_12883,N_12027,N_12436);
or U12884 (N_12884,N_12133,N_12132);
and U12885 (N_12885,N_12130,N_12326);
nand U12886 (N_12886,N_12037,N_12362);
or U12887 (N_12887,N_12100,N_12068);
or U12888 (N_12888,N_12252,N_12397);
nand U12889 (N_12889,N_12085,N_12240);
nor U12890 (N_12890,N_12393,N_12257);
nor U12891 (N_12891,N_12437,N_12347);
and U12892 (N_12892,N_12429,N_12182);
xnor U12893 (N_12893,N_12093,N_12387);
xnor U12894 (N_12894,N_12111,N_12323);
or U12895 (N_12895,N_12176,N_12441);
or U12896 (N_12896,N_12023,N_12050);
and U12897 (N_12897,N_12147,N_12484);
nor U12898 (N_12898,N_12056,N_12405);
nand U12899 (N_12899,N_12270,N_12499);
nand U12900 (N_12900,N_12335,N_12172);
or U12901 (N_12901,N_12464,N_12243);
xnor U12902 (N_12902,N_12192,N_12370);
nor U12903 (N_12903,N_12186,N_12022);
or U12904 (N_12904,N_12032,N_12361);
and U12905 (N_12905,N_12049,N_12223);
or U12906 (N_12906,N_12307,N_12104);
xor U12907 (N_12907,N_12180,N_12156);
nand U12908 (N_12908,N_12259,N_12024);
nand U12909 (N_12909,N_12404,N_12396);
and U12910 (N_12910,N_12116,N_12326);
or U12911 (N_12911,N_12441,N_12282);
nor U12912 (N_12912,N_12145,N_12264);
and U12913 (N_12913,N_12062,N_12246);
and U12914 (N_12914,N_12142,N_12366);
nor U12915 (N_12915,N_12283,N_12225);
and U12916 (N_12916,N_12144,N_12310);
nor U12917 (N_12917,N_12265,N_12217);
or U12918 (N_12918,N_12124,N_12070);
nand U12919 (N_12919,N_12017,N_12162);
xor U12920 (N_12920,N_12102,N_12400);
nor U12921 (N_12921,N_12268,N_12068);
and U12922 (N_12922,N_12275,N_12273);
xnor U12923 (N_12923,N_12270,N_12441);
or U12924 (N_12924,N_12461,N_12204);
nor U12925 (N_12925,N_12159,N_12262);
nor U12926 (N_12926,N_12262,N_12340);
nor U12927 (N_12927,N_12291,N_12099);
nor U12928 (N_12928,N_12353,N_12404);
xor U12929 (N_12929,N_12049,N_12130);
or U12930 (N_12930,N_12460,N_12494);
and U12931 (N_12931,N_12302,N_12413);
or U12932 (N_12932,N_12049,N_12194);
nor U12933 (N_12933,N_12107,N_12141);
xor U12934 (N_12934,N_12244,N_12422);
and U12935 (N_12935,N_12440,N_12404);
nand U12936 (N_12936,N_12007,N_12325);
nand U12937 (N_12937,N_12184,N_12303);
and U12938 (N_12938,N_12106,N_12130);
or U12939 (N_12939,N_12201,N_12083);
nor U12940 (N_12940,N_12292,N_12366);
and U12941 (N_12941,N_12358,N_12449);
or U12942 (N_12942,N_12088,N_12269);
or U12943 (N_12943,N_12199,N_12115);
xnor U12944 (N_12944,N_12091,N_12324);
nand U12945 (N_12945,N_12043,N_12476);
and U12946 (N_12946,N_12016,N_12487);
xnor U12947 (N_12947,N_12337,N_12390);
or U12948 (N_12948,N_12072,N_12166);
nor U12949 (N_12949,N_12158,N_12086);
or U12950 (N_12950,N_12493,N_12199);
or U12951 (N_12951,N_12222,N_12048);
or U12952 (N_12952,N_12069,N_12323);
or U12953 (N_12953,N_12230,N_12497);
xor U12954 (N_12954,N_12352,N_12078);
and U12955 (N_12955,N_12476,N_12159);
nand U12956 (N_12956,N_12448,N_12055);
nor U12957 (N_12957,N_12210,N_12488);
or U12958 (N_12958,N_12491,N_12300);
nand U12959 (N_12959,N_12400,N_12111);
nor U12960 (N_12960,N_12416,N_12362);
nor U12961 (N_12961,N_12451,N_12309);
nor U12962 (N_12962,N_12495,N_12482);
xor U12963 (N_12963,N_12349,N_12081);
nand U12964 (N_12964,N_12113,N_12297);
or U12965 (N_12965,N_12282,N_12114);
nand U12966 (N_12966,N_12066,N_12062);
xnor U12967 (N_12967,N_12075,N_12390);
nor U12968 (N_12968,N_12147,N_12107);
or U12969 (N_12969,N_12193,N_12385);
or U12970 (N_12970,N_12169,N_12211);
and U12971 (N_12971,N_12086,N_12031);
or U12972 (N_12972,N_12258,N_12261);
and U12973 (N_12973,N_12227,N_12235);
and U12974 (N_12974,N_12359,N_12153);
and U12975 (N_12975,N_12084,N_12472);
nand U12976 (N_12976,N_12348,N_12180);
and U12977 (N_12977,N_12370,N_12015);
nand U12978 (N_12978,N_12060,N_12153);
or U12979 (N_12979,N_12359,N_12243);
nand U12980 (N_12980,N_12210,N_12167);
nand U12981 (N_12981,N_12008,N_12294);
nor U12982 (N_12982,N_12469,N_12492);
nor U12983 (N_12983,N_12167,N_12465);
and U12984 (N_12984,N_12317,N_12383);
or U12985 (N_12985,N_12402,N_12176);
or U12986 (N_12986,N_12254,N_12379);
xnor U12987 (N_12987,N_12191,N_12203);
nand U12988 (N_12988,N_12045,N_12493);
nand U12989 (N_12989,N_12304,N_12313);
or U12990 (N_12990,N_12457,N_12069);
nor U12991 (N_12991,N_12058,N_12222);
xor U12992 (N_12992,N_12482,N_12316);
nor U12993 (N_12993,N_12499,N_12274);
and U12994 (N_12994,N_12112,N_12231);
or U12995 (N_12995,N_12156,N_12256);
nor U12996 (N_12996,N_12155,N_12160);
nor U12997 (N_12997,N_12079,N_12017);
and U12998 (N_12998,N_12384,N_12377);
and U12999 (N_12999,N_12373,N_12086);
nor U13000 (N_13000,N_12712,N_12944);
nand U13001 (N_13001,N_12638,N_12636);
or U13002 (N_13002,N_12879,N_12943);
xnor U13003 (N_13003,N_12974,N_12545);
xnor U13004 (N_13004,N_12582,N_12503);
and U13005 (N_13005,N_12730,N_12886);
and U13006 (N_13006,N_12977,N_12693);
or U13007 (N_13007,N_12597,N_12561);
xnor U13008 (N_13008,N_12722,N_12979);
xnor U13009 (N_13009,N_12992,N_12566);
nor U13010 (N_13010,N_12514,N_12889);
nor U13011 (N_13011,N_12787,N_12764);
and U13012 (N_13012,N_12505,N_12683);
or U13013 (N_13013,N_12904,N_12710);
nor U13014 (N_13014,N_12718,N_12800);
nor U13015 (N_13015,N_12991,N_12867);
nor U13016 (N_13016,N_12610,N_12825);
nand U13017 (N_13017,N_12589,N_12808);
and U13018 (N_13018,N_12608,N_12644);
nand U13019 (N_13019,N_12637,N_12791);
xor U13020 (N_13020,N_12845,N_12624);
nor U13021 (N_13021,N_12674,N_12887);
nand U13022 (N_13022,N_12769,N_12536);
and U13023 (N_13023,N_12571,N_12661);
nor U13024 (N_13024,N_12990,N_12573);
nand U13025 (N_13025,N_12701,N_12531);
nand U13026 (N_13026,N_12690,N_12524);
nor U13027 (N_13027,N_12975,N_12609);
and U13028 (N_13028,N_12828,N_12994);
or U13029 (N_13029,N_12580,N_12546);
xor U13030 (N_13030,N_12960,N_12817);
nor U13031 (N_13031,N_12537,N_12512);
and U13032 (N_13032,N_12568,N_12553);
nand U13033 (N_13033,N_12947,N_12850);
and U13034 (N_13034,N_12923,N_12551);
and U13035 (N_13035,N_12670,N_12918);
and U13036 (N_13036,N_12803,N_12849);
and U13037 (N_13037,N_12875,N_12767);
and U13038 (N_13038,N_12894,N_12749);
or U13039 (N_13039,N_12687,N_12883);
or U13040 (N_13040,N_12898,N_12731);
and U13041 (N_13041,N_12509,N_12824);
and U13042 (N_13042,N_12869,N_12516);
nand U13043 (N_13043,N_12549,N_12550);
and U13044 (N_13044,N_12532,N_12841);
nor U13045 (N_13045,N_12583,N_12627);
or U13046 (N_13046,N_12941,N_12590);
nor U13047 (N_13047,N_12675,N_12654);
or U13048 (N_13048,N_12956,N_12556);
nand U13049 (N_13049,N_12739,N_12607);
or U13050 (N_13050,N_12686,N_12868);
or U13051 (N_13051,N_12506,N_12938);
nor U13052 (N_13052,N_12615,N_12954);
or U13053 (N_13053,N_12720,N_12511);
nand U13054 (N_13054,N_12851,N_12581);
xnor U13055 (N_13055,N_12909,N_12903);
nand U13056 (N_13056,N_12703,N_12577);
nand U13057 (N_13057,N_12570,N_12936);
xnor U13058 (N_13058,N_12927,N_12656);
xnor U13059 (N_13059,N_12659,N_12987);
nor U13060 (N_13060,N_12929,N_12510);
and U13061 (N_13061,N_12935,N_12650);
or U13062 (N_13062,N_12804,N_12707);
or U13063 (N_13063,N_12873,N_12774);
or U13064 (N_13064,N_12959,N_12897);
nor U13065 (N_13065,N_12965,N_12876);
and U13066 (N_13066,N_12572,N_12921);
nor U13067 (N_13067,N_12630,N_12756);
or U13068 (N_13068,N_12950,N_12857);
xnor U13069 (N_13069,N_12777,N_12885);
or U13070 (N_13070,N_12812,N_12657);
xnor U13071 (N_13071,N_12585,N_12734);
or U13072 (N_13072,N_12525,N_12881);
nand U13073 (N_13073,N_12575,N_12815);
nor U13074 (N_13074,N_12667,N_12742);
or U13075 (N_13075,N_12946,N_12908);
nand U13076 (N_13076,N_12539,N_12919);
and U13077 (N_13077,N_12666,N_12829);
xor U13078 (N_13078,N_12942,N_12890);
and U13079 (N_13079,N_12858,N_12939);
or U13080 (N_13080,N_12621,N_12902);
xnor U13081 (N_13081,N_12591,N_12809);
xnor U13082 (N_13082,N_12719,N_12515);
and U13083 (N_13083,N_12662,N_12555);
or U13084 (N_13084,N_12784,N_12911);
nand U13085 (N_13085,N_12934,N_12755);
or U13086 (N_13086,N_12775,N_12642);
xor U13087 (N_13087,N_12925,N_12601);
and U13088 (N_13088,N_12617,N_12518);
or U13089 (N_13089,N_12865,N_12998);
xnor U13090 (N_13090,N_12633,N_12860);
and U13091 (N_13091,N_12928,N_12891);
xnor U13092 (N_13092,N_12626,N_12993);
and U13093 (N_13093,N_12697,N_12584);
and U13094 (N_13094,N_12826,N_12847);
xor U13095 (N_13095,N_12649,N_12966);
and U13096 (N_13096,N_12698,N_12671);
and U13097 (N_13097,N_12527,N_12848);
or U13098 (N_13098,N_12616,N_12785);
nand U13099 (N_13099,N_12738,N_12795);
or U13100 (N_13100,N_12762,N_12844);
and U13101 (N_13101,N_12753,N_12560);
xnor U13102 (N_13102,N_12727,N_12793);
and U13103 (N_13103,N_12827,N_12818);
or U13104 (N_13104,N_12884,N_12677);
nand U13105 (N_13105,N_12595,N_12632);
or U13106 (N_13106,N_12563,N_12872);
or U13107 (N_13107,N_12856,N_12871);
or U13108 (N_13108,N_12507,N_12948);
and U13109 (N_13109,N_12893,N_12535);
nor U13110 (N_13110,N_12972,N_12705);
nand U13111 (N_13111,N_12768,N_12963);
or U13112 (N_13112,N_12988,N_12864);
nor U13113 (N_13113,N_12614,N_12723);
xor U13114 (N_13114,N_12750,N_12688);
nand U13115 (N_13115,N_12878,N_12706);
nand U13116 (N_13116,N_12711,N_12602);
xor U13117 (N_13117,N_12805,N_12761);
or U13118 (N_13118,N_12854,N_12540);
and U13119 (N_13119,N_12840,N_12576);
and U13120 (N_13120,N_12997,N_12645);
nand U13121 (N_13121,N_12830,N_12772);
nor U13122 (N_13122,N_12999,N_12853);
or U13123 (N_13123,N_12866,N_12754);
nor U13124 (N_13124,N_12716,N_12986);
nor U13125 (N_13125,N_12905,N_12631);
xor U13126 (N_13126,N_12736,N_12980);
nand U13127 (N_13127,N_12914,N_12778);
xor U13128 (N_13128,N_12658,N_12564);
or U13129 (N_13129,N_12647,N_12534);
nor U13130 (N_13130,N_12862,N_12985);
or U13131 (N_13131,N_12953,N_12640);
and U13132 (N_13132,N_12766,N_12567);
nor U13133 (N_13133,N_12557,N_12724);
or U13134 (N_13134,N_12870,N_12548);
or U13135 (N_13135,N_12593,N_12973);
nand U13136 (N_13136,N_12838,N_12508);
xnor U13137 (N_13137,N_12554,N_12725);
or U13138 (N_13138,N_12628,N_12874);
and U13139 (N_13139,N_12500,N_12678);
and U13140 (N_13140,N_12821,N_12797);
or U13141 (N_13141,N_12533,N_12618);
or U13142 (N_13142,N_12603,N_12781);
or U13143 (N_13143,N_12790,N_12714);
or U13144 (N_13144,N_12726,N_12932);
xor U13145 (N_13145,N_12746,N_12763);
nor U13146 (N_13146,N_12629,N_12819);
or U13147 (N_13147,N_12964,N_12702);
or U13148 (N_13148,N_12634,N_12517);
nor U13149 (N_13149,N_12691,N_12788);
or U13150 (N_13150,N_12970,N_12920);
nand U13151 (N_13151,N_12733,N_12900);
nand U13152 (N_13152,N_12859,N_12692);
xor U13153 (N_13153,N_12839,N_12660);
nand U13154 (N_13154,N_12699,N_12896);
nand U13155 (N_13155,N_12729,N_12861);
nor U13156 (N_13156,N_12810,N_12913);
xnor U13157 (N_13157,N_12802,N_12522);
xor U13158 (N_13158,N_12747,N_12926);
xnor U13159 (N_13159,N_12813,N_12892);
or U13160 (N_13160,N_12646,N_12569);
nor U13161 (N_13161,N_12620,N_12744);
xor U13162 (N_13162,N_12945,N_12759);
nor U13163 (N_13163,N_12700,N_12728);
and U13164 (N_13164,N_12796,N_12820);
and U13165 (N_13165,N_12673,N_12842);
and U13166 (N_13166,N_12606,N_12922);
nor U13167 (N_13167,N_12619,N_12961);
nor U13168 (N_13168,N_12600,N_12594);
xnor U13169 (N_13169,N_12917,N_12780);
nor U13170 (N_13170,N_12641,N_12831);
and U13171 (N_13171,N_12635,N_12578);
nand U13172 (N_13172,N_12757,N_12924);
xor U13173 (N_13173,N_12915,N_12740);
xor U13174 (N_13174,N_12715,N_12748);
or U13175 (N_13175,N_12835,N_12741);
nand U13176 (N_13176,N_12598,N_12852);
xnor U13177 (N_13177,N_12613,N_12669);
xnor U13178 (N_13178,N_12709,N_12989);
or U13179 (N_13179,N_12528,N_12940);
nand U13180 (N_13180,N_12513,N_12834);
xnor U13181 (N_13181,N_12968,N_12822);
and U13182 (N_13182,N_12639,N_12758);
or U13183 (N_13183,N_12502,N_12910);
nand U13184 (N_13184,N_12541,N_12694);
nor U13185 (N_13185,N_12983,N_12996);
nand U13186 (N_13186,N_12931,N_12651);
xnor U13187 (N_13187,N_12765,N_12832);
or U13188 (N_13188,N_12933,N_12969);
xor U13189 (N_13189,N_12837,N_12745);
and U13190 (N_13190,N_12579,N_12882);
xnor U13191 (N_13191,N_12681,N_12958);
or U13192 (N_13192,N_12562,N_12779);
nand U13193 (N_13193,N_12558,N_12520);
and U13194 (N_13194,N_12836,N_12596);
or U13195 (N_13195,N_12529,N_12542);
nand U13196 (N_13196,N_12521,N_12798);
xor U13197 (N_13197,N_12648,N_12721);
and U13198 (N_13198,N_12906,N_12957);
nand U13199 (N_13199,N_12743,N_12971);
nand U13200 (N_13200,N_12623,N_12770);
nand U13201 (N_13201,N_12912,N_12689);
or U13202 (N_13202,N_12814,N_12622);
xor U13203 (N_13203,N_12574,N_12982);
nand U13204 (N_13204,N_12776,N_12559);
xor U13205 (N_13205,N_12823,N_12794);
nand U13206 (N_13206,N_12751,N_12530);
nand U13207 (N_13207,N_12732,N_12984);
xor U13208 (N_13208,N_12955,N_12592);
nor U13209 (N_13209,N_12586,N_12708);
nand U13210 (N_13210,N_12672,N_12665);
nand U13211 (N_13211,N_12833,N_12519);
nor U13212 (N_13212,N_12653,N_12655);
nor U13213 (N_13213,N_12782,N_12526);
xnor U13214 (N_13214,N_12855,N_12863);
nand U13215 (N_13215,N_12544,N_12737);
nand U13216 (N_13216,N_12888,N_12538);
nor U13217 (N_13217,N_12695,N_12786);
xor U13218 (N_13218,N_12949,N_12676);
nand U13219 (N_13219,N_12930,N_12907);
nor U13220 (N_13220,N_12652,N_12916);
or U13221 (N_13221,N_12604,N_12552);
or U13222 (N_13222,N_12523,N_12612);
and U13223 (N_13223,N_12978,N_12901);
nand U13224 (N_13224,N_12679,N_12952);
or U13225 (N_13225,N_12501,N_12504);
nor U13226 (N_13226,N_12696,N_12713);
and U13227 (N_13227,N_12543,N_12680);
xnor U13228 (N_13228,N_12773,N_12899);
xnor U13229 (N_13229,N_12760,N_12664);
xnor U13230 (N_13230,N_12752,N_12735);
xor U13231 (N_13231,N_12843,N_12605);
nand U13232 (N_13232,N_12807,N_12783);
or U13233 (N_13233,N_12880,N_12895);
nand U13234 (N_13234,N_12588,N_12599);
or U13235 (N_13235,N_12995,N_12976);
nand U13236 (N_13236,N_12625,N_12643);
and U13237 (N_13237,N_12951,N_12811);
nor U13238 (N_13238,N_12717,N_12962);
xor U13239 (N_13239,N_12565,N_12547);
or U13240 (N_13240,N_12684,N_12668);
nor U13241 (N_13241,N_12682,N_12937);
nand U13242 (N_13242,N_12685,N_12801);
or U13243 (N_13243,N_12981,N_12771);
xnor U13244 (N_13244,N_12792,N_12967);
xor U13245 (N_13245,N_12816,N_12806);
nand U13246 (N_13246,N_12799,N_12877);
nand U13247 (N_13247,N_12704,N_12587);
and U13248 (N_13248,N_12846,N_12789);
nor U13249 (N_13249,N_12663,N_12611);
and U13250 (N_13250,N_12780,N_12957);
nand U13251 (N_13251,N_12598,N_12631);
nor U13252 (N_13252,N_12984,N_12838);
nand U13253 (N_13253,N_12933,N_12827);
nor U13254 (N_13254,N_12748,N_12661);
or U13255 (N_13255,N_12941,N_12554);
nor U13256 (N_13256,N_12853,N_12917);
and U13257 (N_13257,N_12900,N_12718);
and U13258 (N_13258,N_12854,N_12562);
nand U13259 (N_13259,N_12634,N_12941);
nor U13260 (N_13260,N_12914,N_12634);
nand U13261 (N_13261,N_12774,N_12711);
nor U13262 (N_13262,N_12537,N_12777);
xnor U13263 (N_13263,N_12865,N_12709);
and U13264 (N_13264,N_12839,N_12872);
or U13265 (N_13265,N_12875,N_12898);
nand U13266 (N_13266,N_12552,N_12759);
and U13267 (N_13267,N_12866,N_12875);
nor U13268 (N_13268,N_12878,N_12903);
nor U13269 (N_13269,N_12896,N_12701);
nand U13270 (N_13270,N_12563,N_12564);
xor U13271 (N_13271,N_12575,N_12578);
nor U13272 (N_13272,N_12538,N_12611);
xnor U13273 (N_13273,N_12954,N_12588);
or U13274 (N_13274,N_12619,N_12817);
xor U13275 (N_13275,N_12605,N_12548);
and U13276 (N_13276,N_12969,N_12606);
or U13277 (N_13277,N_12960,N_12787);
nor U13278 (N_13278,N_12632,N_12761);
xnor U13279 (N_13279,N_12826,N_12706);
nand U13280 (N_13280,N_12823,N_12940);
or U13281 (N_13281,N_12711,N_12728);
or U13282 (N_13282,N_12536,N_12600);
or U13283 (N_13283,N_12668,N_12679);
nor U13284 (N_13284,N_12893,N_12782);
and U13285 (N_13285,N_12921,N_12788);
nand U13286 (N_13286,N_12780,N_12913);
nor U13287 (N_13287,N_12697,N_12668);
and U13288 (N_13288,N_12691,N_12946);
nand U13289 (N_13289,N_12855,N_12872);
nand U13290 (N_13290,N_12994,N_12538);
xor U13291 (N_13291,N_12919,N_12920);
or U13292 (N_13292,N_12890,N_12951);
and U13293 (N_13293,N_12688,N_12585);
and U13294 (N_13294,N_12981,N_12957);
or U13295 (N_13295,N_12902,N_12805);
xor U13296 (N_13296,N_12606,N_12511);
and U13297 (N_13297,N_12615,N_12616);
nor U13298 (N_13298,N_12876,N_12561);
or U13299 (N_13299,N_12998,N_12712);
and U13300 (N_13300,N_12873,N_12813);
xnor U13301 (N_13301,N_12770,N_12687);
xor U13302 (N_13302,N_12558,N_12815);
xor U13303 (N_13303,N_12611,N_12568);
or U13304 (N_13304,N_12797,N_12557);
or U13305 (N_13305,N_12844,N_12747);
nor U13306 (N_13306,N_12655,N_12868);
or U13307 (N_13307,N_12978,N_12856);
and U13308 (N_13308,N_12881,N_12720);
or U13309 (N_13309,N_12585,N_12506);
and U13310 (N_13310,N_12953,N_12755);
xnor U13311 (N_13311,N_12775,N_12944);
nand U13312 (N_13312,N_12903,N_12504);
nor U13313 (N_13313,N_12769,N_12510);
nand U13314 (N_13314,N_12694,N_12670);
nor U13315 (N_13315,N_12700,N_12570);
and U13316 (N_13316,N_12926,N_12999);
nor U13317 (N_13317,N_12747,N_12666);
and U13318 (N_13318,N_12513,N_12782);
and U13319 (N_13319,N_12816,N_12781);
xnor U13320 (N_13320,N_12558,N_12521);
nand U13321 (N_13321,N_12834,N_12659);
or U13322 (N_13322,N_12605,N_12586);
xnor U13323 (N_13323,N_12984,N_12617);
nand U13324 (N_13324,N_12978,N_12851);
nor U13325 (N_13325,N_12926,N_12992);
xor U13326 (N_13326,N_12502,N_12883);
nand U13327 (N_13327,N_12710,N_12913);
nand U13328 (N_13328,N_12585,N_12997);
nor U13329 (N_13329,N_12591,N_12801);
or U13330 (N_13330,N_12873,N_12553);
or U13331 (N_13331,N_12856,N_12592);
or U13332 (N_13332,N_12510,N_12798);
xnor U13333 (N_13333,N_12581,N_12821);
xnor U13334 (N_13334,N_12674,N_12843);
xor U13335 (N_13335,N_12685,N_12599);
nand U13336 (N_13336,N_12749,N_12968);
nor U13337 (N_13337,N_12614,N_12979);
or U13338 (N_13338,N_12856,N_12698);
or U13339 (N_13339,N_12915,N_12854);
nand U13340 (N_13340,N_12979,N_12732);
or U13341 (N_13341,N_12874,N_12503);
nor U13342 (N_13342,N_12884,N_12637);
nor U13343 (N_13343,N_12616,N_12777);
nand U13344 (N_13344,N_12723,N_12838);
and U13345 (N_13345,N_12868,N_12927);
or U13346 (N_13346,N_12669,N_12748);
nor U13347 (N_13347,N_12766,N_12566);
xor U13348 (N_13348,N_12966,N_12884);
xnor U13349 (N_13349,N_12907,N_12612);
or U13350 (N_13350,N_12628,N_12768);
nand U13351 (N_13351,N_12612,N_12789);
and U13352 (N_13352,N_12920,N_12502);
nor U13353 (N_13353,N_12866,N_12699);
or U13354 (N_13354,N_12638,N_12899);
nor U13355 (N_13355,N_12939,N_12908);
nand U13356 (N_13356,N_12622,N_12755);
xor U13357 (N_13357,N_12849,N_12893);
xnor U13358 (N_13358,N_12909,N_12612);
or U13359 (N_13359,N_12566,N_12808);
nor U13360 (N_13360,N_12875,N_12892);
nand U13361 (N_13361,N_12652,N_12846);
and U13362 (N_13362,N_12770,N_12576);
nand U13363 (N_13363,N_12910,N_12608);
nand U13364 (N_13364,N_12832,N_12780);
and U13365 (N_13365,N_12636,N_12847);
nand U13366 (N_13366,N_12556,N_12533);
and U13367 (N_13367,N_12650,N_12512);
xor U13368 (N_13368,N_12894,N_12873);
or U13369 (N_13369,N_12598,N_12573);
or U13370 (N_13370,N_12569,N_12663);
nand U13371 (N_13371,N_12540,N_12763);
nand U13372 (N_13372,N_12588,N_12868);
nand U13373 (N_13373,N_12608,N_12586);
and U13374 (N_13374,N_12891,N_12639);
nand U13375 (N_13375,N_12576,N_12628);
or U13376 (N_13376,N_12565,N_12678);
nor U13377 (N_13377,N_12765,N_12975);
xnor U13378 (N_13378,N_12876,N_12819);
or U13379 (N_13379,N_12619,N_12872);
nor U13380 (N_13380,N_12989,N_12839);
and U13381 (N_13381,N_12950,N_12792);
xnor U13382 (N_13382,N_12809,N_12649);
xor U13383 (N_13383,N_12590,N_12729);
and U13384 (N_13384,N_12764,N_12954);
and U13385 (N_13385,N_12916,N_12895);
xnor U13386 (N_13386,N_12789,N_12829);
nand U13387 (N_13387,N_12651,N_12743);
and U13388 (N_13388,N_12661,N_12900);
nor U13389 (N_13389,N_12527,N_12637);
nand U13390 (N_13390,N_12746,N_12507);
xnor U13391 (N_13391,N_12715,N_12844);
nor U13392 (N_13392,N_12868,N_12537);
nor U13393 (N_13393,N_12972,N_12635);
nor U13394 (N_13394,N_12846,N_12885);
xnor U13395 (N_13395,N_12975,N_12591);
and U13396 (N_13396,N_12512,N_12905);
and U13397 (N_13397,N_12909,N_12889);
or U13398 (N_13398,N_12710,N_12654);
xnor U13399 (N_13399,N_12733,N_12539);
or U13400 (N_13400,N_12684,N_12872);
nand U13401 (N_13401,N_12573,N_12929);
nor U13402 (N_13402,N_12730,N_12605);
nor U13403 (N_13403,N_12924,N_12704);
nand U13404 (N_13404,N_12532,N_12810);
nor U13405 (N_13405,N_12697,N_12943);
nand U13406 (N_13406,N_12951,N_12523);
nor U13407 (N_13407,N_12768,N_12634);
nor U13408 (N_13408,N_12734,N_12934);
nand U13409 (N_13409,N_12902,N_12515);
nor U13410 (N_13410,N_12948,N_12700);
nand U13411 (N_13411,N_12702,N_12612);
xnor U13412 (N_13412,N_12506,N_12597);
nor U13413 (N_13413,N_12501,N_12759);
nand U13414 (N_13414,N_12708,N_12955);
nor U13415 (N_13415,N_12783,N_12590);
or U13416 (N_13416,N_12958,N_12837);
nand U13417 (N_13417,N_12698,N_12881);
and U13418 (N_13418,N_12857,N_12862);
nand U13419 (N_13419,N_12729,N_12684);
nor U13420 (N_13420,N_12767,N_12635);
nand U13421 (N_13421,N_12879,N_12586);
xnor U13422 (N_13422,N_12885,N_12931);
or U13423 (N_13423,N_12553,N_12766);
nor U13424 (N_13424,N_12990,N_12639);
nor U13425 (N_13425,N_12934,N_12687);
and U13426 (N_13426,N_12961,N_12656);
xor U13427 (N_13427,N_12816,N_12874);
nor U13428 (N_13428,N_12587,N_12733);
nand U13429 (N_13429,N_12800,N_12844);
nor U13430 (N_13430,N_12788,N_12604);
xnor U13431 (N_13431,N_12586,N_12747);
xor U13432 (N_13432,N_12941,N_12961);
and U13433 (N_13433,N_12552,N_12774);
xnor U13434 (N_13434,N_12745,N_12972);
xnor U13435 (N_13435,N_12961,N_12689);
nor U13436 (N_13436,N_12629,N_12708);
nand U13437 (N_13437,N_12742,N_12825);
xnor U13438 (N_13438,N_12813,N_12683);
and U13439 (N_13439,N_12827,N_12948);
nor U13440 (N_13440,N_12722,N_12717);
or U13441 (N_13441,N_12703,N_12944);
nand U13442 (N_13442,N_12977,N_12805);
and U13443 (N_13443,N_12678,N_12958);
or U13444 (N_13444,N_12564,N_12920);
nor U13445 (N_13445,N_12737,N_12692);
and U13446 (N_13446,N_12907,N_12865);
nor U13447 (N_13447,N_12714,N_12731);
nand U13448 (N_13448,N_12767,N_12552);
xor U13449 (N_13449,N_12928,N_12551);
xnor U13450 (N_13450,N_12609,N_12836);
and U13451 (N_13451,N_12507,N_12504);
xor U13452 (N_13452,N_12854,N_12764);
xnor U13453 (N_13453,N_12660,N_12683);
nand U13454 (N_13454,N_12659,N_12661);
or U13455 (N_13455,N_12691,N_12835);
nor U13456 (N_13456,N_12927,N_12756);
or U13457 (N_13457,N_12667,N_12859);
nor U13458 (N_13458,N_12640,N_12556);
nor U13459 (N_13459,N_12879,N_12894);
nor U13460 (N_13460,N_12701,N_12633);
nor U13461 (N_13461,N_12690,N_12698);
xor U13462 (N_13462,N_12613,N_12797);
nand U13463 (N_13463,N_12752,N_12928);
or U13464 (N_13464,N_12887,N_12617);
nor U13465 (N_13465,N_12532,N_12901);
xor U13466 (N_13466,N_12885,N_12611);
or U13467 (N_13467,N_12586,N_12731);
nor U13468 (N_13468,N_12514,N_12746);
or U13469 (N_13469,N_12725,N_12630);
and U13470 (N_13470,N_12589,N_12959);
or U13471 (N_13471,N_12676,N_12537);
and U13472 (N_13472,N_12788,N_12647);
nand U13473 (N_13473,N_12673,N_12728);
nand U13474 (N_13474,N_12879,N_12722);
nor U13475 (N_13475,N_12674,N_12976);
xnor U13476 (N_13476,N_12750,N_12507);
or U13477 (N_13477,N_12757,N_12631);
or U13478 (N_13478,N_12529,N_12827);
xor U13479 (N_13479,N_12823,N_12564);
nand U13480 (N_13480,N_12860,N_12513);
and U13481 (N_13481,N_12923,N_12673);
xor U13482 (N_13482,N_12910,N_12513);
or U13483 (N_13483,N_12547,N_12523);
nand U13484 (N_13484,N_12538,N_12789);
nand U13485 (N_13485,N_12690,N_12897);
nor U13486 (N_13486,N_12837,N_12563);
xnor U13487 (N_13487,N_12863,N_12743);
or U13488 (N_13488,N_12691,N_12793);
or U13489 (N_13489,N_12544,N_12899);
and U13490 (N_13490,N_12899,N_12876);
nand U13491 (N_13491,N_12950,N_12750);
nand U13492 (N_13492,N_12954,N_12894);
nand U13493 (N_13493,N_12865,N_12745);
and U13494 (N_13494,N_12872,N_12672);
and U13495 (N_13495,N_12815,N_12943);
xor U13496 (N_13496,N_12517,N_12953);
xnor U13497 (N_13497,N_12532,N_12564);
and U13498 (N_13498,N_12522,N_12796);
and U13499 (N_13499,N_12825,N_12939);
nor U13500 (N_13500,N_13211,N_13376);
nand U13501 (N_13501,N_13446,N_13384);
or U13502 (N_13502,N_13404,N_13142);
nor U13503 (N_13503,N_13362,N_13472);
nand U13504 (N_13504,N_13412,N_13326);
nand U13505 (N_13505,N_13174,N_13455);
xor U13506 (N_13506,N_13271,N_13347);
nor U13507 (N_13507,N_13284,N_13344);
nor U13508 (N_13508,N_13409,N_13037);
and U13509 (N_13509,N_13015,N_13125);
and U13510 (N_13510,N_13117,N_13439);
xor U13511 (N_13511,N_13110,N_13112);
and U13512 (N_13512,N_13396,N_13169);
and U13513 (N_13513,N_13264,N_13137);
or U13514 (N_13514,N_13474,N_13471);
xnor U13515 (N_13515,N_13225,N_13432);
or U13516 (N_13516,N_13163,N_13028);
and U13517 (N_13517,N_13013,N_13134);
or U13518 (N_13518,N_13490,N_13452);
or U13519 (N_13519,N_13034,N_13051);
and U13520 (N_13520,N_13005,N_13031);
xnor U13521 (N_13521,N_13058,N_13088);
and U13522 (N_13522,N_13178,N_13094);
xnor U13523 (N_13523,N_13065,N_13305);
xor U13524 (N_13524,N_13437,N_13341);
or U13525 (N_13525,N_13444,N_13221);
and U13526 (N_13526,N_13286,N_13235);
xor U13527 (N_13527,N_13045,N_13183);
nand U13528 (N_13528,N_13310,N_13147);
or U13529 (N_13529,N_13441,N_13380);
nand U13530 (N_13530,N_13268,N_13241);
nor U13531 (N_13531,N_13154,N_13230);
or U13532 (N_13532,N_13064,N_13228);
and U13533 (N_13533,N_13208,N_13055);
nand U13534 (N_13534,N_13018,N_13408);
or U13535 (N_13535,N_13070,N_13066);
and U13536 (N_13536,N_13102,N_13056);
xnor U13537 (N_13537,N_13022,N_13373);
nor U13538 (N_13538,N_13085,N_13243);
or U13539 (N_13539,N_13378,N_13379);
nor U13540 (N_13540,N_13090,N_13390);
and U13541 (N_13541,N_13126,N_13000);
or U13542 (N_13542,N_13014,N_13124);
xor U13543 (N_13543,N_13349,N_13003);
and U13544 (N_13544,N_13468,N_13352);
or U13545 (N_13545,N_13012,N_13411);
nor U13546 (N_13546,N_13196,N_13374);
or U13547 (N_13547,N_13114,N_13122);
xor U13548 (N_13548,N_13410,N_13371);
nor U13549 (N_13549,N_13247,N_13044);
and U13550 (N_13550,N_13329,N_13431);
and U13551 (N_13551,N_13233,N_13303);
nand U13552 (N_13552,N_13316,N_13086);
or U13553 (N_13553,N_13442,N_13074);
xor U13554 (N_13554,N_13033,N_13089);
nand U13555 (N_13555,N_13041,N_13350);
and U13556 (N_13556,N_13423,N_13027);
or U13557 (N_13557,N_13291,N_13486);
nor U13558 (N_13558,N_13072,N_13418);
nor U13559 (N_13559,N_13207,N_13226);
and U13560 (N_13560,N_13210,N_13130);
nor U13561 (N_13561,N_13111,N_13091);
xor U13562 (N_13562,N_13253,N_13222);
and U13563 (N_13563,N_13195,N_13375);
xnor U13564 (N_13564,N_13175,N_13068);
or U13565 (N_13565,N_13436,N_13076);
or U13566 (N_13566,N_13330,N_13280);
nand U13567 (N_13567,N_13239,N_13465);
or U13568 (N_13568,N_13340,N_13244);
nor U13569 (N_13569,N_13389,N_13189);
xnor U13570 (N_13570,N_13367,N_13052);
and U13571 (N_13571,N_13319,N_13081);
nand U13572 (N_13572,N_13042,N_13295);
nor U13573 (N_13573,N_13298,N_13359);
nor U13574 (N_13574,N_13311,N_13156);
or U13575 (N_13575,N_13393,N_13201);
and U13576 (N_13576,N_13236,N_13097);
xnor U13577 (N_13577,N_13495,N_13278);
nand U13578 (N_13578,N_13383,N_13182);
xnor U13579 (N_13579,N_13198,N_13323);
nor U13580 (N_13580,N_13498,N_13216);
or U13581 (N_13581,N_13433,N_13108);
nor U13582 (N_13582,N_13395,N_13277);
nand U13583 (N_13583,N_13494,N_13496);
nor U13584 (N_13584,N_13145,N_13036);
nand U13585 (N_13585,N_13219,N_13479);
and U13586 (N_13586,N_13499,N_13484);
nand U13587 (N_13587,N_13351,N_13204);
nand U13588 (N_13588,N_13077,N_13478);
nor U13589 (N_13589,N_13463,N_13132);
nor U13590 (N_13590,N_13205,N_13242);
and U13591 (N_13591,N_13458,N_13129);
nand U13592 (N_13592,N_13335,N_13141);
nor U13593 (N_13593,N_13152,N_13149);
or U13594 (N_13594,N_13366,N_13109);
or U13595 (N_13595,N_13331,N_13165);
nand U13596 (N_13596,N_13318,N_13158);
or U13597 (N_13597,N_13053,N_13238);
nand U13598 (N_13598,N_13203,N_13257);
nor U13599 (N_13599,N_13360,N_13429);
xor U13600 (N_13600,N_13144,N_13231);
nor U13601 (N_13601,N_13427,N_13357);
and U13602 (N_13602,N_13040,N_13385);
or U13603 (N_13603,N_13099,N_13063);
or U13604 (N_13604,N_13260,N_13067);
or U13605 (N_13605,N_13092,N_13100);
or U13606 (N_13606,N_13128,N_13250);
xnor U13607 (N_13607,N_13237,N_13008);
xnor U13608 (N_13608,N_13240,N_13173);
xor U13609 (N_13609,N_13449,N_13309);
or U13610 (N_13610,N_13202,N_13007);
and U13611 (N_13611,N_13197,N_13140);
nand U13612 (N_13612,N_13394,N_13177);
nor U13613 (N_13613,N_13425,N_13200);
nand U13614 (N_13614,N_13026,N_13146);
nor U13615 (N_13615,N_13263,N_13101);
and U13616 (N_13616,N_13413,N_13229);
nor U13617 (N_13617,N_13011,N_13467);
nand U13618 (N_13618,N_13297,N_13180);
and U13619 (N_13619,N_13282,N_13274);
nor U13620 (N_13620,N_13083,N_13107);
nor U13621 (N_13621,N_13029,N_13289);
or U13622 (N_13622,N_13397,N_13120);
xnor U13623 (N_13623,N_13131,N_13377);
nor U13624 (N_13624,N_13262,N_13215);
nand U13625 (N_13625,N_13181,N_13157);
or U13626 (N_13626,N_13285,N_13450);
and U13627 (N_13627,N_13317,N_13459);
xnor U13628 (N_13628,N_13160,N_13294);
nor U13629 (N_13629,N_13296,N_13127);
and U13630 (N_13630,N_13023,N_13401);
and U13631 (N_13631,N_13453,N_13438);
or U13632 (N_13632,N_13030,N_13403);
nand U13633 (N_13633,N_13489,N_13388);
nand U13634 (N_13634,N_13333,N_13392);
or U13635 (N_13635,N_13492,N_13346);
nor U13636 (N_13636,N_13354,N_13312);
nor U13637 (N_13637,N_13258,N_13267);
or U13638 (N_13638,N_13246,N_13348);
nor U13639 (N_13639,N_13416,N_13299);
and U13640 (N_13640,N_13400,N_13161);
nand U13641 (N_13641,N_13324,N_13342);
or U13642 (N_13642,N_13206,N_13159);
nand U13643 (N_13643,N_13186,N_13482);
and U13644 (N_13644,N_13434,N_13473);
nor U13645 (N_13645,N_13422,N_13368);
xor U13646 (N_13646,N_13301,N_13115);
xnor U13647 (N_13647,N_13171,N_13080);
and U13648 (N_13648,N_13475,N_13372);
xnor U13649 (N_13649,N_13456,N_13491);
or U13650 (N_13650,N_13084,N_13287);
or U13651 (N_13651,N_13462,N_13106);
nor U13652 (N_13652,N_13402,N_13304);
and U13653 (N_13653,N_13001,N_13251);
nor U13654 (N_13654,N_13497,N_13188);
or U13655 (N_13655,N_13143,N_13069);
nor U13656 (N_13656,N_13232,N_13071);
and U13657 (N_13657,N_13061,N_13382);
xor U13658 (N_13658,N_13095,N_13481);
xor U13659 (N_13659,N_13424,N_13009);
nor U13660 (N_13660,N_13321,N_13430);
nand U13661 (N_13661,N_13224,N_13136);
nand U13662 (N_13662,N_13098,N_13047);
nand U13663 (N_13663,N_13358,N_13220);
nor U13664 (N_13664,N_13314,N_13279);
nand U13665 (N_13665,N_13488,N_13139);
nand U13666 (N_13666,N_13038,N_13113);
nand U13667 (N_13667,N_13212,N_13315);
and U13668 (N_13668,N_13148,N_13292);
and U13669 (N_13669,N_13199,N_13153);
nand U13670 (N_13670,N_13016,N_13415);
xnor U13671 (N_13671,N_13002,N_13364);
xnor U13672 (N_13672,N_13405,N_13176);
or U13673 (N_13673,N_13328,N_13327);
nor U13674 (N_13674,N_13062,N_13054);
and U13675 (N_13675,N_13477,N_13414);
nor U13676 (N_13676,N_13179,N_13020);
nor U13677 (N_13677,N_13355,N_13320);
xor U13678 (N_13678,N_13363,N_13337);
nand U13679 (N_13679,N_13313,N_13223);
and U13680 (N_13680,N_13259,N_13308);
or U13681 (N_13681,N_13448,N_13060);
and U13682 (N_13682,N_13105,N_13164);
or U13683 (N_13683,N_13075,N_13116);
xnor U13684 (N_13684,N_13048,N_13025);
or U13685 (N_13685,N_13194,N_13184);
nand U13686 (N_13686,N_13435,N_13386);
or U13687 (N_13687,N_13283,N_13187);
nor U13688 (N_13688,N_13461,N_13338);
xnor U13689 (N_13689,N_13276,N_13281);
and U13690 (N_13690,N_13272,N_13133);
nand U13691 (N_13691,N_13391,N_13006);
and U13692 (N_13692,N_13302,N_13227);
nor U13693 (N_13693,N_13353,N_13035);
nor U13694 (N_13694,N_13192,N_13440);
nor U13695 (N_13695,N_13032,N_13356);
or U13696 (N_13696,N_13306,N_13214);
nor U13697 (N_13697,N_13428,N_13217);
nor U13698 (N_13698,N_13234,N_13361);
nand U13699 (N_13699,N_13454,N_13046);
and U13700 (N_13700,N_13336,N_13370);
and U13701 (N_13701,N_13103,N_13082);
or U13702 (N_13702,N_13050,N_13447);
and U13703 (N_13703,N_13343,N_13104);
nand U13704 (N_13704,N_13079,N_13339);
and U13705 (N_13705,N_13420,N_13256);
nor U13706 (N_13706,N_13162,N_13254);
and U13707 (N_13707,N_13172,N_13151);
xnor U13708 (N_13708,N_13073,N_13121);
nand U13709 (N_13709,N_13213,N_13261);
nand U13710 (N_13710,N_13460,N_13039);
nand U13711 (N_13711,N_13270,N_13480);
and U13712 (N_13712,N_13168,N_13406);
and U13713 (N_13713,N_13381,N_13445);
nand U13714 (N_13714,N_13476,N_13119);
or U13715 (N_13715,N_13248,N_13255);
and U13716 (N_13716,N_13334,N_13387);
and U13717 (N_13717,N_13369,N_13193);
xnor U13718 (N_13718,N_13123,N_13487);
nand U13719 (N_13719,N_13059,N_13024);
and U13720 (N_13720,N_13096,N_13470);
xor U13721 (N_13721,N_13275,N_13307);
and U13722 (N_13722,N_13483,N_13266);
or U13723 (N_13723,N_13087,N_13293);
or U13724 (N_13724,N_13300,N_13170);
xnor U13725 (N_13725,N_13325,N_13190);
xor U13726 (N_13726,N_13078,N_13464);
and U13727 (N_13727,N_13043,N_13218);
and U13728 (N_13728,N_13150,N_13245);
and U13729 (N_13729,N_13421,N_13451);
or U13730 (N_13730,N_13118,N_13345);
xor U13731 (N_13731,N_13273,N_13407);
xnor U13732 (N_13732,N_13269,N_13167);
xnor U13733 (N_13733,N_13290,N_13365);
xnor U13734 (N_13734,N_13426,N_13252);
xor U13735 (N_13735,N_13019,N_13443);
nand U13736 (N_13736,N_13049,N_13419);
nor U13737 (N_13737,N_13185,N_13417);
or U13738 (N_13738,N_13332,N_13485);
nand U13739 (N_13739,N_13249,N_13399);
nand U13740 (N_13740,N_13466,N_13138);
and U13741 (N_13741,N_13166,N_13021);
nor U13742 (N_13742,N_13469,N_13191);
or U13743 (N_13743,N_13493,N_13093);
xor U13744 (N_13744,N_13135,N_13288);
nor U13745 (N_13745,N_13457,N_13322);
and U13746 (N_13746,N_13398,N_13017);
or U13747 (N_13747,N_13057,N_13265);
nor U13748 (N_13748,N_13209,N_13155);
xor U13749 (N_13749,N_13004,N_13010);
xnor U13750 (N_13750,N_13153,N_13007);
xor U13751 (N_13751,N_13104,N_13242);
nor U13752 (N_13752,N_13263,N_13415);
xnor U13753 (N_13753,N_13064,N_13320);
or U13754 (N_13754,N_13458,N_13132);
xnor U13755 (N_13755,N_13270,N_13015);
nor U13756 (N_13756,N_13362,N_13113);
and U13757 (N_13757,N_13416,N_13257);
nor U13758 (N_13758,N_13118,N_13053);
or U13759 (N_13759,N_13405,N_13147);
nor U13760 (N_13760,N_13032,N_13364);
xor U13761 (N_13761,N_13226,N_13029);
or U13762 (N_13762,N_13250,N_13089);
nor U13763 (N_13763,N_13453,N_13110);
nand U13764 (N_13764,N_13255,N_13212);
nand U13765 (N_13765,N_13458,N_13411);
and U13766 (N_13766,N_13199,N_13057);
xor U13767 (N_13767,N_13208,N_13466);
and U13768 (N_13768,N_13044,N_13341);
nor U13769 (N_13769,N_13112,N_13447);
or U13770 (N_13770,N_13109,N_13007);
xor U13771 (N_13771,N_13054,N_13163);
nor U13772 (N_13772,N_13024,N_13096);
xnor U13773 (N_13773,N_13145,N_13499);
nand U13774 (N_13774,N_13053,N_13027);
and U13775 (N_13775,N_13018,N_13211);
and U13776 (N_13776,N_13401,N_13353);
or U13777 (N_13777,N_13052,N_13387);
nand U13778 (N_13778,N_13414,N_13179);
xnor U13779 (N_13779,N_13077,N_13494);
or U13780 (N_13780,N_13170,N_13488);
and U13781 (N_13781,N_13277,N_13183);
and U13782 (N_13782,N_13318,N_13065);
and U13783 (N_13783,N_13380,N_13145);
nor U13784 (N_13784,N_13061,N_13102);
nand U13785 (N_13785,N_13185,N_13344);
nor U13786 (N_13786,N_13066,N_13450);
and U13787 (N_13787,N_13327,N_13159);
and U13788 (N_13788,N_13113,N_13305);
nor U13789 (N_13789,N_13004,N_13065);
nand U13790 (N_13790,N_13257,N_13007);
xor U13791 (N_13791,N_13135,N_13470);
nand U13792 (N_13792,N_13103,N_13072);
nand U13793 (N_13793,N_13078,N_13228);
nor U13794 (N_13794,N_13292,N_13014);
or U13795 (N_13795,N_13141,N_13043);
nand U13796 (N_13796,N_13370,N_13429);
and U13797 (N_13797,N_13010,N_13378);
xnor U13798 (N_13798,N_13305,N_13248);
xor U13799 (N_13799,N_13405,N_13394);
or U13800 (N_13800,N_13255,N_13245);
xnor U13801 (N_13801,N_13153,N_13346);
or U13802 (N_13802,N_13127,N_13004);
nor U13803 (N_13803,N_13067,N_13315);
nand U13804 (N_13804,N_13038,N_13294);
nand U13805 (N_13805,N_13388,N_13387);
nor U13806 (N_13806,N_13069,N_13280);
nand U13807 (N_13807,N_13423,N_13441);
and U13808 (N_13808,N_13052,N_13294);
or U13809 (N_13809,N_13461,N_13362);
xor U13810 (N_13810,N_13465,N_13154);
nand U13811 (N_13811,N_13172,N_13480);
xnor U13812 (N_13812,N_13248,N_13428);
or U13813 (N_13813,N_13117,N_13240);
nand U13814 (N_13814,N_13192,N_13268);
or U13815 (N_13815,N_13423,N_13280);
xor U13816 (N_13816,N_13056,N_13496);
and U13817 (N_13817,N_13043,N_13278);
and U13818 (N_13818,N_13400,N_13463);
nor U13819 (N_13819,N_13088,N_13400);
xor U13820 (N_13820,N_13196,N_13000);
or U13821 (N_13821,N_13220,N_13292);
nand U13822 (N_13822,N_13380,N_13386);
nor U13823 (N_13823,N_13125,N_13456);
or U13824 (N_13824,N_13239,N_13324);
nand U13825 (N_13825,N_13373,N_13443);
nor U13826 (N_13826,N_13363,N_13227);
and U13827 (N_13827,N_13191,N_13440);
and U13828 (N_13828,N_13238,N_13490);
and U13829 (N_13829,N_13488,N_13273);
or U13830 (N_13830,N_13437,N_13242);
xor U13831 (N_13831,N_13081,N_13013);
or U13832 (N_13832,N_13223,N_13057);
xnor U13833 (N_13833,N_13428,N_13448);
nor U13834 (N_13834,N_13168,N_13085);
nor U13835 (N_13835,N_13378,N_13020);
and U13836 (N_13836,N_13255,N_13400);
nor U13837 (N_13837,N_13474,N_13371);
xor U13838 (N_13838,N_13218,N_13046);
xnor U13839 (N_13839,N_13246,N_13404);
and U13840 (N_13840,N_13013,N_13140);
nand U13841 (N_13841,N_13480,N_13492);
xor U13842 (N_13842,N_13260,N_13212);
or U13843 (N_13843,N_13445,N_13098);
nand U13844 (N_13844,N_13083,N_13251);
or U13845 (N_13845,N_13027,N_13025);
and U13846 (N_13846,N_13098,N_13198);
xnor U13847 (N_13847,N_13341,N_13452);
nand U13848 (N_13848,N_13460,N_13267);
nor U13849 (N_13849,N_13425,N_13380);
xor U13850 (N_13850,N_13454,N_13437);
and U13851 (N_13851,N_13176,N_13002);
and U13852 (N_13852,N_13090,N_13187);
xnor U13853 (N_13853,N_13285,N_13002);
xor U13854 (N_13854,N_13066,N_13412);
and U13855 (N_13855,N_13326,N_13266);
and U13856 (N_13856,N_13363,N_13107);
nor U13857 (N_13857,N_13425,N_13484);
nand U13858 (N_13858,N_13398,N_13238);
or U13859 (N_13859,N_13395,N_13365);
xnor U13860 (N_13860,N_13411,N_13187);
nand U13861 (N_13861,N_13471,N_13099);
and U13862 (N_13862,N_13011,N_13324);
or U13863 (N_13863,N_13043,N_13142);
xor U13864 (N_13864,N_13247,N_13288);
or U13865 (N_13865,N_13492,N_13117);
nor U13866 (N_13866,N_13487,N_13170);
and U13867 (N_13867,N_13082,N_13201);
nand U13868 (N_13868,N_13241,N_13328);
xnor U13869 (N_13869,N_13305,N_13418);
or U13870 (N_13870,N_13133,N_13343);
nor U13871 (N_13871,N_13302,N_13132);
or U13872 (N_13872,N_13220,N_13026);
nor U13873 (N_13873,N_13470,N_13073);
and U13874 (N_13874,N_13437,N_13019);
xnor U13875 (N_13875,N_13060,N_13233);
and U13876 (N_13876,N_13219,N_13067);
and U13877 (N_13877,N_13080,N_13345);
nand U13878 (N_13878,N_13142,N_13125);
xor U13879 (N_13879,N_13234,N_13331);
xnor U13880 (N_13880,N_13160,N_13201);
and U13881 (N_13881,N_13305,N_13189);
nand U13882 (N_13882,N_13310,N_13119);
and U13883 (N_13883,N_13233,N_13476);
nand U13884 (N_13884,N_13325,N_13000);
nor U13885 (N_13885,N_13183,N_13084);
or U13886 (N_13886,N_13359,N_13482);
nand U13887 (N_13887,N_13414,N_13392);
and U13888 (N_13888,N_13362,N_13423);
xnor U13889 (N_13889,N_13035,N_13470);
or U13890 (N_13890,N_13445,N_13179);
nor U13891 (N_13891,N_13179,N_13325);
nor U13892 (N_13892,N_13443,N_13055);
and U13893 (N_13893,N_13290,N_13330);
xor U13894 (N_13894,N_13200,N_13286);
and U13895 (N_13895,N_13418,N_13458);
nor U13896 (N_13896,N_13271,N_13453);
nor U13897 (N_13897,N_13170,N_13342);
nand U13898 (N_13898,N_13148,N_13107);
nor U13899 (N_13899,N_13208,N_13043);
and U13900 (N_13900,N_13223,N_13006);
xor U13901 (N_13901,N_13271,N_13450);
nor U13902 (N_13902,N_13054,N_13219);
nor U13903 (N_13903,N_13044,N_13343);
xor U13904 (N_13904,N_13256,N_13236);
xor U13905 (N_13905,N_13092,N_13408);
and U13906 (N_13906,N_13219,N_13087);
and U13907 (N_13907,N_13466,N_13137);
nand U13908 (N_13908,N_13295,N_13262);
xnor U13909 (N_13909,N_13335,N_13339);
xnor U13910 (N_13910,N_13386,N_13223);
nor U13911 (N_13911,N_13048,N_13351);
or U13912 (N_13912,N_13116,N_13341);
xor U13913 (N_13913,N_13423,N_13287);
or U13914 (N_13914,N_13071,N_13237);
nor U13915 (N_13915,N_13129,N_13184);
nor U13916 (N_13916,N_13059,N_13409);
and U13917 (N_13917,N_13477,N_13178);
or U13918 (N_13918,N_13253,N_13261);
and U13919 (N_13919,N_13048,N_13355);
and U13920 (N_13920,N_13242,N_13308);
nand U13921 (N_13921,N_13180,N_13113);
or U13922 (N_13922,N_13273,N_13380);
and U13923 (N_13923,N_13044,N_13372);
nor U13924 (N_13924,N_13438,N_13049);
xor U13925 (N_13925,N_13211,N_13222);
nand U13926 (N_13926,N_13049,N_13397);
nand U13927 (N_13927,N_13423,N_13068);
and U13928 (N_13928,N_13392,N_13189);
nor U13929 (N_13929,N_13387,N_13013);
or U13930 (N_13930,N_13171,N_13357);
xor U13931 (N_13931,N_13423,N_13306);
nor U13932 (N_13932,N_13022,N_13179);
nand U13933 (N_13933,N_13294,N_13237);
nor U13934 (N_13934,N_13040,N_13296);
and U13935 (N_13935,N_13113,N_13332);
nor U13936 (N_13936,N_13468,N_13126);
xor U13937 (N_13937,N_13392,N_13229);
or U13938 (N_13938,N_13100,N_13037);
nand U13939 (N_13939,N_13142,N_13250);
nor U13940 (N_13940,N_13386,N_13147);
and U13941 (N_13941,N_13017,N_13191);
xnor U13942 (N_13942,N_13374,N_13204);
xnor U13943 (N_13943,N_13182,N_13117);
nand U13944 (N_13944,N_13317,N_13398);
nand U13945 (N_13945,N_13433,N_13361);
or U13946 (N_13946,N_13354,N_13483);
and U13947 (N_13947,N_13329,N_13164);
xor U13948 (N_13948,N_13112,N_13132);
xor U13949 (N_13949,N_13326,N_13057);
and U13950 (N_13950,N_13292,N_13397);
and U13951 (N_13951,N_13082,N_13163);
nand U13952 (N_13952,N_13113,N_13196);
xor U13953 (N_13953,N_13325,N_13320);
nand U13954 (N_13954,N_13458,N_13030);
and U13955 (N_13955,N_13071,N_13233);
nor U13956 (N_13956,N_13329,N_13165);
or U13957 (N_13957,N_13070,N_13145);
xnor U13958 (N_13958,N_13102,N_13345);
nand U13959 (N_13959,N_13236,N_13246);
or U13960 (N_13960,N_13427,N_13119);
xor U13961 (N_13961,N_13107,N_13468);
nor U13962 (N_13962,N_13389,N_13460);
and U13963 (N_13963,N_13190,N_13422);
nor U13964 (N_13964,N_13096,N_13455);
and U13965 (N_13965,N_13205,N_13449);
nor U13966 (N_13966,N_13194,N_13420);
nand U13967 (N_13967,N_13030,N_13376);
nor U13968 (N_13968,N_13482,N_13138);
or U13969 (N_13969,N_13222,N_13380);
xnor U13970 (N_13970,N_13212,N_13074);
xor U13971 (N_13971,N_13019,N_13351);
nor U13972 (N_13972,N_13400,N_13368);
or U13973 (N_13973,N_13252,N_13130);
nand U13974 (N_13974,N_13035,N_13181);
or U13975 (N_13975,N_13291,N_13382);
xnor U13976 (N_13976,N_13208,N_13396);
or U13977 (N_13977,N_13308,N_13026);
and U13978 (N_13978,N_13251,N_13016);
nand U13979 (N_13979,N_13482,N_13261);
xor U13980 (N_13980,N_13269,N_13096);
or U13981 (N_13981,N_13258,N_13070);
nand U13982 (N_13982,N_13379,N_13300);
xnor U13983 (N_13983,N_13151,N_13108);
or U13984 (N_13984,N_13124,N_13142);
and U13985 (N_13985,N_13014,N_13246);
nor U13986 (N_13986,N_13128,N_13308);
xnor U13987 (N_13987,N_13226,N_13250);
nor U13988 (N_13988,N_13146,N_13270);
nand U13989 (N_13989,N_13049,N_13292);
xnor U13990 (N_13990,N_13104,N_13454);
and U13991 (N_13991,N_13268,N_13012);
nor U13992 (N_13992,N_13139,N_13330);
and U13993 (N_13993,N_13494,N_13453);
nor U13994 (N_13994,N_13319,N_13465);
nor U13995 (N_13995,N_13334,N_13416);
xnor U13996 (N_13996,N_13349,N_13268);
nand U13997 (N_13997,N_13126,N_13372);
nand U13998 (N_13998,N_13471,N_13302);
nand U13999 (N_13999,N_13253,N_13315);
nand U14000 (N_14000,N_13942,N_13768);
and U14001 (N_14001,N_13597,N_13918);
and U14002 (N_14002,N_13874,N_13781);
or U14003 (N_14003,N_13542,N_13527);
nor U14004 (N_14004,N_13878,N_13714);
and U14005 (N_14005,N_13790,N_13538);
or U14006 (N_14006,N_13723,N_13706);
xor U14007 (N_14007,N_13530,N_13823);
and U14008 (N_14008,N_13633,N_13951);
or U14009 (N_14009,N_13883,N_13871);
or U14010 (N_14010,N_13931,N_13970);
and U14011 (N_14011,N_13812,N_13519);
xor U14012 (N_14012,N_13701,N_13943);
xor U14013 (N_14013,N_13602,N_13989);
or U14014 (N_14014,N_13501,N_13939);
or U14015 (N_14015,N_13867,N_13570);
nor U14016 (N_14016,N_13741,N_13980);
nor U14017 (N_14017,N_13832,N_13656);
or U14018 (N_14018,N_13627,N_13872);
or U14019 (N_14019,N_13803,N_13712);
xor U14020 (N_14020,N_13668,N_13699);
nand U14021 (N_14021,N_13652,N_13583);
nand U14022 (N_14022,N_13830,N_13503);
nor U14023 (N_14023,N_13685,N_13740);
nor U14024 (N_14024,N_13692,N_13808);
nor U14025 (N_14025,N_13585,N_13581);
and U14026 (N_14026,N_13713,N_13601);
nor U14027 (N_14027,N_13885,N_13654);
nor U14028 (N_14028,N_13716,N_13935);
and U14029 (N_14029,N_13901,N_13956);
or U14030 (N_14030,N_13502,N_13590);
xnor U14031 (N_14031,N_13750,N_13689);
and U14032 (N_14032,N_13974,N_13531);
and U14033 (N_14033,N_13695,N_13578);
and U14034 (N_14034,N_13975,N_13926);
nor U14035 (N_14035,N_13797,N_13947);
and U14036 (N_14036,N_13743,N_13671);
or U14037 (N_14037,N_13659,N_13670);
or U14038 (N_14038,N_13655,N_13893);
and U14039 (N_14039,N_13933,N_13968);
and U14040 (N_14040,N_13576,N_13981);
nor U14041 (N_14041,N_13603,N_13908);
nand U14042 (N_14042,N_13810,N_13988);
or U14043 (N_14043,N_13866,N_13860);
and U14044 (N_14044,N_13841,N_13573);
and U14045 (N_14045,N_13562,N_13802);
xnor U14046 (N_14046,N_13754,N_13653);
xnor U14047 (N_14047,N_13642,N_13928);
or U14048 (N_14048,N_13535,N_13514);
nor U14049 (N_14049,N_13813,N_13709);
and U14050 (N_14050,N_13911,N_13814);
nor U14051 (N_14051,N_13651,N_13500);
and U14052 (N_14052,N_13842,N_13611);
or U14053 (N_14053,N_13715,N_13846);
or U14054 (N_14054,N_13676,N_13595);
xnor U14055 (N_14055,N_13669,N_13824);
and U14056 (N_14056,N_13887,N_13621);
or U14057 (N_14057,N_13745,N_13752);
and U14058 (N_14058,N_13698,N_13532);
and U14059 (N_14059,N_13959,N_13732);
or U14060 (N_14060,N_13879,N_13641);
nand U14061 (N_14061,N_13835,N_13977);
and U14062 (N_14062,N_13792,N_13575);
xor U14063 (N_14063,N_13884,N_13877);
nand U14064 (N_14064,N_13799,N_13748);
and U14065 (N_14065,N_13609,N_13546);
nor U14066 (N_14066,N_13663,N_13529);
nand U14067 (N_14067,N_13906,N_13693);
or U14068 (N_14068,N_13782,N_13675);
and U14069 (N_14069,N_13735,N_13628);
or U14070 (N_14070,N_13869,N_13617);
nand U14071 (N_14071,N_13775,N_13967);
nor U14072 (N_14072,N_13518,N_13862);
and U14073 (N_14073,N_13978,N_13673);
xor U14074 (N_14074,N_13798,N_13684);
nor U14075 (N_14075,N_13647,N_13734);
nand U14076 (N_14076,N_13858,N_13553);
nor U14077 (N_14077,N_13672,N_13572);
or U14078 (N_14078,N_13686,N_13955);
nor U14079 (N_14079,N_13786,N_13904);
and U14080 (N_14080,N_13929,N_13515);
xnor U14081 (N_14081,N_13800,N_13596);
and U14082 (N_14082,N_13919,N_13605);
and U14083 (N_14083,N_13854,N_13594);
nor U14084 (N_14084,N_13600,N_13963);
xor U14085 (N_14085,N_13667,N_13536);
and U14086 (N_14086,N_13848,N_13707);
or U14087 (N_14087,N_13746,N_13767);
and U14088 (N_14088,N_13725,N_13625);
nor U14089 (N_14089,N_13571,N_13779);
xnor U14090 (N_14090,N_13903,N_13526);
xor U14091 (N_14091,N_13944,N_13751);
xor U14092 (N_14092,N_13839,N_13843);
nand U14093 (N_14093,N_13704,N_13623);
nand U14094 (N_14094,N_13856,N_13837);
or U14095 (N_14095,N_13662,N_13639);
nor U14096 (N_14096,N_13722,N_13622);
xnor U14097 (N_14097,N_13691,N_13569);
nand U14098 (N_14098,N_13785,N_13838);
or U14099 (N_14099,N_13508,N_13936);
xor U14100 (N_14100,N_13731,N_13938);
nor U14101 (N_14101,N_13550,N_13637);
nand U14102 (N_14102,N_13993,N_13923);
nor U14103 (N_14103,N_13624,N_13630);
nor U14104 (N_14104,N_13859,N_13608);
xnor U14105 (N_14105,N_13506,N_13907);
or U14106 (N_14106,N_13773,N_13537);
nor U14107 (N_14107,N_13765,N_13934);
and U14108 (N_14108,N_13520,N_13729);
xor U14109 (N_14109,N_13787,N_13916);
or U14110 (N_14110,N_13836,N_13755);
nor U14111 (N_14111,N_13645,N_13940);
and U14112 (N_14112,N_13636,N_13616);
and U14113 (N_14113,N_13969,N_13772);
nor U14114 (N_14114,N_13552,N_13761);
xnor U14115 (N_14115,N_13703,N_13644);
xnor U14116 (N_14116,N_13849,N_13949);
or U14117 (N_14117,N_13966,N_13852);
or U14118 (N_14118,N_13718,N_13945);
or U14119 (N_14119,N_13646,N_13991);
and U14120 (N_14120,N_13795,N_13957);
nor U14121 (N_14121,N_13793,N_13658);
or U14122 (N_14122,N_13868,N_13778);
nand U14123 (N_14123,N_13902,N_13556);
and U14124 (N_14124,N_13894,N_13829);
xor U14125 (N_14125,N_13899,N_13555);
or U14126 (N_14126,N_13598,N_13816);
nand U14127 (N_14127,N_13998,N_13632);
xor U14128 (N_14128,N_13547,N_13626);
nand U14129 (N_14129,N_13864,N_13584);
or U14130 (N_14130,N_13720,N_13891);
xnor U14131 (N_14131,N_13582,N_13548);
nand U14132 (N_14132,N_13777,N_13612);
and U14133 (N_14133,N_13567,N_13540);
and U14134 (N_14134,N_13726,N_13888);
or U14135 (N_14135,N_13995,N_13912);
nor U14136 (N_14136,N_13560,N_13972);
or U14137 (N_14137,N_13523,N_13807);
xor U14138 (N_14138,N_13946,N_13660);
nor U14139 (N_14139,N_13880,N_13640);
nand U14140 (N_14140,N_13589,N_13804);
xnor U14141 (N_14141,N_13805,N_13861);
and U14142 (N_14142,N_13833,N_13948);
xor U14143 (N_14143,N_13564,N_13756);
nand U14144 (N_14144,N_13965,N_13516);
or U14145 (N_14145,N_13764,N_13840);
nand U14146 (N_14146,N_13610,N_13788);
nor U14147 (N_14147,N_13762,N_13818);
nand U14148 (N_14148,N_13976,N_13952);
nand U14149 (N_14149,N_13924,N_13747);
and U14150 (N_14150,N_13789,N_13638);
or U14151 (N_14151,N_13753,N_13758);
or U14152 (N_14152,N_13708,N_13607);
nor U14153 (N_14153,N_13844,N_13763);
nor U14154 (N_14154,N_13736,N_13511);
and U14155 (N_14155,N_13791,N_13834);
nor U14156 (N_14156,N_13766,N_13950);
or U14157 (N_14157,N_13588,N_13574);
or U14158 (N_14158,N_13558,N_13524);
nand U14159 (N_14159,N_13727,N_13504);
nand U14160 (N_14160,N_13634,N_13982);
and U14161 (N_14161,N_13629,N_13681);
xor U14162 (N_14162,N_13784,N_13661);
and U14163 (N_14163,N_13865,N_13831);
or U14164 (N_14164,N_13910,N_13643);
nor U14165 (N_14165,N_13783,N_13739);
nand U14166 (N_14166,N_13717,N_13987);
or U14167 (N_14167,N_13618,N_13921);
nand U14168 (N_14168,N_13566,N_13683);
nor U14169 (N_14169,N_13730,N_13892);
or U14170 (N_14170,N_13870,N_13915);
and U14171 (N_14171,N_13507,N_13724);
xor U14172 (N_14172,N_13677,N_13996);
nor U14173 (N_14173,N_13544,N_13826);
nand U14174 (N_14174,N_13897,N_13528);
or U14175 (N_14175,N_13710,N_13593);
and U14176 (N_14176,N_13809,N_13577);
or U14177 (N_14177,N_13682,N_13889);
xnor U14178 (N_14178,N_13999,N_13845);
xor U14179 (N_14179,N_13979,N_13759);
nand U14180 (N_14180,N_13591,N_13971);
nor U14181 (N_14181,N_13563,N_13780);
nor U14182 (N_14182,N_13983,N_13925);
xnor U14183 (N_14183,N_13522,N_13875);
nor U14184 (N_14184,N_13757,N_13819);
nand U14185 (N_14185,N_13992,N_13954);
and U14186 (N_14186,N_13962,N_13895);
or U14187 (N_14187,N_13650,N_13820);
or U14188 (N_14188,N_13850,N_13517);
nor U14189 (N_14189,N_13737,N_13909);
xnor U14190 (N_14190,N_13941,N_13690);
nand U14191 (N_14191,N_13886,N_13985);
xor U14192 (N_14192,N_13964,N_13990);
nor U14193 (N_14193,N_13890,N_13917);
or U14194 (N_14194,N_13873,N_13657);
nand U14195 (N_14195,N_13920,N_13525);
xnor U14196 (N_14196,N_13680,N_13635);
nand U14197 (N_14197,N_13801,N_13696);
and U14198 (N_14198,N_13711,N_13827);
xnor U14199 (N_14199,N_13825,N_13847);
nor U14200 (N_14200,N_13559,N_13688);
nand U14201 (N_14201,N_13619,N_13705);
nand U14202 (N_14202,N_13769,N_13543);
and U14203 (N_14203,N_13606,N_13937);
or U14204 (N_14204,N_13822,N_13953);
or U14205 (N_14205,N_13545,N_13579);
xor U14206 (N_14206,N_13586,N_13534);
or U14207 (N_14207,N_13927,N_13876);
nor U14208 (N_14208,N_13742,N_13719);
and U14209 (N_14209,N_13994,N_13817);
nor U14210 (N_14210,N_13986,N_13881);
nor U14211 (N_14211,N_13806,N_13700);
xnor U14212 (N_14212,N_13749,N_13896);
xnor U14213 (N_14213,N_13811,N_13674);
and U14214 (N_14214,N_13580,N_13679);
xnor U14215 (N_14215,N_13549,N_13561);
or U14216 (N_14216,N_13771,N_13855);
xor U14217 (N_14217,N_13554,N_13857);
nor U14218 (N_14218,N_13851,N_13760);
xor U14219 (N_14219,N_13882,N_13853);
and U14220 (N_14220,N_13512,N_13551);
nand U14221 (N_14221,N_13702,N_13678);
and U14222 (N_14222,N_13649,N_13922);
nand U14223 (N_14223,N_13863,N_13620);
nor U14224 (N_14224,N_13694,N_13541);
and U14225 (N_14225,N_13592,N_13905);
nand U14226 (N_14226,N_13900,N_13776);
nor U14227 (N_14227,N_13973,N_13587);
xor U14228 (N_14228,N_13599,N_13774);
or U14229 (N_14229,N_13664,N_13614);
or U14230 (N_14230,N_13697,N_13568);
or U14231 (N_14231,N_13932,N_13539);
and U14232 (N_14232,N_13557,N_13721);
nor U14233 (N_14233,N_13509,N_13533);
or U14234 (N_14234,N_13665,N_13821);
nand U14235 (N_14235,N_13666,N_13794);
xnor U14236 (N_14236,N_13505,N_13958);
or U14237 (N_14237,N_13898,N_13648);
and U14238 (N_14238,N_13997,N_13738);
xor U14239 (N_14239,N_13961,N_13510);
nor U14240 (N_14240,N_13913,N_13728);
nor U14241 (N_14241,N_13828,N_13613);
xnor U14242 (N_14242,N_13815,N_13914);
or U14243 (N_14243,N_13565,N_13604);
xnor U14244 (N_14244,N_13770,N_13631);
xor U14245 (N_14245,N_13984,N_13960);
nor U14246 (N_14246,N_13744,N_13687);
nand U14247 (N_14247,N_13733,N_13513);
xnor U14248 (N_14248,N_13615,N_13521);
or U14249 (N_14249,N_13796,N_13930);
xnor U14250 (N_14250,N_13986,N_13889);
and U14251 (N_14251,N_13646,N_13615);
nor U14252 (N_14252,N_13743,N_13742);
or U14253 (N_14253,N_13868,N_13934);
nor U14254 (N_14254,N_13535,N_13721);
xnor U14255 (N_14255,N_13533,N_13581);
or U14256 (N_14256,N_13812,N_13697);
xnor U14257 (N_14257,N_13795,N_13931);
nand U14258 (N_14258,N_13507,N_13692);
nor U14259 (N_14259,N_13616,N_13980);
nor U14260 (N_14260,N_13606,N_13645);
xor U14261 (N_14261,N_13732,N_13874);
nor U14262 (N_14262,N_13716,N_13544);
nand U14263 (N_14263,N_13694,N_13761);
or U14264 (N_14264,N_13646,N_13544);
nor U14265 (N_14265,N_13568,N_13716);
xor U14266 (N_14266,N_13999,N_13585);
xor U14267 (N_14267,N_13825,N_13869);
nand U14268 (N_14268,N_13991,N_13892);
nand U14269 (N_14269,N_13891,N_13822);
and U14270 (N_14270,N_13837,N_13984);
and U14271 (N_14271,N_13632,N_13690);
and U14272 (N_14272,N_13824,N_13522);
or U14273 (N_14273,N_13574,N_13744);
xnor U14274 (N_14274,N_13892,N_13863);
and U14275 (N_14275,N_13598,N_13892);
and U14276 (N_14276,N_13929,N_13502);
or U14277 (N_14277,N_13581,N_13907);
nand U14278 (N_14278,N_13724,N_13675);
and U14279 (N_14279,N_13842,N_13824);
xnor U14280 (N_14280,N_13776,N_13548);
or U14281 (N_14281,N_13534,N_13713);
xor U14282 (N_14282,N_13552,N_13660);
xnor U14283 (N_14283,N_13890,N_13676);
xnor U14284 (N_14284,N_13547,N_13589);
xor U14285 (N_14285,N_13661,N_13933);
and U14286 (N_14286,N_13759,N_13646);
and U14287 (N_14287,N_13739,N_13908);
and U14288 (N_14288,N_13822,N_13713);
nor U14289 (N_14289,N_13596,N_13938);
xnor U14290 (N_14290,N_13880,N_13579);
xnor U14291 (N_14291,N_13694,N_13988);
or U14292 (N_14292,N_13855,N_13635);
nor U14293 (N_14293,N_13642,N_13636);
nor U14294 (N_14294,N_13804,N_13590);
and U14295 (N_14295,N_13856,N_13589);
xnor U14296 (N_14296,N_13757,N_13754);
or U14297 (N_14297,N_13884,N_13813);
xor U14298 (N_14298,N_13894,N_13908);
nor U14299 (N_14299,N_13618,N_13865);
nand U14300 (N_14300,N_13787,N_13820);
xor U14301 (N_14301,N_13854,N_13816);
or U14302 (N_14302,N_13744,N_13853);
or U14303 (N_14303,N_13895,N_13745);
nor U14304 (N_14304,N_13541,N_13501);
or U14305 (N_14305,N_13975,N_13660);
nand U14306 (N_14306,N_13552,N_13998);
or U14307 (N_14307,N_13975,N_13508);
nor U14308 (N_14308,N_13899,N_13986);
nor U14309 (N_14309,N_13955,N_13893);
xnor U14310 (N_14310,N_13712,N_13665);
nor U14311 (N_14311,N_13662,N_13661);
nand U14312 (N_14312,N_13956,N_13615);
nand U14313 (N_14313,N_13671,N_13581);
or U14314 (N_14314,N_13898,N_13754);
and U14315 (N_14315,N_13655,N_13540);
nand U14316 (N_14316,N_13994,N_13689);
nor U14317 (N_14317,N_13500,N_13965);
nand U14318 (N_14318,N_13670,N_13688);
or U14319 (N_14319,N_13804,N_13756);
xor U14320 (N_14320,N_13743,N_13588);
nand U14321 (N_14321,N_13719,N_13991);
and U14322 (N_14322,N_13552,N_13773);
nand U14323 (N_14323,N_13818,N_13566);
nand U14324 (N_14324,N_13554,N_13537);
nand U14325 (N_14325,N_13560,N_13724);
xor U14326 (N_14326,N_13783,N_13646);
or U14327 (N_14327,N_13889,N_13669);
nor U14328 (N_14328,N_13623,N_13672);
nor U14329 (N_14329,N_13823,N_13852);
xor U14330 (N_14330,N_13900,N_13815);
nor U14331 (N_14331,N_13925,N_13765);
and U14332 (N_14332,N_13999,N_13888);
or U14333 (N_14333,N_13879,N_13978);
xnor U14334 (N_14334,N_13500,N_13803);
nand U14335 (N_14335,N_13938,N_13554);
nand U14336 (N_14336,N_13596,N_13522);
or U14337 (N_14337,N_13872,N_13890);
xnor U14338 (N_14338,N_13792,N_13571);
or U14339 (N_14339,N_13586,N_13738);
nor U14340 (N_14340,N_13559,N_13810);
or U14341 (N_14341,N_13525,N_13631);
nand U14342 (N_14342,N_13518,N_13687);
nand U14343 (N_14343,N_13657,N_13623);
xor U14344 (N_14344,N_13983,N_13652);
and U14345 (N_14345,N_13731,N_13877);
and U14346 (N_14346,N_13673,N_13945);
nand U14347 (N_14347,N_13984,N_13802);
or U14348 (N_14348,N_13706,N_13745);
xnor U14349 (N_14349,N_13880,N_13733);
and U14350 (N_14350,N_13926,N_13595);
nor U14351 (N_14351,N_13582,N_13689);
or U14352 (N_14352,N_13659,N_13710);
or U14353 (N_14353,N_13756,N_13801);
xnor U14354 (N_14354,N_13797,N_13989);
nor U14355 (N_14355,N_13753,N_13558);
or U14356 (N_14356,N_13935,N_13886);
nor U14357 (N_14357,N_13679,N_13748);
and U14358 (N_14358,N_13706,N_13883);
and U14359 (N_14359,N_13649,N_13696);
nand U14360 (N_14360,N_13891,N_13863);
nor U14361 (N_14361,N_13615,N_13698);
nand U14362 (N_14362,N_13826,N_13594);
nand U14363 (N_14363,N_13535,N_13598);
nand U14364 (N_14364,N_13854,N_13538);
or U14365 (N_14365,N_13786,N_13547);
nand U14366 (N_14366,N_13795,N_13543);
and U14367 (N_14367,N_13766,N_13923);
or U14368 (N_14368,N_13997,N_13893);
and U14369 (N_14369,N_13522,N_13799);
nor U14370 (N_14370,N_13901,N_13795);
nand U14371 (N_14371,N_13848,N_13613);
nand U14372 (N_14372,N_13576,N_13835);
or U14373 (N_14373,N_13987,N_13974);
nor U14374 (N_14374,N_13669,N_13793);
or U14375 (N_14375,N_13564,N_13929);
and U14376 (N_14376,N_13900,N_13705);
xnor U14377 (N_14377,N_13885,N_13672);
xnor U14378 (N_14378,N_13564,N_13995);
xor U14379 (N_14379,N_13916,N_13659);
or U14380 (N_14380,N_13618,N_13745);
and U14381 (N_14381,N_13717,N_13752);
nand U14382 (N_14382,N_13721,N_13889);
and U14383 (N_14383,N_13658,N_13970);
nor U14384 (N_14384,N_13823,N_13983);
xor U14385 (N_14385,N_13682,N_13643);
nand U14386 (N_14386,N_13892,N_13729);
or U14387 (N_14387,N_13536,N_13764);
nor U14388 (N_14388,N_13733,N_13947);
nand U14389 (N_14389,N_13501,N_13720);
nand U14390 (N_14390,N_13622,N_13964);
nor U14391 (N_14391,N_13594,N_13993);
or U14392 (N_14392,N_13898,N_13585);
and U14393 (N_14393,N_13836,N_13712);
or U14394 (N_14394,N_13581,N_13595);
nor U14395 (N_14395,N_13900,N_13653);
nand U14396 (N_14396,N_13640,N_13996);
xor U14397 (N_14397,N_13516,N_13739);
nor U14398 (N_14398,N_13830,N_13670);
or U14399 (N_14399,N_13523,N_13647);
nand U14400 (N_14400,N_13510,N_13982);
and U14401 (N_14401,N_13700,N_13747);
nand U14402 (N_14402,N_13824,N_13948);
nor U14403 (N_14403,N_13503,N_13776);
or U14404 (N_14404,N_13832,N_13776);
and U14405 (N_14405,N_13930,N_13791);
and U14406 (N_14406,N_13620,N_13887);
and U14407 (N_14407,N_13738,N_13807);
or U14408 (N_14408,N_13672,N_13968);
xor U14409 (N_14409,N_13699,N_13767);
nand U14410 (N_14410,N_13603,N_13566);
nor U14411 (N_14411,N_13878,N_13620);
nor U14412 (N_14412,N_13881,N_13988);
or U14413 (N_14413,N_13560,N_13538);
or U14414 (N_14414,N_13590,N_13558);
xnor U14415 (N_14415,N_13774,N_13675);
and U14416 (N_14416,N_13671,N_13744);
and U14417 (N_14417,N_13607,N_13852);
nor U14418 (N_14418,N_13594,N_13858);
and U14419 (N_14419,N_13796,N_13786);
xnor U14420 (N_14420,N_13909,N_13849);
xnor U14421 (N_14421,N_13860,N_13926);
nand U14422 (N_14422,N_13846,N_13969);
nand U14423 (N_14423,N_13886,N_13635);
and U14424 (N_14424,N_13794,N_13942);
nand U14425 (N_14425,N_13661,N_13739);
nand U14426 (N_14426,N_13560,N_13519);
nand U14427 (N_14427,N_13606,N_13970);
nand U14428 (N_14428,N_13922,N_13682);
nor U14429 (N_14429,N_13657,N_13848);
and U14430 (N_14430,N_13665,N_13541);
nand U14431 (N_14431,N_13730,N_13625);
and U14432 (N_14432,N_13722,N_13691);
nand U14433 (N_14433,N_13979,N_13559);
xor U14434 (N_14434,N_13745,N_13977);
nand U14435 (N_14435,N_13672,N_13992);
and U14436 (N_14436,N_13577,N_13668);
nor U14437 (N_14437,N_13803,N_13510);
xor U14438 (N_14438,N_13577,N_13843);
nor U14439 (N_14439,N_13930,N_13915);
nor U14440 (N_14440,N_13504,N_13511);
nor U14441 (N_14441,N_13576,N_13992);
and U14442 (N_14442,N_13930,N_13514);
nand U14443 (N_14443,N_13855,N_13721);
and U14444 (N_14444,N_13777,N_13770);
and U14445 (N_14445,N_13768,N_13508);
nand U14446 (N_14446,N_13970,N_13785);
nor U14447 (N_14447,N_13874,N_13690);
and U14448 (N_14448,N_13533,N_13948);
and U14449 (N_14449,N_13587,N_13721);
nor U14450 (N_14450,N_13612,N_13875);
and U14451 (N_14451,N_13579,N_13687);
nor U14452 (N_14452,N_13770,N_13997);
or U14453 (N_14453,N_13558,N_13898);
nand U14454 (N_14454,N_13518,N_13542);
nand U14455 (N_14455,N_13784,N_13528);
and U14456 (N_14456,N_13837,N_13881);
or U14457 (N_14457,N_13692,N_13867);
and U14458 (N_14458,N_13906,N_13699);
nand U14459 (N_14459,N_13622,N_13848);
or U14460 (N_14460,N_13993,N_13778);
nor U14461 (N_14461,N_13993,N_13883);
nand U14462 (N_14462,N_13510,N_13518);
and U14463 (N_14463,N_13831,N_13570);
or U14464 (N_14464,N_13839,N_13603);
nand U14465 (N_14465,N_13501,N_13619);
nor U14466 (N_14466,N_13605,N_13521);
xnor U14467 (N_14467,N_13543,N_13906);
nand U14468 (N_14468,N_13761,N_13978);
and U14469 (N_14469,N_13948,N_13958);
or U14470 (N_14470,N_13826,N_13548);
nor U14471 (N_14471,N_13575,N_13992);
nand U14472 (N_14472,N_13582,N_13924);
and U14473 (N_14473,N_13834,N_13652);
xnor U14474 (N_14474,N_13940,N_13990);
or U14475 (N_14475,N_13501,N_13786);
and U14476 (N_14476,N_13576,N_13936);
nor U14477 (N_14477,N_13579,N_13575);
and U14478 (N_14478,N_13939,N_13967);
nor U14479 (N_14479,N_13970,N_13723);
nor U14480 (N_14480,N_13875,N_13666);
nor U14481 (N_14481,N_13830,N_13971);
nand U14482 (N_14482,N_13547,N_13700);
nor U14483 (N_14483,N_13545,N_13777);
and U14484 (N_14484,N_13592,N_13558);
nor U14485 (N_14485,N_13655,N_13501);
nand U14486 (N_14486,N_13661,N_13840);
xor U14487 (N_14487,N_13787,N_13625);
and U14488 (N_14488,N_13672,N_13704);
or U14489 (N_14489,N_13562,N_13936);
and U14490 (N_14490,N_13800,N_13700);
nand U14491 (N_14491,N_13897,N_13618);
and U14492 (N_14492,N_13763,N_13988);
and U14493 (N_14493,N_13589,N_13964);
and U14494 (N_14494,N_13690,N_13612);
nand U14495 (N_14495,N_13762,N_13926);
nor U14496 (N_14496,N_13917,N_13901);
nor U14497 (N_14497,N_13818,N_13758);
nand U14498 (N_14498,N_13870,N_13612);
or U14499 (N_14499,N_13700,N_13519);
and U14500 (N_14500,N_14380,N_14464);
nand U14501 (N_14501,N_14484,N_14303);
or U14502 (N_14502,N_14289,N_14461);
nor U14503 (N_14503,N_14496,N_14131);
xor U14504 (N_14504,N_14450,N_14233);
nand U14505 (N_14505,N_14291,N_14349);
nand U14506 (N_14506,N_14389,N_14049);
and U14507 (N_14507,N_14061,N_14469);
nand U14508 (N_14508,N_14155,N_14135);
or U14509 (N_14509,N_14494,N_14407);
xor U14510 (N_14510,N_14322,N_14101);
nand U14511 (N_14511,N_14035,N_14255);
xor U14512 (N_14512,N_14421,N_14042);
and U14513 (N_14513,N_14180,N_14300);
or U14514 (N_14514,N_14246,N_14331);
or U14515 (N_14515,N_14040,N_14344);
or U14516 (N_14516,N_14495,N_14189);
or U14517 (N_14517,N_14041,N_14236);
nand U14518 (N_14518,N_14091,N_14498);
and U14519 (N_14519,N_14362,N_14038);
nand U14520 (N_14520,N_14002,N_14161);
xnor U14521 (N_14521,N_14266,N_14273);
and U14522 (N_14522,N_14446,N_14005);
nand U14523 (N_14523,N_14259,N_14036);
and U14524 (N_14524,N_14373,N_14125);
xnor U14525 (N_14525,N_14491,N_14309);
or U14526 (N_14526,N_14395,N_14237);
and U14527 (N_14527,N_14126,N_14326);
and U14528 (N_14528,N_14466,N_14102);
and U14529 (N_14529,N_14010,N_14197);
xnor U14530 (N_14530,N_14020,N_14472);
nand U14531 (N_14531,N_14134,N_14011);
nor U14532 (N_14532,N_14258,N_14384);
nor U14533 (N_14533,N_14033,N_14415);
and U14534 (N_14534,N_14245,N_14471);
or U14535 (N_14535,N_14286,N_14453);
and U14536 (N_14536,N_14256,N_14100);
nor U14537 (N_14537,N_14463,N_14084);
xor U14538 (N_14538,N_14071,N_14375);
and U14539 (N_14539,N_14054,N_14398);
xnor U14540 (N_14540,N_14391,N_14442);
nor U14541 (N_14541,N_14120,N_14132);
nand U14542 (N_14542,N_14327,N_14149);
or U14543 (N_14543,N_14347,N_14356);
nor U14544 (N_14544,N_14402,N_14119);
or U14545 (N_14545,N_14108,N_14148);
xor U14546 (N_14546,N_14439,N_14295);
xnor U14547 (N_14547,N_14017,N_14048);
and U14548 (N_14548,N_14357,N_14008);
nand U14549 (N_14549,N_14117,N_14165);
nand U14550 (N_14550,N_14064,N_14441);
nor U14551 (N_14551,N_14488,N_14336);
nand U14552 (N_14552,N_14269,N_14417);
nand U14553 (N_14553,N_14107,N_14271);
xor U14554 (N_14554,N_14051,N_14308);
nand U14555 (N_14555,N_14000,N_14001);
and U14556 (N_14556,N_14090,N_14490);
nor U14557 (N_14557,N_14133,N_14432);
and U14558 (N_14558,N_14306,N_14006);
or U14559 (N_14559,N_14234,N_14350);
nand U14560 (N_14560,N_14078,N_14288);
nor U14561 (N_14561,N_14487,N_14114);
and U14562 (N_14562,N_14328,N_14195);
and U14563 (N_14563,N_14159,N_14473);
xnor U14564 (N_14564,N_14368,N_14199);
xor U14565 (N_14565,N_14096,N_14482);
nor U14566 (N_14566,N_14156,N_14351);
and U14567 (N_14567,N_14379,N_14196);
nand U14568 (N_14568,N_14105,N_14462);
nand U14569 (N_14569,N_14278,N_14445);
nor U14570 (N_14570,N_14136,N_14315);
nor U14571 (N_14571,N_14468,N_14184);
nor U14572 (N_14572,N_14050,N_14211);
nand U14573 (N_14573,N_14039,N_14062);
or U14574 (N_14574,N_14264,N_14212);
and U14575 (N_14575,N_14217,N_14325);
xor U14576 (N_14576,N_14403,N_14055);
xor U14577 (N_14577,N_14283,N_14329);
or U14578 (N_14578,N_14168,N_14143);
nor U14579 (N_14579,N_14014,N_14141);
and U14580 (N_14580,N_14457,N_14279);
or U14581 (N_14581,N_14169,N_14140);
nand U14582 (N_14582,N_14173,N_14378);
and U14583 (N_14583,N_14167,N_14024);
xnor U14584 (N_14584,N_14338,N_14434);
and U14585 (N_14585,N_14323,N_14082);
or U14586 (N_14586,N_14438,N_14047);
xnor U14587 (N_14587,N_14274,N_14037);
xor U14588 (N_14588,N_14376,N_14242);
and U14589 (N_14589,N_14252,N_14076);
or U14590 (N_14590,N_14282,N_14174);
nand U14591 (N_14591,N_14359,N_14254);
or U14592 (N_14592,N_14177,N_14367);
xnor U14593 (N_14593,N_14243,N_14066);
nand U14594 (N_14594,N_14477,N_14383);
nand U14595 (N_14595,N_14146,N_14112);
and U14596 (N_14596,N_14364,N_14247);
or U14597 (N_14597,N_14163,N_14467);
nand U14598 (N_14598,N_14301,N_14238);
nand U14599 (N_14599,N_14154,N_14221);
nand U14600 (N_14600,N_14124,N_14190);
nor U14601 (N_14601,N_14123,N_14345);
or U14602 (N_14602,N_14302,N_14183);
xnor U14603 (N_14603,N_14414,N_14228);
xnor U14604 (N_14604,N_14281,N_14276);
or U14605 (N_14605,N_14192,N_14352);
nor U14606 (N_14606,N_14244,N_14410);
nor U14607 (N_14607,N_14390,N_14436);
nor U14608 (N_14608,N_14485,N_14489);
and U14609 (N_14609,N_14070,N_14202);
or U14610 (N_14610,N_14297,N_14377);
nand U14611 (N_14611,N_14387,N_14111);
nor U14612 (N_14612,N_14486,N_14022);
nand U14613 (N_14613,N_14144,N_14068);
and U14614 (N_14614,N_14092,N_14287);
nand U14615 (N_14615,N_14257,N_14069);
xnor U14616 (N_14616,N_14479,N_14121);
nand U14617 (N_14617,N_14200,N_14455);
and U14618 (N_14618,N_14290,N_14435);
nand U14619 (N_14619,N_14251,N_14009);
xor U14620 (N_14620,N_14162,N_14015);
and U14621 (N_14621,N_14012,N_14103);
nand U14622 (N_14622,N_14366,N_14260);
and U14623 (N_14623,N_14460,N_14201);
xnor U14624 (N_14624,N_14056,N_14388);
or U14625 (N_14625,N_14227,N_14393);
nand U14626 (N_14626,N_14369,N_14430);
nand U14627 (N_14627,N_14294,N_14339);
or U14628 (N_14628,N_14209,N_14128);
and U14629 (N_14629,N_14151,N_14348);
xor U14630 (N_14630,N_14346,N_14044);
nor U14631 (N_14631,N_14353,N_14314);
xor U14632 (N_14632,N_14458,N_14474);
nand U14633 (N_14633,N_14232,N_14019);
nor U14634 (N_14634,N_14229,N_14444);
nor U14635 (N_14635,N_14094,N_14045);
and U14636 (N_14636,N_14299,N_14334);
xor U14637 (N_14637,N_14213,N_14275);
nor U14638 (N_14638,N_14305,N_14240);
nor U14639 (N_14639,N_14077,N_14492);
nand U14640 (N_14640,N_14371,N_14493);
nor U14641 (N_14641,N_14138,N_14317);
and U14642 (N_14642,N_14267,N_14116);
nor U14643 (N_14643,N_14052,N_14072);
or U14644 (N_14644,N_14265,N_14231);
or U14645 (N_14645,N_14465,N_14158);
nor U14646 (N_14646,N_14418,N_14164);
nand U14647 (N_14647,N_14433,N_14272);
xor U14648 (N_14648,N_14110,N_14263);
or U14649 (N_14649,N_14063,N_14425);
nor U14650 (N_14650,N_14324,N_14422);
and U14651 (N_14651,N_14130,N_14179);
or U14652 (N_14652,N_14059,N_14447);
xnor U14653 (N_14653,N_14152,N_14067);
nand U14654 (N_14654,N_14075,N_14476);
or U14655 (N_14655,N_14320,N_14007);
xor U14656 (N_14656,N_14404,N_14060);
nand U14657 (N_14657,N_14385,N_14337);
or U14658 (N_14658,N_14304,N_14193);
nand U14659 (N_14659,N_14394,N_14034);
or U14660 (N_14660,N_14046,N_14225);
nor U14661 (N_14661,N_14206,N_14186);
nand U14662 (N_14662,N_14113,N_14449);
xor U14663 (N_14663,N_14437,N_14181);
or U14664 (N_14664,N_14409,N_14032);
nor U14665 (N_14665,N_14443,N_14408);
or U14666 (N_14666,N_14451,N_14157);
and U14667 (N_14667,N_14426,N_14166);
or U14668 (N_14668,N_14270,N_14400);
and U14669 (N_14669,N_14420,N_14086);
or U14670 (N_14670,N_14145,N_14480);
xor U14671 (N_14671,N_14249,N_14153);
xnor U14672 (N_14672,N_14292,N_14427);
and U14673 (N_14673,N_14440,N_14030);
nand U14674 (N_14674,N_14080,N_14215);
xnor U14675 (N_14675,N_14087,N_14003);
or U14676 (N_14676,N_14023,N_14031);
or U14677 (N_14677,N_14239,N_14083);
nand U14678 (N_14678,N_14318,N_14285);
or U14679 (N_14679,N_14313,N_14419);
and U14680 (N_14680,N_14248,N_14284);
nor U14681 (N_14681,N_14218,N_14191);
nor U14682 (N_14682,N_14170,N_14029);
or U14683 (N_14683,N_14321,N_14330);
xnor U14684 (N_14684,N_14065,N_14483);
nand U14685 (N_14685,N_14198,N_14456);
nand U14686 (N_14686,N_14098,N_14185);
or U14687 (N_14687,N_14203,N_14470);
nor U14688 (N_14688,N_14093,N_14250);
nand U14689 (N_14689,N_14210,N_14027);
nand U14690 (N_14690,N_14497,N_14382);
nor U14691 (N_14691,N_14413,N_14214);
nor U14692 (N_14692,N_14099,N_14332);
xor U14693 (N_14693,N_14187,N_14109);
nand U14694 (N_14694,N_14095,N_14171);
nor U14695 (N_14695,N_14293,N_14431);
or U14696 (N_14696,N_14175,N_14230);
or U14697 (N_14697,N_14406,N_14341);
nor U14698 (N_14698,N_14396,N_14454);
or U14699 (N_14699,N_14147,N_14088);
xnor U14700 (N_14700,N_14261,N_14310);
xnor U14701 (N_14701,N_14205,N_14115);
nor U14702 (N_14702,N_14223,N_14397);
or U14703 (N_14703,N_14089,N_14381);
or U14704 (N_14704,N_14208,N_14172);
or U14705 (N_14705,N_14277,N_14365);
xor U14706 (N_14706,N_14013,N_14429);
and U14707 (N_14707,N_14182,N_14004);
xnor U14708 (N_14708,N_14386,N_14150);
xor U14709 (N_14709,N_14204,N_14399);
nand U14710 (N_14710,N_14081,N_14311);
and U14711 (N_14711,N_14316,N_14424);
nor U14712 (N_14712,N_14342,N_14073);
xnor U14713 (N_14713,N_14057,N_14220);
nor U14714 (N_14714,N_14475,N_14262);
nand U14715 (N_14715,N_14481,N_14363);
nor U14716 (N_14716,N_14127,N_14188);
nand U14717 (N_14717,N_14333,N_14355);
xor U14718 (N_14718,N_14374,N_14224);
or U14719 (N_14719,N_14142,N_14452);
xnor U14720 (N_14720,N_14176,N_14085);
nand U14721 (N_14721,N_14226,N_14058);
or U14722 (N_14722,N_14222,N_14448);
nor U14723 (N_14723,N_14354,N_14296);
nand U14724 (N_14724,N_14358,N_14499);
or U14725 (N_14725,N_14343,N_14104);
or U14726 (N_14726,N_14139,N_14459);
nor U14727 (N_14727,N_14392,N_14416);
nor U14728 (N_14728,N_14028,N_14241);
nand U14729 (N_14729,N_14219,N_14079);
or U14730 (N_14730,N_14307,N_14025);
and U14731 (N_14731,N_14340,N_14160);
and U14732 (N_14732,N_14043,N_14312);
nor U14733 (N_14733,N_14360,N_14016);
xnor U14734 (N_14734,N_14053,N_14097);
nand U14735 (N_14735,N_14370,N_14106);
xnor U14736 (N_14736,N_14372,N_14361);
and U14737 (N_14737,N_14118,N_14412);
nand U14738 (N_14738,N_14018,N_14280);
nor U14739 (N_14739,N_14268,N_14405);
xnor U14740 (N_14740,N_14319,N_14253);
xnor U14741 (N_14741,N_14216,N_14401);
xnor U14742 (N_14742,N_14207,N_14235);
and U14743 (N_14743,N_14428,N_14423);
xor U14744 (N_14744,N_14026,N_14021);
and U14745 (N_14745,N_14137,N_14178);
nand U14746 (N_14746,N_14335,N_14478);
nand U14747 (N_14747,N_14194,N_14298);
or U14748 (N_14748,N_14129,N_14074);
or U14749 (N_14749,N_14122,N_14411);
nand U14750 (N_14750,N_14057,N_14047);
nor U14751 (N_14751,N_14240,N_14252);
and U14752 (N_14752,N_14077,N_14173);
nand U14753 (N_14753,N_14151,N_14426);
xnor U14754 (N_14754,N_14381,N_14284);
nor U14755 (N_14755,N_14482,N_14248);
xnor U14756 (N_14756,N_14050,N_14239);
nor U14757 (N_14757,N_14113,N_14144);
nand U14758 (N_14758,N_14015,N_14402);
nor U14759 (N_14759,N_14300,N_14129);
nand U14760 (N_14760,N_14289,N_14070);
nand U14761 (N_14761,N_14442,N_14254);
and U14762 (N_14762,N_14226,N_14001);
xnor U14763 (N_14763,N_14153,N_14103);
nand U14764 (N_14764,N_14241,N_14443);
xnor U14765 (N_14765,N_14246,N_14469);
nand U14766 (N_14766,N_14481,N_14234);
nor U14767 (N_14767,N_14017,N_14135);
or U14768 (N_14768,N_14129,N_14470);
xor U14769 (N_14769,N_14052,N_14068);
and U14770 (N_14770,N_14195,N_14139);
and U14771 (N_14771,N_14167,N_14303);
or U14772 (N_14772,N_14294,N_14095);
or U14773 (N_14773,N_14233,N_14184);
nor U14774 (N_14774,N_14251,N_14257);
nor U14775 (N_14775,N_14345,N_14060);
nand U14776 (N_14776,N_14232,N_14183);
or U14777 (N_14777,N_14390,N_14463);
nor U14778 (N_14778,N_14478,N_14211);
and U14779 (N_14779,N_14045,N_14386);
nand U14780 (N_14780,N_14490,N_14268);
or U14781 (N_14781,N_14293,N_14396);
xnor U14782 (N_14782,N_14334,N_14232);
and U14783 (N_14783,N_14282,N_14063);
and U14784 (N_14784,N_14109,N_14384);
xnor U14785 (N_14785,N_14117,N_14471);
nand U14786 (N_14786,N_14308,N_14441);
xor U14787 (N_14787,N_14003,N_14067);
or U14788 (N_14788,N_14499,N_14350);
and U14789 (N_14789,N_14080,N_14439);
nand U14790 (N_14790,N_14141,N_14443);
nor U14791 (N_14791,N_14051,N_14017);
and U14792 (N_14792,N_14433,N_14192);
xor U14793 (N_14793,N_14307,N_14473);
xor U14794 (N_14794,N_14450,N_14396);
nor U14795 (N_14795,N_14318,N_14360);
nand U14796 (N_14796,N_14078,N_14206);
and U14797 (N_14797,N_14177,N_14494);
xor U14798 (N_14798,N_14044,N_14185);
xnor U14799 (N_14799,N_14455,N_14035);
nor U14800 (N_14800,N_14385,N_14327);
xnor U14801 (N_14801,N_14271,N_14149);
or U14802 (N_14802,N_14319,N_14468);
nor U14803 (N_14803,N_14099,N_14354);
nor U14804 (N_14804,N_14255,N_14265);
and U14805 (N_14805,N_14423,N_14316);
xor U14806 (N_14806,N_14285,N_14236);
xnor U14807 (N_14807,N_14488,N_14159);
nor U14808 (N_14808,N_14428,N_14030);
xor U14809 (N_14809,N_14250,N_14089);
and U14810 (N_14810,N_14270,N_14494);
and U14811 (N_14811,N_14178,N_14328);
nor U14812 (N_14812,N_14003,N_14194);
or U14813 (N_14813,N_14328,N_14228);
xor U14814 (N_14814,N_14019,N_14063);
xor U14815 (N_14815,N_14155,N_14460);
and U14816 (N_14816,N_14292,N_14450);
xor U14817 (N_14817,N_14310,N_14185);
or U14818 (N_14818,N_14109,N_14330);
nand U14819 (N_14819,N_14081,N_14477);
xnor U14820 (N_14820,N_14343,N_14166);
xor U14821 (N_14821,N_14069,N_14272);
or U14822 (N_14822,N_14427,N_14477);
or U14823 (N_14823,N_14475,N_14220);
nor U14824 (N_14824,N_14373,N_14274);
nand U14825 (N_14825,N_14013,N_14153);
nand U14826 (N_14826,N_14122,N_14394);
nor U14827 (N_14827,N_14325,N_14410);
and U14828 (N_14828,N_14468,N_14175);
and U14829 (N_14829,N_14173,N_14354);
nand U14830 (N_14830,N_14085,N_14082);
nor U14831 (N_14831,N_14413,N_14252);
nor U14832 (N_14832,N_14361,N_14428);
nand U14833 (N_14833,N_14245,N_14479);
or U14834 (N_14834,N_14105,N_14355);
nand U14835 (N_14835,N_14012,N_14272);
xor U14836 (N_14836,N_14248,N_14457);
nor U14837 (N_14837,N_14256,N_14060);
xnor U14838 (N_14838,N_14186,N_14012);
or U14839 (N_14839,N_14048,N_14021);
xor U14840 (N_14840,N_14474,N_14409);
nand U14841 (N_14841,N_14483,N_14302);
or U14842 (N_14842,N_14208,N_14071);
or U14843 (N_14843,N_14300,N_14450);
xor U14844 (N_14844,N_14050,N_14285);
and U14845 (N_14845,N_14372,N_14456);
and U14846 (N_14846,N_14298,N_14457);
xnor U14847 (N_14847,N_14020,N_14128);
nand U14848 (N_14848,N_14179,N_14474);
nor U14849 (N_14849,N_14413,N_14491);
and U14850 (N_14850,N_14419,N_14394);
nor U14851 (N_14851,N_14304,N_14063);
or U14852 (N_14852,N_14314,N_14441);
xor U14853 (N_14853,N_14354,N_14035);
or U14854 (N_14854,N_14290,N_14166);
nor U14855 (N_14855,N_14003,N_14453);
and U14856 (N_14856,N_14212,N_14363);
and U14857 (N_14857,N_14059,N_14099);
and U14858 (N_14858,N_14459,N_14269);
or U14859 (N_14859,N_14128,N_14088);
or U14860 (N_14860,N_14388,N_14485);
or U14861 (N_14861,N_14403,N_14070);
nor U14862 (N_14862,N_14435,N_14384);
xor U14863 (N_14863,N_14342,N_14066);
xor U14864 (N_14864,N_14110,N_14396);
and U14865 (N_14865,N_14325,N_14130);
or U14866 (N_14866,N_14201,N_14328);
and U14867 (N_14867,N_14383,N_14020);
nand U14868 (N_14868,N_14022,N_14435);
xnor U14869 (N_14869,N_14395,N_14281);
nor U14870 (N_14870,N_14413,N_14052);
xnor U14871 (N_14871,N_14085,N_14348);
xor U14872 (N_14872,N_14027,N_14388);
nor U14873 (N_14873,N_14058,N_14212);
and U14874 (N_14874,N_14452,N_14092);
and U14875 (N_14875,N_14381,N_14364);
and U14876 (N_14876,N_14146,N_14339);
nor U14877 (N_14877,N_14101,N_14430);
or U14878 (N_14878,N_14130,N_14157);
or U14879 (N_14879,N_14409,N_14451);
xor U14880 (N_14880,N_14356,N_14377);
nor U14881 (N_14881,N_14333,N_14210);
nand U14882 (N_14882,N_14154,N_14051);
nor U14883 (N_14883,N_14211,N_14070);
and U14884 (N_14884,N_14395,N_14426);
nand U14885 (N_14885,N_14102,N_14110);
nand U14886 (N_14886,N_14411,N_14360);
nor U14887 (N_14887,N_14184,N_14264);
and U14888 (N_14888,N_14256,N_14079);
or U14889 (N_14889,N_14292,N_14254);
xnor U14890 (N_14890,N_14463,N_14105);
or U14891 (N_14891,N_14350,N_14262);
nand U14892 (N_14892,N_14282,N_14096);
nand U14893 (N_14893,N_14037,N_14396);
nor U14894 (N_14894,N_14317,N_14047);
and U14895 (N_14895,N_14268,N_14180);
and U14896 (N_14896,N_14497,N_14099);
xnor U14897 (N_14897,N_14344,N_14115);
xnor U14898 (N_14898,N_14088,N_14430);
nand U14899 (N_14899,N_14264,N_14481);
nor U14900 (N_14900,N_14414,N_14116);
nor U14901 (N_14901,N_14312,N_14060);
nor U14902 (N_14902,N_14141,N_14155);
or U14903 (N_14903,N_14277,N_14001);
and U14904 (N_14904,N_14461,N_14469);
and U14905 (N_14905,N_14347,N_14146);
and U14906 (N_14906,N_14350,N_14184);
and U14907 (N_14907,N_14437,N_14213);
and U14908 (N_14908,N_14156,N_14056);
xnor U14909 (N_14909,N_14459,N_14152);
nor U14910 (N_14910,N_14375,N_14003);
nor U14911 (N_14911,N_14224,N_14341);
or U14912 (N_14912,N_14430,N_14024);
and U14913 (N_14913,N_14333,N_14278);
or U14914 (N_14914,N_14447,N_14261);
and U14915 (N_14915,N_14309,N_14297);
or U14916 (N_14916,N_14417,N_14467);
nor U14917 (N_14917,N_14080,N_14109);
nor U14918 (N_14918,N_14147,N_14384);
or U14919 (N_14919,N_14358,N_14218);
nand U14920 (N_14920,N_14156,N_14053);
and U14921 (N_14921,N_14242,N_14399);
or U14922 (N_14922,N_14075,N_14152);
or U14923 (N_14923,N_14431,N_14240);
and U14924 (N_14924,N_14128,N_14113);
xnor U14925 (N_14925,N_14255,N_14135);
and U14926 (N_14926,N_14119,N_14071);
nand U14927 (N_14927,N_14053,N_14135);
xor U14928 (N_14928,N_14272,N_14244);
xor U14929 (N_14929,N_14247,N_14310);
xnor U14930 (N_14930,N_14450,N_14073);
or U14931 (N_14931,N_14203,N_14430);
and U14932 (N_14932,N_14363,N_14010);
nor U14933 (N_14933,N_14020,N_14078);
nand U14934 (N_14934,N_14458,N_14472);
xnor U14935 (N_14935,N_14365,N_14160);
nand U14936 (N_14936,N_14290,N_14206);
nand U14937 (N_14937,N_14160,N_14351);
nor U14938 (N_14938,N_14007,N_14370);
and U14939 (N_14939,N_14170,N_14483);
xor U14940 (N_14940,N_14357,N_14086);
or U14941 (N_14941,N_14147,N_14190);
nor U14942 (N_14942,N_14406,N_14276);
nand U14943 (N_14943,N_14120,N_14363);
nand U14944 (N_14944,N_14119,N_14494);
xnor U14945 (N_14945,N_14174,N_14002);
nand U14946 (N_14946,N_14396,N_14279);
or U14947 (N_14947,N_14420,N_14396);
xor U14948 (N_14948,N_14464,N_14168);
and U14949 (N_14949,N_14452,N_14289);
nor U14950 (N_14950,N_14015,N_14360);
or U14951 (N_14951,N_14493,N_14291);
and U14952 (N_14952,N_14159,N_14495);
xnor U14953 (N_14953,N_14043,N_14381);
or U14954 (N_14954,N_14004,N_14300);
nor U14955 (N_14955,N_14122,N_14416);
and U14956 (N_14956,N_14034,N_14038);
nor U14957 (N_14957,N_14058,N_14064);
nor U14958 (N_14958,N_14385,N_14051);
and U14959 (N_14959,N_14042,N_14147);
nand U14960 (N_14960,N_14412,N_14164);
nand U14961 (N_14961,N_14067,N_14425);
nand U14962 (N_14962,N_14032,N_14051);
or U14963 (N_14963,N_14130,N_14245);
nor U14964 (N_14964,N_14484,N_14020);
and U14965 (N_14965,N_14270,N_14484);
nor U14966 (N_14966,N_14465,N_14194);
or U14967 (N_14967,N_14197,N_14376);
nand U14968 (N_14968,N_14461,N_14312);
xor U14969 (N_14969,N_14456,N_14420);
nor U14970 (N_14970,N_14139,N_14033);
and U14971 (N_14971,N_14020,N_14001);
xnor U14972 (N_14972,N_14200,N_14137);
or U14973 (N_14973,N_14475,N_14032);
nor U14974 (N_14974,N_14395,N_14384);
or U14975 (N_14975,N_14304,N_14484);
or U14976 (N_14976,N_14449,N_14068);
or U14977 (N_14977,N_14281,N_14368);
xor U14978 (N_14978,N_14011,N_14463);
and U14979 (N_14979,N_14049,N_14091);
nor U14980 (N_14980,N_14281,N_14471);
nand U14981 (N_14981,N_14027,N_14420);
xnor U14982 (N_14982,N_14169,N_14162);
xor U14983 (N_14983,N_14181,N_14049);
and U14984 (N_14984,N_14094,N_14281);
xor U14985 (N_14985,N_14155,N_14238);
nor U14986 (N_14986,N_14407,N_14325);
nor U14987 (N_14987,N_14219,N_14242);
and U14988 (N_14988,N_14179,N_14204);
nor U14989 (N_14989,N_14235,N_14302);
or U14990 (N_14990,N_14298,N_14039);
nor U14991 (N_14991,N_14035,N_14347);
nor U14992 (N_14992,N_14205,N_14119);
and U14993 (N_14993,N_14461,N_14194);
nor U14994 (N_14994,N_14412,N_14162);
nor U14995 (N_14995,N_14478,N_14016);
or U14996 (N_14996,N_14303,N_14316);
nor U14997 (N_14997,N_14182,N_14268);
nor U14998 (N_14998,N_14224,N_14179);
xor U14999 (N_14999,N_14323,N_14474);
nand U15000 (N_15000,N_14867,N_14741);
or U15001 (N_15001,N_14813,N_14619);
and U15002 (N_15002,N_14983,N_14666);
and U15003 (N_15003,N_14963,N_14912);
xnor U15004 (N_15004,N_14579,N_14926);
nor U15005 (N_15005,N_14976,N_14773);
xor U15006 (N_15006,N_14540,N_14986);
xnor U15007 (N_15007,N_14947,N_14736);
or U15008 (N_15008,N_14626,N_14653);
or U15009 (N_15009,N_14878,N_14995);
nand U15010 (N_15010,N_14975,N_14921);
or U15011 (N_15011,N_14643,N_14980);
xnor U15012 (N_15012,N_14636,N_14907);
and U15013 (N_15013,N_14827,N_14633);
xor U15014 (N_15014,N_14823,N_14507);
nor U15015 (N_15015,N_14782,N_14593);
xor U15016 (N_15016,N_14638,N_14835);
nand U15017 (N_15017,N_14639,N_14537);
nor U15018 (N_15018,N_14974,N_14502);
nor U15019 (N_15019,N_14992,N_14882);
xor U15020 (N_15020,N_14886,N_14599);
and U15021 (N_15021,N_14716,N_14923);
nor U15022 (N_15022,N_14575,N_14645);
and U15023 (N_15023,N_14706,N_14874);
xnor U15024 (N_15024,N_14936,N_14777);
xor U15025 (N_15025,N_14800,N_14763);
xor U15026 (N_15026,N_14808,N_14945);
nand U15027 (N_15027,N_14534,N_14602);
or U15028 (N_15028,N_14756,N_14739);
xnor U15029 (N_15029,N_14804,N_14817);
nand U15030 (N_15030,N_14862,N_14560);
xor U15031 (N_15031,N_14541,N_14860);
nand U15032 (N_15032,N_14851,N_14880);
and U15033 (N_15033,N_14972,N_14863);
xor U15034 (N_15034,N_14637,N_14696);
nand U15035 (N_15035,N_14610,N_14853);
nand U15036 (N_15036,N_14762,N_14686);
and U15037 (N_15037,N_14994,N_14546);
and U15038 (N_15038,N_14999,N_14829);
or U15039 (N_15039,N_14572,N_14725);
and U15040 (N_15040,N_14962,N_14893);
nor U15041 (N_15041,N_14641,N_14977);
and U15042 (N_15042,N_14832,N_14953);
nor U15043 (N_15043,N_14908,N_14791);
nor U15044 (N_15044,N_14803,N_14771);
and U15045 (N_15045,N_14590,N_14911);
xnor U15046 (N_15046,N_14877,N_14951);
nand U15047 (N_15047,N_14738,N_14997);
xor U15048 (N_15048,N_14830,N_14865);
or U15049 (N_15049,N_14868,N_14818);
nor U15050 (N_15050,N_14535,N_14634);
xnor U15051 (N_15051,N_14723,N_14793);
nor U15052 (N_15052,N_14646,N_14583);
nor U15053 (N_15053,N_14917,N_14663);
xnor U15054 (N_15054,N_14855,N_14720);
xnor U15055 (N_15055,N_14678,N_14734);
and U15056 (N_15056,N_14523,N_14526);
nor U15057 (N_15057,N_14846,N_14884);
xnor U15058 (N_15058,N_14631,N_14891);
and U15059 (N_15059,N_14551,N_14859);
and U15060 (N_15060,N_14801,N_14938);
and U15061 (N_15061,N_14973,N_14718);
xor U15062 (N_15062,N_14611,N_14858);
and U15063 (N_15063,N_14730,N_14752);
nor U15064 (N_15064,N_14520,N_14881);
nand U15065 (N_15065,N_14747,N_14927);
or U15066 (N_15066,N_14650,N_14950);
nor U15067 (N_15067,N_14757,N_14900);
or U15068 (N_15068,N_14514,N_14841);
or U15069 (N_15069,N_14697,N_14679);
xnor U15070 (N_15070,N_14895,N_14627);
nand U15071 (N_15071,N_14866,N_14814);
nand U15072 (N_15072,N_14667,N_14872);
and U15073 (N_15073,N_14568,N_14573);
nand U15074 (N_15074,N_14635,N_14576);
nor U15075 (N_15075,N_14613,N_14525);
nor U15076 (N_15076,N_14515,N_14993);
and U15077 (N_15077,N_14543,N_14929);
nor U15078 (N_15078,N_14713,N_14766);
xor U15079 (N_15079,N_14620,N_14733);
nor U15080 (N_15080,N_14839,N_14510);
nand U15081 (N_15081,N_14794,N_14618);
nor U15082 (N_15082,N_14664,N_14849);
and U15083 (N_15083,N_14699,N_14532);
nand U15084 (N_15084,N_14584,N_14815);
nand U15085 (N_15085,N_14609,N_14796);
nand U15086 (N_15086,N_14749,N_14533);
and U15087 (N_15087,N_14624,N_14674);
nand U15088 (N_15088,N_14854,N_14847);
or U15089 (N_15089,N_14675,N_14587);
nand U15090 (N_15090,N_14565,N_14961);
xor U15091 (N_15091,N_14876,N_14754);
nor U15092 (N_15092,N_14591,N_14668);
or U15093 (N_15093,N_14970,N_14614);
xor U15094 (N_15094,N_14828,N_14988);
nor U15095 (N_15095,N_14850,N_14758);
xnor U15096 (N_15096,N_14967,N_14948);
nor U15097 (N_15097,N_14659,N_14728);
xnor U15098 (N_15098,N_14955,N_14776);
nor U15099 (N_15099,N_14952,N_14647);
nand U15100 (N_15100,N_14968,N_14623);
xnor U15101 (N_15101,N_14842,N_14531);
nor U15102 (N_15102,N_14949,N_14563);
or U15103 (N_15103,N_14562,N_14712);
or U15104 (N_15104,N_14982,N_14632);
or U15105 (N_15105,N_14856,N_14831);
nand U15106 (N_15106,N_14744,N_14608);
xnor U15107 (N_15107,N_14934,N_14745);
nand U15108 (N_15108,N_14629,N_14597);
xor U15109 (N_15109,N_14998,N_14964);
xor U15110 (N_15110,N_14769,N_14790);
xor U15111 (N_15111,N_14630,N_14665);
nor U15112 (N_15112,N_14922,N_14670);
and U15113 (N_15113,N_14621,N_14505);
or U15114 (N_15114,N_14985,N_14698);
nor U15115 (N_15115,N_14598,N_14705);
and U15116 (N_15116,N_14930,N_14774);
nand U15117 (N_15117,N_14661,N_14506);
and U15118 (N_15118,N_14658,N_14802);
nor U15119 (N_15119,N_14707,N_14864);
nor U15120 (N_15120,N_14662,N_14656);
nor U15121 (N_15121,N_14795,N_14913);
xor U15122 (N_15122,N_14750,N_14941);
xnor U15123 (N_15123,N_14906,N_14848);
and U15124 (N_15124,N_14596,N_14996);
nor U15125 (N_15125,N_14935,N_14969);
or U15126 (N_15126,N_14806,N_14990);
nor U15127 (N_15127,N_14991,N_14581);
nor U15128 (N_15128,N_14552,N_14574);
and U15129 (N_15129,N_14722,N_14909);
nand U15130 (N_15130,N_14924,N_14810);
or U15131 (N_15131,N_14742,N_14612);
nor U15132 (N_15132,N_14558,N_14887);
nor U15133 (N_15133,N_14740,N_14530);
nand U15134 (N_15134,N_14873,N_14772);
and U15135 (N_15135,N_14737,N_14617);
or U15136 (N_15136,N_14688,N_14861);
xor U15137 (N_15137,N_14654,N_14657);
xor U15138 (N_15138,N_14694,N_14899);
nor U15139 (N_15139,N_14710,N_14651);
nand U15140 (N_15140,N_14845,N_14640);
and U15141 (N_15141,N_14799,N_14735);
nand U15142 (N_15142,N_14932,N_14601);
or U15143 (N_15143,N_14622,N_14690);
nand U15144 (N_15144,N_14946,N_14748);
nor U15145 (N_15145,N_14836,N_14511);
nand U15146 (N_15146,N_14751,N_14914);
or U15147 (N_15147,N_14711,N_14902);
and U15148 (N_15148,N_14578,N_14903);
or U15149 (N_15149,N_14984,N_14701);
and U15150 (N_15150,N_14978,N_14605);
nor U15151 (N_15151,N_14673,N_14883);
or U15152 (N_15152,N_14919,N_14504);
xor U15153 (N_15153,N_14959,N_14729);
or U15154 (N_15154,N_14569,N_14592);
and U15155 (N_15155,N_14683,N_14965);
nand U15156 (N_15156,N_14557,N_14943);
and U15157 (N_15157,N_14539,N_14896);
nand U15158 (N_15158,N_14732,N_14682);
nor U15159 (N_15159,N_14731,N_14628);
nand U15160 (N_15160,N_14580,N_14979);
and U15161 (N_15161,N_14594,N_14759);
nand U15162 (N_15162,N_14564,N_14779);
nand U15163 (N_15163,N_14516,N_14792);
and U15164 (N_15164,N_14844,N_14536);
nor U15165 (N_15165,N_14518,N_14559);
and U15166 (N_15166,N_14840,N_14652);
or U15167 (N_15167,N_14727,N_14809);
nand U15168 (N_15168,N_14513,N_14798);
xnor U15169 (N_15169,N_14826,N_14685);
nand U15170 (N_15170,N_14797,N_14821);
or U15171 (N_15171,N_14781,N_14655);
and U15172 (N_15172,N_14916,N_14700);
nand U15173 (N_15173,N_14784,N_14527);
xor U15174 (N_15174,N_14554,N_14888);
xnor U15175 (N_15175,N_14607,N_14582);
nor U15176 (N_15176,N_14719,N_14671);
nor U15177 (N_15177,N_14825,N_14692);
or U15178 (N_15178,N_14588,N_14501);
nor U15179 (N_15179,N_14521,N_14807);
xnor U15180 (N_15180,N_14918,N_14755);
xor U15181 (N_15181,N_14760,N_14904);
xnor U15182 (N_15182,N_14517,N_14857);
or U15183 (N_15183,N_14561,N_14702);
nand U15184 (N_15184,N_14549,N_14743);
nand U15185 (N_15185,N_14571,N_14957);
or U15186 (N_15186,N_14889,N_14786);
nand U15187 (N_15187,N_14939,N_14894);
nor U15188 (N_15188,N_14689,N_14585);
xnor U15189 (N_15189,N_14508,N_14649);
nand U15190 (N_15190,N_14570,N_14960);
or U15191 (N_15191,N_14567,N_14717);
or U15192 (N_15192,N_14905,N_14761);
xnor U15193 (N_15193,N_14625,N_14788);
nor U15194 (N_15194,N_14871,N_14838);
and U15195 (N_15195,N_14724,N_14765);
or U15196 (N_15196,N_14954,N_14524);
nor U15197 (N_15197,N_14956,N_14684);
and U15198 (N_15198,N_14648,N_14837);
xor U15199 (N_15199,N_14925,N_14833);
and U15200 (N_15200,N_14500,N_14547);
or U15201 (N_15201,N_14542,N_14709);
nand U15202 (N_15202,N_14715,N_14616);
xnor U15203 (N_15203,N_14870,N_14898);
or U15204 (N_15204,N_14901,N_14885);
xor U15205 (N_15205,N_14834,N_14528);
nor U15206 (N_15206,N_14615,N_14595);
nand U15207 (N_15207,N_14681,N_14556);
nand U15208 (N_15208,N_14672,N_14812);
and U15209 (N_15209,N_14604,N_14869);
nor U15210 (N_15210,N_14695,N_14775);
nand U15211 (N_15211,N_14805,N_14764);
nand U15212 (N_15212,N_14726,N_14971);
nand U15213 (N_15213,N_14989,N_14553);
xor U15214 (N_15214,N_14811,N_14503);
nor U15215 (N_15215,N_14677,N_14586);
xor U15216 (N_15216,N_14522,N_14910);
nand U15217 (N_15217,N_14783,N_14897);
or U15218 (N_15218,N_14879,N_14824);
nor U15219 (N_15219,N_14746,N_14987);
and U15220 (N_15220,N_14875,N_14703);
or U15221 (N_15221,N_14933,N_14577);
nand U15222 (N_15222,N_14566,N_14915);
xor U15223 (N_15223,N_14603,N_14669);
and U15224 (N_15224,N_14940,N_14958);
nand U15225 (N_15225,N_14550,N_14937);
or U15226 (N_15226,N_14966,N_14721);
nand U15227 (N_15227,N_14942,N_14822);
and U15228 (N_15228,N_14890,N_14589);
xor U15229 (N_15229,N_14708,N_14714);
xnor U15230 (N_15230,N_14928,N_14944);
nand U15231 (N_15231,N_14509,N_14680);
nor U15232 (N_15232,N_14691,N_14981);
xor U15233 (N_15233,N_14767,N_14660);
nor U15234 (N_15234,N_14642,N_14816);
and U15235 (N_15235,N_14545,N_14787);
nor U15236 (N_15236,N_14780,N_14819);
nand U15237 (N_15237,N_14544,N_14753);
nand U15238 (N_15238,N_14519,N_14555);
and U15239 (N_15239,N_14644,N_14606);
nor U15240 (N_15240,N_14920,N_14538);
xor U15241 (N_15241,N_14600,N_14529);
and U15242 (N_15242,N_14548,N_14789);
or U15243 (N_15243,N_14843,N_14931);
and U15244 (N_15244,N_14676,N_14852);
or U15245 (N_15245,N_14768,N_14820);
and U15246 (N_15246,N_14770,N_14785);
nor U15247 (N_15247,N_14778,N_14687);
nand U15248 (N_15248,N_14704,N_14892);
nor U15249 (N_15249,N_14512,N_14693);
nand U15250 (N_15250,N_14568,N_14947);
xnor U15251 (N_15251,N_14951,N_14706);
xnor U15252 (N_15252,N_14707,N_14914);
or U15253 (N_15253,N_14802,N_14710);
or U15254 (N_15254,N_14945,N_14920);
and U15255 (N_15255,N_14606,N_14970);
and U15256 (N_15256,N_14901,N_14568);
xnor U15257 (N_15257,N_14796,N_14502);
xnor U15258 (N_15258,N_14943,N_14823);
or U15259 (N_15259,N_14882,N_14863);
and U15260 (N_15260,N_14696,N_14663);
nor U15261 (N_15261,N_14982,N_14812);
nand U15262 (N_15262,N_14624,N_14619);
nor U15263 (N_15263,N_14585,N_14635);
xor U15264 (N_15264,N_14669,N_14784);
or U15265 (N_15265,N_14681,N_14670);
nand U15266 (N_15266,N_14785,N_14780);
and U15267 (N_15267,N_14904,N_14711);
nand U15268 (N_15268,N_14781,N_14614);
nor U15269 (N_15269,N_14710,N_14585);
or U15270 (N_15270,N_14556,N_14770);
or U15271 (N_15271,N_14903,N_14735);
and U15272 (N_15272,N_14642,N_14900);
nand U15273 (N_15273,N_14545,N_14531);
nand U15274 (N_15274,N_14905,N_14546);
nor U15275 (N_15275,N_14820,N_14826);
nor U15276 (N_15276,N_14775,N_14591);
nand U15277 (N_15277,N_14780,N_14577);
or U15278 (N_15278,N_14823,N_14996);
nor U15279 (N_15279,N_14597,N_14609);
and U15280 (N_15280,N_14614,N_14947);
or U15281 (N_15281,N_14669,N_14608);
nor U15282 (N_15282,N_14986,N_14756);
or U15283 (N_15283,N_14699,N_14631);
nand U15284 (N_15284,N_14830,N_14791);
and U15285 (N_15285,N_14972,N_14685);
nand U15286 (N_15286,N_14860,N_14639);
nand U15287 (N_15287,N_14863,N_14920);
xnor U15288 (N_15288,N_14884,N_14511);
and U15289 (N_15289,N_14930,N_14685);
and U15290 (N_15290,N_14569,N_14986);
nand U15291 (N_15291,N_14794,N_14934);
and U15292 (N_15292,N_14540,N_14804);
nor U15293 (N_15293,N_14870,N_14885);
or U15294 (N_15294,N_14893,N_14727);
and U15295 (N_15295,N_14672,N_14810);
or U15296 (N_15296,N_14941,N_14928);
and U15297 (N_15297,N_14721,N_14986);
and U15298 (N_15298,N_14756,N_14972);
or U15299 (N_15299,N_14945,N_14840);
and U15300 (N_15300,N_14508,N_14521);
and U15301 (N_15301,N_14697,N_14808);
or U15302 (N_15302,N_14822,N_14533);
nor U15303 (N_15303,N_14553,N_14615);
and U15304 (N_15304,N_14593,N_14841);
or U15305 (N_15305,N_14913,N_14831);
xnor U15306 (N_15306,N_14528,N_14949);
nand U15307 (N_15307,N_14607,N_14519);
nand U15308 (N_15308,N_14934,N_14951);
nand U15309 (N_15309,N_14827,N_14801);
and U15310 (N_15310,N_14787,N_14886);
nor U15311 (N_15311,N_14842,N_14583);
or U15312 (N_15312,N_14512,N_14643);
nor U15313 (N_15313,N_14728,N_14807);
nor U15314 (N_15314,N_14724,N_14538);
and U15315 (N_15315,N_14665,N_14910);
and U15316 (N_15316,N_14583,N_14790);
xor U15317 (N_15317,N_14888,N_14850);
xor U15318 (N_15318,N_14584,N_14634);
xnor U15319 (N_15319,N_14982,N_14980);
nand U15320 (N_15320,N_14665,N_14753);
or U15321 (N_15321,N_14937,N_14851);
xnor U15322 (N_15322,N_14612,N_14961);
or U15323 (N_15323,N_14730,N_14521);
nor U15324 (N_15324,N_14532,N_14990);
xor U15325 (N_15325,N_14687,N_14605);
xor U15326 (N_15326,N_14938,N_14796);
or U15327 (N_15327,N_14590,N_14936);
and U15328 (N_15328,N_14970,N_14518);
nor U15329 (N_15329,N_14602,N_14858);
xor U15330 (N_15330,N_14752,N_14511);
or U15331 (N_15331,N_14691,N_14780);
nor U15332 (N_15332,N_14969,N_14555);
or U15333 (N_15333,N_14842,N_14781);
xor U15334 (N_15334,N_14880,N_14965);
or U15335 (N_15335,N_14982,N_14728);
xor U15336 (N_15336,N_14742,N_14877);
nand U15337 (N_15337,N_14669,N_14731);
and U15338 (N_15338,N_14939,N_14702);
and U15339 (N_15339,N_14592,N_14647);
nor U15340 (N_15340,N_14978,N_14947);
nand U15341 (N_15341,N_14849,N_14502);
xor U15342 (N_15342,N_14706,N_14631);
or U15343 (N_15343,N_14577,N_14641);
xor U15344 (N_15344,N_14849,N_14685);
nor U15345 (N_15345,N_14735,N_14795);
nand U15346 (N_15346,N_14950,N_14982);
or U15347 (N_15347,N_14638,N_14977);
xor U15348 (N_15348,N_14514,N_14944);
nand U15349 (N_15349,N_14647,N_14706);
nor U15350 (N_15350,N_14858,N_14612);
or U15351 (N_15351,N_14927,N_14726);
nor U15352 (N_15352,N_14635,N_14893);
nor U15353 (N_15353,N_14622,N_14548);
xnor U15354 (N_15354,N_14840,N_14705);
xnor U15355 (N_15355,N_14777,N_14859);
or U15356 (N_15356,N_14524,N_14592);
xor U15357 (N_15357,N_14591,N_14981);
or U15358 (N_15358,N_14948,N_14657);
or U15359 (N_15359,N_14866,N_14535);
nor U15360 (N_15360,N_14896,N_14555);
nand U15361 (N_15361,N_14694,N_14838);
or U15362 (N_15362,N_14777,N_14515);
xnor U15363 (N_15363,N_14816,N_14937);
and U15364 (N_15364,N_14989,N_14522);
nand U15365 (N_15365,N_14899,N_14738);
nor U15366 (N_15366,N_14541,N_14836);
nand U15367 (N_15367,N_14796,N_14708);
and U15368 (N_15368,N_14910,N_14602);
nor U15369 (N_15369,N_14601,N_14822);
nand U15370 (N_15370,N_14708,N_14526);
xor U15371 (N_15371,N_14827,N_14680);
nor U15372 (N_15372,N_14669,N_14761);
and U15373 (N_15373,N_14913,N_14651);
xnor U15374 (N_15374,N_14727,N_14604);
xnor U15375 (N_15375,N_14930,N_14520);
nor U15376 (N_15376,N_14594,N_14832);
and U15377 (N_15377,N_14530,N_14506);
xnor U15378 (N_15378,N_14645,N_14886);
nand U15379 (N_15379,N_14634,N_14667);
or U15380 (N_15380,N_14658,N_14992);
and U15381 (N_15381,N_14560,N_14921);
or U15382 (N_15382,N_14746,N_14992);
nand U15383 (N_15383,N_14655,N_14961);
xnor U15384 (N_15384,N_14513,N_14746);
and U15385 (N_15385,N_14927,N_14883);
or U15386 (N_15386,N_14694,N_14866);
and U15387 (N_15387,N_14592,N_14671);
xnor U15388 (N_15388,N_14923,N_14737);
and U15389 (N_15389,N_14595,N_14912);
and U15390 (N_15390,N_14744,N_14625);
nand U15391 (N_15391,N_14863,N_14770);
and U15392 (N_15392,N_14759,N_14613);
and U15393 (N_15393,N_14774,N_14557);
and U15394 (N_15394,N_14500,N_14957);
or U15395 (N_15395,N_14518,N_14756);
nand U15396 (N_15396,N_14721,N_14617);
and U15397 (N_15397,N_14712,N_14853);
nor U15398 (N_15398,N_14833,N_14556);
and U15399 (N_15399,N_14726,N_14514);
xnor U15400 (N_15400,N_14894,N_14574);
or U15401 (N_15401,N_14672,N_14581);
or U15402 (N_15402,N_14850,N_14946);
xor U15403 (N_15403,N_14733,N_14522);
xnor U15404 (N_15404,N_14797,N_14829);
nand U15405 (N_15405,N_14687,N_14712);
nand U15406 (N_15406,N_14893,N_14724);
or U15407 (N_15407,N_14511,N_14914);
nand U15408 (N_15408,N_14606,N_14510);
and U15409 (N_15409,N_14580,N_14806);
xor U15410 (N_15410,N_14967,N_14574);
or U15411 (N_15411,N_14530,N_14712);
nand U15412 (N_15412,N_14909,N_14554);
or U15413 (N_15413,N_14912,N_14949);
nor U15414 (N_15414,N_14804,N_14915);
nor U15415 (N_15415,N_14975,N_14543);
nor U15416 (N_15416,N_14720,N_14732);
and U15417 (N_15417,N_14752,N_14585);
xnor U15418 (N_15418,N_14749,N_14625);
xor U15419 (N_15419,N_14757,N_14926);
xnor U15420 (N_15420,N_14858,N_14904);
and U15421 (N_15421,N_14829,N_14643);
nor U15422 (N_15422,N_14589,N_14619);
nor U15423 (N_15423,N_14950,N_14507);
nor U15424 (N_15424,N_14843,N_14663);
xor U15425 (N_15425,N_14683,N_14809);
or U15426 (N_15426,N_14940,N_14523);
or U15427 (N_15427,N_14661,N_14635);
xor U15428 (N_15428,N_14606,N_14651);
nor U15429 (N_15429,N_14750,N_14694);
nor U15430 (N_15430,N_14701,N_14563);
or U15431 (N_15431,N_14918,N_14658);
nor U15432 (N_15432,N_14633,N_14667);
and U15433 (N_15433,N_14682,N_14661);
or U15434 (N_15434,N_14808,N_14899);
nor U15435 (N_15435,N_14995,N_14538);
or U15436 (N_15436,N_14676,N_14564);
and U15437 (N_15437,N_14822,N_14730);
nand U15438 (N_15438,N_14867,N_14619);
nand U15439 (N_15439,N_14775,N_14885);
nor U15440 (N_15440,N_14602,N_14575);
nor U15441 (N_15441,N_14744,N_14821);
xor U15442 (N_15442,N_14683,N_14974);
or U15443 (N_15443,N_14954,N_14999);
or U15444 (N_15444,N_14597,N_14637);
nand U15445 (N_15445,N_14507,N_14553);
and U15446 (N_15446,N_14618,N_14986);
and U15447 (N_15447,N_14897,N_14676);
or U15448 (N_15448,N_14854,N_14848);
nand U15449 (N_15449,N_14565,N_14578);
nand U15450 (N_15450,N_14989,N_14928);
and U15451 (N_15451,N_14598,N_14755);
and U15452 (N_15452,N_14606,N_14998);
nand U15453 (N_15453,N_14845,N_14904);
and U15454 (N_15454,N_14668,N_14585);
xor U15455 (N_15455,N_14655,N_14942);
or U15456 (N_15456,N_14513,N_14653);
and U15457 (N_15457,N_14777,N_14898);
xnor U15458 (N_15458,N_14557,N_14712);
nor U15459 (N_15459,N_14872,N_14590);
and U15460 (N_15460,N_14901,N_14999);
nand U15461 (N_15461,N_14673,N_14837);
and U15462 (N_15462,N_14676,N_14925);
nor U15463 (N_15463,N_14689,N_14732);
nand U15464 (N_15464,N_14912,N_14539);
nand U15465 (N_15465,N_14753,N_14565);
nor U15466 (N_15466,N_14743,N_14796);
nand U15467 (N_15467,N_14583,N_14573);
or U15468 (N_15468,N_14907,N_14789);
nand U15469 (N_15469,N_14908,N_14884);
nor U15470 (N_15470,N_14811,N_14648);
nand U15471 (N_15471,N_14715,N_14603);
or U15472 (N_15472,N_14673,N_14608);
xnor U15473 (N_15473,N_14748,N_14911);
nor U15474 (N_15474,N_14957,N_14834);
or U15475 (N_15475,N_14506,N_14838);
nand U15476 (N_15476,N_14872,N_14512);
xnor U15477 (N_15477,N_14674,N_14561);
nand U15478 (N_15478,N_14625,N_14709);
xnor U15479 (N_15479,N_14662,N_14949);
nor U15480 (N_15480,N_14747,N_14827);
nand U15481 (N_15481,N_14502,N_14855);
xnor U15482 (N_15482,N_14520,N_14912);
nand U15483 (N_15483,N_14519,N_14636);
nor U15484 (N_15484,N_14638,N_14531);
or U15485 (N_15485,N_14872,N_14789);
nand U15486 (N_15486,N_14628,N_14809);
xor U15487 (N_15487,N_14887,N_14973);
nand U15488 (N_15488,N_14814,N_14835);
and U15489 (N_15489,N_14698,N_14656);
nor U15490 (N_15490,N_14873,N_14679);
and U15491 (N_15491,N_14930,N_14783);
nor U15492 (N_15492,N_14753,N_14561);
nand U15493 (N_15493,N_14664,N_14904);
and U15494 (N_15494,N_14744,N_14597);
nand U15495 (N_15495,N_14820,N_14755);
xor U15496 (N_15496,N_14712,N_14509);
nand U15497 (N_15497,N_14734,N_14871);
nor U15498 (N_15498,N_14929,N_14724);
nand U15499 (N_15499,N_14633,N_14967);
or U15500 (N_15500,N_15462,N_15335);
or U15501 (N_15501,N_15048,N_15470);
or U15502 (N_15502,N_15294,N_15004);
and U15503 (N_15503,N_15028,N_15402);
xor U15504 (N_15504,N_15258,N_15245);
and U15505 (N_15505,N_15367,N_15083);
or U15506 (N_15506,N_15151,N_15366);
nor U15507 (N_15507,N_15092,N_15097);
nor U15508 (N_15508,N_15293,N_15042);
xor U15509 (N_15509,N_15128,N_15044);
nor U15510 (N_15510,N_15168,N_15051);
or U15511 (N_15511,N_15306,N_15389);
nor U15512 (N_15512,N_15291,N_15019);
xor U15513 (N_15513,N_15208,N_15252);
nand U15514 (N_15514,N_15447,N_15164);
xnor U15515 (N_15515,N_15326,N_15103);
nor U15516 (N_15516,N_15463,N_15435);
nand U15517 (N_15517,N_15399,N_15279);
xor U15518 (N_15518,N_15388,N_15322);
nor U15519 (N_15519,N_15095,N_15417);
xnor U15520 (N_15520,N_15041,N_15085);
or U15521 (N_15521,N_15328,N_15045);
nand U15522 (N_15522,N_15337,N_15008);
nand U15523 (N_15523,N_15263,N_15400);
nand U15524 (N_15524,N_15397,N_15458);
nor U15525 (N_15525,N_15407,N_15285);
and U15526 (N_15526,N_15405,N_15016);
or U15527 (N_15527,N_15066,N_15432);
or U15528 (N_15528,N_15251,N_15375);
xor U15529 (N_15529,N_15370,N_15466);
nand U15530 (N_15530,N_15473,N_15010);
and U15531 (N_15531,N_15341,N_15018);
and U15532 (N_15532,N_15060,N_15346);
xor U15533 (N_15533,N_15136,N_15319);
nand U15534 (N_15534,N_15012,N_15132);
and U15535 (N_15535,N_15104,N_15025);
nand U15536 (N_15536,N_15054,N_15234);
or U15537 (N_15537,N_15376,N_15209);
and U15538 (N_15538,N_15394,N_15213);
nand U15539 (N_15539,N_15149,N_15377);
nand U15540 (N_15540,N_15070,N_15476);
and U15541 (N_15541,N_15098,N_15429);
nor U15542 (N_15542,N_15225,N_15372);
nand U15543 (N_15543,N_15365,N_15492);
nand U15544 (N_15544,N_15109,N_15179);
or U15545 (N_15545,N_15090,N_15061);
nor U15546 (N_15546,N_15301,N_15112);
and U15547 (N_15547,N_15193,N_15284);
nand U15548 (N_15548,N_15155,N_15451);
nor U15549 (N_15549,N_15441,N_15310);
xor U15550 (N_15550,N_15250,N_15487);
or U15551 (N_15551,N_15434,N_15224);
xnor U15552 (N_15552,N_15127,N_15262);
nor U15553 (N_15553,N_15498,N_15099);
or U15554 (N_15554,N_15295,N_15409);
and U15555 (N_15555,N_15243,N_15320);
xnor U15556 (N_15556,N_15415,N_15032);
nor U15557 (N_15557,N_15353,N_15232);
nor U15558 (N_15558,N_15390,N_15031);
nor U15559 (N_15559,N_15137,N_15486);
xnor U15560 (N_15560,N_15049,N_15256);
nand U15561 (N_15561,N_15312,N_15069);
or U15562 (N_15562,N_15236,N_15253);
or U15563 (N_15563,N_15167,N_15229);
or U15564 (N_15564,N_15349,N_15246);
nand U15565 (N_15565,N_15182,N_15283);
xor U15566 (N_15566,N_15471,N_15218);
nand U15567 (N_15567,N_15348,N_15043);
and U15568 (N_15568,N_15309,N_15126);
and U15569 (N_15569,N_15361,N_15057);
xor U15570 (N_15570,N_15379,N_15489);
nor U15571 (N_15571,N_15427,N_15276);
nor U15572 (N_15572,N_15459,N_15091);
or U15573 (N_15573,N_15001,N_15238);
nor U15574 (N_15574,N_15383,N_15391);
xnor U15575 (N_15575,N_15134,N_15260);
and U15576 (N_15576,N_15248,N_15161);
nor U15577 (N_15577,N_15403,N_15443);
nor U15578 (N_15578,N_15003,N_15172);
nand U15579 (N_15579,N_15360,N_15106);
or U15580 (N_15580,N_15327,N_15196);
or U15581 (N_15581,N_15211,N_15497);
and U15582 (N_15582,N_15005,N_15411);
nor U15583 (N_15583,N_15053,N_15176);
or U15584 (N_15584,N_15318,N_15189);
or U15585 (N_15585,N_15425,N_15135);
nor U15586 (N_15586,N_15290,N_15449);
nand U15587 (N_15587,N_15040,N_15445);
and U15588 (N_15588,N_15364,N_15261);
or U15589 (N_15589,N_15495,N_15423);
nor U15590 (N_15590,N_15108,N_15114);
and U15591 (N_15591,N_15133,N_15257);
or U15592 (N_15592,N_15185,N_15485);
and U15593 (N_15593,N_15347,N_15442);
and U15594 (N_15594,N_15385,N_15000);
or U15595 (N_15595,N_15204,N_15289);
nor U15596 (N_15596,N_15436,N_15047);
and U15597 (N_15597,N_15152,N_15147);
nor U15598 (N_15598,N_15195,N_15223);
nand U15599 (N_15599,N_15329,N_15359);
xnor U15600 (N_15600,N_15214,N_15052);
nand U15601 (N_15601,N_15007,N_15288);
nand U15602 (N_15602,N_15171,N_15490);
xnor U15603 (N_15603,N_15292,N_15222);
or U15604 (N_15604,N_15418,N_15075);
nor U15605 (N_15605,N_15015,N_15215);
nand U15606 (N_15606,N_15480,N_15159);
nand U15607 (N_15607,N_15446,N_15472);
or U15608 (N_15608,N_15452,N_15267);
nor U15609 (N_15609,N_15094,N_15055);
or U15610 (N_15610,N_15333,N_15268);
xnor U15611 (N_15611,N_15191,N_15068);
nand U15612 (N_15612,N_15358,N_15062);
nand U15613 (N_15613,N_15424,N_15474);
or U15614 (N_15614,N_15249,N_15461);
xnor U15615 (N_15615,N_15079,N_15113);
nand U15616 (N_15616,N_15146,N_15180);
and U15617 (N_15617,N_15100,N_15494);
and U15618 (N_15618,N_15227,N_15324);
or U15619 (N_15619,N_15380,N_15130);
nand U15620 (N_15620,N_15174,N_15111);
nor U15621 (N_15621,N_15426,N_15316);
nor U15622 (N_15622,N_15422,N_15190);
nor U15623 (N_15623,N_15428,N_15404);
or U15624 (N_15624,N_15455,N_15493);
nand U15625 (N_15625,N_15039,N_15050);
xor U15626 (N_15626,N_15482,N_15266);
or U15627 (N_15627,N_15124,N_15207);
xor U15628 (N_15628,N_15082,N_15265);
nand U15629 (N_15629,N_15065,N_15200);
nor U15630 (N_15630,N_15125,N_15080);
nand U15631 (N_15631,N_15163,N_15338);
nand U15632 (N_15632,N_15036,N_15469);
or U15633 (N_15633,N_15431,N_15339);
xor U15634 (N_15634,N_15242,N_15244);
and U15635 (N_15635,N_15302,N_15384);
nand U15636 (N_15636,N_15323,N_15173);
and U15637 (N_15637,N_15101,N_15142);
nand U15638 (N_15638,N_15226,N_15074);
xnor U15639 (N_15639,N_15145,N_15064);
nor U15640 (N_15640,N_15181,N_15027);
xor U15641 (N_15641,N_15084,N_15491);
xor U15642 (N_15642,N_15314,N_15465);
xor U15643 (N_15643,N_15175,N_15107);
or U15644 (N_15644,N_15440,N_15002);
and U15645 (N_15645,N_15307,N_15131);
or U15646 (N_15646,N_15340,N_15378);
or U15647 (N_15647,N_15033,N_15274);
and U15648 (N_15648,N_15475,N_15186);
and U15649 (N_15649,N_15437,N_15479);
or U15650 (N_15650,N_15350,N_15321);
and U15651 (N_15651,N_15264,N_15058);
xnor U15652 (N_15652,N_15371,N_15281);
or U15653 (N_15653,N_15356,N_15138);
or U15654 (N_15654,N_15071,N_15072);
and U15655 (N_15655,N_15140,N_15011);
nor U15656 (N_15656,N_15115,N_15014);
nor U15657 (N_15657,N_15221,N_15331);
xor U15658 (N_15658,N_15240,N_15153);
or U15659 (N_15659,N_15278,N_15230);
xor U15660 (N_15660,N_15121,N_15355);
nand U15661 (N_15661,N_15122,N_15086);
and U15662 (N_15662,N_15296,N_15026);
nor U15663 (N_15663,N_15216,N_15017);
or U15664 (N_15664,N_15160,N_15484);
nor U15665 (N_15665,N_15282,N_15336);
xor U15666 (N_15666,N_15464,N_15165);
nor U15667 (N_15667,N_15387,N_15270);
and U15668 (N_15668,N_15139,N_15219);
and U15669 (N_15669,N_15202,N_15170);
and U15670 (N_15670,N_15363,N_15344);
nand U15671 (N_15671,N_15158,N_15408);
nand U15672 (N_15672,N_15420,N_15343);
nand U15673 (N_15673,N_15352,N_15374);
xnor U15674 (N_15674,N_15067,N_15034);
and U15675 (N_15675,N_15305,N_15406);
nor U15676 (N_15676,N_15119,N_15096);
nand U15677 (N_15677,N_15154,N_15298);
nor U15678 (N_15678,N_15395,N_15228);
nand U15679 (N_15679,N_15414,N_15313);
nand U15680 (N_15680,N_15037,N_15241);
and U15681 (N_15681,N_15259,N_15035);
xnor U15682 (N_15682,N_15203,N_15089);
xnor U15683 (N_15683,N_15330,N_15198);
xnor U15684 (N_15684,N_15239,N_15334);
nor U15685 (N_15685,N_15117,N_15450);
or U15686 (N_15686,N_15141,N_15460);
xnor U15687 (N_15687,N_15396,N_15392);
xnor U15688 (N_15688,N_15477,N_15448);
or U15689 (N_15689,N_15169,N_15499);
xnor U15690 (N_15690,N_15201,N_15233);
or U15691 (N_15691,N_15369,N_15373);
and U15692 (N_15692,N_15304,N_15059);
nor U15693 (N_15693,N_15453,N_15038);
nor U15694 (N_15694,N_15287,N_15188);
and U15695 (N_15695,N_15433,N_15087);
nand U15696 (N_15696,N_15362,N_15217);
nor U15697 (N_15697,N_15046,N_15013);
and U15698 (N_15698,N_15299,N_15156);
and U15699 (N_15699,N_15162,N_15020);
or U15700 (N_15700,N_15212,N_15496);
nand U15701 (N_15701,N_15093,N_15237);
and U15702 (N_15702,N_15247,N_15029);
and U15703 (N_15703,N_15342,N_15430);
nor U15704 (N_15704,N_15177,N_15178);
nor U15705 (N_15705,N_15351,N_15076);
or U15706 (N_15706,N_15467,N_15199);
nor U15707 (N_15707,N_15009,N_15220);
nand U15708 (N_15708,N_15468,N_15192);
nand U15709 (N_15709,N_15118,N_15006);
nand U15710 (N_15710,N_15315,N_15439);
xor U15711 (N_15711,N_15024,N_15308);
or U15712 (N_15712,N_15269,N_15102);
xnor U15713 (N_15713,N_15286,N_15303);
and U15714 (N_15714,N_15271,N_15393);
and U15715 (N_15715,N_15254,N_15078);
xor U15716 (N_15716,N_15325,N_15275);
or U15717 (N_15717,N_15157,N_15022);
nor U15718 (N_15718,N_15235,N_15077);
and U15719 (N_15719,N_15144,N_15401);
nand U15720 (N_15720,N_15277,N_15116);
xor U15721 (N_15721,N_15483,N_15381);
xor U15722 (N_15722,N_15368,N_15166);
nor U15723 (N_15723,N_15297,N_15129);
xnor U15724 (N_15724,N_15311,N_15210);
xnor U15725 (N_15725,N_15021,N_15272);
and U15726 (N_15726,N_15150,N_15063);
xor U15727 (N_15727,N_15481,N_15143);
nand U15728 (N_15728,N_15187,N_15410);
or U15729 (N_15729,N_15184,N_15056);
and U15730 (N_15730,N_15357,N_15317);
and U15731 (N_15731,N_15123,N_15457);
and U15732 (N_15732,N_15345,N_15197);
and U15733 (N_15733,N_15300,N_15194);
or U15734 (N_15734,N_15183,N_15206);
or U15735 (N_15735,N_15354,N_15273);
or U15736 (N_15736,N_15205,N_15456);
or U15737 (N_15737,N_15231,N_15421);
or U15738 (N_15738,N_15332,N_15105);
xor U15739 (N_15739,N_15023,N_15088);
nor U15740 (N_15740,N_15412,N_15382);
and U15741 (N_15741,N_15444,N_15386);
or U15742 (N_15742,N_15255,N_15413);
xnor U15743 (N_15743,N_15030,N_15488);
nor U15744 (N_15744,N_15416,N_15438);
and U15745 (N_15745,N_15280,N_15110);
xnor U15746 (N_15746,N_15120,N_15478);
xnor U15747 (N_15747,N_15398,N_15148);
nor U15748 (N_15748,N_15419,N_15454);
or U15749 (N_15749,N_15081,N_15073);
or U15750 (N_15750,N_15224,N_15303);
nor U15751 (N_15751,N_15330,N_15463);
nor U15752 (N_15752,N_15447,N_15339);
nor U15753 (N_15753,N_15183,N_15392);
and U15754 (N_15754,N_15301,N_15160);
or U15755 (N_15755,N_15222,N_15481);
nor U15756 (N_15756,N_15329,N_15440);
or U15757 (N_15757,N_15318,N_15448);
or U15758 (N_15758,N_15219,N_15073);
xnor U15759 (N_15759,N_15280,N_15044);
nor U15760 (N_15760,N_15132,N_15464);
nor U15761 (N_15761,N_15104,N_15112);
or U15762 (N_15762,N_15085,N_15175);
xor U15763 (N_15763,N_15267,N_15081);
nand U15764 (N_15764,N_15384,N_15182);
and U15765 (N_15765,N_15087,N_15287);
xor U15766 (N_15766,N_15119,N_15395);
and U15767 (N_15767,N_15242,N_15489);
nor U15768 (N_15768,N_15412,N_15231);
or U15769 (N_15769,N_15465,N_15265);
and U15770 (N_15770,N_15293,N_15180);
nor U15771 (N_15771,N_15463,N_15306);
nand U15772 (N_15772,N_15112,N_15054);
or U15773 (N_15773,N_15070,N_15164);
and U15774 (N_15774,N_15435,N_15460);
nand U15775 (N_15775,N_15231,N_15463);
and U15776 (N_15776,N_15430,N_15264);
or U15777 (N_15777,N_15036,N_15306);
nor U15778 (N_15778,N_15156,N_15470);
and U15779 (N_15779,N_15025,N_15278);
xor U15780 (N_15780,N_15361,N_15099);
xnor U15781 (N_15781,N_15002,N_15196);
and U15782 (N_15782,N_15020,N_15211);
nor U15783 (N_15783,N_15280,N_15214);
nor U15784 (N_15784,N_15326,N_15143);
or U15785 (N_15785,N_15152,N_15341);
nand U15786 (N_15786,N_15190,N_15321);
xor U15787 (N_15787,N_15278,N_15015);
nand U15788 (N_15788,N_15497,N_15095);
xor U15789 (N_15789,N_15254,N_15467);
nor U15790 (N_15790,N_15436,N_15018);
nor U15791 (N_15791,N_15287,N_15059);
nor U15792 (N_15792,N_15276,N_15386);
or U15793 (N_15793,N_15394,N_15140);
nand U15794 (N_15794,N_15300,N_15338);
nand U15795 (N_15795,N_15144,N_15223);
or U15796 (N_15796,N_15141,N_15135);
and U15797 (N_15797,N_15276,N_15259);
nand U15798 (N_15798,N_15060,N_15026);
or U15799 (N_15799,N_15308,N_15475);
or U15800 (N_15800,N_15494,N_15021);
xor U15801 (N_15801,N_15163,N_15167);
nor U15802 (N_15802,N_15201,N_15142);
xnor U15803 (N_15803,N_15240,N_15431);
xor U15804 (N_15804,N_15208,N_15265);
nor U15805 (N_15805,N_15385,N_15484);
xor U15806 (N_15806,N_15235,N_15361);
xor U15807 (N_15807,N_15280,N_15194);
and U15808 (N_15808,N_15323,N_15368);
nor U15809 (N_15809,N_15340,N_15237);
xor U15810 (N_15810,N_15402,N_15428);
or U15811 (N_15811,N_15404,N_15280);
and U15812 (N_15812,N_15090,N_15035);
xor U15813 (N_15813,N_15306,N_15184);
and U15814 (N_15814,N_15267,N_15374);
xor U15815 (N_15815,N_15370,N_15231);
nor U15816 (N_15816,N_15446,N_15318);
xor U15817 (N_15817,N_15145,N_15173);
nand U15818 (N_15818,N_15070,N_15404);
or U15819 (N_15819,N_15279,N_15481);
nor U15820 (N_15820,N_15203,N_15387);
nor U15821 (N_15821,N_15381,N_15376);
xnor U15822 (N_15822,N_15409,N_15379);
or U15823 (N_15823,N_15162,N_15157);
nand U15824 (N_15824,N_15315,N_15402);
nor U15825 (N_15825,N_15362,N_15194);
nor U15826 (N_15826,N_15434,N_15429);
nor U15827 (N_15827,N_15105,N_15320);
and U15828 (N_15828,N_15391,N_15247);
and U15829 (N_15829,N_15236,N_15217);
xor U15830 (N_15830,N_15290,N_15224);
nand U15831 (N_15831,N_15322,N_15034);
and U15832 (N_15832,N_15492,N_15334);
nor U15833 (N_15833,N_15109,N_15427);
or U15834 (N_15834,N_15207,N_15468);
and U15835 (N_15835,N_15362,N_15266);
xnor U15836 (N_15836,N_15062,N_15453);
xor U15837 (N_15837,N_15228,N_15412);
nor U15838 (N_15838,N_15197,N_15170);
or U15839 (N_15839,N_15484,N_15339);
nand U15840 (N_15840,N_15286,N_15243);
xnor U15841 (N_15841,N_15207,N_15156);
nor U15842 (N_15842,N_15240,N_15342);
nor U15843 (N_15843,N_15217,N_15345);
and U15844 (N_15844,N_15317,N_15119);
nand U15845 (N_15845,N_15478,N_15274);
nand U15846 (N_15846,N_15204,N_15243);
nor U15847 (N_15847,N_15477,N_15425);
nor U15848 (N_15848,N_15008,N_15493);
and U15849 (N_15849,N_15473,N_15490);
nand U15850 (N_15850,N_15321,N_15424);
or U15851 (N_15851,N_15208,N_15148);
and U15852 (N_15852,N_15227,N_15234);
nor U15853 (N_15853,N_15226,N_15049);
and U15854 (N_15854,N_15281,N_15122);
xor U15855 (N_15855,N_15011,N_15251);
nand U15856 (N_15856,N_15194,N_15308);
and U15857 (N_15857,N_15131,N_15140);
and U15858 (N_15858,N_15344,N_15399);
nor U15859 (N_15859,N_15469,N_15244);
nor U15860 (N_15860,N_15385,N_15160);
or U15861 (N_15861,N_15295,N_15243);
or U15862 (N_15862,N_15354,N_15291);
nor U15863 (N_15863,N_15172,N_15006);
nand U15864 (N_15864,N_15257,N_15018);
or U15865 (N_15865,N_15086,N_15245);
or U15866 (N_15866,N_15159,N_15037);
or U15867 (N_15867,N_15050,N_15324);
and U15868 (N_15868,N_15409,N_15476);
or U15869 (N_15869,N_15426,N_15415);
nand U15870 (N_15870,N_15127,N_15292);
nand U15871 (N_15871,N_15478,N_15396);
and U15872 (N_15872,N_15334,N_15439);
nand U15873 (N_15873,N_15454,N_15202);
or U15874 (N_15874,N_15140,N_15086);
or U15875 (N_15875,N_15437,N_15175);
xnor U15876 (N_15876,N_15157,N_15437);
xnor U15877 (N_15877,N_15175,N_15389);
or U15878 (N_15878,N_15427,N_15250);
nand U15879 (N_15879,N_15454,N_15361);
nor U15880 (N_15880,N_15110,N_15427);
nand U15881 (N_15881,N_15133,N_15319);
nand U15882 (N_15882,N_15222,N_15067);
nand U15883 (N_15883,N_15463,N_15396);
or U15884 (N_15884,N_15133,N_15042);
nor U15885 (N_15885,N_15490,N_15379);
nand U15886 (N_15886,N_15227,N_15288);
and U15887 (N_15887,N_15400,N_15055);
and U15888 (N_15888,N_15294,N_15047);
nor U15889 (N_15889,N_15324,N_15016);
and U15890 (N_15890,N_15055,N_15445);
or U15891 (N_15891,N_15493,N_15097);
nand U15892 (N_15892,N_15207,N_15421);
xor U15893 (N_15893,N_15499,N_15467);
xnor U15894 (N_15894,N_15417,N_15259);
or U15895 (N_15895,N_15406,N_15415);
nand U15896 (N_15896,N_15259,N_15373);
or U15897 (N_15897,N_15262,N_15463);
nor U15898 (N_15898,N_15138,N_15480);
nor U15899 (N_15899,N_15286,N_15057);
xor U15900 (N_15900,N_15322,N_15207);
or U15901 (N_15901,N_15063,N_15382);
nand U15902 (N_15902,N_15277,N_15039);
nand U15903 (N_15903,N_15101,N_15012);
xor U15904 (N_15904,N_15412,N_15437);
nor U15905 (N_15905,N_15415,N_15164);
nor U15906 (N_15906,N_15305,N_15427);
nand U15907 (N_15907,N_15428,N_15177);
or U15908 (N_15908,N_15297,N_15318);
xnor U15909 (N_15909,N_15377,N_15439);
nor U15910 (N_15910,N_15352,N_15327);
xor U15911 (N_15911,N_15465,N_15383);
nand U15912 (N_15912,N_15134,N_15443);
nand U15913 (N_15913,N_15464,N_15387);
nand U15914 (N_15914,N_15392,N_15485);
xnor U15915 (N_15915,N_15327,N_15288);
nand U15916 (N_15916,N_15090,N_15208);
or U15917 (N_15917,N_15382,N_15100);
or U15918 (N_15918,N_15269,N_15487);
nand U15919 (N_15919,N_15494,N_15173);
nand U15920 (N_15920,N_15495,N_15317);
and U15921 (N_15921,N_15339,N_15457);
nor U15922 (N_15922,N_15134,N_15069);
or U15923 (N_15923,N_15147,N_15055);
and U15924 (N_15924,N_15089,N_15389);
and U15925 (N_15925,N_15230,N_15071);
nor U15926 (N_15926,N_15422,N_15246);
or U15927 (N_15927,N_15108,N_15086);
nand U15928 (N_15928,N_15448,N_15323);
nand U15929 (N_15929,N_15249,N_15203);
nor U15930 (N_15930,N_15084,N_15301);
nor U15931 (N_15931,N_15213,N_15464);
or U15932 (N_15932,N_15169,N_15489);
or U15933 (N_15933,N_15291,N_15199);
xor U15934 (N_15934,N_15084,N_15363);
nand U15935 (N_15935,N_15099,N_15235);
xnor U15936 (N_15936,N_15487,N_15413);
xnor U15937 (N_15937,N_15292,N_15386);
nand U15938 (N_15938,N_15483,N_15184);
nand U15939 (N_15939,N_15452,N_15432);
nand U15940 (N_15940,N_15414,N_15407);
nand U15941 (N_15941,N_15443,N_15279);
nand U15942 (N_15942,N_15213,N_15457);
xor U15943 (N_15943,N_15345,N_15419);
nand U15944 (N_15944,N_15031,N_15133);
and U15945 (N_15945,N_15320,N_15384);
nand U15946 (N_15946,N_15323,N_15382);
nor U15947 (N_15947,N_15209,N_15127);
nor U15948 (N_15948,N_15239,N_15179);
xor U15949 (N_15949,N_15251,N_15252);
nand U15950 (N_15950,N_15174,N_15178);
xnor U15951 (N_15951,N_15043,N_15203);
and U15952 (N_15952,N_15264,N_15015);
or U15953 (N_15953,N_15354,N_15038);
nand U15954 (N_15954,N_15148,N_15340);
nor U15955 (N_15955,N_15305,N_15311);
and U15956 (N_15956,N_15119,N_15070);
xnor U15957 (N_15957,N_15264,N_15416);
and U15958 (N_15958,N_15149,N_15166);
nor U15959 (N_15959,N_15100,N_15176);
and U15960 (N_15960,N_15001,N_15124);
and U15961 (N_15961,N_15223,N_15062);
nor U15962 (N_15962,N_15102,N_15065);
and U15963 (N_15963,N_15111,N_15277);
xor U15964 (N_15964,N_15221,N_15212);
nor U15965 (N_15965,N_15424,N_15392);
and U15966 (N_15966,N_15160,N_15098);
xor U15967 (N_15967,N_15027,N_15439);
or U15968 (N_15968,N_15017,N_15386);
nand U15969 (N_15969,N_15395,N_15261);
nand U15970 (N_15970,N_15407,N_15100);
or U15971 (N_15971,N_15496,N_15314);
nand U15972 (N_15972,N_15092,N_15474);
nand U15973 (N_15973,N_15367,N_15225);
nor U15974 (N_15974,N_15254,N_15218);
nand U15975 (N_15975,N_15274,N_15165);
or U15976 (N_15976,N_15016,N_15375);
and U15977 (N_15977,N_15380,N_15265);
xor U15978 (N_15978,N_15067,N_15454);
nand U15979 (N_15979,N_15087,N_15488);
and U15980 (N_15980,N_15401,N_15164);
nand U15981 (N_15981,N_15019,N_15455);
xnor U15982 (N_15982,N_15298,N_15230);
xor U15983 (N_15983,N_15067,N_15019);
nand U15984 (N_15984,N_15107,N_15253);
xor U15985 (N_15985,N_15358,N_15410);
nor U15986 (N_15986,N_15258,N_15209);
nor U15987 (N_15987,N_15278,N_15478);
xor U15988 (N_15988,N_15481,N_15475);
nand U15989 (N_15989,N_15297,N_15446);
xnor U15990 (N_15990,N_15410,N_15139);
nand U15991 (N_15991,N_15362,N_15208);
and U15992 (N_15992,N_15370,N_15191);
and U15993 (N_15993,N_15415,N_15261);
or U15994 (N_15994,N_15487,N_15482);
nand U15995 (N_15995,N_15336,N_15195);
or U15996 (N_15996,N_15401,N_15448);
and U15997 (N_15997,N_15275,N_15084);
nor U15998 (N_15998,N_15025,N_15426);
or U15999 (N_15999,N_15376,N_15491);
xor U16000 (N_16000,N_15946,N_15779);
and U16001 (N_16001,N_15603,N_15855);
xor U16002 (N_16002,N_15715,N_15961);
nor U16003 (N_16003,N_15842,N_15546);
xor U16004 (N_16004,N_15765,N_15767);
or U16005 (N_16005,N_15852,N_15692);
nand U16006 (N_16006,N_15722,N_15955);
nand U16007 (N_16007,N_15689,N_15510);
xor U16008 (N_16008,N_15557,N_15799);
nand U16009 (N_16009,N_15783,N_15817);
nor U16010 (N_16010,N_15820,N_15846);
nand U16011 (N_16011,N_15578,N_15571);
nor U16012 (N_16012,N_15832,N_15993);
nand U16013 (N_16013,N_15834,N_15534);
nor U16014 (N_16014,N_15562,N_15587);
nor U16015 (N_16015,N_15579,N_15784);
nand U16016 (N_16016,N_15851,N_15536);
and U16017 (N_16017,N_15941,N_15978);
and U16018 (N_16018,N_15705,N_15959);
or U16019 (N_16019,N_15998,N_15980);
or U16020 (N_16020,N_15861,N_15547);
nor U16021 (N_16021,N_15964,N_15836);
xnor U16022 (N_16022,N_15828,N_15673);
or U16023 (N_16023,N_15592,N_15633);
or U16024 (N_16024,N_15677,N_15656);
nor U16025 (N_16025,N_15801,N_15804);
nor U16026 (N_16026,N_15653,N_15521);
nor U16027 (N_16027,N_15843,N_15598);
nor U16028 (N_16028,N_15973,N_15771);
nand U16029 (N_16029,N_15872,N_15732);
or U16030 (N_16030,N_15582,N_15781);
or U16031 (N_16031,N_15697,N_15920);
and U16032 (N_16032,N_15654,N_15753);
xnor U16033 (N_16033,N_15948,N_15627);
and U16034 (N_16034,N_15687,N_15594);
nand U16035 (N_16035,N_15965,N_15962);
nor U16036 (N_16036,N_15706,N_15601);
nand U16037 (N_16037,N_15791,N_15577);
xnor U16038 (N_16038,N_15937,N_15927);
and U16039 (N_16039,N_15680,N_15575);
nor U16040 (N_16040,N_15768,N_15635);
nand U16041 (N_16041,N_15981,N_15874);
nand U16042 (N_16042,N_15584,N_15651);
nor U16043 (N_16043,N_15777,N_15803);
and U16044 (N_16044,N_15664,N_15714);
nor U16045 (N_16045,N_15985,N_15793);
or U16046 (N_16046,N_15674,N_15728);
or U16047 (N_16047,N_15869,N_15859);
or U16048 (N_16048,N_15759,N_15772);
or U16049 (N_16049,N_15883,N_15616);
and U16050 (N_16050,N_15602,N_15926);
nand U16051 (N_16051,N_15886,N_15966);
nor U16052 (N_16052,N_15888,N_15929);
xnor U16053 (N_16053,N_15893,N_15967);
nor U16054 (N_16054,N_15539,N_15750);
xnor U16055 (N_16055,N_15632,N_15560);
nand U16056 (N_16056,N_15770,N_15506);
nand U16057 (N_16057,N_15847,N_15625);
nor U16058 (N_16058,N_15502,N_15503);
or U16059 (N_16059,N_15566,N_15766);
xnor U16060 (N_16060,N_15564,N_15716);
and U16061 (N_16061,N_15897,N_15911);
nor U16062 (N_16062,N_15942,N_15544);
xor U16063 (N_16063,N_15563,N_15902);
nand U16064 (N_16064,N_15854,N_15565);
nand U16065 (N_16065,N_15830,N_15554);
or U16066 (N_16066,N_15821,N_15933);
nand U16067 (N_16067,N_15637,N_15943);
nor U16068 (N_16068,N_15761,N_15889);
and U16069 (N_16069,N_15829,N_15958);
xor U16070 (N_16070,N_15800,N_15658);
xnor U16071 (N_16071,N_15763,N_15556);
and U16072 (N_16072,N_15553,N_15516);
xnor U16073 (N_16073,N_15994,N_15811);
xnor U16074 (N_16074,N_15940,N_15909);
and U16075 (N_16075,N_15641,N_15990);
and U16076 (N_16076,N_15736,N_15605);
and U16077 (N_16077,N_15682,N_15744);
and U16078 (N_16078,N_15899,N_15528);
or U16079 (N_16079,N_15600,N_15758);
and U16080 (N_16080,N_15729,N_15691);
and U16081 (N_16081,N_15809,N_15936);
xnor U16082 (N_16082,N_15860,N_15754);
nor U16083 (N_16083,N_15535,N_15631);
or U16084 (N_16084,N_15573,N_15794);
or U16085 (N_16085,N_15552,N_15514);
and U16086 (N_16086,N_15660,N_15504);
and U16087 (N_16087,N_15662,N_15898);
nand U16088 (N_16088,N_15649,N_15645);
nor U16089 (N_16089,N_15796,N_15996);
nor U16090 (N_16090,N_15953,N_15922);
or U16091 (N_16091,N_15717,N_15576);
xnor U16092 (N_16092,N_15963,N_15650);
or U16093 (N_16093,N_15885,N_15542);
nand U16094 (N_16094,N_15919,N_15760);
nand U16095 (N_16095,N_15976,N_15591);
or U16096 (N_16096,N_15707,N_15526);
and U16097 (N_16097,N_15731,N_15630);
nand U16098 (N_16098,N_15703,N_15895);
or U16099 (N_16099,N_15686,N_15730);
xnor U16100 (N_16100,N_15853,N_15696);
or U16101 (N_16101,N_15815,N_15537);
or U16102 (N_16102,N_15798,N_15585);
xor U16103 (N_16103,N_15999,N_15621);
or U16104 (N_16104,N_15988,N_15873);
and U16105 (N_16105,N_15904,N_15570);
or U16106 (N_16106,N_15708,N_15727);
or U16107 (N_16107,N_15841,N_15887);
xor U16108 (N_16108,N_15702,N_15878);
xor U16109 (N_16109,N_15524,N_15550);
or U16110 (N_16110,N_15529,N_15835);
xnor U16111 (N_16111,N_15523,N_15548);
nand U16112 (N_16112,N_15527,N_15757);
xor U16113 (N_16113,N_15833,N_15808);
or U16114 (N_16114,N_15620,N_15741);
nor U16115 (N_16115,N_15541,N_15956);
and U16116 (N_16116,N_15979,N_15655);
nor U16117 (N_16117,N_15839,N_15928);
nor U16118 (N_16118,N_15814,N_15877);
xor U16119 (N_16119,N_15675,N_15905);
and U16120 (N_16120,N_15991,N_15995);
xnor U16121 (N_16121,N_15572,N_15950);
nor U16122 (N_16122,N_15824,N_15612);
and U16123 (N_16123,N_15915,N_15825);
and U16124 (N_16124,N_15826,N_15756);
and U16125 (N_16125,N_15989,N_15509);
nand U16126 (N_16126,N_15543,N_15951);
nor U16127 (N_16127,N_15501,N_15567);
and U16128 (N_16128,N_15642,N_15609);
or U16129 (N_16129,N_15983,N_15780);
or U16130 (N_16130,N_15969,N_15850);
xnor U16131 (N_16131,N_15634,N_15845);
and U16132 (N_16132,N_15644,N_15734);
nor U16133 (N_16133,N_15975,N_15623);
and U16134 (N_16134,N_15685,N_15724);
or U16135 (N_16135,N_15711,N_15738);
nor U16136 (N_16136,N_15595,N_15607);
nor U16137 (N_16137,N_15619,N_15880);
and U16138 (N_16138,N_15792,N_15788);
and U16139 (N_16139,N_15661,N_15856);
or U16140 (N_16140,N_15617,N_15517);
or U16141 (N_16141,N_15701,N_15533);
and U16142 (N_16142,N_15522,N_15789);
and U16143 (N_16143,N_15752,N_15790);
nor U16144 (N_16144,N_15626,N_15984);
and U16145 (N_16145,N_15508,N_15912);
and U16146 (N_16146,N_15906,N_15806);
and U16147 (N_16147,N_15676,N_15900);
xnor U16148 (N_16148,N_15666,N_15913);
xnor U16149 (N_16149,N_15511,N_15597);
nand U16150 (N_16150,N_15986,N_15818);
xnor U16151 (N_16151,N_15745,N_15870);
and U16152 (N_16152,N_15785,N_15774);
or U16153 (N_16153,N_15954,N_15723);
nand U16154 (N_16154,N_15797,N_15775);
nand U16155 (N_16155,N_15823,N_15987);
nand U16156 (N_16156,N_15901,N_15590);
or U16157 (N_16157,N_15862,N_15588);
nor U16158 (N_16158,N_15709,N_15669);
xor U16159 (N_16159,N_15949,N_15879);
and U16160 (N_16160,N_15581,N_15652);
nor U16161 (N_16161,N_15810,N_15944);
nor U16162 (N_16162,N_15740,N_15606);
nand U16163 (N_16163,N_15646,N_15586);
nor U16164 (N_16164,N_15871,N_15518);
nand U16165 (N_16165,N_15977,N_15934);
and U16166 (N_16166,N_15917,N_15907);
and U16167 (N_16167,N_15840,N_15742);
nor U16168 (N_16168,N_15894,N_15891);
nor U16169 (N_16169,N_15684,N_15678);
nor U16170 (N_16170,N_15671,N_15938);
and U16171 (N_16171,N_15726,N_15787);
or U16172 (N_16172,N_15713,N_15749);
nor U16173 (N_16173,N_15735,N_15694);
nand U16174 (N_16174,N_15663,N_15935);
and U16175 (N_16175,N_15532,N_15599);
nand U16176 (N_16176,N_15712,N_15764);
nand U16177 (N_16177,N_15812,N_15589);
nand U16178 (N_16178,N_15849,N_15704);
and U16179 (N_16179,N_15515,N_15875);
nor U16180 (N_16180,N_15569,N_15970);
nor U16181 (N_16181,N_15568,N_15972);
xor U16182 (N_16182,N_15921,N_15957);
nand U16183 (N_16183,N_15838,N_15672);
or U16184 (N_16184,N_15884,N_15903);
and U16185 (N_16185,N_15540,N_15876);
nor U16186 (N_16186,N_15580,N_15558);
nand U16187 (N_16187,N_15507,N_15992);
nand U16188 (N_16188,N_15545,N_15802);
nand U16189 (N_16189,N_15593,N_15866);
and U16190 (N_16190,N_15688,N_15916);
or U16191 (N_16191,N_15968,N_15925);
xor U16192 (N_16192,N_15939,N_15512);
xnor U16193 (N_16193,N_15604,N_15683);
nand U16194 (N_16194,N_15947,N_15746);
nand U16195 (N_16195,N_15743,N_15699);
or U16196 (N_16196,N_15538,N_15690);
or U16197 (N_16197,N_15945,N_15908);
nand U16198 (N_16198,N_15596,N_15881);
nand U16199 (N_16199,N_15882,N_15896);
nand U16200 (N_16200,N_15613,N_15618);
or U16201 (N_16201,N_15762,N_15831);
xor U16202 (N_16202,N_15932,N_15561);
or U16203 (N_16203,N_15681,N_15863);
xnor U16204 (N_16204,N_15721,N_15776);
nor U16205 (N_16205,N_15782,N_15747);
or U16206 (N_16206,N_15519,N_15622);
nand U16207 (N_16207,N_15816,N_15748);
xor U16208 (N_16208,N_15807,N_15555);
nand U16209 (N_16209,N_15559,N_15648);
or U16210 (N_16210,N_15813,N_15773);
or U16211 (N_16211,N_15647,N_15868);
xor U16212 (N_16212,N_15638,N_15710);
and U16213 (N_16213,N_15520,N_15629);
nor U16214 (N_16214,N_15525,N_15615);
and U16215 (N_16215,N_15924,N_15914);
xor U16216 (N_16216,N_15574,N_15657);
nand U16217 (N_16217,N_15551,N_15864);
or U16218 (N_16218,N_15695,N_15670);
nand U16219 (N_16219,N_15837,N_15805);
xor U16220 (N_16220,N_15890,N_15720);
or U16221 (N_16221,N_15931,N_15718);
and U16222 (N_16222,N_15997,N_15930);
nor U16223 (N_16223,N_15659,N_15624);
and U16224 (N_16224,N_15739,N_15865);
nor U16225 (N_16225,N_15858,N_15500);
xnor U16226 (N_16226,N_15733,N_15918);
or U16227 (N_16227,N_15698,N_15530);
or U16228 (N_16228,N_15549,N_15639);
or U16229 (N_16229,N_15923,N_15892);
nand U16230 (N_16230,N_15700,N_15819);
xnor U16231 (N_16231,N_15971,N_15667);
nand U16232 (N_16232,N_15668,N_15867);
nand U16233 (N_16233,N_15628,N_15614);
or U16234 (N_16234,N_15725,N_15844);
nand U16235 (N_16235,N_15505,N_15778);
nand U16236 (N_16236,N_15531,N_15719);
xor U16237 (N_16237,N_15737,N_15848);
or U16238 (N_16238,N_15822,N_15769);
xor U16239 (N_16239,N_15583,N_15952);
and U16240 (N_16240,N_15636,N_15640);
nand U16241 (N_16241,N_15960,N_15982);
nor U16242 (N_16242,N_15610,N_15974);
and U16243 (N_16243,N_15513,N_15608);
and U16244 (N_16244,N_15643,N_15679);
nor U16245 (N_16245,N_15786,N_15795);
xor U16246 (N_16246,N_15857,N_15665);
and U16247 (N_16247,N_15827,N_15755);
or U16248 (N_16248,N_15693,N_15751);
and U16249 (N_16249,N_15611,N_15910);
xnor U16250 (N_16250,N_15772,N_15566);
or U16251 (N_16251,N_15584,N_15662);
or U16252 (N_16252,N_15642,N_15554);
or U16253 (N_16253,N_15916,N_15553);
or U16254 (N_16254,N_15853,N_15765);
xnor U16255 (N_16255,N_15795,N_15565);
nand U16256 (N_16256,N_15712,N_15901);
xnor U16257 (N_16257,N_15762,N_15965);
and U16258 (N_16258,N_15672,N_15904);
nand U16259 (N_16259,N_15765,N_15638);
or U16260 (N_16260,N_15977,N_15600);
nand U16261 (N_16261,N_15629,N_15563);
xor U16262 (N_16262,N_15758,N_15977);
or U16263 (N_16263,N_15982,N_15869);
nand U16264 (N_16264,N_15741,N_15821);
nor U16265 (N_16265,N_15812,N_15780);
and U16266 (N_16266,N_15902,N_15748);
nor U16267 (N_16267,N_15785,N_15968);
and U16268 (N_16268,N_15891,N_15957);
xnor U16269 (N_16269,N_15643,N_15879);
nor U16270 (N_16270,N_15868,N_15927);
or U16271 (N_16271,N_15828,N_15647);
nor U16272 (N_16272,N_15817,N_15865);
nor U16273 (N_16273,N_15942,N_15502);
nor U16274 (N_16274,N_15700,N_15714);
or U16275 (N_16275,N_15616,N_15556);
nor U16276 (N_16276,N_15987,N_15801);
and U16277 (N_16277,N_15820,N_15879);
nor U16278 (N_16278,N_15833,N_15650);
and U16279 (N_16279,N_15707,N_15952);
nor U16280 (N_16280,N_15571,N_15597);
nor U16281 (N_16281,N_15733,N_15539);
nand U16282 (N_16282,N_15882,N_15759);
and U16283 (N_16283,N_15733,N_15805);
or U16284 (N_16284,N_15859,N_15513);
and U16285 (N_16285,N_15716,N_15625);
nor U16286 (N_16286,N_15818,N_15648);
xor U16287 (N_16287,N_15544,N_15892);
and U16288 (N_16288,N_15860,N_15561);
nor U16289 (N_16289,N_15805,N_15657);
xnor U16290 (N_16290,N_15841,N_15806);
xor U16291 (N_16291,N_15762,N_15766);
nand U16292 (N_16292,N_15561,N_15913);
nor U16293 (N_16293,N_15633,N_15818);
and U16294 (N_16294,N_15668,N_15932);
nor U16295 (N_16295,N_15801,N_15755);
or U16296 (N_16296,N_15758,N_15980);
nand U16297 (N_16297,N_15926,N_15569);
nand U16298 (N_16298,N_15702,N_15951);
and U16299 (N_16299,N_15933,N_15612);
or U16300 (N_16300,N_15973,N_15669);
or U16301 (N_16301,N_15730,N_15949);
xnor U16302 (N_16302,N_15813,N_15741);
or U16303 (N_16303,N_15870,N_15705);
nand U16304 (N_16304,N_15619,N_15884);
or U16305 (N_16305,N_15602,N_15674);
xor U16306 (N_16306,N_15755,N_15747);
xnor U16307 (N_16307,N_15819,N_15781);
and U16308 (N_16308,N_15857,N_15602);
xor U16309 (N_16309,N_15998,N_15945);
nand U16310 (N_16310,N_15777,N_15517);
and U16311 (N_16311,N_15851,N_15609);
and U16312 (N_16312,N_15757,N_15840);
xor U16313 (N_16313,N_15742,N_15868);
nand U16314 (N_16314,N_15882,N_15641);
nor U16315 (N_16315,N_15583,N_15942);
xor U16316 (N_16316,N_15848,N_15883);
nor U16317 (N_16317,N_15914,N_15695);
nand U16318 (N_16318,N_15541,N_15729);
or U16319 (N_16319,N_15804,N_15943);
or U16320 (N_16320,N_15919,N_15889);
nor U16321 (N_16321,N_15918,N_15796);
nand U16322 (N_16322,N_15721,N_15507);
xnor U16323 (N_16323,N_15555,N_15863);
and U16324 (N_16324,N_15851,N_15598);
and U16325 (N_16325,N_15816,N_15963);
nand U16326 (N_16326,N_15613,N_15767);
nor U16327 (N_16327,N_15703,N_15999);
and U16328 (N_16328,N_15843,N_15899);
xnor U16329 (N_16329,N_15559,N_15594);
nor U16330 (N_16330,N_15802,N_15816);
xnor U16331 (N_16331,N_15649,N_15705);
or U16332 (N_16332,N_15564,N_15868);
nand U16333 (N_16333,N_15609,N_15636);
and U16334 (N_16334,N_15974,N_15526);
nand U16335 (N_16335,N_15810,N_15563);
or U16336 (N_16336,N_15932,N_15956);
and U16337 (N_16337,N_15910,N_15882);
nor U16338 (N_16338,N_15705,N_15603);
and U16339 (N_16339,N_15524,N_15972);
or U16340 (N_16340,N_15575,N_15936);
nand U16341 (N_16341,N_15506,N_15879);
or U16342 (N_16342,N_15769,N_15615);
or U16343 (N_16343,N_15770,N_15514);
and U16344 (N_16344,N_15804,N_15544);
and U16345 (N_16345,N_15807,N_15998);
nor U16346 (N_16346,N_15522,N_15783);
nor U16347 (N_16347,N_15610,N_15756);
nand U16348 (N_16348,N_15679,N_15955);
nand U16349 (N_16349,N_15788,N_15728);
or U16350 (N_16350,N_15661,N_15919);
nor U16351 (N_16351,N_15595,N_15816);
nand U16352 (N_16352,N_15518,N_15517);
xnor U16353 (N_16353,N_15737,N_15812);
nand U16354 (N_16354,N_15614,N_15931);
and U16355 (N_16355,N_15633,N_15973);
nand U16356 (N_16356,N_15916,N_15635);
nor U16357 (N_16357,N_15759,N_15634);
and U16358 (N_16358,N_15727,N_15917);
or U16359 (N_16359,N_15974,N_15920);
xnor U16360 (N_16360,N_15823,N_15787);
nand U16361 (N_16361,N_15701,N_15583);
nand U16362 (N_16362,N_15709,N_15852);
and U16363 (N_16363,N_15828,N_15676);
nand U16364 (N_16364,N_15886,N_15742);
or U16365 (N_16365,N_15782,N_15899);
nand U16366 (N_16366,N_15699,N_15584);
and U16367 (N_16367,N_15805,N_15868);
and U16368 (N_16368,N_15859,N_15607);
or U16369 (N_16369,N_15659,N_15592);
or U16370 (N_16370,N_15672,N_15996);
nor U16371 (N_16371,N_15672,N_15689);
nor U16372 (N_16372,N_15979,N_15717);
or U16373 (N_16373,N_15576,N_15671);
nor U16374 (N_16374,N_15577,N_15712);
or U16375 (N_16375,N_15545,N_15690);
nand U16376 (N_16376,N_15516,N_15724);
nor U16377 (N_16377,N_15606,N_15984);
nor U16378 (N_16378,N_15987,N_15860);
and U16379 (N_16379,N_15586,N_15848);
nor U16380 (N_16380,N_15769,N_15573);
or U16381 (N_16381,N_15996,N_15879);
xnor U16382 (N_16382,N_15580,N_15676);
xnor U16383 (N_16383,N_15786,N_15631);
or U16384 (N_16384,N_15670,N_15851);
nor U16385 (N_16385,N_15679,N_15642);
and U16386 (N_16386,N_15557,N_15603);
and U16387 (N_16387,N_15778,N_15684);
nand U16388 (N_16388,N_15543,N_15744);
nor U16389 (N_16389,N_15917,N_15795);
nor U16390 (N_16390,N_15683,N_15851);
nor U16391 (N_16391,N_15628,N_15753);
nand U16392 (N_16392,N_15639,N_15576);
xnor U16393 (N_16393,N_15998,N_15882);
and U16394 (N_16394,N_15714,N_15638);
nor U16395 (N_16395,N_15936,N_15854);
and U16396 (N_16396,N_15888,N_15547);
xnor U16397 (N_16397,N_15820,N_15866);
nand U16398 (N_16398,N_15750,N_15992);
and U16399 (N_16399,N_15510,N_15682);
and U16400 (N_16400,N_15858,N_15880);
nor U16401 (N_16401,N_15608,N_15952);
and U16402 (N_16402,N_15835,N_15649);
xor U16403 (N_16403,N_15767,N_15539);
nand U16404 (N_16404,N_15703,N_15567);
and U16405 (N_16405,N_15855,N_15589);
nand U16406 (N_16406,N_15693,N_15878);
nor U16407 (N_16407,N_15645,N_15856);
nand U16408 (N_16408,N_15520,N_15567);
nand U16409 (N_16409,N_15594,N_15601);
nor U16410 (N_16410,N_15693,N_15533);
nor U16411 (N_16411,N_15777,N_15686);
and U16412 (N_16412,N_15889,N_15781);
xnor U16413 (N_16413,N_15907,N_15711);
nor U16414 (N_16414,N_15936,N_15704);
or U16415 (N_16415,N_15696,N_15902);
nand U16416 (N_16416,N_15808,N_15555);
and U16417 (N_16417,N_15723,N_15711);
nand U16418 (N_16418,N_15728,N_15916);
xnor U16419 (N_16419,N_15527,N_15611);
and U16420 (N_16420,N_15831,N_15808);
and U16421 (N_16421,N_15638,N_15855);
or U16422 (N_16422,N_15772,N_15560);
nor U16423 (N_16423,N_15634,N_15853);
nand U16424 (N_16424,N_15915,N_15550);
and U16425 (N_16425,N_15581,N_15899);
or U16426 (N_16426,N_15888,N_15783);
and U16427 (N_16427,N_15844,N_15878);
and U16428 (N_16428,N_15667,N_15785);
or U16429 (N_16429,N_15974,N_15783);
xor U16430 (N_16430,N_15561,N_15556);
xnor U16431 (N_16431,N_15889,N_15521);
nand U16432 (N_16432,N_15628,N_15671);
nand U16433 (N_16433,N_15906,N_15514);
nand U16434 (N_16434,N_15943,N_15675);
xnor U16435 (N_16435,N_15811,N_15950);
nand U16436 (N_16436,N_15897,N_15965);
or U16437 (N_16437,N_15956,N_15689);
nand U16438 (N_16438,N_15928,N_15509);
and U16439 (N_16439,N_15765,N_15581);
nand U16440 (N_16440,N_15836,N_15919);
and U16441 (N_16441,N_15965,N_15693);
nand U16442 (N_16442,N_15816,N_15753);
nand U16443 (N_16443,N_15759,N_15860);
nand U16444 (N_16444,N_15936,N_15715);
nor U16445 (N_16445,N_15709,N_15513);
or U16446 (N_16446,N_15592,N_15632);
and U16447 (N_16447,N_15659,N_15586);
xnor U16448 (N_16448,N_15668,N_15603);
xnor U16449 (N_16449,N_15865,N_15921);
or U16450 (N_16450,N_15903,N_15708);
nand U16451 (N_16451,N_15964,N_15556);
nor U16452 (N_16452,N_15824,N_15712);
and U16453 (N_16453,N_15570,N_15852);
xor U16454 (N_16454,N_15914,N_15771);
or U16455 (N_16455,N_15678,N_15865);
xnor U16456 (N_16456,N_15793,N_15518);
nor U16457 (N_16457,N_15950,N_15645);
and U16458 (N_16458,N_15912,N_15564);
nand U16459 (N_16459,N_15563,N_15610);
nand U16460 (N_16460,N_15577,N_15618);
nor U16461 (N_16461,N_15537,N_15991);
xnor U16462 (N_16462,N_15530,N_15884);
and U16463 (N_16463,N_15974,N_15734);
or U16464 (N_16464,N_15506,N_15576);
nand U16465 (N_16465,N_15644,N_15874);
and U16466 (N_16466,N_15947,N_15564);
xnor U16467 (N_16467,N_15684,N_15528);
nor U16468 (N_16468,N_15576,N_15841);
xnor U16469 (N_16469,N_15978,N_15677);
nor U16470 (N_16470,N_15626,N_15962);
or U16471 (N_16471,N_15730,N_15931);
and U16472 (N_16472,N_15650,N_15867);
or U16473 (N_16473,N_15738,N_15687);
nand U16474 (N_16474,N_15713,N_15903);
nor U16475 (N_16475,N_15943,N_15998);
and U16476 (N_16476,N_15831,N_15972);
nand U16477 (N_16477,N_15532,N_15535);
nand U16478 (N_16478,N_15976,N_15550);
nand U16479 (N_16479,N_15688,N_15647);
nand U16480 (N_16480,N_15850,N_15659);
or U16481 (N_16481,N_15730,N_15651);
xnor U16482 (N_16482,N_15882,N_15965);
xnor U16483 (N_16483,N_15889,N_15597);
nor U16484 (N_16484,N_15511,N_15658);
xor U16485 (N_16485,N_15500,N_15741);
and U16486 (N_16486,N_15579,N_15510);
and U16487 (N_16487,N_15680,N_15706);
nand U16488 (N_16488,N_15596,N_15890);
or U16489 (N_16489,N_15856,N_15892);
nand U16490 (N_16490,N_15783,N_15623);
and U16491 (N_16491,N_15752,N_15881);
nor U16492 (N_16492,N_15699,N_15891);
and U16493 (N_16493,N_15570,N_15501);
or U16494 (N_16494,N_15508,N_15959);
xnor U16495 (N_16495,N_15673,N_15738);
nor U16496 (N_16496,N_15600,N_15566);
nor U16497 (N_16497,N_15681,N_15975);
xor U16498 (N_16498,N_15620,N_15575);
xor U16499 (N_16499,N_15508,N_15934);
nor U16500 (N_16500,N_16371,N_16270);
xnor U16501 (N_16501,N_16059,N_16286);
nand U16502 (N_16502,N_16476,N_16093);
nand U16503 (N_16503,N_16195,N_16063);
nand U16504 (N_16504,N_16216,N_16243);
nand U16505 (N_16505,N_16478,N_16061);
or U16506 (N_16506,N_16322,N_16277);
or U16507 (N_16507,N_16126,N_16365);
and U16508 (N_16508,N_16235,N_16328);
nor U16509 (N_16509,N_16483,N_16289);
nor U16510 (N_16510,N_16383,N_16450);
or U16511 (N_16511,N_16074,N_16143);
nand U16512 (N_16512,N_16395,N_16340);
or U16513 (N_16513,N_16106,N_16229);
nor U16514 (N_16514,N_16454,N_16125);
nand U16515 (N_16515,N_16141,N_16110);
or U16516 (N_16516,N_16276,N_16342);
nand U16517 (N_16517,N_16188,N_16288);
nor U16518 (N_16518,N_16209,N_16344);
nand U16519 (N_16519,N_16248,N_16055);
xor U16520 (N_16520,N_16267,N_16274);
or U16521 (N_16521,N_16396,N_16298);
nor U16522 (N_16522,N_16048,N_16088);
nand U16523 (N_16523,N_16256,N_16439);
or U16524 (N_16524,N_16182,N_16479);
xnor U16525 (N_16525,N_16324,N_16217);
nor U16526 (N_16526,N_16201,N_16473);
nor U16527 (N_16527,N_16482,N_16013);
nand U16528 (N_16528,N_16161,N_16004);
and U16529 (N_16529,N_16017,N_16131);
xnor U16530 (N_16530,N_16357,N_16127);
or U16531 (N_16531,N_16121,N_16087);
xor U16532 (N_16532,N_16065,N_16242);
and U16533 (N_16533,N_16260,N_16046);
or U16534 (N_16534,N_16435,N_16296);
nand U16535 (N_16535,N_16347,N_16230);
nand U16536 (N_16536,N_16374,N_16358);
nor U16537 (N_16537,N_16052,N_16490);
and U16538 (N_16538,N_16191,N_16255);
and U16539 (N_16539,N_16429,N_16027);
xnor U16540 (N_16540,N_16175,N_16354);
or U16541 (N_16541,N_16149,N_16254);
and U16542 (N_16542,N_16169,N_16067);
nor U16543 (N_16543,N_16107,N_16453);
xor U16544 (N_16544,N_16163,N_16001);
or U16545 (N_16545,N_16146,N_16128);
nor U16546 (N_16546,N_16299,N_16071);
nor U16547 (N_16547,N_16484,N_16292);
xor U16548 (N_16548,N_16335,N_16011);
nor U16549 (N_16549,N_16204,N_16398);
or U16550 (N_16550,N_16041,N_16302);
or U16551 (N_16551,N_16236,N_16238);
nand U16552 (N_16552,N_16372,N_16198);
xnor U16553 (N_16553,N_16040,N_16311);
xnor U16554 (N_16554,N_16069,N_16233);
or U16555 (N_16555,N_16221,N_16187);
and U16556 (N_16556,N_16232,N_16389);
xnor U16557 (N_16557,N_16464,N_16376);
xnor U16558 (N_16558,N_16100,N_16437);
and U16559 (N_16559,N_16446,N_16316);
nor U16560 (N_16560,N_16142,N_16402);
xnor U16561 (N_16561,N_16317,N_16393);
nor U16562 (N_16562,N_16291,N_16321);
nor U16563 (N_16563,N_16045,N_16240);
nand U16564 (N_16564,N_16047,N_16377);
nand U16565 (N_16565,N_16480,N_16179);
nand U16566 (N_16566,N_16370,N_16152);
xor U16567 (N_16567,N_16250,N_16207);
and U16568 (N_16568,N_16213,N_16012);
xor U16569 (N_16569,N_16290,N_16266);
xnor U16570 (N_16570,N_16010,N_16083);
nor U16571 (N_16571,N_16475,N_16186);
nand U16572 (N_16572,N_16094,N_16352);
or U16573 (N_16573,N_16024,N_16447);
xnor U16574 (N_16574,N_16399,N_16463);
xnor U16575 (N_16575,N_16105,N_16481);
nand U16576 (N_16576,N_16486,N_16005);
nor U16577 (N_16577,N_16109,N_16026);
or U16578 (N_16578,N_16456,N_16190);
and U16579 (N_16579,N_16348,N_16058);
and U16580 (N_16580,N_16408,N_16387);
xnor U16581 (N_16581,N_16323,N_16303);
and U16582 (N_16582,N_16325,N_16409);
xnor U16583 (N_16583,N_16223,N_16102);
nor U16584 (N_16584,N_16258,N_16029);
nor U16585 (N_16585,N_16155,N_16444);
nor U16586 (N_16586,N_16022,N_16312);
or U16587 (N_16587,N_16440,N_16037);
xor U16588 (N_16588,N_16438,N_16042);
nand U16589 (N_16589,N_16313,N_16097);
or U16590 (N_16590,N_16412,N_16355);
nand U16591 (N_16591,N_16382,N_16319);
nor U16592 (N_16592,N_16060,N_16489);
xor U16593 (N_16593,N_16451,N_16452);
or U16594 (N_16594,N_16492,N_16305);
or U16595 (N_16595,N_16318,N_16044);
xor U16596 (N_16596,N_16089,N_16193);
or U16597 (N_16597,N_16346,N_16062);
nand U16598 (N_16598,N_16417,N_16057);
nor U16599 (N_16599,N_16096,N_16337);
xor U16600 (N_16600,N_16279,N_16332);
xnor U16601 (N_16601,N_16420,N_16368);
nor U16602 (N_16602,N_16210,N_16173);
and U16603 (N_16603,N_16016,N_16356);
xnor U16604 (N_16604,N_16028,N_16416);
or U16605 (N_16605,N_16499,N_16261);
or U16606 (N_16606,N_16252,N_16111);
nor U16607 (N_16607,N_16075,N_16426);
or U16608 (N_16608,N_16158,N_16113);
nand U16609 (N_16609,N_16397,N_16284);
nand U16610 (N_16610,N_16234,N_16474);
nor U16611 (N_16611,N_16331,N_16135);
xnor U16612 (N_16612,N_16414,N_16369);
nand U16613 (N_16613,N_16086,N_16036);
or U16614 (N_16614,N_16390,N_16225);
nand U16615 (N_16615,N_16461,N_16345);
xnor U16616 (N_16616,N_16167,N_16031);
xor U16617 (N_16617,N_16441,N_16310);
nand U16618 (N_16618,N_16467,N_16206);
nand U16619 (N_16619,N_16320,N_16156);
nor U16620 (N_16620,N_16386,N_16278);
xor U16621 (N_16621,N_16264,N_16160);
nor U16622 (N_16622,N_16053,N_16080);
nand U16623 (N_16623,N_16251,N_16419);
nor U16624 (N_16624,N_16038,N_16023);
xnor U16625 (N_16625,N_16073,N_16066);
nor U16626 (N_16626,N_16424,N_16388);
nand U16627 (N_16627,N_16306,N_16498);
and U16628 (N_16628,N_16297,N_16485);
and U16629 (N_16629,N_16431,N_16039);
nand U16630 (N_16630,N_16007,N_16018);
and U16631 (N_16631,N_16090,N_16129);
xor U16632 (N_16632,N_16140,N_16147);
or U16633 (N_16633,N_16470,N_16380);
or U16634 (N_16634,N_16082,N_16008);
xor U16635 (N_16635,N_16427,N_16084);
xor U16636 (N_16636,N_16384,N_16137);
xnor U16637 (N_16637,N_16469,N_16391);
and U16638 (N_16638,N_16448,N_16488);
nor U16639 (N_16639,N_16425,N_16361);
and U16640 (N_16640,N_16056,N_16253);
nor U16641 (N_16641,N_16280,N_16123);
nand U16642 (N_16642,N_16285,N_16034);
xor U16643 (N_16643,N_16339,N_16184);
or U16644 (N_16644,N_16363,N_16268);
or U16645 (N_16645,N_16226,N_16237);
and U16646 (N_16646,N_16367,N_16085);
xnor U16647 (N_16647,N_16176,N_16049);
or U16648 (N_16648,N_16199,N_16019);
and U16649 (N_16649,N_16466,N_16183);
or U16650 (N_16650,N_16436,N_16154);
nor U16651 (N_16651,N_16406,N_16117);
nor U16652 (N_16652,N_16433,N_16170);
and U16653 (N_16653,N_16468,N_16497);
nand U16654 (N_16654,N_16304,N_16457);
xor U16655 (N_16655,N_16445,N_16212);
nor U16656 (N_16656,N_16403,N_16244);
xnor U16657 (N_16657,N_16079,N_16021);
or U16658 (N_16658,N_16112,N_16178);
and U16659 (N_16659,N_16458,N_16118);
nor U16660 (N_16660,N_16373,N_16275);
nor U16661 (N_16661,N_16308,N_16145);
nand U16662 (N_16662,N_16000,N_16157);
xor U16663 (N_16663,N_16078,N_16379);
nor U16664 (N_16664,N_16231,N_16465);
or U16665 (N_16665,N_16164,N_16491);
and U16666 (N_16666,N_16300,N_16050);
xnor U16667 (N_16667,N_16460,N_16459);
nor U16668 (N_16668,N_16366,N_16418);
and U16669 (N_16669,N_16189,N_16002);
and U16670 (N_16670,N_16407,N_16385);
xnor U16671 (N_16671,N_16185,N_16272);
xnor U16672 (N_16672,N_16428,N_16294);
xor U16673 (N_16673,N_16330,N_16177);
and U16674 (N_16674,N_16077,N_16220);
and U16675 (N_16675,N_16421,N_16341);
nand U16676 (N_16676,N_16401,N_16430);
nand U16677 (N_16677,N_16181,N_16477);
nor U16678 (N_16678,N_16130,N_16032);
nor U16679 (N_16679,N_16283,N_16334);
nand U16680 (N_16680,N_16494,N_16196);
or U16681 (N_16681,N_16434,N_16133);
nand U16682 (N_16682,N_16104,N_16114);
nand U16683 (N_16683,N_16134,N_16336);
nand U16684 (N_16684,N_16314,N_16168);
or U16685 (N_16685,N_16215,N_16350);
or U16686 (N_16686,N_16211,N_16092);
xnor U16687 (N_16687,N_16122,N_16404);
nand U16688 (N_16688,N_16263,N_16159);
and U16689 (N_16689,N_16455,N_16151);
nand U16690 (N_16690,N_16072,N_16076);
or U16691 (N_16691,N_16394,N_16360);
and U16692 (N_16692,N_16315,N_16364);
nand U16693 (N_16693,N_16003,N_16124);
nor U16694 (N_16694,N_16172,N_16165);
nand U16695 (N_16695,N_16194,N_16353);
nor U16696 (N_16696,N_16224,N_16015);
nand U16697 (N_16697,N_16033,N_16192);
or U16698 (N_16698,N_16043,N_16246);
nor U16699 (N_16699,N_16281,N_16095);
or U16700 (N_16700,N_16228,N_16171);
nor U16701 (N_16701,N_16472,N_16293);
nor U16702 (N_16702,N_16262,N_16116);
xnor U16703 (N_16703,N_16271,N_16227);
xnor U16704 (N_16704,N_16257,N_16423);
and U16705 (N_16705,N_16265,N_16282);
or U16706 (N_16706,N_16241,N_16139);
xnor U16707 (N_16707,N_16343,N_16239);
nand U16708 (N_16708,N_16120,N_16245);
xnor U16709 (N_16709,N_16349,N_16411);
nor U16710 (N_16710,N_16020,N_16442);
or U16711 (N_16711,N_16070,N_16351);
nand U16712 (N_16712,N_16327,N_16108);
or U16713 (N_16713,N_16115,N_16091);
xnor U16714 (N_16714,N_16051,N_16030);
xor U16715 (N_16715,N_16392,N_16400);
or U16716 (N_16716,N_16247,N_16099);
or U16717 (N_16717,N_16259,N_16362);
xnor U16718 (N_16718,N_16410,N_16014);
nand U16719 (N_16719,N_16449,N_16148);
xor U16720 (N_16720,N_16025,N_16068);
or U16721 (N_16721,N_16203,N_16214);
nand U16722 (N_16722,N_16375,N_16219);
nand U16723 (N_16723,N_16101,N_16132);
nand U16724 (N_16724,N_16103,N_16218);
or U16725 (N_16725,N_16471,N_16208);
xor U16726 (N_16726,N_16415,N_16180);
or U16727 (N_16727,N_16153,N_16307);
and U16728 (N_16728,N_16197,N_16035);
xnor U16729 (N_16729,N_16249,N_16162);
and U16730 (N_16730,N_16144,N_16496);
nor U16731 (N_16731,N_16287,N_16333);
nand U16732 (N_16732,N_16487,N_16295);
and U16733 (N_16733,N_16405,N_16202);
nor U16734 (N_16734,N_16150,N_16301);
nor U16735 (N_16735,N_16098,N_16054);
nor U16736 (N_16736,N_16081,N_16495);
and U16737 (N_16737,N_16200,N_16329);
nand U16738 (N_16738,N_16338,N_16422);
and U16739 (N_16739,N_16378,N_16443);
or U16740 (N_16740,N_16359,N_16273);
and U16741 (N_16741,N_16413,N_16174);
or U16742 (N_16742,N_16326,N_16381);
nor U16743 (N_16743,N_16493,N_16009);
xnor U16744 (N_16744,N_16119,N_16432);
and U16745 (N_16745,N_16136,N_16205);
nor U16746 (N_16746,N_16138,N_16166);
or U16747 (N_16747,N_16462,N_16222);
or U16748 (N_16748,N_16269,N_16309);
xor U16749 (N_16749,N_16064,N_16006);
xnor U16750 (N_16750,N_16336,N_16484);
nor U16751 (N_16751,N_16194,N_16339);
or U16752 (N_16752,N_16361,N_16259);
nor U16753 (N_16753,N_16254,N_16316);
or U16754 (N_16754,N_16163,N_16478);
nor U16755 (N_16755,N_16322,N_16245);
xor U16756 (N_16756,N_16160,N_16493);
nor U16757 (N_16757,N_16125,N_16132);
or U16758 (N_16758,N_16391,N_16435);
and U16759 (N_16759,N_16425,N_16002);
nor U16760 (N_16760,N_16193,N_16248);
and U16761 (N_16761,N_16263,N_16049);
and U16762 (N_16762,N_16159,N_16459);
nor U16763 (N_16763,N_16189,N_16418);
nand U16764 (N_16764,N_16326,N_16289);
nor U16765 (N_16765,N_16381,N_16323);
nand U16766 (N_16766,N_16323,N_16396);
and U16767 (N_16767,N_16090,N_16168);
nor U16768 (N_16768,N_16452,N_16098);
nor U16769 (N_16769,N_16269,N_16346);
and U16770 (N_16770,N_16120,N_16367);
or U16771 (N_16771,N_16230,N_16063);
nor U16772 (N_16772,N_16355,N_16324);
xor U16773 (N_16773,N_16111,N_16054);
nor U16774 (N_16774,N_16243,N_16252);
nand U16775 (N_16775,N_16103,N_16475);
or U16776 (N_16776,N_16238,N_16428);
and U16777 (N_16777,N_16420,N_16352);
or U16778 (N_16778,N_16396,N_16184);
or U16779 (N_16779,N_16399,N_16165);
or U16780 (N_16780,N_16079,N_16167);
nand U16781 (N_16781,N_16355,N_16466);
nand U16782 (N_16782,N_16467,N_16257);
nor U16783 (N_16783,N_16351,N_16141);
nor U16784 (N_16784,N_16495,N_16241);
nor U16785 (N_16785,N_16313,N_16403);
nand U16786 (N_16786,N_16165,N_16030);
and U16787 (N_16787,N_16028,N_16337);
nand U16788 (N_16788,N_16294,N_16104);
xnor U16789 (N_16789,N_16364,N_16427);
nor U16790 (N_16790,N_16093,N_16386);
nand U16791 (N_16791,N_16084,N_16263);
and U16792 (N_16792,N_16216,N_16382);
nor U16793 (N_16793,N_16498,N_16467);
and U16794 (N_16794,N_16474,N_16391);
and U16795 (N_16795,N_16159,N_16363);
nor U16796 (N_16796,N_16177,N_16333);
or U16797 (N_16797,N_16415,N_16174);
xor U16798 (N_16798,N_16471,N_16265);
xor U16799 (N_16799,N_16324,N_16201);
nor U16800 (N_16800,N_16308,N_16373);
or U16801 (N_16801,N_16002,N_16433);
and U16802 (N_16802,N_16060,N_16479);
nand U16803 (N_16803,N_16367,N_16119);
nand U16804 (N_16804,N_16477,N_16152);
nor U16805 (N_16805,N_16050,N_16012);
and U16806 (N_16806,N_16314,N_16207);
xnor U16807 (N_16807,N_16101,N_16368);
xor U16808 (N_16808,N_16197,N_16338);
and U16809 (N_16809,N_16330,N_16022);
xor U16810 (N_16810,N_16463,N_16366);
nor U16811 (N_16811,N_16244,N_16320);
nand U16812 (N_16812,N_16089,N_16199);
nand U16813 (N_16813,N_16382,N_16184);
xnor U16814 (N_16814,N_16282,N_16098);
and U16815 (N_16815,N_16387,N_16020);
nor U16816 (N_16816,N_16487,N_16441);
nand U16817 (N_16817,N_16249,N_16150);
and U16818 (N_16818,N_16031,N_16293);
or U16819 (N_16819,N_16249,N_16052);
or U16820 (N_16820,N_16493,N_16247);
and U16821 (N_16821,N_16095,N_16259);
xnor U16822 (N_16822,N_16011,N_16364);
nand U16823 (N_16823,N_16178,N_16314);
xnor U16824 (N_16824,N_16078,N_16420);
nand U16825 (N_16825,N_16023,N_16367);
and U16826 (N_16826,N_16084,N_16301);
or U16827 (N_16827,N_16044,N_16357);
nor U16828 (N_16828,N_16343,N_16443);
and U16829 (N_16829,N_16039,N_16340);
nand U16830 (N_16830,N_16272,N_16229);
or U16831 (N_16831,N_16410,N_16163);
or U16832 (N_16832,N_16335,N_16443);
or U16833 (N_16833,N_16313,N_16142);
and U16834 (N_16834,N_16304,N_16126);
xnor U16835 (N_16835,N_16032,N_16316);
and U16836 (N_16836,N_16388,N_16288);
nor U16837 (N_16837,N_16219,N_16162);
nor U16838 (N_16838,N_16146,N_16280);
nand U16839 (N_16839,N_16117,N_16027);
or U16840 (N_16840,N_16285,N_16021);
xor U16841 (N_16841,N_16392,N_16300);
and U16842 (N_16842,N_16324,N_16428);
xnor U16843 (N_16843,N_16432,N_16349);
and U16844 (N_16844,N_16138,N_16357);
xnor U16845 (N_16845,N_16304,N_16082);
xnor U16846 (N_16846,N_16476,N_16473);
nand U16847 (N_16847,N_16458,N_16346);
nor U16848 (N_16848,N_16384,N_16329);
xnor U16849 (N_16849,N_16421,N_16127);
xnor U16850 (N_16850,N_16391,N_16422);
nor U16851 (N_16851,N_16400,N_16423);
nor U16852 (N_16852,N_16216,N_16399);
xnor U16853 (N_16853,N_16232,N_16188);
nor U16854 (N_16854,N_16472,N_16376);
nand U16855 (N_16855,N_16247,N_16034);
nand U16856 (N_16856,N_16320,N_16043);
xor U16857 (N_16857,N_16141,N_16022);
or U16858 (N_16858,N_16304,N_16315);
nor U16859 (N_16859,N_16172,N_16084);
and U16860 (N_16860,N_16280,N_16219);
nand U16861 (N_16861,N_16321,N_16391);
nand U16862 (N_16862,N_16411,N_16072);
xor U16863 (N_16863,N_16150,N_16115);
xnor U16864 (N_16864,N_16228,N_16294);
or U16865 (N_16865,N_16461,N_16265);
or U16866 (N_16866,N_16191,N_16140);
and U16867 (N_16867,N_16460,N_16390);
nor U16868 (N_16868,N_16130,N_16393);
xnor U16869 (N_16869,N_16125,N_16105);
or U16870 (N_16870,N_16020,N_16422);
xnor U16871 (N_16871,N_16019,N_16391);
and U16872 (N_16872,N_16496,N_16364);
nor U16873 (N_16873,N_16454,N_16195);
or U16874 (N_16874,N_16331,N_16306);
nand U16875 (N_16875,N_16357,N_16079);
or U16876 (N_16876,N_16271,N_16080);
or U16877 (N_16877,N_16348,N_16030);
xnor U16878 (N_16878,N_16001,N_16073);
and U16879 (N_16879,N_16098,N_16334);
xor U16880 (N_16880,N_16163,N_16160);
nand U16881 (N_16881,N_16464,N_16237);
nor U16882 (N_16882,N_16184,N_16062);
or U16883 (N_16883,N_16469,N_16208);
nand U16884 (N_16884,N_16018,N_16072);
or U16885 (N_16885,N_16329,N_16210);
nand U16886 (N_16886,N_16441,N_16340);
nand U16887 (N_16887,N_16303,N_16352);
nor U16888 (N_16888,N_16445,N_16494);
nand U16889 (N_16889,N_16418,N_16169);
or U16890 (N_16890,N_16258,N_16050);
and U16891 (N_16891,N_16315,N_16055);
or U16892 (N_16892,N_16231,N_16446);
and U16893 (N_16893,N_16217,N_16446);
or U16894 (N_16894,N_16492,N_16441);
xnor U16895 (N_16895,N_16271,N_16083);
or U16896 (N_16896,N_16491,N_16471);
xor U16897 (N_16897,N_16034,N_16302);
xnor U16898 (N_16898,N_16404,N_16035);
xnor U16899 (N_16899,N_16391,N_16044);
nor U16900 (N_16900,N_16215,N_16240);
or U16901 (N_16901,N_16173,N_16062);
xnor U16902 (N_16902,N_16101,N_16112);
nor U16903 (N_16903,N_16160,N_16183);
nor U16904 (N_16904,N_16049,N_16092);
and U16905 (N_16905,N_16073,N_16359);
nor U16906 (N_16906,N_16414,N_16149);
and U16907 (N_16907,N_16188,N_16313);
or U16908 (N_16908,N_16267,N_16283);
nor U16909 (N_16909,N_16492,N_16309);
nor U16910 (N_16910,N_16217,N_16214);
or U16911 (N_16911,N_16327,N_16134);
nor U16912 (N_16912,N_16286,N_16118);
xnor U16913 (N_16913,N_16251,N_16443);
and U16914 (N_16914,N_16141,N_16232);
or U16915 (N_16915,N_16172,N_16116);
and U16916 (N_16916,N_16012,N_16321);
or U16917 (N_16917,N_16494,N_16055);
xnor U16918 (N_16918,N_16444,N_16187);
nor U16919 (N_16919,N_16175,N_16245);
nor U16920 (N_16920,N_16055,N_16246);
or U16921 (N_16921,N_16493,N_16399);
nand U16922 (N_16922,N_16187,N_16300);
nor U16923 (N_16923,N_16458,N_16197);
nor U16924 (N_16924,N_16311,N_16144);
nand U16925 (N_16925,N_16445,N_16113);
nand U16926 (N_16926,N_16368,N_16416);
xnor U16927 (N_16927,N_16023,N_16473);
or U16928 (N_16928,N_16103,N_16284);
and U16929 (N_16929,N_16277,N_16065);
xor U16930 (N_16930,N_16008,N_16429);
and U16931 (N_16931,N_16435,N_16036);
xor U16932 (N_16932,N_16069,N_16411);
nand U16933 (N_16933,N_16453,N_16339);
xnor U16934 (N_16934,N_16426,N_16212);
xnor U16935 (N_16935,N_16416,N_16335);
xor U16936 (N_16936,N_16152,N_16473);
nor U16937 (N_16937,N_16226,N_16068);
nand U16938 (N_16938,N_16039,N_16129);
and U16939 (N_16939,N_16283,N_16309);
nand U16940 (N_16940,N_16280,N_16490);
or U16941 (N_16941,N_16231,N_16034);
nand U16942 (N_16942,N_16450,N_16171);
xnor U16943 (N_16943,N_16362,N_16070);
nor U16944 (N_16944,N_16112,N_16073);
nand U16945 (N_16945,N_16316,N_16356);
or U16946 (N_16946,N_16308,N_16470);
xor U16947 (N_16947,N_16095,N_16017);
nor U16948 (N_16948,N_16032,N_16039);
and U16949 (N_16949,N_16146,N_16036);
and U16950 (N_16950,N_16233,N_16433);
and U16951 (N_16951,N_16411,N_16071);
nand U16952 (N_16952,N_16221,N_16266);
nor U16953 (N_16953,N_16261,N_16220);
xnor U16954 (N_16954,N_16286,N_16379);
nand U16955 (N_16955,N_16124,N_16317);
and U16956 (N_16956,N_16115,N_16222);
and U16957 (N_16957,N_16437,N_16312);
and U16958 (N_16958,N_16174,N_16143);
or U16959 (N_16959,N_16426,N_16320);
nand U16960 (N_16960,N_16147,N_16348);
or U16961 (N_16961,N_16231,N_16398);
and U16962 (N_16962,N_16183,N_16298);
or U16963 (N_16963,N_16091,N_16035);
or U16964 (N_16964,N_16230,N_16237);
xor U16965 (N_16965,N_16427,N_16151);
nand U16966 (N_16966,N_16437,N_16220);
and U16967 (N_16967,N_16419,N_16306);
or U16968 (N_16968,N_16351,N_16225);
nand U16969 (N_16969,N_16467,N_16225);
nand U16970 (N_16970,N_16258,N_16407);
nor U16971 (N_16971,N_16236,N_16131);
nand U16972 (N_16972,N_16095,N_16153);
nor U16973 (N_16973,N_16260,N_16179);
nand U16974 (N_16974,N_16045,N_16158);
and U16975 (N_16975,N_16442,N_16274);
nand U16976 (N_16976,N_16015,N_16231);
xor U16977 (N_16977,N_16423,N_16438);
or U16978 (N_16978,N_16199,N_16300);
nand U16979 (N_16979,N_16405,N_16476);
and U16980 (N_16980,N_16128,N_16267);
nand U16981 (N_16981,N_16335,N_16434);
nor U16982 (N_16982,N_16252,N_16155);
xor U16983 (N_16983,N_16017,N_16228);
or U16984 (N_16984,N_16272,N_16387);
nand U16985 (N_16985,N_16365,N_16421);
and U16986 (N_16986,N_16418,N_16322);
nor U16987 (N_16987,N_16307,N_16273);
or U16988 (N_16988,N_16443,N_16286);
xnor U16989 (N_16989,N_16176,N_16243);
xnor U16990 (N_16990,N_16156,N_16104);
xnor U16991 (N_16991,N_16337,N_16209);
nand U16992 (N_16992,N_16009,N_16020);
nand U16993 (N_16993,N_16254,N_16383);
nand U16994 (N_16994,N_16094,N_16286);
nand U16995 (N_16995,N_16408,N_16021);
or U16996 (N_16996,N_16402,N_16030);
nand U16997 (N_16997,N_16446,N_16031);
or U16998 (N_16998,N_16366,N_16259);
xor U16999 (N_16999,N_16206,N_16401);
nor U17000 (N_17000,N_16650,N_16772);
xor U17001 (N_17001,N_16985,N_16717);
or U17002 (N_17002,N_16852,N_16581);
and U17003 (N_17003,N_16600,N_16590);
nand U17004 (N_17004,N_16915,N_16745);
and U17005 (N_17005,N_16758,N_16707);
nor U17006 (N_17006,N_16769,N_16813);
and U17007 (N_17007,N_16934,N_16766);
nand U17008 (N_17008,N_16843,N_16604);
or U17009 (N_17009,N_16674,N_16797);
or U17010 (N_17010,N_16595,N_16950);
nand U17011 (N_17011,N_16690,N_16853);
nand U17012 (N_17012,N_16618,N_16641);
nor U17013 (N_17013,N_16735,N_16592);
xnor U17014 (N_17014,N_16856,N_16685);
xor U17015 (N_17015,N_16507,N_16622);
nor U17016 (N_17016,N_16890,N_16996);
xor U17017 (N_17017,N_16871,N_16623);
and U17018 (N_17018,N_16504,N_16887);
xor U17019 (N_17019,N_16921,N_16886);
or U17020 (N_17020,N_16543,N_16978);
or U17021 (N_17021,N_16913,N_16651);
or U17022 (N_17022,N_16806,N_16998);
nor U17023 (N_17023,N_16607,N_16520);
or U17024 (N_17024,N_16937,N_16644);
nor U17025 (N_17025,N_16855,N_16633);
nand U17026 (N_17026,N_16624,N_16694);
xor U17027 (N_17027,N_16764,N_16566);
or U17028 (N_17028,N_16736,N_16837);
xor U17029 (N_17029,N_16829,N_16796);
or U17030 (N_17030,N_16879,N_16561);
nand U17031 (N_17031,N_16669,N_16961);
and U17032 (N_17032,N_16818,N_16602);
nand U17033 (N_17033,N_16596,N_16778);
and U17034 (N_17034,N_16626,N_16771);
or U17035 (N_17035,N_16662,N_16822);
nor U17036 (N_17036,N_16611,N_16916);
nor U17037 (N_17037,N_16597,N_16671);
nor U17038 (N_17038,N_16866,N_16820);
nor U17039 (N_17039,N_16533,N_16817);
or U17040 (N_17040,N_16683,N_16609);
or U17041 (N_17041,N_16749,N_16876);
xnor U17042 (N_17042,N_16786,N_16975);
or U17043 (N_17043,N_16713,N_16724);
and U17044 (N_17044,N_16734,N_16579);
nor U17045 (N_17045,N_16750,N_16727);
xnor U17046 (N_17046,N_16576,N_16708);
or U17047 (N_17047,N_16560,N_16909);
nand U17048 (N_17048,N_16687,N_16722);
nor U17049 (N_17049,N_16785,N_16941);
or U17050 (N_17050,N_16914,N_16911);
nand U17051 (N_17051,N_16833,N_16804);
xor U17052 (N_17052,N_16842,N_16865);
nand U17053 (N_17053,N_16582,N_16574);
and U17054 (N_17054,N_16621,N_16518);
or U17055 (N_17055,N_16688,N_16858);
xnor U17056 (N_17056,N_16591,N_16794);
nor U17057 (N_17057,N_16986,N_16827);
xor U17058 (N_17058,N_16728,N_16629);
xor U17059 (N_17059,N_16739,N_16679);
xnor U17060 (N_17060,N_16552,N_16619);
or U17061 (N_17061,N_16698,N_16841);
xnor U17062 (N_17062,N_16712,N_16555);
or U17063 (N_17063,N_16828,N_16652);
and U17064 (N_17064,N_16696,N_16680);
xnor U17065 (N_17065,N_16558,N_16725);
nand U17066 (N_17066,N_16899,N_16925);
nor U17067 (N_17067,N_16747,N_16895);
nor U17068 (N_17068,N_16705,N_16968);
nand U17069 (N_17069,N_16516,N_16744);
xor U17070 (N_17070,N_16657,N_16862);
xor U17071 (N_17071,N_16501,N_16891);
or U17072 (N_17072,N_16616,N_16535);
nand U17073 (N_17073,N_16798,N_16594);
nor U17074 (N_17074,N_16663,N_16952);
nor U17075 (N_17075,N_16664,N_16919);
xor U17076 (N_17076,N_16539,N_16906);
nor U17077 (N_17077,N_16885,N_16900);
xor U17078 (N_17078,N_16716,N_16718);
and U17079 (N_17079,N_16640,N_16880);
or U17080 (N_17080,N_16759,N_16816);
or U17081 (N_17081,N_16765,N_16661);
and U17082 (N_17082,N_16704,N_16636);
and U17083 (N_17083,N_16940,N_16848);
or U17084 (N_17084,N_16810,N_16695);
nor U17085 (N_17085,N_16601,N_16684);
and U17086 (N_17086,N_16763,N_16991);
xor U17087 (N_17087,N_16976,N_16930);
or U17088 (N_17088,N_16614,N_16999);
and U17089 (N_17089,N_16922,N_16805);
nand U17090 (N_17090,N_16973,N_16628);
xnor U17091 (N_17091,N_16655,N_16874);
xnor U17092 (N_17092,N_16956,N_16953);
or U17093 (N_17093,N_16997,N_16568);
or U17094 (N_17094,N_16748,N_16839);
and U17095 (N_17095,N_16846,N_16572);
and U17096 (N_17096,N_16859,N_16672);
and U17097 (N_17097,N_16559,N_16892);
xnor U17098 (N_17098,N_16894,N_16944);
nand U17099 (N_17099,N_16746,N_16788);
nor U17100 (N_17100,N_16742,N_16795);
nor U17101 (N_17101,N_16924,N_16993);
xnor U17102 (N_17102,N_16923,N_16957);
nand U17103 (N_17103,N_16815,N_16814);
nor U17104 (N_17104,N_16770,N_16675);
xnor U17105 (N_17105,N_16525,N_16834);
xor U17106 (N_17106,N_16710,N_16936);
and U17107 (N_17107,N_16992,N_16645);
or U17108 (N_17108,N_16942,N_16711);
nand U17109 (N_17109,N_16738,N_16955);
nand U17110 (N_17110,N_16638,N_16912);
nor U17111 (N_17111,N_16665,N_16586);
nand U17112 (N_17112,N_16939,N_16612);
nand U17113 (N_17113,N_16835,N_16541);
or U17114 (N_17114,N_16562,N_16929);
nand U17115 (N_17115,N_16830,N_16974);
or U17116 (N_17116,N_16699,N_16500);
and U17117 (N_17117,N_16966,N_16656);
nor U17118 (N_17118,N_16723,N_16731);
nor U17119 (N_17119,N_16868,N_16808);
and U17120 (N_17120,N_16767,N_16511);
nor U17121 (N_17121,N_16536,N_16864);
and U17122 (N_17122,N_16838,N_16754);
and U17123 (N_17123,N_16701,N_16989);
nor U17124 (N_17124,N_16753,N_16775);
nand U17125 (N_17125,N_16983,N_16793);
nor U17126 (N_17126,N_16954,N_16948);
nor U17127 (N_17127,N_16585,N_16519);
and U17128 (N_17128,N_16643,N_16733);
xnor U17129 (N_17129,N_16803,N_16857);
xnor U17130 (N_17130,N_16823,N_16888);
xor U17131 (N_17131,N_16969,N_16740);
or U17132 (N_17132,N_16583,N_16920);
xor U17133 (N_17133,N_16938,N_16529);
nand U17134 (N_17134,N_16964,N_16980);
or U17135 (N_17135,N_16777,N_16762);
and U17136 (N_17136,N_16606,N_16781);
or U17137 (N_17137,N_16654,N_16902);
nand U17138 (N_17138,N_16821,N_16608);
nand U17139 (N_17139,N_16811,N_16570);
nand U17140 (N_17140,N_16826,N_16792);
xnor U17141 (N_17141,N_16673,N_16951);
nand U17142 (N_17142,N_16901,N_16538);
xor U17143 (N_17143,N_16931,N_16615);
nor U17144 (N_17144,N_16984,N_16860);
or U17145 (N_17145,N_16741,N_16668);
nor U17146 (N_17146,N_16598,N_16553);
nor U17147 (N_17147,N_16667,N_16577);
and U17148 (N_17148,N_16521,N_16564);
or U17149 (N_17149,N_16587,N_16620);
and U17150 (N_17150,N_16971,N_16927);
nand U17151 (N_17151,N_16875,N_16653);
nor U17152 (N_17152,N_16702,N_16557);
or U17153 (N_17153,N_16720,N_16540);
xnor U17154 (N_17154,N_16751,N_16505);
nor U17155 (N_17155,N_16584,N_16715);
or U17156 (N_17156,N_16905,N_16844);
nor U17157 (N_17157,N_16571,N_16897);
and U17158 (N_17158,N_16565,N_16773);
nand U17159 (N_17159,N_16768,N_16760);
nand U17160 (N_17160,N_16824,N_16659);
xnor U17161 (N_17161,N_16569,N_16873);
nor U17162 (N_17162,N_16898,N_16515);
nand U17163 (N_17163,N_16646,N_16779);
or U17164 (N_17164,N_16782,N_16756);
and U17165 (N_17165,N_16706,N_16677);
or U17166 (N_17166,N_16700,N_16580);
and U17167 (N_17167,N_16981,N_16863);
or U17168 (N_17168,N_16726,N_16851);
xor U17169 (N_17169,N_16691,N_16554);
or U17170 (N_17170,N_16836,N_16647);
or U17171 (N_17171,N_16528,N_16926);
nor U17172 (N_17172,N_16512,N_16681);
nand U17173 (N_17173,N_16903,N_16630);
or U17174 (N_17174,N_16861,N_16625);
or U17175 (N_17175,N_16575,N_16589);
nand U17176 (N_17176,N_16648,N_16730);
or U17177 (N_17177,N_16972,N_16634);
nor U17178 (N_17178,N_16752,N_16506);
nor U17179 (N_17179,N_16849,N_16884);
or U17180 (N_17180,N_16660,N_16508);
nor U17181 (N_17181,N_16599,N_16721);
or U17182 (N_17182,N_16831,N_16578);
nor U17183 (N_17183,N_16544,N_16550);
nand U17184 (N_17184,N_16531,N_16603);
xor U17185 (N_17185,N_16547,N_16947);
and U17186 (N_17186,N_16801,N_16960);
nor U17187 (N_17187,N_16588,N_16542);
and U17188 (N_17188,N_16867,N_16686);
or U17189 (N_17189,N_16605,N_16845);
xnor U17190 (N_17190,N_16503,N_16932);
xnor U17191 (N_17191,N_16963,N_16878);
and U17192 (N_17192,N_16697,N_16563);
and U17193 (N_17193,N_16613,N_16593);
nand U17194 (N_17194,N_16994,N_16908);
and U17195 (N_17195,N_16784,N_16949);
xor U17196 (N_17196,N_16502,N_16524);
xor U17197 (N_17197,N_16757,N_16990);
nand U17198 (N_17198,N_16791,N_16877);
nor U17199 (N_17199,N_16967,N_16910);
nand U17200 (N_17200,N_16802,N_16825);
and U17201 (N_17201,N_16549,N_16666);
nor U17202 (N_17202,N_16907,N_16807);
or U17203 (N_17203,N_16776,N_16869);
and U17204 (N_17204,N_16573,N_16928);
or U17205 (N_17205,N_16979,N_16918);
xnor U17206 (N_17206,N_16882,N_16787);
nand U17207 (N_17207,N_16790,N_16780);
nor U17208 (N_17208,N_16635,N_16904);
or U17209 (N_17209,N_16832,N_16556);
xnor U17210 (N_17210,N_16761,N_16523);
or U17211 (N_17211,N_16649,N_16774);
or U17212 (N_17212,N_16509,N_16658);
nor U17213 (N_17213,N_16893,N_16854);
or U17214 (N_17214,N_16514,N_16678);
or U17215 (N_17215,N_16642,N_16935);
or U17216 (N_17216,N_16783,N_16917);
xnor U17217 (N_17217,N_16639,N_16800);
and U17218 (N_17218,N_16933,N_16537);
or U17219 (N_17219,N_16840,N_16789);
nor U17220 (N_17220,N_16870,N_16982);
nand U17221 (N_17221,N_16551,N_16977);
nand U17222 (N_17222,N_16627,N_16676);
or U17223 (N_17223,N_16513,N_16719);
or U17224 (N_17224,N_16703,N_16965);
and U17225 (N_17225,N_16510,N_16812);
nor U17226 (N_17226,N_16799,N_16872);
nand U17227 (N_17227,N_16958,N_16945);
or U17228 (N_17228,N_16545,N_16962);
xnor U17229 (N_17229,N_16743,N_16526);
nor U17230 (N_17230,N_16546,N_16732);
nor U17231 (N_17231,N_16617,N_16567);
and U17232 (N_17232,N_16548,N_16995);
and U17233 (N_17233,N_16522,N_16714);
or U17234 (N_17234,N_16959,N_16632);
nand U17235 (N_17235,N_16883,N_16970);
xor U17236 (N_17236,N_16847,N_16850);
or U17237 (N_17237,N_16946,N_16943);
nand U17238 (N_17238,N_16729,N_16527);
or U17239 (N_17239,N_16530,N_16682);
or U17240 (N_17240,N_16889,N_16693);
xor U17241 (N_17241,N_16737,N_16637);
and U17242 (N_17242,N_16692,N_16987);
xnor U17243 (N_17243,N_16709,N_16631);
nor U17244 (N_17244,N_16819,N_16517);
or U17245 (N_17245,N_16755,N_16988);
nor U17246 (N_17246,N_16534,N_16610);
xor U17247 (N_17247,N_16670,N_16896);
nand U17248 (N_17248,N_16689,N_16532);
and U17249 (N_17249,N_16809,N_16881);
or U17250 (N_17250,N_16733,N_16648);
xnor U17251 (N_17251,N_16855,N_16689);
nand U17252 (N_17252,N_16976,N_16601);
and U17253 (N_17253,N_16781,N_16549);
and U17254 (N_17254,N_16868,N_16988);
nand U17255 (N_17255,N_16549,N_16718);
nand U17256 (N_17256,N_16696,N_16973);
nor U17257 (N_17257,N_16741,N_16930);
nand U17258 (N_17258,N_16588,N_16722);
nand U17259 (N_17259,N_16506,N_16992);
nand U17260 (N_17260,N_16666,N_16803);
or U17261 (N_17261,N_16812,N_16737);
nand U17262 (N_17262,N_16623,N_16539);
xor U17263 (N_17263,N_16641,N_16905);
nand U17264 (N_17264,N_16572,N_16586);
or U17265 (N_17265,N_16627,N_16784);
nor U17266 (N_17266,N_16734,N_16624);
xnor U17267 (N_17267,N_16915,N_16514);
xor U17268 (N_17268,N_16619,N_16729);
and U17269 (N_17269,N_16889,N_16773);
and U17270 (N_17270,N_16554,N_16908);
xor U17271 (N_17271,N_16642,N_16836);
xnor U17272 (N_17272,N_16977,N_16905);
or U17273 (N_17273,N_16977,N_16658);
xnor U17274 (N_17274,N_16943,N_16982);
nand U17275 (N_17275,N_16791,N_16766);
or U17276 (N_17276,N_16619,N_16800);
and U17277 (N_17277,N_16616,N_16860);
and U17278 (N_17278,N_16948,N_16500);
nand U17279 (N_17279,N_16586,N_16727);
or U17280 (N_17280,N_16643,N_16645);
nand U17281 (N_17281,N_16946,N_16978);
and U17282 (N_17282,N_16929,N_16588);
nor U17283 (N_17283,N_16721,N_16546);
and U17284 (N_17284,N_16559,N_16824);
nor U17285 (N_17285,N_16899,N_16926);
nand U17286 (N_17286,N_16543,N_16518);
nor U17287 (N_17287,N_16573,N_16821);
xor U17288 (N_17288,N_16895,N_16626);
xor U17289 (N_17289,N_16738,N_16765);
nand U17290 (N_17290,N_16681,N_16854);
or U17291 (N_17291,N_16738,N_16932);
and U17292 (N_17292,N_16628,N_16805);
and U17293 (N_17293,N_16507,N_16569);
xnor U17294 (N_17294,N_16840,N_16992);
xor U17295 (N_17295,N_16544,N_16827);
nand U17296 (N_17296,N_16760,N_16836);
and U17297 (N_17297,N_16529,N_16809);
and U17298 (N_17298,N_16916,N_16507);
xor U17299 (N_17299,N_16631,N_16759);
and U17300 (N_17300,N_16708,N_16772);
or U17301 (N_17301,N_16935,N_16663);
and U17302 (N_17302,N_16541,N_16846);
nor U17303 (N_17303,N_16951,N_16731);
or U17304 (N_17304,N_16618,N_16823);
nor U17305 (N_17305,N_16683,N_16679);
xor U17306 (N_17306,N_16951,N_16662);
nand U17307 (N_17307,N_16706,N_16536);
xor U17308 (N_17308,N_16832,N_16836);
nand U17309 (N_17309,N_16793,N_16992);
nand U17310 (N_17310,N_16686,N_16926);
and U17311 (N_17311,N_16907,N_16696);
nand U17312 (N_17312,N_16820,N_16914);
and U17313 (N_17313,N_16942,N_16655);
nor U17314 (N_17314,N_16623,N_16683);
nor U17315 (N_17315,N_16999,N_16567);
and U17316 (N_17316,N_16656,N_16877);
xnor U17317 (N_17317,N_16725,N_16862);
nand U17318 (N_17318,N_16505,N_16877);
and U17319 (N_17319,N_16850,N_16574);
or U17320 (N_17320,N_16891,N_16857);
or U17321 (N_17321,N_16861,N_16754);
nor U17322 (N_17322,N_16955,N_16627);
or U17323 (N_17323,N_16654,N_16799);
nor U17324 (N_17324,N_16847,N_16945);
or U17325 (N_17325,N_16977,N_16848);
nor U17326 (N_17326,N_16526,N_16895);
or U17327 (N_17327,N_16598,N_16946);
xor U17328 (N_17328,N_16922,N_16568);
and U17329 (N_17329,N_16939,N_16586);
nand U17330 (N_17330,N_16690,N_16657);
xor U17331 (N_17331,N_16569,N_16742);
nand U17332 (N_17332,N_16805,N_16595);
nand U17333 (N_17333,N_16590,N_16706);
xnor U17334 (N_17334,N_16547,N_16741);
xor U17335 (N_17335,N_16990,N_16508);
nand U17336 (N_17336,N_16679,N_16673);
and U17337 (N_17337,N_16535,N_16782);
or U17338 (N_17338,N_16812,N_16649);
nand U17339 (N_17339,N_16707,N_16692);
xor U17340 (N_17340,N_16576,N_16614);
xnor U17341 (N_17341,N_16793,N_16525);
nor U17342 (N_17342,N_16542,N_16702);
nor U17343 (N_17343,N_16584,N_16578);
nor U17344 (N_17344,N_16768,N_16830);
or U17345 (N_17345,N_16874,N_16983);
or U17346 (N_17346,N_16972,N_16843);
xnor U17347 (N_17347,N_16549,N_16559);
or U17348 (N_17348,N_16848,N_16660);
xor U17349 (N_17349,N_16902,N_16813);
or U17350 (N_17350,N_16764,N_16877);
and U17351 (N_17351,N_16629,N_16661);
and U17352 (N_17352,N_16900,N_16652);
xnor U17353 (N_17353,N_16964,N_16601);
nor U17354 (N_17354,N_16505,N_16532);
nor U17355 (N_17355,N_16596,N_16786);
nand U17356 (N_17356,N_16781,N_16556);
and U17357 (N_17357,N_16997,N_16966);
xnor U17358 (N_17358,N_16562,N_16593);
and U17359 (N_17359,N_16670,N_16846);
nor U17360 (N_17360,N_16783,N_16940);
or U17361 (N_17361,N_16504,N_16711);
xnor U17362 (N_17362,N_16928,N_16720);
or U17363 (N_17363,N_16531,N_16643);
xor U17364 (N_17364,N_16520,N_16537);
nand U17365 (N_17365,N_16638,N_16959);
nand U17366 (N_17366,N_16585,N_16923);
or U17367 (N_17367,N_16684,N_16513);
xnor U17368 (N_17368,N_16551,N_16532);
or U17369 (N_17369,N_16566,N_16511);
and U17370 (N_17370,N_16705,N_16668);
nor U17371 (N_17371,N_16506,N_16583);
or U17372 (N_17372,N_16810,N_16864);
nor U17373 (N_17373,N_16686,N_16551);
nand U17374 (N_17374,N_16874,N_16867);
and U17375 (N_17375,N_16997,N_16653);
nor U17376 (N_17376,N_16921,N_16920);
and U17377 (N_17377,N_16760,N_16667);
nor U17378 (N_17378,N_16551,N_16660);
nor U17379 (N_17379,N_16660,N_16838);
nor U17380 (N_17380,N_16880,N_16819);
or U17381 (N_17381,N_16529,N_16796);
xor U17382 (N_17382,N_16948,N_16598);
and U17383 (N_17383,N_16783,N_16792);
nor U17384 (N_17384,N_16772,N_16743);
nand U17385 (N_17385,N_16569,N_16805);
xnor U17386 (N_17386,N_16764,N_16571);
nand U17387 (N_17387,N_16689,N_16794);
and U17388 (N_17388,N_16855,N_16557);
or U17389 (N_17389,N_16867,N_16653);
nand U17390 (N_17390,N_16988,N_16689);
or U17391 (N_17391,N_16878,N_16803);
and U17392 (N_17392,N_16547,N_16906);
nand U17393 (N_17393,N_16526,N_16614);
or U17394 (N_17394,N_16910,N_16868);
nor U17395 (N_17395,N_16648,N_16928);
xor U17396 (N_17396,N_16999,N_16743);
nor U17397 (N_17397,N_16575,N_16857);
and U17398 (N_17398,N_16779,N_16969);
xnor U17399 (N_17399,N_16874,N_16858);
nand U17400 (N_17400,N_16782,N_16613);
or U17401 (N_17401,N_16997,N_16550);
xnor U17402 (N_17402,N_16682,N_16689);
and U17403 (N_17403,N_16788,N_16511);
xor U17404 (N_17404,N_16833,N_16656);
or U17405 (N_17405,N_16542,N_16824);
and U17406 (N_17406,N_16958,N_16778);
or U17407 (N_17407,N_16622,N_16749);
and U17408 (N_17408,N_16523,N_16705);
nor U17409 (N_17409,N_16500,N_16732);
xnor U17410 (N_17410,N_16750,N_16557);
or U17411 (N_17411,N_16719,N_16635);
nand U17412 (N_17412,N_16694,N_16680);
or U17413 (N_17413,N_16972,N_16606);
and U17414 (N_17414,N_16904,N_16851);
xnor U17415 (N_17415,N_16626,N_16711);
and U17416 (N_17416,N_16857,N_16812);
or U17417 (N_17417,N_16672,N_16544);
and U17418 (N_17418,N_16792,N_16837);
and U17419 (N_17419,N_16731,N_16847);
or U17420 (N_17420,N_16838,N_16533);
and U17421 (N_17421,N_16608,N_16873);
xnor U17422 (N_17422,N_16612,N_16960);
and U17423 (N_17423,N_16858,N_16775);
or U17424 (N_17424,N_16917,N_16668);
xnor U17425 (N_17425,N_16866,N_16882);
nor U17426 (N_17426,N_16783,N_16741);
and U17427 (N_17427,N_16861,N_16935);
and U17428 (N_17428,N_16687,N_16616);
xor U17429 (N_17429,N_16608,N_16532);
xnor U17430 (N_17430,N_16591,N_16888);
or U17431 (N_17431,N_16931,N_16908);
nand U17432 (N_17432,N_16832,N_16727);
nor U17433 (N_17433,N_16594,N_16926);
nor U17434 (N_17434,N_16722,N_16523);
nand U17435 (N_17435,N_16930,N_16880);
nor U17436 (N_17436,N_16788,N_16672);
and U17437 (N_17437,N_16559,N_16952);
or U17438 (N_17438,N_16575,N_16867);
or U17439 (N_17439,N_16750,N_16931);
xnor U17440 (N_17440,N_16562,N_16846);
nand U17441 (N_17441,N_16628,N_16560);
nor U17442 (N_17442,N_16884,N_16547);
and U17443 (N_17443,N_16847,N_16747);
or U17444 (N_17444,N_16909,N_16533);
nand U17445 (N_17445,N_16996,N_16960);
or U17446 (N_17446,N_16673,N_16819);
nor U17447 (N_17447,N_16650,N_16815);
or U17448 (N_17448,N_16964,N_16563);
nand U17449 (N_17449,N_16879,N_16865);
nand U17450 (N_17450,N_16554,N_16986);
nor U17451 (N_17451,N_16628,N_16633);
nand U17452 (N_17452,N_16612,N_16919);
and U17453 (N_17453,N_16690,N_16660);
xor U17454 (N_17454,N_16702,N_16960);
or U17455 (N_17455,N_16675,N_16889);
nand U17456 (N_17456,N_16883,N_16686);
nor U17457 (N_17457,N_16632,N_16649);
or U17458 (N_17458,N_16840,N_16591);
and U17459 (N_17459,N_16906,N_16840);
and U17460 (N_17460,N_16534,N_16583);
and U17461 (N_17461,N_16847,N_16675);
and U17462 (N_17462,N_16739,N_16970);
nand U17463 (N_17463,N_16764,N_16803);
nor U17464 (N_17464,N_16727,N_16661);
nand U17465 (N_17465,N_16728,N_16531);
and U17466 (N_17466,N_16549,N_16828);
or U17467 (N_17467,N_16544,N_16915);
nand U17468 (N_17468,N_16759,N_16620);
nor U17469 (N_17469,N_16869,N_16885);
or U17470 (N_17470,N_16573,N_16510);
xnor U17471 (N_17471,N_16578,N_16715);
and U17472 (N_17472,N_16989,N_16986);
nand U17473 (N_17473,N_16650,N_16868);
and U17474 (N_17474,N_16745,N_16682);
xnor U17475 (N_17475,N_16648,N_16722);
or U17476 (N_17476,N_16835,N_16837);
or U17477 (N_17477,N_16922,N_16624);
nand U17478 (N_17478,N_16736,N_16882);
or U17479 (N_17479,N_16880,N_16511);
and U17480 (N_17480,N_16821,N_16876);
xor U17481 (N_17481,N_16989,N_16703);
and U17482 (N_17482,N_16819,N_16514);
nand U17483 (N_17483,N_16933,N_16760);
nand U17484 (N_17484,N_16892,N_16590);
nor U17485 (N_17485,N_16613,N_16542);
nand U17486 (N_17486,N_16835,N_16901);
nor U17487 (N_17487,N_16947,N_16628);
xnor U17488 (N_17488,N_16921,N_16516);
or U17489 (N_17489,N_16989,N_16606);
xor U17490 (N_17490,N_16831,N_16731);
xor U17491 (N_17491,N_16577,N_16704);
and U17492 (N_17492,N_16580,N_16784);
or U17493 (N_17493,N_16789,N_16908);
nor U17494 (N_17494,N_16674,N_16971);
nor U17495 (N_17495,N_16561,N_16880);
nor U17496 (N_17496,N_16929,N_16525);
and U17497 (N_17497,N_16700,N_16851);
nand U17498 (N_17498,N_16801,N_16656);
nor U17499 (N_17499,N_16689,N_16953);
nand U17500 (N_17500,N_17238,N_17364);
nor U17501 (N_17501,N_17309,N_17143);
nor U17502 (N_17502,N_17409,N_17225);
nand U17503 (N_17503,N_17389,N_17315);
nand U17504 (N_17504,N_17060,N_17417);
and U17505 (N_17505,N_17075,N_17144);
and U17506 (N_17506,N_17290,N_17304);
xnor U17507 (N_17507,N_17092,N_17473);
and U17508 (N_17508,N_17283,N_17188);
or U17509 (N_17509,N_17124,N_17470);
or U17510 (N_17510,N_17197,N_17317);
nor U17511 (N_17511,N_17475,N_17168);
or U17512 (N_17512,N_17125,N_17151);
xnor U17513 (N_17513,N_17160,N_17268);
and U17514 (N_17514,N_17014,N_17138);
nor U17515 (N_17515,N_17469,N_17301);
and U17516 (N_17516,N_17205,N_17215);
nor U17517 (N_17517,N_17491,N_17208);
or U17518 (N_17518,N_17049,N_17085);
or U17519 (N_17519,N_17286,N_17093);
and U17520 (N_17520,N_17045,N_17267);
nor U17521 (N_17521,N_17111,N_17146);
nand U17522 (N_17522,N_17436,N_17156);
nand U17523 (N_17523,N_17010,N_17278);
and U17524 (N_17524,N_17008,N_17349);
and U17525 (N_17525,N_17058,N_17372);
xor U17526 (N_17526,N_17166,N_17173);
or U17527 (N_17527,N_17171,N_17280);
nor U17528 (N_17528,N_17257,N_17303);
and U17529 (N_17529,N_17441,N_17292);
xor U17530 (N_17530,N_17438,N_17416);
xor U17531 (N_17531,N_17019,N_17312);
nor U17532 (N_17532,N_17451,N_17313);
nand U17533 (N_17533,N_17499,N_17204);
xor U17534 (N_17534,N_17408,N_17424);
xor U17535 (N_17535,N_17172,N_17359);
or U17536 (N_17536,N_17229,N_17161);
or U17537 (N_17537,N_17202,N_17114);
nor U17538 (N_17538,N_17291,N_17159);
xnor U17539 (N_17539,N_17134,N_17034);
nor U17540 (N_17540,N_17064,N_17331);
or U17541 (N_17541,N_17360,N_17355);
or U17542 (N_17542,N_17285,N_17320);
nor U17543 (N_17543,N_17232,N_17153);
and U17544 (N_17544,N_17235,N_17090);
or U17545 (N_17545,N_17494,N_17220);
xnor U17546 (N_17546,N_17484,N_17425);
xnor U17547 (N_17547,N_17270,N_17463);
and U17548 (N_17548,N_17383,N_17209);
nor U17549 (N_17549,N_17490,N_17239);
and U17550 (N_17550,N_17017,N_17284);
nand U17551 (N_17551,N_17094,N_17422);
xnor U17552 (N_17552,N_17460,N_17420);
or U17553 (N_17553,N_17057,N_17023);
nand U17554 (N_17554,N_17015,N_17190);
xor U17555 (N_17555,N_17071,N_17405);
nand U17556 (N_17556,N_17224,N_17080);
nor U17557 (N_17557,N_17454,N_17311);
nand U17558 (N_17558,N_17376,N_17103);
or U17559 (N_17559,N_17261,N_17082);
xor U17560 (N_17560,N_17002,N_17192);
xor U17561 (N_17561,N_17180,N_17065);
nand U17562 (N_17562,N_17401,N_17236);
or U17563 (N_17563,N_17339,N_17427);
xor U17564 (N_17564,N_17423,N_17222);
and U17565 (N_17565,N_17402,N_17147);
nand U17566 (N_17566,N_17009,N_17186);
and U17567 (N_17567,N_17025,N_17377);
xnor U17568 (N_17568,N_17366,N_17458);
xor U17569 (N_17569,N_17345,N_17411);
or U17570 (N_17570,N_17245,N_17437);
nor U17571 (N_17571,N_17101,N_17478);
nor U17572 (N_17572,N_17467,N_17293);
and U17573 (N_17573,N_17145,N_17480);
and U17574 (N_17574,N_17382,N_17096);
or U17575 (N_17575,N_17018,N_17052);
nand U17576 (N_17576,N_17026,N_17195);
and U17577 (N_17577,N_17200,N_17353);
nand U17578 (N_17578,N_17474,N_17260);
nand U17579 (N_17579,N_17048,N_17234);
nor U17580 (N_17580,N_17007,N_17005);
nor U17581 (N_17581,N_17373,N_17165);
or U17582 (N_17582,N_17051,N_17477);
or U17583 (N_17583,N_17403,N_17374);
xor U17584 (N_17584,N_17078,N_17148);
nand U17585 (N_17585,N_17446,N_17095);
nand U17586 (N_17586,N_17252,N_17227);
nand U17587 (N_17587,N_17479,N_17448);
nand U17588 (N_17588,N_17350,N_17242);
nor U17589 (N_17589,N_17219,N_17191);
or U17590 (N_17590,N_17329,N_17097);
xor U17591 (N_17591,N_17184,N_17126);
nand U17592 (N_17592,N_17340,N_17249);
nand U17593 (N_17593,N_17336,N_17496);
nand U17594 (N_17594,N_17091,N_17120);
nand U17595 (N_17595,N_17117,N_17039);
nor U17596 (N_17596,N_17321,N_17136);
nor U17597 (N_17597,N_17170,N_17447);
nor U17598 (N_17598,N_17476,N_17206);
or U17599 (N_17599,N_17119,N_17063);
nand U17600 (N_17600,N_17237,N_17110);
or U17601 (N_17601,N_17073,N_17352);
nor U17602 (N_17602,N_17388,N_17187);
xor U17603 (N_17603,N_17356,N_17419);
or U17604 (N_17604,N_17387,N_17378);
and U17605 (N_17605,N_17397,N_17324);
or U17606 (N_17606,N_17489,N_17011);
xnor U17607 (N_17607,N_17358,N_17322);
nor U17608 (N_17608,N_17036,N_17047);
nand U17609 (N_17609,N_17129,N_17294);
xnor U17610 (N_17610,N_17053,N_17406);
nor U17611 (N_17611,N_17128,N_17337);
and U17612 (N_17612,N_17254,N_17139);
xnor U17613 (N_17613,N_17410,N_17158);
nand U17614 (N_17614,N_17105,N_17141);
or U17615 (N_17615,N_17299,N_17455);
and U17616 (N_17616,N_17282,N_17330);
and U17617 (N_17617,N_17287,N_17230);
xnor U17618 (N_17618,N_17354,N_17497);
or U17619 (N_17619,N_17182,N_17308);
or U17620 (N_17620,N_17107,N_17177);
nor U17621 (N_17621,N_17203,N_17346);
and U17622 (N_17622,N_17465,N_17189);
xor U17623 (N_17623,N_17279,N_17109);
nand U17624 (N_17624,N_17162,N_17115);
or U17625 (N_17625,N_17462,N_17342);
and U17626 (N_17626,N_17127,N_17248);
nand U17627 (N_17627,N_17174,N_17307);
xnor U17628 (N_17628,N_17046,N_17264);
and U17629 (N_17629,N_17233,N_17179);
and U17630 (N_17630,N_17196,N_17440);
nor U17631 (N_17631,N_17483,N_17221);
nor U17632 (N_17632,N_17000,N_17368);
or U17633 (N_17633,N_17262,N_17338);
xor U17634 (N_17634,N_17083,N_17271);
nor U17635 (N_17635,N_17256,N_17181);
nor U17636 (N_17636,N_17449,N_17013);
and U17637 (N_17637,N_17185,N_17343);
nor U17638 (N_17638,N_17472,N_17394);
nor U17639 (N_17639,N_17488,N_17296);
xnor U17640 (N_17640,N_17032,N_17067);
nand U17641 (N_17641,N_17391,N_17390);
and U17642 (N_17642,N_17487,N_17006);
nand U17643 (N_17643,N_17395,N_17361);
nand U17644 (N_17644,N_17061,N_17211);
or U17645 (N_17645,N_17421,N_17108);
or U17646 (N_17646,N_17121,N_17041);
nand U17647 (N_17647,N_17485,N_17439);
and U17648 (N_17648,N_17131,N_17258);
or U17649 (N_17649,N_17042,N_17323);
or U17650 (N_17650,N_17468,N_17210);
and U17651 (N_17651,N_17297,N_17194);
xor U17652 (N_17652,N_17123,N_17444);
or U17653 (N_17653,N_17266,N_17302);
nor U17654 (N_17654,N_17415,N_17021);
nor U17655 (N_17655,N_17265,N_17231);
and U17656 (N_17656,N_17244,N_17399);
xor U17657 (N_17657,N_17432,N_17152);
xnor U17658 (N_17658,N_17466,N_17433);
or U17659 (N_17659,N_17223,N_17251);
nor U17660 (N_17660,N_17459,N_17167);
or U17661 (N_17661,N_17426,N_17450);
or U17662 (N_17662,N_17149,N_17347);
or U17663 (N_17663,N_17498,N_17443);
and U17664 (N_17664,N_17493,N_17068);
nor U17665 (N_17665,N_17319,N_17250);
nor U17666 (N_17666,N_17272,N_17089);
or U17667 (N_17667,N_17456,N_17298);
nand U17668 (N_17668,N_17164,N_17059);
xor U17669 (N_17669,N_17481,N_17122);
nor U17670 (N_17670,N_17098,N_17038);
and U17671 (N_17671,N_17022,N_17012);
xnor U17672 (N_17672,N_17275,N_17412);
nand U17673 (N_17673,N_17207,N_17461);
and U17674 (N_17674,N_17132,N_17326);
xor U17675 (N_17675,N_17193,N_17431);
nand U17676 (N_17676,N_17453,N_17169);
nor U17677 (N_17677,N_17418,N_17385);
and U17678 (N_17678,N_17327,N_17037);
nor U17679 (N_17679,N_17367,N_17216);
and U17680 (N_17680,N_17056,N_17375);
and U17681 (N_17681,N_17281,N_17079);
nor U17682 (N_17682,N_17076,N_17043);
or U17683 (N_17683,N_17163,N_17135);
nor U17684 (N_17684,N_17226,N_17001);
and U17685 (N_17685,N_17428,N_17381);
nor U17686 (N_17686,N_17365,N_17457);
xor U17687 (N_17687,N_17404,N_17253);
or U17688 (N_17688,N_17066,N_17393);
nor U17689 (N_17689,N_17031,N_17054);
or U17690 (N_17690,N_17102,N_17396);
and U17691 (N_17691,N_17295,N_17178);
xnor U17692 (N_17692,N_17198,N_17118);
nor U17693 (N_17693,N_17314,N_17482);
nor U17694 (N_17694,N_17062,N_17269);
nand U17695 (N_17695,N_17407,N_17333);
nand U17696 (N_17696,N_17112,N_17199);
nand U17697 (N_17697,N_17429,N_17310);
nor U17698 (N_17698,N_17289,N_17100);
xnor U17699 (N_17699,N_17113,N_17104);
nor U17700 (N_17700,N_17243,N_17072);
and U17701 (N_17701,N_17413,N_17212);
xor U17702 (N_17702,N_17150,N_17398);
nand U17703 (N_17703,N_17069,N_17247);
nor U17704 (N_17704,N_17070,N_17471);
and U17705 (N_17705,N_17228,N_17130);
and U17706 (N_17706,N_17142,N_17318);
and U17707 (N_17707,N_17028,N_17334);
or U17708 (N_17708,N_17306,N_17035);
nand U17709 (N_17709,N_17328,N_17445);
or U17710 (N_17710,N_17081,N_17380);
nor U17711 (N_17711,N_17074,N_17087);
nand U17712 (N_17712,N_17040,N_17213);
xnor U17713 (N_17713,N_17442,N_17116);
xnor U17714 (N_17714,N_17003,N_17240);
and U17715 (N_17715,N_17217,N_17348);
or U17716 (N_17716,N_17435,N_17273);
and U17717 (N_17717,N_17175,N_17176);
or U17718 (N_17718,N_17369,N_17452);
xnor U17719 (N_17719,N_17029,N_17392);
or U17720 (N_17720,N_17430,N_17020);
or U17721 (N_17721,N_17332,N_17084);
xor U17722 (N_17722,N_17379,N_17400);
and U17723 (N_17723,N_17140,N_17274);
nor U17724 (N_17724,N_17033,N_17183);
or U17725 (N_17725,N_17434,N_17414);
xnor U17726 (N_17726,N_17106,N_17486);
and U17727 (N_17727,N_17316,N_17464);
or U17728 (N_17728,N_17154,N_17086);
nand U17729 (N_17729,N_17344,N_17351);
nor U17730 (N_17730,N_17495,N_17218);
nand U17731 (N_17731,N_17004,N_17370);
nand U17732 (N_17732,N_17214,N_17246);
xnor U17733 (N_17733,N_17362,N_17288);
xnor U17734 (N_17734,N_17357,N_17024);
or U17735 (N_17735,N_17305,N_17077);
nor U17736 (N_17736,N_17099,N_17325);
and U17737 (N_17737,N_17044,N_17055);
nand U17738 (N_17738,N_17335,N_17137);
nand U17739 (N_17739,N_17276,N_17371);
and U17740 (N_17740,N_17133,N_17157);
nor U17741 (N_17741,N_17386,N_17492);
nor U17742 (N_17742,N_17050,N_17027);
or U17743 (N_17743,N_17263,N_17201);
and U17744 (N_17744,N_17241,N_17259);
nand U17745 (N_17745,N_17341,N_17030);
xnor U17746 (N_17746,N_17088,N_17255);
nand U17747 (N_17747,N_17277,N_17155);
or U17748 (N_17748,N_17016,N_17363);
and U17749 (N_17749,N_17300,N_17384);
and U17750 (N_17750,N_17033,N_17184);
nand U17751 (N_17751,N_17344,N_17436);
nor U17752 (N_17752,N_17444,N_17352);
or U17753 (N_17753,N_17127,N_17074);
and U17754 (N_17754,N_17472,N_17182);
or U17755 (N_17755,N_17203,N_17268);
nand U17756 (N_17756,N_17439,N_17284);
nor U17757 (N_17757,N_17280,N_17198);
or U17758 (N_17758,N_17032,N_17231);
nand U17759 (N_17759,N_17111,N_17245);
and U17760 (N_17760,N_17193,N_17039);
and U17761 (N_17761,N_17190,N_17042);
and U17762 (N_17762,N_17095,N_17261);
nand U17763 (N_17763,N_17108,N_17498);
xnor U17764 (N_17764,N_17257,N_17004);
nand U17765 (N_17765,N_17158,N_17101);
nor U17766 (N_17766,N_17332,N_17091);
nand U17767 (N_17767,N_17117,N_17146);
or U17768 (N_17768,N_17190,N_17082);
and U17769 (N_17769,N_17409,N_17447);
nor U17770 (N_17770,N_17129,N_17184);
nand U17771 (N_17771,N_17190,N_17268);
or U17772 (N_17772,N_17097,N_17451);
and U17773 (N_17773,N_17362,N_17153);
nor U17774 (N_17774,N_17431,N_17350);
nor U17775 (N_17775,N_17425,N_17045);
and U17776 (N_17776,N_17160,N_17390);
and U17777 (N_17777,N_17340,N_17148);
nand U17778 (N_17778,N_17407,N_17395);
xor U17779 (N_17779,N_17491,N_17426);
or U17780 (N_17780,N_17047,N_17486);
xnor U17781 (N_17781,N_17302,N_17108);
nor U17782 (N_17782,N_17253,N_17132);
nand U17783 (N_17783,N_17437,N_17206);
nor U17784 (N_17784,N_17202,N_17490);
and U17785 (N_17785,N_17188,N_17338);
and U17786 (N_17786,N_17099,N_17366);
and U17787 (N_17787,N_17450,N_17111);
and U17788 (N_17788,N_17217,N_17417);
or U17789 (N_17789,N_17265,N_17287);
and U17790 (N_17790,N_17084,N_17278);
nor U17791 (N_17791,N_17156,N_17191);
nor U17792 (N_17792,N_17244,N_17184);
and U17793 (N_17793,N_17111,N_17186);
nand U17794 (N_17794,N_17206,N_17421);
nor U17795 (N_17795,N_17403,N_17122);
xnor U17796 (N_17796,N_17217,N_17177);
and U17797 (N_17797,N_17341,N_17313);
and U17798 (N_17798,N_17117,N_17140);
xnor U17799 (N_17799,N_17428,N_17293);
or U17800 (N_17800,N_17365,N_17275);
nor U17801 (N_17801,N_17043,N_17282);
nor U17802 (N_17802,N_17106,N_17376);
nand U17803 (N_17803,N_17387,N_17202);
xor U17804 (N_17804,N_17189,N_17323);
nand U17805 (N_17805,N_17029,N_17210);
nor U17806 (N_17806,N_17236,N_17025);
nand U17807 (N_17807,N_17064,N_17202);
and U17808 (N_17808,N_17292,N_17084);
xnor U17809 (N_17809,N_17370,N_17284);
xor U17810 (N_17810,N_17252,N_17089);
and U17811 (N_17811,N_17456,N_17186);
xor U17812 (N_17812,N_17117,N_17240);
and U17813 (N_17813,N_17068,N_17454);
nand U17814 (N_17814,N_17176,N_17179);
or U17815 (N_17815,N_17320,N_17371);
nor U17816 (N_17816,N_17442,N_17096);
and U17817 (N_17817,N_17253,N_17474);
xnor U17818 (N_17818,N_17135,N_17383);
or U17819 (N_17819,N_17102,N_17049);
nand U17820 (N_17820,N_17176,N_17397);
or U17821 (N_17821,N_17190,N_17168);
nand U17822 (N_17822,N_17202,N_17374);
and U17823 (N_17823,N_17055,N_17119);
xnor U17824 (N_17824,N_17276,N_17159);
xor U17825 (N_17825,N_17097,N_17423);
or U17826 (N_17826,N_17331,N_17444);
nor U17827 (N_17827,N_17064,N_17081);
or U17828 (N_17828,N_17326,N_17038);
nor U17829 (N_17829,N_17011,N_17410);
nor U17830 (N_17830,N_17494,N_17117);
or U17831 (N_17831,N_17199,N_17455);
nor U17832 (N_17832,N_17159,N_17043);
xor U17833 (N_17833,N_17194,N_17166);
nor U17834 (N_17834,N_17240,N_17370);
nand U17835 (N_17835,N_17267,N_17362);
xor U17836 (N_17836,N_17249,N_17377);
xor U17837 (N_17837,N_17043,N_17419);
nand U17838 (N_17838,N_17169,N_17137);
nand U17839 (N_17839,N_17483,N_17161);
xnor U17840 (N_17840,N_17399,N_17470);
nor U17841 (N_17841,N_17291,N_17317);
and U17842 (N_17842,N_17121,N_17196);
or U17843 (N_17843,N_17416,N_17425);
or U17844 (N_17844,N_17330,N_17366);
or U17845 (N_17845,N_17235,N_17434);
nor U17846 (N_17846,N_17276,N_17060);
nand U17847 (N_17847,N_17117,N_17083);
xnor U17848 (N_17848,N_17401,N_17157);
and U17849 (N_17849,N_17395,N_17061);
or U17850 (N_17850,N_17179,N_17349);
and U17851 (N_17851,N_17013,N_17335);
and U17852 (N_17852,N_17244,N_17379);
nor U17853 (N_17853,N_17165,N_17498);
and U17854 (N_17854,N_17142,N_17255);
nand U17855 (N_17855,N_17325,N_17219);
or U17856 (N_17856,N_17411,N_17263);
or U17857 (N_17857,N_17427,N_17296);
and U17858 (N_17858,N_17250,N_17018);
nand U17859 (N_17859,N_17081,N_17474);
xnor U17860 (N_17860,N_17149,N_17013);
xor U17861 (N_17861,N_17132,N_17356);
or U17862 (N_17862,N_17203,N_17237);
nor U17863 (N_17863,N_17463,N_17478);
and U17864 (N_17864,N_17426,N_17088);
nor U17865 (N_17865,N_17413,N_17070);
nand U17866 (N_17866,N_17339,N_17195);
and U17867 (N_17867,N_17441,N_17280);
nand U17868 (N_17868,N_17433,N_17147);
and U17869 (N_17869,N_17181,N_17257);
xor U17870 (N_17870,N_17213,N_17003);
nand U17871 (N_17871,N_17388,N_17030);
xor U17872 (N_17872,N_17432,N_17414);
xnor U17873 (N_17873,N_17427,N_17096);
nor U17874 (N_17874,N_17295,N_17094);
or U17875 (N_17875,N_17008,N_17288);
xor U17876 (N_17876,N_17093,N_17253);
nor U17877 (N_17877,N_17164,N_17212);
nand U17878 (N_17878,N_17222,N_17254);
xor U17879 (N_17879,N_17185,N_17132);
xor U17880 (N_17880,N_17047,N_17178);
nand U17881 (N_17881,N_17159,N_17122);
and U17882 (N_17882,N_17348,N_17129);
or U17883 (N_17883,N_17037,N_17366);
xnor U17884 (N_17884,N_17354,N_17050);
xnor U17885 (N_17885,N_17384,N_17047);
nand U17886 (N_17886,N_17132,N_17357);
nand U17887 (N_17887,N_17423,N_17403);
or U17888 (N_17888,N_17277,N_17116);
and U17889 (N_17889,N_17424,N_17082);
and U17890 (N_17890,N_17265,N_17013);
xor U17891 (N_17891,N_17441,N_17040);
nor U17892 (N_17892,N_17093,N_17369);
or U17893 (N_17893,N_17050,N_17306);
and U17894 (N_17894,N_17153,N_17292);
nand U17895 (N_17895,N_17333,N_17018);
xor U17896 (N_17896,N_17254,N_17421);
or U17897 (N_17897,N_17281,N_17137);
xor U17898 (N_17898,N_17453,N_17355);
nand U17899 (N_17899,N_17328,N_17446);
or U17900 (N_17900,N_17139,N_17140);
or U17901 (N_17901,N_17215,N_17001);
nand U17902 (N_17902,N_17317,N_17446);
or U17903 (N_17903,N_17305,N_17324);
nor U17904 (N_17904,N_17083,N_17130);
or U17905 (N_17905,N_17285,N_17454);
xor U17906 (N_17906,N_17343,N_17384);
and U17907 (N_17907,N_17323,N_17296);
or U17908 (N_17908,N_17108,N_17427);
nand U17909 (N_17909,N_17404,N_17179);
nand U17910 (N_17910,N_17495,N_17312);
or U17911 (N_17911,N_17379,N_17351);
nor U17912 (N_17912,N_17339,N_17014);
xnor U17913 (N_17913,N_17131,N_17115);
and U17914 (N_17914,N_17387,N_17148);
and U17915 (N_17915,N_17210,N_17338);
nand U17916 (N_17916,N_17072,N_17434);
xor U17917 (N_17917,N_17278,N_17192);
and U17918 (N_17918,N_17228,N_17060);
and U17919 (N_17919,N_17423,N_17253);
and U17920 (N_17920,N_17425,N_17304);
xnor U17921 (N_17921,N_17394,N_17192);
nor U17922 (N_17922,N_17080,N_17095);
nand U17923 (N_17923,N_17456,N_17210);
and U17924 (N_17924,N_17174,N_17421);
xor U17925 (N_17925,N_17292,N_17379);
or U17926 (N_17926,N_17345,N_17262);
nor U17927 (N_17927,N_17448,N_17209);
and U17928 (N_17928,N_17484,N_17405);
nor U17929 (N_17929,N_17045,N_17375);
xor U17930 (N_17930,N_17019,N_17176);
xnor U17931 (N_17931,N_17476,N_17456);
nor U17932 (N_17932,N_17027,N_17358);
nor U17933 (N_17933,N_17107,N_17231);
and U17934 (N_17934,N_17378,N_17423);
nor U17935 (N_17935,N_17263,N_17412);
xnor U17936 (N_17936,N_17356,N_17193);
and U17937 (N_17937,N_17156,N_17383);
or U17938 (N_17938,N_17381,N_17102);
nor U17939 (N_17939,N_17471,N_17230);
xor U17940 (N_17940,N_17061,N_17175);
nand U17941 (N_17941,N_17437,N_17372);
nand U17942 (N_17942,N_17029,N_17045);
nand U17943 (N_17943,N_17113,N_17305);
nand U17944 (N_17944,N_17277,N_17446);
and U17945 (N_17945,N_17415,N_17404);
xnor U17946 (N_17946,N_17477,N_17374);
and U17947 (N_17947,N_17142,N_17025);
nor U17948 (N_17948,N_17345,N_17498);
nor U17949 (N_17949,N_17157,N_17454);
xor U17950 (N_17950,N_17374,N_17110);
nand U17951 (N_17951,N_17493,N_17222);
xor U17952 (N_17952,N_17324,N_17374);
xnor U17953 (N_17953,N_17051,N_17453);
xor U17954 (N_17954,N_17108,N_17219);
or U17955 (N_17955,N_17254,N_17123);
or U17956 (N_17956,N_17279,N_17236);
or U17957 (N_17957,N_17453,N_17070);
nor U17958 (N_17958,N_17054,N_17058);
nand U17959 (N_17959,N_17061,N_17322);
and U17960 (N_17960,N_17076,N_17277);
and U17961 (N_17961,N_17007,N_17355);
nand U17962 (N_17962,N_17210,N_17108);
nand U17963 (N_17963,N_17408,N_17059);
nand U17964 (N_17964,N_17113,N_17016);
nor U17965 (N_17965,N_17375,N_17414);
and U17966 (N_17966,N_17365,N_17498);
xor U17967 (N_17967,N_17002,N_17046);
or U17968 (N_17968,N_17208,N_17016);
and U17969 (N_17969,N_17105,N_17290);
and U17970 (N_17970,N_17431,N_17334);
nor U17971 (N_17971,N_17275,N_17174);
and U17972 (N_17972,N_17314,N_17403);
and U17973 (N_17973,N_17041,N_17498);
nor U17974 (N_17974,N_17008,N_17187);
nand U17975 (N_17975,N_17259,N_17103);
nor U17976 (N_17976,N_17284,N_17083);
and U17977 (N_17977,N_17211,N_17286);
or U17978 (N_17978,N_17455,N_17248);
and U17979 (N_17979,N_17073,N_17264);
and U17980 (N_17980,N_17188,N_17218);
xnor U17981 (N_17981,N_17241,N_17432);
and U17982 (N_17982,N_17335,N_17325);
xor U17983 (N_17983,N_17348,N_17074);
and U17984 (N_17984,N_17137,N_17492);
nand U17985 (N_17985,N_17217,N_17086);
nor U17986 (N_17986,N_17419,N_17378);
xor U17987 (N_17987,N_17051,N_17376);
and U17988 (N_17988,N_17176,N_17169);
and U17989 (N_17989,N_17225,N_17156);
nand U17990 (N_17990,N_17397,N_17392);
or U17991 (N_17991,N_17273,N_17192);
nor U17992 (N_17992,N_17090,N_17428);
nand U17993 (N_17993,N_17021,N_17338);
and U17994 (N_17994,N_17489,N_17116);
and U17995 (N_17995,N_17031,N_17475);
or U17996 (N_17996,N_17071,N_17450);
or U17997 (N_17997,N_17127,N_17466);
and U17998 (N_17998,N_17301,N_17152);
nand U17999 (N_17999,N_17108,N_17284);
xnor U18000 (N_18000,N_17695,N_17766);
xor U18001 (N_18001,N_17760,N_17761);
xnor U18002 (N_18002,N_17911,N_17827);
nor U18003 (N_18003,N_17910,N_17600);
xor U18004 (N_18004,N_17670,N_17717);
and U18005 (N_18005,N_17691,N_17625);
nand U18006 (N_18006,N_17606,N_17664);
xnor U18007 (N_18007,N_17641,N_17627);
or U18008 (N_18008,N_17500,N_17979);
xor U18009 (N_18009,N_17992,N_17983);
and U18010 (N_18010,N_17531,N_17968);
or U18011 (N_18011,N_17564,N_17604);
xnor U18012 (N_18012,N_17607,N_17608);
and U18013 (N_18013,N_17700,N_17730);
xor U18014 (N_18014,N_17689,N_17503);
and U18015 (N_18015,N_17648,N_17985);
nor U18016 (N_18016,N_17643,N_17721);
and U18017 (N_18017,N_17950,N_17711);
or U18018 (N_18018,N_17559,N_17501);
xnor U18019 (N_18019,N_17969,N_17954);
and U18020 (N_18020,N_17757,N_17510);
or U18021 (N_18021,N_17772,N_17962);
nor U18022 (N_18022,N_17779,N_17519);
xnor U18023 (N_18023,N_17633,N_17795);
xnor U18024 (N_18024,N_17907,N_17538);
and U18025 (N_18025,N_17862,N_17617);
or U18026 (N_18026,N_17666,N_17602);
nor U18027 (N_18027,N_17785,N_17556);
nor U18028 (N_18028,N_17642,N_17825);
and U18029 (N_18029,N_17994,N_17879);
or U18030 (N_18030,N_17770,N_17776);
nand U18031 (N_18031,N_17736,N_17850);
or U18032 (N_18032,N_17599,N_17735);
or U18033 (N_18033,N_17914,N_17566);
or U18034 (N_18034,N_17558,N_17596);
xor U18035 (N_18035,N_17589,N_17814);
nor U18036 (N_18036,N_17913,N_17810);
nor U18037 (N_18037,N_17886,N_17672);
xnor U18038 (N_18038,N_17540,N_17842);
nor U18039 (N_18039,N_17553,N_17680);
xnor U18040 (N_18040,N_17650,N_17588);
xnor U18041 (N_18041,N_17967,N_17533);
xor U18042 (N_18042,N_17763,N_17991);
nor U18043 (N_18043,N_17861,N_17720);
nand U18044 (N_18044,N_17819,N_17733);
xor U18045 (N_18045,N_17514,N_17561);
and U18046 (N_18046,N_17637,N_17848);
nor U18047 (N_18047,N_17527,N_17507);
nor U18048 (N_18048,N_17667,N_17894);
xor U18049 (N_18049,N_17509,N_17880);
or U18050 (N_18050,N_17806,N_17638);
xnor U18051 (N_18051,N_17869,N_17807);
nor U18052 (N_18052,N_17535,N_17833);
or U18053 (N_18053,N_17937,N_17528);
nor U18054 (N_18054,N_17669,N_17959);
or U18055 (N_18055,N_17927,N_17657);
or U18056 (N_18056,N_17934,N_17928);
or U18057 (N_18057,N_17512,N_17621);
or U18058 (N_18058,N_17921,N_17836);
or U18059 (N_18059,N_17671,N_17876);
and U18060 (N_18060,N_17645,N_17694);
or U18061 (N_18061,N_17984,N_17925);
and U18062 (N_18062,N_17539,N_17773);
or U18063 (N_18063,N_17636,N_17811);
or U18064 (N_18064,N_17947,N_17567);
xnor U18065 (N_18065,N_17919,N_17892);
xnor U18066 (N_18066,N_17997,N_17552);
xor U18067 (N_18067,N_17603,N_17788);
nor U18068 (N_18068,N_17723,N_17605);
nand U18069 (N_18069,N_17874,N_17809);
xnor U18070 (N_18070,N_17595,N_17804);
xnor U18071 (N_18071,N_17549,N_17826);
nor U18072 (N_18072,N_17956,N_17935);
nor U18073 (N_18073,N_17777,N_17629);
xor U18074 (N_18074,N_17731,N_17631);
nor U18075 (N_18075,N_17855,N_17727);
and U18076 (N_18076,N_17745,N_17513);
xor U18077 (N_18077,N_17893,N_17725);
xor U18078 (N_18078,N_17949,N_17601);
or U18079 (N_18079,N_17975,N_17854);
nor U18080 (N_18080,N_17565,N_17523);
and U18081 (N_18081,N_17762,N_17891);
nand U18082 (N_18082,N_17652,N_17882);
or U18083 (N_18083,N_17787,N_17563);
xor U18084 (N_18084,N_17976,N_17915);
or U18085 (N_18085,N_17775,N_17574);
nand U18086 (N_18086,N_17570,N_17930);
xor U18087 (N_18087,N_17831,N_17734);
or U18088 (N_18088,N_17708,N_17709);
nand U18089 (N_18089,N_17665,N_17737);
nor U18090 (N_18090,N_17767,N_17659);
xor U18091 (N_18091,N_17557,N_17783);
nor U18092 (N_18092,N_17612,N_17995);
and U18093 (N_18093,N_17703,N_17774);
or U18094 (N_18094,N_17635,N_17634);
nor U18095 (N_18095,N_17578,N_17722);
nor U18096 (N_18096,N_17800,N_17678);
nand U18097 (N_18097,N_17609,N_17903);
and U18098 (N_18098,N_17820,N_17525);
and U18099 (N_18099,N_17957,N_17646);
nor U18100 (N_18100,N_17865,N_17802);
nor U18101 (N_18101,N_17614,N_17916);
and U18102 (N_18102,N_17545,N_17698);
nor U18103 (N_18103,N_17632,N_17996);
nand U18104 (N_18104,N_17555,N_17912);
nor U18105 (N_18105,N_17890,N_17920);
nor U18106 (N_18106,N_17948,N_17719);
nor U18107 (N_18107,N_17958,N_17541);
nand U18108 (N_18108,N_17579,N_17768);
and U18109 (N_18109,N_17748,N_17943);
nor U18110 (N_18110,N_17712,N_17577);
or U18111 (N_18111,N_17581,N_17778);
nor U18112 (N_18112,N_17989,N_17834);
or U18113 (N_18113,N_17562,N_17977);
nand U18114 (N_18114,N_17750,N_17789);
or U18115 (N_18115,N_17987,N_17837);
nand U18116 (N_18116,N_17841,N_17863);
nand U18117 (N_18117,N_17679,N_17917);
nand U18118 (N_18118,N_17803,N_17573);
xor U18119 (N_18119,N_17591,N_17551);
nor U18120 (N_18120,N_17839,N_17530);
nand U18121 (N_18121,N_17792,N_17981);
nand U18122 (N_18122,N_17986,N_17630);
nor U18123 (N_18123,N_17988,N_17815);
nand U18124 (N_18124,N_17851,N_17704);
or U18125 (N_18125,N_17529,N_17728);
or U18126 (N_18126,N_17952,N_17522);
or U18127 (N_18127,N_17686,N_17790);
nand U18128 (N_18128,N_17859,N_17547);
xnor U18129 (N_18129,N_17868,N_17951);
nor U18130 (N_18130,N_17676,N_17906);
or U18131 (N_18131,N_17857,N_17755);
and U18132 (N_18132,N_17515,N_17856);
or U18133 (N_18133,N_17924,N_17715);
nand U18134 (N_18134,N_17931,N_17942);
xnor U18135 (N_18135,N_17816,N_17946);
nor U18136 (N_18136,N_17569,N_17813);
nand U18137 (N_18137,N_17812,N_17938);
xor U18138 (N_18138,N_17651,N_17590);
nand U18139 (N_18139,N_17502,N_17918);
or U18140 (N_18140,N_17830,N_17724);
or U18141 (N_18141,N_17696,N_17970);
nand U18142 (N_18142,N_17611,N_17939);
and U18143 (N_18143,N_17808,N_17554);
nand U18144 (N_18144,N_17990,N_17878);
nor U18145 (N_18145,N_17845,N_17585);
xor U18146 (N_18146,N_17751,N_17858);
nor U18147 (N_18147,N_17697,N_17619);
and U18148 (N_18148,N_17662,N_17526);
nor U18149 (N_18149,N_17941,N_17622);
nand U18150 (N_18150,N_17687,N_17754);
nor U18151 (N_18151,N_17998,N_17944);
xnor U18152 (N_18152,N_17571,N_17899);
xor U18153 (N_18153,N_17705,N_17904);
nand U18154 (N_18154,N_17508,N_17888);
or U18155 (N_18155,N_17644,N_17654);
nand U18156 (N_18156,N_17884,N_17542);
nand U18157 (N_18157,N_17866,N_17769);
nor U18158 (N_18158,N_17932,N_17871);
and U18159 (N_18159,N_17823,N_17628);
xor U18160 (N_18160,N_17506,N_17692);
and U18161 (N_18161,N_17690,N_17681);
nand U18162 (N_18162,N_17505,N_17517);
xor U18163 (N_18163,N_17797,N_17647);
or U18164 (N_18164,N_17765,N_17901);
nor U18165 (N_18165,N_17504,N_17875);
nand U18166 (N_18166,N_17738,N_17610);
or U18167 (N_18167,N_17896,N_17818);
nor U18168 (N_18168,N_17518,N_17560);
nand U18169 (N_18169,N_17582,N_17753);
xnor U18170 (N_18170,N_17844,N_17592);
nand U18171 (N_18171,N_17598,N_17516);
xnor U18172 (N_18172,N_17713,N_17781);
xor U18173 (N_18173,N_17999,N_17618);
or U18174 (N_18174,N_17973,N_17534);
nand U18175 (N_18175,N_17974,N_17511);
nand U18176 (N_18176,N_17707,N_17674);
xor U18177 (N_18177,N_17828,N_17673);
xnor U18178 (N_18178,N_17744,N_17902);
xor U18179 (N_18179,N_17639,N_17758);
or U18180 (N_18180,N_17743,N_17624);
nor U18181 (N_18181,N_17840,N_17964);
nand U18182 (N_18182,N_17821,N_17759);
nor U18183 (N_18183,N_17798,N_17685);
and U18184 (N_18184,N_17701,N_17663);
xnor U18185 (N_18185,N_17764,N_17580);
xnor U18186 (N_18186,N_17955,N_17544);
xnor U18187 (N_18187,N_17742,N_17794);
nor U18188 (N_18188,N_17923,N_17747);
nor U18189 (N_18189,N_17796,N_17784);
or U18190 (N_18190,N_17960,N_17718);
nand U18191 (N_18191,N_17971,N_17817);
and U18192 (N_18192,N_17714,N_17849);
nor U18193 (N_18193,N_17829,N_17661);
xnor U18194 (N_18194,N_17702,N_17846);
and U18195 (N_18195,N_17749,N_17741);
and U18196 (N_18196,N_17791,N_17900);
or U18197 (N_18197,N_17576,N_17872);
or U18198 (N_18198,N_17867,N_17963);
or U18199 (N_18199,N_17655,N_17594);
or U18200 (N_18200,N_17572,N_17660);
xnor U18201 (N_18201,N_17961,N_17980);
and U18202 (N_18202,N_17739,N_17726);
or U18203 (N_18203,N_17877,N_17716);
nor U18204 (N_18204,N_17870,N_17940);
nand U18205 (N_18205,N_17583,N_17537);
xnor U18206 (N_18206,N_17546,N_17616);
and U18207 (N_18207,N_17847,N_17897);
and U18208 (N_18208,N_17682,N_17883);
xor U18209 (N_18209,N_17683,N_17587);
xnor U18210 (N_18210,N_17793,N_17568);
and U18211 (N_18211,N_17584,N_17675);
nand U18212 (N_18212,N_17688,N_17771);
and U18213 (N_18213,N_17905,N_17864);
nor U18214 (N_18214,N_17873,N_17597);
nand U18215 (N_18215,N_17684,N_17656);
nor U18216 (N_18216,N_17887,N_17699);
or U18217 (N_18217,N_17521,N_17752);
nor U18218 (N_18218,N_17832,N_17972);
nor U18219 (N_18219,N_17710,N_17860);
nor U18220 (N_18220,N_17732,N_17729);
nand U18221 (N_18221,N_17740,N_17922);
nand U18222 (N_18222,N_17575,N_17929);
nor U18223 (N_18223,N_17978,N_17966);
and U18224 (N_18224,N_17668,N_17926);
nand U18225 (N_18225,N_17805,N_17835);
xnor U18226 (N_18226,N_17586,N_17824);
and U18227 (N_18227,N_17693,N_17909);
and U18228 (N_18228,N_17780,N_17543);
nand U18229 (N_18229,N_17853,N_17653);
nand U18230 (N_18230,N_17898,N_17843);
xnor U18231 (N_18231,N_17953,N_17613);
xnor U18232 (N_18232,N_17548,N_17982);
and U18233 (N_18233,N_17801,N_17933);
and U18234 (N_18234,N_17623,N_17889);
nand U18235 (N_18235,N_17799,N_17852);
or U18236 (N_18236,N_17908,N_17649);
xnor U18237 (N_18237,N_17677,N_17626);
and U18238 (N_18238,N_17640,N_17786);
or U18239 (N_18239,N_17965,N_17615);
nand U18240 (N_18240,N_17706,N_17532);
nor U18241 (N_18241,N_17620,N_17756);
nor U18242 (N_18242,N_17881,N_17993);
nor U18243 (N_18243,N_17746,N_17838);
and U18244 (N_18244,N_17822,N_17936);
and U18245 (N_18245,N_17895,N_17520);
and U18246 (N_18246,N_17885,N_17536);
nor U18247 (N_18247,N_17593,N_17945);
and U18248 (N_18248,N_17550,N_17524);
nor U18249 (N_18249,N_17658,N_17782);
nand U18250 (N_18250,N_17709,N_17994);
nand U18251 (N_18251,N_17897,N_17798);
or U18252 (N_18252,N_17696,N_17884);
xnor U18253 (N_18253,N_17892,N_17883);
nor U18254 (N_18254,N_17525,N_17899);
xnor U18255 (N_18255,N_17854,N_17634);
nand U18256 (N_18256,N_17933,N_17903);
nand U18257 (N_18257,N_17903,N_17690);
xor U18258 (N_18258,N_17621,N_17818);
nor U18259 (N_18259,N_17513,N_17823);
nand U18260 (N_18260,N_17533,N_17826);
xnor U18261 (N_18261,N_17944,N_17627);
xnor U18262 (N_18262,N_17715,N_17991);
nand U18263 (N_18263,N_17695,N_17985);
nor U18264 (N_18264,N_17735,N_17502);
nor U18265 (N_18265,N_17576,N_17942);
nor U18266 (N_18266,N_17519,N_17767);
xnor U18267 (N_18267,N_17815,N_17594);
or U18268 (N_18268,N_17603,N_17542);
or U18269 (N_18269,N_17899,N_17770);
nand U18270 (N_18270,N_17684,N_17937);
or U18271 (N_18271,N_17790,N_17660);
and U18272 (N_18272,N_17697,N_17676);
nor U18273 (N_18273,N_17984,N_17675);
and U18274 (N_18274,N_17864,N_17685);
nor U18275 (N_18275,N_17705,N_17612);
and U18276 (N_18276,N_17771,N_17926);
nand U18277 (N_18277,N_17553,N_17591);
xnor U18278 (N_18278,N_17818,N_17987);
nor U18279 (N_18279,N_17789,N_17766);
or U18280 (N_18280,N_17727,N_17549);
nor U18281 (N_18281,N_17987,N_17966);
nand U18282 (N_18282,N_17775,N_17702);
xor U18283 (N_18283,N_17870,N_17944);
and U18284 (N_18284,N_17550,N_17600);
nor U18285 (N_18285,N_17581,N_17712);
xor U18286 (N_18286,N_17958,N_17869);
and U18287 (N_18287,N_17702,N_17730);
and U18288 (N_18288,N_17954,N_17960);
or U18289 (N_18289,N_17948,N_17833);
nand U18290 (N_18290,N_17821,N_17789);
xnor U18291 (N_18291,N_17858,N_17827);
nand U18292 (N_18292,N_17606,N_17697);
nor U18293 (N_18293,N_17901,N_17589);
nand U18294 (N_18294,N_17882,N_17619);
nor U18295 (N_18295,N_17870,N_17951);
or U18296 (N_18296,N_17703,N_17997);
or U18297 (N_18297,N_17910,N_17956);
xor U18298 (N_18298,N_17840,N_17745);
or U18299 (N_18299,N_17811,N_17923);
nor U18300 (N_18300,N_17868,N_17569);
or U18301 (N_18301,N_17894,N_17550);
nor U18302 (N_18302,N_17907,N_17840);
and U18303 (N_18303,N_17634,N_17965);
xor U18304 (N_18304,N_17666,N_17937);
or U18305 (N_18305,N_17914,N_17798);
and U18306 (N_18306,N_17908,N_17934);
nor U18307 (N_18307,N_17655,N_17922);
nand U18308 (N_18308,N_17767,N_17916);
nor U18309 (N_18309,N_17932,N_17767);
nor U18310 (N_18310,N_17847,N_17523);
and U18311 (N_18311,N_17689,N_17887);
nand U18312 (N_18312,N_17683,N_17523);
nor U18313 (N_18313,N_17667,N_17649);
nor U18314 (N_18314,N_17781,N_17519);
nor U18315 (N_18315,N_17635,N_17936);
and U18316 (N_18316,N_17980,N_17664);
nand U18317 (N_18317,N_17799,N_17712);
xor U18318 (N_18318,N_17529,N_17976);
nand U18319 (N_18319,N_17503,N_17986);
xnor U18320 (N_18320,N_17517,N_17590);
or U18321 (N_18321,N_17877,N_17698);
or U18322 (N_18322,N_17548,N_17813);
nand U18323 (N_18323,N_17693,N_17612);
xnor U18324 (N_18324,N_17914,N_17822);
nand U18325 (N_18325,N_17815,N_17622);
nor U18326 (N_18326,N_17614,N_17615);
or U18327 (N_18327,N_17747,N_17582);
and U18328 (N_18328,N_17967,N_17509);
xnor U18329 (N_18329,N_17910,N_17646);
nand U18330 (N_18330,N_17711,N_17918);
nor U18331 (N_18331,N_17681,N_17746);
nor U18332 (N_18332,N_17713,N_17582);
xnor U18333 (N_18333,N_17506,N_17591);
or U18334 (N_18334,N_17691,N_17525);
or U18335 (N_18335,N_17504,N_17581);
and U18336 (N_18336,N_17670,N_17704);
xnor U18337 (N_18337,N_17784,N_17768);
nor U18338 (N_18338,N_17528,N_17684);
xnor U18339 (N_18339,N_17867,N_17841);
xnor U18340 (N_18340,N_17810,N_17835);
or U18341 (N_18341,N_17971,N_17855);
and U18342 (N_18342,N_17963,N_17598);
nor U18343 (N_18343,N_17737,N_17756);
nor U18344 (N_18344,N_17865,N_17721);
and U18345 (N_18345,N_17881,N_17606);
nand U18346 (N_18346,N_17844,N_17768);
nand U18347 (N_18347,N_17676,N_17824);
xor U18348 (N_18348,N_17507,N_17915);
or U18349 (N_18349,N_17889,N_17650);
nand U18350 (N_18350,N_17589,N_17858);
and U18351 (N_18351,N_17845,N_17680);
or U18352 (N_18352,N_17893,N_17903);
nand U18353 (N_18353,N_17833,N_17648);
or U18354 (N_18354,N_17838,N_17909);
nor U18355 (N_18355,N_17636,N_17957);
nor U18356 (N_18356,N_17538,N_17979);
or U18357 (N_18357,N_17551,N_17707);
nand U18358 (N_18358,N_17583,N_17752);
xor U18359 (N_18359,N_17512,N_17927);
xor U18360 (N_18360,N_17845,N_17836);
or U18361 (N_18361,N_17820,N_17719);
and U18362 (N_18362,N_17845,N_17719);
nand U18363 (N_18363,N_17661,N_17514);
nor U18364 (N_18364,N_17533,N_17721);
xnor U18365 (N_18365,N_17987,N_17958);
and U18366 (N_18366,N_17984,N_17815);
nand U18367 (N_18367,N_17863,N_17805);
or U18368 (N_18368,N_17548,N_17635);
or U18369 (N_18369,N_17738,N_17927);
xor U18370 (N_18370,N_17881,N_17925);
nand U18371 (N_18371,N_17568,N_17733);
xnor U18372 (N_18372,N_17846,N_17778);
nand U18373 (N_18373,N_17503,N_17925);
nor U18374 (N_18374,N_17919,N_17909);
and U18375 (N_18375,N_17940,N_17948);
xnor U18376 (N_18376,N_17682,N_17923);
xor U18377 (N_18377,N_17930,N_17745);
and U18378 (N_18378,N_17838,N_17598);
xor U18379 (N_18379,N_17984,N_17937);
or U18380 (N_18380,N_17976,N_17726);
xor U18381 (N_18381,N_17535,N_17960);
and U18382 (N_18382,N_17873,N_17662);
nor U18383 (N_18383,N_17609,N_17519);
nand U18384 (N_18384,N_17606,N_17872);
nand U18385 (N_18385,N_17828,N_17860);
or U18386 (N_18386,N_17653,N_17601);
and U18387 (N_18387,N_17911,N_17592);
nand U18388 (N_18388,N_17698,N_17537);
nand U18389 (N_18389,N_17916,N_17830);
nor U18390 (N_18390,N_17706,N_17775);
xnor U18391 (N_18391,N_17731,N_17817);
xnor U18392 (N_18392,N_17873,N_17892);
or U18393 (N_18393,N_17543,N_17591);
xnor U18394 (N_18394,N_17807,N_17692);
nand U18395 (N_18395,N_17774,N_17570);
or U18396 (N_18396,N_17790,N_17548);
and U18397 (N_18397,N_17709,N_17907);
nand U18398 (N_18398,N_17939,N_17632);
nor U18399 (N_18399,N_17818,N_17949);
or U18400 (N_18400,N_17900,N_17562);
xor U18401 (N_18401,N_17792,N_17518);
nand U18402 (N_18402,N_17966,N_17516);
xor U18403 (N_18403,N_17994,N_17826);
nor U18404 (N_18404,N_17995,N_17813);
and U18405 (N_18405,N_17805,N_17954);
nor U18406 (N_18406,N_17921,N_17911);
and U18407 (N_18407,N_17598,N_17779);
nand U18408 (N_18408,N_17648,N_17598);
nor U18409 (N_18409,N_17671,N_17994);
nand U18410 (N_18410,N_17668,N_17794);
or U18411 (N_18411,N_17824,N_17998);
xor U18412 (N_18412,N_17603,N_17831);
nor U18413 (N_18413,N_17608,N_17799);
and U18414 (N_18414,N_17625,N_17751);
or U18415 (N_18415,N_17538,N_17744);
or U18416 (N_18416,N_17951,N_17854);
or U18417 (N_18417,N_17593,N_17826);
nor U18418 (N_18418,N_17647,N_17570);
and U18419 (N_18419,N_17853,N_17518);
nor U18420 (N_18420,N_17522,N_17604);
xnor U18421 (N_18421,N_17591,N_17531);
nor U18422 (N_18422,N_17821,N_17847);
xor U18423 (N_18423,N_17707,N_17603);
xnor U18424 (N_18424,N_17926,N_17988);
xnor U18425 (N_18425,N_17611,N_17718);
nor U18426 (N_18426,N_17523,N_17873);
and U18427 (N_18427,N_17865,N_17898);
and U18428 (N_18428,N_17759,N_17914);
nand U18429 (N_18429,N_17937,N_17596);
or U18430 (N_18430,N_17675,N_17660);
nor U18431 (N_18431,N_17976,N_17570);
xor U18432 (N_18432,N_17847,N_17738);
or U18433 (N_18433,N_17525,N_17738);
nor U18434 (N_18434,N_17968,N_17953);
nor U18435 (N_18435,N_17578,N_17812);
xor U18436 (N_18436,N_17713,N_17569);
or U18437 (N_18437,N_17942,N_17637);
nor U18438 (N_18438,N_17637,N_17722);
xor U18439 (N_18439,N_17693,N_17959);
and U18440 (N_18440,N_17923,N_17612);
or U18441 (N_18441,N_17803,N_17626);
and U18442 (N_18442,N_17500,N_17567);
xor U18443 (N_18443,N_17890,N_17744);
or U18444 (N_18444,N_17774,N_17561);
or U18445 (N_18445,N_17977,N_17777);
xor U18446 (N_18446,N_17990,N_17989);
or U18447 (N_18447,N_17662,N_17638);
xor U18448 (N_18448,N_17987,N_17976);
xor U18449 (N_18449,N_17813,N_17720);
xor U18450 (N_18450,N_17764,N_17545);
or U18451 (N_18451,N_17558,N_17815);
and U18452 (N_18452,N_17541,N_17778);
and U18453 (N_18453,N_17764,N_17971);
or U18454 (N_18454,N_17902,N_17574);
nor U18455 (N_18455,N_17921,N_17599);
nor U18456 (N_18456,N_17662,N_17986);
nor U18457 (N_18457,N_17510,N_17693);
nor U18458 (N_18458,N_17791,N_17534);
nor U18459 (N_18459,N_17827,N_17796);
nand U18460 (N_18460,N_17901,N_17871);
xnor U18461 (N_18461,N_17520,N_17706);
nand U18462 (N_18462,N_17856,N_17913);
nand U18463 (N_18463,N_17605,N_17803);
and U18464 (N_18464,N_17806,N_17846);
xnor U18465 (N_18465,N_17856,N_17634);
nor U18466 (N_18466,N_17950,N_17937);
xnor U18467 (N_18467,N_17551,N_17648);
xor U18468 (N_18468,N_17608,N_17865);
nand U18469 (N_18469,N_17800,N_17891);
or U18470 (N_18470,N_17841,N_17554);
nor U18471 (N_18471,N_17511,N_17745);
xnor U18472 (N_18472,N_17901,N_17926);
nor U18473 (N_18473,N_17923,N_17956);
nor U18474 (N_18474,N_17802,N_17915);
nor U18475 (N_18475,N_17941,N_17858);
and U18476 (N_18476,N_17908,N_17637);
nand U18477 (N_18477,N_17695,N_17874);
and U18478 (N_18478,N_17545,N_17712);
or U18479 (N_18479,N_17828,N_17969);
nor U18480 (N_18480,N_17717,N_17697);
nor U18481 (N_18481,N_17989,N_17695);
nand U18482 (N_18482,N_17886,N_17758);
and U18483 (N_18483,N_17741,N_17866);
nand U18484 (N_18484,N_17839,N_17837);
and U18485 (N_18485,N_17793,N_17648);
or U18486 (N_18486,N_17810,N_17843);
or U18487 (N_18487,N_17592,N_17871);
and U18488 (N_18488,N_17701,N_17696);
nor U18489 (N_18489,N_17868,N_17962);
nor U18490 (N_18490,N_17715,N_17909);
nand U18491 (N_18491,N_17913,N_17828);
or U18492 (N_18492,N_17836,N_17648);
nor U18493 (N_18493,N_17807,N_17767);
or U18494 (N_18494,N_17675,N_17732);
and U18495 (N_18495,N_17590,N_17522);
or U18496 (N_18496,N_17587,N_17632);
nand U18497 (N_18497,N_17657,N_17664);
nor U18498 (N_18498,N_17928,N_17722);
nor U18499 (N_18499,N_17822,N_17796);
nor U18500 (N_18500,N_18171,N_18039);
nand U18501 (N_18501,N_18016,N_18454);
nor U18502 (N_18502,N_18479,N_18348);
and U18503 (N_18503,N_18223,N_18188);
and U18504 (N_18504,N_18218,N_18117);
nand U18505 (N_18505,N_18014,N_18338);
or U18506 (N_18506,N_18419,N_18429);
xor U18507 (N_18507,N_18265,N_18167);
nand U18508 (N_18508,N_18090,N_18238);
nand U18509 (N_18509,N_18203,N_18376);
xnor U18510 (N_18510,N_18369,N_18333);
and U18511 (N_18511,N_18222,N_18433);
nor U18512 (N_18512,N_18032,N_18465);
and U18513 (N_18513,N_18396,N_18295);
or U18514 (N_18514,N_18066,N_18283);
or U18515 (N_18515,N_18056,N_18183);
or U18516 (N_18516,N_18097,N_18316);
nor U18517 (N_18517,N_18439,N_18389);
nor U18518 (N_18518,N_18064,N_18105);
xor U18519 (N_18519,N_18133,N_18289);
and U18520 (N_18520,N_18372,N_18052);
and U18521 (N_18521,N_18233,N_18401);
xnor U18522 (N_18522,N_18166,N_18494);
or U18523 (N_18523,N_18418,N_18451);
xnor U18524 (N_18524,N_18336,N_18147);
nand U18525 (N_18525,N_18434,N_18368);
nand U18526 (N_18526,N_18431,N_18214);
xnor U18527 (N_18527,N_18163,N_18426);
and U18528 (N_18528,N_18024,N_18319);
nand U18529 (N_18529,N_18402,N_18449);
or U18530 (N_18530,N_18006,N_18169);
nand U18531 (N_18531,N_18252,N_18130);
and U18532 (N_18532,N_18109,N_18428);
or U18533 (N_18533,N_18144,N_18269);
nor U18534 (N_18534,N_18351,N_18312);
nand U18535 (N_18535,N_18489,N_18152);
or U18536 (N_18536,N_18335,N_18080);
and U18537 (N_18537,N_18123,N_18255);
nand U18538 (N_18538,N_18161,N_18185);
xor U18539 (N_18539,N_18371,N_18422);
xnor U18540 (N_18540,N_18356,N_18370);
xnor U18541 (N_18541,N_18301,N_18060);
nand U18542 (N_18542,N_18287,N_18211);
nor U18543 (N_18543,N_18089,N_18044);
or U18544 (N_18544,N_18483,N_18087);
xor U18545 (N_18545,N_18137,N_18326);
xnor U18546 (N_18546,N_18436,N_18033);
xnor U18547 (N_18547,N_18325,N_18441);
nand U18548 (N_18548,N_18180,N_18456);
nand U18549 (N_18549,N_18308,N_18142);
nand U18550 (N_18550,N_18119,N_18047);
nand U18551 (N_18551,N_18225,N_18278);
or U18552 (N_18552,N_18069,N_18395);
xor U18553 (N_18553,N_18413,N_18377);
nor U18554 (N_18554,N_18084,N_18182);
xor U18555 (N_18555,N_18003,N_18186);
and U18556 (N_18556,N_18217,N_18317);
nor U18557 (N_18557,N_18010,N_18198);
or U18558 (N_18558,N_18281,N_18261);
xnor U18559 (N_18559,N_18030,N_18212);
nand U18560 (N_18560,N_18228,N_18096);
xnor U18561 (N_18561,N_18366,N_18264);
xnor U18562 (N_18562,N_18447,N_18239);
nor U18563 (N_18563,N_18143,N_18469);
nand U18564 (N_18564,N_18328,N_18048);
xnor U18565 (N_18565,N_18496,N_18165);
and U18566 (N_18566,N_18231,N_18002);
nor U18567 (N_18567,N_18288,N_18468);
nor U18568 (N_18568,N_18004,N_18135);
xor U18569 (N_18569,N_18086,N_18246);
nor U18570 (N_18570,N_18059,N_18303);
nand U18571 (N_18571,N_18474,N_18062);
nor U18572 (N_18572,N_18072,N_18248);
xnor U18573 (N_18573,N_18311,N_18394);
nand U18574 (N_18574,N_18018,N_18442);
or U18575 (N_18575,N_18029,N_18227);
or U18576 (N_18576,N_18355,N_18407);
nor U18577 (N_18577,N_18362,N_18365);
and U18578 (N_18578,N_18092,N_18124);
nand U18579 (N_18579,N_18001,N_18164);
nor U18580 (N_18580,N_18127,N_18388);
nand U18581 (N_18581,N_18153,N_18268);
xnor U18582 (N_18582,N_18297,N_18495);
xnor U18583 (N_18583,N_18277,N_18346);
or U18584 (N_18584,N_18076,N_18384);
nor U18585 (N_18585,N_18435,N_18463);
or U18586 (N_18586,N_18294,N_18196);
nor U18587 (N_18587,N_18458,N_18404);
or U18588 (N_18588,N_18329,N_18000);
and U18589 (N_18589,N_18154,N_18015);
xnor U18590 (N_18590,N_18050,N_18397);
and U18591 (N_18591,N_18156,N_18204);
nor U18592 (N_18592,N_18009,N_18412);
nand U18593 (N_18593,N_18405,N_18337);
and U18594 (N_18594,N_18199,N_18245);
or U18595 (N_18595,N_18149,N_18475);
xor U18596 (N_18596,N_18058,N_18162);
and U18597 (N_18597,N_18128,N_18031);
xnor U18598 (N_18598,N_18102,N_18041);
and U18599 (N_18599,N_18318,N_18221);
nand U18600 (N_18600,N_18381,N_18440);
nand U18601 (N_18601,N_18074,N_18497);
nand U18602 (N_18602,N_18061,N_18045);
or U18603 (N_18603,N_18379,N_18085);
or U18604 (N_18604,N_18067,N_18481);
nor U18605 (N_18605,N_18068,N_18181);
nor U18606 (N_18606,N_18464,N_18460);
nand U18607 (N_18607,N_18195,N_18499);
and U18608 (N_18608,N_18094,N_18417);
nor U18609 (N_18609,N_18172,N_18110);
xor U18610 (N_18610,N_18391,N_18487);
nand U18611 (N_18611,N_18380,N_18254);
xor U18612 (N_18612,N_18352,N_18423);
or U18613 (N_18613,N_18453,N_18491);
xor U18614 (N_18614,N_18293,N_18070);
nand U18615 (N_18615,N_18158,N_18408);
and U18616 (N_18616,N_18190,N_18274);
or U18617 (N_18617,N_18392,N_18339);
nand U18618 (N_18618,N_18490,N_18157);
or U18619 (N_18619,N_18266,N_18305);
nand U18620 (N_18620,N_18399,N_18359);
or U18621 (N_18621,N_18013,N_18091);
nor U18622 (N_18622,N_18034,N_18107);
nor U18623 (N_18623,N_18390,N_18035);
nand U18624 (N_18624,N_18358,N_18364);
xor U18625 (N_18625,N_18173,N_18321);
or U18626 (N_18626,N_18098,N_18310);
nor U18627 (N_18627,N_18350,N_18279);
nor U18628 (N_18628,N_18270,N_18267);
xnor U18629 (N_18629,N_18360,N_18208);
or U18630 (N_18630,N_18315,N_18020);
nor U18631 (N_18631,N_18324,N_18410);
or U18632 (N_18632,N_18249,N_18340);
and U18633 (N_18633,N_18151,N_18466);
xor U18634 (N_18634,N_18322,N_18409);
or U18635 (N_18635,N_18073,N_18046);
nand U18636 (N_18636,N_18411,N_18140);
xnor U18637 (N_18637,N_18282,N_18236);
xor U18638 (N_18638,N_18260,N_18242);
nor U18639 (N_18639,N_18375,N_18007);
or U18640 (N_18640,N_18403,N_18349);
nand U18641 (N_18641,N_18146,N_18189);
and U18642 (N_18642,N_18028,N_18353);
xnor U18643 (N_18643,N_18306,N_18296);
nand U18644 (N_18644,N_18229,N_18057);
or U18645 (N_18645,N_18065,N_18111);
or U18646 (N_18646,N_18226,N_18457);
nand U18647 (N_18647,N_18493,N_18421);
nor U18648 (N_18648,N_18284,N_18291);
nand U18649 (N_18649,N_18425,N_18159);
or U18650 (N_18650,N_18477,N_18343);
xor U18651 (N_18651,N_18443,N_18112);
nand U18652 (N_18652,N_18101,N_18027);
xor U18653 (N_18653,N_18472,N_18304);
nand U18654 (N_18654,N_18484,N_18176);
nand U18655 (N_18655,N_18290,N_18373);
nor U18656 (N_18656,N_18342,N_18250);
xnor U18657 (N_18657,N_18385,N_18197);
or U18658 (N_18658,N_18095,N_18202);
nand U18659 (N_18659,N_18235,N_18077);
xnor U18660 (N_18660,N_18093,N_18141);
and U18661 (N_18661,N_18448,N_18113);
and U18662 (N_18662,N_18285,N_18446);
xnor U18663 (N_18663,N_18302,N_18415);
or U18664 (N_18664,N_18482,N_18406);
and U18665 (N_18665,N_18374,N_18055);
and U18666 (N_18666,N_18271,N_18416);
nand U18667 (N_18667,N_18115,N_18462);
or U18668 (N_18668,N_18191,N_18131);
nor U18669 (N_18669,N_18378,N_18083);
xor U18670 (N_18670,N_18126,N_18139);
xor U18671 (N_18671,N_18054,N_18344);
xor U18672 (N_18672,N_18021,N_18082);
xnor U18673 (N_18673,N_18104,N_18470);
or U18674 (N_18674,N_18262,N_18367);
nand U18675 (N_18675,N_18053,N_18253);
and U18676 (N_18676,N_18251,N_18275);
nand U18677 (N_18677,N_18129,N_18243);
and U18678 (N_18678,N_18420,N_18108);
xor U18679 (N_18679,N_18177,N_18008);
or U18680 (N_18680,N_18363,N_18452);
or U18681 (N_18681,N_18219,N_18272);
nor U18682 (N_18682,N_18256,N_18134);
nand U18683 (N_18683,N_18184,N_18387);
nor U18684 (N_18684,N_18049,N_18476);
nand U18685 (N_18685,N_18323,N_18237);
and U18686 (N_18686,N_18320,N_18026);
nand U18687 (N_18687,N_18234,N_18232);
and U18688 (N_18688,N_18150,N_18230);
xnor U18689 (N_18689,N_18445,N_18259);
xor U18690 (N_18690,N_18012,N_18179);
nor U18691 (N_18691,N_18071,N_18201);
and U18692 (N_18692,N_18307,N_18492);
xnor U18693 (N_18693,N_18040,N_18118);
xnor U18694 (N_18694,N_18099,N_18168);
nor U18695 (N_18695,N_18148,N_18430);
xnor U18696 (N_18696,N_18498,N_18078);
or U18697 (N_18697,N_18206,N_18063);
or U18698 (N_18698,N_18400,N_18486);
nor U18699 (N_18699,N_18037,N_18299);
xnor U18700 (N_18700,N_18332,N_18100);
or U18701 (N_18701,N_18081,N_18438);
nor U18702 (N_18702,N_18247,N_18025);
nor U18703 (N_18703,N_18088,N_18357);
xor U18704 (N_18704,N_18075,N_18210);
and U18705 (N_18705,N_18314,N_18309);
and U18706 (N_18706,N_18478,N_18215);
nand U18707 (N_18707,N_18361,N_18145);
xor U18708 (N_18708,N_18038,N_18444);
and U18709 (N_18709,N_18042,N_18213);
nand U18710 (N_18710,N_18398,N_18175);
or U18711 (N_18711,N_18459,N_18488);
nand U18712 (N_18712,N_18286,N_18313);
or U18713 (N_18713,N_18480,N_18216);
xnor U18714 (N_18714,N_18432,N_18138);
xor U18715 (N_18715,N_18292,N_18178);
and U18716 (N_18716,N_18414,N_18122);
nand U18717 (N_18717,N_18194,N_18187);
or U18718 (N_18718,N_18393,N_18280);
nor U18719 (N_18719,N_18022,N_18192);
or U18720 (N_18720,N_18258,N_18136);
nor U18721 (N_18721,N_18036,N_18354);
nand U18722 (N_18722,N_18116,N_18386);
or U18723 (N_18723,N_18079,N_18455);
or U18724 (N_18724,N_18011,N_18170);
and U18725 (N_18725,N_18341,N_18120);
and U18726 (N_18726,N_18257,N_18174);
nor U18727 (N_18727,N_18132,N_18019);
and U18728 (N_18728,N_18334,N_18017);
xor U18729 (N_18729,N_18114,N_18347);
or U18730 (N_18730,N_18005,N_18155);
and U18731 (N_18731,N_18023,N_18160);
xor U18732 (N_18732,N_18471,N_18331);
or U18733 (N_18733,N_18200,N_18106);
and U18734 (N_18734,N_18485,N_18437);
xor U18735 (N_18735,N_18121,N_18051);
nand U18736 (N_18736,N_18327,N_18244);
nor U18737 (N_18737,N_18240,N_18276);
nor U18738 (N_18738,N_18263,N_18424);
nand U18739 (N_18739,N_18450,N_18383);
nand U18740 (N_18740,N_18467,N_18473);
nor U18741 (N_18741,N_18224,N_18193);
xnor U18742 (N_18742,N_18427,N_18330);
nor U18743 (N_18743,N_18300,N_18205);
and U18744 (N_18744,N_18209,N_18241);
nand U18745 (N_18745,N_18043,N_18207);
and U18746 (N_18746,N_18298,N_18345);
nand U18747 (N_18747,N_18273,N_18461);
and U18748 (N_18748,N_18382,N_18125);
and U18749 (N_18749,N_18103,N_18220);
and U18750 (N_18750,N_18025,N_18139);
nand U18751 (N_18751,N_18319,N_18467);
nand U18752 (N_18752,N_18152,N_18304);
nor U18753 (N_18753,N_18393,N_18193);
nand U18754 (N_18754,N_18008,N_18036);
and U18755 (N_18755,N_18012,N_18424);
xor U18756 (N_18756,N_18279,N_18454);
nor U18757 (N_18757,N_18011,N_18118);
xor U18758 (N_18758,N_18069,N_18458);
nand U18759 (N_18759,N_18486,N_18426);
xor U18760 (N_18760,N_18397,N_18095);
xor U18761 (N_18761,N_18291,N_18120);
xnor U18762 (N_18762,N_18380,N_18176);
or U18763 (N_18763,N_18492,N_18152);
nand U18764 (N_18764,N_18079,N_18118);
or U18765 (N_18765,N_18168,N_18198);
xor U18766 (N_18766,N_18011,N_18042);
or U18767 (N_18767,N_18285,N_18255);
and U18768 (N_18768,N_18281,N_18489);
or U18769 (N_18769,N_18194,N_18149);
nand U18770 (N_18770,N_18266,N_18075);
and U18771 (N_18771,N_18019,N_18309);
nor U18772 (N_18772,N_18264,N_18110);
and U18773 (N_18773,N_18109,N_18274);
or U18774 (N_18774,N_18115,N_18441);
nor U18775 (N_18775,N_18356,N_18277);
or U18776 (N_18776,N_18234,N_18480);
xnor U18777 (N_18777,N_18247,N_18219);
or U18778 (N_18778,N_18424,N_18005);
xnor U18779 (N_18779,N_18062,N_18490);
nor U18780 (N_18780,N_18460,N_18272);
or U18781 (N_18781,N_18022,N_18368);
nand U18782 (N_18782,N_18374,N_18490);
and U18783 (N_18783,N_18242,N_18343);
and U18784 (N_18784,N_18257,N_18417);
nand U18785 (N_18785,N_18400,N_18206);
nor U18786 (N_18786,N_18231,N_18422);
xnor U18787 (N_18787,N_18261,N_18413);
nand U18788 (N_18788,N_18114,N_18272);
xnor U18789 (N_18789,N_18036,N_18454);
or U18790 (N_18790,N_18310,N_18487);
nand U18791 (N_18791,N_18316,N_18399);
nand U18792 (N_18792,N_18296,N_18331);
or U18793 (N_18793,N_18278,N_18460);
nor U18794 (N_18794,N_18472,N_18048);
nor U18795 (N_18795,N_18375,N_18407);
nor U18796 (N_18796,N_18374,N_18426);
and U18797 (N_18797,N_18071,N_18471);
nand U18798 (N_18798,N_18249,N_18207);
nor U18799 (N_18799,N_18083,N_18346);
nand U18800 (N_18800,N_18290,N_18297);
xnor U18801 (N_18801,N_18084,N_18069);
nand U18802 (N_18802,N_18192,N_18416);
or U18803 (N_18803,N_18016,N_18040);
nand U18804 (N_18804,N_18439,N_18013);
or U18805 (N_18805,N_18479,N_18175);
xnor U18806 (N_18806,N_18032,N_18237);
nand U18807 (N_18807,N_18439,N_18184);
nand U18808 (N_18808,N_18113,N_18479);
and U18809 (N_18809,N_18025,N_18382);
nor U18810 (N_18810,N_18408,N_18388);
nor U18811 (N_18811,N_18491,N_18168);
nor U18812 (N_18812,N_18166,N_18452);
xnor U18813 (N_18813,N_18094,N_18264);
nor U18814 (N_18814,N_18251,N_18165);
nand U18815 (N_18815,N_18167,N_18401);
and U18816 (N_18816,N_18017,N_18353);
or U18817 (N_18817,N_18150,N_18292);
xor U18818 (N_18818,N_18069,N_18189);
xor U18819 (N_18819,N_18365,N_18263);
nor U18820 (N_18820,N_18348,N_18386);
xnor U18821 (N_18821,N_18060,N_18297);
nor U18822 (N_18822,N_18492,N_18216);
nand U18823 (N_18823,N_18293,N_18080);
or U18824 (N_18824,N_18208,N_18473);
nor U18825 (N_18825,N_18184,N_18030);
nand U18826 (N_18826,N_18470,N_18445);
or U18827 (N_18827,N_18112,N_18001);
nor U18828 (N_18828,N_18308,N_18458);
or U18829 (N_18829,N_18174,N_18070);
nor U18830 (N_18830,N_18037,N_18449);
or U18831 (N_18831,N_18188,N_18234);
xnor U18832 (N_18832,N_18082,N_18273);
nand U18833 (N_18833,N_18473,N_18064);
and U18834 (N_18834,N_18472,N_18175);
or U18835 (N_18835,N_18296,N_18481);
nand U18836 (N_18836,N_18149,N_18307);
nand U18837 (N_18837,N_18371,N_18145);
nand U18838 (N_18838,N_18188,N_18054);
or U18839 (N_18839,N_18312,N_18107);
and U18840 (N_18840,N_18109,N_18414);
nor U18841 (N_18841,N_18370,N_18186);
nor U18842 (N_18842,N_18440,N_18212);
xnor U18843 (N_18843,N_18414,N_18317);
xor U18844 (N_18844,N_18442,N_18343);
or U18845 (N_18845,N_18298,N_18295);
or U18846 (N_18846,N_18019,N_18417);
xor U18847 (N_18847,N_18034,N_18357);
and U18848 (N_18848,N_18174,N_18016);
and U18849 (N_18849,N_18232,N_18226);
and U18850 (N_18850,N_18223,N_18306);
nor U18851 (N_18851,N_18215,N_18458);
and U18852 (N_18852,N_18437,N_18438);
nand U18853 (N_18853,N_18344,N_18226);
or U18854 (N_18854,N_18206,N_18460);
and U18855 (N_18855,N_18271,N_18431);
nor U18856 (N_18856,N_18290,N_18378);
and U18857 (N_18857,N_18027,N_18116);
xor U18858 (N_18858,N_18408,N_18005);
or U18859 (N_18859,N_18265,N_18450);
and U18860 (N_18860,N_18031,N_18117);
nand U18861 (N_18861,N_18445,N_18472);
or U18862 (N_18862,N_18454,N_18293);
nand U18863 (N_18863,N_18486,N_18307);
nor U18864 (N_18864,N_18357,N_18295);
or U18865 (N_18865,N_18055,N_18310);
and U18866 (N_18866,N_18019,N_18061);
nor U18867 (N_18867,N_18353,N_18435);
nor U18868 (N_18868,N_18286,N_18141);
nand U18869 (N_18869,N_18202,N_18384);
nand U18870 (N_18870,N_18208,N_18264);
nand U18871 (N_18871,N_18160,N_18112);
xor U18872 (N_18872,N_18151,N_18113);
nand U18873 (N_18873,N_18164,N_18103);
nand U18874 (N_18874,N_18145,N_18075);
nor U18875 (N_18875,N_18163,N_18199);
xnor U18876 (N_18876,N_18117,N_18429);
nand U18877 (N_18877,N_18323,N_18136);
nor U18878 (N_18878,N_18279,N_18403);
xor U18879 (N_18879,N_18297,N_18283);
nor U18880 (N_18880,N_18226,N_18288);
or U18881 (N_18881,N_18183,N_18284);
nand U18882 (N_18882,N_18091,N_18142);
xor U18883 (N_18883,N_18088,N_18163);
xnor U18884 (N_18884,N_18069,N_18225);
xor U18885 (N_18885,N_18233,N_18032);
xor U18886 (N_18886,N_18385,N_18182);
xnor U18887 (N_18887,N_18228,N_18322);
or U18888 (N_18888,N_18289,N_18217);
xnor U18889 (N_18889,N_18057,N_18270);
xor U18890 (N_18890,N_18363,N_18427);
or U18891 (N_18891,N_18230,N_18019);
or U18892 (N_18892,N_18181,N_18339);
or U18893 (N_18893,N_18456,N_18173);
xnor U18894 (N_18894,N_18352,N_18187);
or U18895 (N_18895,N_18389,N_18086);
or U18896 (N_18896,N_18454,N_18329);
xor U18897 (N_18897,N_18176,N_18345);
nor U18898 (N_18898,N_18091,N_18084);
nor U18899 (N_18899,N_18182,N_18496);
nand U18900 (N_18900,N_18109,N_18156);
nand U18901 (N_18901,N_18118,N_18444);
or U18902 (N_18902,N_18093,N_18169);
nand U18903 (N_18903,N_18075,N_18073);
nand U18904 (N_18904,N_18320,N_18369);
or U18905 (N_18905,N_18211,N_18246);
nand U18906 (N_18906,N_18044,N_18109);
or U18907 (N_18907,N_18443,N_18380);
xnor U18908 (N_18908,N_18119,N_18188);
nor U18909 (N_18909,N_18012,N_18322);
xor U18910 (N_18910,N_18258,N_18268);
xor U18911 (N_18911,N_18475,N_18088);
xor U18912 (N_18912,N_18393,N_18489);
nand U18913 (N_18913,N_18163,N_18181);
nand U18914 (N_18914,N_18233,N_18362);
xor U18915 (N_18915,N_18390,N_18359);
nand U18916 (N_18916,N_18245,N_18131);
and U18917 (N_18917,N_18449,N_18088);
nor U18918 (N_18918,N_18295,N_18356);
nand U18919 (N_18919,N_18342,N_18041);
nand U18920 (N_18920,N_18196,N_18088);
xor U18921 (N_18921,N_18347,N_18445);
xor U18922 (N_18922,N_18143,N_18020);
and U18923 (N_18923,N_18485,N_18023);
and U18924 (N_18924,N_18168,N_18424);
xor U18925 (N_18925,N_18385,N_18471);
nand U18926 (N_18926,N_18454,N_18072);
nand U18927 (N_18927,N_18157,N_18228);
nand U18928 (N_18928,N_18464,N_18218);
or U18929 (N_18929,N_18276,N_18130);
or U18930 (N_18930,N_18481,N_18253);
nand U18931 (N_18931,N_18071,N_18062);
nand U18932 (N_18932,N_18303,N_18251);
nand U18933 (N_18933,N_18304,N_18455);
nand U18934 (N_18934,N_18150,N_18497);
or U18935 (N_18935,N_18356,N_18367);
nor U18936 (N_18936,N_18479,N_18153);
nor U18937 (N_18937,N_18018,N_18134);
nor U18938 (N_18938,N_18161,N_18096);
xor U18939 (N_18939,N_18280,N_18358);
and U18940 (N_18940,N_18070,N_18362);
or U18941 (N_18941,N_18456,N_18288);
and U18942 (N_18942,N_18282,N_18486);
nor U18943 (N_18943,N_18273,N_18180);
nor U18944 (N_18944,N_18239,N_18110);
and U18945 (N_18945,N_18120,N_18343);
nand U18946 (N_18946,N_18159,N_18409);
nand U18947 (N_18947,N_18234,N_18036);
nand U18948 (N_18948,N_18072,N_18275);
nor U18949 (N_18949,N_18057,N_18477);
or U18950 (N_18950,N_18417,N_18176);
and U18951 (N_18951,N_18436,N_18387);
xor U18952 (N_18952,N_18181,N_18344);
nor U18953 (N_18953,N_18060,N_18459);
xor U18954 (N_18954,N_18461,N_18497);
xor U18955 (N_18955,N_18216,N_18040);
or U18956 (N_18956,N_18381,N_18143);
nor U18957 (N_18957,N_18438,N_18073);
xor U18958 (N_18958,N_18416,N_18378);
and U18959 (N_18959,N_18254,N_18436);
and U18960 (N_18960,N_18419,N_18170);
nor U18961 (N_18961,N_18021,N_18490);
nand U18962 (N_18962,N_18058,N_18118);
nor U18963 (N_18963,N_18429,N_18317);
nor U18964 (N_18964,N_18114,N_18235);
nand U18965 (N_18965,N_18317,N_18154);
nand U18966 (N_18966,N_18493,N_18377);
nand U18967 (N_18967,N_18176,N_18493);
nor U18968 (N_18968,N_18429,N_18363);
nor U18969 (N_18969,N_18209,N_18136);
nor U18970 (N_18970,N_18367,N_18499);
nor U18971 (N_18971,N_18432,N_18082);
or U18972 (N_18972,N_18268,N_18287);
and U18973 (N_18973,N_18085,N_18055);
xnor U18974 (N_18974,N_18038,N_18212);
nand U18975 (N_18975,N_18044,N_18354);
nor U18976 (N_18976,N_18253,N_18250);
and U18977 (N_18977,N_18275,N_18304);
xnor U18978 (N_18978,N_18031,N_18434);
nor U18979 (N_18979,N_18248,N_18054);
nor U18980 (N_18980,N_18450,N_18010);
nor U18981 (N_18981,N_18180,N_18335);
and U18982 (N_18982,N_18309,N_18052);
nand U18983 (N_18983,N_18277,N_18303);
nand U18984 (N_18984,N_18144,N_18258);
xor U18985 (N_18985,N_18162,N_18046);
and U18986 (N_18986,N_18137,N_18023);
nand U18987 (N_18987,N_18201,N_18229);
or U18988 (N_18988,N_18071,N_18229);
or U18989 (N_18989,N_18093,N_18274);
xor U18990 (N_18990,N_18130,N_18209);
and U18991 (N_18991,N_18306,N_18327);
or U18992 (N_18992,N_18074,N_18362);
xor U18993 (N_18993,N_18232,N_18363);
xnor U18994 (N_18994,N_18074,N_18111);
or U18995 (N_18995,N_18465,N_18108);
xnor U18996 (N_18996,N_18035,N_18043);
xor U18997 (N_18997,N_18200,N_18030);
nor U18998 (N_18998,N_18460,N_18443);
nor U18999 (N_18999,N_18341,N_18441);
and U19000 (N_19000,N_18633,N_18763);
and U19001 (N_19001,N_18671,N_18949);
and U19002 (N_19002,N_18872,N_18675);
and U19003 (N_19003,N_18814,N_18863);
and U19004 (N_19004,N_18860,N_18909);
or U19005 (N_19005,N_18648,N_18977);
xor U19006 (N_19006,N_18843,N_18870);
nor U19007 (N_19007,N_18713,N_18947);
and U19008 (N_19008,N_18710,N_18901);
nand U19009 (N_19009,N_18862,N_18958);
nand U19010 (N_19010,N_18845,N_18748);
nor U19011 (N_19011,N_18795,N_18935);
nor U19012 (N_19012,N_18698,N_18720);
nand U19013 (N_19013,N_18667,N_18782);
nor U19014 (N_19014,N_18867,N_18746);
or U19015 (N_19015,N_18767,N_18712);
and U19016 (N_19016,N_18547,N_18598);
or U19017 (N_19017,N_18809,N_18786);
xor U19018 (N_19018,N_18808,N_18605);
and U19019 (N_19019,N_18785,N_18573);
and U19020 (N_19020,N_18695,N_18575);
nor U19021 (N_19021,N_18638,N_18537);
nor U19022 (N_19022,N_18742,N_18706);
and U19023 (N_19023,N_18662,N_18516);
xnor U19024 (N_19024,N_18738,N_18597);
and U19025 (N_19025,N_18511,N_18697);
nor U19026 (N_19026,N_18716,N_18915);
xnor U19027 (N_19027,N_18812,N_18770);
and U19028 (N_19028,N_18571,N_18664);
or U19029 (N_19029,N_18944,N_18688);
xnor U19030 (N_19030,N_18635,N_18801);
and U19031 (N_19031,N_18848,N_18868);
nor U19032 (N_19032,N_18779,N_18853);
or U19033 (N_19033,N_18881,N_18778);
nor U19034 (N_19034,N_18834,N_18832);
nand U19035 (N_19035,N_18890,N_18956);
and U19036 (N_19036,N_18941,N_18887);
or U19037 (N_19037,N_18888,N_18608);
and U19038 (N_19038,N_18623,N_18886);
and U19039 (N_19039,N_18772,N_18762);
nand U19040 (N_19040,N_18907,N_18620);
nor U19041 (N_19041,N_18517,N_18589);
nor U19042 (N_19042,N_18936,N_18681);
nor U19043 (N_19043,N_18963,N_18611);
or U19044 (N_19044,N_18578,N_18747);
xnor U19045 (N_19045,N_18728,N_18616);
nor U19046 (N_19046,N_18727,N_18789);
nor U19047 (N_19047,N_18669,N_18854);
nor U19048 (N_19048,N_18594,N_18980);
nand U19049 (N_19049,N_18668,N_18791);
or U19050 (N_19050,N_18810,N_18799);
xor U19051 (N_19051,N_18714,N_18976);
nor U19052 (N_19052,N_18521,N_18736);
nand U19053 (N_19053,N_18683,N_18904);
nor U19054 (N_19054,N_18550,N_18565);
nand U19055 (N_19055,N_18548,N_18524);
nand U19056 (N_19056,N_18940,N_18817);
nor U19057 (N_19057,N_18532,N_18583);
nor U19058 (N_19058,N_18806,N_18942);
nor U19059 (N_19059,N_18892,N_18570);
or U19060 (N_19060,N_18512,N_18733);
or U19061 (N_19061,N_18766,N_18829);
and U19062 (N_19062,N_18566,N_18735);
xnor U19063 (N_19063,N_18593,N_18588);
or U19064 (N_19064,N_18614,N_18562);
xnor U19065 (N_19065,N_18555,N_18678);
or U19066 (N_19066,N_18509,N_18750);
or U19067 (N_19067,N_18626,N_18811);
nor U19068 (N_19068,N_18918,N_18549);
or U19069 (N_19069,N_18525,N_18676);
nand U19070 (N_19070,N_18670,N_18705);
or U19071 (N_19071,N_18531,N_18897);
or U19072 (N_19072,N_18729,N_18579);
nand U19073 (N_19073,N_18663,N_18928);
or U19074 (N_19074,N_18787,N_18953);
or U19075 (N_19075,N_18592,N_18938);
nand U19076 (N_19076,N_18696,N_18653);
and U19077 (N_19077,N_18715,N_18986);
nand U19078 (N_19078,N_18534,N_18798);
nor U19079 (N_19079,N_18687,N_18518);
xor U19080 (N_19080,N_18866,N_18777);
or U19081 (N_19081,N_18691,N_18576);
nand U19082 (N_19082,N_18841,N_18711);
xnor U19083 (N_19083,N_18679,N_18725);
nand U19084 (N_19084,N_18722,N_18768);
or U19085 (N_19085,N_18931,N_18970);
and U19086 (N_19086,N_18837,N_18873);
and U19087 (N_19087,N_18959,N_18783);
nor U19088 (N_19088,N_18718,N_18739);
nor U19089 (N_19089,N_18939,N_18558);
or U19090 (N_19090,N_18932,N_18503);
nor U19091 (N_19091,N_18730,N_18895);
and U19092 (N_19092,N_18629,N_18969);
or U19093 (N_19093,N_18618,N_18621);
or U19094 (N_19094,N_18526,N_18924);
or U19095 (N_19095,N_18771,N_18615);
and U19096 (N_19096,N_18673,N_18946);
and U19097 (N_19097,N_18846,N_18794);
or U19098 (N_19098,N_18535,N_18805);
nand U19099 (N_19099,N_18833,N_18514);
or U19100 (N_19100,N_18553,N_18913);
or U19101 (N_19101,N_18822,N_18726);
and U19102 (N_19102,N_18709,N_18585);
nor U19103 (N_19103,N_18978,N_18916);
xor U19104 (N_19104,N_18745,N_18646);
nor U19105 (N_19105,N_18689,N_18922);
nor U19106 (N_19106,N_18855,N_18917);
xnor U19107 (N_19107,N_18654,N_18802);
and U19108 (N_19108,N_18741,N_18984);
or U19109 (N_19109,N_18876,N_18912);
and U19110 (N_19110,N_18828,N_18641);
nand U19111 (N_19111,N_18820,N_18607);
or U19112 (N_19112,N_18983,N_18647);
xor U19113 (N_19113,N_18744,N_18769);
xnor U19114 (N_19114,N_18965,N_18634);
nor U19115 (N_19115,N_18545,N_18755);
and U19116 (N_19116,N_18879,N_18797);
or U19117 (N_19117,N_18985,N_18740);
nand U19118 (N_19118,N_18898,N_18560);
nand U19119 (N_19119,N_18813,N_18754);
and U19120 (N_19120,N_18827,N_18905);
nand U19121 (N_19121,N_18586,N_18721);
nand U19122 (N_19122,N_18567,N_18650);
nor U19123 (N_19123,N_18559,N_18756);
and U19124 (N_19124,N_18930,N_18657);
or U19125 (N_19125,N_18502,N_18536);
or U19126 (N_19126,N_18758,N_18911);
and U19127 (N_19127,N_18604,N_18776);
xnor U19128 (N_19128,N_18875,N_18825);
nand U19129 (N_19129,N_18974,N_18600);
nand U19130 (N_19130,N_18541,N_18617);
nand U19131 (N_19131,N_18851,N_18666);
and U19132 (N_19132,N_18856,N_18816);
nor U19133 (N_19133,N_18753,N_18543);
or U19134 (N_19134,N_18554,N_18577);
nor U19135 (N_19135,N_18765,N_18665);
xnor U19136 (N_19136,N_18551,N_18831);
and U19137 (N_19137,N_18950,N_18864);
or U19138 (N_19138,N_18520,N_18569);
nand U19139 (N_19139,N_18542,N_18538);
or U19140 (N_19140,N_18702,N_18973);
or U19141 (N_19141,N_18590,N_18780);
nor U19142 (N_19142,N_18724,N_18743);
and U19143 (N_19143,N_18639,N_18943);
and U19144 (N_19144,N_18557,N_18530);
and U19145 (N_19145,N_18672,N_18500);
or U19146 (N_19146,N_18891,N_18640);
and U19147 (N_19147,N_18644,N_18906);
and U19148 (N_19148,N_18800,N_18998);
and U19149 (N_19149,N_18656,N_18539);
or U19150 (N_19150,N_18850,N_18572);
nor U19151 (N_19151,N_18835,N_18723);
xor U19152 (N_19152,N_18749,N_18921);
and U19153 (N_19153,N_18540,N_18752);
xnor U19154 (N_19154,N_18630,N_18877);
or U19155 (N_19155,N_18510,N_18582);
or U19156 (N_19156,N_18584,N_18788);
nand U19157 (N_19157,N_18775,N_18849);
nor U19158 (N_19158,N_18859,N_18732);
and U19159 (N_19159,N_18994,N_18926);
nand U19160 (N_19160,N_18948,N_18708);
nand U19161 (N_19161,N_18601,N_18910);
or U19162 (N_19162,N_18568,N_18880);
nor U19163 (N_19163,N_18587,N_18636);
nor U19164 (N_19164,N_18903,N_18971);
nand U19165 (N_19165,N_18818,N_18684);
xnor U19166 (N_19166,N_18527,N_18734);
or U19167 (N_19167,N_18761,N_18842);
xor U19168 (N_19168,N_18836,N_18964);
nor U19169 (N_19169,N_18929,N_18899);
and U19170 (N_19170,N_18645,N_18528);
and U19171 (N_19171,N_18519,N_18627);
nand U19172 (N_19172,N_18649,N_18882);
nand U19173 (N_19173,N_18642,N_18945);
xnor U19174 (N_19174,N_18505,N_18612);
nand U19175 (N_19175,N_18865,N_18619);
nor U19176 (N_19176,N_18692,N_18564);
xor U19177 (N_19177,N_18599,N_18680);
xor U19178 (N_19178,N_18651,N_18933);
or U19179 (N_19179,N_18591,N_18815);
nand U19180 (N_19180,N_18632,N_18504);
or U19181 (N_19181,N_18751,N_18596);
and U19182 (N_19182,N_18717,N_18966);
nor U19183 (N_19183,N_18513,N_18919);
xnor U19184 (N_19184,N_18937,N_18580);
xnor U19185 (N_19185,N_18603,N_18613);
and U19186 (N_19186,N_18652,N_18852);
nor U19187 (N_19187,N_18803,N_18914);
nand U19188 (N_19188,N_18685,N_18804);
or U19189 (N_19189,N_18990,N_18838);
or U19190 (N_19190,N_18896,N_18796);
and U19191 (N_19191,N_18823,N_18523);
xor U19192 (N_19192,N_18871,N_18561);
nand U19193 (N_19193,N_18840,N_18900);
and U19194 (N_19194,N_18699,N_18830);
nor U19195 (N_19195,N_18508,N_18552);
xor U19196 (N_19196,N_18658,N_18624);
nor U19197 (N_19197,N_18764,N_18923);
or U19198 (N_19198,N_18847,N_18884);
or U19199 (N_19199,N_18883,N_18979);
and U19200 (N_19200,N_18694,N_18686);
or U19201 (N_19201,N_18622,N_18957);
nor U19202 (N_19202,N_18701,N_18874);
and U19203 (N_19203,N_18507,N_18628);
and U19204 (N_19204,N_18774,N_18975);
nor U19205 (N_19205,N_18556,N_18533);
nor U19206 (N_19206,N_18858,N_18757);
nor U19207 (N_19207,N_18595,N_18824);
nand U19208 (N_19208,N_18988,N_18889);
xnor U19209 (N_19209,N_18581,N_18826);
and U19210 (N_19210,N_18819,N_18703);
or U19211 (N_19211,N_18606,N_18661);
and U19212 (N_19212,N_18704,N_18643);
and U19213 (N_19213,N_18677,N_18544);
xor U19214 (N_19214,N_18885,N_18999);
nor U19215 (N_19215,N_18737,N_18790);
and U19216 (N_19216,N_18807,N_18515);
or U19217 (N_19217,N_18972,N_18878);
or U19218 (N_19218,N_18574,N_18682);
nor U19219 (N_19219,N_18719,N_18960);
xnor U19220 (N_19220,N_18690,N_18968);
or U19221 (N_19221,N_18792,N_18955);
nor U19222 (N_19222,N_18773,N_18821);
or U19223 (N_19223,N_18610,N_18951);
or U19224 (N_19224,N_18700,N_18693);
nand U19225 (N_19225,N_18659,N_18961);
or U19226 (N_19226,N_18996,N_18707);
nand U19227 (N_19227,N_18637,N_18869);
nor U19228 (N_19228,N_18546,N_18927);
xor U19229 (N_19229,N_18674,N_18631);
nor U19230 (N_19230,N_18781,N_18908);
and U19231 (N_19231,N_18925,N_18655);
and U19232 (N_19232,N_18844,N_18893);
xor U19233 (N_19233,N_18759,N_18660);
nand U19234 (N_19234,N_18760,N_18952);
or U19235 (N_19235,N_18506,N_18987);
and U19236 (N_19236,N_18967,N_18920);
nor U19237 (N_19237,N_18625,N_18991);
and U19238 (N_19238,N_18563,N_18995);
nand U19239 (N_19239,N_18954,N_18793);
nor U19240 (N_19240,N_18609,N_18731);
nor U19241 (N_19241,N_18992,N_18894);
and U19242 (N_19242,N_18902,N_18989);
or U19243 (N_19243,N_18529,N_18962);
nor U19244 (N_19244,N_18522,N_18997);
nand U19245 (N_19245,N_18839,N_18934);
or U19246 (N_19246,N_18981,N_18784);
nand U19247 (N_19247,N_18993,N_18982);
and U19248 (N_19248,N_18602,N_18861);
nand U19249 (N_19249,N_18857,N_18501);
xor U19250 (N_19250,N_18782,N_18764);
nand U19251 (N_19251,N_18735,N_18792);
xnor U19252 (N_19252,N_18574,N_18941);
or U19253 (N_19253,N_18916,N_18945);
and U19254 (N_19254,N_18573,N_18921);
xor U19255 (N_19255,N_18786,N_18992);
or U19256 (N_19256,N_18513,N_18654);
or U19257 (N_19257,N_18731,N_18944);
and U19258 (N_19258,N_18558,N_18820);
or U19259 (N_19259,N_18861,N_18681);
nor U19260 (N_19260,N_18546,N_18705);
or U19261 (N_19261,N_18996,N_18522);
xor U19262 (N_19262,N_18979,N_18843);
nand U19263 (N_19263,N_18578,N_18504);
nor U19264 (N_19264,N_18778,N_18722);
and U19265 (N_19265,N_18616,N_18722);
xnor U19266 (N_19266,N_18753,N_18556);
xnor U19267 (N_19267,N_18905,N_18999);
nand U19268 (N_19268,N_18915,N_18717);
and U19269 (N_19269,N_18923,N_18688);
xor U19270 (N_19270,N_18591,N_18618);
and U19271 (N_19271,N_18798,N_18647);
nor U19272 (N_19272,N_18783,N_18842);
xor U19273 (N_19273,N_18642,N_18641);
xnor U19274 (N_19274,N_18510,N_18976);
nand U19275 (N_19275,N_18931,N_18705);
nor U19276 (N_19276,N_18567,N_18759);
nor U19277 (N_19277,N_18657,N_18900);
xnor U19278 (N_19278,N_18858,N_18971);
or U19279 (N_19279,N_18935,N_18841);
nor U19280 (N_19280,N_18503,N_18872);
or U19281 (N_19281,N_18931,N_18541);
xor U19282 (N_19282,N_18941,N_18856);
xor U19283 (N_19283,N_18527,N_18825);
or U19284 (N_19284,N_18970,N_18514);
and U19285 (N_19285,N_18615,N_18783);
and U19286 (N_19286,N_18542,N_18913);
and U19287 (N_19287,N_18897,N_18802);
xor U19288 (N_19288,N_18948,N_18592);
nand U19289 (N_19289,N_18642,N_18778);
and U19290 (N_19290,N_18591,N_18977);
nand U19291 (N_19291,N_18926,N_18864);
nand U19292 (N_19292,N_18775,N_18632);
and U19293 (N_19293,N_18814,N_18833);
and U19294 (N_19294,N_18947,N_18842);
nor U19295 (N_19295,N_18589,N_18663);
xnor U19296 (N_19296,N_18733,N_18549);
or U19297 (N_19297,N_18768,N_18547);
and U19298 (N_19298,N_18550,N_18539);
xnor U19299 (N_19299,N_18940,N_18687);
nor U19300 (N_19300,N_18652,N_18612);
and U19301 (N_19301,N_18723,N_18742);
or U19302 (N_19302,N_18731,N_18856);
nor U19303 (N_19303,N_18648,N_18580);
xor U19304 (N_19304,N_18808,N_18600);
xor U19305 (N_19305,N_18931,N_18788);
and U19306 (N_19306,N_18981,N_18944);
xor U19307 (N_19307,N_18999,N_18679);
xor U19308 (N_19308,N_18512,N_18567);
xnor U19309 (N_19309,N_18599,N_18769);
or U19310 (N_19310,N_18756,N_18886);
xnor U19311 (N_19311,N_18887,N_18726);
xnor U19312 (N_19312,N_18689,N_18559);
nand U19313 (N_19313,N_18704,N_18708);
xnor U19314 (N_19314,N_18555,N_18511);
xnor U19315 (N_19315,N_18656,N_18561);
and U19316 (N_19316,N_18547,N_18732);
and U19317 (N_19317,N_18641,N_18821);
nand U19318 (N_19318,N_18931,N_18694);
and U19319 (N_19319,N_18709,N_18973);
xnor U19320 (N_19320,N_18775,N_18641);
xor U19321 (N_19321,N_18713,N_18648);
and U19322 (N_19322,N_18768,N_18732);
xnor U19323 (N_19323,N_18724,N_18501);
nand U19324 (N_19324,N_18629,N_18678);
xor U19325 (N_19325,N_18550,N_18724);
xnor U19326 (N_19326,N_18552,N_18854);
and U19327 (N_19327,N_18873,N_18809);
or U19328 (N_19328,N_18645,N_18660);
xnor U19329 (N_19329,N_18684,N_18756);
or U19330 (N_19330,N_18595,N_18811);
or U19331 (N_19331,N_18927,N_18815);
nor U19332 (N_19332,N_18926,N_18767);
nor U19333 (N_19333,N_18916,N_18746);
and U19334 (N_19334,N_18665,N_18606);
nor U19335 (N_19335,N_18509,N_18573);
or U19336 (N_19336,N_18841,N_18672);
nand U19337 (N_19337,N_18511,N_18514);
nor U19338 (N_19338,N_18802,N_18935);
nand U19339 (N_19339,N_18625,N_18549);
nand U19340 (N_19340,N_18994,N_18760);
and U19341 (N_19341,N_18987,N_18821);
and U19342 (N_19342,N_18613,N_18821);
nor U19343 (N_19343,N_18772,N_18722);
nand U19344 (N_19344,N_18747,N_18992);
and U19345 (N_19345,N_18683,N_18527);
nand U19346 (N_19346,N_18605,N_18565);
and U19347 (N_19347,N_18780,N_18818);
xnor U19348 (N_19348,N_18503,N_18811);
or U19349 (N_19349,N_18961,N_18954);
xor U19350 (N_19350,N_18723,N_18570);
or U19351 (N_19351,N_18622,N_18718);
and U19352 (N_19352,N_18750,N_18684);
and U19353 (N_19353,N_18725,N_18884);
nand U19354 (N_19354,N_18677,N_18930);
nor U19355 (N_19355,N_18878,N_18884);
nor U19356 (N_19356,N_18594,N_18906);
xnor U19357 (N_19357,N_18589,N_18707);
nand U19358 (N_19358,N_18684,N_18817);
xor U19359 (N_19359,N_18886,N_18717);
nand U19360 (N_19360,N_18992,N_18566);
nor U19361 (N_19361,N_18592,N_18923);
nand U19362 (N_19362,N_18566,N_18962);
and U19363 (N_19363,N_18674,N_18687);
xor U19364 (N_19364,N_18674,N_18571);
nand U19365 (N_19365,N_18899,N_18832);
and U19366 (N_19366,N_18792,N_18668);
nor U19367 (N_19367,N_18804,N_18500);
nor U19368 (N_19368,N_18984,N_18790);
nand U19369 (N_19369,N_18655,N_18844);
and U19370 (N_19370,N_18616,N_18854);
nand U19371 (N_19371,N_18592,N_18746);
xnor U19372 (N_19372,N_18958,N_18720);
nand U19373 (N_19373,N_18619,N_18861);
and U19374 (N_19374,N_18529,N_18862);
nand U19375 (N_19375,N_18534,N_18575);
xor U19376 (N_19376,N_18555,N_18860);
nor U19377 (N_19377,N_18551,N_18852);
nand U19378 (N_19378,N_18536,N_18535);
nand U19379 (N_19379,N_18539,N_18897);
and U19380 (N_19380,N_18856,N_18682);
xnor U19381 (N_19381,N_18768,N_18553);
nand U19382 (N_19382,N_18707,N_18516);
or U19383 (N_19383,N_18821,N_18544);
nand U19384 (N_19384,N_18508,N_18708);
nor U19385 (N_19385,N_18804,N_18503);
xnor U19386 (N_19386,N_18630,N_18815);
xor U19387 (N_19387,N_18709,N_18763);
xnor U19388 (N_19388,N_18744,N_18896);
nand U19389 (N_19389,N_18604,N_18903);
nor U19390 (N_19390,N_18734,N_18619);
or U19391 (N_19391,N_18594,N_18562);
nand U19392 (N_19392,N_18597,N_18562);
or U19393 (N_19393,N_18800,N_18596);
nand U19394 (N_19394,N_18590,N_18652);
xor U19395 (N_19395,N_18760,N_18547);
and U19396 (N_19396,N_18792,N_18588);
nand U19397 (N_19397,N_18779,N_18719);
and U19398 (N_19398,N_18732,N_18515);
xnor U19399 (N_19399,N_18906,N_18710);
xor U19400 (N_19400,N_18891,N_18632);
nor U19401 (N_19401,N_18936,N_18783);
and U19402 (N_19402,N_18576,N_18706);
or U19403 (N_19403,N_18670,N_18801);
xnor U19404 (N_19404,N_18969,N_18704);
nor U19405 (N_19405,N_18575,N_18958);
nand U19406 (N_19406,N_18780,N_18826);
xor U19407 (N_19407,N_18729,N_18954);
xnor U19408 (N_19408,N_18931,N_18729);
nor U19409 (N_19409,N_18527,N_18663);
nor U19410 (N_19410,N_18799,N_18545);
or U19411 (N_19411,N_18907,N_18736);
xor U19412 (N_19412,N_18960,N_18559);
or U19413 (N_19413,N_18870,N_18976);
nor U19414 (N_19414,N_18934,N_18891);
nor U19415 (N_19415,N_18991,N_18737);
nor U19416 (N_19416,N_18510,N_18987);
xor U19417 (N_19417,N_18634,N_18952);
nor U19418 (N_19418,N_18880,N_18573);
or U19419 (N_19419,N_18515,N_18856);
or U19420 (N_19420,N_18585,N_18671);
nand U19421 (N_19421,N_18789,N_18882);
nor U19422 (N_19422,N_18755,N_18716);
or U19423 (N_19423,N_18738,N_18993);
and U19424 (N_19424,N_18713,N_18624);
xor U19425 (N_19425,N_18523,N_18870);
or U19426 (N_19426,N_18779,N_18797);
nor U19427 (N_19427,N_18917,N_18682);
nand U19428 (N_19428,N_18681,N_18606);
or U19429 (N_19429,N_18932,N_18614);
and U19430 (N_19430,N_18976,N_18980);
and U19431 (N_19431,N_18950,N_18945);
nor U19432 (N_19432,N_18906,N_18790);
or U19433 (N_19433,N_18794,N_18747);
and U19434 (N_19434,N_18698,N_18823);
or U19435 (N_19435,N_18628,N_18640);
and U19436 (N_19436,N_18888,N_18907);
nand U19437 (N_19437,N_18565,N_18761);
nor U19438 (N_19438,N_18587,N_18915);
and U19439 (N_19439,N_18796,N_18747);
nand U19440 (N_19440,N_18817,N_18793);
and U19441 (N_19441,N_18922,N_18781);
nor U19442 (N_19442,N_18761,N_18830);
or U19443 (N_19443,N_18945,N_18524);
and U19444 (N_19444,N_18990,N_18892);
nor U19445 (N_19445,N_18925,N_18967);
xnor U19446 (N_19446,N_18726,N_18525);
or U19447 (N_19447,N_18827,N_18943);
xnor U19448 (N_19448,N_18597,N_18590);
and U19449 (N_19449,N_18867,N_18556);
xnor U19450 (N_19450,N_18502,N_18942);
or U19451 (N_19451,N_18890,N_18614);
or U19452 (N_19452,N_18901,N_18917);
nand U19453 (N_19453,N_18549,N_18795);
nor U19454 (N_19454,N_18865,N_18969);
xor U19455 (N_19455,N_18774,N_18696);
nor U19456 (N_19456,N_18540,N_18642);
or U19457 (N_19457,N_18618,N_18697);
xnor U19458 (N_19458,N_18859,N_18865);
or U19459 (N_19459,N_18804,N_18596);
or U19460 (N_19460,N_18916,N_18808);
nand U19461 (N_19461,N_18587,N_18957);
xnor U19462 (N_19462,N_18512,N_18915);
nand U19463 (N_19463,N_18765,N_18688);
nor U19464 (N_19464,N_18936,N_18550);
and U19465 (N_19465,N_18563,N_18707);
and U19466 (N_19466,N_18951,N_18960);
or U19467 (N_19467,N_18620,N_18598);
and U19468 (N_19468,N_18882,N_18691);
and U19469 (N_19469,N_18708,N_18884);
xor U19470 (N_19470,N_18905,N_18682);
nand U19471 (N_19471,N_18851,N_18994);
xor U19472 (N_19472,N_18920,N_18894);
nand U19473 (N_19473,N_18544,N_18565);
or U19474 (N_19474,N_18910,N_18703);
xor U19475 (N_19475,N_18862,N_18584);
nor U19476 (N_19476,N_18574,N_18934);
and U19477 (N_19477,N_18607,N_18929);
or U19478 (N_19478,N_18533,N_18630);
nand U19479 (N_19479,N_18769,N_18534);
nor U19480 (N_19480,N_18836,N_18504);
nor U19481 (N_19481,N_18630,N_18963);
nor U19482 (N_19482,N_18777,N_18938);
and U19483 (N_19483,N_18923,N_18841);
nor U19484 (N_19484,N_18930,N_18766);
nand U19485 (N_19485,N_18693,N_18884);
and U19486 (N_19486,N_18577,N_18540);
nor U19487 (N_19487,N_18873,N_18564);
nor U19488 (N_19488,N_18716,N_18715);
or U19489 (N_19489,N_18830,N_18561);
or U19490 (N_19490,N_18737,N_18825);
nor U19491 (N_19491,N_18656,N_18563);
and U19492 (N_19492,N_18963,N_18751);
xnor U19493 (N_19493,N_18610,N_18602);
xnor U19494 (N_19494,N_18864,N_18901);
or U19495 (N_19495,N_18674,N_18755);
nand U19496 (N_19496,N_18687,N_18677);
nand U19497 (N_19497,N_18627,N_18974);
or U19498 (N_19498,N_18984,N_18800);
nor U19499 (N_19499,N_18680,N_18872);
nand U19500 (N_19500,N_19449,N_19447);
and U19501 (N_19501,N_19046,N_19400);
or U19502 (N_19502,N_19142,N_19191);
nand U19503 (N_19503,N_19481,N_19389);
xnor U19504 (N_19504,N_19440,N_19165);
and U19505 (N_19505,N_19458,N_19099);
nor U19506 (N_19506,N_19118,N_19081);
or U19507 (N_19507,N_19164,N_19214);
nor U19508 (N_19508,N_19235,N_19073);
nor U19509 (N_19509,N_19336,N_19473);
nand U19510 (N_19510,N_19104,N_19024);
or U19511 (N_19511,N_19415,N_19326);
xor U19512 (N_19512,N_19064,N_19213);
or U19513 (N_19513,N_19428,N_19451);
xor U19514 (N_19514,N_19391,N_19055);
or U19515 (N_19515,N_19395,N_19450);
nand U19516 (N_19516,N_19373,N_19479);
nor U19517 (N_19517,N_19338,N_19343);
or U19518 (N_19518,N_19075,N_19207);
or U19519 (N_19519,N_19319,N_19052);
xor U19520 (N_19520,N_19102,N_19009);
or U19521 (N_19521,N_19334,N_19025);
and U19522 (N_19522,N_19433,N_19443);
or U19523 (N_19523,N_19444,N_19129);
nand U19524 (N_19524,N_19196,N_19240);
nand U19525 (N_19525,N_19166,N_19227);
nand U19526 (N_19526,N_19237,N_19072);
nand U19527 (N_19527,N_19362,N_19303);
and U19528 (N_19528,N_19304,N_19393);
nand U19529 (N_19529,N_19162,N_19051);
xnor U19530 (N_19530,N_19154,N_19257);
xnor U19531 (N_19531,N_19098,N_19267);
nand U19532 (N_19532,N_19000,N_19374);
xnor U19533 (N_19533,N_19288,N_19232);
xnor U19534 (N_19534,N_19403,N_19406);
nand U19535 (N_19535,N_19396,N_19271);
xor U19536 (N_19536,N_19140,N_19039);
nor U19537 (N_19537,N_19048,N_19120);
or U19538 (N_19538,N_19454,N_19020);
nand U19539 (N_19539,N_19408,N_19351);
xnor U19540 (N_19540,N_19144,N_19347);
or U19541 (N_19541,N_19471,N_19372);
and U19542 (N_19542,N_19094,N_19381);
nand U19543 (N_19543,N_19115,N_19302);
and U19544 (N_19544,N_19382,N_19202);
nor U19545 (N_19545,N_19050,N_19241);
nor U19546 (N_19546,N_19483,N_19180);
nand U19547 (N_19547,N_19284,N_19044);
or U19548 (N_19548,N_19173,N_19058);
nand U19549 (N_19549,N_19457,N_19199);
xor U19550 (N_19550,N_19490,N_19033);
nand U19551 (N_19551,N_19226,N_19439);
nor U19552 (N_19552,N_19323,N_19184);
xnor U19553 (N_19553,N_19476,N_19434);
or U19554 (N_19554,N_19015,N_19459);
xnor U19555 (N_19555,N_19385,N_19187);
nand U19556 (N_19556,N_19455,N_19054);
nand U19557 (N_19557,N_19276,N_19268);
nor U19558 (N_19558,N_19088,N_19464);
xnor U19559 (N_19559,N_19363,N_19038);
nor U19560 (N_19560,N_19090,N_19156);
xnor U19561 (N_19561,N_19378,N_19280);
and U19562 (N_19562,N_19040,N_19059);
xor U19563 (N_19563,N_19157,N_19300);
and U19564 (N_19564,N_19273,N_19113);
and U19565 (N_19565,N_19469,N_19126);
xnor U19566 (N_19566,N_19265,N_19127);
or U19567 (N_19567,N_19390,N_19200);
nand U19568 (N_19568,N_19082,N_19225);
xor U19569 (N_19569,N_19239,N_19100);
or U19570 (N_19570,N_19007,N_19489);
or U19571 (N_19571,N_19361,N_19143);
or U19572 (N_19572,N_19315,N_19124);
and U19573 (N_19573,N_19233,N_19321);
xnor U19574 (N_19574,N_19308,N_19078);
nor U19575 (N_19575,N_19001,N_19410);
or U19576 (N_19576,N_19172,N_19117);
and U19577 (N_19577,N_19096,N_19367);
nor U19578 (N_19578,N_19085,N_19478);
or U19579 (N_19579,N_19460,N_19356);
xnor U19580 (N_19580,N_19138,N_19488);
nand U19581 (N_19581,N_19087,N_19339);
nand U19582 (N_19582,N_19270,N_19247);
nor U19583 (N_19583,N_19296,N_19204);
xnor U19584 (N_19584,N_19206,N_19008);
and U19585 (N_19585,N_19417,N_19132);
or U19586 (N_19586,N_19245,N_19371);
xnor U19587 (N_19587,N_19168,N_19375);
and U19588 (N_19588,N_19305,N_19155);
xnor U19589 (N_19589,N_19077,N_19224);
nor U19590 (N_19590,N_19452,N_19324);
and U19591 (N_19591,N_19217,N_19063);
and U19592 (N_19592,N_19397,N_19071);
or U19593 (N_19593,N_19092,N_19432);
nand U19594 (N_19594,N_19466,N_19448);
xnor U19595 (N_19595,N_19218,N_19335);
or U19596 (N_19596,N_19364,N_19125);
nand U19597 (N_19597,N_19491,N_19269);
and U19598 (N_19598,N_19274,N_19176);
nand U19599 (N_19599,N_19170,N_19262);
nor U19600 (N_19600,N_19145,N_19005);
nor U19601 (N_19601,N_19135,N_19057);
nand U19602 (N_19602,N_19353,N_19116);
nor U19603 (N_19603,N_19027,N_19492);
and U19604 (N_19604,N_19016,N_19175);
or U19605 (N_19605,N_19482,N_19146);
nor U19606 (N_19606,N_19197,N_19211);
xnor U19607 (N_19607,N_19256,N_19462);
nor U19608 (N_19608,N_19034,N_19086);
nand U19609 (N_19609,N_19183,N_19309);
or U19610 (N_19610,N_19287,N_19139);
nand U19611 (N_19611,N_19035,N_19472);
or U19612 (N_19612,N_19107,N_19272);
and U19613 (N_19613,N_19074,N_19163);
xnor U19614 (N_19614,N_19043,N_19178);
nand U19615 (N_19615,N_19453,N_19091);
nand U19616 (N_19616,N_19108,N_19003);
nand U19617 (N_19617,N_19203,N_19341);
or U19618 (N_19618,N_19133,N_19350);
nand U19619 (N_19619,N_19147,N_19498);
and U19620 (N_19620,N_19292,N_19243);
or U19621 (N_19621,N_19076,N_19251);
nor U19622 (N_19622,N_19402,N_19419);
and U19623 (N_19623,N_19194,N_19437);
nor U19624 (N_19624,N_19426,N_19463);
nand U19625 (N_19625,N_19179,N_19101);
xor U19626 (N_19626,N_19006,N_19424);
xor U19627 (N_19627,N_19030,N_19456);
nand U19628 (N_19628,N_19312,N_19185);
nand U19629 (N_19629,N_19357,N_19429);
nand U19630 (N_19630,N_19327,N_19366);
nand U19631 (N_19631,N_19413,N_19103);
or U19632 (N_19632,N_19340,N_19369);
or U19633 (N_19633,N_19320,N_19499);
and U19634 (N_19634,N_19332,N_19106);
xnor U19635 (N_19635,N_19401,N_19109);
nor U19636 (N_19636,N_19134,N_19136);
nand U19637 (N_19637,N_19249,N_19061);
or U19638 (N_19638,N_19392,N_19310);
and U19639 (N_19639,N_19119,N_19209);
xor U19640 (N_19640,N_19438,N_19407);
and U19641 (N_19641,N_19151,N_19167);
nor U19642 (N_19642,N_19285,N_19198);
nand U19643 (N_19643,N_19067,N_19021);
nor U19644 (N_19644,N_19474,N_19289);
and U19645 (N_19645,N_19279,N_19377);
and U19646 (N_19646,N_19255,N_19148);
nor U19647 (N_19647,N_19445,N_19355);
and U19648 (N_19648,N_19311,N_19299);
nand U19649 (N_19649,N_19089,N_19468);
nor U19650 (N_19650,N_19123,N_19023);
or U19651 (N_19651,N_19066,N_19246);
nand U19652 (N_19652,N_19045,N_19242);
xnor U19653 (N_19653,N_19494,N_19149);
or U19654 (N_19654,N_19193,N_19370);
nor U19655 (N_19655,N_19158,N_19354);
and U19656 (N_19656,N_19275,N_19250);
nand U19657 (N_19657,N_19398,N_19263);
nand U19658 (N_19658,N_19037,N_19253);
nand U19659 (N_19659,N_19436,N_19261);
or U19660 (N_19660,N_19153,N_19314);
or U19661 (N_19661,N_19301,N_19348);
nand U19662 (N_19662,N_19475,N_19002);
xor U19663 (N_19663,N_19084,N_19095);
nor U19664 (N_19664,N_19031,N_19306);
or U19665 (N_19665,N_19496,N_19049);
or U19666 (N_19666,N_19137,N_19152);
xor U19667 (N_19667,N_19497,N_19248);
xor U19668 (N_19668,N_19441,N_19386);
nand U19669 (N_19669,N_19110,N_19365);
or U19670 (N_19670,N_19079,N_19461);
nand U19671 (N_19671,N_19019,N_19430);
nand U19672 (N_19672,N_19368,N_19223);
and U19673 (N_19673,N_19036,N_19421);
or U19674 (N_19674,N_19388,N_19022);
and U19675 (N_19675,N_19254,N_19328);
or U19676 (N_19676,N_19412,N_19277);
or U19677 (N_19677,N_19062,N_19345);
xnor U19678 (N_19678,N_19486,N_19159);
nand U19679 (N_19679,N_19283,N_19220);
and U19680 (N_19680,N_19404,N_19219);
or U19681 (N_19681,N_19068,N_19212);
nor U19682 (N_19682,N_19346,N_19290);
xnor U19683 (N_19683,N_19480,N_19174);
nand U19684 (N_19684,N_19161,N_19231);
xnor U19685 (N_19685,N_19416,N_19411);
nor U19686 (N_19686,N_19422,N_19383);
and U19687 (N_19687,N_19012,N_19011);
and U19688 (N_19688,N_19358,N_19337);
xnor U19689 (N_19689,N_19189,N_19186);
nand U19690 (N_19690,N_19083,N_19069);
xor U19691 (N_19691,N_19181,N_19208);
and U19692 (N_19692,N_19465,N_19041);
nor U19693 (N_19693,N_19216,N_19405);
and U19694 (N_19694,N_19294,N_19318);
and U19695 (N_19695,N_19316,N_19418);
xor U19696 (N_19696,N_19435,N_19032);
or U19697 (N_19697,N_19360,N_19210);
or U19698 (N_19698,N_19177,N_19286);
and U19699 (N_19699,N_19010,N_19234);
or U19700 (N_19700,N_19493,N_19150);
nand U19701 (N_19701,N_19409,N_19260);
nand U19702 (N_19702,N_19359,N_19477);
and U19703 (N_19703,N_19013,N_19379);
and U19704 (N_19704,N_19384,N_19238);
or U19705 (N_19705,N_19278,N_19349);
nand U19706 (N_19706,N_19331,N_19188);
or U19707 (N_19707,N_19128,N_19282);
and U19708 (N_19708,N_19442,N_19112);
or U19709 (N_19709,N_19295,N_19431);
xnor U19710 (N_19710,N_19467,N_19169);
and U19711 (N_19711,N_19291,N_19171);
or U19712 (N_19712,N_19495,N_19047);
xor U19713 (N_19713,N_19229,N_19121);
or U19714 (N_19714,N_19322,N_19026);
nor U19715 (N_19715,N_19230,N_19221);
and U19716 (N_19716,N_19293,N_19065);
nand U19717 (N_19717,N_19258,N_19425);
xnor U19718 (N_19718,N_19266,N_19329);
and U19719 (N_19719,N_19080,N_19004);
xor U19720 (N_19720,N_19333,N_19122);
xor U19721 (N_19721,N_19053,N_19427);
xor U19722 (N_19722,N_19195,N_19205);
nor U19723 (N_19723,N_19192,N_19330);
nand U19724 (N_19724,N_19376,N_19160);
and U19725 (N_19725,N_19281,N_19259);
xnor U19726 (N_19726,N_19060,N_19042);
nor U19727 (N_19727,N_19017,N_19093);
or U19728 (N_19728,N_19414,N_19352);
xnor U19729 (N_19729,N_19297,N_19111);
nand U19730 (N_19730,N_19244,N_19317);
nor U19731 (N_19731,N_19313,N_19446);
or U19732 (N_19732,N_19028,N_19342);
nand U19733 (N_19733,N_19190,N_19056);
nand U19734 (N_19734,N_19097,N_19387);
and U19735 (N_19735,N_19298,N_19236);
or U19736 (N_19736,N_19070,N_19307);
or U19737 (N_19737,N_19344,N_19029);
xor U19738 (N_19738,N_19182,N_19325);
nor U19739 (N_19739,N_19487,N_19420);
or U19740 (N_19740,N_19252,N_19201);
nor U19741 (N_19741,N_19114,N_19380);
and U19742 (N_19742,N_19105,N_19485);
or U19743 (N_19743,N_19131,N_19141);
or U19744 (N_19744,N_19215,N_19470);
nor U19745 (N_19745,N_19264,N_19014);
xnor U19746 (N_19746,N_19018,N_19423);
nand U19747 (N_19747,N_19484,N_19399);
and U19748 (N_19748,N_19228,N_19394);
nand U19749 (N_19749,N_19130,N_19222);
nand U19750 (N_19750,N_19218,N_19312);
nor U19751 (N_19751,N_19280,N_19028);
xnor U19752 (N_19752,N_19132,N_19166);
nand U19753 (N_19753,N_19438,N_19280);
nor U19754 (N_19754,N_19150,N_19302);
nand U19755 (N_19755,N_19000,N_19251);
or U19756 (N_19756,N_19135,N_19062);
xnor U19757 (N_19757,N_19297,N_19136);
xnor U19758 (N_19758,N_19014,N_19105);
and U19759 (N_19759,N_19324,N_19083);
and U19760 (N_19760,N_19237,N_19171);
nor U19761 (N_19761,N_19007,N_19284);
nor U19762 (N_19762,N_19433,N_19351);
and U19763 (N_19763,N_19465,N_19025);
and U19764 (N_19764,N_19110,N_19147);
xor U19765 (N_19765,N_19275,N_19405);
or U19766 (N_19766,N_19029,N_19145);
nor U19767 (N_19767,N_19024,N_19020);
nand U19768 (N_19768,N_19272,N_19195);
xor U19769 (N_19769,N_19259,N_19378);
nand U19770 (N_19770,N_19075,N_19477);
or U19771 (N_19771,N_19167,N_19121);
or U19772 (N_19772,N_19013,N_19405);
xnor U19773 (N_19773,N_19366,N_19195);
nand U19774 (N_19774,N_19020,N_19145);
nor U19775 (N_19775,N_19338,N_19026);
or U19776 (N_19776,N_19299,N_19147);
nand U19777 (N_19777,N_19248,N_19423);
nor U19778 (N_19778,N_19428,N_19295);
xor U19779 (N_19779,N_19024,N_19298);
xnor U19780 (N_19780,N_19218,N_19316);
and U19781 (N_19781,N_19432,N_19459);
xor U19782 (N_19782,N_19470,N_19102);
nand U19783 (N_19783,N_19266,N_19200);
and U19784 (N_19784,N_19296,N_19110);
and U19785 (N_19785,N_19288,N_19220);
or U19786 (N_19786,N_19168,N_19129);
xnor U19787 (N_19787,N_19217,N_19205);
nand U19788 (N_19788,N_19497,N_19267);
nor U19789 (N_19789,N_19121,N_19299);
xor U19790 (N_19790,N_19052,N_19469);
xor U19791 (N_19791,N_19157,N_19115);
or U19792 (N_19792,N_19473,N_19090);
xnor U19793 (N_19793,N_19426,N_19314);
nor U19794 (N_19794,N_19464,N_19013);
and U19795 (N_19795,N_19308,N_19350);
and U19796 (N_19796,N_19400,N_19268);
or U19797 (N_19797,N_19111,N_19417);
and U19798 (N_19798,N_19323,N_19338);
or U19799 (N_19799,N_19152,N_19409);
or U19800 (N_19800,N_19146,N_19256);
and U19801 (N_19801,N_19353,N_19175);
or U19802 (N_19802,N_19025,N_19057);
nand U19803 (N_19803,N_19367,N_19235);
nand U19804 (N_19804,N_19313,N_19189);
and U19805 (N_19805,N_19069,N_19444);
and U19806 (N_19806,N_19460,N_19232);
or U19807 (N_19807,N_19016,N_19423);
nand U19808 (N_19808,N_19460,N_19037);
nor U19809 (N_19809,N_19376,N_19295);
nand U19810 (N_19810,N_19046,N_19094);
or U19811 (N_19811,N_19338,N_19340);
nand U19812 (N_19812,N_19293,N_19476);
and U19813 (N_19813,N_19176,N_19470);
xnor U19814 (N_19814,N_19310,N_19358);
nand U19815 (N_19815,N_19264,N_19361);
or U19816 (N_19816,N_19154,N_19206);
and U19817 (N_19817,N_19093,N_19324);
xnor U19818 (N_19818,N_19101,N_19012);
or U19819 (N_19819,N_19472,N_19153);
xor U19820 (N_19820,N_19198,N_19391);
and U19821 (N_19821,N_19101,N_19358);
nor U19822 (N_19822,N_19097,N_19060);
xnor U19823 (N_19823,N_19266,N_19410);
nor U19824 (N_19824,N_19403,N_19197);
or U19825 (N_19825,N_19033,N_19340);
nor U19826 (N_19826,N_19200,N_19335);
xnor U19827 (N_19827,N_19238,N_19084);
nand U19828 (N_19828,N_19206,N_19119);
xor U19829 (N_19829,N_19249,N_19271);
or U19830 (N_19830,N_19361,N_19281);
or U19831 (N_19831,N_19274,N_19334);
xnor U19832 (N_19832,N_19208,N_19094);
nor U19833 (N_19833,N_19368,N_19168);
xnor U19834 (N_19834,N_19086,N_19243);
or U19835 (N_19835,N_19090,N_19414);
nor U19836 (N_19836,N_19016,N_19034);
nand U19837 (N_19837,N_19318,N_19121);
or U19838 (N_19838,N_19014,N_19476);
or U19839 (N_19839,N_19258,N_19494);
and U19840 (N_19840,N_19223,N_19194);
nand U19841 (N_19841,N_19229,N_19264);
nand U19842 (N_19842,N_19443,N_19066);
nand U19843 (N_19843,N_19471,N_19468);
and U19844 (N_19844,N_19188,N_19486);
or U19845 (N_19845,N_19229,N_19332);
or U19846 (N_19846,N_19021,N_19031);
xnor U19847 (N_19847,N_19084,N_19015);
nand U19848 (N_19848,N_19048,N_19067);
xor U19849 (N_19849,N_19018,N_19468);
or U19850 (N_19850,N_19394,N_19089);
xor U19851 (N_19851,N_19477,N_19110);
xnor U19852 (N_19852,N_19060,N_19073);
nor U19853 (N_19853,N_19137,N_19403);
nor U19854 (N_19854,N_19351,N_19218);
nor U19855 (N_19855,N_19126,N_19319);
and U19856 (N_19856,N_19205,N_19238);
xnor U19857 (N_19857,N_19058,N_19405);
or U19858 (N_19858,N_19097,N_19103);
or U19859 (N_19859,N_19061,N_19311);
or U19860 (N_19860,N_19329,N_19001);
nor U19861 (N_19861,N_19422,N_19369);
nor U19862 (N_19862,N_19373,N_19328);
xor U19863 (N_19863,N_19469,N_19379);
nand U19864 (N_19864,N_19361,N_19229);
nor U19865 (N_19865,N_19034,N_19322);
nor U19866 (N_19866,N_19035,N_19160);
and U19867 (N_19867,N_19467,N_19000);
and U19868 (N_19868,N_19355,N_19439);
nor U19869 (N_19869,N_19016,N_19203);
and U19870 (N_19870,N_19130,N_19304);
nand U19871 (N_19871,N_19037,N_19144);
xnor U19872 (N_19872,N_19395,N_19081);
and U19873 (N_19873,N_19232,N_19161);
xor U19874 (N_19874,N_19333,N_19234);
and U19875 (N_19875,N_19065,N_19329);
nand U19876 (N_19876,N_19207,N_19283);
xor U19877 (N_19877,N_19262,N_19258);
or U19878 (N_19878,N_19198,N_19150);
nor U19879 (N_19879,N_19476,N_19300);
nand U19880 (N_19880,N_19380,N_19015);
nor U19881 (N_19881,N_19068,N_19194);
or U19882 (N_19882,N_19198,N_19444);
nand U19883 (N_19883,N_19286,N_19316);
and U19884 (N_19884,N_19186,N_19076);
and U19885 (N_19885,N_19042,N_19237);
nand U19886 (N_19886,N_19497,N_19119);
and U19887 (N_19887,N_19301,N_19485);
nand U19888 (N_19888,N_19223,N_19437);
nand U19889 (N_19889,N_19200,N_19230);
or U19890 (N_19890,N_19373,N_19317);
or U19891 (N_19891,N_19422,N_19438);
nor U19892 (N_19892,N_19004,N_19219);
nand U19893 (N_19893,N_19158,N_19293);
and U19894 (N_19894,N_19465,N_19108);
xor U19895 (N_19895,N_19153,N_19140);
or U19896 (N_19896,N_19418,N_19176);
nor U19897 (N_19897,N_19198,N_19074);
nand U19898 (N_19898,N_19238,N_19392);
nor U19899 (N_19899,N_19238,N_19461);
nand U19900 (N_19900,N_19353,N_19216);
nor U19901 (N_19901,N_19467,N_19342);
nand U19902 (N_19902,N_19204,N_19008);
xnor U19903 (N_19903,N_19361,N_19044);
nor U19904 (N_19904,N_19418,N_19132);
nor U19905 (N_19905,N_19027,N_19385);
nor U19906 (N_19906,N_19012,N_19286);
nand U19907 (N_19907,N_19088,N_19293);
xnor U19908 (N_19908,N_19493,N_19073);
and U19909 (N_19909,N_19311,N_19264);
nor U19910 (N_19910,N_19280,N_19302);
xnor U19911 (N_19911,N_19074,N_19343);
xor U19912 (N_19912,N_19073,N_19472);
or U19913 (N_19913,N_19193,N_19416);
nand U19914 (N_19914,N_19499,N_19134);
xor U19915 (N_19915,N_19345,N_19494);
xnor U19916 (N_19916,N_19093,N_19146);
xnor U19917 (N_19917,N_19497,N_19087);
or U19918 (N_19918,N_19245,N_19153);
nand U19919 (N_19919,N_19318,N_19498);
and U19920 (N_19920,N_19433,N_19324);
or U19921 (N_19921,N_19189,N_19276);
or U19922 (N_19922,N_19278,N_19049);
xor U19923 (N_19923,N_19077,N_19236);
nand U19924 (N_19924,N_19488,N_19311);
nand U19925 (N_19925,N_19020,N_19311);
and U19926 (N_19926,N_19337,N_19071);
nor U19927 (N_19927,N_19064,N_19413);
xnor U19928 (N_19928,N_19330,N_19124);
and U19929 (N_19929,N_19363,N_19128);
or U19930 (N_19930,N_19134,N_19127);
and U19931 (N_19931,N_19020,N_19228);
nor U19932 (N_19932,N_19215,N_19334);
xor U19933 (N_19933,N_19050,N_19464);
and U19934 (N_19934,N_19126,N_19239);
and U19935 (N_19935,N_19111,N_19084);
xor U19936 (N_19936,N_19271,N_19032);
nand U19937 (N_19937,N_19007,N_19281);
and U19938 (N_19938,N_19202,N_19135);
nand U19939 (N_19939,N_19306,N_19004);
nand U19940 (N_19940,N_19010,N_19431);
xor U19941 (N_19941,N_19181,N_19192);
nor U19942 (N_19942,N_19467,N_19383);
and U19943 (N_19943,N_19078,N_19174);
nor U19944 (N_19944,N_19145,N_19305);
nor U19945 (N_19945,N_19063,N_19344);
nor U19946 (N_19946,N_19092,N_19331);
xor U19947 (N_19947,N_19491,N_19365);
nand U19948 (N_19948,N_19334,N_19048);
and U19949 (N_19949,N_19139,N_19031);
or U19950 (N_19950,N_19061,N_19185);
and U19951 (N_19951,N_19009,N_19303);
or U19952 (N_19952,N_19076,N_19462);
nor U19953 (N_19953,N_19222,N_19407);
or U19954 (N_19954,N_19458,N_19477);
nand U19955 (N_19955,N_19492,N_19275);
or U19956 (N_19956,N_19432,N_19313);
or U19957 (N_19957,N_19400,N_19213);
or U19958 (N_19958,N_19224,N_19294);
nand U19959 (N_19959,N_19308,N_19272);
xor U19960 (N_19960,N_19363,N_19254);
xnor U19961 (N_19961,N_19234,N_19485);
nor U19962 (N_19962,N_19182,N_19464);
or U19963 (N_19963,N_19268,N_19093);
and U19964 (N_19964,N_19378,N_19456);
and U19965 (N_19965,N_19372,N_19310);
or U19966 (N_19966,N_19431,N_19003);
or U19967 (N_19967,N_19371,N_19168);
nand U19968 (N_19968,N_19256,N_19394);
nor U19969 (N_19969,N_19121,N_19070);
nor U19970 (N_19970,N_19450,N_19368);
nor U19971 (N_19971,N_19403,N_19290);
nor U19972 (N_19972,N_19358,N_19100);
xor U19973 (N_19973,N_19118,N_19225);
and U19974 (N_19974,N_19113,N_19306);
xnor U19975 (N_19975,N_19471,N_19205);
or U19976 (N_19976,N_19102,N_19390);
or U19977 (N_19977,N_19232,N_19401);
and U19978 (N_19978,N_19195,N_19088);
and U19979 (N_19979,N_19253,N_19426);
and U19980 (N_19980,N_19307,N_19310);
nor U19981 (N_19981,N_19359,N_19316);
and U19982 (N_19982,N_19415,N_19045);
xnor U19983 (N_19983,N_19227,N_19416);
xor U19984 (N_19984,N_19475,N_19089);
xor U19985 (N_19985,N_19458,N_19329);
nor U19986 (N_19986,N_19432,N_19376);
nor U19987 (N_19987,N_19158,N_19487);
nand U19988 (N_19988,N_19003,N_19341);
nor U19989 (N_19989,N_19137,N_19271);
nor U19990 (N_19990,N_19195,N_19006);
and U19991 (N_19991,N_19480,N_19103);
xnor U19992 (N_19992,N_19032,N_19081);
and U19993 (N_19993,N_19335,N_19405);
nor U19994 (N_19994,N_19201,N_19314);
nor U19995 (N_19995,N_19255,N_19164);
nor U19996 (N_19996,N_19368,N_19190);
or U19997 (N_19997,N_19008,N_19345);
nand U19998 (N_19998,N_19495,N_19457);
or U19999 (N_19999,N_19341,N_19190);
nor U20000 (N_20000,N_19851,N_19753);
or U20001 (N_20001,N_19668,N_19715);
xor U20002 (N_20002,N_19676,N_19747);
nand U20003 (N_20003,N_19734,N_19654);
or U20004 (N_20004,N_19873,N_19742);
nand U20005 (N_20005,N_19822,N_19605);
nand U20006 (N_20006,N_19616,N_19512);
nor U20007 (N_20007,N_19876,N_19545);
or U20008 (N_20008,N_19701,N_19729);
and U20009 (N_20009,N_19641,N_19696);
or U20010 (N_20010,N_19798,N_19840);
nor U20011 (N_20011,N_19749,N_19765);
xnor U20012 (N_20012,N_19553,N_19607);
nand U20013 (N_20013,N_19967,N_19856);
xor U20014 (N_20014,N_19965,N_19969);
or U20015 (N_20015,N_19580,N_19933);
and U20016 (N_20016,N_19841,N_19863);
nand U20017 (N_20017,N_19702,N_19835);
nand U20018 (N_20018,N_19651,N_19532);
or U20019 (N_20019,N_19789,N_19975);
nor U20020 (N_20020,N_19591,N_19511);
nor U20021 (N_20021,N_19501,N_19977);
or U20022 (N_20022,N_19963,N_19735);
or U20023 (N_20023,N_19821,N_19530);
nand U20024 (N_20024,N_19976,N_19684);
and U20025 (N_20025,N_19554,N_19935);
xor U20026 (N_20026,N_19859,N_19535);
xor U20027 (N_20027,N_19636,N_19884);
nand U20028 (N_20028,N_19795,N_19836);
nand U20029 (N_20029,N_19722,N_19907);
nor U20030 (N_20030,N_19630,N_19877);
xnor U20031 (N_20031,N_19693,N_19912);
or U20032 (N_20032,N_19883,N_19891);
nand U20033 (N_20033,N_19783,N_19540);
nor U20034 (N_20034,N_19612,N_19970);
xnor U20035 (N_20035,N_19908,N_19714);
or U20036 (N_20036,N_19584,N_19737);
or U20037 (N_20037,N_19522,N_19770);
nor U20038 (N_20038,N_19806,N_19611);
or U20039 (N_20039,N_19646,N_19999);
nand U20040 (N_20040,N_19872,N_19746);
nor U20041 (N_20041,N_19927,N_19763);
nor U20042 (N_20042,N_19647,N_19643);
or U20043 (N_20043,N_19586,N_19582);
nor U20044 (N_20044,N_19675,N_19953);
and U20045 (N_20045,N_19812,N_19538);
or U20046 (N_20046,N_19791,N_19960);
or U20047 (N_20047,N_19968,N_19743);
nand U20048 (N_20048,N_19906,N_19569);
or U20049 (N_20049,N_19921,N_19725);
nor U20050 (N_20050,N_19762,N_19982);
or U20051 (N_20051,N_19780,N_19561);
or U20052 (N_20052,N_19815,N_19857);
and U20053 (N_20053,N_19614,N_19817);
nor U20054 (N_20054,N_19936,N_19593);
nand U20055 (N_20055,N_19740,N_19677);
xnor U20056 (N_20056,N_19916,N_19871);
nand U20057 (N_20057,N_19931,N_19825);
and U20058 (N_20058,N_19576,N_19588);
nor U20059 (N_20059,N_19955,N_19750);
nor U20060 (N_20060,N_19978,N_19704);
xor U20061 (N_20061,N_19682,N_19502);
or U20062 (N_20062,N_19920,N_19519);
nor U20063 (N_20063,N_19830,N_19659);
nor U20064 (N_20064,N_19796,N_19577);
nor U20065 (N_20065,N_19596,N_19813);
or U20066 (N_20066,N_19855,N_19503);
and U20067 (N_20067,N_19673,N_19666);
nor U20068 (N_20068,N_19504,N_19686);
and U20069 (N_20069,N_19619,N_19680);
or U20070 (N_20070,N_19984,N_19900);
nand U20071 (N_20071,N_19555,N_19784);
or U20072 (N_20072,N_19698,N_19544);
xor U20073 (N_20073,N_19837,N_19515);
and U20074 (N_20074,N_19990,N_19957);
nor U20075 (N_20075,N_19951,N_19950);
xnor U20076 (N_20076,N_19772,N_19758);
or U20077 (N_20077,N_19664,N_19602);
xor U20078 (N_20078,N_19560,N_19550);
nand U20079 (N_20079,N_19928,N_19868);
nor U20080 (N_20080,N_19697,N_19542);
or U20081 (N_20081,N_19639,N_19741);
and U20082 (N_20082,N_19958,N_19521);
xnor U20083 (N_20083,N_19624,N_19803);
xor U20084 (N_20084,N_19991,N_19635);
xor U20085 (N_20085,N_19531,N_19961);
xor U20086 (N_20086,N_19962,N_19709);
or U20087 (N_20087,N_19681,N_19939);
nor U20088 (N_20088,N_19942,N_19730);
xnor U20089 (N_20089,N_19838,N_19988);
and U20090 (N_20090,N_19774,N_19756);
or U20091 (N_20091,N_19513,N_19843);
or U20092 (N_20092,N_19563,N_19606);
or U20093 (N_20093,N_19518,N_19979);
and U20094 (N_20094,N_19947,N_19570);
or U20095 (N_20095,N_19731,N_19685);
xor U20096 (N_20096,N_19880,N_19896);
nand U20097 (N_20097,N_19801,N_19925);
nor U20098 (N_20098,N_19674,N_19574);
and U20099 (N_20099,N_19833,N_19946);
xor U20100 (N_20100,N_19971,N_19543);
nor U20101 (N_20101,N_19745,N_19728);
nor U20102 (N_20102,N_19768,N_19887);
xnor U20103 (N_20103,N_19794,N_19679);
nor U20104 (N_20104,N_19670,N_19759);
or U20105 (N_20105,N_19541,N_19993);
nor U20106 (N_20106,N_19583,N_19648);
nand U20107 (N_20107,N_19599,N_19549);
xnor U20108 (N_20108,N_19726,N_19736);
or U20109 (N_20109,N_19621,N_19754);
xnor U20110 (N_20110,N_19779,N_19592);
xnor U20111 (N_20111,N_19536,N_19655);
xor U20112 (N_20112,N_19909,N_19886);
or U20113 (N_20113,N_19827,N_19802);
nand U20114 (N_20114,N_19618,N_19687);
or U20115 (N_20115,N_19678,N_19524);
nand U20116 (N_20116,N_19790,N_19776);
and U20117 (N_20117,N_19787,N_19769);
and U20118 (N_20118,N_19778,N_19994);
xor U20119 (N_20119,N_19601,N_19878);
or U20120 (N_20120,N_19706,N_19566);
and U20121 (N_20121,N_19672,N_19819);
nand U20122 (N_20122,N_19667,N_19954);
and U20123 (N_20123,N_19915,N_19854);
nor U20124 (N_20124,N_19792,N_19898);
nor U20125 (N_20125,N_19785,N_19914);
nor U20126 (N_20126,N_19869,N_19913);
or U20127 (N_20127,N_19797,N_19923);
and U20128 (N_20128,N_19849,N_19949);
and U20129 (N_20129,N_19810,N_19807);
and U20130 (N_20130,N_19842,N_19829);
or U20131 (N_20131,N_19665,N_19692);
and U20132 (N_20132,N_19874,N_19809);
or U20133 (N_20133,N_19505,N_19608);
nor U20134 (N_20134,N_19587,N_19864);
nor U20135 (N_20135,N_19889,N_19782);
or U20136 (N_20136,N_19805,N_19831);
nand U20137 (N_20137,N_19890,N_19567);
xor U20138 (N_20138,N_19788,N_19980);
or U20139 (N_20139,N_19562,N_19860);
and U20140 (N_20140,N_19721,N_19930);
and U20141 (N_20141,N_19650,N_19617);
xnor U20142 (N_20142,N_19767,N_19610);
or U20143 (N_20143,N_19552,N_19534);
nor U20144 (N_20144,N_19852,N_19671);
and U20145 (N_20145,N_19633,N_19564);
nor U20146 (N_20146,N_19568,N_19903);
xor U20147 (N_20147,N_19811,N_19661);
nand U20148 (N_20148,N_19517,N_19653);
xnor U20149 (N_20149,N_19516,N_19508);
or U20150 (N_20150,N_19964,N_19800);
nor U20151 (N_20151,N_19997,N_19594);
nand U20152 (N_20152,N_19645,N_19700);
xor U20153 (N_20153,N_19724,N_19952);
or U20154 (N_20154,N_19509,N_19711);
xnor U20155 (N_20155,N_19656,N_19764);
nor U20156 (N_20156,N_19657,N_19848);
nand U20157 (N_20157,N_19893,N_19823);
and U20158 (N_20158,N_19732,N_19966);
and U20159 (N_20159,N_19885,N_19558);
nor U20160 (N_20160,N_19603,N_19691);
xor U20161 (N_20161,N_19705,N_19649);
and U20162 (N_20162,N_19985,N_19717);
nor U20163 (N_20163,N_19695,N_19941);
nor U20164 (N_20164,N_19755,N_19590);
or U20165 (N_20165,N_19853,N_19622);
and U20166 (N_20166,N_19981,N_19926);
xnor U20167 (N_20167,N_19634,N_19986);
or U20168 (N_20168,N_19720,N_19771);
xnor U20169 (N_20169,N_19631,N_19609);
nor U20170 (N_20170,N_19895,N_19845);
or U20171 (N_20171,N_19760,N_19520);
xnor U20172 (N_20172,N_19944,N_19808);
nand U20173 (N_20173,N_19751,N_19500);
nor U20174 (N_20174,N_19904,N_19738);
nor U20175 (N_20175,N_19644,N_19559);
and U20176 (N_20176,N_19992,N_19620);
nand U20177 (N_20177,N_19866,N_19551);
nor U20178 (N_20178,N_19793,N_19959);
xor U20179 (N_20179,N_19556,N_19716);
nand U20180 (N_20180,N_19847,N_19713);
xnor U20181 (N_20181,N_19727,N_19652);
nand U20182 (N_20182,N_19781,N_19637);
xnor U20183 (N_20183,N_19526,N_19761);
and U20184 (N_20184,N_19589,N_19604);
or U20185 (N_20185,N_19699,N_19989);
nor U20186 (N_20186,N_19919,N_19998);
and U20187 (N_20187,N_19861,N_19956);
xor U20188 (N_20188,N_19694,N_19839);
xor U20189 (N_20189,N_19703,N_19879);
xnor U20190 (N_20190,N_19565,N_19688);
and U20191 (N_20191,N_19826,N_19973);
nor U20192 (N_20192,N_19718,N_19902);
or U20193 (N_20193,N_19940,N_19707);
and U20194 (N_20194,N_19897,N_19548);
or U20195 (N_20195,N_19929,N_19932);
or U20196 (N_20196,N_19660,N_19816);
or U20197 (N_20197,N_19917,N_19875);
xnor U20198 (N_20198,N_19892,N_19938);
nand U20199 (N_20199,N_19514,N_19527);
nand U20200 (N_20200,N_19537,N_19804);
nand U20201 (N_20201,N_19744,N_19640);
or U20202 (N_20202,N_19628,N_19623);
and U20203 (N_20203,N_19748,N_19882);
or U20204 (N_20204,N_19905,N_19525);
and U20205 (N_20205,N_19934,N_19547);
and U20206 (N_20206,N_19777,N_19996);
nor U20207 (N_20207,N_19862,N_19571);
nand U20208 (N_20208,N_19662,N_19578);
xor U20209 (N_20209,N_19625,N_19824);
or U20210 (N_20210,N_19597,N_19775);
or U20211 (N_20211,N_19899,N_19773);
or U20212 (N_20212,N_19894,N_19865);
nand U20213 (N_20213,N_19658,N_19757);
or U20214 (N_20214,N_19799,N_19948);
or U20215 (N_20215,N_19850,N_19881);
nor U20216 (N_20216,N_19867,N_19638);
nand U20217 (N_20217,N_19888,N_19708);
nand U20218 (N_20218,N_19585,N_19710);
or U20219 (N_20219,N_19663,N_19572);
nand U20220 (N_20220,N_19595,N_19814);
nor U20221 (N_20221,N_19910,N_19507);
or U20222 (N_20222,N_19669,N_19974);
xor U20223 (N_20223,N_19712,N_19828);
nor U20224 (N_20224,N_19786,N_19846);
xnor U20225 (N_20225,N_19858,N_19924);
nor U20226 (N_20226,N_19598,N_19573);
xnor U20227 (N_20227,N_19937,N_19943);
nand U20228 (N_20228,N_19870,N_19983);
and U20229 (N_20229,N_19752,N_19689);
nand U20230 (N_20230,N_19766,N_19834);
xor U20231 (N_20231,N_19546,N_19510);
nor U20232 (N_20232,N_19627,N_19818);
xor U20233 (N_20233,N_19901,N_19911);
xor U20234 (N_20234,N_19820,N_19690);
nand U20235 (N_20235,N_19972,N_19613);
xor U20236 (N_20236,N_19575,N_19615);
and U20237 (N_20237,N_19945,N_19506);
nand U20238 (N_20238,N_19719,N_19918);
and U20239 (N_20239,N_19995,N_19581);
or U20240 (N_20240,N_19600,N_19528);
and U20241 (N_20241,N_19557,N_19642);
xnor U20242 (N_20242,N_19579,N_19844);
or U20243 (N_20243,N_19922,N_19723);
and U20244 (N_20244,N_19683,N_19533);
nor U20245 (N_20245,N_19733,N_19539);
or U20246 (N_20246,N_19626,N_19632);
and U20247 (N_20247,N_19739,N_19629);
nand U20248 (N_20248,N_19529,N_19832);
xor U20249 (N_20249,N_19987,N_19523);
or U20250 (N_20250,N_19962,N_19787);
xor U20251 (N_20251,N_19645,N_19511);
xor U20252 (N_20252,N_19628,N_19894);
nor U20253 (N_20253,N_19937,N_19645);
nor U20254 (N_20254,N_19855,N_19793);
nor U20255 (N_20255,N_19565,N_19529);
nand U20256 (N_20256,N_19645,N_19834);
and U20257 (N_20257,N_19704,N_19671);
nand U20258 (N_20258,N_19751,N_19773);
nor U20259 (N_20259,N_19522,N_19525);
or U20260 (N_20260,N_19641,N_19785);
or U20261 (N_20261,N_19539,N_19605);
nand U20262 (N_20262,N_19708,N_19743);
and U20263 (N_20263,N_19534,N_19787);
nand U20264 (N_20264,N_19586,N_19584);
nor U20265 (N_20265,N_19798,N_19672);
and U20266 (N_20266,N_19843,N_19547);
xor U20267 (N_20267,N_19796,N_19914);
and U20268 (N_20268,N_19602,N_19571);
and U20269 (N_20269,N_19974,N_19706);
nand U20270 (N_20270,N_19649,N_19753);
nor U20271 (N_20271,N_19888,N_19525);
and U20272 (N_20272,N_19525,N_19699);
nand U20273 (N_20273,N_19879,N_19888);
xnor U20274 (N_20274,N_19744,N_19657);
or U20275 (N_20275,N_19929,N_19857);
or U20276 (N_20276,N_19645,N_19681);
nand U20277 (N_20277,N_19880,N_19762);
nor U20278 (N_20278,N_19528,N_19931);
nor U20279 (N_20279,N_19747,N_19576);
xor U20280 (N_20280,N_19737,N_19901);
xor U20281 (N_20281,N_19519,N_19570);
xnor U20282 (N_20282,N_19923,N_19912);
xor U20283 (N_20283,N_19906,N_19726);
or U20284 (N_20284,N_19795,N_19722);
and U20285 (N_20285,N_19591,N_19940);
or U20286 (N_20286,N_19507,N_19918);
and U20287 (N_20287,N_19588,N_19543);
and U20288 (N_20288,N_19589,N_19776);
nor U20289 (N_20289,N_19815,N_19597);
xor U20290 (N_20290,N_19680,N_19815);
or U20291 (N_20291,N_19670,N_19651);
nand U20292 (N_20292,N_19840,N_19622);
and U20293 (N_20293,N_19849,N_19979);
xnor U20294 (N_20294,N_19522,N_19933);
xor U20295 (N_20295,N_19771,N_19967);
or U20296 (N_20296,N_19627,N_19864);
nor U20297 (N_20297,N_19657,N_19691);
and U20298 (N_20298,N_19819,N_19839);
nor U20299 (N_20299,N_19917,N_19763);
nand U20300 (N_20300,N_19733,N_19797);
nor U20301 (N_20301,N_19841,N_19538);
nor U20302 (N_20302,N_19816,N_19872);
xnor U20303 (N_20303,N_19871,N_19854);
nand U20304 (N_20304,N_19870,N_19634);
or U20305 (N_20305,N_19547,N_19561);
nor U20306 (N_20306,N_19975,N_19829);
nor U20307 (N_20307,N_19965,N_19696);
nand U20308 (N_20308,N_19801,N_19862);
nand U20309 (N_20309,N_19583,N_19755);
and U20310 (N_20310,N_19554,N_19548);
and U20311 (N_20311,N_19911,N_19597);
nand U20312 (N_20312,N_19596,N_19670);
xor U20313 (N_20313,N_19887,N_19689);
or U20314 (N_20314,N_19597,N_19620);
xnor U20315 (N_20315,N_19554,N_19543);
nor U20316 (N_20316,N_19636,N_19585);
and U20317 (N_20317,N_19912,N_19529);
nor U20318 (N_20318,N_19736,N_19544);
nor U20319 (N_20319,N_19545,N_19518);
nor U20320 (N_20320,N_19616,N_19663);
or U20321 (N_20321,N_19852,N_19704);
and U20322 (N_20322,N_19655,N_19696);
or U20323 (N_20323,N_19940,N_19535);
xor U20324 (N_20324,N_19851,N_19856);
nand U20325 (N_20325,N_19957,N_19883);
or U20326 (N_20326,N_19761,N_19669);
xor U20327 (N_20327,N_19922,N_19801);
nor U20328 (N_20328,N_19879,N_19772);
nand U20329 (N_20329,N_19638,N_19799);
or U20330 (N_20330,N_19771,N_19965);
nor U20331 (N_20331,N_19811,N_19537);
xor U20332 (N_20332,N_19547,N_19993);
or U20333 (N_20333,N_19894,N_19839);
nor U20334 (N_20334,N_19802,N_19974);
and U20335 (N_20335,N_19907,N_19924);
and U20336 (N_20336,N_19877,N_19782);
nand U20337 (N_20337,N_19732,N_19528);
or U20338 (N_20338,N_19573,N_19883);
xor U20339 (N_20339,N_19991,N_19753);
or U20340 (N_20340,N_19846,N_19882);
and U20341 (N_20341,N_19614,N_19782);
xnor U20342 (N_20342,N_19718,N_19712);
xor U20343 (N_20343,N_19669,N_19580);
nand U20344 (N_20344,N_19798,N_19567);
and U20345 (N_20345,N_19650,N_19603);
or U20346 (N_20346,N_19613,N_19839);
nor U20347 (N_20347,N_19598,N_19729);
nand U20348 (N_20348,N_19983,N_19831);
xnor U20349 (N_20349,N_19514,N_19517);
nand U20350 (N_20350,N_19961,N_19536);
or U20351 (N_20351,N_19901,N_19806);
xnor U20352 (N_20352,N_19801,N_19687);
nor U20353 (N_20353,N_19889,N_19858);
nor U20354 (N_20354,N_19847,N_19718);
or U20355 (N_20355,N_19624,N_19875);
or U20356 (N_20356,N_19689,N_19778);
xnor U20357 (N_20357,N_19554,N_19961);
nand U20358 (N_20358,N_19704,N_19849);
and U20359 (N_20359,N_19680,N_19647);
nor U20360 (N_20360,N_19555,N_19795);
and U20361 (N_20361,N_19748,N_19778);
xor U20362 (N_20362,N_19838,N_19741);
nand U20363 (N_20363,N_19883,N_19524);
nand U20364 (N_20364,N_19660,N_19843);
or U20365 (N_20365,N_19830,N_19684);
nor U20366 (N_20366,N_19834,N_19563);
nand U20367 (N_20367,N_19838,N_19800);
or U20368 (N_20368,N_19531,N_19863);
nand U20369 (N_20369,N_19896,N_19943);
xor U20370 (N_20370,N_19673,N_19880);
nand U20371 (N_20371,N_19862,N_19793);
nand U20372 (N_20372,N_19871,N_19576);
and U20373 (N_20373,N_19872,N_19725);
xnor U20374 (N_20374,N_19538,N_19965);
nand U20375 (N_20375,N_19809,N_19763);
nand U20376 (N_20376,N_19618,N_19952);
nand U20377 (N_20377,N_19905,N_19983);
nand U20378 (N_20378,N_19848,N_19527);
and U20379 (N_20379,N_19504,N_19997);
nor U20380 (N_20380,N_19824,N_19669);
nand U20381 (N_20381,N_19551,N_19845);
nor U20382 (N_20382,N_19758,N_19704);
nand U20383 (N_20383,N_19605,N_19527);
nand U20384 (N_20384,N_19941,N_19582);
xnor U20385 (N_20385,N_19898,N_19540);
nand U20386 (N_20386,N_19612,N_19813);
xnor U20387 (N_20387,N_19931,N_19926);
nor U20388 (N_20388,N_19792,N_19983);
or U20389 (N_20389,N_19553,N_19672);
or U20390 (N_20390,N_19842,N_19832);
nor U20391 (N_20391,N_19635,N_19536);
xnor U20392 (N_20392,N_19517,N_19564);
xnor U20393 (N_20393,N_19812,N_19931);
nor U20394 (N_20394,N_19708,N_19751);
xnor U20395 (N_20395,N_19889,N_19506);
nand U20396 (N_20396,N_19673,N_19986);
and U20397 (N_20397,N_19828,N_19913);
nor U20398 (N_20398,N_19974,N_19573);
xnor U20399 (N_20399,N_19690,N_19655);
nor U20400 (N_20400,N_19828,N_19623);
or U20401 (N_20401,N_19870,N_19990);
and U20402 (N_20402,N_19901,N_19525);
or U20403 (N_20403,N_19796,N_19862);
and U20404 (N_20404,N_19673,N_19524);
and U20405 (N_20405,N_19817,N_19784);
nor U20406 (N_20406,N_19506,N_19618);
nand U20407 (N_20407,N_19575,N_19803);
xor U20408 (N_20408,N_19837,N_19775);
nor U20409 (N_20409,N_19839,N_19544);
and U20410 (N_20410,N_19517,N_19842);
xor U20411 (N_20411,N_19588,N_19887);
xor U20412 (N_20412,N_19837,N_19840);
xnor U20413 (N_20413,N_19673,N_19916);
nand U20414 (N_20414,N_19981,N_19894);
nand U20415 (N_20415,N_19512,N_19975);
or U20416 (N_20416,N_19911,N_19817);
and U20417 (N_20417,N_19863,N_19623);
or U20418 (N_20418,N_19707,N_19866);
and U20419 (N_20419,N_19674,N_19931);
xnor U20420 (N_20420,N_19528,N_19970);
nor U20421 (N_20421,N_19884,N_19861);
nand U20422 (N_20422,N_19659,N_19677);
nand U20423 (N_20423,N_19726,N_19900);
nand U20424 (N_20424,N_19721,N_19949);
nor U20425 (N_20425,N_19686,N_19710);
or U20426 (N_20426,N_19535,N_19730);
and U20427 (N_20427,N_19910,N_19871);
and U20428 (N_20428,N_19586,N_19583);
xnor U20429 (N_20429,N_19919,N_19615);
xor U20430 (N_20430,N_19537,N_19821);
and U20431 (N_20431,N_19665,N_19703);
or U20432 (N_20432,N_19628,N_19640);
nand U20433 (N_20433,N_19645,N_19670);
nor U20434 (N_20434,N_19620,N_19976);
nand U20435 (N_20435,N_19913,N_19502);
nor U20436 (N_20436,N_19926,N_19755);
nor U20437 (N_20437,N_19970,N_19960);
nor U20438 (N_20438,N_19576,N_19729);
and U20439 (N_20439,N_19578,N_19911);
xnor U20440 (N_20440,N_19996,N_19712);
xnor U20441 (N_20441,N_19792,N_19515);
or U20442 (N_20442,N_19724,N_19518);
nor U20443 (N_20443,N_19570,N_19505);
nand U20444 (N_20444,N_19868,N_19857);
or U20445 (N_20445,N_19694,N_19669);
and U20446 (N_20446,N_19882,N_19667);
and U20447 (N_20447,N_19596,N_19647);
or U20448 (N_20448,N_19874,N_19903);
nand U20449 (N_20449,N_19650,N_19705);
and U20450 (N_20450,N_19576,N_19632);
or U20451 (N_20451,N_19563,N_19755);
nand U20452 (N_20452,N_19556,N_19824);
nor U20453 (N_20453,N_19943,N_19521);
xnor U20454 (N_20454,N_19866,N_19531);
nor U20455 (N_20455,N_19715,N_19685);
or U20456 (N_20456,N_19540,N_19664);
nand U20457 (N_20457,N_19597,N_19829);
xor U20458 (N_20458,N_19882,N_19926);
and U20459 (N_20459,N_19603,N_19633);
xor U20460 (N_20460,N_19814,N_19960);
and U20461 (N_20461,N_19706,N_19748);
or U20462 (N_20462,N_19570,N_19611);
and U20463 (N_20463,N_19530,N_19670);
nor U20464 (N_20464,N_19806,N_19931);
or U20465 (N_20465,N_19735,N_19848);
and U20466 (N_20466,N_19799,N_19968);
nand U20467 (N_20467,N_19751,N_19576);
nand U20468 (N_20468,N_19972,N_19763);
nand U20469 (N_20469,N_19781,N_19511);
or U20470 (N_20470,N_19777,N_19969);
xnor U20471 (N_20471,N_19624,N_19536);
or U20472 (N_20472,N_19965,N_19526);
nor U20473 (N_20473,N_19654,N_19603);
nand U20474 (N_20474,N_19823,N_19830);
xnor U20475 (N_20475,N_19808,N_19868);
or U20476 (N_20476,N_19752,N_19703);
nand U20477 (N_20477,N_19543,N_19937);
and U20478 (N_20478,N_19891,N_19631);
xnor U20479 (N_20479,N_19634,N_19559);
xnor U20480 (N_20480,N_19574,N_19906);
nand U20481 (N_20481,N_19878,N_19896);
nand U20482 (N_20482,N_19519,N_19975);
and U20483 (N_20483,N_19662,N_19843);
nand U20484 (N_20484,N_19731,N_19805);
xnor U20485 (N_20485,N_19913,N_19949);
and U20486 (N_20486,N_19896,N_19578);
nand U20487 (N_20487,N_19899,N_19649);
or U20488 (N_20488,N_19929,N_19673);
xnor U20489 (N_20489,N_19682,N_19579);
nand U20490 (N_20490,N_19714,N_19644);
xor U20491 (N_20491,N_19568,N_19716);
xnor U20492 (N_20492,N_19860,N_19786);
nor U20493 (N_20493,N_19624,N_19920);
nor U20494 (N_20494,N_19595,N_19881);
nor U20495 (N_20495,N_19756,N_19870);
nor U20496 (N_20496,N_19584,N_19938);
and U20497 (N_20497,N_19723,N_19954);
and U20498 (N_20498,N_19900,N_19915);
and U20499 (N_20499,N_19975,N_19768);
nand U20500 (N_20500,N_20034,N_20179);
nand U20501 (N_20501,N_20459,N_20381);
and U20502 (N_20502,N_20343,N_20045);
nor U20503 (N_20503,N_20051,N_20256);
nand U20504 (N_20504,N_20139,N_20199);
nand U20505 (N_20505,N_20353,N_20077);
and U20506 (N_20506,N_20328,N_20317);
and U20507 (N_20507,N_20074,N_20475);
xnor U20508 (N_20508,N_20333,N_20265);
nor U20509 (N_20509,N_20141,N_20050);
nand U20510 (N_20510,N_20183,N_20364);
and U20511 (N_20511,N_20425,N_20274);
nand U20512 (N_20512,N_20231,N_20053);
or U20513 (N_20513,N_20230,N_20347);
nand U20514 (N_20514,N_20498,N_20040);
nor U20515 (N_20515,N_20126,N_20217);
nor U20516 (N_20516,N_20196,N_20262);
nor U20517 (N_20517,N_20167,N_20398);
nand U20518 (N_20518,N_20487,N_20411);
or U20519 (N_20519,N_20214,N_20122);
nor U20520 (N_20520,N_20041,N_20131);
nand U20521 (N_20521,N_20293,N_20497);
or U20522 (N_20522,N_20361,N_20470);
xor U20523 (N_20523,N_20363,N_20029);
nand U20524 (N_20524,N_20039,N_20158);
and U20525 (N_20525,N_20268,N_20491);
nor U20526 (N_20526,N_20107,N_20289);
nor U20527 (N_20527,N_20061,N_20002);
xor U20528 (N_20528,N_20253,N_20073);
nor U20529 (N_20529,N_20148,N_20430);
nor U20530 (N_20530,N_20338,N_20447);
xnor U20531 (N_20531,N_20474,N_20031);
xor U20532 (N_20532,N_20127,N_20089);
xnor U20533 (N_20533,N_20365,N_20070);
xnor U20534 (N_20534,N_20480,N_20489);
and U20535 (N_20535,N_20278,N_20204);
or U20536 (N_20536,N_20134,N_20008);
and U20537 (N_20537,N_20477,N_20086);
nor U20538 (N_20538,N_20358,N_20027);
nand U20539 (N_20539,N_20090,N_20151);
and U20540 (N_20540,N_20266,N_20111);
nor U20541 (N_20541,N_20083,N_20337);
xnor U20542 (N_20542,N_20412,N_20479);
xor U20543 (N_20543,N_20420,N_20377);
or U20544 (N_20544,N_20012,N_20119);
or U20545 (N_20545,N_20250,N_20311);
or U20546 (N_20546,N_20322,N_20401);
and U20547 (N_20547,N_20427,N_20024);
or U20548 (N_20548,N_20387,N_20155);
nor U20549 (N_20549,N_20004,N_20057);
nand U20550 (N_20550,N_20055,N_20368);
nor U20551 (N_20551,N_20300,N_20354);
xnor U20552 (N_20552,N_20193,N_20048);
or U20553 (N_20553,N_20345,N_20146);
and U20554 (N_20554,N_20340,N_20424);
or U20555 (N_20555,N_20465,N_20306);
xor U20556 (N_20556,N_20021,N_20038);
or U20557 (N_20557,N_20128,N_20110);
and U20558 (N_20558,N_20207,N_20215);
nor U20559 (N_20559,N_20383,N_20476);
xnor U20560 (N_20560,N_20150,N_20097);
nor U20561 (N_20561,N_20101,N_20032);
nor U20562 (N_20562,N_20376,N_20466);
xor U20563 (N_20563,N_20344,N_20005);
nor U20564 (N_20564,N_20117,N_20094);
or U20565 (N_20565,N_20314,N_20174);
or U20566 (N_20566,N_20209,N_20299);
and U20567 (N_20567,N_20147,N_20185);
xnor U20568 (N_20568,N_20145,N_20351);
and U20569 (N_20569,N_20442,N_20091);
and U20570 (N_20570,N_20049,N_20301);
and U20571 (N_20571,N_20013,N_20330);
nand U20572 (N_20572,N_20218,N_20190);
nand U20573 (N_20573,N_20009,N_20244);
xor U20574 (N_20574,N_20198,N_20348);
or U20575 (N_20575,N_20432,N_20393);
or U20576 (N_20576,N_20332,N_20279);
nor U20577 (N_20577,N_20187,N_20241);
nand U20578 (N_20578,N_20087,N_20372);
xnor U20579 (N_20579,N_20177,N_20473);
nand U20580 (N_20580,N_20052,N_20288);
and U20581 (N_20581,N_20054,N_20451);
nand U20582 (N_20582,N_20403,N_20114);
nor U20583 (N_20583,N_20191,N_20220);
nor U20584 (N_20584,N_20437,N_20325);
or U20585 (N_20585,N_20120,N_20416);
nor U20586 (N_20586,N_20211,N_20036);
or U20587 (N_20587,N_20342,N_20017);
nand U20588 (N_20588,N_20302,N_20494);
or U20589 (N_20589,N_20271,N_20224);
nor U20590 (N_20590,N_20227,N_20273);
or U20591 (N_20591,N_20312,N_20249);
nand U20592 (N_20592,N_20104,N_20406);
xor U20593 (N_20593,N_20238,N_20349);
nor U20594 (N_20594,N_20113,N_20388);
nand U20595 (N_20595,N_20135,N_20153);
nand U20596 (N_20596,N_20162,N_20176);
nand U20597 (N_20597,N_20023,N_20413);
xnor U20598 (N_20598,N_20285,N_20492);
nand U20599 (N_20599,N_20258,N_20367);
xnor U20600 (N_20600,N_20402,N_20064);
nor U20601 (N_20601,N_20251,N_20163);
nand U20602 (N_20602,N_20431,N_20272);
and U20603 (N_20603,N_20389,N_20189);
or U20604 (N_20604,N_20356,N_20275);
and U20605 (N_20605,N_20105,N_20390);
xor U20606 (N_20606,N_20281,N_20294);
or U20607 (N_20607,N_20173,N_20448);
or U20608 (N_20608,N_20205,N_20267);
and U20609 (N_20609,N_20071,N_20248);
and U20610 (N_20610,N_20240,N_20316);
nand U20611 (N_20611,N_20092,N_20096);
and U20612 (N_20612,N_20161,N_20234);
nor U20613 (N_20613,N_20103,N_20252);
xnor U20614 (N_20614,N_20108,N_20461);
nand U20615 (N_20615,N_20458,N_20144);
nor U20616 (N_20616,N_20010,N_20011);
nand U20617 (N_20617,N_20493,N_20047);
or U20618 (N_20618,N_20125,N_20006);
or U20619 (N_20619,N_20043,N_20331);
nand U20620 (N_20620,N_20060,N_20391);
or U20621 (N_20621,N_20371,N_20197);
xnor U20622 (N_20622,N_20374,N_20438);
nor U20623 (N_20623,N_20478,N_20419);
and U20624 (N_20624,N_20310,N_20025);
and U20625 (N_20625,N_20042,N_20429);
nor U20626 (N_20626,N_20219,N_20082);
xor U20627 (N_20627,N_20378,N_20007);
or U20628 (N_20628,N_20015,N_20168);
and U20629 (N_20629,N_20315,N_20308);
xnor U20630 (N_20630,N_20022,N_20320);
and U20631 (N_20631,N_20433,N_20026);
or U20632 (N_20632,N_20186,N_20072);
or U20633 (N_20633,N_20000,N_20418);
xor U20634 (N_20634,N_20235,N_20467);
or U20635 (N_20635,N_20323,N_20321);
nand U20636 (N_20636,N_20399,N_20346);
and U20637 (N_20637,N_20123,N_20414);
and U20638 (N_20638,N_20297,N_20078);
xor U20639 (N_20639,N_20386,N_20203);
xor U20640 (N_20640,N_20166,N_20341);
nor U20641 (N_20641,N_20172,N_20257);
and U20642 (N_20642,N_20138,N_20201);
or U20643 (N_20643,N_20407,N_20225);
nand U20644 (N_20644,N_20446,N_20370);
or U20645 (N_20645,N_20069,N_20450);
and U20646 (N_20646,N_20067,N_20366);
xor U20647 (N_20647,N_20495,N_20408);
nand U20648 (N_20648,N_20109,N_20260);
or U20649 (N_20649,N_20362,N_20254);
xnor U20650 (N_20650,N_20415,N_20129);
nor U20651 (N_20651,N_20212,N_20384);
xor U20652 (N_20652,N_20350,N_20202);
and U20653 (N_20653,N_20453,N_20093);
xnor U20654 (N_20654,N_20084,N_20284);
nor U20655 (N_20655,N_20304,N_20352);
nand U20656 (N_20656,N_20460,N_20280);
nor U20657 (N_20657,N_20436,N_20132);
or U20658 (N_20658,N_20178,N_20065);
nand U20659 (N_20659,N_20454,N_20395);
nor U20660 (N_20660,N_20417,N_20276);
and U20661 (N_20661,N_20357,N_20062);
nor U20662 (N_20662,N_20160,N_20359);
nand U20663 (N_20663,N_20355,N_20206);
nor U20664 (N_20664,N_20392,N_20223);
or U20665 (N_20665,N_20428,N_20449);
nand U20666 (N_20666,N_20472,N_20044);
or U20667 (N_20667,N_20484,N_20059);
xnor U20668 (N_20668,N_20194,N_20295);
nor U20669 (N_20669,N_20259,N_20490);
nor U20670 (N_20670,N_20441,N_20255);
nor U20671 (N_20671,N_20226,N_20222);
nor U20672 (N_20672,N_20499,N_20075);
nand U20673 (N_20673,N_20099,N_20016);
xnor U20674 (N_20674,N_20133,N_20270);
nor U20675 (N_20675,N_20319,N_20379);
xor U20676 (N_20676,N_20014,N_20313);
and U20677 (N_20677,N_20124,N_20339);
nor U20678 (N_20678,N_20137,N_20360);
xnor U20679 (N_20679,N_20030,N_20434);
nand U20680 (N_20680,N_20243,N_20159);
nor U20681 (N_20681,N_20462,N_20307);
or U20682 (N_20682,N_20143,N_20112);
xor U20683 (N_20683,N_20095,N_20182);
or U20684 (N_20684,N_20118,N_20396);
and U20685 (N_20685,N_20181,N_20033);
nand U20686 (N_20686,N_20154,N_20422);
nor U20687 (N_20687,N_20200,N_20169);
and U20688 (N_20688,N_20385,N_20210);
or U20689 (N_20689,N_20213,N_20242);
or U20690 (N_20690,N_20003,N_20239);
and U20691 (N_20691,N_20157,N_20152);
xnor U20692 (N_20692,N_20076,N_20247);
nand U20693 (N_20693,N_20171,N_20245);
nand U20694 (N_20694,N_20236,N_20056);
nor U20695 (N_20695,N_20496,N_20326);
xor U20696 (N_20696,N_20232,N_20318);
or U20697 (N_20697,N_20290,N_20400);
and U20698 (N_20698,N_20063,N_20115);
nand U20699 (N_20699,N_20404,N_20456);
nor U20700 (N_20700,N_20263,N_20375);
and U20701 (N_20701,N_20394,N_20121);
or U20702 (N_20702,N_20019,N_20440);
or U20703 (N_20703,N_20149,N_20409);
nand U20704 (N_20704,N_20028,N_20046);
xor U20705 (N_20705,N_20098,N_20068);
xor U20706 (N_20706,N_20471,N_20081);
xnor U20707 (N_20707,N_20164,N_20269);
or U20708 (N_20708,N_20291,N_20102);
or U20709 (N_20709,N_20106,N_20373);
nand U20710 (N_20710,N_20445,N_20100);
or U20711 (N_20711,N_20327,N_20463);
and U20712 (N_20712,N_20485,N_20296);
or U20713 (N_20713,N_20180,N_20208);
nand U20714 (N_20714,N_20221,N_20324);
or U20715 (N_20715,N_20080,N_20283);
xor U20716 (N_20716,N_20469,N_20001);
nand U20717 (N_20717,N_20405,N_20426);
nor U20718 (N_20718,N_20292,N_20035);
or U20719 (N_20719,N_20468,N_20136);
xor U20720 (N_20720,N_20079,N_20303);
or U20721 (N_20721,N_20443,N_20421);
xnor U20722 (N_20722,N_20192,N_20184);
nor U20723 (N_20723,N_20195,N_20261);
or U20724 (N_20724,N_20140,N_20282);
nor U20725 (N_20725,N_20329,N_20058);
xor U20726 (N_20726,N_20481,N_20287);
and U20727 (N_20727,N_20170,N_20088);
nand U20728 (N_20728,N_20457,N_20237);
nor U20729 (N_20729,N_20188,N_20486);
or U20730 (N_20730,N_20423,N_20455);
nor U20731 (N_20731,N_20264,N_20435);
and U20732 (N_20732,N_20334,N_20216);
nor U20733 (N_20733,N_20085,N_20175);
nand U20734 (N_20734,N_20246,N_20397);
or U20735 (N_20735,N_20298,N_20439);
or U20736 (N_20736,N_20483,N_20309);
nor U20737 (N_20737,N_20165,N_20380);
nand U20738 (N_20738,N_20382,N_20020);
nand U20739 (N_20739,N_20305,N_20277);
nor U20740 (N_20740,N_20488,N_20018);
or U20741 (N_20741,N_20335,N_20369);
xnor U20742 (N_20742,N_20156,N_20037);
nor U20743 (N_20743,N_20116,N_20233);
xnor U20744 (N_20744,N_20444,N_20410);
nand U20745 (N_20745,N_20336,N_20229);
xnor U20746 (N_20746,N_20286,N_20142);
or U20747 (N_20747,N_20066,N_20482);
or U20748 (N_20748,N_20228,N_20464);
nand U20749 (N_20749,N_20130,N_20452);
nand U20750 (N_20750,N_20056,N_20374);
or U20751 (N_20751,N_20484,N_20166);
nor U20752 (N_20752,N_20107,N_20167);
nor U20753 (N_20753,N_20303,N_20155);
or U20754 (N_20754,N_20350,N_20472);
nor U20755 (N_20755,N_20199,N_20315);
and U20756 (N_20756,N_20465,N_20008);
or U20757 (N_20757,N_20057,N_20110);
nand U20758 (N_20758,N_20332,N_20077);
nand U20759 (N_20759,N_20359,N_20398);
and U20760 (N_20760,N_20434,N_20072);
or U20761 (N_20761,N_20188,N_20107);
and U20762 (N_20762,N_20337,N_20301);
and U20763 (N_20763,N_20199,N_20330);
or U20764 (N_20764,N_20234,N_20148);
nand U20765 (N_20765,N_20432,N_20489);
or U20766 (N_20766,N_20338,N_20339);
nor U20767 (N_20767,N_20405,N_20427);
nor U20768 (N_20768,N_20107,N_20403);
and U20769 (N_20769,N_20344,N_20072);
nor U20770 (N_20770,N_20348,N_20060);
or U20771 (N_20771,N_20044,N_20247);
xor U20772 (N_20772,N_20420,N_20036);
nor U20773 (N_20773,N_20256,N_20084);
xor U20774 (N_20774,N_20273,N_20155);
nor U20775 (N_20775,N_20219,N_20098);
and U20776 (N_20776,N_20464,N_20003);
xnor U20777 (N_20777,N_20494,N_20175);
xor U20778 (N_20778,N_20284,N_20016);
or U20779 (N_20779,N_20214,N_20330);
xor U20780 (N_20780,N_20139,N_20361);
xnor U20781 (N_20781,N_20426,N_20222);
xor U20782 (N_20782,N_20294,N_20237);
and U20783 (N_20783,N_20378,N_20393);
nand U20784 (N_20784,N_20369,N_20135);
xnor U20785 (N_20785,N_20288,N_20421);
xor U20786 (N_20786,N_20229,N_20465);
xor U20787 (N_20787,N_20140,N_20055);
nand U20788 (N_20788,N_20121,N_20481);
nand U20789 (N_20789,N_20244,N_20488);
nand U20790 (N_20790,N_20020,N_20349);
or U20791 (N_20791,N_20088,N_20460);
xor U20792 (N_20792,N_20133,N_20442);
xor U20793 (N_20793,N_20191,N_20100);
nand U20794 (N_20794,N_20136,N_20372);
nor U20795 (N_20795,N_20105,N_20385);
nand U20796 (N_20796,N_20233,N_20171);
nor U20797 (N_20797,N_20212,N_20343);
and U20798 (N_20798,N_20480,N_20115);
nor U20799 (N_20799,N_20283,N_20350);
and U20800 (N_20800,N_20183,N_20166);
nand U20801 (N_20801,N_20243,N_20470);
xor U20802 (N_20802,N_20001,N_20496);
or U20803 (N_20803,N_20138,N_20162);
nor U20804 (N_20804,N_20379,N_20417);
and U20805 (N_20805,N_20473,N_20454);
xor U20806 (N_20806,N_20203,N_20340);
xnor U20807 (N_20807,N_20132,N_20330);
and U20808 (N_20808,N_20195,N_20433);
xor U20809 (N_20809,N_20157,N_20452);
xor U20810 (N_20810,N_20406,N_20155);
nor U20811 (N_20811,N_20063,N_20307);
or U20812 (N_20812,N_20160,N_20117);
nand U20813 (N_20813,N_20238,N_20211);
and U20814 (N_20814,N_20414,N_20292);
and U20815 (N_20815,N_20481,N_20236);
nand U20816 (N_20816,N_20213,N_20150);
or U20817 (N_20817,N_20191,N_20162);
xnor U20818 (N_20818,N_20186,N_20476);
xor U20819 (N_20819,N_20035,N_20466);
nand U20820 (N_20820,N_20189,N_20352);
nand U20821 (N_20821,N_20374,N_20280);
or U20822 (N_20822,N_20337,N_20465);
nor U20823 (N_20823,N_20066,N_20355);
xor U20824 (N_20824,N_20304,N_20075);
nor U20825 (N_20825,N_20492,N_20026);
or U20826 (N_20826,N_20489,N_20479);
nor U20827 (N_20827,N_20212,N_20027);
xor U20828 (N_20828,N_20391,N_20489);
nand U20829 (N_20829,N_20382,N_20467);
or U20830 (N_20830,N_20416,N_20223);
xor U20831 (N_20831,N_20267,N_20419);
and U20832 (N_20832,N_20461,N_20228);
nand U20833 (N_20833,N_20091,N_20377);
and U20834 (N_20834,N_20197,N_20134);
nand U20835 (N_20835,N_20292,N_20314);
and U20836 (N_20836,N_20274,N_20144);
nor U20837 (N_20837,N_20310,N_20190);
and U20838 (N_20838,N_20291,N_20138);
nand U20839 (N_20839,N_20130,N_20394);
xnor U20840 (N_20840,N_20227,N_20148);
xor U20841 (N_20841,N_20107,N_20295);
or U20842 (N_20842,N_20326,N_20251);
nand U20843 (N_20843,N_20469,N_20173);
nor U20844 (N_20844,N_20089,N_20330);
or U20845 (N_20845,N_20300,N_20396);
nor U20846 (N_20846,N_20465,N_20024);
or U20847 (N_20847,N_20257,N_20057);
and U20848 (N_20848,N_20187,N_20136);
and U20849 (N_20849,N_20042,N_20378);
xnor U20850 (N_20850,N_20184,N_20262);
or U20851 (N_20851,N_20278,N_20458);
or U20852 (N_20852,N_20073,N_20267);
nand U20853 (N_20853,N_20072,N_20307);
nand U20854 (N_20854,N_20466,N_20225);
or U20855 (N_20855,N_20074,N_20478);
xnor U20856 (N_20856,N_20069,N_20355);
and U20857 (N_20857,N_20051,N_20280);
and U20858 (N_20858,N_20325,N_20400);
nand U20859 (N_20859,N_20297,N_20103);
xor U20860 (N_20860,N_20444,N_20175);
xor U20861 (N_20861,N_20297,N_20351);
or U20862 (N_20862,N_20114,N_20351);
nand U20863 (N_20863,N_20373,N_20475);
xor U20864 (N_20864,N_20275,N_20113);
xnor U20865 (N_20865,N_20396,N_20122);
nand U20866 (N_20866,N_20247,N_20228);
xor U20867 (N_20867,N_20096,N_20491);
xnor U20868 (N_20868,N_20003,N_20107);
nor U20869 (N_20869,N_20286,N_20366);
nand U20870 (N_20870,N_20023,N_20051);
nor U20871 (N_20871,N_20041,N_20397);
xor U20872 (N_20872,N_20012,N_20141);
and U20873 (N_20873,N_20446,N_20204);
nand U20874 (N_20874,N_20455,N_20448);
or U20875 (N_20875,N_20371,N_20041);
and U20876 (N_20876,N_20496,N_20373);
nand U20877 (N_20877,N_20177,N_20443);
or U20878 (N_20878,N_20125,N_20344);
or U20879 (N_20879,N_20325,N_20303);
nand U20880 (N_20880,N_20295,N_20398);
or U20881 (N_20881,N_20050,N_20486);
nand U20882 (N_20882,N_20208,N_20004);
xnor U20883 (N_20883,N_20307,N_20278);
or U20884 (N_20884,N_20404,N_20088);
xnor U20885 (N_20885,N_20241,N_20139);
or U20886 (N_20886,N_20014,N_20180);
nand U20887 (N_20887,N_20133,N_20410);
nor U20888 (N_20888,N_20281,N_20081);
nand U20889 (N_20889,N_20027,N_20274);
and U20890 (N_20890,N_20347,N_20248);
nor U20891 (N_20891,N_20081,N_20111);
or U20892 (N_20892,N_20228,N_20026);
or U20893 (N_20893,N_20090,N_20447);
and U20894 (N_20894,N_20426,N_20259);
or U20895 (N_20895,N_20469,N_20109);
nor U20896 (N_20896,N_20321,N_20334);
xor U20897 (N_20897,N_20170,N_20176);
nand U20898 (N_20898,N_20489,N_20429);
xnor U20899 (N_20899,N_20039,N_20130);
or U20900 (N_20900,N_20066,N_20233);
and U20901 (N_20901,N_20133,N_20021);
nand U20902 (N_20902,N_20135,N_20191);
and U20903 (N_20903,N_20482,N_20048);
nand U20904 (N_20904,N_20241,N_20026);
nor U20905 (N_20905,N_20094,N_20258);
and U20906 (N_20906,N_20216,N_20168);
nor U20907 (N_20907,N_20273,N_20219);
xor U20908 (N_20908,N_20053,N_20398);
and U20909 (N_20909,N_20449,N_20054);
xnor U20910 (N_20910,N_20060,N_20434);
or U20911 (N_20911,N_20033,N_20225);
and U20912 (N_20912,N_20078,N_20466);
and U20913 (N_20913,N_20225,N_20075);
or U20914 (N_20914,N_20491,N_20222);
nand U20915 (N_20915,N_20047,N_20495);
nand U20916 (N_20916,N_20088,N_20112);
nand U20917 (N_20917,N_20411,N_20205);
and U20918 (N_20918,N_20274,N_20036);
nand U20919 (N_20919,N_20449,N_20375);
xor U20920 (N_20920,N_20255,N_20451);
xnor U20921 (N_20921,N_20328,N_20209);
nand U20922 (N_20922,N_20269,N_20155);
and U20923 (N_20923,N_20012,N_20423);
and U20924 (N_20924,N_20052,N_20108);
xor U20925 (N_20925,N_20342,N_20339);
nand U20926 (N_20926,N_20102,N_20194);
nor U20927 (N_20927,N_20260,N_20193);
or U20928 (N_20928,N_20306,N_20010);
nor U20929 (N_20929,N_20099,N_20244);
or U20930 (N_20930,N_20171,N_20253);
nor U20931 (N_20931,N_20223,N_20202);
nand U20932 (N_20932,N_20019,N_20439);
and U20933 (N_20933,N_20334,N_20159);
or U20934 (N_20934,N_20146,N_20059);
nor U20935 (N_20935,N_20495,N_20071);
nand U20936 (N_20936,N_20145,N_20209);
or U20937 (N_20937,N_20219,N_20358);
or U20938 (N_20938,N_20070,N_20130);
and U20939 (N_20939,N_20414,N_20234);
or U20940 (N_20940,N_20472,N_20262);
xnor U20941 (N_20941,N_20121,N_20137);
nor U20942 (N_20942,N_20095,N_20423);
nor U20943 (N_20943,N_20047,N_20334);
nand U20944 (N_20944,N_20163,N_20356);
xor U20945 (N_20945,N_20368,N_20198);
nor U20946 (N_20946,N_20213,N_20088);
xnor U20947 (N_20947,N_20163,N_20101);
nand U20948 (N_20948,N_20487,N_20179);
nor U20949 (N_20949,N_20022,N_20312);
xnor U20950 (N_20950,N_20018,N_20416);
nor U20951 (N_20951,N_20177,N_20235);
nand U20952 (N_20952,N_20088,N_20278);
nand U20953 (N_20953,N_20482,N_20136);
nor U20954 (N_20954,N_20382,N_20017);
and U20955 (N_20955,N_20222,N_20051);
and U20956 (N_20956,N_20361,N_20173);
xor U20957 (N_20957,N_20374,N_20128);
xnor U20958 (N_20958,N_20111,N_20148);
and U20959 (N_20959,N_20224,N_20471);
and U20960 (N_20960,N_20440,N_20164);
xnor U20961 (N_20961,N_20457,N_20452);
nand U20962 (N_20962,N_20323,N_20479);
nor U20963 (N_20963,N_20260,N_20212);
or U20964 (N_20964,N_20313,N_20479);
xnor U20965 (N_20965,N_20018,N_20477);
nand U20966 (N_20966,N_20048,N_20204);
nand U20967 (N_20967,N_20272,N_20498);
nor U20968 (N_20968,N_20075,N_20324);
and U20969 (N_20969,N_20361,N_20231);
xor U20970 (N_20970,N_20289,N_20378);
nor U20971 (N_20971,N_20394,N_20277);
nor U20972 (N_20972,N_20199,N_20468);
xnor U20973 (N_20973,N_20127,N_20244);
nand U20974 (N_20974,N_20216,N_20045);
or U20975 (N_20975,N_20125,N_20156);
nor U20976 (N_20976,N_20201,N_20158);
xor U20977 (N_20977,N_20359,N_20075);
or U20978 (N_20978,N_20369,N_20181);
xor U20979 (N_20979,N_20478,N_20488);
xnor U20980 (N_20980,N_20028,N_20074);
xor U20981 (N_20981,N_20421,N_20019);
and U20982 (N_20982,N_20220,N_20442);
nand U20983 (N_20983,N_20332,N_20459);
nand U20984 (N_20984,N_20109,N_20040);
or U20985 (N_20985,N_20237,N_20478);
nor U20986 (N_20986,N_20217,N_20428);
nor U20987 (N_20987,N_20492,N_20336);
or U20988 (N_20988,N_20109,N_20271);
nor U20989 (N_20989,N_20194,N_20320);
nand U20990 (N_20990,N_20053,N_20275);
and U20991 (N_20991,N_20360,N_20188);
and U20992 (N_20992,N_20185,N_20364);
and U20993 (N_20993,N_20215,N_20046);
xnor U20994 (N_20994,N_20293,N_20136);
xor U20995 (N_20995,N_20103,N_20099);
or U20996 (N_20996,N_20393,N_20128);
nor U20997 (N_20997,N_20377,N_20119);
nor U20998 (N_20998,N_20190,N_20161);
nand U20999 (N_20999,N_20412,N_20457);
nand U21000 (N_21000,N_20508,N_20635);
nand U21001 (N_21001,N_20564,N_20990);
xor U21002 (N_21002,N_20578,N_20815);
nor U21003 (N_21003,N_20548,N_20796);
or U21004 (N_21004,N_20643,N_20772);
or U21005 (N_21005,N_20863,N_20916);
xnor U21006 (N_21006,N_20761,N_20962);
xnor U21007 (N_21007,N_20785,N_20788);
xor U21008 (N_21008,N_20541,N_20514);
xnor U21009 (N_21009,N_20717,N_20610);
or U21010 (N_21010,N_20851,N_20773);
xor U21011 (N_21011,N_20666,N_20620);
or U21012 (N_21012,N_20664,N_20611);
xnor U21013 (N_21013,N_20752,N_20901);
xnor U21014 (N_21014,N_20707,N_20952);
xnor U21015 (N_21015,N_20905,N_20708);
nor U21016 (N_21016,N_20517,N_20600);
nand U21017 (N_21017,N_20812,N_20934);
xor U21018 (N_21018,N_20813,N_20532);
nand U21019 (N_21019,N_20994,N_20747);
nor U21020 (N_21020,N_20599,N_20999);
or U21021 (N_21021,N_20669,N_20650);
nand U21022 (N_21022,N_20911,N_20545);
or U21023 (N_21023,N_20582,N_20547);
nand U21024 (N_21024,N_20799,N_20728);
nor U21025 (N_21025,N_20959,N_20891);
xnor U21026 (N_21026,N_20646,N_20917);
xor U21027 (N_21027,N_20769,N_20876);
or U21028 (N_21028,N_20802,N_20766);
nor U21029 (N_21029,N_20682,N_20974);
and U21030 (N_21030,N_20725,N_20720);
or U21031 (N_21031,N_20843,N_20846);
nor U21032 (N_21032,N_20819,N_20888);
or U21033 (N_21033,N_20626,N_20976);
xnor U21034 (N_21034,N_20731,N_20544);
or U21035 (N_21035,N_20762,N_20982);
nor U21036 (N_21036,N_20783,N_20518);
or U21037 (N_21037,N_20632,N_20521);
or U21038 (N_21038,N_20886,N_20755);
xor U21039 (N_21039,N_20794,N_20693);
nand U21040 (N_21040,N_20734,N_20535);
nand U21041 (N_21041,N_20906,N_20557);
or U21042 (N_21042,N_20560,N_20726);
and U21043 (N_21043,N_20536,N_20505);
nor U21044 (N_21044,N_20581,N_20506);
nor U21045 (N_21045,N_20638,N_20998);
xor U21046 (N_21046,N_20692,N_20672);
or U21047 (N_21047,N_20604,N_20838);
nand U21048 (N_21048,N_20854,N_20507);
or U21049 (N_21049,N_20588,N_20567);
xor U21050 (N_21050,N_20782,N_20951);
or U21051 (N_21051,N_20943,N_20698);
and U21052 (N_21052,N_20679,N_20647);
nor U21053 (N_21053,N_20885,N_20964);
xor U21054 (N_21054,N_20842,N_20922);
nand U21055 (N_21055,N_20841,N_20711);
nand U21056 (N_21056,N_20691,N_20558);
or U21057 (N_21057,N_20655,N_20686);
nor U21058 (N_21058,N_20713,N_20520);
xnor U21059 (N_21059,N_20733,N_20798);
xor U21060 (N_21060,N_20939,N_20572);
xnor U21061 (N_21061,N_20821,N_20844);
nand U21062 (N_21062,N_20570,N_20942);
xor U21063 (N_21063,N_20897,N_20631);
or U21064 (N_21064,N_20742,N_20674);
nand U21065 (N_21065,N_20770,N_20628);
nor U21066 (N_21066,N_20884,N_20937);
and U21067 (N_21067,N_20516,N_20856);
or U21068 (N_21068,N_20966,N_20676);
xnor U21069 (N_21069,N_20525,N_20853);
nand U21070 (N_21070,N_20907,N_20503);
or U21071 (N_21071,N_20940,N_20639);
nand U21072 (N_21072,N_20661,N_20818);
nand U21073 (N_21073,N_20850,N_20721);
nand U21074 (N_21074,N_20530,N_20957);
nor U21075 (N_21075,N_20991,N_20613);
or U21076 (N_21076,N_20997,N_20584);
xor U21077 (N_21077,N_20849,N_20790);
nor U21078 (N_21078,N_20804,N_20831);
nor U21079 (N_21079,N_20967,N_20662);
and U21080 (N_21080,N_20660,N_20774);
xor U21081 (N_21081,N_20836,N_20590);
nor U21082 (N_21082,N_20882,N_20552);
nor U21083 (N_21083,N_20828,N_20542);
xor U21084 (N_21084,N_20781,N_20630);
or U21085 (N_21085,N_20933,N_20984);
and U21086 (N_21086,N_20980,N_20824);
nand U21087 (N_21087,N_20685,N_20642);
and U21088 (N_21088,N_20670,N_20866);
xor U21089 (N_21089,N_20816,N_20887);
nand U21090 (N_21090,N_20603,N_20701);
and U21091 (N_21091,N_20502,N_20736);
nand U21092 (N_21092,N_20681,N_20894);
nor U21093 (N_21093,N_20528,N_20986);
or U21094 (N_21094,N_20741,N_20823);
nand U21095 (N_21095,N_20871,N_20577);
or U21096 (N_21096,N_20948,N_20680);
nor U21097 (N_21097,N_20743,N_20554);
nand U21098 (N_21098,N_20673,N_20924);
nand U21099 (N_21099,N_20878,N_20738);
xnor U21100 (N_21100,N_20716,N_20935);
and U21101 (N_21101,N_20931,N_20960);
and U21102 (N_21102,N_20754,N_20775);
nor U21103 (N_21103,N_20864,N_20874);
or U21104 (N_21104,N_20988,N_20549);
or U21105 (N_21105,N_20969,N_20807);
nand U21106 (N_21106,N_20744,N_20973);
or U21107 (N_21107,N_20709,N_20597);
and U21108 (N_21108,N_20877,N_20817);
xnor U21109 (N_21109,N_20710,N_20677);
xor U21110 (N_21110,N_20537,N_20511);
and U21111 (N_21111,N_20657,N_20873);
nand U21112 (N_21112,N_20546,N_20792);
and U21113 (N_21113,N_20751,N_20524);
or U21114 (N_21114,N_20822,N_20668);
and U21115 (N_21115,N_20615,N_20579);
or U21116 (N_21116,N_20658,N_20621);
or U21117 (N_21117,N_20909,N_20757);
or U21118 (N_21118,N_20875,N_20765);
or U21119 (N_21119,N_20983,N_20714);
or U21120 (N_21120,N_20618,N_20789);
xor U21121 (N_21121,N_20637,N_20634);
or U21122 (N_21122,N_20921,N_20832);
and U21123 (N_21123,N_20543,N_20705);
xor U21124 (N_21124,N_20636,N_20833);
xnor U21125 (N_21125,N_20580,N_20791);
or U21126 (N_21126,N_20746,N_20972);
nand U21127 (N_21127,N_20501,N_20719);
nor U21128 (N_21128,N_20663,N_20566);
and U21129 (N_21129,N_20616,N_20756);
or U21130 (N_21130,N_20947,N_20992);
nor U21131 (N_21131,N_20779,N_20704);
and U21132 (N_21132,N_20859,N_20510);
xor U21133 (N_21133,N_20562,N_20732);
or U21134 (N_21134,N_20830,N_20624);
nor U21135 (N_21135,N_20767,N_20981);
or U21136 (N_21136,N_20556,N_20608);
xnor U21137 (N_21137,N_20869,N_20644);
nor U21138 (N_21138,N_20920,N_20550);
nand U21139 (N_21139,N_20827,N_20574);
nor U21140 (N_21140,N_20847,N_20649);
or U21141 (N_21141,N_20919,N_20946);
nand U21142 (N_21142,N_20868,N_20763);
nor U21143 (N_21143,N_20699,N_20504);
nand U21144 (N_21144,N_20723,N_20955);
nor U21145 (N_21145,N_20923,N_20979);
nor U21146 (N_21146,N_20977,N_20712);
nor U21147 (N_21147,N_20784,N_20927);
and U21148 (N_21148,N_20764,N_20961);
and U21149 (N_21149,N_20617,N_20696);
and U21150 (N_21150,N_20848,N_20722);
and U21151 (N_21151,N_20531,N_20879);
nor U21152 (N_21152,N_20750,N_20534);
or U21153 (N_21153,N_20809,N_20619);
nor U21154 (N_21154,N_20892,N_20857);
or U21155 (N_21155,N_20527,N_20801);
nor U21156 (N_21156,N_20653,N_20622);
or U21157 (N_21157,N_20926,N_20697);
xor U21158 (N_21158,N_20786,N_20695);
and U21159 (N_21159,N_20936,N_20768);
nor U21160 (N_21160,N_20865,N_20623);
and U21161 (N_21161,N_20739,N_20978);
and U21162 (N_21162,N_20573,N_20576);
and U21163 (N_21163,N_20589,N_20987);
or U21164 (N_21164,N_20860,N_20509);
nand U21165 (N_21165,N_20749,N_20513);
nand U21166 (N_21166,N_20512,N_20820);
and U21167 (N_21167,N_20727,N_20759);
or U21168 (N_21168,N_20687,N_20526);
xor U21169 (N_21169,N_20835,N_20729);
nor U21170 (N_21170,N_20963,N_20596);
and U21171 (N_21171,N_20845,N_20592);
nand U21172 (N_21172,N_20678,N_20654);
nand U21173 (N_21173,N_20591,N_20932);
and U21174 (N_21174,N_20667,N_20814);
and U21175 (N_21175,N_20870,N_20553);
xnor U21176 (N_21176,N_20910,N_20715);
and U21177 (N_21177,N_20702,N_20938);
xor U21178 (N_21178,N_20671,N_20797);
nor U21179 (N_21179,N_20918,N_20971);
nand U21180 (N_21180,N_20777,N_20595);
and U21181 (N_21181,N_20970,N_20694);
or U21182 (N_21182,N_20928,N_20855);
xor U21183 (N_21183,N_20995,N_20586);
nor U21184 (N_21184,N_20640,N_20500);
or U21185 (N_21185,N_20583,N_20771);
or U21186 (N_21186,N_20780,N_20800);
and U21187 (N_21187,N_20825,N_20861);
xor U21188 (N_21188,N_20568,N_20703);
and U21189 (N_21189,N_20985,N_20605);
xnor U21190 (N_21190,N_20645,N_20883);
xnor U21191 (N_21191,N_20522,N_20601);
nor U21192 (N_21192,N_20941,N_20593);
or U21193 (N_21193,N_20609,N_20880);
nand U21194 (N_21194,N_20895,N_20810);
and U21195 (N_21195,N_20718,N_20958);
xor U21196 (N_21196,N_20858,N_20993);
nand U21197 (N_21197,N_20837,N_20648);
nor U21198 (N_21198,N_20925,N_20614);
xnor U21199 (N_21199,N_20569,N_20559);
or U21200 (N_21200,N_20758,N_20902);
xor U21201 (N_21201,N_20659,N_20519);
nand U21202 (N_21202,N_20538,N_20598);
and U21203 (N_21203,N_20949,N_20683);
nor U21204 (N_21204,N_20730,N_20629);
xnor U21205 (N_21205,N_20806,N_20551);
xor U21206 (N_21206,N_20760,N_20915);
and U21207 (N_21207,N_20795,N_20914);
or U21208 (N_21208,N_20834,N_20690);
and U21209 (N_21209,N_20808,N_20585);
or U21210 (N_21210,N_20867,N_20896);
nor U21211 (N_21211,N_20803,N_20555);
nand U21212 (N_21212,N_20571,N_20811);
or U21213 (N_21213,N_20594,N_20627);
nor U21214 (N_21214,N_20529,N_20633);
nor U21215 (N_21215,N_20606,N_20956);
xor U21216 (N_21216,N_20904,N_20953);
and U21217 (N_21217,N_20929,N_20872);
or U21218 (N_21218,N_20665,N_20700);
xor U21219 (N_21219,N_20740,N_20996);
nor U21220 (N_21220,N_20539,N_20523);
nand U21221 (N_21221,N_20903,N_20745);
and U21222 (N_21222,N_20533,N_20913);
or U21223 (N_21223,N_20689,N_20735);
nand U21224 (N_21224,N_20563,N_20651);
and U21225 (N_21225,N_20625,N_20968);
nor U21226 (N_21226,N_20893,N_20840);
nand U21227 (N_21227,N_20944,N_20565);
xnor U21228 (N_21228,N_20688,N_20805);
nor U21229 (N_21229,N_20965,N_20826);
nor U21230 (N_21230,N_20975,N_20898);
nand U21231 (N_21231,N_20908,N_20641);
and U21232 (N_21232,N_20656,N_20652);
and U21233 (N_21233,N_20787,N_20540);
or U21234 (N_21234,N_20793,N_20612);
or U21235 (N_21235,N_20684,N_20889);
and U21236 (N_21236,N_20899,N_20737);
nand U21237 (N_21237,N_20950,N_20561);
and U21238 (N_21238,N_20575,N_20839);
and U21239 (N_21239,N_20724,N_20912);
nor U21240 (N_21240,N_20881,N_20954);
nor U21241 (N_21241,N_20602,N_20945);
nor U21242 (N_21242,N_20706,N_20862);
and U21243 (N_21243,N_20829,N_20753);
or U21244 (N_21244,N_20778,N_20748);
or U21245 (N_21245,N_20776,N_20515);
nor U21246 (N_21246,N_20852,N_20607);
xor U21247 (N_21247,N_20989,N_20900);
xnor U21248 (N_21248,N_20890,N_20930);
xor U21249 (N_21249,N_20587,N_20675);
nand U21250 (N_21250,N_20836,N_20608);
or U21251 (N_21251,N_20891,N_20681);
and U21252 (N_21252,N_20692,N_20795);
nand U21253 (N_21253,N_20888,N_20530);
and U21254 (N_21254,N_20746,N_20783);
nand U21255 (N_21255,N_20967,N_20996);
nor U21256 (N_21256,N_20763,N_20929);
xor U21257 (N_21257,N_20513,N_20527);
or U21258 (N_21258,N_20500,N_20778);
or U21259 (N_21259,N_20917,N_20753);
nand U21260 (N_21260,N_20849,N_20672);
or U21261 (N_21261,N_20691,N_20660);
or U21262 (N_21262,N_20815,N_20770);
nor U21263 (N_21263,N_20775,N_20731);
xor U21264 (N_21264,N_20826,N_20586);
or U21265 (N_21265,N_20718,N_20740);
or U21266 (N_21266,N_20656,N_20569);
and U21267 (N_21267,N_20842,N_20557);
or U21268 (N_21268,N_20525,N_20980);
xnor U21269 (N_21269,N_20851,N_20517);
nor U21270 (N_21270,N_20773,N_20770);
xnor U21271 (N_21271,N_20545,N_20977);
or U21272 (N_21272,N_20904,N_20623);
xor U21273 (N_21273,N_20661,N_20836);
nand U21274 (N_21274,N_20896,N_20711);
xnor U21275 (N_21275,N_20700,N_20835);
or U21276 (N_21276,N_20678,N_20524);
xnor U21277 (N_21277,N_20654,N_20698);
nor U21278 (N_21278,N_20862,N_20694);
or U21279 (N_21279,N_20760,N_20688);
nand U21280 (N_21280,N_20546,N_20970);
and U21281 (N_21281,N_20796,N_20857);
and U21282 (N_21282,N_20948,N_20775);
nand U21283 (N_21283,N_20618,N_20723);
or U21284 (N_21284,N_20551,N_20774);
nand U21285 (N_21285,N_20787,N_20524);
nand U21286 (N_21286,N_20532,N_20512);
nor U21287 (N_21287,N_20762,N_20879);
nor U21288 (N_21288,N_20507,N_20872);
nand U21289 (N_21289,N_20544,N_20604);
nand U21290 (N_21290,N_20592,N_20602);
nor U21291 (N_21291,N_20892,N_20920);
or U21292 (N_21292,N_20960,N_20656);
and U21293 (N_21293,N_20573,N_20524);
nor U21294 (N_21294,N_20670,N_20755);
nor U21295 (N_21295,N_20992,N_20753);
and U21296 (N_21296,N_20629,N_20754);
nor U21297 (N_21297,N_20828,N_20870);
nand U21298 (N_21298,N_20646,N_20968);
nand U21299 (N_21299,N_20746,N_20579);
or U21300 (N_21300,N_20629,N_20510);
nor U21301 (N_21301,N_20903,N_20726);
nor U21302 (N_21302,N_20866,N_20591);
and U21303 (N_21303,N_20544,N_20641);
or U21304 (N_21304,N_20922,N_20594);
nand U21305 (N_21305,N_20577,N_20933);
or U21306 (N_21306,N_20646,N_20598);
nand U21307 (N_21307,N_20536,N_20836);
nand U21308 (N_21308,N_20652,N_20541);
nand U21309 (N_21309,N_20705,N_20874);
nand U21310 (N_21310,N_20650,N_20823);
and U21311 (N_21311,N_20645,N_20977);
nand U21312 (N_21312,N_20508,N_20793);
or U21313 (N_21313,N_20596,N_20519);
and U21314 (N_21314,N_20909,N_20594);
nor U21315 (N_21315,N_20997,N_20760);
nor U21316 (N_21316,N_20566,N_20813);
and U21317 (N_21317,N_20734,N_20610);
xnor U21318 (N_21318,N_20721,N_20863);
xnor U21319 (N_21319,N_20935,N_20962);
and U21320 (N_21320,N_20740,N_20648);
and U21321 (N_21321,N_20724,N_20513);
and U21322 (N_21322,N_20971,N_20549);
and U21323 (N_21323,N_20611,N_20693);
nand U21324 (N_21324,N_20658,N_20997);
and U21325 (N_21325,N_20939,N_20874);
nor U21326 (N_21326,N_20897,N_20671);
or U21327 (N_21327,N_20846,N_20891);
or U21328 (N_21328,N_20992,N_20541);
or U21329 (N_21329,N_20849,N_20510);
xor U21330 (N_21330,N_20797,N_20789);
xnor U21331 (N_21331,N_20611,N_20981);
nand U21332 (N_21332,N_20770,N_20715);
or U21333 (N_21333,N_20892,N_20769);
nor U21334 (N_21334,N_20638,N_20547);
nor U21335 (N_21335,N_20790,N_20925);
and U21336 (N_21336,N_20550,N_20738);
xor U21337 (N_21337,N_20854,N_20819);
nand U21338 (N_21338,N_20696,N_20534);
or U21339 (N_21339,N_20591,N_20822);
nand U21340 (N_21340,N_20515,N_20549);
nor U21341 (N_21341,N_20693,N_20979);
xnor U21342 (N_21342,N_20509,N_20781);
or U21343 (N_21343,N_20954,N_20806);
nand U21344 (N_21344,N_20806,N_20622);
nand U21345 (N_21345,N_20769,N_20578);
nor U21346 (N_21346,N_20550,N_20993);
nor U21347 (N_21347,N_20814,N_20521);
nand U21348 (N_21348,N_20523,N_20997);
nand U21349 (N_21349,N_20789,N_20857);
or U21350 (N_21350,N_20997,N_20894);
nand U21351 (N_21351,N_20579,N_20988);
nor U21352 (N_21352,N_20791,N_20677);
or U21353 (N_21353,N_20765,N_20822);
and U21354 (N_21354,N_20719,N_20520);
nand U21355 (N_21355,N_20771,N_20741);
nand U21356 (N_21356,N_20886,N_20787);
nand U21357 (N_21357,N_20869,N_20745);
and U21358 (N_21358,N_20645,N_20713);
nor U21359 (N_21359,N_20620,N_20538);
and U21360 (N_21360,N_20768,N_20591);
xor U21361 (N_21361,N_20957,N_20585);
or U21362 (N_21362,N_20882,N_20802);
xnor U21363 (N_21363,N_20546,N_20597);
and U21364 (N_21364,N_20714,N_20786);
nand U21365 (N_21365,N_20903,N_20597);
nand U21366 (N_21366,N_20570,N_20664);
and U21367 (N_21367,N_20894,N_20754);
and U21368 (N_21368,N_20979,N_20654);
xnor U21369 (N_21369,N_20851,N_20730);
and U21370 (N_21370,N_20890,N_20831);
nor U21371 (N_21371,N_20678,N_20964);
xnor U21372 (N_21372,N_20768,N_20795);
nand U21373 (N_21373,N_20687,N_20996);
and U21374 (N_21374,N_20982,N_20880);
and U21375 (N_21375,N_20549,N_20809);
nand U21376 (N_21376,N_20762,N_20728);
nor U21377 (N_21377,N_20682,N_20726);
nor U21378 (N_21378,N_20824,N_20842);
nor U21379 (N_21379,N_20853,N_20632);
and U21380 (N_21380,N_20694,N_20713);
and U21381 (N_21381,N_20990,N_20729);
and U21382 (N_21382,N_20629,N_20733);
nor U21383 (N_21383,N_20802,N_20881);
or U21384 (N_21384,N_20847,N_20906);
or U21385 (N_21385,N_20708,N_20580);
and U21386 (N_21386,N_20662,N_20736);
nor U21387 (N_21387,N_20576,N_20555);
or U21388 (N_21388,N_20939,N_20919);
xnor U21389 (N_21389,N_20743,N_20520);
or U21390 (N_21390,N_20622,N_20984);
or U21391 (N_21391,N_20561,N_20582);
or U21392 (N_21392,N_20721,N_20719);
nor U21393 (N_21393,N_20704,N_20874);
or U21394 (N_21394,N_20754,N_20505);
nor U21395 (N_21395,N_20590,N_20606);
and U21396 (N_21396,N_20804,N_20516);
or U21397 (N_21397,N_20938,N_20655);
nor U21398 (N_21398,N_20584,N_20713);
xor U21399 (N_21399,N_20792,N_20840);
and U21400 (N_21400,N_20673,N_20915);
nand U21401 (N_21401,N_20877,N_20893);
or U21402 (N_21402,N_20765,N_20987);
and U21403 (N_21403,N_20927,N_20596);
xor U21404 (N_21404,N_20962,N_20807);
or U21405 (N_21405,N_20529,N_20591);
nand U21406 (N_21406,N_20872,N_20533);
nand U21407 (N_21407,N_20968,N_20621);
xnor U21408 (N_21408,N_20781,N_20939);
or U21409 (N_21409,N_20922,N_20823);
xor U21410 (N_21410,N_20858,N_20516);
nand U21411 (N_21411,N_20582,N_20811);
xnor U21412 (N_21412,N_20798,N_20742);
or U21413 (N_21413,N_20765,N_20580);
and U21414 (N_21414,N_20666,N_20636);
xor U21415 (N_21415,N_20839,N_20603);
or U21416 (N_21416,N_20710,N_20662);
and U21417 (N_21417,N_20899,N_20745);
or U21418 (N_21418,N_20753,N_20633);
and U21419 (N_21419,N_20953,N_20933);
nor U21420 (N_21420,N_20650,N_20648);
or U21421 (N_21421,N_20818,N_20521);
or U21422 (N_21422,N_20502,N_20866);
nor U21423 (N_21423,N_20650,N_20509);
and U21424 (N_21424,N_20689,N_20839);
xnor U21425 (N_21425,N_20501,N_20671);
nor U21426 (N_21426,N_20918,N_20682);
xnor U21427 (N_21427,N_20984,N_20922);
nand U21428 (N_21428,N_20896,N_20772);
nor U21429 (N_21429,N_20941,N_20818);
and U21430 (N_21430,N_20981,N_20699);
nor U21431 (N_21431,N_20542,N_20968);
or U21432 (N_21432,N_20893,N_20917);
nor U21433 (N_21433,N_20923,N_20556);
and U21434 (N_21434,N_20969,N_20876);
nand U21435 (N_21435,N_20783,N_20639);
xor U21436 (N_21436,N_20933,N_20551);
xnor U21437 (N_21437,N_20525,N_20830);
nand U21438 (N_21438,N_20871,N_20775);
xor U21439 (N_21439,N_20819,N_20660);
xnor U21440 (N_21440,N_20558,N_20626);
nor U21441 (N_21441,N_20745,N_20949);
xnor U21442 (N_21442,N_20990,N_20513);
and U21443 (N_21443,N_20997,N_20830);
and U21444 (N_21444,N_20891,N_20828);
nand U21445 (N_21445,N_20939,N_20898);
xnor U21446 (N_21446,N_20882,N_20663);
and U21447 (N_21447,N_20784,N_20930);
xor U21448 (N_21448,N_20896,N_20835);
or U21449 (N_21449,N_20856,N_20779);
nor U21450 (N_21450,N_20516,N_20965);
nor U21451 (N_21451,N_20765,N_20532);
nand U21452 (N_21452,N_20788,N_20799);
xnor U21453 (N_21453,N_20512,N_20878);
and U21454 (N_21454,N_20705,N_20809);
and U21455 (N_21455,N_20633,N_20942);
xnor U21456 (N_21456,N_20700,N_20851);
or U21457 (N_21457,N_20695,N_20616);
nor U21458 (N_21458,N_20525,N_20694);
xor U21459 (N_21459,N_20700,N_20520);
xnor U21460 (N_21460,N_20628,N_20956);
nand U21461 (N_21461,N_20538,N_20896);
nor U21462 (N_21462,N_20963,N_20741);
and U21463 (N_21463,N_20731,N_20629);
nand U21464 (N_21464,N_20632,N_20704);
nand U21465 (N_21465,N_20726,N_20889);
and U21466 (N_21466,N_20625,N_20785);
nand U21467 (N_21467,N_20832,N_20650);
and U21468 (N_21468,N_20608,N_20987);
and U21469 (N_21469,N_20545,N_20992);
and U21470 (N_21470,N_20516,N_20787);
nand U21471 (N_21471,N_20714,N_20683);
nand U21472 (N_21472,N_20851,N_20720);
xor U21473 (N_21473,N_20866,N_20500);
or U21474 (N_21474,N_20596,N_20797);
nand U21475 (N_21475,N_20965,N_20730);
and U21476 (N_21476,N_20767,N_20726);
nand U21477 (N_21477,N_20854,N_20596);
and U21478 (N_21478,N_20665,N_20518);
nor U21479 (N_21479,N_20576,N_20672);
or U21480 (N_21480,N_20690,N_20878);
nand U21481 (N_21481,N_20768,N_20817);
nand U21482 (N_21482,N_20594,N_20515);
nor U21483 (N_21483,N_20531,N_20794);
and U21484 (N_21484,N_20658,N_20788);
nand U21485 (N_21485,N_20897,N_20951);
xor U21486 (N_21486,N_20617,N_20755);
nand U21487 (N_21487,N_20541,N_20537);
nand U21488 (N_21488,N_20942,N_20577);
and U21489 (N_21489,N_20969,N_20842);
or U21490 (N_21490,N_20890,N_20686);
xor U21491 (N_21491,N_20742,N_20711);
nand U21492 (N_21492,N_20993,N_20755);
or U21493 (N_21493,N_20916,N_20556);
xnor U21494 (N_21494,N_20765,N_20913);
nor U21495 (N_21495,N_20554,N_20952);
or U21496 (N_21496,N_20767,N_20902);
or U21497 (N_21497,N_20668,N_20939);
nor U21498 (N_21498,N_20803,N_20556);
nand U21499 (N_21499,N_20632,N_20625);
or U21500 (N_21500,N_21258,N_21133);
xnor U21501 (N_21501,N_21186,N_21227);
nor U21502 (N_21502,N_21047,N_21490);
nand U21503 (N_21503,N_21156,N_21089);
or U21504 (N_21504,N_21287,N_21494);
nor U21505 (N_21505,N_21348,N_21074);
xor U21506 (N_21506,N_21273,N_21106);
xor U21507 (N_21507,N_21040,N_21275);
nor U21508 (N_21508,N_21470,N_21192);
nand U21509 (N_21509,N_21063,N_21367);
or U21510 (N_21510,N_21230,N_21324);
nor U21511 (N_21511,N_21184,N_21366);
and U21512 (N_21512,N_21267,N_21244);
and U21513 (N_21513,N_21263,N_21140);
nor U21514 (N_21514,N_21034,N_21315);
nor U21515 (N_21515,N_21412,N_21319);
xor U21516 (N_21516,N_21357,N_21262);
or U21517 (N_21517,N_21487,N_21188);
nor U21518 (N_21518,N_21172,N_21045);
nand U21519 (N_21519,N_21334,N_21284);
nand U21520 (N_21520,N_21007,N_21092);
xor U21521 (N_21521,N_21223,N_21243);
or U21522 (N_21522,N_21392,N_21087);
xor U21523 (N_21523,N_21467,N_21277);
or U21524 (N_21524,N_21351,N_21143);
nand U21525 (N_21525,N_21113,N_21157);
or U21526 (N_21526,N_21163,N_21030);
and U21527 (N_21527,N_21228,N_21199);
xor U21528 (N_21528,N_21441,N_21096);
nor U21529 (N_21529,N_21265,N_21046);
or U21530 (N_21530,N_21354,N_21397);
and U21531 (N_21531,N_21497,N_21373);
xor U21532 (N_21532,N_21274,N_21110);
xor U21533 (N_21533,N_21136,N_21235);
or U21534 (N_21534,N_21291,N_21396);
or U21535 (N_21535,N_21406,N_21128);
nand U21536 (N_21536,N_21158,N_21003);
nand U21537 (N_21537,N_21342,N_21290);
or U21538 (N_21538,N_21031,N_21381);
or U21539 (N_21539,N_21299,N_21219);
xor U21540 (N_21540,N_21304,N_21463);
or U21541 (N_21541,N_21292,N_21245);
and U21542 (N_21542,N_21439,N_21403);
or U21543 (N_21543,N_21043,N_21481);
and U21544 (N_21544,N_21356,N_21402);
xnor U21545 (N_21545,N_21401,N_21187);
nor U21546 (N_21546,N_21075,N_21301);
and U21547 (N_21547,N_21122,N_21177);
xor U21548 (N_21548,N_21281,N_21496);
nand U21549 (N_21549,N_21100,N_21293);
or U21550 (N_21550,N_21220,N_21196);
and U21551 (N_21551,N_21314,N_21430);
and U21552 (N_21552,N_21460,N_21035);
and U21553 (N_21553,N_21057,N_21221);
xnor U21554 (N_21554,N_21288,N_21384);
and U21555 (N_21555,N_21021,N_21005);
nor U21556 (N_21556,N_21261,N_21447);
xor U21557 (N_21557,N_21414,N_21058);
nand U21558 (N_21558,N_21056,N_21099);
or U21559 (N_21559,N_21339,N_21138);
and U21560 (N_21560,N_21112,N_21103);
nand U21561 (N_21561,N_21251,N_21226);
and U21562 (N_21562,N_21377,N_21407);
nor U21563 (N_21563,N_21194,N_21480);
xor U21564 (N_21564,N_21395,N_21182);
nand U21565 (N_21565,N_21476,N_21197);
xor U21566 (N_21566,N_21130,N_21474);
or U21567 (N_21567,N_21424,N_21294);
xnor U21568 (N_21568,N_21359,N_21303);
nor U21569 (N_21569,N_21264,N_21149);
nor U21570 (N_21570,N_21067,N_21323);
xnor U21571 (N_21571,N_21239,N_21446);
or U21572 (N_21572,N_21038,N_21069);
and U21573 (N_21573,N_21093,N_21449);
nand U21574 (N_21574,N_21091,N_21493);
nand U21575 (N_21575,N_21062,N_21410);
xnor U21576 (N_21576,N_21012,N_21164);
or U21577 (N_21577,N_21152,N_21204);
xnor U21578 (N_21578,N_21327,N_21451);
or U21579 (N_21579,N_21079,N_21380);
or U21580 (N_21580,N_21455,N_21139);
xor U21581 (N_21581,N_21166,N_21066);
nor U21582 (N_21582,N_21499,N_21257);
xnor U21583 (N_21583,N_21161,N_21020);
xnor U21584 (N_21584,N_21478,N_21145);
nor U21585 (N_21585,N_21232,N_21286);
and U21586 (N_21586,N_21346,N_21160);
nand U21587 (N_21587,N_21417,N_21428);
nor U21588 (N_21588,N_21162,N_21159);
nor U21589 (N_21589,N_21386,N_21173);
or U21590 (N_21590,N_21071,N_21391);
nor U21591 (N_21591,N_21083,N_21489);
nor U21592 (N_21592,N_21084,N_21080);
nor U21593 (N_21593,N_21378,N_21408);
xnor U21594 (N_21594,N_21015,N_21124);
xnor U21595 (N_21595,N_21036,N_21399);
xor U21596 (N_21596,N_21060,N_21114);
and U21597 (N_21597,N_21423,N_21437);
and U21598 (N_21598,N_21216,N_21416);
or U21599 (N_21599,N_21049,N_21448);
nand U21600 (N_21600,N_21340,N_21413);
nand U21601 (N_21601,N_21338,N_21374);
xor U21602 (N_21602,N_21129,N_21026);
or U21603 (N_21603,N_21210,N_21425);
or U21604 (N_21604,N_21300,N_21024);
nor U21605 (N_21605,N_21125,N_21253);
xor U21606 (N_21606,N_21311,N_21462);
or U21607 (N_21607,N_21330,N_21211);
xor U21608 (N_21608,N_21233,N_21120);
nor U21609 (N_21609,N_21217,N_21440);
and U21610 (N_21610,N_21055,N_21006);
and U21611 (N_21611,N_21370,N_21222);
nor U21612 (N_21612,N_21104,N_21332);
nor U21613 (N_21613,N_21061,N_21382);
nor U21614 (N_21614,N_21247,N_21102);
and U21615 (N_21615,N_21355,N_21432);
nand U21616 (N_21616,N_21353,N_21337);
xor U21617 (N_21617,N_21132,N_21486);
and U21618 (N_21618,N_21011,N_21419);
xor U21619 (N_21619,N_21385,N_21242);
nand U21620 (N_21620,N_21297,N_21023);
xnor U21621 (N_21621,N_21053,N_21450);
nor U21622 (N_21622,N_21185,N_21404);
nor U21623 (N_21623,N_21051,N_21420);
nor U21624 (N_21624,N_21014,N_21305);
nor U21625 (N_21625,N_21405,N_21485);
xnor U21626 (N_21626,N_21170,N_21224);
or U21627 (N_21627,N_21065,N_21289);
or U21628 (N_21628,N_21189,N_21333);
xor U21629 (N_21629,N_21059,N_21434);
or U21630 (N_21630,N_21318,N_21421);
xor U21631 (N_21631,N_21119,N_21218);
or U21632 (N_21632,N_21167,N_21109);
or U21633 (N_21633,N_21394,N_21002);
or U21634 (N_21634,N_21042,N_21376);
and U21635 (N_21635,N_21190,N_21271);
and U21636 (N_21636,N_21438,N_21176);
nor U21637 (N_21637,N_21256,N_21295);
or U21638 (N_21638,N_21017,N_21302);
nand U21639 (N_21639,N_21238,N_21459);
or U21640 (N_21640,N_21081,N_21442);
and U21641 (N_21641,N_21313,N_21389);
and U21642 (N_21642,N_21360,N_21473);
or U21643 (N_21643,N_21078,N_21212);
xor U21644 (N_21644,N_21214,N_21453);
nor U21645 (N_21645,N_21137,N_21350);
or U21646 (N_21646,N_21019,N_21475);
nand U21647 (N_21647,N_21008,N_21308);
and U21648 (N_21648,N_21483,N_21431);
and U21649 (N_21649,N_21082,N_21037);
nand U21650 (N_21650,N_21252,N_21387);
and U21651 (N_21651,N_21362,N_21029);
xnor U21652 (N_21652,N_21200,N_21269);
nand U21653 (N_21653,N_21076,N_21179);
nand U21654 (N_21654,N_21321,N_21072);
nand U21655 (N_21655,N_21142,N_21155);
or U21656 (N_21656,N_21325,N_21458);
or U21657 (N_21657,N_21372,N_21181);
nor U21658 (N_21658,N_21183,N_21205);
and U21659 (N_21659,N_21168,N_21436);
or U21660 (N_21660,N_21379,N_21369);
nor U21661 (N_21661,N_21280,N_21479);
xnor U21662 (N_21662,N_21326,N_21443);
xnor U21663 (N_21663,N_21203,N_21328);
xnor U21664 (N_21664,N_21296,N_21260);
and U21665 (N_21665,N_21121,N_21016);
and U21666 (N_21666,N_21468,N_21010);
nor U21667 (N_21667,N_21285,N_21236);
or U21668 (N_21668,N_21371,N_21118);
and U21669 (N_21669,N_21278,N_21141);
and U21670 (N_21670,N_21433,N_21202);
and U21671 (N_21671,N_21033,N_21209);
or U21672 (N_21672,N_21070,N_21495);
or U21673 (N_21673,N_21469,N_21178);
or U21674 (N_21674,N_21364,N_21358);
xor U21675 (N_21675,N_21231,N_21270);
xor U21676 (N_21676,N_21312,N_21477);
and U21677 (N_21677,N_21482,N_21409);
xor U21678 (N_21678,N_21268,N_21101);
nand U21679 (N_21679,N_21307,N_21094);
and U21680 (N_21680,N_21427,N_21426);
and U21681 (N_21681,N_21259,N_21054);
nand U21682 (N_21682,N_21279,N_21422);
nand U21683 (N_21683,N_21208,N_21498);
or U21684 (N_21684,N_21464,N_21491);
nand U21685 (N_21685,N_21175,N_21393);
nand U21686 (N_21686,N_21435,N_21388);
and U21687 (N_21687,N_21456,N_21098);
nor U21688 (N_21688,N_21336,N_21365);
nand U21689 (N_21689,N_21452,N_21032);
nor U21690 (N_21690,N_21317,N_21335);
or U21691 (N_21691,N_21241,N_21283);
or U21692 (N_21692,N_21400,N_21329);
xnor U21693 (N_21693,N_21115,N_21193);
and U21694 (N_21694,N_21492,N_21028);
nor U21695 (N_21695,N_21225,N_21272);
nor U21696 (N_21696,N_21174,N_21255);
xnor U21697 (N_21697,N_21249,N_21151);
nand U21698 (N_21698,N_21086,N_21383);
and U21699 (N_21699,N_21237,N_21198);
nand U21700 (N_21700,N_21165,N_21107);
or U21701 (N_21701,N_21309,N_21466);
and U21702 (N_21702,N_21316,N_21363);
or U21703 (N_21703,N_21331,N_21123);
xor U21704 (N_21704,N_21310,N_21117);
nor U21705 (N_21705,N_21146,N_21429);
nor U21706 (N_21706,N_21052,N_21013);
nor U21707 (N_21707,N_21484,N_21009);
and U21708 (N_21708,N_21077,N_21215);
and U21709 (N_21709,N_21134,N_21108);
xor U21710 (N_21710,N_21144,N_21105);
nor U21711 (N_21711,N_21097,N_21457);
nand U21712 (N_21712,N_21191,N_21068);
xnor U21713 (N_21713,N_21116,N_21488);
and U21714 (N_21714,N_21344,N_21111);
nand U21715 (N_21715,N_21246,N_21298);
and U21716 (N_21716,N_21085,N_21411);
nor U21717 (N_21717,N_21126,N_21254);
xor U21718 (N_21718,N_21169,N_21234);
and U21719 (N_21719,N_21361,N_21090);
xor U21720 (N_21720,N_21154,N_21282);
nand U21721 (N_21721,N_21000,N_21150);
nand U21722 (N_21722,N_21050,N_21064);
and U21723 (N_21723,N_21320,N_21375);
nor U21724 (N_21724,N_21472,N_21127);
and U21725 (N_21725,N_21471,N_21347);
xor U21726 (N_21726,N_21195,N_21206);
or U21727 (N_21727,N_21343,N_21322);
xnor U21728 (N_21728,N_21153,N_21004);
and U21729 (N_21729,N_21341,N_21018);
or U21730 (N_21730,N_21465,N_21131);
or U21731 (N_21731,N_21171,N_21418);
nand U21732 (N_21732,N_21135,N_21445);
or U21733 (N_21733,N_21461,N_21266);
xor U21734 (N_21734,N_21276,N_21454);
nand U21735 (N_21735,N_21088,N_21027);
or U21736 (N_21736,N_21044,N_21001);
and U21737 (N_21737,N_21390,N_21398);
or U21738 (N_21738,N_21240,N_21095);
xor U21739 (N_21739,N_21345,N_21147);
nand U21740 (N_21740,N_21250,N_21349);
and U21741 (N_21741,N_21415,N_21041);
nand U21742 (N_21742,N_21352,N_21207);
and U21743 (N_21743,N_21368,N_21025);
nand U21744 (N_21744,N_21201,N_21229);
or U21745 (N_21745,N_21180,N_21444);
or U21746 (N_21746,N_21306,N_21248);
xnor U21747 (N_21747,N_21022,N_21039);
nand U21748 (N_21748,N_21048,N_21148);
xor U21749 (N_21749,N_21073,N_21213);
nand U21750 (N_21750,N_21450,N_21003);
nand U21751 (N_21751,N_21364,N_21210);
or U21752 (N_21752,N_21322,N_21175);
and U21753 (N_21753,N_21340,N_21251);
and U21754 (N_21754,N_21467,N_21037);
or U21755 (N_21755,N_21473,N_21314);
and U21756 (N_21756,N_21330,N_21439);
and U21757 (N_21757,N_21198,N_21348);
xor U21758 (N_21758,N_21499,N_21071);
nand U21759 (N_21759,N_21005,N_21220);
nand U21760 (N_21760,N_21188,N_21466);
nand U21761 (N_21761,N_21405,N_21158);
or U21762 (N_21762,N_21423,N_21265);
or U21763 (N_21763,N_21127,N_21014);
nor U21764 (N_21764,N_21077,N_21247);
nand U21765 (N_21765,N_21319,N_21282);
xnor U21766 (N_21766,N_21407,N_21428);
xnor U21767 (N_21767,N_21333,N_21474);
xnor U21768 (N_21768,N_21488,N_21233);
xor U21769 (N_21769,N_21184,N_21079);
or U21770 (N_21770,N_21487,N_21456);
or U21771 (N_21771,N_21339,N_21394);
nand U21772 (N_21772,N_21312,N_21277);
nor U21773 (N_21773,N_21303,N_21127);
nand U21774 (N_21774,N_21023,N_21078);
xnor U21775 (N_21775,N_21011,N_21481);
nor U21776 (N_21776,N_21153,N_21301);
or U21777 (N_21777,N_21400,N_21360);
nor U21778 (N_21778,N_21168,N_21351);
nor U21779 (N_21779,N_21296,N_21319);
or U21780 (N_21780,N_21274,N_21001);
xor U21781 (N_21781,N_21487,N_21060);
nand U21782 (N_21782,N_21131,N_21026);
nand U21783 (N_21783,N_21054,N_21196);
xor U21784 (N_21784,N_21138,N_21247);
or U21785 (N_21785,N_21035,N_21264);
and U21786 (N_21786,N_21036,N_21491);
or U21787 (N_21787,N_21407,N_21190);
nor U21788 (N_21788,N_21119,N_21283);
and U21789 (N_21789,N_21225,N_21421);
nand U21790 (N_21790,N_21381,N_21465);
xor U21791 (N_21791,N_21118,N_21047);
xnor U21792 (N_21792,N_21378,N_21362);
xnor U21793 (N_21793,N_21467,N_21044);
xnor U21794 (N_21794,N_21169,N_21250);
xor U21795 (N_21795,N_21107,N_21409);
and U21796 (N_21796,N_21221,N_21198);
and U21797 (N_21797,N_21085,N_21366);
nand U21798 (N_21798,N_21412,N_21464);
nand U21799 (N_21799,N_21109,N_21118);
nor U21800 (N_21800,N_21353,N_21189);
nor U21801 (N_21801,N_21105,N_21461);
nand U21802 (N_21802,N_21291,N_21023);
nand U21803 (N_21803,N_21475,N_21063);
nor U21804 (N_21804,N_21405,N_21027);
nor U21805 (N_21805,N_21237,N_21323);
and U21806 (N_21806,N_21339,N_21232);
nand U21807 (N_21807,N_21101,N_21266);
nor U21808 (N_21808,N_21265,N_21019);
nor U21809 (N_21809,N_21103,N_21402);
xor U21810 (N_21810,N_21306,N_21253);
or U21811 (N_21811,N_21030,N_21302);
and U21812 (N_21812,N_21463,N_21407);
nand U21813 (N_21813,N_21178,N_21248);
nand U21814 (N_21814,N_21100,N_21159);
and U21815 (N_21815,N_21027,N_21434);
nand U21816 (N_21816,N_21432,N_21383);
nand U21817 (N_21817,N_21431,N_21375);
xnor U21818 (N_21818,N_21089,N_21225);
and U21819 (N_21819,N_21274,N_21439);
and U21820 (N_21820,N_21292,N_21074);
nand U21821 (N_21821,N_21099,N_21067);
nand U21822 (N_21822,N_21321,N_21250);
nand U21823 (N_21823,N_21481,N_21444);
nor U21824 (N_21824,N_21371,N_21134);
or U21825 (N_21825,N_21477,N_21017);
or U21826 (N_21826,N_21102,N_21410);
or U21827 (N_21827,N_21084,N_21019);
or U21828 (N_21828,N_21258,N_21456);
xnor U21829 (N_21829,N_21392,N_21318);
or U21830 (N_21830,N_21385,N_21437);
nor U21831 (N_21831,N_21114,N_21083);
nand U21832 (N_21832,N_21259,N_21020);
and U21833 (N_21833,N_21046,N_21378);
nor U21834 (N_21834,N_21462,N_21123);
nor U21835 (N_21835,N_21111,N_21440);
or U21836 (N_21836,N_21498,N_21020);
nor U21837 (N_21837,N_21044,N_21158);
nand U21838 (N_21838,N_21367,N_21175);
nand U21839 (N_21839,N_21153,N_21354);
or U21840 (N_21840,N_21455,N_21321);
xnor U21841 (N_21841,N_21294,N_21276);
nor U21842 (N_21842,N_21305,N_21363);
and U21843 (N_21843,N_21030,N_21258);
nand U21844 (N_21844,N_21405,N_21338);
or U21845 (N_21845,N_21373,N_21165);
nand U21846 (N_21846,N_21342,N_21352);
xnor U21847 (N_21847,N_21203,N_21111);
nand U21848 (N_21848,N_21125,N_21049);
or U21849 (N_21849,N_21467,N_21003);
and U21850 (N_21850,N_21126,N_21120);
xnor U21851 (N_21851,N_21106,N_21168);
nand U21852 (N_21852,N_21264,N_21196);
and U21853 (N_21853,N_21434,N_21072);
xnor U21854 (N_21854,N_21249,N_21038);
nor U21855 (N_21855,N_21048,N_21179);
and U21856 (N_21856,N_21071,N_21431);
xor U21857 (N_21857,N_21465,N_21481);
or U21858 (N_21858,N_21128,N_21078);
nor U21859 (N_21859,N_21204,N_21248);
nor U21860 (N_21860,N_21162,N_21431);
and U21861 (N_21861,N_21094,N_21244);
or U21862 (N_21862,N_21497,N_21167);
nand U21863 (N_21863,N_21455,N_21077);
and U21864 (N_21864,N_21384,N_21337);
and U21865 (N_21865,N_21023,N_21471);
nor U21866 (N_21866,N_21467,N_21429);
xnor U21867 (N_21867,N_21430,N_21388);
nand U21868 (N_21868,N_21384,N_21356);
and U21869 (N_21869,N_21459,N_21273);
nor U21870 (N_21870,N_21475,N_21406);
and U21871 (N_21871,N_21383,N_21148);
nor U21872 (N_21872,N_21223,N_21006);
nand U21873 (N_21873,N_21152,N_21112);
and U21874 (N_21874,N_21427,N_21421);
xor U21875 (N_21875,N_21158,N_21157);
nand U21876 (N_21876,N_21118,N_21466);
nor U21877 (N_21877,N_21343,N_21279);
and U21878 (N_21878,N_21496,N_21009);
or U21879 (N_21879,N_21356,N_21212);
nand U21880 (N_21880,N_21362,N_21409);
or U21881 (N_21881,N_21498,N_21258);
nor U21882 (N_21882,N_21225,N_21118);
and U21883 (N_21883,N_21219,N_21245);
xnor U21884 (N_21884,N_21406,N_21126);
and U21885 (N_21885,N_21122,N_21239);
xnor U21886 (N_21886,N_21111,N_21126);
nand U21887 (N_21887,N_21484,N_21358);
or U21888 (N_21888,N_21419,N_21347);
xnor U21889 (N_21889,N_21409,N_21474);
nor U21890 (N_21890,N_21046,N_21254);
or U21891 (N_21891,N_21202,N_21258);
nand U21892 (N_21892,N_21383,N_21205);
xnor U21893 (N_21893,N_21197,N_21115);
xor U21894 (N_21894,N_21129,N_21359);
xnor U21895 (N_21895,N_21346,N_21126);
nor U21896 (N_21896,N_21461,N_21406);
or U21897 (N_21897,N_21432,N_21137);
xnor U21898 (N_21898,N_21357,N_21405);
and U21899 (N_21899,N_21444,N_21220);
and U21900 (N_21900,N_21103,N_21392);
or U21901 (N_21901,N_21240,N_21158);
or U21902 (N_21902,N_21403,N_21324);
xor U21903 (N_21903,N_21262,N_21044);
nand U21904 (N_21904,N_21491,N_21288);
nor U21905 (N_21905,N_21240,N_21384);
xor U21906 (N_21906,N_21129,N_21211);
and U21907 (N_21907,N_21291,N_21269);
or U21908 (N_21908,N_21314,N_21300);
and U21909 (N_21909,N_21438,N_21187);
or U21910 (N_21910,N_21376,N_21161);
nand U21911 (N_21911,N_21343,N_21495);
or U21912 (N_21912,N_21248,N_21197);
nor U21913 (N_21913,N_21103,N_21044);
xnor U21914 (N_21914,N_21056,N_21483);
nand U21915 (N_21915,N_21294,N_21286);
xor U21916 (N_21916,N_21023,N_21152);
or U21917 (N_21917,N_21389,N_21201);
nor U21918 (N_21918,N_21206,N_21273);
nor U21919 (N_21919,N_21203,N_21469);
xnor U21920 (N_21920,N_21279,N_21209);
and U21921 (N_21921,N_21169,N_21325);
xnor U21922 (N_21922,N_21320,N_21152);
or U21923 (N_21923,N_21386,N_21451);
and U21924 (N_21924,N_21360,N_21009);
or U21925 (N_21925,N_21225,N_21492);
and U21926 (N_21926,N_21228,N_21305);
or U21927 (N_21927,N_21307,N_21435);
or U21928 (N_21928,N_21433,N_21240);
nor U21929 (N_21929,N_21126,N_21495);
nor U21930 (N_21930,N_21038,N_21131);
or U21931 (N_21931,N_21353,N_21417);
and U21932 (N_21932,N_21180,N_21135);
and U21933 (N_21933,N_21298,N_21343);
xor U21934 (N_21934,N_21049,N_21072);
xor U21935 (N_21935,N_21118,N_21032);
nor U21936 (N_21936,N_21337,N_21155);
and U21937 (N_21937,N_21019,N_21043);
nand U21938 (N_21938,N_21010,N_21185);
or U21939 (N_21939,N_21302,N_21435);
nand U21940 (N_21940,N_21473,N_21380);
or U21941 (N_21941,N_21345,N_21154);
nand U21942 (N_21942,N_21006,N_21451);
or U21943 (N_21943,N_21439,N_21326);
and U21944 (N_21944,N_21162,N_21225);
nand U21945 (N_21945,N_21212,N_21436);
and U21946 (N_21946,N_21489,N_21068);
and U21947 (N_21947,N_21412,N_21269);
xnor U21948 (N_21948,N_21302,N_21485);
or U21949 (N_21949,N_21038,N_21117);
and U21950 (N_21950,N_21184,N_21492);
and U21951 (N_21951,N_21149,N_21292);
nand U21952 (N_21952,N_21295,N_21467);
and U21953 (N_21953,N_21249,N_21480);
nor U21954 (N_21954,N_21365,N_21183);
nor U21955 (N_21955,N_21017,N_21056);
and U21956 (N_21956,N_21120,N_21141);
or U21957 (N_21957,N_21168,N_21298);
and U21958 (N_21958,N_21035,N_21044);
nand U21959 (N_21959,N_21249,N_21054);
nand U21960 (N_21960,N_21170,N_21281);
nor U21961 (N_21961,N_21036,N_21489);
nand U21962 (N_21962,N_21000,N_21493);
nand U21963 (N_21963,N_21008,N_21066);
and U21964 (N_21964,N_21254,N_21319);
or U21965 (N_21965,N_21350,N_21434);
and U21966 (N_21966,N_21491,N_21424);
nor U21967 (N_21967,N_21124,N_21341);
xnor U21968 (N_21968,N_21499,N_21214);
nand U21969 (N_21969,N_21409,N_21329);
or U21970 (N_21970,N_21438,N_21049);
or U21971 (N_21971,N_21378,N_21139);
xnor U21972 (N_21972,N_21165,N_21398);
or U21973 (N_21973,N_21219,N_21139);
nor U21974 (N_21974,N_21433,N_21061);
nor U21975 (N_21975,N_21138,N_21415);
or U21976 (N_21976,N_21013,N_21257);
and U21977 (N_21977,N_21234,N_21032);
nor U21978 (N_21978,N_21116,N_21315);
nor U21979 (N_21979,N_21159,N_21054);
xor U21980 (N_21980,N_21444,N_21428);
nand U21981 (N_21981,N_21015,N_21051);
xnor U21982 (N_21982,N_21365,N_21011);
and U21983 (N_21983,N_21077,N_21376);
nand U21984 (N_21984,N_21107,N_21357);
and U21985 (N_21985,N_21111,N_21350);
nand U21986 (N_21986,N_21226,N_21308);
xnor U21987 (N_21987,N_21491,N_21414);
nand U21988 (N_21988,N_21402,N_21106);
nor U21989 (N_21989,N_21411,N_21090);
nor U21990 (N_21990,N_21413,N_21230);
and U21991 (N_21991,N_21301,N_21167);
nor U21992 (N_21992,N_21190,N_21334);
nand U21993 (N_21993,N_21356,N_21337);
or U21994 (N_21994,N_21063,N_21257);
nand U21995 (N_21995,N_21070,N_21076);
xor U21996 (N_21996,N_21174,N_21433);
xnor U21997 (N_21997,N_21365,N_21467);
nand U21998 (N_21998,N_21458,N_21316);
xnor U21999 (N_21999,N_21055,N_21287);
xnor U22000 (N_22000,N_21892,N_21901);
xnor U22001 (N_22001,N_21916,N_21598);
or U22002 (N_22002,N_21702,N_21987);
xor U22003 (N_22003,N_21692,N_21971);
xor U22004 (N_22004,N_21801,N_21739);
or U22005 (N_22005,N_21504,N_21796);
or U22006 (N_22006,N_21605,N_21622);
nor U22007 (N_22007,N_21663,N_21867);
nand U22008 (N_22008,N_21929,N_21868);
or U22009 (N_22009,N_21920,N_21958);
xor U22010 (N_22010,N_21675,N_21523);
nor U22011 (N_22011,N_21764,N_21545);
and U22012 (N_22012,N_21679,N_21777);
and U22013 (N_22013,N_21577,N_21888);
nor U22014 (N_22014,N_21625,N_21891);
or U22015 (N_22015,N_21590,N_21832);
nor U22016 (N_22016,N_21544,N_21695);
xor U22017 (N_22017,N_21610,N_21951);
and U22018 (N_22018,N_21861,N_21542);
and U22019 (N_22019,N_21696,N_21841);
xnor U22020 (N_22020,N_21503,N_21532);
xnor U22021 (N_22021,N_21849,N_21816);
nor U22022 (N_22022,N_21961,N_21694);
or U22023 (N_22023,N_21875,N_21838);
nor U22024 (N_22024,N_21613,N_21923);
nand U22025 (N_22025,N_21632,N_21895);
nand U22026 (N_22026,N_21986,N_21509);
nor U22027 (N_22027,N_21778,N_21771);
nand U22028 (N_22028,N_21927,N_21877);
xor U22029 (N_22029,N_21755,N_21941);
or U22030 (N_22030,N_21546,N_21568);
nor U22031 (N_22031,N_21804,N_21900);
nand U22032 (N_22032,N_21786,N_21751);
nor U22033 (N_22033,N_21797,N_21818);
xor U22034 (N_22034,N_21713,N_21752);
xnor U22035 (N_22035,N_21767,N_21683);
or U22036 (N_22036,N_21904,N_21762);
and U22037 (N_22037,N_21670,N_21588);
or U22038 (N_22038,N_21745,N_21833);
nor U22039 (N_22039,N_21788,N_21933);
nand U22040 (N_22040,N_21894,N_21700);
and U22041 (N_22041,N_21939,N_21729);
nand U22042 (N_22042,N_21822,N_21530);
and U22043 (N_22043,N_21705,N_21826);
nor U22044 (N_22044,N_21698,N_21650);
nor U22045 (N_22045,N_21671,N_21528);
xnor U22046 (N_22046,N_21918,N_21960);
nor U22047 (N_22047,N_21585,N_21810);
or U22048 (N_22048,N_21653,N_21554);
and U22049 (N_22049,N_21737,N_21773);
nand U22050 (N_22050,N_21828,N_21708);
nor U22051 (N_22051,N_21899,N_21648);
and U22052 (N_22052,N_21850,N_21594);
nand U22053 (N_22053,N_21903,N_21743);
nor U22054 (N_22054,N_21944,N_21834);
nor U22055 (N_22055,N_21835,N_21732);
nor U22056 (N_22056,N_21586,N_21946);
nand U22057 (N_22057,N_21574,N_21725);
xnor U22058 (N_22058,N_21534,N_21657);
nor U22059 (N_22059,N_21748,N_21945);
xor U22060 (N_22060,N_21689,N_21513);
and U22061 (N_22061,N_21765,N_21561);
and U22062 (N_22062,N_21703,N_21995);
or U22063 (N_22063,N_21589,N_21966);
and U22064 (N_22064,N_21953,N_21690);
and U22065 (N_22065,N_21618,N_21579);
nand U22066 (N_22066,N_21550,N_21631);
nor U22067 (N_22067,N_21831,N_21520);
nand U22068 (N_22068,N_21514,N_21967);
xor U22069 (N_22069,N_21993,N_21516);
and U22070 (N_22070,N_21769,N_21515);
and U22071 (N_22071,N_21932,N_21608);
xnor U22072 (N_22072,N_21790,N_21633);
and U22073 (N_22073,N_21569,N_21580);
nand U22074 (N_22074,N_21720,N_21910);
nand U22075 (N_22075,N_21518,N_21936);
nand U22076 (N_22076,N_21726,N_21662);
nand U22077 (N_22077,N_21872,N_21972);
and U22078 (N_22078,N_21836,N_21807);
nor U22079 (N_22079,N_21661,N_21922);
xnor U22080 (N_22080,N_21623,N_21738);
or U22081 (N_22081,N_21697,N_21510);
nand U22082 (N_22082,N_21549,N_21652);
nor U22083 (N_22083,N_21915,N_21768);
and U22084 (N_22084,N_21978,N_21604);
or U22085 (N_22085,N_21666,N_21913);
nor U22086 (N_22086,N_21638,N_21563);
nor U22087 (N_22087,N_21969,N_21815);
nor U22088 (N_22088,N_21844,N_21667);
and U22089 (N_22089,N_21674,N_21654);
nand U22090 (N_22090,N_21805,N_21879);
or U22091 (N_22091,N_21687,N_21820);
and U22092 (N_22092,N_21706,N_21587);
nand U22093 (N_22093,N_21621,N_21656);
xnor U22094 (N_22094,N_21791,N_21583);
xor U22095 (N_22095,N_21814,N_21572);
nand U22096 (N_22096,N_21789,N_21780);
xnor U22097 (N_22097,N_21505,N_21741);
nand U22098 (N_22098,N_21564,N_21887);
xor U22099 (N_22099,N_21880,N_21883);
nand U22100 (N_22100,N_21606,N_21691);
nand U22101 (N_22101,N_21540,N_21859);
and U22102 (N_22102,N_21924,N_21938);
and U22103 (N_22103,N_21824,N_21851);
nor U22104 (N_22104,N_21957,N_21723);
xor U22105 (N_22105,N_21931,N_21792);
or U22106 (N_22106,N_21533,N_21535);
or U22107 (N_22107,N_21842,N_21658);
nand U22108 (N_22108,N_21827,N_21673);
or U22109 (N_22109,N_21556,N_21878);
xnor U22110 (N_22110,N_21750,N_21857);
nor U22111 (N_22111,N_21906,N_21940);
and U22112 (N_22112,N_21963,N_21862);
xor U22113 (N_22113,N_21665,N_21521);
and U22114 (N_22114,N_21812,N_21949);
xnor U22115 (N_22115,N_21717,N_21562);
or U22116 (N_22116,N_21800,N_21507);
nor U22117 (N_22117,N_21529,N_21893);
and U22118 (N_22118,N_21512,N_21950);
and U22119 (N_22119,N_21813,N_21886);
or U22120 (N_22120,N_21640,N_21964);
nor U22121 (N_22121,N_21624,N_21566);
and U22122 (N_22122,N_21871,N_21643);
nand U22123 (N_22123,N_21716,N_21655);
xnor U22124 (N_22124,N_21526,N_21746);
xor U22125 (N_22125,N_21710,N_21537);
xor U22126 (N_22126,N_21912,N_21798);
or U22127 (N_22127,N_21869,N_21576);
nand U22128 (N_22128,N_21582,N_21669);
xnor U22129 (N_22129,N_21551,N_21500);
or U22130 (N_22130,N_21926,N_21793);
xor U22131 (N_22131,N_21553,N_21991);
nand U22132 (N_22132,N_21601,N_21609);
or U22133 (N_22133,N_21845,N_21627);
and U22134 (N_22134,N_21517,N_21629);
nor U22135 (N_22135,N_21506,N_21644);
nor U22136 (N_22136,N_21909,N_21712);
nor U22137 (N_22137,N_21763,N_21637);
xor U22138 (N_22138,N_21955,N_21602);
nor U22139 (N_22139,N_21616,N_21681);
nor U22140 (N_22140,N_21908,N_21635);
nor U22141 (N_22141,N_21928,N_21647);
xor U22142 (N_22142,N_21715,N_21646);
xnor U22143 (N_22143,N_21704,N_21885);
or U22144 (N_22144,N_21890,N_21809);
or U22145 (N_22145,N_21701,N_21942);
nor U22146 (N_22146,N_21573,N_21558);
and U22147 (N_22147,N_21758,N_21848);
nand U22148 (N_22148,N_21559,N_21853);
nor U22149 (N_22149,N_21668,N_21817);
nand U22150 (N_22150,N_21593,N_21992);
nand U22151 (N_22151,N_21952,N_21921);
or U22152 (N_22152,N_21840,N_21592);
and U22153 (N_22153,N_21795,N_21688);
nand U22154 (N_22154,N_21947,N_21975);
or U22155 (N_22155,N_21979,N_21787);
nor U22156 (N_22156,N_21754,N_21782);
nor U22157 (N_22157,N_21854,N_21897);
nand U22158 (N_22158,N_21808,N_21578);
xor U22159 (N_22159,N_21742,N_21989);
nand U22160 (N_22160,N_21990,N_21772);
or U22161 (N_22161,N_21948,N_21902);
or U22162 (N_22162,N_21898,N_21676);
nand U22163 (N_22163,N_21959,N_21736);
and U22164 (N_22164,N_21996,N_21802);
nor U22165 (N_22165,N_21628,N_21930);
nor U22166 (N_22166,N_21855,N_21649);
nor U22167 (N_22167,N_21994,N_21599);
nand U22168 (N_22168,N_21719,N_21502);
or U22169 (N_22169,N_21718,N_21508);
or U22170 (N_22170,N_21956,N_21735);
nand U22171 (N_22171,N_21864,N_21722);
nand U22172 (N_22172,N_21686,N_21976);
nor U22173 (N_22173,N_21775,N_21575);
or U22174 (N_22174,N_21884,N_21794);
nand U22175 (N_22175,N_21714,N_21660);
nand U22176 (N_22176,N_21830,N_21760);
nand U22177 (N_22177,N_21837,N_21596);
xnor U22178 (N_22178,N_21759,N_21527);
and U22179 (N_22179,N_21501,N_21757);
and U22180 (N_22180,N_21611,N_21684);
xor U22181 (N_22181,N_21614,N_21829);
nand U22182 (N_22182,N_21783,N_21779);
nand U22183 (N_22183,N_21981,N_21825);
or U22184 (N_22184,N_21803,N_21724);
nand U22185 (N_22185,N_21749,N_21597);
or U22186 (N_22186,N_21615,N_21731);
nand U22187 (N_22187,N_21651,N_21744);
nand U22188 (N_22188,N_21531,N_21595);
or U22189 (N_22189,N_21962,N_21896);
nand U22190 (N_22190,N_21699,N_21522);
and U22191 (N_22191,N_21619,N_21740);
and U22192 (N_22192,N_21678,N_21581);
nand U22193 (N_22193,N_21860,N_21747);
and U22194 (N_22194,N_21876,N_21873);
and U22195 (N_22195,N_21911,N_21858);
or U22196 (N_22196,N_21983,N_21823);
nand U22197 (N_22197,N_21811,N_21645);
nand U22198 (N_22198,N_21543,N_21784);
nor U22199 (N_22199,N_21847,N_21766);
and U22200 (N_22200,N_21620,N_21727);
xor U22201 (N_22201,N_21734,N_21925);
or U22202 (N_22202,N_21584,N_21753);
nand U22203 (N_22203,N_21756,N_21560);
or U22204 (N_22204,N_21914,N_21852);
xnor U22205 (N_22205,N_21856,N_21607);
or U22206 (N_22206,N_21672,N_21685);
nor U22207 (N_22207,N_21863,N_21998);
and U22208 (N_22208,N_21571,N_21821);
nand U22209 (N_22209,N_21709,N_21907);
and U22210 (N_22210,N_21935,N_21642);
and U22211 (N_22211,N_21677,N_21937);
and U22212 (N_22212,N_21603,N_21866);
or U22213 (N_22213,N_21693,N_21819);
nand U22214 (N_22214,N_21973,N_21565);
nor U22215 (N_22215,N_21557,N_21519);
nor U22216 (N_22216,N_21785,N_21846);
nor U22217 (N_22217,N_21617,N_21555);
or U22218 (N_22218,N_21980,N_21774);
nand U22219 (N_22219,N_21511,N_21659);
or U22220 (N_22220,N_21707,N_21770);
xnor U22221 (N_22221,N_21977,N_21634);
or U22222 (N_22222,N_21881,N_21965);
and U22223 (N_22223,N_21970,N_21968);
nand U22224 (N_22224,N_21626,N_21711);
or U22225 (N_22225,N_21999,N_21974);
or U22226 (N_22226,N_21641,N_21548);
nand U22227 (N_22227,N_21882,N_21539);
or U22228 (N_22228,N_21761,N_21728);
nand U22229 (N_22229,N_21874,N_21843);
xor U22230 (N_22230,N_21547,N_21567);
xor U22231 (N_22231,N_21591,N_21954);
nand U22232 (N_22232,N_21917,N_21730);
or U22233 (N_22233,N_21682,N_21781);
xor U22234 (N_22234,N_21541,N_21538);
xor U22235 (N_22235,N_21985,N_21919);
nor U22236 (N_22236,N_21664,N_21889);
or U22237 (N_22237,N_21612,N_21905);
nor U22238 (N_22238,N_21680,N_21733);
nand U22239 (N_22239,N_21865,N_21870);
nand U22240 (N_22240,N_21570,N_21639);
nor U22241 (N_22241,N_21636,N_21630);
and U22242 (N_22242,N_21552,N_21600);
or U22243 (N_22243,N_21934,N_21943);
or U22244 (N_22244,N_21988,N_21839);
or U22245 (N_22245,N_21997,N_21721);
xnor U22246 (N_22246,N_21536,N_21984);
or U22247 (N_22247,N_21524,N_21982);
nand U22248 (N_22248,N_21806,N_21799);
xnor U22249 (N_22249,N_21776,N_21525);
nand U22250 (N_22250,N_21576,N_21504);
xor U22251 (N_22251,N_21535,N_21755);
nor U22252 (N_22252,N_21517,N_21692);
and U22253 (N_22253,N_21924,N_21515);
and U22254 (N_22254,N_21511,N_21562);
or U22255 (N_22255,N_21686,N_21764);
nor U22256 (N_22256,N_21579,N_21837);
nand U22257 (N_22257,N_21745,N_21735);
xnor U22258 (N_22258,N_21561,N_21848);
or U22259 (N_22259,N_21898,N_21513);
nor U22260 (N_22260,N_21561,N_21927);
and U22261 (N_22261,N_21621,N_21748);
nand U22262 (N_22262,N_21562,N_21555);
nor U22263 (N_22263,N_21949,N_21679);
or U22264 (N_22264,N_21565,N_21601);
nor U22265 (N_22265,N_21717,N_21667);
xor U22266 (N_22266,N_21671,N_21793);
nor U22267 (N_22267,N_21711,N_21566);
and U22268 (N_22268,N_21649,N_21780);
or U22269 (N_22269,N_21916,N_21836);
and U22270 (N_22270,N_21666,N_21598);
nor U22271 (N_22271,N_21534,N_21565);
xor U22272 (N_22272,N_21855,N_21751);
nor U22273 (N_22273,N_21851,N_21720);
or U22274 (N_22274,N_21706,N_21920);
or U22275 (N_22275,N_21509,N_21703);
and U22276 (N_22276,N_21573,N_21879);
or U22277 (N_22277,N_21924,N_21816);
and U22278 (N_22278,N_21689,N_21657);
nor U22279 (N_22279,N_21997,N_21632);
or U22280 (N_22280,N_21879,N_21803);
nand U22281 (N_22281,N_21726,N_21583);
or U22282 (N_22282,N_21836,N_21629);
xnor U22283 (N_22283,N_21525,N_21683);
nor U22284 (N_22284,N_21994,N_21766);
xnor U22285 (N_22285,N_21846,N_21550);
xnor U22286 (N_22286,N_21738,N_21927);
nand U22287 (N_22287,N_21684,N_21709);
or U22288 (N_22288,N_21914,N_21925);
nor U22289 (N_22289,N_21587,N_21698);
or U22290 (N_22290,N_21928,N_21733);
or U22291 (N_22291,N_21958,N_21876);
nor U22292 (N_22292,N_21658,N_21716);
and U22293 (N_22293,N_21760,N_21647);
or U22294 (N_22294,N_21836,N_21856);
nand U22295 (N_22295,N_21847,N_21784);
and U22296 (N_22296,N_21544,N_21700);
and U22297 (N_22297,N_21502,N_21863);
or U22298 (N_22298,N_21589,N_21700);
xnor U22299 (N_22299,N_21508,N_21827);
nand U22300 (N_22300,N_21527,N_21895);
xor U22301 (N_22301,N_21705,N_21877);
nand U22302 (N_22302,N_21739,N_21913);
xnor U22303 (N_22303,N_21505,N_21986);
nor U22304 (N_22304,N_21750,N_21877);
or U22305 (N_22305,N_21956,N_21999);
and U22306 (N_22306,N_21845,N_21849);
xor U22307 (N_22307,N_21904,N_21673);
xor U22308 (N_22308,N_21635,N_21992);
xnor U22309 (N_22309,N_21925,N_21905);
nor U22310 (N_22310,N_21581,N_21949);
or U22311 (N_22311,N_21514,N_21795);
nor U22312 (N_22312,N_21598,N_21701);
nand U22313 (N_22313,N_21870,N_21800);
or U22314 (N_22314,N_21888,N_21908);
nand U22315 (N_22315,N_21903,N_21672);
or U22316 (N_22316,N_21985,N_21548);
xor U22317 (N_22317,N_21683,N_21687);
nand U22318 (N_22318,N_21654,N_21521);
nand U22319 (N_22319,N_21877,N_21800);
and U22320 (N_22320,N_21808,N_21926);
xnor U22321 (N_22321,N_21787,N_21690);
and U22322 (N_22322,N_21949,N_21676);
nand U22323 (N_22323,N_21741,N_21967);
nor U22324 (N_22324,N_21816,N_21808);
nand U22325 (N_22325,N_21731,N_21928);
and U22326 (N_22326,N_21530,N_21556);
nand U22327 (N_22327,N_21510,N_21574);
xnor U22328 (N_22328,N_21960,N_21911);
or U22329 (N_22329,N_21993,N_21663);
or U22330 (N_22330,N_21646,N_21832);
and U22331 (N_22331,N_21755,N_21748);
nor U22332 (N_22332,N_21946,N_21672);
nand U22333 (N_22333,N_21739,N_21598);
xnor U22334 (N_22334,N_21670,N_21600);
and U22335 (N_22335,N_21914,N_21978);
nor U22336 (N_22336,N_21916,N_21944);
nand U22337 (N_22337,N_21688,N_21926);
xor U22338 (N_22338,N_21603,N_21632);
or U22339 (N_22339,N_21938,N_21592);
xnor U22340 (N_22340,N_21825,N_21655);
and U22341 (N_22341,N_21950,N_21883);
and U22342 (N_22342,N_21695,N_21955);
nor U22343 (N_22343,N_21929,N_21562);
or U22344 (N_22344,N_21502,N_21902);
nand U22345 (N_22345,N_21846,N_21679);
and U22346 (N_22346,N_21612,N_21968);
nand U22347 (N_22347,N_21737,N_21748);
and U22348 (N_22348,N_21983,N_21906);
nand U22349 (N_22349,N_21944,N_21780);
nor U22350 (N_22350,N_21954,N_21569);
or U22351 (N_22351,N_21828,N_21838);
nand U22352 (N_22352,N_21861,N_21740);
nand U22353 (N_22353,N_21572,N_21885);
nor U22354 (N_22354,N_21728,N_21647);
and U22355 (N_22355,N_21896,N_21698);
nor U22356 (N_22356,N_21561,N_21836);
and U22357 (N_22357,N_21534,N_21602);
nand U22358 (N_22358,N_21964,N_21782);
nor U22359 (N_22359,N_21669,N_21539);
xor U22360 (N_22360,N_21951,N_21521);
or U22361 (N_22361,N_21600,N_21529);
nand U22362 (N_22362,N_21708,N_21606);
or U22363 (N_22363,N_21704,N_21844);
nor U22364 (N_22364,N_21680,N_21804);
nor U22365 (N_22365,N_21850,N_21815);
or U22366 (N_22366,N_21625,N_21989);
nand U22367 (N_22367,N_21921,N_21639);
xor U22368 (N_22368,N_21688,N_21778);
or U22369 (N_22369,N_21544,N_21731);
nand U22370 (N_22370,N_21881,N_21525);
and U22371 (N_22371,N_21901,N_21803);
and U22372 (N_22372,N_21949,N_21941);
nand U22373 (N_22373,N_21798,N_21541);
and U22374 (N_22374,N_21767,N_21745);
or U22375 (N_22375,N_21633,N_21602);
nand U22376 (N_22376,N_21713,N_21783);
or U22377 (N_22377,N_21742,N_21771);
or U22378 (N_22378,N_21627,N_21879);
nand U22379 (N_22379,N_21596,N_21988);
nor U22380 (N_22380,N_21603,N_21586);
nand U22381 (N_22381,N_21886,N_21515);
nor U22382 (N_22382,N_21818,N_21724);
or U22383 (N_22383,N_21505,N_21842);
xor U22384 (N_22384,N_21982,N_21954);
and U22385 (N_22385,N_21818,N_21563);
nor U22386 (N_22386,N_21562,N_21534);
nor U22387 (N_22387,N_21618,N_21529);
xor U22388 (N_22388,N_21658,N_21893);
and U22389 (N_22389,N_21730,N_21626);
nor U22390 (N_22390,N_21837,N_21782);
nor U22391 (N_22391,N_21928,N_21792);
or U22392 (N_22392,N_21765,N_21589);
xnor U22393 (N_22393,N_21792,N_21791);
and U22394 (N_22394,N_21944,N_21532);
or U22395 (N_22395,N_21537,N_21771);
or U22396 (N_22396,N_21518,N_21555);
or U22397 (N_22397,N_21646,N_21876);
and U22398 (N_22398,N_21922,N_21923);
or U22399 (N_22399,N_21872,N_21706);
or U22400 (N_22400,N_21673,N_21540);
xor U22401 (N_22401,N_21663,N_21756);
xnor U22402 (N_22402,N_21962,N_21805);
nand U22403 (N_22403,N_21515,N_21652);
or U22404 (N_22404,N_21697,N_21965);
xor U22405 (N_22405,N_21691,N_21969);
nor U22406 (N_22406,N_21923,N_21563);
or U22407 (N_22407,N_21757,N_21992);
xor U22408 (N_22408,N_21629,N_21916);
nor U22409 (N_22409,N_21686,N_21803);
nor U22410 (N_22410,N_21952,N_21795);
xnor U22411 (N_22411,N_21542,N_21555);
nor U22412 (N_22412,N_21843,N_21934);
nor U22413 (N_22413,N_21957,N_21582);
xnor U22414 (N_22414,N_21863,N_21790);
nand U22415 (N_22415,N_21663,N_21556);
or U22416 (N_22416,N_21845,N_21936);
or U22417 (N_22417,N_21992,N_21535);
and U22418 (N_22418,N_21760,N_21808);
xnor U22419 (N_22419,N_21736,N_21605);
and U22420 (N_22420,N_21896,N_21629);
xnor U22421 (N_22421,N_21839,N_21538);
or U22422 (N_22422,N_21919,N_21570);
and U22423 (N_22423,N_21924,N_21931);
and U22424 (N_22424,N_21847,N_21874);
nor U22425 (N_22425,N_21683,N_21551);
or U22426 (N_22426,N_21550,N_21807);
or U22427 (N_22427,N_21712,N_21667);
xor U22428 (N_22428,N_21727,N_21759);
xnor U22429 (N_22429,N_21933,N_21508);
nand U22430 (N_22430,N_21516,N_21563);
and U22431 (N_22431,N_21997,N_21881);
nor U22432 (N_22432,N_21505,N_21973);
nand U22433 (N_22433,N_21625,N_21788);
nand U22434 (N_22434,N_21920,N_21916);
nor U22435 (N_22435,N_21910,N_21953);
nor U22436 (N_22436,N_21602,N_21860);
and U22437 (N_22437,N_21911,N_21673);
nand U22438 (N_22438,N_21736,N_21849);
nand U22439 (N_22439,N_21813,N_21806);
or U22440 (N_22440,N_21849,N_21920);
nand U22441 (N_22441,N_21860,N_21705);
and U22442 (N_22442,N_21885,N_21643);
xnor U22443 (N_22443,N_21927,N_21605);
and U22444 (N_22444,N_21967,N_21765);
nor U22445 (N_22445,N_21936,N_21649);
and U22446 (N_22446,N_21968,N_21999);
nand U22447 (N_22447,N_21605,N_21785);
nor U22448 (N_22448,N_21684,N_21575);
nor U22449 (N_22449,N_21688,N_21843);
xor U22450 (N_22450,N_21661,N_21586);
nand U22451 (N_22451,N_21796,N_21961);
nor U22452 (N_22452,N_21895,N_21755);
xnor U22453 (N_22453,N_21860,N_21881);
and U22454 (N_22454,N_21502,N_21528);
nand U22455 (N_22455,N_21682,N_21771);
nor U22456 (N_22456,N_21845,N_21590);
or U22457 (N_22457,N_21657,N_21665);
nor U22458 (N_22458,N_21781,N_21690);
nor U22459 (N_22459,N_21577,N_21532);
nor U22460 (N_22460,N_21973,N_21643);
or U22461 (N_22461,N_21917,N_21615);
and U22462 (N_22462,N_21979,N_21533);
or U22463 (N_22463,N_21971,N_21736);
or U22464 (N_22464,N_21887,N_21538);
or U22465 (N_22465,N_21680,N_21792);
nand U22466 (N_22466,N_21815,N_21994);
or U22467 (N_22467,N_21810,N_21881);
or U22468 (N_22468,N_21951,N_21767);
nor U22469 (N_22469,N_21518,N_21880);
xnor U22470 (N_22470,N_21941,N_21743);
or U22471 (N_22471,N_21557,N_21835);
xor U22472 (N_22472,N_21938,N_21733);
or U22473 (N_22473,N_21565,N_21926);
and U22474 (N_22474,N_21764,N_21750);
or U22475 (N_22475,N_21711,N_21953);
or U22476 (N_22476,N_21963,N_21590);
nand U22477 (N_22477,N_21706,N_21954);
xnor U22478 (N_22478,N_21703,N_21715);
nor U22479 (N_22479,N_21674,N_21845);
xor U22480 (N_22480,N_21917,N_21724);
nor U22481 (N_22481,N_21829,N_21678);
xnor U22482 (N_22482,N_21853,N_21974);
and U22483 (N_22483,N_21628,N_21695);
nor U22484 (N_22484,N_21686,N_21772);
xnor U22485 (N_22485,N_21823,N_21569);
or U22486 (N_22486,N_21927,N_21884);
nand U22487 (N_22487,N_21571,N_21797);
or U22488 (N_22488,N_21657,N_21693);
xnor U22489 (N_22489,N_21764,N_21691);
nand U22490 (N_22490,N_21897,N_21768);
xor U22491 (N_22491,N_21770,N_21746);
xnor U22492 (N_22492,N_21652,N_21979);
or U22493 (N_22493,N_21718,N_21590);
nor U22494 (N_22494,N_21829,N_21954);
nand U22495 (N_22495,N_21984,N_21568);
xor U22496 (N_22496,N_21525,N_21852);
nand U22497 (N_22497,N_21619,N_21970);
xor U22498 (N_22498,N_21583,N_21664);
and U22499 (N_22499,N_21563,N_21969);
xnor U22500 (N_22500,N_22173,N_22050);
nand U22501 (N_22501,N_22051,N_22264);
or U22502 (N_22502,N_22117,N_22407);
nor U22503 (N_22503,N_22289,N_22018);
nand U22504 (N_22504,N_22368,N_22203);
nand U22505 (N_22505,N_22095,N_22155);
xnor U22506 (N_22506,N_22209,N_22040);
or U22507 (N_22507,N_22333,N_22312);
and U22508 (N_22508,N_22358,N_22265);
nand U22509 (N_22509,N_22398,N_22186);
xnor U22510 (N_22510,N_22255,N_22410);
or U22511 (N_22511,N_22032,N_22100);
nor U22512 (N_22512,N_22359,N_22401);
nand U22513 (N_22513,N_22011,N_22239);
nand U22514 (N_22514,N_22268,N_22411);
or U22515 (N_22515,N_22482,N_22384);
nand U22516 (N_22516,N_22053,N_22212);
and U22517 (N_22517,N_22062,N_22092);
or U22518 (N_22518,N_22338,N_22252);
xor U22519 (N_22519,N_22184,N_22473);
nand U22520 (N_22520,N_22066,N_22034);
xnor U22521 (N_22521,N_22025,N_22116);
xnor U22522 (N_22522,N_22329,N_22048);
nand U22523 (N_22523,N_22142,N_22425);
or U22524 (N_22524,N_22306,N_22055);
or U22525 (N_22525,N_22493,N_22190);
or U22526 (N_22526,N_22456,N_22156);
or U22527 (N_22527,N_22375,N_22185);
and U22528 (N_22528,N_22376,N_22499);
xnor U22529 (N_22529,N_22158,N_22144);
nor U22530 (N_22530,N_22346,N_22123);
nor U22531 (N_22531,N_22068,N_22325);
nor U22532 (N_22532,N_22310,N_22481);
nor U22533 (N_22533,N_22253,N_22172);
nor U22534 (N_22534,N_22403,N_22487);
nand U22535 (N_22535,N_22213,N_22463);
nor U22536 (N_22536,N_22107,N_22081);
nand U22537 (N_22537,N_22134,N_22019);
nor U22538 (N_22538,N_22098,N_22337);
xnor U22539 (N_22539,N_22187,N_22220);
and U22540 (N_22540,N_22026,N_22163);
xnor U22541 (N_22541,N_22469,N_22274);
nor U22542 (N_22542,N_22417,N_22273);
xor U22543 (N_22543,N_22112,N_22448);
nor U22544 (N_22544,N_22089,N_22443);
or U22545 (N_22545,N_22096,N_22041);
nand U22546 (N_22546,N_22106,N_22351);
and U22547 (N_22547,N_22372,N_22299);
nor U22548 (N_22548,N_22397,N_22243);
and U22549 (N_22549,N_22498,N_22340);
nand U22550 (N_22550,N_22354,N_22148);
xor U22551 (N_22551,N_22444,N_22205);
and U22552 (N_22552,N_22435,N_22269);
nor U22553 (N_22553,N_22028,N_22216);
xor U22554 (N_22554,N_22222,N_22439);
nor U22555 (N_22555,N_22491,N_22168);
or U22556 (N_22556,N_22064,N_22249);
and U22557 (N_22557,N_22402,N_22073);
xor U22558 (N_22558,N_22366,N_22447);
nor U22559 (N_22559,N_22294,N_22360);
and U22560 (N_22560,N_22094,N_22462);
nand U22561 (N_22561,N_22226,N_22323);
nand U22562 (N_22562,N_22450,N_22006);
xor U22563 (N_22563,N_22334,N_22084);
xor U22564 (N_22564,N_22387,N_22159);
or U22565 (N_22565,N_22371,N_22065);
and U22566 (N_22566,N_22342,N_22474);
and U22567 (N_22567,N_22234,N_22478);
and U22568 (N_22568,N_22301,N_22309);
or U22569 (N_22569,N_22017,N_22176);
or U22570 (N_22570,N_22101,N_22374);
nand U22571 (N_22571,N_22286,N_22389);
nor U22572 (N_22572,N_22150,N_22152);
nor U22573 (N_22573,N_22361,N_22151);
nor U22574 (N_22574,N_22464,N_22395);
nand U22575 (N_22575,N_22396,N_22426);
nor U22576 (N_22576,N_22189,N_22385);
xor U22577 (N_22577,N_22131,N_22157);
nor U22578 (N_22578,N_22319,N_22208);
nand U22579 (N_22579,N_22419,N_22167);
xnor U22580 (N_22580,N_22335,N_22317);
nand U22581 (N_22581,N_22353,N_22029);
or U22582 (N_22582,N_22115,N_22221);
nand U22583 (N_22583,N_22386,N_22494);
xor U22584 (N_22584,N_22078,N_22214);
nand U22585 (N_22585,N_22316,N_22196);
xor U22586 (N_22586,N_22297,N_22293);
nor U22587 (N_22587,N_22490,N_22153);
nor U22588 (N_22588,N_22496,N_22012);
and U22589 (N_22589,N_22348,N_22180);
or U22590 (N_22590,N_22010,N_22000);
nand U22591 (N_22591,N_22341,N_22432);
or U22592 (N_22592,N_22305,N_22383);
and U22593 (N_22593,N_22031,N_22271);
and U22594 (N_22594,N_22232,N_22457);
or U22595 (N_22595,N_22015,N_22304);
nor U22596 (N_22596,N_22364,N_22278);
xor U22597 (N_22597,N_22060,N_22087);
and U22598 (N_22598,N_22380,N_22270);
nand U22599 (N_22599,N_22008,N_22223);
nand U22600 (N_22600,N_22298,N_22016);
or U22601 (N_22601,N_22489,N_22200);
nand U22602 (N_22602,N_22001,N_22113);
or U22603 (N_22603,N_22072,N_22467);
or U22604 (N_22604,N_22327,N_22245);
nor U22605 (N_22605,N_22059,N_22313);
and U22606 (N_22606,N_22356,N_22345);
and U22607 (N_22607,N_22388,N_22074);
xnor U22608 (N_22608,N_22170,N_22460);
or U22609 (N_22609,N_22229,N_22138);
xor U22610 (N_22610,N_22171,N_22174);
nand U22611 (N_22611,N_22237,N_22405);
nand U22612 (N_22612,N_22391,N_22178);
xor U22613 (N_22613,N_22246,N_22262);
nor U22614 (N_22614,N_22166,N_22350);
xor U22615 (N_22615,N_22429,N_22412);
nand U22616 (N_22616,N_22242,N_22347);
or U22617 (N_22617,N_22191,N_22169);
or U22618 (N_22618,N_22283,N_22037);
nor U22619 (N_22619,N_22303,N_22033);
or U22620 (N_22620,N_22488,N_22126);
nand U22621 (N_22621,N_22254,N_22466);
and U22622 (N_22622,N_22192,N_22077);
or U22623 (N_22623,N_22322,N_22483);
and U22624 (N_22624,N_22045,N_22408);
and U22625 (N_22625,N_22014,N_22109);
nor U22626 (N_22626,N_22206,N_22227);
and U22627 (N_22627,N_22406,N_22465);
nand U22628 (N_22628,N_22195,N_22118);
and U22629 (N_22629,N_22224,N_22328);
nor U22630 (N_22630,N_22458,N_22141);
xnor U22631 (N_22631,N_22320,N_22165);
nor U22632 (N_22632,N_22230,N_22266);
nor U22633 (N_22633,N_22287,N_22315);
nand U22634 (N_22634,N_22326,N_22217);
or U22635 (N_22635,N_22003,N_22258);
or U22636 (N_22636,N_22461,N_22132);
nor U22637 (N_22637,N_22244,N_22042);
nor U22638 (N_22638,N_22218,N_22378);
nand U22639 (N_22639,N_22193,N_22377);
nand U22640 (N_22640,N_22470,N_22370);
or U22641 (N_22641,N_22104,N_22296);
nor U22642 (N_22642,N_22440,N_22423);
xnor U22643 (N_22643,N_22211,N_22357);
nand U22644 (N_22644,N_22275,N_22183);
xnor U22645 (N_22645,N_22129,N_22046);
and U22646 (N_22646,N_22004,N_22251);
nand U22647 (N_22647,N_22256,N_22280);
nand U22648 (N_22648,N_22197,N_22056);
and U22649 (N_22649,N_22061,N_22344);
and U22650 (N_22650,N_22035,N_22071);
xnor U22651 (N_22651,N_22133,N_22424);
and U22652 (N_22652,N_22143,N_22382);
nand U22653 (N_22653,N_22154,N_22495);
nor U22654 (N_22654,N_22441,N_22076);
and U22655 (N_22655,N_22324,N_22485);
and U22656 (N_22656,N_22393,N_22261);
nor U22657 (N_22657,N_22421,N_22075);
or U22658 (N_22658,N_22302,N_22414);
nand U22659 (N_22659,N_22330,N_22121);
or U22660 (N_22660,N_22369,N_22137);
nand U22661 (N_22661,N_22453,N_22091);
nand U22662 (N_22662,N_22161,N_22009);
and U22663 (N_22663,N_22002,N_22308);
nand U22664 (N_22664,N_22128,N_22108);
and U22665 (N_22665,N_22147,N_22355);
xnor U22666 (N_22666,N_22039,N_22314);
xnor U22667 (N_22667,N_22404,N_22210);
xor U22668 (N_22668,N_22149,N_22363);
and U22669 (N_22669,N_22436,N_22367);
and U22670 (N_22670,N_22020,N_22400);
xor U22671 (N_22671,N_22177,N_22427);
nor U22672 (N_22672,N_22022,N_22069);
nor U22673 (N_22673,N_22124,N_22390);
or U22674 (N_22674,N_22130,N_22175);
nand U22675 (N_22675,N_22451,N_22428);
or U22676 (N_22676,N_22445,N_22162);
nand U22677 (N_22677,N_22311,N_22418);
and U22678 (N_22678,N_22023,N_22024);
nand U22679 (N_22679,N_22257,N_22036);
xnor U22680 (N_22680,N_22492,N_22373);
or U22681 (N_22681,N_22235,N_22468);
or U22682 (N_22682,N_22477,N_22279);
xnor U22683 (N_22683,N_22103,N_22497);
nor U22684 (N_22684,N_22083,N_22263);
nand U22685 (N_22685,N_22090,N_22431);
nor U22686 (N_22686,N_22442,N_22476);
nand U22687 (N_22687,N_22446,N_22392);
or U22688 (N_22688,N_22260,N_22136);
xor U22689 (N_22689,N_22139,N_22318);
nor U22690 (N_22690,N_22430,N_22336);
xor U22691 (N_22691,N_22365,N_22199);
nand U22692 (N_22692,N_22332,N_22452);
or U22693 (N_22693,N_22285,N_22295);
nor U22694 (N_22694,N_22343,N_22145);
xor U22695 (N_22695,N_22052,N_22250);
nor U22696 (N_22696,N_22058,N_22454);
nand U22697 (N_22697,N_22282,N_22122);
nand U22698 (N_22698,N_22160,N_22379);
and U22699 (N_22699,N_22182,N_22281);
or U22700 (N_22700,N_22321,N_22110);
and U22701 (N_22701,N_22486,N_22204);
nor U22702 (N_22702,N_22267,N_22277);
or U22703 (N_22703,N_22043,N_22479);
nor U22704 (N_22704,N_22088,N_22459);
and U22705 (N_22705,N_22284,N_22114);
or U22706 (N_22706,N_22349,N_22480);
or U22707 (N_22707,N_22238,N_22472);
nand U22708 (N_22708,N_22125,N_22415);
and U22709 (N_22709,N_22231,N_22111);
xnor U22710 (N_22710,N_22399,N_22484);
nor U22711 (N_22711,N_22416,N_22207);
and U22712 (N_22712,N_22013,N_22198);
nor U22713 (N_22713,N_22140,N_22449);
and U22714 (N_22714,N_22005,N_22027);
xnor U22715 (N_22715,N_22352,N_22063);
and U22716 (N_22716,N_22339,N_22135);
nand U22717 (N_22717,N_22086,N_22422);
or U22718 (N_22718,N_22085,N_22475);
or U22719 (N_22719,N_22079,N_22331);
nor U22720 (N_22720,N_22082,N_22433);
nor U22721 (N_22721,N_22248,N_22188);
nor U22722 (N_22722,N_22290,N_22292);
or U22723 (N_22723,N_22120,N_22164);
nand U22724 (N_22724,N_22099,N_22307);
or U22725 (N_22725,N_22225,N_22054);
and U22726 (N_22726,N_22241,N_22105);
xor U22727 (N_22727,N_22215,N_22228);
and U22728 (N_22728,N_22381,N_22394);
xor U22729 (N_22729,N_22038,N_22219);
nor U22730 (N_22730,N_22080,N_22102);
nand U22731 (N_22731,N_22067,N_22420);
and U22732 (N_22732,N_22272,N_22202);
nor U22733 (N_22733,N_22057,N_22047);
xor U22734 (N_22734,N_22093,N_22455);
or U22735 (N_22735,N_22471,N_22179);
xor U22736 (N_22736,N_22021,N_22300);
or U22737 (N_22737,N_22119,N_22181);
and U22738 (N_22738,N_22291,N_22236);
and U22739 (N_22739,N_22413,N_22049);
nand U22740 (N_22740,N_22201,N_22240);
and U22741 (N_22741,N_22030,N_22437);
and U22742 (N_22742,N_22070,N_22276);
or U22743 (N_22743,N_22146,N_22194);
nor U22744 (N_22744,N_22127,N_22233);
nand U22745 (N_22745,N_22409,N_22007);
and U22746 (N_22746,N_22259,N_22097);
or U22747 (N_22747,N_22044,N_22247);
or U22748 (N_22748,N_22438,N_22434);
xor U22749 (N_22749,N_22288,N_22362);
nor U22750 (N_22750,N_22414,N_22164);
nand U22751 (N_22751,N_22177,N_22234);
and U22752 (N_22752,N_22128,N_22177);
xnor U22753 (N_22753,N_22131,N_22103);
nor U22754 (N_22754,N_22327,N_22217);
xor U22755 (N_22755,N_22153,N_22077);
or U22756 (N_22756,N_22328,N_22222);
and U22757 (N_22757,N_22498,N_22336);
xnor U22758 (N_22758,N_22441,N_22280);
nor U22759 (N_22759,N_22046,N_22381);
and U22760 (N_22760,N_22491,N_22189);
or U22761 (N_22761,N_22426,N_22480);
nor U22762 (N_22762,N_22093,N_22210);
xor U22763 (N_22763,N_22280,N_22135);
xor U22764 (N_22764,N_22370,N_22093);
xnor U22765 (N_22765,N_22455,N_22337);
and U22766 (N_22766,N_22156,N_22071);
nor U22767 (N_22767,N_22478,N_22304);
or U22768 (N_22768,N_22064,N_22312);
nand U22769 (N_22769,N_22464,N_22103);
and U22770 (N_22770,N_22168,N_22451);
nor U22771 (N_22771,N_22499,N_22239);
and U22772 (N_22772,N_22412,N_22445);
nor U22773 (N_22773,N_22483,N_22097);
or U22774 (N_22774,N_22070,N_22057);
or U22775 (N_22775,N_22475,N_22323);
nand U22776 (N_22776,N_22032,N_22099);
or U22777 (N_22777,N_22191,N_22327);
xnor U22778 (N_22778,N_22413,N_22221);
and U22779 (N_22779,N_22452,N_22283);
or U22780 (N_22780,N_22089,N_22344);
xor U22781 (N_22781,N_22330,N_22215);
xor U22782 (N_22782,N_22111,N_22045);
and U22783 (N_22783,N_22240,N_22134);
nand U22784 (N_22784,N_22165,N_22062);
xnor U22785 (N_22785,N_22282,N_22019);
nor U22786 (N_22786,N_22286,N_22439);
nand U22787 (N_22787,N_22123,N_22334);
and U22788 (N_22788,N_22248,N_22366);
nor U22789 (N_22789,N_22286,N_22258);
and U22790 (N_22790,N_22319,N_22168);
xnor U22791 (N_22791,N_22041,N_22465);
and U22792 (N_22792,N_22114,N_22334);
xnor U22793 (N_22793,N_22339,N_22286);
or U22794 (N_22794,N_22314,N_22401);
nor U22795 (N_22795,N_22047,N_22220);
nand U22796 (N_22796,N_22142,N_22384);
or U22797 (N_22797,N_22261,N_22008);
nor U22798 (N_22798,N_22005,N_22297);
xor U22799 (N_22799,N_22067,N_22341);
nand U22800 (N_22800,N_22101,N_22118);
nor U22801 (N_22801,N_22315,N_22245);
or U22802 (N_22802,N_22209,N_22360);
or U22803 (N_22803,N_22369,N_22024);
and U22804 (N_22804,N_22238,N_22140);
or U22805 (N_22805,N_22188,N_22132);
nor U22806 (N_22806,N_22200,N_22323);
nand U22807 (N_22807,N_22035,N_22263);
xnor U22808 (N_22808,N_22433,N_22326);
nor U22809 (N_22809,N_22283,N_22410);
or U22810 (N_22810,N_22386,N_22047);
and U22811 (N_22811,N_22415,N_22013);
and U22812 (N_22812,N_22008,N_22348);
xor U22813 (N_22813,N_22355,N_22096);
and U22814 (N_22814,N_22112,N_22163);
and U22815 (N_22815,N_22311,N_22149);
nand U22816 (N_22816,N_22452,N_22001);
and U22817 (N_22817,N_22444,N_22049);
xor U22818 (N_22818,N_22029,N_22016);
nor U22819 (N_22819,N_22232,N_22194);
xnor U22820 (N_22820,N_22099,N_22080);
nor U22821 (N_22821,N_22363,N_22421);
nor U22822 (N_22822,N_22256,N_22377);
or U22823 (N_22823,N_22308,N_22153);
xor U22824 (N_22824,N_22181,N_22247);
nor U22825 (N_22825,N_22433,N_22164);
nor U22826 (N_22826,N_22044,N_22179);
and U22827 (N_22827,N_22362,N_22036);
and U22828 (N_22828,N_22028,N_22048);
and U22829 (N_22829,N_22279,N_22167);
nand U22830 (N_22830,N_22163,N_22311);
and U22831 (N_22831,N_22421,N_22298);
xor U22832 (N_22832,N_22108,N_22161);
nor U22833 (N_22833,N_22459,N_22321);
nand U22834 (N_22834,N_22070,N_22330);
nor U22835 (N_22835,N_22407,N_22414);
nor U22836 (N_22836,N_22336,N_22244);
and U22837 (N_22837,N_22281,N_22377);
xor U22838 (N_22838,N_22048,N_22461);
nor U22839 (N_22839,N_22362,N_22136);
or U22840 (N_22840,N_22182,N_22009);
and U22841 (N_22841,N_22040,N_22447);
and U22842 (N_22842,N_22031,N_22168);
and U22843 (N_22843,N_22109,N_22335);
and U22844 (N_22844,N_22029,N_22131);
xnor U22845 (N_22845,N_22237,N_22166);
and U22846 (N_22846,N_22229,N_22103);
nand U22847 (N_22847,N_22065,N_22290);
and U22848 (N_22848,N_22218,N_22486);
and U22849 (N_22849,N_22355,N_22131);
nand U22850 (N_22850,N_22219,N_22425);
and U22851 (N_22851,N_22321,N_22020);
xnor U22852 (N_22852,N_22452,N_22203);
and U22853 (N_22853,N_22472,N_22368);
or U22854 (N_22854,N_22158,N_22462);
nor U22855 (N_22855,N_22091,N_22467);
nor U22856 (N_22856,N_22348,N_22283);
and U22857 (N_22857,N_22150,N_22409);
and U22858 (N_22858,N_22313,N_22259);
xor U22859 (N_22859,N_22236,N_22199);
and U22860 (N_22860,N_22465,N_22053);
or U22861 (N_22861,N_22169,N_22372);
nor U22862 (N_22862,N_22284,N_22049);
or U22863 (N_22863,N_22146,N_22316);
nand U22864 (N_22864,N_22249,N_22479);
nor U22865 (N_22865,N_22299,N_22459);
xnor U22866 (N_22866,N_22362,N_22308);
and U22867 (N_22867,N_22238,N_22399);
and U22868 (N_22868,N_22257,N_22137);
or U22869 (N_22869,N_22172,N_22333);
nand U22870 (N_22870,N_22421,N_22121);
or U22871 (N_22871,N_22185,N_22485);
nor U22872 (N_22872,N_22172,N_22411);
and U22873 (N_22873,N_22040,N_22153);
and U22874 (N_22874,N_22096,N_22378);
or U22875 (N_22875,N_22034,N_22409);
nor U22876 (N_22876,N_22268,N_22439);
nand U22877 (N_22877,N_22124,N_22011);
and U22878 (N_22878,N_22154,N_22180);
nor U22879 (N_22879,N_22056,N_22303);
and U22880 (N_22880,N_22230,N_22104);
or U22881 (N_22881,N_22168,N_22162);
nand U22882 (N_22882,N_22143,N_22191);
nand U22883 (N_22883,N_22431,N_22408);
or U22884 (N_22884,N_22466,N_22082);
or U22885 (N_22885,N_22204,N_22268);
and U22886 (N_22886,N_22406,N_22025);
or U22887 (N_22887,N_22046,N_22094);
nand U22888 (N_22888,N_22460,N_22387);
nor U22889 (N_22889,N_22233,N_22430);
or U22890 (N_22890,N_22258,N_22221);
nor U22891 (N_22891,N_22311,N_22103);
nor U22892 (N_22892,N_22051,N_22406);
xor U22893 (N_22893,N_22066,N_22165);
nand U22894 (N_22894,N_22292,N_22081);
or U22895 (N_22895,N_22222,N_22431);
xor U22896 (N_22896,N_22373,N_22311);
or U22897 (N_22897,N_22063,N_22148);
nor U22898 (N_22898,N_22309,N_22192);
and U22899 (N_22899,N_22280,N_22392);
nand U22900 (N_22900,N_22263,N_22465);
and U22901 (N_22901,N_22205,N_22019);
nand U22902 (N_22902,N_22011,N_22041);
nand U22903 (N_22903,N_22147,N_22374);
nand U22904 (N_22904,N_22217,N_22103);
nor U22905 (N_22905,N_22074,N_22022);
or U22906 (N_22906,N_22408,N_22167);
and U22907 (N_22907,N_22169,N_22189);
xnor U22908 (N_22908,N_22082,N_22403);
xnor U22909 (N_22909,N_22229,N_22195);
xor U22910 (N_22910,N_22207,N_22295);
nor U22911 (N_22911,N_22427,N_22248);
nor U22912 (N_22912,N_22141,N_22067);
nor U22913 (N_22913,N_22445,N_22158);
nor U22914 (N_22914,N_22122,N_22026);
and U22915 (N_22915,N_22414,N_22340);
and U22916 (N_22916,N_22126,N_22490);
xor U22917 (N_22917,N_22354,N_22406);
nor U22918 (N_22918,N_22166,N_22310);
nor U22919 (N_22919,N_22355,N_22203);
and U22920 (N_22920,N_22476,N_22133);
and U22921 (N_22921,N_22300,N_22172);
and U22922 (N_22922,N_22222,N_22074);
nor U22923 (N_22923,N_22278,N_22363);
and U22924 (N_22924,N_22127,N_22391);
nor U22925 (N_22925,N_22206,N_22346);
and U22926 (N_22926,N_22028,N_22153);
nor U22927 (N_22927,N_22308,N_22256);
xnor U22928 (N_22928,N_22273,N_22296);
or U22929 (N_22929,N_22028,N_22042);
or U22930 (N_22930,N_22189,N_22382);
and U22931 (N_22931,N_22198,N_22047);
xnor U22932 (N_22932,N_22134,N_22272);
nor U22933 (N_22933,N_22009,N_22290);
or U22934 (N_22934,N_22402,N_22363);
and U22935 (N_22935,N_22404,N_22192);
and U22936 (N_22936,N_22424,N_22032);
nand U22937 (N_22937,N_22181,N_22369);
nor U22938 (N_22938,N_22418,N_22172);
or U22939 (N_22939,N_22090,N_22316);
or U22940 (N_22940,N_22382,N_22237);
or U22941 (N_22941,N_22041,N_22070);
xnor U22942 (N_22942,N_22038,N_22280);
xor U22943 (N_22943,N_22339,N_22055);
or U22944 (N_22944,N_22063,N_22463);
nand U22945 (N_22945,N_22165,N_22203);
or U22946 (N_22946,N_22037,N_22281);
and U22947 (N_22947,N_22200,N_22336);
or U22948 (N_22948,N_22494,N_22284);
nand U22949 (N_22949,N_22008,N_22189);
nor U22950 (N_22950,N_22387,N_22058);
nor U22951 (N_22951,N_22221,N_22456);
and U22952 (N_22952,N_22022,N_22400);
or U22953 (N_22953,N_22247,N_22406);
xor U22954 (N_22954,N_22062,N_22045);
xnor U22955 (N_22955,N_22323,N_22136);
or U22956 (N_22956,N_22193,N_22029);
nand U22957 (N_22957,N_22378,N_22044);
nand U22958 (N_22958,N_22380,N_22156);
or U22959 (N_22959,N_22097,N_22282);
and U22960 (N_22960,N_22327,N_22485);
and U22961 (N_22961,N_22206,N_22441);
nor U22962 (N_22962,N_22205,N_22265);
xor U22963 (N_22963,N_22476,N_22446);
nor U22964 (N_22964,N_22317,N_22285);
nand U22965 (N_22965,N_22069,N_22190);
and U22966 (N_22966,N_22336,N_22011);
or U22967 (N_22967,N_22015,N_22306);
or U22968 (N_22968,N_22425,N_22078);
xnor U22969 (N_22969,N_22164,N_22032);
and U22970 (N_22970,N_22065,N_22238);
nor U22971 (N_22971,N_22331,N_22323);
xor U22972 (N_22972,N_22402,N_22292);
nor U22973 (N_22973,N_22481,N_22362);
or U22974 (N_22974,N_22075,N_22025);
xor U22975 (N_22975,N_22319,N_22114);
nor U22976 (N_22976,N_22066,N_22495);
and U22977 (N_22977,N_22026,N_22384);
and U22978 (N_22978,N_22178,N_22129);
xor U22979 (N_22979,N_22349,N_22355);
or U22980 (N_22980,N_22010,N_22303);
and U22981 (N_22981,N_22031,N_22403);
xor U22982 (N_22982,N_22064,N_22187);
xor U22983 (N_22983,N_22295,N_22252);
nand U22984 (N_22984,N_22014,N_22470);
and U22985 (N_22985,N_22074,N_22295);
nand U22986 (N_22986,N_22268,N_22318);
nor U22987 (N_22987,N_22486,N_22460);
or U22988 (N_22988,N_22275,N_22221);
xor U22989 (N_22989,N_22086,N_22277);
xor U22990 (N_22990,N_22200,N_22095);
nor U22991 (N_22991,N_22154,N_22076);
nor U22992 (N_22992,N_22426,N_22296);
nand U22993 (N_22993,N_22337,N_22451);
nor U22994 (N_22994,N_22411,N_22263);
nor U22995 (N_22995,N_22344,N_22179);
nand U22996 (N_22996,N_22160,N_22383);
nor U22997 (N_22997,N_22464,N_22086);
xnor U22998 (N_22998,N_22494,N_22492);
and U22999 (N_22999,N_22079,N_22301);
xnor U23000 (N_23000,N_22502,N_22851);
xor U23001 (N_23001,N_22749,N_22858);
and U23002 (N_23002,N_22910,N_22946);
and U23003 (N_23003,N_22517,N_22692);
nand U23004 (N_23004,N_22846,N_22809);
nand U23005 (N_23005,N_22936,N_22700);
nand U23006 (N_23006,N_22816,N_22867);
nand U23007 (N_23007,N_22532,N_22754);
or U23008 (N_23008,N_22651,N_22630);
nor U23009 (N_23009,N_22689,N_22892);
xnor U23010 (N_23010,N_22584,N_22732);
or U23011 (N_23011,N_22801,N_22557);
or U23012 (N_23012,N_22827,N_22725);
nand U23013 (N_23013,N_22666,N_22739);
nor U23014 (N_23014,N_22769,N_22930);
nand U23015 (N_23015,N_22575,N_22586);
xor U23016 (N_23016,N_22695,N_22702);
nand U23017 (N_23017,N_22991,N_22632);
and U23018 (N_23018,N_22639,N_22648);
and U23019 (N_23019,N_22529,N_22800);
nor U23020 (N_23020,N_22992,N_22719);
nand U23021 (N_23021,N_22984,N_22789);
or U23022 (N_23022,N_22876,N_22519);
and U23023 (N_23023,N_22540,N_22574);
and U23024 (N_23024,N_22665,N_22768);
xor U23025 (N_23025,N_22803,N_22658);
and U23026 (N_23026,N_22514,N_22747);
nand U23027 (N_23027,N_22958,N_22585);
or U23028 (N_23028,N_22799,N_22677);
or U23029 (N_23029,N_22833,N_22706);
or U23030 (N_23030,N_22786,N_22905);
nand U23031 (N_23031,N_22731,N_22569);
xor U23032 (N_23032,N_22948,N_22746);
and U23033 (N_23033,N_22937,N_22782);
nor U23034 (N_23034,N_22638,N_22712);
or U23035 (N_23035,N_22815,N_22776);
nand U23036 (N_23036,N_22734,N_22811);
nand U23037 (N_23037,N_22860,N_22602);
xor U23038 (N_23038,N_22608,N_22878);
nand U23039 (N_23039,N_22850,N_22622);
xnor U23040 (N_23040,N_22952,N_22647);
xnor U23041 (N_23041,N_22837,N_22922);
xor U23042 (N_23042,N_22843,N_22976);
nand U23043 (N_23043,N_22520,N_22889);
and U23044 (N_23044,N_22883,N_22927);
xnor U23045 (N_23045,N_22556,N_22977);
xor U23046 (N_23046,N_22591,N_22761);
xnor U23047 (N_23047,N_22758,N_22756);
and U23048 (N_23048,N_22753,N_22545);
nor U23049 (N_23049,N_22999,N_22982);
nand U23050 (N_23050,N_22711,N_22573);
or U23051 (N_23051,N_22604,N_22845);
or U23052 (N_23052,N_22671,N_22821);
nand U23053 (N_23053,N_22757,N_22684);
and U23054 (N_23054,N_22953,N_22628);
nor U23055 (N_23055,N_22752,N_22765);
xor U23056 (N_23056,N_22595,N_22656);
nand U23057 (N_23057,N_22884,N_22537);
xnor U23058 (N_23058,N_22510,N_22770);
and U23059 (N_23059,N_22903,N_22567);
xor U23060 (N_23060,N_22680,N_22920);
nor U23061 (N_23061,N_22634,N_22565);
or U23062 (N_23062,N_22642,N_22544);
xor U23063 (N_23063,N_22555,N_22863);
xnor U23064 (N_23064,N_22812,N_22610);
nand U23065 (N_23065,N_22531,N_22830);
xnor U23066 (N_23066,N_22566,N_22645);
nand U23067 (N_23067,N_22576,N_22662);
xnor U23068 (N_23068,N_22716,N_22560);
xor U23069 (N_23069,N_22944,N_22871);
or U23070 (N_23070,N_22637,N_22969);
or U23071 (N_23071,N_22663,N_22998);
and U23072 (N_23072,N_22996,N_22613);
nand U23073 (N_23073,N_22553,N_22854);
nor U23074 (N_23074,N_22793,N_22543);
and U23075 (N_23075,N_22699,N_22774);
or U23076 (N_23076,N_22820,N_22694);
xnor U23077 (N_23077,N_22902,N_22947);
nand U23078 (N_23078,N_22729,N_22924);
nand U23079 (N_23079,N_22538,N_22881);
nand U23080 (N_23080,N_22641,N_22908);
nand U23081 (N_23081,N_22986,N_22940);
xor U23082 (N_23082,N_22814,N_22755);
nor U23083 (N_23083,N_22709,N_22857);
and U23084 (N_23084,N_22703,N_22743);
or U23085 (N_23085,N_22597,N_22945);
nand U23086 (N_23086,N_22650,N_22562);
nand U23087 (N_23087,N_22640,N_22988);
or U23088 (N_23088,N_22733,N_22558);
and U23089 (N_23089,N_22720,N_22693);
nand U23090 (N_23090,N_22633,N_22580);
or U23091 (N_23091,N_22631,N_22527);
and U23092 (N_23092,N_22764,N_22862);
or U23093 (N_23093,N_22649,N_22503);
and U23094 (N_23094,N_22701,N_22714);
xnor U23095 (N_23095,N_22505,N_22831);
or U23096 (N_23096,N_22890,N_22721);
xor U23097 (N_23097,N_22750,N_22823);
nand U23098 (N_23098,N_22524,N_22810);
or U23099 (N_23099,N_22523,N_22931);
xor U23100 (N_23100,N_22941,N_22978);
nor U23101 (N_23101,N_22909,N_22783);
or U23102 (N_23102,N_22873,N_22698);
nand U23103 (N_23103,N_22659,N_22906);
nor U23104 (N_23104,N_22668,N_22588);
xnor U23105 (N_23105,N_22727,N_22990);
nor U23106 (N_23106,N_22621,N_22934);
nor U23107 (N_23107,N_22723,N_22893);
or U23108 (N_23108,N_22744,N_22880);
nor U23109 (N_23109,N_22802,N_22598);
nand U23110 (N_23110,N_22707,N_22797);
nand U23111 (N_23111,N_22772,N_22773);
nor U23112 (N_23112,N_22935,N_22943);
xnor U23113 (N_23113,N_22796,N_22636);
nor U23114 (N_23114,N_22859,N_22696);
and U23115 (N_23115,N_22968,N_22738);
and U23116 (N_23116,N_22913,N_22675);
and U23117 (N_23117,N_22748,N_22518);
or U23118 (N_23118,N_22506,N_22577);
or U23119 (N_23119,N_22829,N_22644);
xnor U23120 (N_23120,N_22635,N_22819);
xor U23121 (N_23121,N_22875,N_22511);
and U23122 (N_23122,N_22563,N_22885);
xnor U23123 (N_23123,N_22886,N_22603);
and U23124 (N_23124,N_22856,N_22840);
and U23125 (N_23125,N_22550,N_22735);
or U23126 (N_23126,N_22963,N_22987);
or U23127 (N_23127,N_22643,N_22708);
nor U23128 (N_23128,N_22791,N_22687);
nor U23129 (N_23129,N_22683,N_22818);
and U23130 (N_23130,N_22981,N_22713);
and U23131 (N_23131,N_22795,N_22921);
nor U23132 (N_23132,N_22778,N_22777);
nand U23133 (N_23133,N_22691,N_22861);
or U23134 (N_23134,N_22975,N_22805);
xor U23135 (N_23135,N_22688,N_22997);
nor U23136 (N_23136,N_22836,N_22513);
or U23137 (N_23137,N_22539,N_22798);
nand U23138 (N_23138,N_22839,N_22607);
nor U23139 (N_23139,N_22781,N_22847);
xnor U23140 (N_23140,N_22521,N_22918);
xnor U23141 (N_23141,N_22616,N_22932);
and U23142 (N_23142,N_22611,N_22629);
and U23143 (N_23143,N_22919,N_22760);
or U23144 (N_23144,N_22925,N_22654);
or U23145 (N_23145,N_22877,N_22915);
xnor U23146 (N_23146,N_22955,N_22678);
nor U23147 (N_23147,N_22718,N_22504);
or U23148 (N_23148,N_22686,N_22899);
nor U23149 (N_23149,N_22985,N_22736);
or U23150 (N_23150,N_22966,N_22813);
nand U23151 (N_23151,N_22600,N_22530);
and U23152 (N_23152,N_22682,N_22594);
xor U23153 (N_23153,N_22685,N_22785);
nor U23154 (N_23154,N_22742,N_22826);
nand U23155 (N_23155,N_22561,N_22564);
and U23156 (N_23156,N_22784,N_22869);
nand U23157 (N_23157,N_22933,N_22950);
and U23158 (N_23158,N_22509,N_22835);
or U23159 (N_23159,N_22762,N_22942);
and U23160 (N_23160,N_22740,N_22620);
xor U23161 (N_23161,N_22661,N_22994);
xor U23162 (N_23162,N_22972,N_22715);
nand U23163 (N_23163,N_22842,N_22974);
nand U23164 (N_23164,N_22825,N_22817);
and U23165 (N_23165,N_22779,N_22501);
nor U23166 (N_23166,N_22737,N_22849);
nor U23167 (N_23167,N_22896,N_22792);
nand U23168 (N_23168,N_22891,N_22929);
xor U23169 (N_23169,N_22790,N_22853);
xnor U23170 (N_23170,N_22592,N_22612);
nor U23171 (N_23171,N_22967,N_22559);
xnor U23172 (N_23172,N_22938,N_22674);
or U23173 (N_23173,N_22895,N_22579);
nor U23174 (N_23174,N_22570,N_22667);
nor U23175 (N_23175,N_22522,N_22832);
nor U23176 (N_23176,N_22887,N_22788);
xor U23177 (N_23177,N_22995,N_22808);
or U23178 (N_23178,N_22549,N_22615);
or U23179 (N_23179,N_22587,N_22759);
or U23180 (N_23180,N_22690,N_22970);
nor U23181 (N_23181,N_22865,N_22672);
nand U23182 (N_23182,N_22535,N_22624);
nor U23183 (N_23183,N_22547,N_22957);
xnor U23184 (N_23184,N_22528,N_22741);
or U23185 (N_23185,N_22618,N_22824);
xor U23186 (N_23186,N_22652,N_22500);
and U23187 (N_23187,N_22828,N_22879);
xor U23188 (N_23188,N_22848,N_22572);
nor U23189 (N_23189,N_22646,N_22855);
xor U23190 (N_23190,N_22960,N_22722);
xnor U23191 (N_23191,N_22625,N_22745);
nor U23192 (N_23192,N_22923,N_22911);
nor U23193 (N_23193,N_22804,N_22894);
xnor U23194 (N_23194,N_22917,N_22979);
nor U23195 (N_23195,N_22676,N_22864);
xor U23196 (N_23196,N_22508,N_22787);
xnor U23197 (N_23197,N_22904,N_22704);
xor U23198 (N_23198,N_22627,N_22548);
xor U23199 (N_23199,N_22551,N_22578);
or U23200 (N_23200,N_22898,N_22590);
nor U23201 (N_23201,N_22897,N_22601);
xor U23202 (N_23202,N_22962,N_22679);
xnor U23203 (N_23203,N_22673,N_22949);
nor U23204 (N_23204,N_22763,N_22807);
xnor U23205 (N_23205,N_22664,N_22939);
or U23206 (N_23206,N_22730,N_22771);
and U23207 (N_23207,N_22844,N_22961);
xor U23208 (N_23208,N_22697,N_22526);
nor U23209 (N_23209,N_22605,N_22841);
xor U23210 (N_23210,N_22914,N_22900);
or U23211 (N_23211,N_22965,N_22515);
or U23212 (N_23212,N_22852,N_22838);
and U23213 (N_23213,N_22717,N_22724);
or U23214 (N_23214,N_22912,N_22866);
and U23215 (N_23215,N_22870,N_22583);
nand U23216 (N_23216,N_22928,N_22546);
nor U23217 (N_23217,N_22512,N_22582);
xor U23218 (N_23218,N_22868,N_22541);
nand U23219 (N_23219,N_22874,N_22623);
nand U23220 (N_23220,N_22907,N_22767);
nand U23221 (N_23221,N_22681,N_22626);
nor U23222 (N_23222,N_22916,N_22766);
and U23223 (N_23223,N_22926,N_22669);
xor U23224 (N_23224,N_22552,N_22589);
xor U23225 (N_23225,N_22954,N_22593);
nand U23226 (N_23226,N_22983,N_22993);
xnor U23227 (N_23227,N_22617,N_22705);
or U23228 (N_23228,N_22542,N_22534);
and U23229 (N_23229,N_22507,N_22973);
or U23230 (N_23230,N_22822,N_22599);
xor U23231 (N_23231,N_22834,N_22554);
nand U23232 (N_23232,N_22670,N_22989);
or U23233 (N_23233,N_22596,N_22606);
nor U23234 (N_23234,N_22525,N_22980);
nor U23235 (N_23235,N_22533,N_22568);
or U23236 (N_23236,N_22780,N_22882);
nand U23237 (N_23237,N_22710,N_22964);
xor U23238 (N_23238,N_22775,N_22751);
or U23239 (N_23239,N_22655,N_22956);
xnor U23240 (N_23240,N_22872,N_22794);
or U23241 (N_23241,N_22581,N_22660);
nand U23242 (N_23242,N_22516,N_22726);
nor U23243 (N_23243,N_22614,N_22971);
or U23244 (N_23244,N_22657,N_22728);
or U23245 (N_23245,N_22571,N_22901);
or U23246 (N_23246,N_22806,N_22609);
or U23247 (N_23247,N_22653,N_22619);
nand U23248 (N_23248,N_22959,N_22888);
and U23249 (N_23249,N_22536,N_22951);
or U23250 (N_23250,N_22689,N_22780);
nand U23251 (N_23251,N_22590,N_22730);
and U23252 (N_23252,N_22890,N_22935);
nor U23253 (N_23253,N_22684,N_22915);
nor U23254 (N_23254,N_22945,N_22867);
and U23255 (N_23255,N_22934,N_22807);
xor U23256 (N_23256,N_22869,N_22719);
nor U23257 (N_23257,N_22872,N_22510);
nor U23258 (N_23258,N_22781,N_22731);
nor U23259 (N_23259,N_22571,N_22664);
nor U23260 (N_23260,N_22627,N_22765);
or U23261 (N_23261,N_22845,N_22962);
xor U23262 (N_23262,N_22671,N_22679);
nand U23263 (N_23263,N_22552,N_22771);
nand U23264 (N_23264,N_22913,N_22896);
or U23265 (N_23265,N_22820,N_22510);
nor U23266 (N_23266,N_22650,N_22975);
xor U23267 (N_23267,N_22932,N_22891);
and U23268 (N_23268,N_22666,N_22574);
nand U23269 (N_23269,N_22794,N_22657);
and U23270 (N_23270,N_22953,N_22541);
nand U23271 (N_23271,N_22813,N_22706);
xnor U23272 (N_23272,N_22856,N_22791);
nand U23273 (N_23273,N_22963,N_22624);
or U23274 (N_23274,N_22639,N_22520);
nor U23275 (N_23275,N_22752,N_22944);
or U23276 (N_23276,N_22915,N_22779);
nand U23277 (N_23277,N_22983,N_22835);
or U23278 (N_23278,N_22808,N_22665);
xor U23279 (N_23279,N_22667,N_22655);
and U23280 (N_23280,N_22809,N_22569);
nand U23281 (N_23281,N_22631,N_22829);
nand U23282 (N_23282,N_22669,N_22578);
nand U23283 (N_23283,N_22763,N_22553);
and U23284 (N_23284,N_22970,N_22575);
and U23285 (N_23285,N_22670,N_22674);
nor U23286 (N_23286,N_22974,N_22694);
and U23287 (N_23287,N_22533,N_22818);
nand U23288 (N_23288,N_22799,N_22858);
and U23289 (N_23289,N_22580,N_22749);
or U23290 (N_23290,N_22715,N_22773);
xor U23291 (N_23291,N_22655,N_22628);
xnor U23292 (N_23292,N_22994,N_22691);
and U23293 (N_23293,N_22888,N_22678);
nor U23294 (N_23294,N_22525,N_22852);
and U23295 (N_23295,N_22923,N_22522);
nand U23296 (N_23296,N_22712,N_22923);
xnor U23297 (N_23297,N_22530,N_22811);
or U23298 (N_23298,N_22614,N_22524);
nand U23299 (N_23299,N_22814,N_22549);
nor U23300 (N_23300,N_22732,N_22517);
and U23301 (N_23301,N_22721,N_22807);
or U23302 (N_23302,N_22505,N_22958);
nand U23303 (N_23303,N_22583,N_22590);
nand U23304 (N_23304,N_22613,N_22516);
or U23305 (N_23305,N_22697,N_22793);
xor U23306 (N_23306,N_22711,N_22525);
nor U23307 (N_23307,N_22534,N_22862);
xor U23308 (N_23308,N_22911,N_22767);
nand U23309 (N_23309,N_22758,N_22626);
or U23310 (N_23310,N_22878,N_22665);
nand U23311 (N_23311,N_22574,N_22636);
nor U23312 (N_23312,N_22935,N_22749);
and U23313 (N_23313,N_22838,N_22510);
or U23314 (N_23314,N_22730,N_22736);
and U23315 (N_23315,N_22790,N_22814);
nand U23316 (N_23316,N_22595,N_22536);
xnor U23317 (N_23317,N_22605,N_22972);
and U23318 (N_23318,N_22777,N_22599);
and U23319 (N_23319,N_22715,N_22697);
xnor U23320 (N_23320,N_22542,N_22707);
nand U23321 (N_23321,N_22541,N_22791);
nand U23322 (N_23322,N_22511,N_22682);
or U23323 (N_23323,N_22739,N_22793);
or U23324 (N_23324,N_22853,N_22640);
nor U23325 (N_23325,N_22697,N_22632);
xnor U23326 (N_23326,N_22509,N_22727);
or U23327 (N_23327,N_22510,N_22746);
or U23328 (N_23328,N_22506,N_22962);
nand U23329 (N_23329,N_22509,N_22611);
nand U23330 (N_23330,N_22941,N_22988);
nand U23331 (N_23331,N_22866,N_22624);
or U23332 (N_23332,N_22857,N_22701);
xnor U23333 (N_23333,N_22514,N_22789);
or U23334 (N_23334,N_22848,N_22988);
xor U23335 (N_23335,N_22781,N_22928);
nor U23336 (N_23336,N_22971,N_22945);
nand U23337 (N_23337,N_22756,N_22568);
and U23338 (N_23338,N_22803,N_22662);
nand U23339 (N_23339,N_22887,N_22640);
and U23340 (N_23340,N_22734,N_22973);
nor U23341 (N_23341,N_22711,N_22543);
nor U23342 (N_23342,N_22979,N_22787);
and U23343 (N_23343,N_22583,N_22818);
or U23344 (N_23344,N_22640,N_22980);
xnor U23345 (N_23345,N_22515,N_22721);
and U23346 (N_23346,N_22790,N_22965);
xnor U23347 (N_23347,N_22819,N_22562);
nor U23348 (N_23348,N_22907,N_22757);
nor U23349 (N_23349,N_22788,N_22660);
or U23350 (N_23350,N_22648,N_22811);
nor U23351 (N_23351,N_22775,N_22913);
xor U23352 (N_23352,N_22892,N_22741);
or U23353 (N_23353,N_22692,N_22964);
xnor U23354 (N_23354,N_22807,N_22700);
and U23355 (N_23355,N_22908,N_22660);
or U23356 (N_23356,N_22620,N_22503);
and U23357 (N_23357,N_22865,N_22794);
nand U23358 (N_23358,N_22689,N_22556);
nand U23359 (N_23359,N_22713,N_22765);
or U23360 (N_23360,N_22752,N_22640);
nand U23361 (N_23361,N_22714,N_22663);
or U23362 (N_23362,N_22781,N_22803);
nor U23363 (N_23363,N_22880,N_22506);
and U23364 (N_23364,N_22861,N_22544);
and U23365 (N_23365,N_22856,N_22962);
or U23366 (N_23366,N_22547,N_22658);
xnor U23367 (N_23367,N_22941,N_22873);
and U23368 (N_23368,N_22647,N_22928);
and U23369 (N_23369,N_22746,N_22829);
or U23370 (N_23370,N_22985,N_22997);
nand U23371 (N_23371,N_22720,N_22525);
or U23372 (N_23372,N_22548,N_22950);
nand U23373 (N_23373,N_22674,N_22838);
xnor U23374 (N_23374,N_22962,N_22942);
nand U23375 (N_23375,N_22516,N_22999);
nand U23376 (N_23376,N_22895,N_22542);
xor U23377 (N_23377,N_22780,N_22865);
nor U23378 (N_23378,N_22777,N_22639);
and U23379 (N_23379,N_22913,N_22915);
and U23380 (N_23380,N_22839,N_22852);
nor U23381 (N_23381,N_22764,N_22549);
or U23382 (N_23382,N_22961,N_22589);
or U23383 (N_23383,N_22660,N_22636);
nor U23384 (N_23384,N_22902,N_22745);
nand U23385 (N_23385,N_22864,N_22956);
nand U23386 (N_23386,N_22852,N_22679);
nor U23387 (N_23387,N_22543,N_22873);
nand U23388 (N_23388,N_22562,N_22521);
nor U23389 (N_23389,N_22832,N_22689);
xnor U23390 (N_23390,N_22710,N_22682);
nand U23391 (N_23391,N_22722,N_22723);
xor U23392 (N_23392,N_22758,N_22511);
nor U23393 (N_23393,N_22633,N_22509);
or U23394 (N_23394,N_22854,N_22731);
nand U23395 (N_23395,N_22894,N_22522);
nand U23396 (N_23396,N_22687,N_22528);
or U23397 (N_23397,N_22664,N_22612);
nor U23398 (N_23398,N_22940,N_22921);
nand U23399 (N_23399,N_22801,N_22771);
nand U23400 (N_23400,N_22739,N_22787);
and U23401 (N_23401,N_22991,N_22586);
xor U23402 (N_23402,N_22805,N_22514);
xnor U23403 (N_23403,N_22693,N_22910);
and U23404 (N_23404,N_22501,N_22936);
xor U23405 (N_23405,N_22877,N_22658);
nor U23406 (N_23406,N_22778,N_22728);
nand U23407 (N_23407,N_22957,N_22795);
nor U23408 (N_23408,N_22920,N_22860);
xnor U23409 (N_23409,N_22907,N_22937);
nor U23410 (N_23410,N_22600,N_22679);
nor U23411 (N_23411,N_22649,N_22910);
and U23412 (N_23412,N_22860,N_22835);
and U23413 (N_23413,N_22863,N_22611);
or U23414 (N_23414,N_22572,N_22809);
or U23415 (N_23415,N_22532,N_22836);
xnor U23416 (N_23416,N_22582,N_22915);
or U23417 (N_23417,N_22763,N_22753);
nor U23418 (N_23418,N_22980,N_22683);
or U23419 (N_23419,N_22887,N_22659);
or U23420 (N_23420,N_22869,N_22793);
nor U23421 (N_23421,N_22690,N_22958);
xnor U23422 (N_23422,N_22706,N_22794);
nand U23423 (N_23423,N_22882,N_22719);
xnor U23424 (N_23424,N_22792,N_22812);
and U23425 (N_23425,N_22535,N_22886);
xor U23426 (N_23426,N_22669,N_22633);
or U23427 (N_23427,N_22750,N_22575);
nand U23428 (N_23428,N_22781,N_22783);
xnor U23429 (N_23429,N_22954,N_22956);
or U23430 (N_23430,N_22610,N_22738);
xnor U23431 (N_23431,N_22879,N_22544);
nand U23432 (N_23432,N_22567,N_22721);
or U23433 (N_23433,N_22607,N_22863);
and U23434 (N_23434,N_22881,N_22585);
or U23435 (N_23435,N_22573,N_22968);
nor U23436 (N_23436,N_22634,N_22843);
xnor U23437 (N_23437,N_22535,N_22934);
xnor U23438 (N_23438,N_22634,N_22601);
xor U23439 (N_23439,N_22748,N_22507);
or U23440 (N_23440,N_22746,N_22824);
nor U23441 (N_23441,N_22962,N_22719);
xor U23442 (N_23442,N_22626,N_22869);
nor U23443 (N_23443,N_22982,N_22823);
or U23444 (N_23444,N_22867,N_22649);
and U23445 (N_23445,N_22560,N_22906);
and U23446 (N_23446,N_22584,N_22677);
nor U23447 (N_23447,N_22783,N_22575);
nor U23448 (N_23448,N_22915,N_22889);
and U23449 (N_23449,N_22893,N_22677);
nand U23450 (N_23450,N_22541,N_22664);
nor U23451 (N_23451,N_22747,N_22881);
nand U23452 (N_23452,N_22884,N_22950);
nand U23453 (N_23453,N_22548,N_22678);
nor U23454 (N_23454,N_22716,N_22844);
nor U23455 (N_23455,N_22697,N_22750);
xor U23456 (N_23456,N_22644,N_22876);
or U23457 (N_23457,N_22599,N_22816);
and U23458 (N_23458,N_22593,N_22521);
or U23459 (N_23459,N_22858,N_22586);
or U23460 (N_23460,N_22984,N_22653);
or U23461 (N_23461,N_22507,N_22738);
nor U23462 (N_23462,N_22804,N_22979);
nor U23463 (N_23463,N_22787,N_22503);
xnor U23464 (N_23464,N_22648,N_22744);
or U23465 (N_23465,N_22806,N_22643);
or U23466 (N_23466,N_22527,N_22904);
nor U23467 (N_23467,N_22837,N_22817);
or U23468 (N_23468,N_22573,N_22971);
xnor U23469 (N_23469,N_22573,N_22819);
nor U23470 (N_23470,N_22684,N_22658);
and U23471 (N_23471,N_22847,N_22550);
and U23472 (N_23472,N_22831,N_22614);
and U23473 (N_23473,N_22581,N_22945);
nand U23474 (N_23474,N_22709,N_22961);
xor U23475 (N_23475,N_22650,N_22764);
and U23476 (N_23476,N_22710,N_22722);
nor U23477 (N_23477,N_22970,N_22514);
or U23478 (N_23478,N_22798,N_22654);
and U23479 (N_23479,N_22745,N_22839);
and U23480 (N_23480,N_22688,N_22643);
or U23481 (N_23481,N_22673,N_22526);
or U23482 (N_23482,N_22711,N_22932);
and U23483 (N_23483,N_22571,N_22737);
and U23484 (N_23484,N_22775,N_22976);
or U23485 (N_23485,N_22789,N_22817);
or U23486 (N_23486,N_22726,N_22524);
and U23487 (N_23487,N_22662,N_22722);
xor U23488 (N_23488,N_22871,N_22510);
nor U23489 (N_23489,N_22874,N_22841);
xnor U23490 (N_23490,N_22565,N_22898);
nand U23491 (N_23491,N_22694,N_22576);
or U23492 (N_23492,N_22675,N_22833);
xor U23493 (N_23493,N_22720,N_22904);
and U23494 (N_23494,N_22787,N_22518);
or U23495 (N_23495,N_22600,N_22950);
nor U23496 (N_23496,N_22560,N_22605);
nor U23497 (N_23497,N_22958,N_22573);
xnor U23498 (N_23498,N_22943,N_22635);
nand U23499 (N_23499,N_22736,N_22721);
xnor U23500 (N_23500,N_23329,N_23302);
nand U23501 (N_23501,N_23262,N_23250);
xnor U23502 (N_23502,N_23111,N_23089);
and U23503 (N_23503,N_23469,N_23176);
nor U23504 (N_23504,N_23411,N_23104);
nor U23505 (N_23505,N_23152,N_23075);
nor U23506 (N_23506,N_23238,N_23242);
nor U23507 (N_23507,N_23059,N_23015);
nor U23508 (N_23508,N_23119,N_23353);
or U23509 (N_23509,N_23488,N_23009);
or U23510 (N_23510,N_23168,N_23211);
nand U23511 (N_23511,N_23273,N_23379);
xor U23512 (N_23512,N_23494,N_23181);
nor U23513 (N_23513,N_23341,N_23229);
nand U23514 (N_23514,N_23456,N_23451);
xnor U23515 (N_23515,N_23463,N_23122);
nand U23516 (N_23516,N_23333,N_23481);
and U23517 (N_23517,N_23072,N_23438);
or U23518 (N_23518,N_23492,N_23251);
and U23519 (N_23519,N_23140,N_23030);
or U23520 (N_23520,N_23239,N_23345);
nand U23521 (N_23521,N_23188,N_23325);
nor U23522 (N_23522,N_23281,N_23086);
or U23523 (N_23523,N_23269,N_23385);
or U23524 (N_23524,N_23131,N_23311);
nor U23525 (N_23525,N_23163,N_23146);
xnor U23526 (N_23526,N_23169,N_23095);
xor U23527 (N_23527,N_23368,N_23297);
or U23528 (N_23528,N_23381,N_23183);
xor U23529 (N_23529,N_23083,N_23372);
nand U23530 (N_23530,N_23055,N_23355);
xor U23531 (N_23531,N_23424,N_23178);
nor U23532 (N_23532,N_23477,N_23236);
nor U23533 (N_23533,N_23174,N_23461);
nor U23534 (N_23534,N_23051,N_23419);
nand U23535 (N_23535,N_23068,N_23007);
xor U23536 (N_23536,N_23475,N_23081);
nand U23537 (N_23537,N_23416,N_23042);
xor U23538 (N_23538,N_23272,N_23234);
or U23539 (N_23539,N_23450,N_23091);
nand U23540 (N_23540,N_23227,N_23185);
or U23541 (N_23541,N_23123,N_23443);
nor U23542 (N_23542,N_23225,N_23224);
nor U23543 (N_23543,N_23237,N_23374);
nor U23544 (N_23544,N_23328,N_23433);
nand U23545 (N_23545,N_23021,N_23164);
xnor U23546 (N_23546,N_23113,N_23191);
or U23547 (N_23547,N_23196,N_23375);
nor U23548 (N_23548,N_23366,N_23447);
nor U23549 (N_23549,N_23166,N_23357);
xnor U23550 (N_23550,N_23031,N_23029);
or U23551 (N_23551,N_23097,N_23118);
nand U23552 (N_23552,N_23417,N_23263);
nor U23553 (N_23553,N_23202,N_23287);
nand U23554 (N_23554,N_23479,N_23245);
nand U23555 (N_23555,N_23305,N_23421);
and U23556 (N_23556,N_23252,N_23155);
nand U23557 (N_23557,N_23499,N_23098);
xor U23558 (N_23558,N_23173,N_23257);
or U23559 (N_23559,N_23189,N_23066);
and U23560 (N_23560,N_23117,N_23474);
nand U23561 (N_23561,N_23376,N_23332);
or U23562 (N_23562,N_23150,N_23220);
or U23563 (N_23563,N_23393,N_23033);
nand U23564 (N_23564,N_23439,N_23249);
and U23565 (N_23565,N_23156,N_23192);
xnor U23566 (N_23566,N_23077,N_23036);
xor U23567 (N_23567,N_23268,N_23344);
nand U23568 (N_23568,N_23267,N_23006);
nor U23569 (N_23569,N_23258,N_23253);
or U23570 (N_23570,N_23065,N_23274);
nor U23571 (N_23571,N_23067,N_23060);
or U23572 (N_23572,N_23321,N_23276);
nor U23573 (N_23573,N_23254,N_23338);
nand U23574 (N_23574,N_23010,N_23420);
xnor U23575 (N_23575,N_23044,N_23429);
or U23576 (N_23576,N_23145,N_23310);
and U23577 (N_23577,N_23397,N_23294);
xnor U23578 (N_23578,N_23161,N_23412);
nand U23579 (N_23579,N_23124,N_23389);
nor U23580 (N_23580,N_23125,N_23039);
nand U23581 (N_23581,N_23203,N_23478);
and U23582 (N_23582,N_23410,N_23303);
xor U23583 (N_23583,N_23206,N_23316);
nand U23584 (N_23584,N_23323,N_23394);
or U23585 (N_23585,N_23343,N_23370);
or U23586 (N_23586,N_23383,N_23486);
nand U23587 (N_23587,N_23369,N_23318);
nor U23588 (N_23588,N_23057,N_23464);
or U23589 (N_23589,N_23356,N_23354);
xnor U23590 (N_23590,N_23418,N_23043);
nor U23591 (N_23591,N_23476,N_23406);
xnor U23592 (N_23592,N_23003,N_23384);
or U23593 (N_23593,N_23437,N_23398);
nor U23594 (N_23594,N_23226,N_23008);
nor U23595 (N_23595,N_23054,N_23489);
nand U23596 (N_23596,N_23466,N_23280);
xor U23597 (N_23597,N_23304,N_23050);
xor U23598 (N_23598,N_23400,N_23497);
or U23599 (N_23599,N_23326,N_23367);
nor U23600 (N_23600,N_23134,N_23387);
nor U23601 (N_23601,N_23195,N_23243);
and U23602 (N_23602,N_23427,N_23460);
nand U23603 (N_23603,N_23442,N_23232);
nor U23604 (N_23604,N_23014,N_23446);
and U23605 (N_23605,N_23024,N_23483);
and U23606 (N_23606,N_23472,N_23365);
nor U23607 (N_23607,N_23414,N_23088);
nand U23608 (N_23608,N_23363,N_23470);
nand U23609 (N_23609,N_23053,N_23444);
xor U23610 (N_23610,N_23047,N_23284);
nor U23611 (N_23611,N_23348,N_23208);
nand U23612 (N_23612,N_23013,N_23436);
and U23613 (N_23613,N_23214,N_23396);
nor U23614 (N_23614,N_23335,N_23079);
and U23615 (N_23615,N_23435,N_23114);
xor U23616 (N_23616,N_23395,N_23207);
nor U23617 (N_23617,N_23016,N_23193);
xor U23618 (N_23618,N_23132,N_23404);
or U23619 (N_23619,N_23453,N_23158);
and U23620 (N_23620,N_23040,N_23484);
nand U23621 (N_23621,N_23440,N_23023);
nor U23622 (N_23622,N_23327,N_23340);
or U23623 (N_23623,N_23217,N_23100);
and U23624 (N_23624,N_23074,N_23209);
or U23625 (N_23625,N_23144,N_23244);
nor U23626 (N_23626,N_23289,N_23485);
nor U23627 (N_23627,N_23495,N_23336);
xor U23628 (N_23628,N_23361,N_23187);
or U23629 (N_23629,N_23465,N_23022);
or U23630 (N_23630,N_23197,N_23471);
and U23631 (N_23631,N_23141,N_23128);
nand U23632 (N_23632,N_23061,N_23286);
and U23633 (N_23633,N_23093,N_23282);
and U23634 (N_23634,N_23301,N_23292);
or U23635 (N_23635,N_23415,N_23165);
xor U23636 (N_23636,N_23459,N_23147);
nor U23637 (N_23637,N_23019,N_23261);
nor U23638 (N_23638,N_23352,N_23094);
and U23639 (N_23639,N_23482,N_23223);
nand U23640 (N_23640,N_23260,N_23020);
nor U23641 (N_23641,N_23167,N_23080);
or U23642 (N_23642,N_23215,N_23378);
nor U23643 (N_23643,N_23319,N_23112);
nand U23644 (N_23644,N_23182,N_23034);
and U23645 (N_23645,N_23409,N_23002);
or U23646 (N_23646,N_23018,N_23347);
xor U23647 (N_23647,N_23076,N_23313);
and U23648 (N_23648,N_23246,N_23351);
nor U23649 (N_23649,N_23255,N_23402);
nor U23650 (N_23650,N_23180,N_23135);
or U23651 (N_23651,N_23171,N_23290);
and U23652 (N_23652,N_23004,N_23070);
or U23653 (N_23653,N_23247,N_23270);
and U23654 (N_23654,N_23493,N_23380);
and U23655 (N_23655,N_23285,N_23058);
nor U23656 (N_23656,N_23498,N_23231);
xnor U23657 (N_23657,N_23177,N_23360);
and U23658 (N_23658,N_23048,N_23334);
nand U23659 (N_23659,N_23392,N_23186);
nor U23660 (N_23660,N_23279,N_23142);
nand U23661 (N_23661,N_23448,N_23127);
xnor U23662 (N_23662,N_23078,N_23025);
and U23663 (N_23663,N_23458,N_23371);
and U23664 (N_23664,N_23320,N_23063);
nand U23665 (N_23665,N_23350,N_23151);
nand U23666 (N_23666,N_23266,N_23377);
xnor U23667 (N_23667,N_23431,N_23342);
or U23668 (N_23668,N_23071,N_23102);
nand U23669 (N_23669,N_23306,N_23364);
or U23670 (N_23670,N_23108,N_23069);
and U23671 (N_23671,N_23434,N_23265);
and U23672 (N_23672,N_23452,N_23090);
and U23673 (N_23673,N_23064,N_23455);
or U23674 (N_23674,N_23115,N_23092);
xnor U23675 (N_23675,N_23312,N_23230);
or U23676 (N_23676,N_23299,N_23032);
and U23677 (N_23677,N_23293,N_23403);
nor U23678 (N_23678,N_23233,N_23056);
nor U23679 (N_23679,N_23116,N_23441);
xnor U23680 (N_23680,N_23307,N_23084);
and U23681 (N_23681,N_23149,N_23337);
or U23682 (N_23682,N_23045,N_23487);
xnor U23683 (N_23683,N_23259,N_23490);
xnor U23684 (N_23684,N_23153,N_23358);
nand U23685 (N_23685,N_23005,N_23201);
nand U23686 (N_23686,N_23109,N_23085);
nor U23687 (N_23687,N_23046,N_23179);
nor U23688 (N_23688,N_23359,N_23190);
nand U23689 (N_23689,N_23052,N_23216);
nor U23690 (N_23690,N_23199,N_23496);
nand U23691 (N_23691,N_23248,N_23391);
xnor U23692 (N_23692,N_23213,N_23349);
or U23693 (N_23693,N_23184,N_23283);
xor U23694 (N_23694,N_23121,N_23062);
nor U23695 (N_23695,N_23143,N_23026);
xnor U23696 (N_23696,N_23315,N_23425);
and U23697 (N_23697,N_23194,N_23480);
nor U23698 (N_23698,N_23408,N_23324);
and U23699 (N_23699,N_23096,N_23390);
nor U23700 (N_23700,N_23388,N_23126);
or U23701 (N_23701,N_23148,N_23445);
xnor U23702 (N_23702,N_23154,N_23049);
or U23703 (N_23703,N_23278,N_23218);
nand U23704 (N_23704,N_23386,N_23204);
and U23705 (N_23705,N_23277,N_23175);
and U23706 (N_23706,N_23198,N_23133);
xnor U23707 (N_23707,N_23106,N_23330);
nand U23708 (N_23708,N_23139,N_23295);
nand U23709 (N_23709,N_23073,N_23222);
and U23710 (N_23710,N_23428,N_23430);
xnor U23711 (N_23711,N_23000,N_23037);
nand U23712 (N_23712,N_23457,N_23170);
or U23713 (N_23713,N_23291,N_23138);
xnor U23714 (N_23714,N_23157,N_23240);
nand U23715 (N_23715,N_23491,N_23449);
and U23716 (N_23716,N_23035,N_23041);
xnor U23717 (N_23717,N_23017,N_23129);
nand U23718 (N_23718,N_23205,N_23331);
and U23719 (N_23719,N_23264,N_23426);
nand U23720 (N_23720,N_23467,N_23219);
nand U23721 (N_23721,N_23235,N_23382);
nor U23722 (N_23722,N_23288,N_23099);
and U23723 (N_23723,N_23454,N_23296);
nand U23724 (N_23724,N_23462,N_23362);
or U23725 (N_23725,N_23413,N_23308);
nor U23726 (N_23726,N_23107,N_23309);
or U23727 (N_23727,N_23271,N_23300);
or U23728 (N_23728,N_23012,N_23027);
xor U23729 (N_23729,N_23275,N_23346);
nor U23730 (N_23730,N_23373,N_23422);
or U23731 (N_23731,N_23314,N_23339);
nor U23732 (N_23732,N_23110,N_23082);
or U23733 (N_23733,N_23210,N_23105);
or U23734 (N_23734,N_23317,N_23298);
and U23735 (N_23735,N_23212,N_23172);
nor U23736 (N_23736,N_23407,N_23322);
nand U23737 (N_23737,N_23473,N_23256);
or U23738 (N_23738,N_23103,N_23137);
nor U23739 (N_23739,N_23136,N_23228);
nand U23740 (N_23740,N_23405,N_23401);
xor U23741 (N_23741,N_23120,N_23087);
nor U23742 (N_23742,N_23028,N_23432);
nor U23743 (N_23743,N_23001,N_23101);
or U23744 (N_23744,N_23399,N_23011);
and U23745 (N_23745,N_23160,N_23423);
or U23746 (N_23746,N_23162,N_23038);
xnor U23747 (N_23747,N_23241,N_23468);
xor U23748 (N_23748,N_23130,N_23200);
and U23749 (N_23749,N_23221,N_23159);
and U23750 (N_23750,N_23461,N_23496);
nand U23751 (N_23751,N_23091,N_23343);
nand U23752 (N_23752,N_23225,N_23022);
and U23753 (N_23753,N_23400,N_23191);
and U23754 (N_23754,N_23095,N_23313);
or U23755 (N_23755,N_23338,N_23384);
xor U23756 (N_23756,N_23458,N_23487);
nor U23757 (N_23757,N_23256,N_23101);
nor U23758 (N_23758,N_23309,N_23426);
and U23759 (N_23759,N_23128,N_23324);
nor U23760 (N_23760,N_23371,N_23245);
or U23761 (N_23761,N_23225,N_23392);
xor U23762 (N_23762,N_23019,N_23171);
or U23763 (N_23763,N_23060,N_23076);
or U23764 (N_23764,N_23245,N_23094);
xor U23765 (N_23765,N_23447,N_23208);
nor U23766 (N_23766,N_23187,N_23315);
xor U23767 (N_23767,N_23316,N_23114);
or U23768 (N_23768,N_23269,N_23165);
nand U23769 (N_23769,N_23252,N_23174);
or U23770 (N_23770,N_23278,N_23157);
or U23771 (N_23771,N_23072,N_23494);
nor U23772 (N_23772,N_23046,N_23192);
and U23773 (N_23773,N_23496,N_23249);
or U23774 (N_23774,N_23099,N_23455);
xor U23775 (N_23775,N_23398,N_23472);
or U23776 (N_23776,N_23372,N_23307);
nand U23777 (N_23777,N_23272,N_23210);
and U23778 (N_23778,N_23136,N_23270);
xor U23779 (N_23779,N_23134,N_23311);
nor U23780 (N_23780,N_23082,N_23416);
or U23781 (N_23781,N_23474,N_23009);
and U23782 (N_23782,N_23245,N_23144);
nand U23783 (N_23783,N_23118,N_23135);
nand U23784 (N_23784,N_23363,N_23138);
nor U23785 (N_23785,N_23273,N_23011);
nand U23786 (N_23786,N_23340,N_23421);
or U23787 (N_23787,N_23010,N_23057);
and U23788 (N_23788,N_23405,N_23303);
and U23789 (N_23789,N_23230,N_23471);
xor U23790 (N_23790,N_23309,N_23097);
and U23791 (N_23791,N_23188,N_23166);
nor U23792 (N_23792,N_23201,N_23318);
nand U23793 (N_23793,N_23449,N_23157);
or U23794 (N_23794,N_23246,N_23432);
nand U23795 (N_23795,N_23115,N_23302);
nor U23796 (N_23796,N_23365,N_23223);
nand U23797 (N_23797,N_23393,N_23256);
or U23798 (N_23798,N_23417,N_23005);
or U23799 (N_23799,N_23314,N_23327);
nand U23800 (N_23800,N_23327,N_23406);
and U23801 (N_23801,N_23338,N_23326);
xor U23802 (N_23802,N_23490,N_23012);
and U23803 (N_23803,N_23306,N_23079);
xor U23804 (N_23804,N_23291,N_23042);
xnor U23805 (N_23805,N_23117,N_23224);
nand U23806 (N_23806,N_23478,N_23392);
nor U23807 (N_23807,N_23029,N_23011);
nand U23808 (N_23808,N_23460,N_23282);
nor U23809 (N_23809,N_23434,N_23040);
or U23810 (N_23810,N_23118,N_23212);
nand U23811 (N_23811,N_23052,N_23368);
and U23812 (N_23812,N_23264,N_23226);
or U23813 (N_23813,N_23164,N_23410);
and U23814 (N_23814,N_23082,N_23205);
or U23815 (N_23815,N_23146,N_23370);
and U23816 (N_23816,N_23340,N_23082);
and U23817 (N_23817,N_23341,N_23162);
xor U23818 (N_23818,N_23448,N_23260);
nand U23819 (N_23819,N_23379,N_23207);
or U23820 (N_23820,N_23347,N_23300);
and U23821 (N_23821,N_23194,N_23337);
and U23822 (N_23822,N_23256,N_23203);
nand U23823 (N_23823,N_23110,N_23422);
xor U23824 (N_23824,N_23499,N_23326);
xnor U23825 (N_23825,N_23283,N_23498);
nor U23826 (N_23826,N_23374,N_23454);
or U23827 (N_23827,N_23404,N_23103);
nand U23828 (N_23828,N_23012,N_23377);
nand U23829 (N_23829,N_23328,N_23391);
nor U23830 (N_23830,N_23160,N_23422);
nor U23831 (N_23831,N_23065,N_23302);
xnor U23832 (N_23832,N_23426,N_23063);
xnor U23833 (N_23833,N_23101,N_23008);
and U23834 (N_23834,N_23350,N_23154);
nor U23835 (N_23835,N_23059,N_23238);
xnor U23836 (N_23836,N_23181,N_23208);
and U23837 (N_23837,N_23230,N_23175);
xnor U23838 (N_23838,N_23015,N_23006);
xor U23839 (N_23839,N_23120,N_23461);
nor U23840 (N_23840,N_23448,N_23415);
nor U23841 (N_23841,N_23013,N_23069);
or U23842 (N_23842,N_23351,N_23486);
or U23843 (N_23843,N_23049,N_23164);
nand U23844 (N_23844,N_23312,N_23446);
or U23845 (N_23845,N_23308,N_23378);
nand U23846 (N_23846,N_23084,N_23097);
or U23847 (N_23847,N_23053,N_23314);
and U23848 (N_23848,N_23123,N_23371);
nor U23849 (N_23849,N_23132,N_23293);
nor U23850 (N_23850,N_23467,N_23196);
or U23851 (N_23851,N_23173,N_23224);
xnor U23852 (N_23852,N_23363,N_23405);
nor U23853 (N_23853,N_23070,N_23124);
nor U23854 (N_23854,N_23223,N_23394);
nor U23855 (N_23855,N_23294,N_23020);
or U23856 (N_23856,N_23283,N_23193);
nor U23857 (N_23857,N_23401,N_23006);
xor U23858 (N_23858,N_23114,N_23083);
nand U23859 (N_23859,N_23335,N_23005);
and U23860 (N_23860,N_23407,N_23430);
and U23861 (N_23861,N_23340,N_23299);
xor U23862 (N_23862,N_23288,N_23325);
nand U23863 (N_23863,N_23129,N_23387);
and U23864 (N_23864,N_23268,N_23338);
xor U23865 (N_23865,N_23118,N_23259);
nand U23866 (N_23866,N_23437,N_23491);
and U23867 (N_23867,N_23025,N_23179);
and U23868 (N_23868,N_23404,N_23494);
xnor U23869 (N_23869,N_23168,N_23241);
and U23870 (N_23870,N_23196,N_23234);
nor U23871 (N_23871,N_23433,N_23090);
nand U23872 (N_23872,N_23379,N_23089);
xor U23873 (N_23873,N_23200,N_23185);
nor U23874 (N_23874,N_23489,N_23231);
nor U23875 (N_23875,N_23335,N_23091);
nand U23876 (N_23876,N_23185,N_23365);
xnor U23877 (N_23877,N_23039,N_23191);
and U23878 (N_23878,N_23359,N_23291);
or U23879 (N_23879,N_23181,N_23176);
nand U23880 (N_23880,N_23234,N_23376);
xor U23881 (N_23881,N_23407,N_23499);
xor U23882 (N_23882,N_23243,N_23063);
and U23883 (N_23883,N_23385,N_23185);
or U23884 (N_23884,N_23189,N_23227);
nand U23885 (N_23885,N_23490,N_23068);
or U23886 (N_23886,N_23252,N_23440);
and U23887 (N_23887,N_23416,N_23382);
or U23888 (N_23888,N_23056,N_23297);
nand U23889 (N_23889,N_23303,N_23431);
xnor U23890 (N_23890,N_23026,N_23362);
xnor U23891 (N_23891,N_23037,N_23263);
nor U23892 (N_23892,N_23025,N_23238);
or U23893 (N_23893,N_23310,N_23466);
and U23894 (N_23894,N_23422,N_23403);
nand U23895 (N_23895,N_23256,N_23098);
nor U23896 (N_23896,N_23214,N_23162);
or U23897 (N_23897,N_23190,N_23440);
nor U23898 (N_23898,N_23253,N_23343);
nand U23899 (N_23899,N_23133,N_23041);
xor U23900 (N_23900,N_23372,N_23440);
nand U23901 (N_23901,N_23206,N_23460);
nor U23902 (N_23902,N_23123,N_23135);
and U23903 (N_23903,N_23219,N_23070);
and U23904 (N_23904,N_23350,N_23357);
or U23905 (N_23905,N_23386,N_23432);
xnor U23906 (N_23906,N_23072,N_23402);
xor U23907 (N_23907,N_23242,N_23312);
xor U23908 (N_23908,N_23164,N_23334);
and U23909 (N_23909,N_23414,N_23311);
xor U23910 (N_23910,N_23400,N_23063);
nor U23911 (N_23911,N_23150,N_23402);
nand U23912 (N_23912,N_23213,N_23065);
xnor U23913 (N_23913,N_23126,N_23409);
nand U23914 (N_23914,N_23131,N_23108);
and U23915 (N_23915,N_23373,N_23268);
xnor U23916 (N_23916,N_23373,N_23128);
xnor U23917 (N_23917,N_23413,N_23045);
or U23918 (N_23918,N_23271,N_23498);
and U23919 (N_23919,N_23214,N_23366);
nor U23920 (N_23920,N_23312,N_23444);
and U23921 (N_23921,N_23276,N_23421);
xor U23922 (N_23922,N_23165,N_23135);
or U23923 (N_23923,N_23447,N_23290);
xor U23924 (N_23924,N_23486,N_23212);
or U23925 (N_23925,N_23132,N_23005);
and U23926 (N_23926,N_23297,N_23032);
and U23927 (N_23927,N_23444,N_23379);
nand U23928 (N_23928,N_23371,N_23179);
xor U23929 (N_23929,N_23227,N_23226);
and U23930 (N_23930,N_23088,N_23246);
or U23931 (N_23931,N_23096,N_23363);
nand U23932 (N_23932,N_23332,N_23446);
nor U23933 (N_23933,N_23214,N_23147);
nor U23934 (N_23934,N_23087,N_23264);
xnor U23935 (N_23935,N_23276,N_23269);
xnor U23936 (N_23936,N_23018,N_23129);
or U23937 (N_23937,N_23046,N_23160);
xor U23938 (N_23938,N_23149,N_23428);
nand U23939 (N_23939,N_23271,N_23472);
nand U23940 (N_23940,N_23021,N_23320);
or U23941 (N_23941,N_23213,N_23424);
and U23942 (N_23942,N_23376,N_23416);
xnor U23943 (N_23943,N_23310,N_23015);
nor U23944 (N_23944,N_23093,N_23385);
nand U23945 (N_23945,N_23272,N_23021);
or U23946 (N_23946,N_23145,N_23253);
or U23947 (N_23947,N_23324,N_23106);
xnor U23948 (N_23948,N_23475,N_23213);
and U23949 (N_23949,N_23037,N_23188);
nand U23950 (N_23950,N_23080,N_23401);
or U23951 (N_23951,N_23161,N_23070);
and U23952 (N_23952,N_23458,N_23102);
or U23953 (N_23953,N_23222,N_23091);
nand U23954 (N_23954,N_23358,N_23430);
nor U23955 (N_23955,N_23449,N_23308);
and U23956 (N_23956,N_23398,N_23019);
nor U23957 (N_23957,N_23327,N_23089);
or U23958 (N_23958,N_23093,N_23487);
or U23959 (N_23959,N_23094,N_23377);
nor U23960 (N_23960,N_23479,N_23364);
nand U23961 (N_23961,N_23220,N_23305);
and U23962 (N_23962,N_23453,N_23477);
and U23963 (N_23963,N_23295,N_23415);
xnor U23964 (N_23964,N_23451,N_23413);
nor U23965 (N_23965,N_23146,N_23371);
and U23966 (N_23966,N_23033,N_23259);
xor U23967 (N_23967,N_23305,N_23265);
nor U23968 (N_23968,N_23252,N_23369);
and U23969 (N_23969,N_23141,N_23175);
or U23970 (N_23970,N_23253,N_23454);
and U23971 (N_23971,N_23094,N_23016);
and U23972 (N_23972,N_23383,N_23035);
xnor U23973 (N_23973,N_23123,N_23112);
nor U23974 (N_23974,N_23278,N_23437);
xor U23975 (N_23975,N_23148,N_23206);
nor U23976 (N_23976,N_23095,N_23168);
nand U23977 (N_23977,N_23312,N_23062);
or U23978 (N_23978,N_23161,N_23198);
xor U23979 (N_23979,N_23472,N_23161);
xnor U23980 (N_23980,N_23144,N_23145);
nor U23981 (N_23981,N_23373,N_23351);
or U23982 (N_23982,N_23225,N_23461);
xnor U23983 (N_23983,N_23212,N_23287);
nand U23984 (N_23984,N_23236,N_23054);
xnor U23985 (N_23985,N_23049,N_23040);
and U23986 (N_23986,N_23026,N_23281);
and U23987 (N_23987,N_23396,N_23150);
or U23988 (N_23988,N_23088,N_23313);
or U23989 (N_23989,N_23371,N_23005);
or U23990 (N_23990,N_23019,N_23387);
nor U23991 (N_23991,N_23344,N_23131);
and U23992 (N_23992,N_23483,N_23203);
or U23993 (N_23993,N_23461,N_23289);
nor U23994 (N_23994,N_23417,N_23493);
nand U23995 (N_23995,N_23313,N_23360);
or U23996 (N_23996,N_23394,N_23321);
nand U23997 (N_23997,N_23037,N_23412);
xnor U23998 (N_23998,N_23043,N_23244);
and U23999 (N_23999,N_23241,N_23025);
nor U24000 (N_24000,N_23513,N_23500);
nor U24001 (N_24001,N_23675,N_23887);
or U24002 (N_24002,N_23599,N_23951);
and U24003 (N_24003,N_23609,N_23897);
nand U24004 (N_24004,N_23885,N_23526);
nand U24005 (N_24005,N_23909,N_23704);
and U24006 (N_24006,N_23729,N_23875);
and U24007 (N_24007,N_23976,N_23984);
and U24008 (N_24008,N_23737,N_23527);
nor U24009 (N_24009,N_23763,N_23544);
xnor U24010 (N_24010,N_23912,N_23538);
nor U24011 (N_24011,N_23691,N_23840);
or U24012 (N_24012,N_23997,N_23974);
nor U24013 (N_24013,N_23938,N_23834);
and U24014 (N_24014,N_23776,N_23548);
and U24015 (N_24015,N_23781,N_23567);
or U24016 (N_24016,N_23919,N_23750);
nor U24017 (N_24017,N_23606,N_23747);
nand U24018 (N_24018,N_23820,N_23819);
or U24019 (N_24019,N_23673,N_23658);
xnor U24020 (N_24020,N_23643,N_23844);
and U24021 (N_24021,N_23765,N_23593);
nand U24022 (N_24022,N_23577,N_23901);
nor U24023 (N_24023,N_23809,N_23816);
or U24024 (N_24024,N_23983,N_23578);
or U24025 (N_24025,N_23715,N_23724);
and U24026 (N_24026,N_23789,N_23505);
and U24027 (N_24027,N_23672,N_23775);
or U24028 (N_24028,N_23697,N_23648);
nand U24029 (N_24029,N_23972,N_23512);
nor U24030 (N_24030,N_23634,N_23839);
and U24031 (N_24031,N_23662,N_23523);
nor U24032 (N_24032,N_23549,N_23749);
xnor U24033 (N_24033,N_23867,N_23861);
and U24034 (N_24034,N_23908,N_23583);
nor U24035 (N_24035,N_23690,N_23536);
nor U24036 (N_24036,N_23946,N_23980);
and U24037 (N_24037,N_23772,N_23668);
xnor U24038 (N_24038,N_23519,N_23918);
nand U24039 (N_24039,N_23712,N_23702);
xor U24040 (N_24040,N_23812,N_23925);
and U24041 (N_24041,N_23898,N_23682);
nor U24042 (N_24042,N_23687,N_23883);
xnor U24043 (N_24043,N_23773,N_23766);
and U24044 (N_24044,N_23859,N_23735);
or U24045 (N_24045,N_23958,N_23986);
and U24046 (N_24046,N_23568,N_23657);
nand U24047 (N_24047,N_23933,N_23808);
or U24048 (N_24048,N_23771,N_23641);
nand U24049 (N_24049,N_23507,N_23692);
nand U24050 (N_24050,N_23981,N_23625);
nor U24051 (N_24051,N_23565,N_23744);
or U24052 (N_24052,N_23894,N_23823);
nor U24053 (N_24053,N_23963,N_23863);
nand U24054 (N_24054,N_23708,N_23688);
and U24055 (N_24055,N_23939,N_23754);
and U24056 (N_24056,N_23604,N_23917);
nand U24057 (N_24057,N_23922,N_23624);
and U24058 (N_24058,N_23534,N_23790);
nor U24059 (N_24059,N_23971,N_23795);
xnor U24060 (N_24060,N_23993,N_23719);
and U24061 (N_24061,N_23616,N_23597);
xnor U24062 (N_24062,N_23761,N_23752);
nand U24063 (N_24063,N_23934,N_23562);
nand U24064 (N_24064,N_23770,N_23684);
nor U24065 (N_24065,N_23764,N_23829);
and U24066 (N_24066,N_23612,N_23890);
or U24067 (N_24067,N_23502,N_23791);
or U24068 (N_24068,N_23681,N_23659);
xnor U24069 (N_24069,N_23928,N_23920);
xor U24070 (N_24070,N_23913,N_23555);
nor U24071 (N_24071,N_23835,N_23585);
xor U24072 (N_24072,N_23982,N_23547);
nand U24073 (N_24073,N_23999,N_23798);
nor U24074 (N_24074,N_23650,N_23889);
or U24075 (N_24075,N_23746,N_23996);
xor U24076 (N_24076,N_23960,N_23924);
or U24077 (N_24077,N_23845,N_23869);
and U24078 (N_24078,N_23669,N_23734);
nor U24079 (N_24079,N_23930,N_23838);
or U24080 (N_24080,N_23872,N_23871);
and U24081 (N_24081,N_23953,N_23558);
xnor U24082 (N_24082,N_23814,N_23566);
or U24083 (N_24083,N_23792,N_23560);
and U24084 (N_24084,N_23916,N_23651);
nor U24085 (N_24085,N_23556,N_23945);
xnor U24086 (N_24086,N_23642,N_23892);
and U24087 (N_24087,N_23639,N_23663);
or U24088 (N_24088,N_23646,N_23857);
or U24089 (N_24089,N_23677,N_23927);
or U24090 (N_24090,N_23714,N_23973);
nor U24091 (N_24091,N_23618,N_23743);
and U24092 (N_24092,N_23638,N_23557);
or U24093 (N_24093,N_23978,N_23709);
nand U24094 (N_24094,N_23514,N_23948);
nor U24095 (N_24095,N_23598,N_23803);
and U24096 (N_24096,N_23895,N_23801);
nand U24097 (N_24097,N_23563,N_23621);
and U24098 (N_24098,N_23738,N_23730);
or U24099 (N_24099,N_23666,N_23849);
nor U24100 (N_24100,N_23811,N_23903);
xor U24101 (N_24101,N_23852,N_23674);
xor U24102 (N_24102,N_23874,N_23652);
nand U24103 (N_24103,N_23956,N_23732);
nor U24104 (N_24104,N_23573,N_23782);
xor U24105 (N_24105,N_23998,N_23707);
xnor U24106 (N_24106,N_23914,N_23818);
and U24107 (N_24107,N_23699,N_23990);
xnor U24108 (N_24108,N_23888,N_23531);
and U24109 (N_24109,N_23586,N_23813);
or U24110 (N_24110,N_23509,N_23726);
xnor U24111 (N_24111,N_23508,N_23633);
nand U24112 (N_24112,N_23535,N_23756);
xor U24113 (N_24113,N_23537,N_23602);
or U24114 (N_24114,N_23710,N_23723);
nor U24115 (N_24115,N_23760,N_23590);
xnor U24116 (N_24116,N_23944,N_23579);
xnor U24117 (N_24117,N_23717,N_23899);
nor U24118 (N_24118,N_23979,N_23628);
nand U24119 (N_24119,N_23653,N_23637);
or U24120 (N_24120,N_23571,N_23932);
and U24121 (N_24121,N_23665,N_23745);
and U24122 (N_24122,N_23727,N_23689);
and U24123 (N_24123,N_23518,N_23722);
xnor U24124 (N_24124,N_23968,N_23843);
nor U24125 (N_24125,N_23921,N_23627);
and U24126 (N_24126,N_23521,N_23530);
nor U24127 (N_24127,N_23937,N_23631);
nand U24128 (N_24128,N_23828,N_23629);
xor U24129 (N_24129,N_23995,N_23703);
nand U24130 (N_24130,N_23831,N_23966);
xor U24131 (N_24131,N_23806,N_23854);
and U24132 (N_24132,N_23636,N_23941);
or U24133 (N_24133,N_23842,N_23611);
nand U24134 (N_24134,N_23706,N_23975);
nor U24135 (N_24135,N_23705,N_23626);
nor U24136 (N_24136,N_23929,N_23615);
nand U24137 (N_24137,N_23582,N_23696);
or U24138 (N_24138,N_23554,N_23876);
or U24139 (N_24139,N_23619,N_23753);
nor U24140 (N_24140,N_23893,N_23543);
xnor U24141 (N_24141,N_23533,N_23964);
xnor U24142 (N_24142,N_23851,N_23581);
nand U24143 (N_24143,N_23862,N_23748);
nor U24144 (N_24144,N_23552,N_23794);
or U24145 (N_24145,N_23942,N_23695);
xor U24146 (N_24146,N_23522,N_23667);
nand U24147 (N_24147,N_23825,N_23768);
and U24148 (N_24148,N_23896,N_23904);
or U24149 (N_24149,N_23529,N_23736);
or U24150 (N_24150,N_23961,N_23516);
and U24151 (N_24151,N_23757,N_23926);
nor U24152 (N_24152,N_23994,N_23532);
and U24153 (N_24153,N_23936,N_23949);
nor U24154 (N_24154,N_23676,N_23617);
nand U24155 (N_24155,N_23647,N_23731);
and U24156 (N_24156,N_23685,N_23810);
and U24157 (N_24157,N_23596,N_23864);
nor U24158 (N_24158,N_23610,N_23886);
xor U24159 (N_24159,N_23906,N_23967);
xnor U24160 (N_24160,N_23713,N_23900);
and U24161 (N_24161,N_23517,N_23866);
nand U24162 (N_24162,N_23833,N_23826);
xnor U24163 (N_24163,N_23574,N_23640);
or U24164 (N_24164,N_23796,N_23680);
or U24165 (N_24165,N_23541,N_23540);
xor U24166 (N_24166,N_23817,N_23856);
xnor U24167 (N_24167,N_23935,N_23952);
xnor U24168 (N_24168,N_23780,N_23725);
nor U24169 (N_24169,N_23614,N_23711);
nor U24170 (N_24170,N_23700,N_23807);
and U24171 (N_24171,N_23940,N_23911);
or U24172 (N_24172,N_23686,N_23588);
nor U24173 (N_24173,N_23877,N_23788);
nor U24174 (N_24174,N_23884,N_23601);
nor U24175 (N_24175,N_23720,N_23846);
and U24176 (N_24176,N_23561,N_23546);
nor U24177 (N_24177,N_23800,N_23841);
or U24178 (N_24178,N_23969,N_23860);
nand U24179 (N_24179,N_23644,N_23553);
xor U24180 (N_24180,N_23832,N_23698);
nor U24181 (N_24181,N_23520,N_23955);
nor U24182 (N_24182,N_23915,N_23799);
or U24183 (N_24183,N_23880,N_23767);
xor U24184 (N_24184,N_23539,N_23515);
xnor U24185 (N_24185,N_23836,N_23622);
nand U24186 (N_24186,N_23797,N_23716);
and U24187 (N_24187,N_23510,N_23564);
or U24188 (N_24188,N_23868,N_23551);
and U24189 (N_24189,N_23592,N_23804);
or U24190 (N_24190,N_23977,N_23589);
and U24191 (N_24191,N_23882,N_23524);
and U24192 (N_24192,N_23623,N_23858);
nand U24193 (N_24193,N_23821,N_23784);
nand U24194 (N_24194,N_23721,N_23850);
or U24195 (N_24195,N_23670,N_23907);
or U24196 (N_24196,N_23656,N_23787);
xnor U24197 (N_24197,N_23570,N_23620);
nand U24198 (N_24198,N_23959,N_23575);
nand U24199 (N_24199,N_23603,N_23793);
xnor U24200 (N_24200,N_23525,N_23718);
nor U24201 (N_24201,N_23830,N_23992);
and U24202 (N_24202,N_23545,N_23501);
nand U24203 (N_24203,N_23661,N_23950);
and U24204 (N_24204,N_23591,N_23678);
nand U24205 (N_24205,N_23910,N_23559);
or U24206 (N_24206,N_23569,N_23785);
nor U24207 (N_24207,N_23655,N_23870);
nor U24208 (N_24208,N_23891,N_23576);
xnor U24209 (N_24209,N_23740,N_23595);
and U24210 (N_24210,N_23671,N_23815);
nand U24211 (N_24211,N_23774,N_23600);
xnor U24212 (N_24212,N_23848,N_23824);
nand U24213 (N_24213,N_23822,N_23855);
or U24214 (N_24214,N_23645,N_23879);
or U24215 (N_24215,N_23550,N_23751);
nor U24216 (N_24216,N_23694,N_23905);
xnor U24217 (N_24217,N_23613,N_23632);
nor U24218 (N_24218,N_23957,N_23630);
nand U24219 (N_24219,N_23777,N_23970);
and U24220 (N_24220,N_23755,N_23881);
xnor U24221 (N_24221,N_23635,N_23528);
and U24222 (N_24222,N_23506,N_23783);
nor U24223 (N_24223,N_23802,N_23504);
and U24224 (N_24224,N_23664,N_23742);
nor U24225 (N_24225,N_23762,N_23739);
nor U24226 (N_24226,N_23679,N_23511);
and U24227 (N_24227,N_23988,N_23962);
nand U24228 (N_24228,N_23605,N_23758);
nand U24229 (N_24229,N_23608,N_23728);
and U24230 (N_24230,N_23580,N_23837);
nor U24231 (N_24231,N_23594,N_23584);
or U24232 (N_24232,N_23701,N_23693);
nor U24233 (N_24233,N_23759,N_23991);
or U24234 (N_24234,N_23683,N_23769);
nor U24235 (N_24235,N_23985,N_23954);
nand U24236 (N_24236,N_23923,N_23607);
nand U24237 (N_24237,N_23654,N_23542);
nor U24238 (N_24238,N_23649,N_23902);
or U24239 (N_24239,N_23786,N_23965);
nor U24240 (N_24240,N_23989,N_23587);
or U24241 (N_24241,N_23778,N_23931);
nand U24242 (N_24242,N_23503,N_23878);
nor U24243 (N_24243,N_23827,N_23865);
xor U24244 (N_24244,N_23779,N_23805);
nand U24245 (N_24245,N_23987,N_23943);
xor U24246 (N_24246,N_23847,N_23733);
or U24247 (N_24247,N_23873,N_23853);
and U24248 (N_24248,N_23572,N_23947);
nand U24249 (N_24249,N_23741,N_23660);
and U24250 (N_24250,N_23580,N_23912);
and U24251 (N_24251,N_23729,N_23848);
or U24252 (N_24252,N_23870,N_23669);
or U24253 (N_24253,N_23521,N_23950);
nor U24254 (N_24254,N_23913,N_23922);
nor U24255 (N_24255,N_23880,N_23846);
nand U24256 (N_24256,N_23675,N_23870);
xnor U24257 (N_24257,N_23787,N_23865);
nand U24258 (N_24258,N_23556,N_23778);
nand U24259 (N_24259,N_23759,N_23875);
xnor U24260 (N_24260,N_23618,N_23682);
and U24261 (N_24261,N_23970,N_23896);
or U24262 (N_24262,N_23903,N_23530);
nand U24263 (N_24263,N_23686,N_23967);
or U24264 (N_24264,N_23663,N_23665);
nor U24265 (N_24265,N_23928,N_23606);
and U24266 (N_24266,N_23851,N_23871);
xnor U24267 (N_24267,N_23732,N_23841);
nand U24268 (N_24268,N_23842,N_23946);
and U24269 (N_24269,N_23728,N_23586);
nor U24270 (N_24270,N_23920,N_23590);
nor U24271 (N_24271,N_23754,N_23596);
nand U24272 (N_24272,N_23959,N_23900);
nand U24273 (N_24273,N_23870,N_23695);
or U24274 (N_24274,N_23858,N_23919);
nand U24275 (N_24275,N_23661,N_23538);
and U24276 (N_24276,N_23737,N_23950);
xor U24277 (N_24277,N_23902,N_23662);
nand U24278 (N_24278,N_23630,N_23706);
or U24279 (N_24279,N_23580,N_23604);
nand U24280 (N_24280,N_23794,N_23753);
nand U24281 (N_24281,N_23920,N_23926);
nor U24282 (N_24282,N_23503,N_23735);
or U24283 (N_24283,N_23934,N_23574);
xor U24284 (N_24284,N_23585,N_23545);
and U24285 (N_24285,N_23852,N_23881);
xnor U24286 (N_24286,N_23632,N_23818);
nor U24287 (N_24287,N_23668,N_23953);
xnor U24288 (N_24288,N_23559,N_23686);
nor U24289 (N_24289,N_23847,N_23503);
or U24290 (N_24290,N_23777,N_23994);
or U24291 (N_24291,N_23826,N_23680);
xor U24292 (N_24292,N_23621,N_23630);
nand U24293 (N_24293,N_23754,N_23721);
nor U24294 (N_24294,N_23844,N_23551);
xor U24295 (N_24295,N_23951,N_23604);
and U24296 (N_24296,N_23782,N_23992);
and U24297 (N_24297,N_23832,N_23601);
and U24298 (N_24298,N_23588,N_23920);
and U24299 (N_24299,N_23856,N_23646);
nor U24300 (N_24300,N_23663,N_23574);
nor U24301 (N_24301,N_23553,N_23612);
or U24302 (N_24302,N_23769,N_23606);
and U24303 (N_24303,N_23632,N_23524);
nand U24304 (N_24304,N_23867,N_23630);
or U24305 (N_24305,N_23971,N_23608);
xor U24306 (N_24306,N_23957,N_23983);
nor U24307 (N_24307,N_23547,N_23826);
and U24308 (N_24308,N_23588,N_23974);
or U24309 (N_24309,N_23581,N_23850);
and U24310 (N_24310,N_23682,N_23851);
or U24311 (N_24311,N_23634,N_23918);
xor U24312 (N_24312,N_23501,N_23771);
or U24313 (N_24313,N_23667,N_23799);
xnor U24314 (N_24314,N_23772,N_23749);
and U24315 (N_24315,N_23781,N_23695);
and U24316 (N_24316,N_23836,N_23861);
or U24317 (N_24317,N_23537,N_23636);
or U24318 (N_24318,N_23666,N_23875);
nand U24319 (N_24319,N_23696,N_23716);
xor U24320 (N_24320,N_23724,N_23588);
nor U24321 (N_24321,N_23696,N_23810);
nand U24322 (N_24322,N_23632,N_23865);
nor U24323 (N_24323,N_23700,N_23999);
and U24324 (N_24324,N_23948,N_23877);
or U24325 (N_24325,N_23590,N_23871);
nand U24326 (N_24326,N_23545,N_23986);
nand U24327 (N_24327,N_23691,N_23757);
or U24328 (N_24328,N_23630,N_23547);
and U24329 (N_24329,N_23927,N_23703);
xnor U24330 (N_24330,N_23820,N_23738);
nor U24331 (N_24331,N_23699,N_23628);
nand U24332 (N_24332,N_23528,N_23888);
nor U24333 (N_24333,N_23685,N_23545);
nor U24334 (N_24334,N_23815,N_23778);
and U24335 (N_24335,N_23632,N_23547);
nor U24336 (N_24336,N_23635,N_23644);
nand U24337 (N_24337,N_23804,N_23790);
or U24338 (N_24338,N_23939,N_23876);
or U24339 (N_24339,N_23540,N_23530);
nor U24340 (N_24340,N_23828,N_23702);
nor U24341 (N_24341,N_23597,N_23599);
and U24342 (N_24342,N_23859,N_23920);
and U24343 (N_24343,N_23802,N_23788);
nand U24344 (N_24344,N_23534,N_23565);
nor U24345 (N_24345,N_23553,N_23512);
and U24346 (N_24346,N_23839,N_23970);
xnor U24347 (N_24347,N_23724,N_23878);
or U24348 (N_24348,N_23605,N_23721);
nor U24349 (N_24349,N_23564,N_23880);
nand U24350 (N_24350,N_23888,N_23614);
nor U24351 (N_24351,N_23981,N_23544);
xnor U24352 (N_24352,N_23735,N_23881);
and U24353 (N_24353,N_23946,N_23895);
and U24354 (N_24354,N_23913,N_23634);
nor U24355 (N_24355,N_23685,N_23869);
or U24356 (N_24356,N_23914,N_23512);
and U24357 (N_24357,N_23875,N_23789);
or U24358 (N_24358,N_23500,N_23602);
xnor U24359 (N_24359,N_23970,N_23942);
or U24360 (N_24360,N_23822,N_23549);
xnor U24361 (N_24361,N_23741,N_23707);
nor U24362 (N_24362,N_23831,N_23658);
nand U24363 (N_24363,N_23786,N_23876);
nand U24364 (N_24364,N_23534,N_23918);
xor U24365 (N_24365,N_23596,N_23523);
or U24366 (N_24366,N_23839,N_23895);
and U24367 (N_24367,N_23785,N_23659);
nor U24368 (N_24368,N_23926,N_23624);
xnor U24369 (N_24369,N_23758,N_23628);
nor U24370 (N_24370,N_23987,N_23960);
xnor U24371 (N_24371,N_23949,N_23749);
nor U24372 (N_24372,N_23576,N_23631);
or U24373 (N_24373,N_23612,N_23966);
nor U24374 (N_24374,N_23831,N_23654);
or U24375 (N_24375,N_23722,N_23590);
or U24376 (N_24376,N_23616,N_23662);
and U24377 (N_24377,N_23676,N_23723);
nand U24378 (N_24378,N_23755,N_23506);
nor U24379 (N_24379,N_23900,N_23716);
nor U24380 (N_24380,N_23743,N_23615);
nand U24381 (N_24381,N_23909,N_23910);
nor U24382 (N_24382,N_23993,N_23863);
or U24383 (N_24383,N_23803,N_23734);
or U24384 (N_24384,N_23781,N_23865);
xnor U24385 (N_24385,N_23938,N_23721);
xor U24386 (N_24386,N_23804,N_23547);
xor U24387 (N_24387,N_23995,N_23939);
nand U24388 (N_24388,N_23782,N_23946);
nor U24389 (N_24389,N_23725,N_23841);
or U24390 (N_24390,N_23975,N_23540);
nor U24391 (N_24391,N_23744,N_23710);
nor U24392 (N_24392,N_23734,N_23551);
xor U24393 (N_24393,N_23694,N_23876);
and U24394 (N_24394,N_23923,N_23697);
xnor U24395 (N_24395,N_23867,N_23577);
and U24396 (N_24396,N_23843,N_23514);
or U24397 (N_24397,N_23650,N_23971);
xor U24398 (N_24398,N_23618,N_23664);
and U24399 (N_24399,N_23503,N_23929);
nor U24400 (N_24400,N_23809,N_23529);
nor U24401 (N_24401,N_23706,N_23946);
nor U24402 (N_24402,N_23661,N_23642);
or U24403 (N_24403,N_23976,N_23894);
and U24404 (N_24404,N_23798,N_23963);
nand U24405 (N_24405,N_23503,N_23660);
and U24406 (N_24406,N_23864,N_23879);
nor U24407 (N_24407,N_23932,N_23674);
nor U24408 (N_24408,N_23976,N_23505);
nand U24409 (N_24409,N_23532,N_23616);
nand U24410 (N_24410,N_23911,N_23987);
and U24411 (N_24411,N_23833,N_23718);
or U24412 (N_24412,N_23519,N_23634);
and U24413 (N_24413,N_23967,N_23739);
xor U24414 (N_24414,N_23580,N_23907);
and U24415 (N_24415,N_23556,N_23575);
nor U24416 (N_24416,N_23599,N_23865);
and U24417 (N_24417,N_23720,N_23558);
xnor U24418 (N_24418,N_23861,N_23839);
and U24419 (N_24419,N_23879,N_23718);
nand U24420 (N_24420,N_23841,N_23525);
nand U24421 (N_24421,N_23905,N_23937);
xnor U24422 (N_24422,N_23765,N_23877);
or U24423 (N_24423,N_23844,N_23574);
nand U24424 (N_24424,N_23521,N_23701);
or U24425 (N_24425,N_23594,N_23854);
nor U24426 (N_24426,N_23727,N_23814);
or U24427 (N_24427,N_23772,N_23925);
nor U24428 (N_24428,N_23581,N_23821);
or U24429 (N_24429,N_23618,N_23701);
or U24430 (N_24430,N_23933,N_23552);
nor U24431 (N_24431,N_23693,N_23953);
nand U24432 (N_24432,N_23969,N_23918);
nor U24433 (N_24433,N_23990,N_23804);
nand U24434 (N_24434,N_23685,N_23531);
and U24435 (N_24435,N_23657,N_23728);
or U24436 (N_24436,N_23950,N_23589);
and U24437 (N_24437,N_23713,N_23533);
nor U24438 (N_24438,N_23733,N_23543);
nor U24439 (N_24439,N_23782,N_23561);
or U24440 (N_24440,N_23772,N_23752);
and U24441 (N_24441,N_23700,N_23544);
xnor U24442 (N_24442,N_23500,N_23654);
and U24443 (N_24443,N_23651,N_23942);
nand U24444 (N_24444,N_23857,N_23818);
and U24445 (N_24445,N_23641,N_23700);
nand U24446 (N_24446,N_23886,N_23699);
nor U24447 (N_24447,N_23747,N_23706);
xnor U24448 (N_24448,N_23722,N_23678);
nand U24449 (N_24449,N_23759,N_23997);
xor U24450 (N_24450,N_23795,N_23820);
or U24451 (N_24451,N_23714,N_23780);
and U24452 (N_24452,N_23737,N_23938);
nand U24453 (N_24453,N_23861,N_23873);
nor U24454 (N_24454,N_23760,N_23863);
nor U24455 (N_24455,N_23581,N_23667);
nor U24456 (N_24456,N_23766,N_23525);
xnor U24457 (N_24457,N_23812,N_23645);
or U24458 (N_24458,N_23747,N_23611);
nand U24459 (N_24459,N_23696,N_23509);
nor U24460 (N_24460,N_23736,N_23657);
or U24461 (N_24461,N_23586,N_23837);
nor U24462 (N_24462,N_23556,N_23915);
nand U24463 (N_24463,N_23989,N_23562);
xor U24464 (N_24464,N_23716,N_23586);
or U24465 (N_24465,N_23605,N_23993);
and U24466 (N_24466,N_23733,N_23857);
or U24467 (N_24467,N_23832,N_23684);
nand U24468 (N_24468,N_23978,N_23964);
xnor U24469 (N_24469,N_23629,N_23620);
or U24470 (N_24470,N_23663,N_23625);
and U24471 (N_24471,N_23798,N_23625);
nor U24472 (N_24472,N_23949,N_23976);
nor U24473 (N_24473,N_23687,N_23984);
nand U24474 (N_24474,N_23938,N_23710);
or U24475 (N_24475,N_23782,N_23930);
and U24476 (N_24476,N_23954,N_23780);
nand U24477 (N_24477,N_23663,N_23589);
xnor U24478 (N_24478,N_23914,N_23883);
xor U24479 (N_24479,N_23837,N_23895);
nand U24480 (N_24480,N_23990,N_23523);
and U24481 (N_24481,N_23874,N_23795);
nand U24482 (N_24482,N_23750,N_23735);
nand U24483 (N_24483,N_23902,N_23799);
nand U24484 (N_24484,N_23951,N_23637);
nor U24485 (N_24485,N_23806,N_23649);
or U24486 (N_24486,N_23575,N_23616);
xnor U24487 (N_24487,N_23909,N_23861);
and U24488 (N_24488,N_23734,N_23989);
nor U24489 (N_24489,N_23500,N_23707);
nand U24490 (N_24490,N_23933,N_23794);
and U24491 (N_24491,N_23967,N_23642);
nor U24492 (N_24492,N_23633,N_23542);
or U24493 (N_24493,N_23650,N_23605);
xor U24494 (N_24494,N_23501,N_23850);
or U24495 (N_24495,N_23766,N_23749);
nand U24496 (N_24496,N_23866,N_23997);
nand U24497 (N_24497,N_23881,N_23706);
or U24498 (N_24498,N_23684,N_23676);
nor U24499 (N_24499,N_23776,N_23582);
and U24500 (N_24500,N_24378,N_24050);
nand U24501 (N_24501,N_24462,N_24293);
nand U24502 (N_24502,N_24047,N_24495);
or U24503 (N_24503,N_24305,N_24239);
and U24504 (N_24504,N_24242,N_24023);
xnor U24505 (N_24505,N_24272,N_24363);
xor U24506 (N_24506,N_24318,N_24193);
nor U24507 (N_24507,N_24077,N_24081);
nand U24508 (N_24508,N_24038,N_24446);
xor U24509 (N_24509,N_24046,N_24031);
xor U24510 (N_24510,N_24048,N_24475);
and U24511 (N_24511,N_24376,N_24492);
xor U24512 (N_24512,N_24054,N_24278);
or U24513 (N_24513,N_24063,N_24306);
and U24514 (N_24514,N_24301,N_24480);
or U24515 (N_24515,N_24146,N_24033);
or U24516 (N_24516,N_24257,N_24094);
nand U24517 (N_24517,N_24066,N_24157);
xnor U24518 (N_24518,N_24120,N_24255);
nand U24519 (N_24519,N_24061,N_24247);
and U24520 (N_24520,N_24088,N_24017);
nor U24521 (N_24521,N_24147,N_24384);
nand U24522 (N_24522,N_24471,N_24307);
nand U24523 (N_24523,N_24130,N_24248);
or U24524 (N_24524,N_24134,N_24175);
nor U24525 (N_24525,N_24014,N_24434);
or U24526 (N_24526,N_24347,N_24365);
nand U24527 (N_24527,N_24435,N_24029);
or U24528 (N_24528,N_24362,N_24490);
xnor U24529 (N_24529,N_24282,N_24401);
and U24530 (N_24530,N_24470,N_24106);
nand U24531 (N_24531,N_24177,N_24056);
nand U24532 (N_24532,N_24009,N_24332);
nor U24533 (N_24533,N_24155,N_24249);
and U24534 (N_24534,N_24268,N_24374);
xor U24535 (N_24535,N_24223,N_24299);
and U24536 (N_24536,N_24141,N_24427);
and U24537 (N_24537,N_24452,N_24364);
nand U24538 (N_24538,N_24270,N_24034);
and U24539 (N_24539,N_24375,N_24349);
nor U24540 (N_24540,N_24226,N_24181);
and U24541 (N_24541,N_24327,N_24197);
nand U24542 (N_24542,N_24005,N_24458);
nor U24543 (N_24543,N_24412,N_24296);
nand U24544 (N_24544,N_24032,N_24075);
xnor U24545 (N_24545,N_24489,N_24190);
nor U24546 (N_24546,N_24208,N_24224);
nor U24547 (N_24547,N_24290,N_24086);
nor U24548 (N_24548,N_24154,N_24240);
xnor U24549 (N_24549,N_24041,N_24361);
nor U24550 (N_24550,N_24402,N_24124);
nand U24551 (N_24551,N_24222,N_24289);
xnor U24552 (N_24552,N_24300,N_24122);
xor U24553 (N_24553,N_24108,N_24386);
and U24554 (N_24554,N_24180,N_24346);
and U24555 (N_24555,N_24260,N_24131);
and U24556 (N_24556,N_24128,N_24092);
nand U24557 (N_24557,N_24304,N_24123);
xnor U24558 (N_24558,N_24498,N_24043);
nand U24559 (N_24559,N_24065,N_24214);
and U24560 (N_24560,N_24430,N_24125);
and U24561 (N_24561,N_24042,N_24174);
nor U24562 (N_24562,N_24057,N_24126);
or U24563 (N_24563,N_24303,N_24411);
and U24564 (N_24564,N_24479,N_24256);
or U24565 (N_24565,N_24269,N_24285);
and U24566 (N_24566,N_24449,N_24159);
nand U24567 (N_24567,N_24409,N_24469);
and U24568 (N_24568,N_24432,N_24276);
or U24569 (N_24569,N_24233,N_24113);
nor U24570 (N_24570,N_24463,N_24232);
and U24571 (N_24571,N_24227,N_24025);
nor U24572 (N_24572,N_24339,N_24216);
nor U24573 (N_24573,N_24399,N_24100);
nand U24574 (N_24574,N_24336,N_24145);
or U24575 (N_24575,N_24472,N_24234);
nor U24576 (N_24576,N_24439,N_24450);
and U24577 (N_24577,N_24001,N_24419);
and U24578 (N_24578,N_24442,N_24002);
and U24579 (N_24579,N_24085,N_24201);
nor U24580 (N_24580,N_24184,N_24230);
or U24581 (N_24581,N_24039,N_24425);
nand U24582 (N_24582,N_24445,N_24073);
nand U24583 (N_24583,N_24231,N_24135);
nor U24584 (N_24584,N_24312,N_24398);
xnor U24585 (N_24585,N_24018,N_24058);
nand U24586 (N_24586,N_24191,N_24444);
and U24587 (N_24587,N_24024,N_24297);
xnor U24588 (N_24588,N_24275,N_24137);
and U24589 (N_24589,N_24116,N_24497);
or U24590 (N_24590,N_24357,N_24143);
nand U24591 (N_24591,N_24096,N_24367);
or U24592 (N_24592,N_24252,N_24148);
xnor U24593 (N_24593,N_24422,N_24281);
and U24594 (N_24594,N_24350,N_24359);
nor U24595 (N_24595,N_24313,N_24263);
xnor U24596 (N_24596,N_24140,N_24053);
and U24597 (N_24597,N_24342,N_24314);
nor U24598 (N_24598,N_24486,N_24459);
and U24599 (N_24599,N_24426,N_24210);
nor U24600 (N_24600,N_24265,N_24021);
nand U24601 (N_24601,N_24483,N_24244);
nand U24602 (N_24602,N_24316,N_24460);
xor U24603 (N_24603,N_24064,N_24236);
and U24604 (N_24604,N_24105,N_24280);
and U24605 (N_24605,N_24166,N_24308);
xnor U24606 (N_24606,N_24090,N_24035);
or U24607 (N_24607,N_24245,N_24102);
nand U24608 (N_24608,N_24295,N_24217);
nand U24609 (N_24609,N_24404,N_24338);
nand U24610 (N_24610,N_24084,N_24026);
or U24611 (N_24611,N_24127,N_24218);
xnor U24612 (N_24612,N_24277,N_24182);
or U24613 (N_24613,N_24400,N_24264);
and U24614 (N_24614,N_24454,N_24443);
nand U24615 (N_24615,N_24000,N_24408);
and U24616 (N_24616,N_24324,N_24104);
nor U24617 (N_24617,N_24211,N_24200);
and U24618 (N_24618,N_24366,N_24119);
and U24619 (N_24619,N_24060,N_24170);
or U24620 (N_24620,N_24474,N_24437);
and U24621 (N_24621,N_24111,N_24165);
and U24622 (N_24622,N_24162,N_24267);
and U24623 (N_24623,N_24315,N_24246);
nor U24624 (N_24624,N_24390,N_24292);
and U24625 (N_24625,N_24284,N_24052);
nor U24626 (N_24626,N_24121,N_24317);
or U24627 (N_24627,N_24185,N_24294);
and U24628 (N_24628,N_24169,N_24468);
nand U24629 (N_24629,N_24273,N_24387);
and U24630 (N_24630,N_24251,N_24133);
or U24631 (N_24631,N_24311,N_24352);
or U24632 (N_24632,N_24388,N_24076);
or U24633 (N_24633,N_24028,N_24015);
nor U24634 (N_24634,N_24139,N_24235);
xor U24635 (N_24635,N_24302,N_24109);
or U24636 (N_24636,N_24494,N_24202);
and U24637 (N_24637,N_24206,N_24418);
and U24638 (N_24638,N_24049,N_24380);
or U24639 (N_24639,N_24288,N_24089);
and U24640 (N_24640,N_24407,N_24337);
or U24641 (N_24641,N_24079,N_24478);
nor U24642 (N_24642,N_24358,N_24012);
and U24643 (N_24643,N_24433,N_24353);
and U24644 (N_24644,N_24406,N_24168);
nand U24645 (N_24645,N_24467,N_24004);
or U24646 (N_24646,N_24331,N_24428);
nor U24647 (N_24647,N_24205,N_24457);
xnor U24648 (N_24648,N_24195,N_24391);
nor U24649 (N_24649,N_24499,N_24322);
nor U24650 (N_24650,N_24229,N_24040);
xnor U24651 (N_24651,N_24320,N_24097);
and U24652 (N_24652,N_24330,N_24072);
xnor U24653 (N_24653,N_24183,N_24485);
and U24654 (N_24654,N_24417,N_24477);
nor U24655 (N_24655,N_24321,N_24343);
nand U24656 (N_24656,N_24368,N_24036);
xor U24657 (N_24657,N_24078,N_24207);
nand U24658 (N_24658,N_24225,N_24266);
and U24659 (N_24659,N_24416,N_24186);
nor U24660 (N_24660,N_24325,N_24424);
and U24661 (N_24661,N_24261,N_24083);
and U24662 (N_24662,N_24067,N_24403);
xnor U24663 (N_24663,N_24115,N_24194);
and U24664 (N_24664,N_24383,N_24382);
nand U24665 (N_24665,N_24348,N_24488);
xnor U24666 (N_24666,N_24429,N_24431);
or U24667 (N_24667,N_24259,N_24441);
nand U24668 (N_24668,N_24112,N_24019);
nor U24669 (N_24669,N_24188,N_24377);
xor U24670 (N_24670,N_24493,N_24082);
xnor U24671 (N_24671,N_24006,N_24413);
xor U24672 (N_24672,N_24487,N_24080);
nand U24673 (N_24673,N_24360,N_24414);
nand U24674 (N_24674,N_24381,N_24496);
or U24675 (N_24675,N_24243,N_24187);
xnor U24676 (N_24676,N_24209,N_24286);
nand U24677 (N_24677,N_24152,N_24172);
and U24678 (N_24678,N_24396,N_24310);
and U24679 (N_24679,N_24215,N_24068);
nand U24680 (N_24680,N_24192,N_24448);
nand U24681 (N_24681,N_24405,N_24309);
nand U24682 (N_24682,N_24114,N_24103);
or U24683 (N_24683,N_24164,N_24371);
or U24684 (N_24684,N_24095,N_24394);
nand U24685 (N_24685,N_24334,N_24328);
and U24686 (N_24686,N_24228,N_24051);
and U24687 (N_24687,N_24101,N_24393);
nand U24688 (N_24688,N_24385,N_24451);
xnor U24689 (N_24689,N_24011,N_24022);
xnor U24690 (N_24690,N_24142,N_24287);
nand U24691 (N_24691,N_24220,N_24132);
or U24692 (N_24692,N_24389,N_24117);
or U24693 (N_24693,N_24199,N_24274);
nand U24694 (N_24694,N_24481,N_24020);
nand U24695 (N_24695,N_24074,N_24356);
nor U24696 (N_24696,N_24153,N_24007);
nand U24697 (N_24697,N_24351,N_24045);
nor U24698 (N_24698,N_24370,N_24071);
nor U24699 (N_24699,N_24455,N_24238);
xor U24700 (N_24700,N_24319,N_24250);
nor U24701 (N_24701,N_24397,N_24093);
or U24702 (N_24702,N_24464,N_24179);
or U24703 (N_24703,N_24010,N_24271);
nand U24704 (N_24704,N_24167,N_24138);
and U24705 (N_24705,N_24158,N_24379);
and U24706 (N_24706,N_24087,N_24196);
and U24707 (N_24707,N_24329,N_24283);
nor U24708 (N_24708,N_24069,N_24453);
xor U24709 (N_24709,N_24369,N_24410);
nor U24710 (N_24710,N_24258,N_24037);
nor U24711 (N_24711,N_24415,N_24161);
or U24712 (N_24712,N_24098,N_24016);
nor U24713 (N_24713,N_24456,N_24423);
nor U24714 (N_24714,N_24173,N_24003);
nor U24715 (N_24715,N_24438,N_24279);
or U24716 (N_24716,N_24340,N_24160);
or U24717 (N_24717,N_24198,N_24163);
or U24718 (N_24718,N_24345,N_24091);
or U24719 (N_24719,N_24107,N_24118);
or U24720 (N_24720,N_24136,N_24484);
or U24721 (N_24721,N_24221,N_24341);
or U24722 (N_24722,N_24062,N_24204);
nand U24723 (N_24723,N_24344,N_24070);
nand U24724 (N_24724,N_24421,N_24144);
or U24725 (N_24725,N_24213,N_24253);
and U24726 (N_24726,N_24335,N_24333);
nand U24727 (N_24727,N_24059,N_24013);
xnor U24728 (N_24728,N_24027,N_24241);
and U24729 (N_24729,N_24055,N_24373);
xnor U24730 (N_24730,N_24354,N_24473);
and U24731 (N_24731,N_24491,N_24008);
nor U24732 (N_24732,N_24420,N_24171);
or U24733 (N_24733,N_24237,N_24030);
and U24734 (N_24734,N_24150,N_24044);
and U24735 (N_24735,N_24323,N_24254);
and U24736 (N_24736,N_24291,N_24110);
xor U24737 (N_24737,N_24465,N_24466);
nand U24738 (N_24738,N_24212,N_24476);
xor U24739 (N_24739,N_24099,N_24178);
and U24740 (N_24740,N_24482,N_24189);
or U24741 (N_24741,N_24326,N_24129);
nor U24742 (N_24742,N_24395,N_24461);
or U24743 (N_24743,N_24440,N_24262);
xor U24744 (N_24744,N_24447,N_24176);
and U24745 (N_24745,N_24203,N_24151);
nor U24746 (N_24746,N_24355,N_24156);
or U24747 (N_24747,N_24298,N_24392);
or U24748 (N_24748,N_24149,N_24372);
and U24749 (N_24749,N_24436,N_24219);
nor U24750 (N_24750,N_24317,N_24001);
or U24751 (N_24751,N_24406,N_24150);
and U24752 (N_24752,N_24172,N_24263);
or U24753 (N_24753,N_24449,N_24383);
and U24754 (N_24754,N_24082,N_24358);
and U24755 (N_24755,N_24234,N_24364);
or U24756 (N_24756,N_24496,N_24368);
nand U24757 (N_24757,N_24092,N_24402);
xor U24758 (N_24758,N_24065,N_24311);
and U24759 (N_24759,N_24138,N_24233);
nor U24760 (N_24760,N_24019,N_24320);
nor U24761 (N_24761,N_24178,N_24310);
and U24762 (N_24762,N_24328,N_24083);
xor U24763 (N_24763,N_24449,N_24433);
xnor U24764 (N_24764,N_24160,N_24380);
or U24765 (N_24765,N_24352,N_24165);
nor U24766 (N_24766,N_24456,N_24310);
or U24767 (N_24767,N_24369,N_24057);
xor U24768 (N_24768,N_24167,N_24022);
and U24769 (N_24769,N_24313,N_24111);
xnor U24770 (N_24770,N_24066,N_24375);
or U24771 (N_24771,N_24337,N_24306);
nand U24772 (N_24772,N_24024,N_24232);
and U24773 (N_24773,N_24181,N_24284);
nand U24774 (N_24774,N_24449,N_24119);
or U24775 (N_24775,N_24035,N_24033);
or U24776 (N_24776,N_24251,N_24483);
and U24777 (N_24777,N_24112,N_24255);
and U24778 (N_24778,N_24433,N_24094);
nand U24779 (N_24779,N_24467,N_24114);
nand U24780 (N_24780,N_24261,N_24499);
nand U24781 (N_24781,N_24021,N_24223);
nand U24782 (N_24782,N_24440,N_24149);
nor U24783 (N_24783,N_24118,N_24000);
nand U24784 (N_24784,N_24430,N_24043);
nand U24785 (N_24785,N_24033,N_24308);
and U24786 (N_24786,N_24128,N_24086);
and U24787 (N_24787,N_24080,N_24113);
nand U24788 (N_24788,N_24258,N_24013);
and U24789 (N_24789,N_24357,N_24034);
nor U24790 (N_24790,N_24137,N_24475);
and U24791 (N_24791,N_24133,N_24276);
xnor U24792 (N_24792,N_24482,N_24179);
or U24793 (N_24793,N_24021,N_24389);
or U24794 (N_24794,N_24302,N_24245);
and U24795 (N_24795,N_24247,N_24484);
nand U24796 (N_24796,N_24095,N_24021);
nand U24797 (N_24797,N_24218,N_24173);
nand U24798 (N_24798,N_24480,N_24100);
xor U24799 (N_24799,N_24232,N_24247);
xor U24800 (N_24800,N_24107,N_24344);
or U24801 (N_24801,N_24188,N_24436);
or U24802 (N_24802,N_24199,N_24323);
nand U24803 (N_24803,N_24217,N_24086);
xnor U24804 (N_24804,N_24098,N_24014);
and U24805 (N_24805,N_24211,N_24158);
xnor U24806 (N_24806,N_24074,N_24000);
xor U24807 (N_24807,N_24186,N_24287);
or U24808 (N_24808,N_24168,N_24307);
or U24809 (N_24809,N_24110,N_24228);
and U24810 (N_24810,N_24377,N_24251);
nand U24811 (N_24811,N_24495,N_24027);
xor U24812 (N_24812,N_24195,N_24413);
and U24813 (N_24813,N_24209,N_24226);
nor U24814 (N_24814,N_24401,N_24225);
nor U24815 (N_24815,N_24184,N_24307);
nand U24816 (N_24816,N_24000,N_24292);
xnor U24817 (N_24817,N_24228,N_24077);
and U24818 (N_24818,N_24447,N_24444);
nand U24819 (N_24819,N_24221,N_24149);
nor U24820 (N_24820,N_24003,N_24147);
xnor U24821 (N_24821,N_24010,N_24496);
xor U24822 (N_24822,N_24095,N_24364);
and U24823 (N_24823,N_24427,N_24142);
or U24824 (N_24824,N_24076,N_24044);
or U24825 (N_24825,N_24268,N_24278);
xor U24826 (N_24826,N_24080,N_24463);
xor U24827 (N_24827,N_24007,N_24020);
or U24828 (N_24828,N_24244,N_24204);
nand U24829 (N_24829,N_24239,N_24140);
or U24830 (N_24830,N_24250,N_24010);
or U24831 (N_24831,N_24114,N_24191);
nand U24832 (N_24832,N_24328,N_24225);
xnor U24833 (N_24833,N_24203,N_24277);
or U24834 (N_24834,N_24399,N_24423);
or U24835 (N_24835,N_24205,N_24409);
and U24836 (N_24836,N_24263,N_24281);
nand U24837 (N_24837,N_24385,N_24329);
or U24838 (N_24838,N_24107,N_24087);
or U24839 (N_24839,N_24207,N_24417);
nor U24840 (N_24840,N_24220,N_24498);
nand U24841 (N_24841,N_24095,N_24186);
nor U24842 (N_24842,N_24416,N_24116);
xnor U24843 (N_24843,N_24445,N_24340);
nand U24844 (N_24844,N_24227,N_24422);
and U24845 (N_24845,N_24390,N_24133);
and U24846 (N_24846,N_24086,N_24402);
and U24847 (N_24847,N_24444,N_24205);
or U24848 (N_24848,N_24009,N_24063);
nor U24849 (N_24849,N_24305,N_24216);
nand U24850 (N_24850,N_24257,N_24169);
xnor U24851 (N_24851,N_24417,N_24336);
and U24852 (N_24852,N_24404,N_24208);
xnor U24853 (N_24853,N_24110,N_24310);
nor U24854 (N_24854,N_24175,N_24043);
and U24855 (N_24855,N_24250,N_24488);
xnor U24856 (N_24856,N_24109,N_24398);
or U24857 (N_24857,N_24460,N_24080);
and U24858 (N_24858,N_24053,N_24415);
nand U24859 (N_24859,N_24007,N_24279);
or U24860 (N_24860,N_24378,N_24319);
xor U24861 (N_24861,N_24335,N_24245);
xor U24862 (N_24862,N_24374,N_24286);
and U24863 (N_24863,N_24184,N_24006);
and U24864 (N_24864,N_24457,N_24263);
nor U24865 (N_24865,N_24154,N_24246);
xnor U24866 (N_24866,N_24301,N_24174);
or U24867 (N_24867,N_24359,N_24014);
nand U24868 (N_24868,N_24336,N_24300);
or U24869 (N_24869,N_24062,N_24478);
xnor U24870 (N_24870,N_24279,N_24392);
or U24871 (N_24871,N_24336,N_24354);
and U24872 (N_24872,N_24327,N_24086);
and U24873 (N_24873,N_24219,N_24357);
or U24874 (N_24874,N_24292,N_24477);
nand U24875 (N_24875,N_24451,N_24024);
and U24876 (N_24876,N_24145,N_24409);
nor U24877 (N_24877,N_24427,N_24070);
or U24878 (N_24878,N_24065,N_24455);
nand U24879 (N_24879,N_24224,N_24214);
or U24880 (N_24880,N_24488,N_24063);
or U24881 (N_24881,N_24409,N_24397);
nand U24882 (N_24882,N_24433,N_24034);
nor U24883 (N_24883,N_24167,N_24253);
and U24884 (N_24884,N_24446,N_24088);
and U24885 (N_24885,N_24442,N_24276);
and U24886 (N_24886,N_24492,N_24316);
xor U24887 (N_24887,N_24217,N_24022);
xnor U24888 (N_24888,N_24428,N_24402);
nand U24889 (N_24889,N_24043,N_24247);
nor U24890 (N_24890,N_24145,N_24129);
or U24891 (N_24891,N_24353,N_24195);
or U24892 (N_24892,N_24360,N_24346);
or U24893 (N_24893,N_24461,N_24464);
xnor U24894 (N_24894,N_24408,N_24347);
nand U24895 (N_24895,N_24269,N_24158);
or U24896 (N_24896,N_24355,N_24163);
xor U24897 (N_24897,N_24296,N_24086);
nand U24898 (N_24898,N_24418,N_24247);
xnor U24899 (N_24899,N_24343,N_24084);
xor U24900 (N_24900,N_24083,N_24286);
and U24901 (N_24901,N_24307,N_24082);
and U24902 (N_24902,N_24127,N_24068);
xnor U24903 (N_24903,N_24463,N_24013);
and U24904 (N_24904,N_24129,N_24195);
nand U24905 (N_24905,N_24098,N_24089);
nand U24906 (N_24906,N_24070,N_24000);
nand U24907 (N_24907,N_24191,N_24203);
nor U24908 (N_24908,N_24210,N_24235);
or U24909 (N_24909,N_24405,N_24473);
or U24910 (N_24910,N_24374,N_24391);
or U24911 (N_24911,N_24459,N_24376);
nor U24912 (N_24912,N_24098,N_24237);
or U24913 (N_24913,N_24302,N_24358);
nor U24914 (N_24914,N_24225,N_24195);
and U24915 (N_24915,N_24087,N_24321);
or U24916 (N_24916,N_24284,N_24359);
nor U24917 (N_24917,N_24237,N_24191);
nor U24918 (N_24918,N_24037,N_24460);
nand U24919 (N_24919,N_24244,N_24288);
nand U24920 (N_24920,N_24324,N_24436);
xnor U24921 (N_24921,N_24253,N_24103);
xnor U24922 (N_24922,N_24200,N_24497);
or U24923 (N_24923,N_24422,N_24248);
xor U24924 (N_24924,N_24464,N_24214);
nand U24925 (N_24925,N_24197,N_24168);
xnor U24926 (N_24926,N_24216,N_24079);
or U24927 (N_24927,N_24411,N_24271);
xor U24928 (N_24928,N_24340,N_24123);
xor U24929 (N_24929,N_24336,N_24127);
nand U24930 (N_24930,N_24129,N_24028);
or U24931 (N_24931,N_24495,N_24479);
and U24932 (N_24932,N_24385,N_24169);
nor U24933 (N_24933,N_24092,N_24439);
nand U24934 (N_24934,N_24060,N_24422);
nor U24935 (N_24935,N_24477,N_24381);
xor U24936 (N_24936,N_24270,N_24118);
nand U24937 (N_24937,N_24249,N_24460);
and U24938 (N_24938,N_24140,N_24375);
xnor U24939 (N_24939,N_24380,N_24358);
and U24940 (N_24940,N_24252,N_24027);
nor U24941 (N_24941,N_24471,N_24275);
xor U24942 (N_24942,N_24114,N_24472);
nand U24943 (N_24943,N_24235,N_24203);
xnor U24944 (N_24944,N_24110,N_24428);
xor U24945 (N_24945,N_24164,N_24423);
and U24946 (N_24946,N_24062,N_24010);
and U24947 (N_24947,N_24420,N_24432);
nor U24948 (N_24948,N_24117,N_24407);
nor U24949 (N_24949,N_24018,N_24258);
and U24950 (N_24950,N_24477,N_24264);
nor U24951 (N_24951,N_24150,N_24353);
or U24952 (N_24952,N_24476,N_24417);
or U24953 (N_24953,N_24109,N_24352);
xnor U24954 (N_24954,N_24389,N_24408);
xor U24955 (N_24955,N_24054,N_24348);
or U24956 (N_24956,N_24103,N_24356);
and U24957 (N_24957,N_24094,N_24191);
and U24958 (N_24958,N_24349,N_24303);
or U24959 (N_24959,N_24274,N_24183);
xor U24960 (N_24960,N_24246,N_24205);
and U24961 (N_24961,N_24002,N_24419);
nand U24962 (N_24962,N_24425,N_24160);
xor U24963 (N_24963,N_24178,N_24385);
nand U24964 (N_24964,N_24243,N_24375);
or U24965 (N_24965,N_24194,N_24079);
xnor U24966 (N_24966,N_24442,N_24066);
or U24967 (N_24967,N_24477,N_24422);
xor U24968 (N_24968,N_24353,N_24272);
and U24969 (N_24969,N_24019,N_24133);
or U24970 (N_24970,N_24225,N_24318);
nor U24971 (N_24971,N_24366,N_24050);
and U24972 (N_24972,N_24482,N_24020);
nand U24973 (N_24973,N_24198,N_24012);
nor U24974 (N_24974,N_24162,N_24479);
nand U24975 (N_24975,N_24473,N_24200);
nand U24976 (N_24976,N_24105,N_24342);
or U24977 (N_24977,N_24012,N_24078);
nand U24978 (N_24978,N_24109,N_24428);
nand U24979 (N_24979,N_24436,N_24135);
or U24980 (N_24980,N_24164,N_24042);
nand U24981 (N_24981,N_24164,N_24122);
nand U24982 (N_24982,N_24024,N_24326);
nand U24983 (N_24983,N_24001,N_24206);
xor U24984 (N_24984,N_24253,N_24422);
nor U24985 (N_24985,N_24024,N_24488);
nand U24986 (N_24986,N_24011,N_24462);
xor U24987 (N_24987,N_24316,N_24266);
nor U24988 (N_24988,N_24199,N_24255);
xor U24989 (N_24989,N_24295,N_24159);
nand U24990 (N_24990,N_24180,N_24412);
nor U24991 (N_24991,N_24057,N_24472);
xor U24992 (N_24992,N_24040,N_24473);
nand U24993 (N_24993,N_24456,N_24437);
or U24994 (N_24994,N_24121,N_24497);
and U24995 (N_24995,N_24377,N_24208);
or U24996 (N_24996,N_24157,N_24329);
and U24997 (N_24997,N_24280,N_24291);
nor U24998 (N_24998,N_24093,N_24494);
nor U24999 (N_24999,N_24132,N_24305);
nor UO_0 (O_0,N_24783,N_24716);
xnor UO_1 (O_1,N_24744,N_24515);
nor UO_2 (O_2,N_24642,N_24750);
or UO_3 (O_3,N_24868,N_24651);
nand UO_4 (O_4,N_24977,N_24964);
nand UO_5 (O_5,N_24724,N_24732);
nor UO_6 (O_6,N_24892,N_24826);
and UO_7 (O_7,N_24796,N_24999);
xor UO_8 (O_8,N_24959,N_24659);
and UO_9 (O_9,N_24710,N_24720);
nor UO_10 (O_10,N_24504,N_24535);
nor UO_11 (O_11,N_24658,N_24996);
xnor UO_12 (O_12,N_24616,N_24987);
and UO_13 (O_13,N_24995,N_24828);
xor UO_14 (O_14,N_24787,N_24564);
and UO_15 (O_15,N_24685,N_24681);
and UO_16 (O_16,N_24972,N_24589);
nand UO_17 (O_17,N_24877,N_24638);
xor UO_18 (O_18,N_24738,N_24981);
or UO_19 (O_19,N_24915,N_24761);
xnor UO_20 (O_20,N_24810,N_24654);
or UO_21 (O_21,N_24852,N_24907);
or UO_22 (O_22,N_24553,N_24676);
or UO_23 (O_23,N_24517,N_24864);
or UO_24 (O_24,N_24530,N_24572);
nor UO_25 (O_25,N_24576,N_24962);
nor UO_26 (O_26,N_24760,N_24719);
and UO_27 (O_27,N_24910,N_24934);
or UO_28 (O_28,N_24832,N_24963);
nor UO_29 (O_29,N_24920,N_24500);
and UO_30 (O_30,N_24578,N_24836);
and UO_31 (O_31,N_24742,N_24938);
and UO_32 (O_32,N_24694,N_24903);
nand UO_33 (O_33,N_24745,N_24729);
xnor UO_34 (O_34,N_24509,N_24524);
nand UO_35 (O_35,N_24667,N_24919);
xnor UO_36 (O_36,N_24876,N_24687);
nand UO_37 (O_37,N_24726,N_24768);
nor UO_38 (O_38,N_24606,N_24725);
nand UO_39 (O_39,N_24649,N_24799);
nor UO_40 (O_40,N_24521,N_24639);
nor UO_41 (O_41,N_24753,N_24717);
xor UO_42 (O_42,N_24974,N_24709);
xnor UO_43 (O_43,N_24603,N_24531);
or UO_44 (O_44,N_24532,N_24645);
and UO_45 (O_45,N_24880,N_24887);
xor UO_46 (O_46,N_24775,N_24680);
and UO_47 (O_47,N_24594,N_24759);
or UO_48 (O_48,N_24611,N_24911);
or UO_49 (O_49,N_24948,N_24714);
xnor UO_50 (O_50,N_24516,N_24954);
xnor UO_51 (O_51,N_24537,N_24854);
nand UO_52 (O_52,N_24627,N_24730);
xnor UO_53 (O_53,N_24733,N_24824);
nor UO_54 (O_54,N_24957,N_24841);
xnor UO_55 (O_55,N_24812,N_24949);
and UO_56 (O_56,N_24794,N_24558);
nor UO_57 (O_57,N_24704,N_24891);
nand UO_58 (O_58,N_24648,N_24825);
nor UO_59 (O_59,N_24830,N_24707);
and UO_60 (O_60,N_24511,N_24644);
or UO_61 (O_61,N_24908,N_24533);
and UO_62 (O_62,N_24966,N_24757);
nor UO_63 (O_63,N_24931,N_24538);
nand UO_64 (O_64,N_24529,N_24984);
and UO_65 (O_65,N_24574,N_24789);
nand UO_66 (O_66,N_24879,N_24874);
or UO_67 (O_67,N_24665,N_24857);
xor UO_68 (O_68,N_24690,N_24613);
and UO_69 (O_69,N_24628,N_24698);
nor UO_70 (O_70,N_24855,N_24608);
or UO_71 (O_71,N_24534,N_24695);
nand UO_72 (O_72,N_24782,N_24711);
nand UO_73 (O_73,N_24850,N_24506);
nand UO_74 (O_74,N_24541,N_24741);
nand UO_75 (O_75,N_24615,N_24814);
and UO_76 (O_76,N_24755,N_24878);
and UO_77 (O_77,N_24942,N_24840);
and UO_78 (O_78,N_24788,N_24839);
and UO_79 (O_79,N_24581,N_24847);
nor UO_80 (O_80,N_24985,N_24833);
xnor UO_81 (O_81,N_24863,N_24860);
xor UO_82 (O_82,N_24663,N_24945);
or UO_83 (O_83,N_24519,N_24604);
and UO_84 (O_84,N_24993,N_24823);
and UO_85 (O_85,N_24944,N_24846);
and UO_86 (O_86,N_24688,N_24899);
nand UO_87 (O_87,N_24595,N_24666);
or UO_88 (O_88,N_24712,N_24890);
and UO_89 (O_89,N_24965,N_24967);
or UO_90 (O_90,N_24804,N_24776);
or UO_91 (O_91,N_24801,N_24583);
nand UO_92 (O_92,N_24937,N_24701);
nor UO_93 (O_93,N_24612,N_24913);
xor UO_94 (O_94,N_24808,N_24731);
nor UO_95 (O_95,N_24629,N_24871);
and UO_96 (O_96,N_24545,N_24893);
xor UO_97 (O_97,N_24691,N_24643);
or UO_98 (O_98,N_24622,N_24684);
xnor UO_99 (O_99,N_24702,N_24718);
xnor UO_100 (O_100,N_24941,N_24542);
and UO_101 (O_101,N_24652,N_24673);
or UO_102 (O_102,N_24609,N_24885);
nand UO_103 (O_103,N_24922,N_24988);
or UO_104 (O_104,N_24669,N_24590);
nor UO_105 (O_105,N_24953,N_24861);
and UO_106 (O_106,N_24565,N_24647);
or UO_107 (O_107,N_24921,N_24559);
xnor UO_108 (O_108,N_24582,N_24822);
nand UO_109 (O_109,N_24528,N_24844);
or UO_110 (O_110,N_24754,N_24924);
xnor UO_111 (O_111,N_24682,N_24932);
nor UO_112 (O_112,N_24633,N_24873);
nand UO_113 (O_113,N_24561,N_24708);
nand UO_114 (O_114,N_24894,N_24930);
nor UO_115 (O_115,N_24765,N_24785);
nand UO_116 (O_116,N_24668,N_24929);
and UO_117 (O_117,N_24939,N_24856);
or UO_118 (O_118,N_24955,N_24512);
or UO_119 (O_119,N_24811,N_24976);
nand UO_120 (O_120,N_24579,N_24816);
or UO_121 (O_121,N_24971,N_24722);
nand UO_122 (O_122,N_24831,N_24563);
and UO_123 (O_123,N_24943,N_24909);
or UO_124 (O_124,N_24715,N_24970);
xor UO_125 (O_125,N_24566,N_24835);
and UO_126 (O_126,N_24961,N_24838);
nand UO_127 (O_127,N_24580,N_24997);
nor UO_128 (O_128,N_24916,N_24900);
and UO_129 (O_129,N_24888,N_24540);
xnor UO_130 (O_130,N_24862,N_24557);
xor UO_131 (O_131,N_24980,N_24853);
and UO_132 (O_132,N_24774,N_24653);
nor UO_133 (O_133,N_24593,N_24912);
and UO_134 (O_134,N_24727,N_24568);
nand UO_135 (O_135,N_24552,N_24706);
xor UO_136 (O_136,N_24544,N_24735);
nor UO_137 (O_137,N_24827,N_24798);
xnor UO_138 (O_138,N_24771,N_24842);
or UO_139 (O_139,N_24905,N_24554);
nor UO_140 (O_140,N_24763,N_24756);
nor UO_141 (O_141,N_24821,N_24983);
nor UO_142 (O_142,N_24562,N_24547);
or UO_143 (O_143,N_24640,N_24619);
xor UO_144 (O_144,N_24518,N_24998);
nor UO_145 (O_145,N_24881,N_24870);
nor UO_146 (O_146,N_24600,N_24591);
or UO_147 (O_147,N_24713,N_24536);
nor UO_148 (O_148,N_24897,N_24992);
xor UO_149 (O_149,N_24661,N_24869);
and UO_150 (O_150,N_24677,N_24940);
nand UO_151 (O_151,N_24752,N_24620);
xnor UO_152 (O_152,N_24797,N_24867);
nor UO_153 (O_153,N_24906,N_24599);
nand UO_154 (O_154,N_24898,N_24587);
nand UO_155 (O_155,N_24660,N_24927);
xnor UO_156 (O_156,N_24889,N_24960);
nand UO_157 (O_157,N_24859,N_24866);
xnor UO_158 (O_158,N_24696,N_24807);
nor UO_159 (O_159,N_24969,N_24630);
or UO_160 (O_160,N_24723,N_24806);
nor UO_161 (O_161,N_24597,N_24560);
nor UO_162 (O_162,N_24692,N_24767);
and UO_163 (O_163,N_24896,N_24555);
nand UO_164 (O_164,N_24770,N_24751);
or UO_165 (O_165,N_24602,N_24994);
xnor UO_166 (O_166,N_24820,N_24664);
and UO_167 (O_167,N_24634,N_24539);
nand UO_168 (O_168,N_24523,N_24918);
xor UO_169 (O_169,N_24721,N_24845);
nand UO_170 (O_170,N_24550,N_24952);
nor UO_171 (O_171,N_24749,N_24543);
xnor UO_172 (O_172,N_24675,N_24739);
nand UO_173 (O_173,N_24872,N_24657);
and UO_174 (O_174,N_24902,N_24784);
and UO_175 (O_175,N_24501,N_24883);
and UO_176 (O_176,N_24989,N_24570);
and UO_177 (O_177,N_24703,N_24503);
nand UO_178 (O_178,N_24809,N_24848);
xor UO_179 (O_179,N_24584,N_24813);
or UO_180 (O_180,N_24646,N_24520);
nor UO_181 (O_181,N_24551,N_24884);
and UO_182 (O_182,N_24607,N_24510);
or UO_183 (O_183,N_24700,N_24546);
and UO_184 (O_184,N_24655,N_24875);
and UO_185 (O_185,N_24746,N_24641);
and UO_186 (O_186,N_24740,N_24849);
xnor UO_187 (O_187,N_24705,N_24777);
nor UO_188 (O_188,N_24513,N_24936);
and UO_189 (O_189,N_24650,N_24548);
xor UO_190 (O_190,N_24951,N_24697);
nor UO_191 (O_191,N_24671,N_24636);
nor UO_192 (O_192,N_24901,N_24508);
nor UO_193 (O_193,N_24973,N_24829);
and UO_194 (O_194,N_24837,N_24780);
nand UO_195 (O_195,N_24772,N_24800);
nand UO_196 (O_196,N_24773,N_24573);
and UO_197 (O_197,N_24736,N_24577);
and UO_198 (O_198,N_24758,N_24699);
and UO_199 (O_199,N_24928,N_24502);
nand UO_200 (O_200,N_24769,N_24689);
nand UO_201 (O_201,N_24527,N_24817);
xnor UO_202 (O_202,N_24851,N_24743);
or UO_203 (O_203,N_24637,N_24882);
and UO_204 (O_204,N_24567,N_24623);
or UO_205 (O_205,N_24764,N_24693);
and UO_206 (O_206,N_24670,N_24815);
xnor UO_207 (O_207,N_24596,N_24786);
or UO_208 (O_208,N_24865,N_24610);
xor UO_209 (O_209,N_24781,N_24991);
and UO_210 (O_210,N_24592,N_24819);
or UO_211 (O_211,N_24686,N_24818);
nor UO_212 (O_212,N_24935,N_24805);
and UO_213 (O_213,N_24762,N_24946);
xnor UO_214 (O_214,N_24923,N_24895);
xor UO_215 (O_215,N_24631,N_24656);
nor UO_216 (O_216,N_24978,N_24979);
xor UO_217 (O_217,N_24626,N_24975);
and UO_218 (O_218,N_24526,N_24926);
nand UO_219 (O_219,N_24625,N_24958);
or UO_220 (O_220,N_24614,N_24575);
xor UO_221 (O_221,N_24933,N_24683);
and UO_222 (O_222,N_24635,N_24621);
and UO_223 (O_223,N_24632,N_24734);
and UO_224 (O_224,N_24522,N_24605);
xnor UO_225 (O_225,N_24858,N_24950);
nor UO_226 (O_226,N_24766,N_24586);
nand UO_227 (O_227,N_24737,N_24779);
nor UO_228 (O_228,N_24514,N_24803);
nor UO_229 (O_229,N_24549,N_24598);
nand UO_230 (O_230,N_24601,N_24505);
and UO_231 (O_231,N_24748,N_24624);
or UO_232 (O_232,N_24507,N_24588);
xor UO_233 (O_233,N_24556,N_24778);
and UO_234 (O_234,N_24982,N_24569);
nand UO_235 (O_235,N_24618,N_24792);
or UO_236 (O_236,N_24674,N_24585);
xnor UO_237 (O_237,N_24917,N_24747);
nand UO_238 (O_238,N_24793,N_24678);
nand UO_239 (O_239,N_24843,N_24802);
nor UO_240 (O_240,N_24791,N_24990);
or UO_241 (O_241,N_24956,N_24790);
and UO_242 (O_242,N_24986,N_24662);
nand UO_243 (O_243,N_24795,N_24525);
nor UO_244 (O_244,N_24728,N_24672);
xor UO_245 (O_245,N_24617,N_24834);
and UO_246 (O_246,N_24914,N_24947);
xor UO_247 (O_247,N_24886,N_24968);
and UO_248 (O_248,N_24571,N_24679);
nand UO_249 (O_249,N_24925,N_24904);
xnor UO_250 (O_250,N_24592,N_24808);
nor UO_251 (O_251,N_24538,N_24541);
nor UO_252 (O_252,N_24961,N_24611);
nand UO_253 (O_253,N_24500,N_24768);
nor UO_254 (O_254,N_24503,N_24551);
xnor UO_255 (O_255,N_24519,N_24592);
xnor UO_256 (O_256,N_24677,N_24795);
xnor UO_257 (O_257,N_24721,N_24653);
nand UO_258 (O_258,N_24983,N_24927);
xor UO_259 (O_259,N_24724,N_24576);
and UO_260 (O_260,N_24947,N_24636);
nor UO_261 (O_261,N_24831,N_24661);
xor UO_262 (O_262,N_24748,N_24812);
and UO_263 (O_263,N_24746,N_24952);
nand UO_264 (O_264,N_24795,N_24948);
nor UO_265 (O_265,N_24807,N_24987);
and UO_266 (O_266,N_24524,N_24640);
or UO_267 (O_267,N_24774,N_24706);
nor UO_268 (O_268,N_24544,N_24778);
nand UO_269 (O_269,N_24885,N_24987);
and UO_270 (O_270,N_24931,N_24789);
nand UO_271 (O_271,N_24633,N_24588);
or UO_272 (O_272,N_24519,N_24607);
and UO_273 (O_273,N_24863,N_24742);
nand UO_274 (O_274,N_24544,N_24955);
nand UO_275 (O_275,N_24619,N_24527);
and UO_276 (O_276,N_24692,N_24995);
nand UO_277 (O_277,N_24752,N_24932);
xor UO_278 (O_278,N_24625,N_24896);
xor UO_279 (O_279,N_24739,N_24898);
and UO_280 (O_280,N_24697,N_24905);
nor UO_281 (O_281,N_24826,N_24776);
or UO_282 (O_282,N_24502,N_24886);
nor UO_283 (O_283,N_24504,N_24541);
nand UO_284 (O_284,N_24603,N_24590);
xnor UO_285 (O_285,N_24546,N_24985);
or UO_286 (O_286,N_24793,N_24596);
nand UO_287 (O_287,N_24517,N_24986);
xnor UO_288 (O_288,N_24732,N_24690);
nor UO_289 (O_289,N_24766,N_24920);
and UO_290 (O_290,N_24774,N_24961);
or UO_291 (O_291,N_24968,N_24887);
and UO_292 (O_292,N_24692,N_24614);
nor UO_293 (O_293,N_24975,N_24574);
and UO_294 (O_294,N_24907,N_24705);
and UO_295 (O_295,N_24742,N_24670);
nand UO_296 (O_296,N_24807,N_24731);
xor UO_297 (O_297,N_24962,N_24667);
nand UO_298 (O_298,N_24821,N_24690);
nor UO_299 (O_299,N_24558,N_24835);
or UO_300 (O_300,N_24651,N_24825);
xor UO_301 (O_301,N_24958,N_24676);
xnor UO_302 (O_302,N_24775,N_24610);
nor UO_303 (O_303,N_24707,N_24550);
or UO_304 (O_304,N_24594,N_24761);
or UO_305 (O_305,N_24615,N_24532);
xor UO_306 (O_306,N_24797,N_24565);
nand UO_307 (O_307,N_24939,N_24845);
and UO_308 (O_308,N_24628,N_24539);
xor UO_309 (O_309,N_24966,N_24942);
or UO_310 (O_310,N_24983,N_24565);
nand UO_311 (O_311,N_24694,N_24660);
and UO_312 (O_312,N_24667,N_24567);
nand UO_313 (O_313,N_24894,N_24999);
xnor UO_314 (O_314,N_24792,N_24520);
nor UO_315 (O_315,N_24835,N_24867);
xnor UO_316 (O_316,N_24959,N_24517);
or UO_317 (O_317,N_24838,N_24790);
nor UO_318 (O_318,N_24880,N_24557);
xnor UO_319 (O_319,N_24644,N_24727);
and UO_320 (O_320,N_24514,N_24913);
nor UO_321 (O_321,N_24530,N_24562);
xnor UO_322 (O_322,N_24562,N_24598);
xor UO_323 (O_323,N_24574,N_24526);
nor UO_324 (O_324,N_24793,N_24839);
nand UO_325 (O_325,N_24853,N_24997);
nor UO_326 (O_326,N_24669,N_24544);
or UO_327 (O_327,N_24738,N_24942);
nor UO_328 (O_328,N_24911,N_24938);
or UO_329 (O_329,N_24921,N_24617);
or UO_330 (O_330,N_24508,N_24737);
and UO_331 (O_331,N_24995,N_24623);
xor UO_332 (O_332,N_24817,N_24828);
xor UO_333 (O_333,N_24963,N_24851);
nand UO_334 (O_334,N_24743,N_24854);
and UO_335 (O_335,N_24815,N_24757);
nor UO_336 (O_336,N_24522,N_24957);
nor UO_337 (O_337,N_24749,N_24941);
or UO_338 (O_338,N_24540,N_24511);
nand UO_339 (O_339,N_24565,N_24894);
xnor UO_340 (O_340,N_24991,N_24922);
nand UO_341 (O_341,N_24904,N_24821);
nor UO_342 (O_342,N_24980,N_24532);
xor UO_343 (O_343,N_24512,N_24802);
nor UO_344 (O_344,N_24768,N_24561);
xnor UO_345 (O_345,N_24894,N_24884);
xnor UO_346 (O_346,N_24559,N_24950);
and UO_347 (O_347,N_24867,N_24718);
and UO_348 (O_348,N_24734,N_24881);
nor UO_349 (O_349,N_24880,N_24818);
and UO_350 (O_350,N_24729,N_24944);
or UO_351 (O_351,N_24944,N_24910);
xor UO_352 (O_352,N_24777,N_24716);
nand UO_353 (O_353,N_24551,N_24648);
nand UO_354 (O_354,N_24866,N_24516);
and UO_355 (O_355,N_24818,N_24783);
nand UO_356 (O_356,N_24712,N_24827);
and UO_357 (O_357,N_24740,N_24941);
nand UO_358 (O_358,N_24691,N_24737);
xnor UO_359 (O_359,N_24638,N_24965);
nor UO_360 (O_360,N_24661,N_24555);
nor UO_361 (O_361,N_24582,N_24958);
or UO_362 (O_362,N_24531,N_24550);
nand UO_363 (O_363,N_24917,N_24757);
or UO_364 (O_364,N_24594,N_24857);
or UO_365 (O_365,N_24536,N_24557);
nor UO_366 (O_366,N_24767,N_24592);
xnor UO_367 (O_367,N_24921,N_24554);
and UO_368 (O_368,N_24757,N_24569);
and UO_369 (O_369,N_24896,N_24728);
nand UO_370 (O_370,N_24637,N_24536);
or UO_371 (O_371,N_24663,N_24810);
xor UO_372 (O_372,N_24761,N_24981);
nor UO_373 (O_373,N_24999,N_24690);
nand UO_374 (O_374,N_24965,N_24692);
nand UO_375 (O_375,N_24578,N_24685);
and UO_376 (O_376,N_24603,N_24681);
nand UO_377 (O_377,N_24511,N_24701);
or UO_378 (O_378,N_24764,N_24537);
or UO_379 (O_379,N_24997,N_24748);
nand UO_380 (O_380,N_24594,N_24696);
or UO_381 (O_381,N_24715,N_24671);
nand UO_382 (O_382,N_24745,N_24934);
nor UO_383 (O_383,N_24545,N_24643);
nor UO_384 (O_384,N_24642,N_24939);
nand UO_385 (O_385,N_24940,N_24599);
nor UO_386 (O_386,N_24866,N_24625);
nand UO_387 (O_387,N_24664,N_24516);
nor UO_388 (O_388,N_24712,N_24634);
nor UO_389 (O_389,N_24696,N_24787);
or UO_390 (O_390,N_24710,N_24686);
and UO_391 (O_391,N_24797,N_24570);
nand UO_392 (O_392,N_24625,N_24886);
and UO_393 (O_393,N_24742,N_24773);
nor UO_394 (O_394,N_24959,N_24793);
nand UO_395 (O_395,N_24564,N_24773);
and UO_396 (O_396,N_24553,N_24767);
and UO_397 (O_397,N_24542,N_24849);
or UO_398 (O_398,N_24734,N_24864);
nor UO_399 (O_399,N_24868,N_24790);
nor UO_400 (O_400,N_24830,N_24760);
xor UO_401 (O_401,N_24987,N_24678);
or UO_402 (O_402,N_24607,N_24733);
and UO_403 (O_403,N_24510,N_24900);
or UO_404 (O_404,N_24983,N_24785);
or UO_405 (O_405,N_24907,N_24760);
and UO_406 (O_406,N_24534,N_24805);
xor UO_407 (O_407,N_24982,N_24898);
nand UO_408 (O_408,N_24553,N_24589);
xor UO_409 (O_409,N_24541,N_24933);
or UO_410 (O_410,N_24772,N_24844);
and UO_411 (O_411,N_24674,N_24549);
nor UO_412 (O_412,N_24630,N_24698);
or UO_413 (O_413,N_24839,N_24935);
xor UO_414 (O_414,N_24920,N_24794);
xor UO_415 (O_415,N_24947,N_24859);
or UO_416 (O_416,N_24833,N_24702);
nor UO_417 (O_417,N_24719,N_24961);
xnor UO_418 (O_418,N_24966,N_24796);
xnor UO_419 (O_419,N_24969,N_24690);
nand UO_420 (O_420,N_24602,N_24916);
or UO_421 (O_421,N_24893,N_24586);
nand UO_422 (O_422,N_24757,N_24764);
or UO_423 (O_423,N_24981,N_24769);
nand UO_424 (O_424,N_24588,N_24635);
nor UO_425 (O_425,N_24758,N_24504);
or UO_426 (O_426,N_24733,N_24671);
nor UO_427 (O_427,N_24773,N_24570);
and UO_428 (O_428,N_24529,N_24710);
and UO_429 (O_429,N_24898,N_24992);
and UO_430 (O_430,N_24602,N_24579);
nor UO_431 (O_431,N_24654,N_24733);
nor UO_432 (O_432,N_24956,N_24686);
or UO_433 (O_433,N_24600,N_24808);
and UO_434 (O_434,N_24980,N_24774);
xor UO_435 (O_435,N_24591,N_24950);
and UO_436 (O_436,N_24929,N_24572);
or UO_437 (O_437,N_24895,N_24590);
or UO_438 (O_438,N_24500,N_24982);
nor UO_439 (O_439,N_24962,N_24927);
xnor UO_440 (O_440,N_24994,N_24683);
and UO_441 (O_441,N_24981,N_24967);
and UO_442 (O_442,N_24890,N_24752);
and UO_443 (O_443,N_24716,N_24653);
nor UO_444 (O_444,N_24664,N_24607);
or UO_445 (O_445,N_24566,N_24689);
xor UO_446 (O_446,N_24887,N_24726);
and UO_447 (O_447,N_24937,N_24516);
nor UO_448 (O_448,N_24897,N_24512);
or UO_449 (O_449,N_24628,N_24917);
or UO_450 (O_450,N_24980,N_24509);
xor UO_451 (O_451,N_24558,N_24743);
xor UO_452 (O_452,N_24795,N_24558);
and UO_453 (O_453,N_24686,N_24537);
or UO_454 (O_454,N_24559,N_24612);
xnor UO_455 (O_455,N_24724,N_24887);
nand UO_456 (O_456,N_24709,N_24738);
and UO_457 (O_457,N_24731,N_24671);
and UO_458 (O_458,N_24903,N_24911);
or UO_459 (O_459,N_24520,N_24505);
or UO_460 (O_460,N_24577,N_24724);
or UO_461 (O_461,N_24620,N_24801);
and UO_462 (O_462,N_24984,N_24774);
or UO_463 (O_463,N_24510,N_24565);
or UO_464 (O_464,N_24893,N_24788);
and UO_465 (O_465,N_24642,N_24584);
xnor UO_466 (O_466,N_24611,N_24958);
and UO_467 (O_467,N_24717,N_24515);
nor UO_468 (O_468,N_24695,N_24599);
nand UO_469 (O_469,N_24937,N_24631);
nand UO_470 (O_470,N_24739,N_24592);
and UO_471 (O_471,N_24884,N_24692);
or UO_472 (O_472,N_24652,N_24832);
and UO_473 (O_473,N_24993,N_24926);
and UO_474 (O_474,N_24976,N_24796);
and UO_475 (O_475,N_24937,N_24675);
xor UO_476 (O_476,N_24744,N_24840);
nor UO_477 (O_477,N_24924,N_24591);
xnor UO_478 (O_478,N_24545,N_24848);
xor UO_479 (O_479,N_24955,N_24555);
or UO_480 (O_480,N_24940,N_24588);
nor UO_481 (O_481,N_24953,N_24603);
nor UO_482 (O_482,N_24886,N_24914);
nor UO_483 (O_483,N_24544,N_24910);
or UO_484 (O_484,N_24672,N_24700);
or UO_485 (O_485,N_24671,N_24831);
nor UO_486 (O_486,N_24989,N_24725);
xnor UO_487 (O_487,N_24910,N_24582);
nand UO_488 (O_488,N_24813,N_24690);
nor UO_489 (O_489,N_24783,N_24974);
nand UO_490 (O_490,N_24507,N_24517);
nor UO_491 (O_491,N_24801,N_24719);
nand UO_492 (O_492,N_24930,N_24987);
nand UO_493 (O_493,N_24706,N_24956);
nand UO_494 (O_494,N_24626,N_24587);
or UO_495 (O_495,N_24828,N_24571);
nand UO_496 (O_496,N_24786,N_24815);
and UO_497 (O_497,N_24845,N_24704);
nor UO_498 (O_498,N_24933,N_24572);
nor UO_499 (O_499,N_24997,N_24999);
xnor UO_500 (O_500,N_24726,N_24779);
nand UO_501 (O_501,N_24824,N_24725);
and UO_502 (O_502,N_24504,N_24645);
nor UO_503 (O_503,N_24563,N_24634);
xnor UO_504 (O_504,N_24874,N_24637);
xor UO_505 (O_505,N_24964,N_24542);
nand UO_506 (O_506,N_24716,N_24911);
or UO_507 (O_507,N_24783,N_24922);
nor UO_508 (O_508,N_24582,N_24867);
or UO_509 (O_509,N_24538,N_24758);
nor UO_510 (O_510,N_24794,N_24711);
and UO_511 (O_511,N_24654,N_24539);
or UO_512 (O_512,N_24530,N_24685);
xor UO_513 (O_513,N_24691,N_24723);
or UO_514 (O_514,N_24932,N_24733);
nand UO_515 (O_515,N_24845,N_24520);
nand UO_516 (O_516,N_24618,N_24760);
xnor UO_517 (O_517,N_24821,N_24590);
nand UO_518 (O_518,N_24983,N_24536);
and UO_519 (O_519,N_24716,N_24587);
nor UO_520 (O_520,N_24783,N_24809);
nand UO_521 (O_521,N_24523,N_24712);
nor UO_522 (O_522,N_24571,N_24797);
and UO_523 (O_523,N_24688,N_24784);
and UO_524 (O_524,N_24968,N_24874);
xnor UO_525 (O_525,N_24540,N_24616);
xor UO_526 (O_526,N_24853,N_24540);
nor UO_527 (O_527,N_24543,N_24684);
or UO_528 (O_528,N_24945,N_24779);
and UO_529 (O_529,N_24672,N_24599);
or UO_530 (O_530,N_24704,N_24546);
nor UO_531 (O_531,N_24698,N_24617);
xor UO_532 (O_532,N_24947,N_24662);
or UO_533 (O_533,N_24739,N_24846);
and UO_534 (O_534,N_24984,N_24626);
xor UO_535 (O_535,N_24677,N_24709);
or UO_536 (O_536,N_24604,N_24809);
nor UO_537 (O_537,N_24538,N_24559);
or UO_538 (O_538,N_24965,N_24818);
or UO_539 (O_539,N_24598,N_24601);
xor UO_540 (O_540,N_24610,N_24617);
or UO_541 (O_541,N_24700,N_24791);
or UO_542 (O_542,N_24979,N_24671);
nor UO_543 (O_543,N_24885,N_24604);
xor UO_544 (O_544,N_24744,N_24539);
nor UO_545 (O_545,N_24874,N_24609);
and UO_546 (O_546,N_24692,N_24904);
nand UO_547 (O_547,N_24685,N_24852);
and UO_548 (O_548,N_24735,N_24667);
nor UO_549 (O_549,N_24852,N_24756);
or UO_550 (O_550,N_24742,N_24666);
nand UO_551 (O_551,N_24816,N_24955);
xnor UO_552 (O_552,N_24600,N_24930);
and UO_553 (O_553,N_24968,N_24916);
or UO_554 (O_554,N_24579,N_24765);
and UO_555 (O_555,N_24714,N_24738);
nand UO_556 (O_556,N_24687,N_24766);
xnor UO_557 (O_557,N_24654,N_24738);
nor UO_558 (O_558,N_24959,N_24804);
nor UO_559 (O_559,N_24960,N_24969);
or UO_560 (O_560,N_24571,N_24605);
nand UO_561 (O_561,N_24658,N_24501);
xnor UO_562 (O_562,N_24872,N_24925);
or UO_563 (O_563,N_24731,N_24888);
or UO_564 (O_564,N_24620,N_24510);
and UO_565 (O_565,N_24967,N_24970);
nand UO_566 (O_566,N_24881,N_24972);
nand UO_567 (O_567,N_24937,N_24557);
xor UO_568 (O_568,N_24722,N_24881);
nand UO_569 (O_569,N_24872,N_24650);
nand UO_570 (O_570,N_24666,N_24788);
and UO_571 (O_571,N_24950,N_24655);
or UO_572 (O_572,N_24733,N_24748);
xor UO_573 (O_573,N_24606,N_24630);
xor UO_574 (O_574,N_24624,N_24668);
nor UO_575 (O_575,N_24717,N_24531);
xnor UO_576 (O_576,N_24661,N_24741);
xor UO_577 (O_577,N_24871,N_24694);
nor UO_578 (O_578,N_24818,N_24901);
nor UO_579 (O_579,N_24880,N_24788);
xor UO_580 (O_580,N_24951,N_24941);
nand UO_581 (O_581,N_24656,N_24799);
xnor UO_582 (O_582,N_24736,N_24842);
and UO_583 (O_583,N_24793,N_24559);
nor UO_584 (O_584,N_24949,N_24749);
xnor UO_585 (O_585,N_24697,N_24902);
and UO_586 (O_586,N_24780,N_24597);
nand UO_587 (O_587,N_24679,N_24622);
or UO_588 (O_588,N_24819,N_24964);
or UO_589 (O_589,N_24648,N_24514);
xnor UO_590 (O_590,N_24854,N_24657);
xnor UO_591 (O_591,N_24515,N_24695);
nor UO_592 (O_592,N_24595,N_24890);
xnor UO_593 (O_593,N_24898,N_24639);
nor UO_594 (O_594,N_24539,N_24694);
nand UO_595 (O_595,N_24789,N_24924);
nor UO_596 (O_596,N_24777,N_24869);
xor UO_597 (O_597,N_24851,N_24784);
or UO_598 (O_598,N_24687,N_24522);
xnor UO_599 (O_599,N_24857,N_24728);
nand UO_600 (O_600,N_24562,N_24920);
or UO_601 (O_601,N_24755,N_24881);
nand UO_602 (O_602,N_24921,N_24700);
xor UO_603 (O_603,N_24776,N_24540);
and UO_604 (O_604,N_24785,N_24707);
nand UO_605 (O_605,N_24593,N_24921);
nor UO_606 (O_606,N_24689,N_24606);
and UO_607 (O_607,N_24945,N_24520);
or UO_608 (O_608,N_24881,N_24635);
or UO_609 (O_609,N_24985,N_24816);
nand UO_610 (O_610,N_24881,N_24551);
nor UO_611 (O_611,N_24991,N_24960);
nand UO_612 (O_612,N_24733,N_24735);
or UO_613 (O_613,N_24965,N_24974);
nor UO_614 (O_614,N_24746,N_24616);
or UO_615 (O_615,N_24725,N_24564);
xnor UO_616 (O_616,N_24502,N_24686);
and UO_617 (O_617,N_24568,N_24524);
and UO_618 (O_618,N_24774,N_24698);
or UO_619 (O_619,N_24974,N_24994);
and UO_620 (O_620,N_24740,N_24663);
nand UO_621 (O_621,N_24973,N_24995);
nand UO_622 (O_622,N_24509,N_24630);
and UO_623 (O_623,N_24515,N_24795);
and UO_624 (O_624,N_24700,N_24749);
xor UO_625 (O_625,N_24856,N_24522);
and UO_626 (O_626,N_24721,N_24960);
nand UO_627 (O_627,N_24996,N_24516);
xnor UO_628 (O_628,N_24721,N_24930);
nor UO_629 (O_629,N_24939,N_24826);
and UO_630 (O_630,N_24837,N_24670);
or UO_631 (O_631,N_24948,N_24578);
or UO_632 (O_632,N_24690,N_24538);
or UO_633 (O_633,N_24954,N_24742);
xor UO_634 (O_634,N_24589,N_24744);
nand UO_635 (O_635,N_24940,N_24512);
nor UO_636 (O_636,N_24660,N_24899);
nand UO_637 (O_637,N_24646,N_24515);
and UO_638 (O_638,N_24992,N_24725);
xor UO_639 (O_639,N_24836,N_24974);
and UO_640 (O_640,N_24856,N_24656);
nor UO_641 (O_641,N_24916,N_24556);
and UO_642 (O_642,N_24639,N_24537);
xor UO_643 (O_643,N_24789,N_24893);
or UO_644 (O_644,N_24747,N_24834);
or UO_645 (O_645,N_24524,N_24536);
xnor UO_646 (O_646,N_24836,N_24860);
and UO_647 (O_647,N_24652,N_24565);
nand UO_648 (O_648,N_24953,N_24672);
or UO_649 (O_649,N_24991,N_24507);
nand UO_650 (O_650,N_24749,N_24836);
xor UO_651 (O_651,N_24786,N_24858);
nand UO_652 (O_652,N_24664,N_24788);
and UO_653 (O_653,N_24692,N_24660);
nor UO_654 (O_654,N_24786,N_24691);
nand UO_655 (O_655,N_24887,N_24896);
or UO_656 (O_656,N_24627,N_24600);
and UO_657 (O_657,N_24850,N_24593);
xnor UO_658 (O_658,N_24566,N_24597);
nand UO_659 (O_659,N_24609,N_24672);
and UO_660 (O_660,N_24658,N_24535);
nand UO_661 (O_661,N_24706,N_24753);
nor UO_662 (O_662,N_24533,N_24506);
nor UO_663 (O_663,N_24846,N_24600);
xnor UO_664 (O_664,N_24651,N_24718);
xor UO_665 (O_665,N_24561,N_24993);
nand UO_666 (O_666,N_24877,N_24531);
and UO_667 (O_667,N_24772,N_24694);
nand UO_668 (O_668,N_24688,N_24851);
nand UO_669 (O_669,N_24538,N_24912);
and UO_670 (O_670,N_24805,N_24812);
or UO_671 (O_671,N_24842,N_24536);
or UO_672 (O_672,N_24579,N_24519);
nor UO_673 (O_673,N_24585,N_24740);
and UO_674 (O_674,N_24602,N_24810);
nand UO_675 (O_675,N_24694,N_24619);
nor UO_676 (O_676,N_24717,N_24631);
nor UO_677 (O_677,N_24704,N_24823);
and UO_678 (O_678,N_24580,N_24648);
nand UO_679 (O_679,N_24677,N_24936);
or UO_680 (O_680,N_24741,N_24968);
xor UO_681 (O_681,N_24542,N_24870);
xnor UO_682 (O_682,N_24918,N_24540);
xor UO_683 (O_683,N_24619,N_24712);
nor UO_684 (O_684,N_24784,N_24982);
and UO_685 (O_685,N_24650,N_24697);
nor UO_686 (O_686,N_24682,N_24772);
nor UO_687 (O_687,N_24642,N_24997);
nor UO_688 (O_688,N_24585,N_24500);
or UO_689 (O_689,N_24514,N_24558);
or UO_690 (O_690,N_24513,N_24905);
nor UO_691 (O_691,N_24924,N_24521);
nor UO_692 (O_692,N_24727,N_24632);
or UO_693 (O_693,N_24984,N_24730);
or UO_694 (O_694,N_24630,N_24761);
and UO_695 (O_695,N_24987,N_24687);
and UO_696 (O_696,N_24519,N_24633);
xor UO_697 (O_697,N_24726,N_24580);
and UO_698 (O_698,N_24751,N_24676);
or UO_699 (O_699,N_24535,N_24828);
and UO_700 (O_700,N_24605,N_24889);
nor UO_701 (O_701,N_24514,N_24804);
xnor UO_702 (O_702,N_24795,N_24544);
nand UO_703 (O_703,N_24939,N_24730);
nor UO_704 (O_704,N_24595,N_24635);
nor UO_705 (O_705,N_24752,N_24939);
nor UO_706 (O_706,N_24643,N_24700);
or UO_707 (O_707,N_24589,N_24969);
or UO_708 (O_708,N_24515,N_24849);
nor UO_709 (O_709,N_24807,N_24983);
nor UO_710 (O_710,N_24966,N_24688);
xor UO_711 (O_711,N_24563,N_24523);
or UO_712 (O_712,N_24577,N_24970);
nor UO_713 (O_713,N_24558,N_24675);
and UO_714 (O_714,N_24639,N_24648);
or UO_715 (O_715,N_24816,N_24827);
or UO_716 (O_716,N_24834,N_24551);
and UO_717 (O_717,N_24661,N_24513);
or UO_718 (O_718,N_24559,N_24929);
nand UO_719 (O_719,N_24597,N_24809);
nor UO_720 (O_720,N_24589,N_24795);
nor UO_721 (O_721,N_24702,N_24735);
xor UO_722 (O_722,N_24714,N_24728);
nand UO_723 (O_723,N_24731,N_24618);
nor UO_724 (O_724,N_24884,N_24989);
xor UO_725 (O_725,N_24775,N_24803);
nor UO_726 (O_726,N_24500,N_24566);
nor UO_727 (O_727,N_24738,N_24972);
and UO_728 (O_728,N_24905,N_24850);
xnor UO_729 (O_729,N_24691,N_24907);
or UO_730 (O_730,N_24778,N_24989);
nor UO_731 (O_731,N_24643,N_24506);
nand UO_732 (O_732,N_24705,N_24828);
or UO_733 (O_733,N_24537,N_24557);
nand UO_734 (O_734,N_24868,N_24655);
or UO_735 (O_735,N_24742,N_24538);
or UO_736 (O_736,N_24654,N_24961);
or UO_737 (O_737,N_24793,N_24626);
nor UO_738 (O_738,N_24512,N_24774);
or UO_739 (O_739,N_24552,N_24634);
nand UO_740 (O_740,N_24940,N_24979);
or UO_741 (O_741,N_24932,N_24981);
nand UO_742 (O_742,N_24855,N_24500);
nor UO_743 (O_743,N_24764,N_24862);
xor UO_744 (O_744,N_24595,N_24530);
or UO_745 (O_745,N_24714,N_24696);
xnor UO_746 (O_746,N_24575,N_24532);
nand UO_747 (O_747,N_24715,N_24667);
nor UO_748 (O_748,N_24517,N_24712);
xor UO_749 (O_749,N_24917,N_24801);
or UO_750 (O_750,N_24640,N_24838);
nand UO_751 (O_751,N_24658,N_24543);
nand UO_752 (O_752,N_24892,N_24852);
and UO_753 (O_753,N_24745,N_24549);
xor UO_754 (O_754,N_24978,N_24793);
and UO_755 (O_755,N_24770,N_24558);
nor UO_756 (O_756,N_24615,N_24823);
nor UO_757 (O_757,N_24732,N_24549);
and UO_758 (O_758,N_24979,N_24855);
nand UO_759 (O_759,N_24582,N_24678);
nor UO_760 (O_760,N_24922,N_24694);
nand UO_761 (O_761,N_24956,N_24501);
xor UO_762 (O_762,N_24719,N_24942);
and UO_763 (O_763,N_24802,N_24788);
xor UO_764 (O_764,N_24859,N_24954);
nand UO_765 (O_765,N_24596,N_24961);
and UO_766 (O_766,N_24575,N_24744);
or UO_767 (O_767,N_24848,N_24857);
xnor UO_768 (O_768,N_24506,N_24653);
nor UO_769 (O_769,N_24981,N_24787);
nor UO_770 (O_770,N_24776,N_24796);
xor UO_771 (O_771,N_24913,N_24990);
or UO_772 (O_772,N_24916,N_24865);
nand UO_773 (O_773,N_24862,N_24610);
xor UO_774 (O_774,N_24760,N_24877);
nor UO_775 (O_775,N_24574,N_24809);
or UO_776 (O_776,N_24787,N_24783);
nor UO_777 (O_777,N_24963,N_24888);
or UO_778 (O_778,N_24612,N_24527);
and UO_779 (O_779,N_24577,N_24610);
xnor UO_780 (O_780,N_24595,N_24585);
or UO_781 (O_781,N_24770,N_24937);
and UO_782 (O_782,N_24752,N_24732);
nor UO_783 (O_783,N_24947,N_24924);
xor UO_784 (O_784,N_24934,N_24568);
nor UO_785 (O_785,N_24902,N_24985);
and UO_786 (O_786,N_24905,N_24765);
nand UO_787 (O_787,N_24863,N_24824);
and UO_788 (O_788,N_24542,N_24695);
nor UO_789 (O_789,N_24977,N_24648);
nor UO_790 (O_790,N_24687,N_24943);
nand UO_791 (O_791,N_24969,N_24730);
nor UO_792 (O_792,N_24673,N_24557);
and UO_793 (O_793,N_24856,N_24507);
nor UO_794 (O_794,N_24676,N_24576);
or UO_795 (O_795,N_24548,N_24995);
xor UO_796 (O_796,N_24700,N_24513);
nand UO_797 (O_797,N_24859,N_24801);
nor UO_798 (O_798,N_24953,N_24823);
nand UO_799 (O_799,N_24776,N_24680);
and UO_800 (O_800,N_24960,N_24655);
or UO_801 (O_801,N_24550,N_24534);
and UO_802 (O_802,N_24522,N_24586);
nor UO_803 (O_803,N_24871,N_24557);
or UO_804 (O_804,N_24671,N_24718);
xnor UO_805 (O_805,N_24945,N_24935);
nor UO_806 (O_806,N_24920,N_24574);
and UO_807 (O_807,N_24637,N_24985);
or UO_808 (O_808,N_24574,N_24834);
and UO_809 (O_809,N_24511,N_24506);
and UO_810 (O_810,N_24533,N_24527);
and UO_811 (O_811,N_24844,N_24799);
nand UO_812 (O_812,N_24800,N_24534);
nand UO_813 (O_813,N_24716,N_24842);
or UO_814 (O_814,N_24815,N_24609);
xor UO_815 (O_815,N_24766,N_24720);
xnor UO_816 (O_816,N_24737,N_24653);
or UO_817 (O_817,N_24765,N_24887);
xor UO_818 (O_818,N_24603,N_24706);
and UO_819 (O_819,N_24868,N_24716);
and UO_820 (O_820,N_24946,N_24765);
nand UO_821 (O_821,N_24706,N_24610);
or UO_822 (O_822,N_24561,N_24901);
or UO_823 (O_823,N_24669,N_24908);
nand UO_824 (O_824,N_24994,N_24531);
xor UO_825 (O_825,N_24904,N_24727);
nand UO_826 (O_826,N_24705,N_24709);
xnor UO_827 (O_827,N_24559,N_24953);
nand UO_828 (O_828,N_24850,N_24537);
and UO_829 (O_829,N_24846,N_24512);
nand UO_830 (O_830,N_24788,N_24900);
and UO_831 (O_831,N_24717,N_24874);
or UO_832 (O_832,N_24902,N_24560);
and UO_833 (O_833,N_24952,N_24545);
nand UO_834 (O_834,N_24670,N_24921);
nor UO_835 (O_835,N_24837,N_24642);
xor UO_836 (O_836,N_24543,N_24668);
or UO_837 (O_837,N_24637,N_24986);
nand UO_838 (O_838,N_24787,N_24639);
and UO_839 (O_839,N_24553,N_24698);
or UO_840 (O_840,N_24882,N_24835);
nor UO_841 (O_841,N_24888,N_24645);
nand UO_842 (O_842,N_24763,N_24724);
or UO_843 (O_843,N_24633,N_24527);
nor UO_844 (O_844,N_24607,N_24618);
xor UO_845 (O_845,N_24525,N_24983);
or UO_846 (O_846,N_24799,N_24837);
nor UO_847 (O_847,N_24873,N_24843);
nor UO_848 (O_848,N_24594,N_24626);
xnor UO_849 (O_849,N_24614,N_24752);
nand UO_850 (O_850,N_24887,N_24974);
and UO_851 (O_851,N_24841,N_24822);
nand UO_852 (O_852,N_24533,N_24763);
nand UO_853 (O_853,N_24987,N_24798);
nor UO_854 (O_854,N_24971,N_24593);
or UO_855 (O_855,N_24750,N_24654);
nor UO_856 (O_856,N_24795,N_24765);
nand UO_857 (O_857,N_24607,N_24876);
nand UO_858 (O_858,N_24711,N_24680);
nand UO_859 (O_859,N_24949,N_24703);
nand UO_860 (O_860,N_24909,N_24563);
and UO_861 (O_861,N_24877,N_24516);
or UO_862 (O_862,N_24529,N_24903);
nand UO_863 (O_863,N_24866,N_24549);
xor UO_864 (O_864,N_24973,N_24904);
nor UO_865 (O_865,N_24554,N_24777);
nor UO_866 (O_866,N_24947,N_24888);
xnor UO_867 (O_867,N_24981,N_24626);
and UO_868 (O_868,N_24762,N_24666);
and UO_869 (O_869,N_24813,N_24866);
nor UO_870 (O_870,N_24518,N_24894);
or UO_871 (O_871,N_24854,N_24950);
and UO_872 (O_872,N_24925,N_24828);
and UO_873 (O_873,N_24680,N_24744);
nor UO_874 (O_874,N_24581,N_24978);
and UO_875 (O_875,N_24844,N_24579);
or UO_876 (O_876,N_24869,N_24720);
xor UO_877 (O_877,N_24874,N_24978);
nand UO_878 (O_878,N_24808,N_24530);
nor UO_879 (O_879,N_24904,N_24513);
xnor UO_880 (O_880,N_24826,N_24616);
xor UO_881 (O_881,N_24843,N_24537);
nand UO_882 (O_882,N_24673,N_24769);
and UO_883 (O_883,N_24856,N_24969);
nand UO_884 (O_884,N_24902,N_24786);
or UO_885 (O_885,N_24953,N_24831);
and UO_886 (O_886,N_24660,N_24509);
and UO_887 (O_887,N_24501,N_24602);
nand UO_888 (O_888,N_24991,N_24737);
nor UO_889 (O_889,N_24822,N_24942);
and UO_890 (O_890,N_24893,N_24688);
and UO_891 (O_891,N_24686,N_24601);
xor UO_892 (O_892,N_24757,N_24556);
and UO_893 (O_893,N_24924,N_24998);
nor UO_894 (O_894,N_24864,N_24771);
xnor UO_895 (O_895,N_24699,N_24827);
nand UO_896 (O_896,N_24576,N_24771);
and UO_897 (O_897,N_24628,N_24975);
nor UO_898 (O_898,N_24855,N_24774);
nand UO_899 (O_899,N_24537,N_24940);
and UO_900 (O_900,N_24958,N_24685);
xor UO_901 (O_901,N_24818,N_24995);
xnor UO_902 (O_902,N_24712,N_24550);
nor UO_903 (O_903,N_24708,N_24590);
nor UO_904 (O_904,N_24554,N_24793);
or UO_905 (O_905,N_24562,N_24924);
and UO_906 (O_906,N_24748,N_24940);
xor UO_907 (O_907,N_24990,N_24959);
or UO_908 (O_908,N_24520,N_24993);
xor UO_909 (O_909,N_24554,N_24744);
nor UO_910 (O_910,N_24519,N_24710);
xnor UO_911 (O_911,N_24708,N_24558);
nor UO_912 (O_912,N_24900,N_24942);
and UO_913 (O_913,N_24635,N_24710);
and UO_914 (O_914,N_24757,N_24571);
xnor UO_915 (O_915,N_24938,N_24565);
nor UO_916 (O_916,N_24600,N_24706);
and UO_917 (O_917,N_24900,N_24909);
nor UO_918 (O_918,N_24999,N_24921);
or UO_919 (O_919,N_24778,N_24960);
nand UO_920 (O_920,N_24663,N_24524);
or UO_921 (O_921,N_24535,N_24858);
nand UO_922 (O_922,N_24727,N_24768);
and UO_923 (O_923,N_24775,N_24832);
and UO_924 (O_924,N_24791,N_24695);
xor UO_925 (O_925,N_24996,N_24523);
xnor UO_926 (O_926,N_24999,N_24577);
xor UO_927 (O_927,N_24951,N_24566);
nor UO_928 (O_928,N_24581,N_24612);
nor UO_929 (O_929,N_24987,N_24745);
and UO_930 (O_930,N_24584,N_24870);
and UO_931 (O_931,N_24944,N_24774);
nor UO_932 (O_932,N_24925,N_24595);
or UO_933 (O_933,N_24611,N_24604);
or UO_934 (O_934,N_24957,N_24715);
or UO_935 (O_935,N_24700,N_24666);
xor UO_936 (O_936,N_24826,N_24793);
nor UO_937 (O_937,N_24947,N_24546);
xnor UO_938 (O_938,N_24839,N_24646);
or UO_939 (O_939,N_24788,N_24971);
nor UO_940 (O_940,N_24876,N_24828);
nand UO_941 (O_941,N_24509,N_24955);
and UO_942 (O_942,N_24739,N_24902);
nand UO_943 (O_943,N_24530,N_24782);
xnor UO_944 (O_944,N_24823,N_24575);
xor UO_945 (O_945,N_24605,N_24689);
nand UO_946 (O_946,N_24749,N_24971);
nor UO_947 (O_947,N_24816,N_24535);
nand UO_948 (O_948,N_24582,N_24954);
xor UO_949 (O_949,N_24824,N_24740);
nor UO_950 (O_950,N_24933,N_24644);
or UO_951 (O_951,N_24892,N_24629);
or UO_952 (O_952,N_24779,N_24556);
nand UO_953 (O_953,N_24579,N_24935);
or UO_954 (O_954,N_24888,N_24936);
nand UO_955 (O_955,N_24947,N_24904);
nor UO_956 (O_956,N_24755,N_24991);
nand UO_957 (O_957,N_24820,N_24943);
nor UO_958 (O_958,N_24790,N_24905);
nand UO_959 (O_959,N_24997,N_24717);
nand UO_960 (O_960,N_24879,N_24645);
or UO_961 (O_961,N_24539,N_24986);
or UO_962 (O_962,N_24567,N_24920);
nor UO_963 (O_963,N_24681,N_24662);
xor UO_964 (O_964,N_24730,N_24850);
or UO_965 (O_965,N_24510,N_24692);
nor UO_966 (O_966,N_24534,N_24700);
and UO_967 (O_967,N_24714,N_24841);
nor UO_968 (O_968,N_24924,N_24523);
and UO_969 (O_969,N_24778,N_24737);
xor UO_970 (O_970,N_24621,N_24769);
and UO_971 (O_971,N_24605,N_24601);
and UO_972 (O_972,N_24875,N_24810);
or UO_973 (O_973,N_24626,N_24790);
nor UO_974 (O_974,N_24698,N_24947);
or UO_975 (O_975,N_24534,N_24915);
nor UO_976 (O_976,N_24628,N_24889);
xnor UO_977 (O_977,N_24560,N_24839);
or UO_978 (O_978,N_24735,N_24992);
and UO_979 (O_979,N_24612,N_24992);
or UO_980 (O_980,N_24898,N_24937);
nor UO_981 (O_981,N_24634,N_24559);
nor UO_982 (O_982,N_24905,N_24574);
or UO_983 (O_983,N_24740,N_24867);
nor UO_984 (O_984,N_24860,N_24677);
and UO_985 (O_985,N_24569,N_24669);
nand UO_986 (O_986,N_24757,N_24590);
nor UO_987 (O_987,N_24544,N_24598);
nand UO_988 (O_988,N_24602,N_24926);
nand UO_989 (O_989,N_24954,N_24677);
xor UO_990 (O_990,N_24767,N_24996);
xor UO_991 (O_991,N_24995,N_24846);
nand UO_992 (O_992,N_24556,N_24789);
xnor UO_993 (O_993,N_24600,N_24713);
xor UO_994 (O_994,N_24568,N_24611);
nand UO_995 (O_995,N_24879,N_24833);
nand UO_996 (O_996,N_24683,N_24621);
or UO_997 (O_997,N_24877,N_24821);
or UO_998 (O_998,N_24657,N_24541);
or UO_999 (O_999,N_24845,N_24765);
or UO_1000 (O_1000,N_24863,N_24576);
nor UO_1001 (O_1001,N_24616,N_24801);
and UO_1002 (O_1002,N_24816,N_24586);
and UO_1003 (O_1003,N_24609,N_24821);
xor UO_1004 (O_1004,N_24969,N_24511);
nor UO_1005 (O_1005,N_24722,N_24978);
nand UO_1006 (O_1006,N_24846,N_24948);
nor UO_1007 (O_1007,N_24507,N_24763);
nand UO_1008 (O_1008,N_24570,N_24977);
xnor UO_1009 (O_1009,N_24750,N_24849);
or UO_1010 (O_1010,N_24655,N_24961);
xor UO_1011 (O_1011,N_24995,N_24998);
and UO_1012 (O_1012,N_24618,N_24664);
nor UO_1013 (O_1013,N_24627,N_24978);
xnor UO_1014 (O_1014,N_24660,N_24679);
nand UO_1015 (O_1015,N_24600,N_24762);
or UO_1016 (O_1016,N_24590,N_24614);
nand UO_1017 (O_1017,N_24668,N_24689);
or UO_1018 (O_1018,N_24726,N_24773);
and UO_1019 (O_1019,N_24965,N_24512);
nand UO_1020 (O_1020,N_24519,N_24814);
nand UO_1021 (O_1021,N_24593,N_24657);
xnor UO_1022 (O_1022,N_24686,N_24912);
xnor UO_1023 (O_1023,N_24778,N_24961);
nand UO_1024 (O_1024,N_24781,N_24843);
and UO_1025 (O_1025,N_24649,N_24749);
or UO_1026 (O_1026,N_24944,N_24758);
nor UO_1027 (O_1027,N_24702,N_24888);
xnor UO_1028 (O_1028,N_24911,N_24530);
and UO_1029 (O_1029,N_24792,N_24923);
nand UO_1030 (O_1030,N_24591,N_24805);
and UO_1031 (O_1031,N_24625,N_24712);
and UO_1032 (O_1032,N_24954,N_24587);
nor UO_1033 (O_1033,N_24999,N_24730);
xor UO_1034 (O_1034,N_24515,N_24527);
nor UO_1035 (O_1035,N_24506,N_24800);
or UO_1036 (O_1036,N_24790,N_24895);
nor UO_1037 (O_1037,N_24745,N_24881);
and UO_1038 (O_1038,N_24880,N_24997);
nand UO_1039 (O_1039,N_24590,N_24557);
nor UO_1040 (O_1040,N_24688,N_24600);
or UO_1041 (O_1041,N_24538,N_24730);
or UO_1042 (O_1042,N_24784,N_24552);
nand UO_1043 (O_1043,N_24987,N_24634);
and UO_1044 (O_1044,N_24729,N_24586);
or UO_1045 (O_1045,N_24620,N_24930);
and UO_1046 (O_1046,N_24779,N_24669);
nand UO_1047 (O_1047,N_24570,N_24550);
nand UO_1048 (O_1048,N_24679,N_24634);
xor UO_1049 (O_1049,N_24542,N_24779);
or UO_1050 (O_1050,N_24886,N_24553);
and UO_1051 (O_1051,N_24578,N_24714);
and UO_1052 (O_1052,N_24802,N_24840);
xnor UO_1053 (O_1053,N_24518,N_24874);
xnor UO_1054 (O_1054,N_24510,N_24775);
nor UO_1055 (O_1055,N_24667,N_24770);
or UO_1056 (O_1056,N_24505,N_24789);
nor UO_1057 (O_1057,N_24766,N_24984);
xnor UO_1058 (O_1058,N_24864,N_24594);
xor UO_1059 (O_1059,N_24635,N_24982);
and UO_1060 (O_1060,N_24509,N_24682);
nor UO_1061 (O_1061,N_24840,N_24739);
or UO_1062 (O_1062,N_24611,N_24760);
xnor UO_1063 (O_1063,N_24951,N_24751);
and UO_1064 (O_1064,N_24949,N_24724);
xor UO_1065 (O_1065,N_24822,N_24760);
and UO_1066 (O_1066,N_24895,N_24893);
xnor UO_1067 (O_1067,N_24969,N_24794);
and UO_1068 (O_1068,N_24848,N_24909);
nor UO_1069 (O_1069,N_24710,N_24814);
nand UO_1070 (O_1070,N_24593,N_24828);
nand UO_1071 (O_1071,N_24620,N_24544);
nor UO_1072 (O_1072,N_24794,N_24546);
or UO_1073 (O_1073,N_24527,N_24697);
and UO_1074 (O_1074,N_24652,N_24583);
nand UO_1075 (O_1075,N_24679,N_24565);
or UO_1076 (O_1076,N_24752,N_24712);
nand UO_1077 (O_1077,N_24860,N_24847);
xnor UO_1078 (O_1078,N_24947,N_24545);
nand UO_1079 (O_1079,N_24865,N_24588);
xor UO_1080 (O_1080,N_24921,N_24804);
xor UO_1081 (O_1081,N_24870,N_24917);
or UO_1082 (O_1082,N_24788,N_24774);
nor UO_1083 (O_1083,N_24589,N_24690);
nor UO_1084 (O_1084,N_24761,N_24943);
xnor UO_1085 (O_1085,N_24893,N_24781);
nor UO_1086 (O_1086,N_24576,N_24521);
nand UO_1087 (O_1087,N_24799,N_24696);
xor UO_1088 (O_1088,N_24562,N_24828);
nor UO_1089 (O_1089,N_24840,N_24936);
nor UO_1090 (O_1090,N_24634,N_24577);
nor UO_1091 (O_1091,N_24534,N_24547);
nand UO_1092 (O_1092,N_24829,N_24508);
and UO_1093 (O_1093,N_24989,N_24974);
nand UO_1094 (O_1094,N_24971,N_24568);
and UO_1095 (O_1095,N_24598,N_24922);
and UO_1096 (O_1096,N_24956,N_24649);
nand UO_1097 (O_1097,N_24893,N_24535);
nand UO_1098 (O_1098,N_24876,N_24979);
nand UO_1099 (O_1099,N_24856,N_24536);
nand UO_1100 (O_1100,N_24851,N_24626);
nand UO_1101 (O_1101,N_24831,N_24511);
xnor UO_1102 (O_1102,N_24846,N_24638);
and UO_1103 (O_1103,N_24892,N_24997);
or UO_1104 (O_1104,N_24999,N_24909);
and UO_1105 (O_1105,N_24708,N_24835);
nor UO_1106 (O_1106,N_24840,N_24683);
nand UO_1107 (O_1107,N_24929,N_24725);
or UO_1108 (O_1108,N_24848,N_24986);
nor UO_1109 (O_1109,N_24801,N_24601);
xor UO_1110 (O_1110,N_24887,N_24602);
nand UO_1111 (O_1111,N_24779,N_24624);
and UO_1112 (O_1112,N_24562,N_24716);
nand UO_1113 (O_1113,N_24506,N_24736);
and UO_1114 (O_1114,N_24860,N_24672);
or UO_1115 (O_1115,N_24608,N_24843);
nand UO_1116 (O_1116,N_24868,N_24947);
xor UO_1117 (O_1117,N_24564,N_24588);
or UO_1118 (O_1118,N_24512,N_24595);
xnor UO_1119 (O_1119,N_24613,N_24743);
and UO_1120 (O_1120,N_24957,N_24656);
nor UO_1121 (O_1121,N_24654,N_24863);
nand UO_1122 (O_1122,N_24879,N_24685);
xnor UO_1123 (O_1123,N_24714,N_24601);
nor UO_1124 (O_1124,N_24563,N_24799);
and UO_1125 (O_1125,N_24931,N_24890);
nor UO_1126 (O_1126,N_24685,N_24552);
and UO_1127 (O_1127,N_24740,N_24900);
nand UO_1128 (O_1128,N_24852,N_24901);
or UO_1129 (O_1129,N_24874,N_24653);
nand UO_1130 (O_1130,N_24527,N_24884);
or UO_1131 (O_1131,N_24946,N_24857);
nand UO_1132 (O_1132,N_24656,N_24797);
nor UO_1133 (O_1133,N_24682,N_24730);
nor UO_1134 (O_1134,N_24813,N_24534);
or UO_1135 (O_1135,N_24679,N_24881);
nand UO_1136 (O_1136,N_24891,N_24722);
and UO_1137 (O_1137,N_24839,N_24605);
nand UO_1138 (O_1138,N_24810,N_24832);
nand UO_1139 (O_1139,N_24806,N_24810);
or UO_1140 (O_1140,N_24702,N_24920);
and UO_1141 (O_1141,N_24709,N_24967);
or UO_1142 (O_1142,N_24779,N_24808);
xnor UO_1143 (O_1143,N_24775,N_24642);
and UO_1144 (O_1144,N_24569,N_24956);
xnor UO_1145 (O_1145,N_24857,N_24659);
nor UO_1146 (O_1146,N_24601,N_24908);
or UO_1147 (O_1147,N_24630,N_24811);
nor UO_1148 (O_1148,N_24640,N_24767);
xor UO_1149 (O_1149,N_24725,N_24722);
xnor UO_1150 (O_1150,N_24557,N_24986);
and UO_1151 (O_1151,N_24650,N_24690);
and UO_1152 (O_1152,N_24759,N_24626);
xor UO_1153 (O_1153,N_24708,N_24532);
nor UO_1154 (O_1154,N_24868,N_24519);
and UO_1155 (O_1155,N_24934,N_24657);
xnor UO_1156 (O_1156,N_24536,N_24889);
xnor UO_1157 (O_1157,N_24815,N_24851);
and UO_1158 (O_1158,N_24645,N_24681);
xnor UO_1159 (O_1159,N_24823,N_24503);
and UO_1160 (O_1160,N_24691,N_24766);
nor UO_1161 (O_1161,N_24641,N_24614);
xnor UO_1162 (O_1162,N_24718,N_24599);
or UO_1163 (O_1163,N_24702,N_24865);
or UO_1164 (O_1164,N_24608,N_24787);
nor UO_1165 (O_1165,N_24846,N_24801);
nand UO_1166 (O_1166,N_24933,N_24543);
nor UO_1167 (O_1167,N_24698,N_24883);
and UO_1168 (O_1168,N_24893,N_24836);
nand UO_1169 (O_1169,N_24756,N_24998);
and UO_1170 (O_1170,N_24822,N_24812);
nand UO_1171 (O_1171,N_24621,N_24674);
or UO_1172 (O_1172,N_24725,N_24568);
or UO_1173 (O_1173,N_24580,N_24525);
nor UO_1174 (O_1174,N_24987,N_24584);
xnor UO_1175 (O_1175,N_24963,N_24623);
or UO_1176 (O_1176,N_24840,N_24766);
nor UO_1177 (O_1177,N_24915,N_24548);
nor UO_1178 (O_1178,N_24631,N_24958);
nand UO_1179 (O_1179,N_24594,N_24789);
xnor UO_1180 (O_1180,N_24795,N_24554);
nor UO_1181 (O_1181,N_24625,N_24520);
xnor UO_1182 (O_1182,N_24886,N_24787);
and UO_1183 (O_1183,N_24899,N_24756);
xor UO_1184 (O_1184,N_24987,N_24521);
nand UO_1185 (O_1185,N_24699,N_24738);
xor UO_1186 (O_1186,N_24529,N_24546);
nor UO_1187 (O_1187,N_24788,N_24683);
xnor UO_1188 (O_1188,N_24984,N_24999);
or UO_1189 (O_1189,N_24768,N_24515);
xor UO_1190 (O_1190,N_24563,N_24586);
and UO_1191 (O_1191,N_24565,N_24744);
nor UO_1192 (O_1192,N_24975,N_24997);
or UO_1193 (O_1193,N_24883,N_24933);
and UO_1194 (O_1194,N_24898,N_24689);
xnor UO_1195 (O_1195,N_24936,N_24809);
and UO_1196 (O_1196,N_24635,N_24834);
nor UO_1197 (O_1197,N_24698,N_24912);
and UO_1198 (O_1198,N_24969,N_24970);
and UO_1199 (O_1199,N_24991,N_24919);
nand UO_1200 (O_1200,N_24886,N_24663);
nor UO_1201 (O_1201,N_24742,N_24835);
nor UO_1202 (O_1202,N_24679,N_24813);
or UO_1203 (O_1203,N_24838,N_24607);
or UO_1204 (O_1204,N_24645,N_24744);
or UO_1205 (O_1205,N_24959,N_24527);
xor UO_1206 (O_1206,N_24532,N_24868);
xor UO_1207 (O_1207,N_24807,N_24722);
xnor UO_1208 (O_1208,N_24746,N_24621);
xnor UO_1209 (O_1209,N_24736,N_24524);
or UO_1210 (O_1210,N_24962,N_24669);
xor UO_1211 (O_1211,N_24850,N_24635);
nand UO_1212 (O_1212,N_24752,N_24606);
nor UO_1213 (O_1213,N_24594,N_24869);
and UO_1214 (O_1214,N_24772,N_24919);
xnor UO_1215 (O_1215,N_24602,N_24531);
or UO_1216 (O_1216,N_24807,N_24918);
nand UO_1217 (O_1217,N_24813,N_24530);
and UO_1218 (O_1218,N_24504,N_24971);
and UO_1219 (O_1219,N_24784,N_24517);
or UO_1220 (O_1220,N_24506,N_24891);
xnor UO_1221 (O_1221,N_24862,N_24568);
nand UO_1222 (O_1222,N_24608,N_24812);
or UO_1223 (O_1223,N_24752,N_24790);
nor UO_1224 (O_1224,N_24661,N_24695);
nor UO_1225 (O_1225,N_24863,N_24806);
and UO_1226 (O_1226,N_24889,N_24820);
nand UO_1227 (O_1227,N_24959,N_24900);
nand UO_1228 (O_1228,N_24779,N_24678);
and UO_1229 (O_1229,N_24754,N_24514);
or UO_1230 (O_1230,N_24847,N_24541);
and UO_1231 (O_1231,N_24683,N_24637);
and UO_1232 (O_1232,N_24970,N_24921);
and UO_1233 (O_1233,N_24749,N_24785);
xor UO_1234 (O_1234,N_24725,N_24553);
xor UO_1235 (O_1235,N_24705,N_24991);
xnor UO_1236 (O_1236,N_24865,N_24628);
nor UO_1237 (O_1237,N_24736,N_24983);
nor UO_1238 (O_1238,N_24513,N_24773);
nor UO_1239 (O_1239,N_24909,N_24755);
nor UO_1240 (O_1240,N_24587,N_24925);
or UO_1241 (O_1241,N_24716,N_24807);
xor UO_1242 (O_1242,N_24931,N_24827);
nor UO_1243 (O_1243,N_24577,N_24696);
or UO_1244 (O_1244,N_24807,N_24720);
xnor UO_1245 (O_1245,N_24592,N_24885);
nor UO_1246 (O_1246,N_24849,N_24881);
xor UO_1247 (O_1247,N_24787,N_24828);
nand UO_1248 (O_1248,N_24600,N_24916);
xnor UO_1249 (O_1249,N_24710,N_24782);
or UO_1250 (O_1250,N_24816,N_24677);
xor UO_1251 (O_1251,N_24598,N_24892);
xor UO_1252 (O_1252,N_24618,N_24632);
nor UO_1253 (O_1253,N_24610,N_24622);
nor UO_1254 (O_1254,N_24695,N_24592);
nand UO_1255 (O_1255,N_24832,N_24527);
and UO_1256 (O_1256,N_24789,N_24969);
nor UO_1257 (O_1257,N_24544,N_24794);
or UO_1258 (O_1258,N_24915,N_24993);
xnor UO_1259 (O_1259,N_24858,N_24722);
and UO_1260 (O_1260,N_24508,N_24959);
xnor UO_1261 (O_1261,N_24850,N_24802);
or UO_1262 (O_1262,N_24804,N_24785);
or UO_1263 (O_1263,N_24815,N_24708);
xor UO_1264 (O_1264,N_24807,N_24986);
xor UO_1265 (O_1265,N_24528,N_24815);
xnor UO_1266 (O_1266,N_24969,N_24871);
xor UO_1267 (O_1267,N_24694,N_24707);
xor UO_1268 (O_1268,N_24892,N_24748);
xor UO_1269 (O_1269,N_24799,N_24652);
xnor UO_1270 (O_1270,N_24511,N_24665);
nor UO_1271 (O_1271,N_24794,N_24589);
or UO_1272 (O_1272,N_24854,N_24536);
nor UO_1273 (O_1273,N_24683,N_24777);
xor UO_1274 (O_1274,N_24655,N_24814);
xor UO_1275 (O_1275,N_24680,N_24926);
nand UO_1276 (O_1276,N_24588,N_24662);
and UO_1277 (O_1277,N_24649,N_24529);
xor UO_1278 (O_1278,N_24704,N_24870);
and UO_1279 (O_1279,N_24822,N_24921);
nand UO_1280 (O_1280,N_24505,N_24746);
and UO_1281 (O_1281,N_24818,N_24508);
xor UO_1282 (O_1282,N_24684,N_24506);
and UO_1283 (O_1283,N_24895,N_24997);
or UO_1284 (O_1284,N_24944,N_24534);
nor UO_1285 (O_1285,N_24753,N_24949);
xor UO_1286 (O_1286,N_24964,N_24642);
xor UO_1287 (O_1287,N_24696,N_24657);
or UO_1288 (O_1288,N_24805,N_24792);
xor UO_1289 (O_1289,N_24804,N_24979);
nor UO_1290 (O_1290,N_24536,N_24838);
nand UO_1291 (O_1291,N_24838,N_24598);
nor UO_1292 (O_1292,N_24592,N_24857);
xor UO_1293 (O_1293,N_24640,N_24604);
and UO_1294 (O_1294,N_24962,N_24771);
xnor UO_1295 (O_1295,N_24618,N_24645);
xnor UO_1296 (O_1296,N_24832,N_24787);
xor UO_1297 (O_1297,N_24504,N_24774);
nand UO_1298 (O_1298,N_24540,N_24566);
nor UO_1299 (O_1299,N_24720,N_24568);
xnor UO_1300 (O_1300,N_24967,N_24870);
nor UO_1301 (O_1301,N_24984,N_24507);
or UO_1302 (O_1302,N_24571,N_24572);
xnor UO_1303 (O_1303,N_24584,N_24757);
nand UO_1304 (O_1304,N_24537,N_24953);
nand UO_1305 (O_1305,N_24908,N_24845);
nor UO_1306 (O_1306,N_24812,N_24520);
or UO_1307 (O_1307,N_24579,N_24621);
and UO_1308 (O_1308,N_24863,N_24773);
nand UO_1309 (O_1309,N_24834,N_24848);
xnor UO_1310 (O_1310,N_24529,N_24739);
xor UO_1311 (O_1311,N_24891,N_24563);
or UO_1312 (O_1312,N_24503,N_24781);
nand UO_1313 (O_1313,N_24520,N_24969);
and UO_1314 (O_1314,N_24630,N_24896);
nor UO_1315 (O_1315,N_24563,N_24626);
nor UO_1316 (O_1316,N_24561,N_24870);
or UO_1317 (O_1317,N_24733,N_24769);
or UO_1318 (O_1318,N_24719,N_24668);
nor UO_1319 (O_1319,N_24840,N_24693);
nor UO_1320 (O_1320,N_24971,N_24958);
nor UO_1321 (O_1321,N_24769,N_24884);
nand UO_1322 (O_1322,N_24962,N_24955);
xnor UO_1323 (O_1323,N_24624,N_24738);
nor UO_1324 (O_1324,N_24768,N_24924);
or UO_1325 (O_1325,N_24868,N_24508);
and UO_1326 (O_1326,N_24687,N_24780);
or UO_1327 (O_1327,N_24695,N_24901);
xnor UO_1328 (O_1328,N_24777,N_24690);
or UO_1329 (O_1329,N_24598,N_24937);
or UO_1330 (O_1330,N_24517,N_24524);
xnor UO_1331 (O_1331,N_24588,N_24887);
xnor UO_1332 (O_1332,N_24652,N_24738);
nor UO_1333 (O_1333,N_24998,N_24569);
xnor UO_1334 (O_1334,N_24892,N_24643);
and UO_1335 (O_1335,N_24604,N_24557);
and UO_1336 (O_1336,N_24866,N_24823);
xnor UO_1337 (O_1337,N_24716,N_24717);
nor UO_1338 (O_1338,N_24901,N_24898);
nand UO_1339 (O_1339,N_24640,N_24602);
and UO_1340 (O_1340,N_24759,N_24787);
nor UO_1341 (O_1341,N_24882,N_24722);
or UO_1342 (O_1342,N_24889,N_24802);
nor UO_1343 (O_1343,N_24545,N_24677);
or UO_1344 (O_1344,N_24552,N_24769);
xor UO_1345 (O_1345,N_24643,N_24754);
nand UO_1346 (O_1346,N_24540,N_24535);
or UO_1347 (O_1347,N_24900,N_24592);
xnor UO_1348 (O_1348,N_24703,N_24874);
xor UO_1349 (O_1349,N_24632,N_24986);
and UO_1350 (O_1350,N_24605,N_24663);
nor UO_1351 (O_1351,N_24533,N_24631);
or UO_1352 (O_1352,N_24543,N_24731);
nand UO_1353 (O_1353,N_24770,N_24758);
xnor UO_1354 (O_1354,N_24921,N_24580);
xor UO_1355 (O_1355,N_24627,N_24895);
nand UO_1356 (O_1356,N_24844,N_24548);
or UO_1357 (O_1357,N_24512,N_24573);
xnor UO_1358 (O_1358,N_24513,N_24757);
xnor UO_1359 (O_1359,N_24691,N_24576);
nand UO_1360 (O_1360,N_24589,N_24903);
xnor UO_1361 (O_1361,N_24788,N_24548);
or UO_1362 (O_1362,N_24597,N_24589);
and UO_1363 (O_1363,N_24857,N_24711);
nor UO_1364 (O_1364,N_24844,N_24828);
nor UO_1365 (O_1365,N_24997,N_24934);
or UO_1366 (O_1366,N_24708,N_24888);
nor UO_1367 (O_1367,N_24718,N_24978);
or UO_1368 (O_1368,N_24633,N_24836);
xor UO_1369 (O_1369,N_24913,N_24818);
xor UO_1370 (O_1370,N_24967,N_24972);
nor UO_1371 (O_1371,N_24706,N_24563);
nor UO_1372 (O_1372,N_24615,N_24787);
or UO_1373 (O_1373,N_24955,N_24692);
xnor UO_1374 (O_1374,N_24946,N_24958);
nor UO_1375 (O_1375,N_24857,N_24556);
xnor UO_1376 (O_1376,N_24817,N_24812);
xnor UO_1377 (O_1377,N_24698,N_24545);
nor UO_1378 (O_1378,N_24543,N_24558);
xnor UO_1379 (O_1379,N_24981,N_24861);
nand UO_1380 (O_1380,N_24868,N_24953);
nand UO_1381 (O_1381,N_24858,N_24717);
and UO_1382 (O_1382,N_24640,N_24842);
and UO_1383 (O_1383,N_24551,N_24539);
nor UO_1384 (O_1384,N_24641,N_24554);
nand UO_1385 (O_1385,N_24862,N_24766);
or UO_1386 (O_1386,N_24806,N_24699);
or UO_1387 (O_1387,N_24691,N_24515);
xor UO_1388 (O_1388,N_24646,N_24763);
and UO_1389 (O_1389,N_24774,N_24940);
nand UO_1390 (O_1390,N_24762,N_24707);
xnor UO_1391 (O_1391,N_24770,N_24709);
nor UO_1392 (O_1392,N_24921,N_24846);
or UO_1393 (O_1393,N_24827,N_24702);
xor UO_1394 (O_1394,N_24800,N_24888);
nand UO_1395 (O_1395,N_24709,N_24713);
and UO_1396 (O_1396,N_24655,N_24708);
and UO_1397 (O_1397,N_24548,N_24557);
nor UO_1398 (O_1398,N_24952,N_24745);
nor UO_1399 (O_1399,N_24554,N_24555);
nand UO_1400 (O_1400,N_24515,N_24675);
and UO_1401 (O_1401,N_24861,N_24513);
nand UO_1402 (O_1402,N_24727,N_24757);
and UO_1403 (O_1403,N_24636,N_24645);
nand UO_1404 (O_1404,N_24670,N_24589);
and UO_1405 (O_1405,N_24558,N_24900);
nand UO_1406 (O_1406,N_24761,N_24801);
nor UO_1407 (O_1407,N_24719,N_24867);
nand UO_1408 (O_1408,N_24696,N_24624);
nand UO_1409 (O_1409,N_24913,N_24780);
and UO_1410 (O_1410,N_24969,N_24662);
nor UO_1411 (O_1411,N_24566,N_24600);
or UO_1412 (O_1412,N_24660,N_24744);
nor UO_1413 (O_1413,N_24826,N_24600);
xor UO_1414 (O_1414,N_24783,N_24608);
or UO_1415 (O_1415,N_24626,N_24585);
xnor UO_1416 (O_1416,N_24649,N_24560);
or UO_1417 (O_1417,N_24823,N_24661);
nand UO_1418 (O_1418,N_24941,N_24751);
nor UO_1419 (O_1419,N_24745,N_24526);
and UO_1420 (O_1420,N_24866,N_24553);
xor UO_1421 (O_1421,N_24690,N_24535);
nor UO_1422 (O_1422,N_24713,N_24697);
xor UO_1423 (O_1423,N_24931,N_24515);
nor UO_1424 (O_1424,N_24709,N_24646);
and UO_1425 (O_1425,N_24692,N_24682);
and UO_1426 (O_1426,N_24600,N_24730);
nand UO_1427 (O_1427,N_24741,N_24844);
or UO_1428 (O_1428,N_24896,N_24612);
xor UO_1429 (O_1429,N_24575,N_24620);
and UO_1430 (O_1430,N_24893,N_24595);
nor UO_1431 (O_1431,N_24638,N_24909);
and UO_1432 (O_1432,N_24849,N_24742);
and UO_1433 (O_1433,N_24513,N_24849);
and UO_1434 (O_1434,N_24605,N_24742);
nor UO_1435 (O_1435,N_24568,N_24834);
and UO_1436 (O_1436,N_24561,N_24687);
xnor UO_1437 (O_1437,N_24706,N_24952);
nand UO_1438 (O_1438,N_24875,N_24858);
nor UO_1439 (O_1439,N_24674,N_24793);
and UO_1440 (O_1440,N_24561,N_24579);
nor UO_1441 (O_1441,N_24807,N_24684);
nor UO_1442 (O_1442,N_24657,N_24599);
and UO_1443 (O_1443,N_24761,N_24716);
xnor UO_1444 (O_1444,N_24819,N_24861);
and UO_1445 (O_1445,N_24628,N_24946);
or UO_1446 (O_1446,N_24527,N_24755);
and UO_1447 (O_1447,N_24689,N_24558);
or UO_1448 (O_1448,N_24791,N_24521);
xor UO_1449 (O_1449,N_24714,N_24776);
and UO_1450 (O_1450,N_24605,N_24562);
nand UO_1451 (O_1451,N_24520,N_24550);
xor UO_1452 (O_1452,N_24587,N_24516);
xnor UO_1453 (O_1453,N_24647,N_24930);
xor UO_1454 (O_1454,N_24683,N_24503);
xor UO_1455 (O_1455,N_24517,N_24654);
nor UO_1456 (O_1456,N_24803,N_24582);
and UO_1457 (O_1457,N_24528,N_24942);
xor UO_1458 (O_1458,N_24968,N_24712);
nand UO_1459 (O_1459,N_24787,N_24522);
nor UO_1460 (O_1460,N_24848,N_24835);
and UO_1461 (O_1461,N_24773,N_24916);
or UO_1462 (O_1462,N_24873,N_24978);
xnor UO_1463 (O_1463,N_24928,N_24601);
nand UO_1464 (O_1464,N_24837,N_24749);
xor UO_1465 (O_1465,N_24796,N_24857);
nor UO_1466 (O_1466,N_24757,N_24543);
xor UO_1467 (O_1467,N_24973,N_24730);
nand UO_1468 (O_1468,N_24707,N_24537);
and UO_1469 (O_1469,N_24768,N_24635);
nor UO_1470 (O_1470,N_24948,N_24650);
and UO_1471 (O_1471,N_24914,N_24952);
nand UO_1472 (O_1472,N_24869,N_24857);
or UO_1473 (O_1473,N_24697,N_24901);
nor UO_1474 (O_1474,N_24836,N_24637);
or UO_1475 (O_1475,N_24990,N_24788);
or UO_1476 (O_1476,N_24994,N_24672);
xor UO_1477 (O_1477,N_24513,N_24956);
xnor UO_1478 (O_1478,N_24628,N_24858);
nand UO_1479 (O_1479,N_24772,N_24605);
nor UO_1480 (O_1480,N_24781,N_24724);
or UO_1481 (O_1481,N_24853,N_24568);
and UO_1482 (O_1482,N_24557,N_24999);
xor UO_1483 (O_1483,N_24764,N_24868);
and UO_1484 (O_1484,N_24610,N_24935);
nand UO_1485 (O_1485,N_24844,N_24948);
or UO_1486 (O_1486,N_24788,N_24885);
or UO_1487 (O_1487,N_24628,N_24886);
or UO_1488 (O_1488,N_24794,N_24799);
and UO_1489 (O_1489,N_24893,N_24550);
xor UO_1490 (O_1490,N_24760,N_24773);
and UO_1491 (O_1491,N_24626,N_24625);
nand UO_1492 (O_1492,N_24927,N_24729);
xnor UO_1493 (O_1493,N_24540,N_24822);
and UO_1494 (O_1494,N_24526,N_24754);
nor UO_1495 (O_1495,N_24596,N_24549);
or UO_1496 (O_1496,N_24746,N_24693);
nand UO_1497 (O_1497,N_24637,N_24913);
and UO_1498 (O_1498,N_24718,N_24948);
nor UO_1499 (O_1499,N_24507,N_24539);
and UO_1500 (O_1500,N_24682,N_24853);
nor UO_1501 (O_1501,N_24507,N_24512);
nor UO_1502 (O_1502,N_24671,N_24590);
nor UO_1503 (O_1503,N_24823,N_24555);
xnor UO_1504 (O_1504,N_24887,N_24763);
nand UO_1505 (O_1505,N_24572,N_24993);
or UO_1506 (O_1506,N_24811,N_24710);
nand UO_1507 (O_1507,N_24910,N_24877);
and UO_1508 (O_1508,N_24869,N_24552);
xnor UO_1509 (O_1509,N_24556,N_24649);
nand UO_1510 (O_1510,N_24880,N_24899);
nor UO_1511 (O_1511,N_24592,N_24950);
or UO_1512 (O_1512,N_24738,N_24895);
nand UO_1513 (O_1513,N_24524,N_24792);
nor UO_1514 (O_1514,N_24963,N_24785);
nand UO_1515 (O_1515,N_24865,N_24679);
xor UO_1516 (O_1516,N_24921,N_24596);
nor UO_1517 (O_1517,N_24843,N_24650);
xor UO_1518 (O_1518,N_24780,N_24858);
nor UO_1519 (O_1519,N_24985,N_24802);
or UO_1520 (O_1520,N_24647,N_24594);
nand UO_1521 (O_1521,N_24837,N_24774);
xnor UO_1522 (O_1522,N_24620,N_24509);
and UO_1523 (O_1523,N_24994,N_24663);
nor UO_1524 (O_1524,N_24623,N_24539);
or UO_1525 (O_1525,N_24840,N_24622);
xnor UO_1526 (O_1526,N_24537,N_24750);
xor UO_1527 (O_1527,N_24691,N_24980);
or UO_1528 (O_1528,N_24640,N_24543);
nor UO_1529 (O_1529,N_24835,N_24943);
or UO_1530 (O_1530,N_24740,N_24817);
and UO_1531 (O_1531,N_24594,N_24565);
xnor UO_1532 (O_1532,N_24508,N_24987);
xnor UO_1533 (O_1533,N_24626,N_24621);
nand UO_1534 (O_1534,N_24832,N_24705);
xor UO_1535 (O_1535,N_24954,N_24746);
nand UO_1536 (O_1536,N_24736,N_24653);
nor UO_1537 (O_1537,N_24519,N_24540);
nor UO_1538 (O_1538,N_24940,N_24942);
xnor UO_1539 (O_1539,N_24982,N_24703);
and UO_1540 (O_1540,N_24847,N_24627);
xnor UO_1541 (O_1541,N_24545,N_24903);
nor UO_1542 (O_1542,N_24797,N_24771);
nor UO_1543 (O_1543,N_24849,N_24829);
nor UO_1544 (O_1544,N_24883,N_24832);
or UO_1545 (O_1545,N_24891,N_24990);
xor UO_1546 (O_1546,N_24728,N_24770);
nand UO_1547 (O_1547,N_24989,N_24558);
nand UO_1548 (O_1548,N_24626,N_24810);
xnor UO_1549 (O_1549,N_24725,N_24825);
nand UO_1550 (O_1550,N_24542,N_24861);
and UO_1551 (O_1551,N_24533,N_24776);
xor UO_1552 (O_1552,N_24621,N_24765);
nand UO_1553 (O_1553,N_24620,N_24770);
nand UO_1554 (O_1554,N_24523,N_24568);
and UO_1555 (O_1555,N_24829,N_24652);
and UO_1556 (O_1556,N_24834,N_24975);
nand UO_1557 (O_1557,N_24522,N_24582);
xor UO_1558 (O_1558,N_24816,N_24919);
and UO_1559 (O_1559,N_24529,N_24755);
nand UO_1560 (O_1560,N_24851,N_24616);
nor UO_1561 (O_1561,N_24751,N_24557);
xor UO_1562 (O_1562,N_24580,N_24941);
and UO_1563 (O_1563,N_24656,N_24790);
or UO_1564 (O_1564,N_24560,N_24983);
and UO_1565 (O_1565,N_24852,N_24810);
nand UO_1566 (O_1566,N_24864,N_24573);
and UO_1567 (O_1567,N_24760,N_24688);
xnor UO_1568 (O_1568,N_24539,N_24575);
xor UO_1569 (O_1569,N_24973,N_24802);
and UO_1570 (O_1570,N_24949,N_24667);
or UO_1571 (O_1571,N_24517,N_24607);
nand UO_1572 (O_1572,N_24672,N_24807);
and UO_1573 (O_1573,N_24662,N_24836);
nand UO_1574 (O_1574,N_24951,N_24732);
and UO_1575 (O_1575,N_24502,N_24730);
nor UO_1576 (O_1576,N_24640,N_24962);
or UO_1577 (O_1577,N_24604,N_24771);
or UO_1578 (O_1578,N_24997,N_24553);
nor UO_1579 (O_1579,N_24911,N_24517);
xor UO_1580 (O_1580,N_24612,N_24558);
xnor UO_1581 (O_1581,N_24917,N_24944);
and UO_1582 (O_1582,N_24877,N_24570);
nor UO_1583 (O_1583,N_24511,N_24784);
or UO_1584 (O_1584,N_24718,N_24704);
nand UO_1585 (O_1585,N_24536,N_24661);
or UO_1586 (O_1586,N_24577,N_24509);
or UO_1587 (O_1587,N_24878,N_24832);
xor UO_1588 (O_1588,N_24868,N_24662);
nand UO_1589 (O_1589,N_24566,N_24955);
or UO_1590 (O_1590,N_24888,N_24884);
xnor UO_1591 (O_1591,N_24643,N_24837);
nor UO_1592 (O_1592,N_24812,N_24882);
xnor UO_1593 (O_1593,N_24530,N_24755);
and UO_1594 (O_1594,N_24750,N_24603);
nand UO_1595 (O_1595,N_24629,N_24895);
xnor UO_1596 (O_1596,N_24515,N_24699);
or UO_1597 (O_1597,N_24580,N_24622);
or UO_1598 (O_1598,N_24830,N_24712);
and UO_1599 (O_1599,N_24741,N_24800);
xor UO_1600 (O_1600,N_24897,N_24626);
or UO_1601 (O_1601,N_24664,N_24838);
and UO_1602 (O_1602,N_24746,N_24762);
xor UO_1603 (O_1603,N_24671,N_24656);
or UO_1604 (O_1604,N_24546,N_24864);
and UO_1605 (O_1605,N_24929,N_24958);
nand UO_1606 (O_1606,N_24526,N_24933);
or UO_1607 (O_1607,N_24829,N_24981);
or UO_1608 (O_1608,N_24744,N_24890);
nand UO_1609 (O_1609,N_24721,N_24886);
or UO_1610 (O_1610,N_24732,N_24842);
nand UO_1611 (O_1611,N_24620,N_24787);
nand UO_1612 (O_1612,N_24576,N_24722);
xnor UO_1613 (O_1613,N_24886,N_24632);
xor UO_1614 (O_1614,N_24651,N_24794);
and UO_1615 (O_1615,N_24734,N_24639);
nand UO_1616 (O_1616,N_24785,N_24918);
nand UO_1617 (O_1617,N_24885,N_24850);
and UO_1618 (O_1618,N_24553,N_24648);
nor UO_1619 (O_1619,N_24562,N_24665);
xor UO_1620 (O_1620,N_24813,N_24642);
xnor UO_1621 (O_1621,N_24956,N_24986);
nor UO_1622 (O_1622,N_24776,N_24845);
nand UO_1623 (O_1623,N_24510,N_24801);
or UO_1624 (O_1624,N_24756,N_24513);
nand UO_1625 (O_1625,N_24719,N_24730);
xor UO_1626 (O_1626,N_24866,N_24620);
nor UO_1627 (O_1627,N_24736,N_24833);
nand UO_1628 (O_1628,N_24724,N_24637);
nor UO_1629 (O_1629,N_24896,N_24740);
nand UO_1630 (O_1630,N_24861,N_24506);
and UO_1631 (O_1631,N_24955,N_24545);
nor UO_1632 (O_1632,N_24572,N_24915);
nand UO_1633 (O_1633,N_24933,N_24764);
nand UO_1634 (O_1634,N_24507,N_24695);
nand UO_1635 (O_1635,N_24812,N_24836);
xor UO_1636 (O_1636,N_24825,N_24767);
nor UO_1637 (O_1637,N_24575,N_24995);
xor UO_1638 (O_1638,N_24813,N_24747);
and UO_1639 (O_1639,N_24876,N_24676);
nor UO_1640 (O_1640,N_24940,N_24639);
nor UO_1641 (O_1641,N_24924,N_24503);
or UO_1642 (O_1642,N_24765,N_24585);
nand UO_1643 (O_1643,N_24965,N_24878);
nand UO_1644 (O_1644,N_24892,N_24960);
nor UO_1645 (O_1645,N_24910,N_24714);
nand UO_1646 (O_1646,N_24851,N_24596);
and UO_1647 (O_1647,N_24897,N_24551);
nand UO_1648 (O_1648,N_24646,N_24800);
or UO_1649 (O_1649,N_24673,N_24773);
nand UO_1650 (O_1650,N_24928,N_24904);
and UO_1651 (O_1651,N_24619,N_24513);
nand UO_1652 (O_1652,N_24734,N_24836);
or UO_1653 (O_1653,N_24625,N_24817);
or UO_1654 (O_1654,N_24562,N_24531);
or UO_1655 (O_1655,N_24893,N_24693);
and UO_1656 (O_1656,N_24822,N_24551);
and UO_1657 (O_1657,N_24763,N_24844);
or UO_1658 (O_1658,N_24559,N_24841);
nand UO_1659 (O_1659,N_24538,N_24854);
xor UO_1660 (O_1660,N_24977,N_24839);
nor UO_1661 (O_1661,N_24885,N_24835);
and UO_1662 (O_1662,N_24502,N_24798);
nand UO_1663 (O_1663,N_24681,N_24526);
and UO_1664 (O_1664,N_24815,N_24542);
nor UO_1665 (O_1665,N_24661,N_24913);
nor UO_1666 (O_1666,N_24824,N_24592);
nand UO_1667 (O_1667,N_24924,N_24796);
nand UO_1668 (O_1668,N_24621,N_24979);
or UO_1669 (O_1669,N_24735,N_24889);
and UO_1670 (O_1670,N_24810,N_24703);
and UO_1671 (O_1671,N_24939,N_24775);
or UO_1672 (O_1672,N_24733,N_24537);
or UO_1673 (O_1673,N_24790,N_24662);
xor UO_1674 (O_1674,N_24765,N_24548);
or UO_1675 (O_1675,N_24860,N_24924);
nand UO_1676 (O_1676,N_24776,N_24564);
nand UO_1677 (O_1677,N_24778,N_24504);
nor UO_1678 (O_1678,N_24564,N_24996);
nor UO_1679 (O_1679,N_24519,N_24615);
and UO_1680 (O_1680,N_24697,N_24597);
nand UO_1681 (O_1681,N_24614,N_24864);
nand UO_1682 (O_1682,N_24968,N_24508);
and UO_1683 (O_1683,N_24504,N_24743);
xnor UO_1684 (O_1684,N_24640,N_24880);
and UO_1685 (O_1685,N_24552,N_24985);
xnor UO_1686 (O_1686,N_24758,N_24607);
nand UO_1687 (O_1687,N_24922,N_24556);
nor UO_1688 (O_1688,N_24533,N_24868);
and UO_1689 (O_1689,N_24992,N_24548);
or UO_1690 (O_1690,N_24596,N_24691);
nor UO_1691 (O_1691,N_24930,N_24871);
nor UO_1692 (O_1692,N_24769,N_24610);
xor UO_1693 (O_1693,N_24897,N_24773);
nand UO_1694 (O_1694,N_24932,N_24604);
nor UO_1695 (O_1695,N_24509,N_24933);
nand UO_1696 (O_1696,N_24931,N_24828);
and UO_1697 (O_1697,N_24531,N_24898);
and UO_1698 (O_1698,N_24751,N_24616);
nor UO_1699 (O_1699,N_24920,N_24555);
and UO_1700 (O_1700,N_24824,N_24904);
xnor UO_1701 (O_1701,N_24835,N_24886);
or UO_1702 (O_1702,N_24698,N_24758);
nor UO_1703 (O_1703,N_24928,N_24679);
xnor UO_1704 (O_1704,N_24815,N_24573);
and UO_1705 (O_1705,N_24669,N_24837);
or UO_1706 (O_1706,N_24997,N_24660);
xor UO_1707 (O_1707,N_24947,N_24567);
or UO_1708 (O_1708,N_24742,N_24950);
nand UO_1709 (O_1709,N_24536,N_24999);
nand UO_1710 (O_1710,N_24842,N_24896);
nor UO_1711 (O_1711,N_24945,N_24579);
nand UO_1712 (O_1712,N_24543,N_24748);
nand UO_1713 (O_1713,N_24759,N_24637);
xnor UO_1714 (O_1714,N_24726,N_24985);
nand UO_1715 (O_1715,N_24612,N_24814);
nand UO_1716 (O_1716,N_24663,N_24863);
nand UO_1717 (O_1717,N_24607,N_24637);
nor UO_1718 (O_1718,N_24626,N_24738);
xnor UO_1719 (O_1719,N_24766,N_24565);
xor UO_1720 (O_1720,N_24789,N_24743);
or UO_1721 (O_1721,N_24639,N_24674);
nor UO_1722 (O_1722,N_24505,N_24915);
or UO_1723 (O_1723,N_24962,N_24847);
nand UO_1724 (O_1724,N_24554,N_24539);
and UO_1725 (O_1725,N_24515,N_24850);
or UO_1726 (O_1726,N_24700,N_24644);
xor UO_1727 (O_1727,N_24795,N_24630);
xnor UO_1728 (O_1728,N_24786,N_24951);
or UO_1729 (O_1729,N_24874,N_24841);
or UO_1730 (O_1730,N_24796,N_24717);
xor UO_1731 (O_1731,N_24997,N_24937);
or UO_1732 (O_1732,N_24871,N_24862);
xnor UO_1733 (O_1733,N_24710,N_24897);
or UO_1734 (O_1734,N_24556,N_24537);
xnor UO_1735 (O_1735,N_24578,N_24838);
nand UO_1736 (O_1736,N_24776,N_24511);
xnor UO_1737 (O_1737,N_24765,N_24528);
nand UO_1738 (O_1738,N_24892,N_24770);
or UO_1739 (O_1739,N_24680,N_24687);
nor UO_1740 (O_1740,N_24794,N_24698);
nand UO_1741 (O_1741,N_24744,N_24768);
xnor UO_1742 (O_1742,N_24537,N_24586);
nand UO_1743 (O_1743,N_24511,N_24658);
or UO_1744 (O_1744,N_24843,N_24504);
nand UO_1745 (O_1745,N_24986,N_24641);
or UO_1746 (O_1746,N_24836,N_24713);
nand UO_1747 (O_1747,N_24848,N_24619);
xnor UO_1748 (O_1748,N_24723,N_24761);
and UO_1749 (O_1749,N_24611,N_24744);
nand UO_1750 (O_1750,N_24640,N_24516);
nor UO_1751 (O_1751,N_24723,N_24993);
or UO_1752 (O_1752,N_24784,N_24923);
nor UO_1753 (O_1753,N_24792,N_24556);
or UO_1754 (O_1754,N_24500,N_24561);
or UO_1755 (O_1755,N_24880,N_24938);
or UO_1756 (O_1756,N_24927,N_24917);
nor UO_1757 (O_1757,N_24545,N_24525);
and UO_1758 (O_1758,N_24943,N_24699);
nand UO_1759 (O_1759,N_24938,N_24655);
nand UO_1760 (O_1760,N_24946,N_24630);
nand UO_1761 (O_1761,N_24984,N_24555);
xor UO_1762 (O_1762,N_24654,N_24947);
or UO_1763 (O_1763,N_24882,N_24522);
and UO_1764 (O_1764,N_24902,N_24750);
and UO_1765 (O_1765,N_24615,N_24662);
xor UO_1766 (O_1766,N_24622,N_24739);
nand UO_1767 (O_1767,N_24769,N_24705);
nor UO_1768 (O_1768,N_24557,N_24910);
or UO_1769 (O_1769,N_24841,N_24601);
nor UO_1770 (O_1770,N_24948,N_24673);
and UO_1771 (O_1771,N_24730,N_24882);
xor UO_1772 (O_1772,N_24731,N_24692);
or UO_1773 (O_1773,N_24535,N_24581);
and UO_1774 (O_1774,N_24660,N_24984);
xnor UO_1775 (O_1775,N_24781,N_24936);
nor UO_1776 (O_1776,N_24720,N_24620);
or UO_1777 (O_1777,N_24522,N_24995);
xnor UO_1778 (O_1778,N_24800,N_24848);
or UO_1779 (O_1779,N_24764,N_24916);
nor UO_1780 (O_1780,N_24892,N_24609);
and UO_1781 (O_1781,N_24867,N_24602);
or UO_1782 (O_1782,N_24754,N_24958);
xnor UO_1783 (O_1783,N_24863,N_24908);
and UO_1784 (O_1784,N_24924,N_24957);
nor UO_1785 (O_1785,N_24582,N_24746);
and UO_1786 (O_1786,N_24596,N_24642);
or UO_1787 (O_1787,N_24794,N_24797);
xor UO_1788 (O_1788,N_24914,N_24528);
nand UO_1789 (O_1789,N_24846,N_24932);
xor UO_1790 (O_1790,N_24643,N_24770);
xor UO_1791 (O_1791,N_24851,N_24556);
xnor UO_1792 (O_1792,N_24959,N_24998);
nand UO_1793 (O_1793,N_24672,N_24730);
xor UO_1794 (O_1794,N_24977,N_24736);
xnor UO_1795 (O_1795,N_24554,N_24783);
nor UO_1796 (O_1796,N_24786,N_24701);
nand UO_1797 (O_1797,N_24916,N_24808);
and UO_1798 (O_1798,N_24732,N_24959);
and UO_1799 (O_1799,N_24843,N_24878);
nand UO_1800 (O_1800,N_24976,N_24801);
nand UO_1801 (O_1801,N_24904,N_24745);
or UO_1802 (O_1802,N_24540,N_24796);
xor UO_1803 (O_1803,N_24512,N_24738);
and UO_1804 (O_1804,N_24906,N_24636);
and UO_1805 (O_1805,N_24928,N_24817);
nand UO_1806 (O_1806,N_24563,N_24720);
and UO_1807 (O_1807,N_24685,N_24766);
xnor UO_1808 (O_1808,N_24626,N_24668);
nor UO_1809 (O_1809,N_24735,N_24865);
and UO_1810 (O_1810,N_24999,N_24701);
nor UO_1811 (O_1811,N_24762,N_24959);
and UO_1812 (O_1812,N_24958,N_24833);
nor UO_1813 (O_1813,N_24973,N_24553);
nor UO_1814 (O_1814,N_24542,N_24746);
xnor UO_1815 (O_1815,N_24628,N_24667);
nor UO_1816 (O_1816,N_24942,N_24980);
and UO_1817 (O_1817,N_24582,N_24715);
or UO_1818 (O_1818,N_24965,N_24652);
nand UO_1819 (O_1819,N_24961,N_24982);
nand UO_1820 (O_1820,N_24566,N_24555);
nand UO_1821 (O_1821,N_24744,N_24770);
xnor UO_1822 (O_1822,N_24596,N_24703);
xor UO_1823 (O_1823,N_24827,N_24771);
and UO_1824 (O_1824,N_24841,N_24670);
nand UO_1825 (O_1825,N_24957,N_24798);
or UO_1826 (O_1826,N_24562,N_24632);
nor UO_1827 (O_1827,N_24829,N_24546);
or UO_1828 (O_1828,N_24757,N_24944);
nor UO_1829 (O_1829,N_24931,N_24875);
and UO_1830 (O_1830,N_24935,N_24944);
or UO_1831 (O_1831,N_24659,N_24842);
or UO_1832 (O_1832,N_24922,N_24883);
and UO_1833 (O_1833,N_24562,N_24705);
and UO_1834 (O_1834,N_24671,N_24774);
nand UO_1835 (O_1835,N_24918,N_24989);
xnor UO_1836 (O_1836,N_24972,N_24501);
xor UO_1837 (O_1837,N_24725,N_24562);
nand UO_1838 (O_1838,N_24785,N_24675);
or UO_1839 (O_1839,N_24944,N_24546);
nor UO_1840 (O_1840,N_24941,N_24513);
nor UO_1841 (O_1841,N_24934,N_24724);
nor UO_1842 (O_1842,N_24963,N_24910);
xnor UO_1843 (O_1843,N_24549,N_24542);
nor UO_1844 (O_1844,N_24639,N_24871);
or UO_1845 (O_1845,N_24880,N_24972);
nand UO_1846 (O_1846,N_24656,N_24628);
nand UO_1847 (O_1847,N_24907,N_24577);
nand UO_1848 (O_1848,N_24586,N_24517);
xnor UO_1849 (O_1849,N_24893,N_24683);
and UO_1850 (O_1850,N_24797,N_24983);
nor UO_1851 (O_1851,N_24627,N_24675);
and UO_1852 (O_1852,N_24678,N_24590);
nand UO_1853 (O_1853,N_24590,N_24582);
and UO_1854 (O_1854,N_24609,N_24843);
nand UO_1855 (O_1855,N_24657,N_24505);
and UO_1856 (O_1856,N_24828,N_24771);
or UO_1857 (O_1857,N_24591,N_24653);
or UO_1858 (O_1858,N_24985,N_24509);
and UO_1859 (O_1859,N_24956,N_24548);
or UO_1860 (O_1860,N_24772,N_24923);
nor UO_1861 (O_1861,N_24790,N_24638);
xor UO_1862 (O_1862,N_24610,N_24754);
or UO_1863 (O_1863,N_24960,N_24796);
or UO_1864 (O_1864,N_24607,N_24992);
and UO_1865 (O_1865,N_24947,N_24777);
or UO_1866 (O_1866,N_24795,N_24875);
nand UO_1867 (O_1867,N_24973,N_24646);
or UO_1868 (O_1868,N_24610,N_24992);
nand UO_1869 (O_1869,N_24585,N_24839);
and UO_1870 (O_1870,N_24996,N_24569);
xor UO_1871 (O_1871,N_24585,N_24893);
nand UO_1872 (O_1872,N_24985,N_24740);
and UO_1873 (O_1873,N_24869,N_24884);
xnor UO_1874 (O_1874,N_24805,N_24550);
xor UO_1875 (O_1875,N_24642,N_24826);
nor UO_1876 (O_1876,N_24692,N_24734);
or UO_1877 (O_1877,N_24629,N_24852);
nor UO_1878 (O_1878,N_24587,N_24836);
xor UO_1879 (O_1879,N_24967,N_24954);
xor UO_1880 (O_1880,N_24933,N_24557);
nor UO_1881 (O_1881,N_24912,N_24951);
nand UO_1882 (O_1882,N_24653,N_24744);
nor UO_1883 (O_1883,N_24570,N_24997);
or UO_1884 (O_1884,N_24638,N_24837);
nor UO_1885 (O_1885,N_24896,N_24880);
nand UO_1886 (O_1886,N_24972,N_24905);
nand UO_1887 (O_1887,N_24550,N_24639);
or UO_1888 (O_1888,N_24569,N_24859);
or UO_1889 (O_1889,N_24643,N_24730);
nor UO_1890 (O_1890,N_24527,N_24723);
nand UO_1891 (O_1891,N_24897,N_24704);
and UO_1892 (O_1892,N_24733,N_24573);
nand UO_1893 (O_1893,N_24948,N_24533);
and UO_1894 (O_1894,N_24818,N_24638);
nor UO_1895 (O_1895,N_24680,N_24739);
nand UO_1896 (O_1896,N_24762,N_24569);
nor UO_1897 (O_1897,N_24563,N_24929);
or UO_1898 (O_1898,N_24861,N_24593);
nand UO_1899 (O_1899,N_24537,N_24642);
and UO_1900 (O_1900,N_24833,N_24648);
xor UO_1901 (O_1901,N_24541,N_24981);
and UO_1902 (O_1902,N_24951,N_24759);
xnor UO_1903 (O_1903,N_24526,N_24698);
nand UO_1904 (O_1904,N_24709,N_24736);
nand UO_1905 (O_1905,N_24749,N_24713);
xor UO_1906 (O_1906,N_24569,N_24899);
xnor UO_1907 (O_1907,N_24924,N_24572);
nor UO_1908 (O_1908,N_24588,N_24781);
nor UO_1909 (O_1909,N_24801,N_24660);
nor UO_1910 (O_1910,N_24658,N_24795);
and UO_1911 (O_1911,N_24822,N_24630);
xnor UO_1912 (O_1912,N_24931,N_24637);
nor UO_1913 (O_1913,N_24873,N_24717);
xnor UO_1914 (O_1914,N_24892,N_24627);
xor UO_1915 (O_1915,N_24686,N_24782);
nor UO_1916 (O_1916,N_24723,N_24643);
nand UO_1917 (O_1917,N_24834,N_24970);
xnor UO_1918 (O_1918,N_24858,N_24561);
nor UO_1919 (O_1919,N_24847,N_24866);
or UO_1920 (O_1920,N_24965,N_24645);
or UO_1921 (O_1921,N_24722,N_24938);
and UO_1922 (O_1922,N_24961,N_24975);
nor UO_1923 (O_1923,N_24732,N_24977);
and UO_1924 (O_1924,N_24603,N_24772);
or UO_1925 (O_1925,N_24734,N_24822);
or UO_1926 (O_1926,N_24918,N_24951);
and UO_1927 (O_1927,N_24781,N_24658);
nor UO_1928 (O_1928,N_24572,N_24952);
nor UO_1929 (O_1929,N_24651,N_24779);
xnor UO_1930 (O_1930,N_24916,N_24989);
nand UO_1931 (O_1931,N_24837,N_24909);
or UO_1932 (O_1932,N_24851,N_24745);
nor UO_1933 (O_1933,N_24799,N_24685);
and UO_1934 (O_1934,N_24611,N_24514);
nor UO_1935 (O_1935,N_24695,N_24660);
nand UO_1936 (O_1936,N_24541,N_24748);
or UO_1937 (O_1937,N_24704,N_24875);
or UO_1938 (O_1938,N_24839,N_24578);
and UO_1939 (O_1939,N_24715,N_24710);
xor UO_1940 (O_1940,N_24797,N_24845);
xnor UO_1941 (O_1941,N_24936,N_24910);
or UO_1942 (O_1942,N_24677,N_24974);
nand UO_1943 (O_1943,N_24525,N_24548);
nor UO_1944 (O_1944,N_24695,N_24619);
or UO_1945 (O_1945,N_24534,N_24637);
and UO_1946 (O_1946,N_24583,N_24544);
nor UO_1947 (O_1947,N_24751,N_24659);
or UO_1948 (O_1948,N_24521,N_24795);
and UO_1949 (O_1949,N_24710,N_24501);
xnor UO_1950 (O_1950,N_24709,N_24513);
nor UO_1951 (O_1951,N_24931,N_24907);
nand UO_1952 (O_1952,N_24847,N_24824);
nand UO_1953 (O_1953,N_24548,N_24965);
nor UO_1954 (O_1954,N_24746,N_24924);
or UO_1955 (O_1955,N_24551,N_24794);
and UO_1956 (O_1956,N_24807,N_24629);
nand UO_1957 (O_1957,N_24836,N_24938);
or UO_1958 (O_1958,N_24861,N_24749);
or UO_1959 (O_1959,N_24626,N_24832);
nand UO_1960 (O_1960,N_24712,N_24939);
nand UO_1961 (O_1961,N_24934,N_24938);
and UO_1962 (O_1962,N_24691,N_24996);
nor UO_1963 (O_1963,N_24742,N_24733);
nand UO_1964 (O_1964,N_24954,N_24543);
nand UO_1965 (O_1965,N_24511,N_24646);
or UO_1966 (O_1966,N_24918,N_24928);
nor UO_1967 (O_1967,N_24628,N_24992);
xnor UO_1968 (O_1968,N_24656,N_24627);
nor UO_1969 (O_1969,N_24805,N_24946);
xnor UO_1970 (O_1970,N_24765,N_24754);
nand UO_1971 (O_1971,N_24503,N_24916);
nor UO_1972 (O_1972,N_24735,N_24835);
nand UO_1973 (O_1973,N_24757,N_24990);
nor UO_1974 (O_1974,N_24605,N_24818);
and UO_1975 (O_1975,N_24559,N_24809);
and UO_1976 (O_1976,N_24695,N_24927);
nand UO_1977 (O_1977,N_24532,N_24906);
xnor UO_1978 (O_1978,N_24950,N_24816);
or UO_1979 (O_1979,N_24797,N_24697);
xor UO_1980 (O_1980,N_24945,N_24587);
or UO_1981 (O_1981,N_24732,N_24594);
and UO_1982 (O_1982,N_24856,N_24741);
xnor UO_1983 (O_1983,N_24924,N_24829);
and UO_1984 (O_1984,N_24854,N_24900);
or UO_1985 (O_1985,N_24956,N_24941);
nand UO_1986 (O_1986,N_24947,N_24877);
nand UO_1987 (O_1987,N_24659,N_24542);
or UO_1988 (O_1988,N_24880,N_24725);
and UO_1989 (O_1989,N_24841,N_24764);
nor UO_1990 (O_1990,N_24942,N_24767);
xor UO_1991 (O_1991,N_24595,N_24952);
xnor UO_1992 (O_1992,N_24738,N_24783);
nand UO_1993 (O_1993,N_24528,N_24672);
nor UO_1994 (O_1994,N_24802,N_24899);
xnor UO_1995 (O_1995,N_24891,N_24757);
xor UO_1996 (O_1996,N_24622,N_24808);
nor UO_1997 (O_1997,N_24532,N_24994);
nor UO_1998 (O_1998,N_24874,N_24709);
and UO_1999 (O_1999,N_24905,N_24524);
xor UO_2000 (O_2000,N_24530,N_24569);
and UO_2001 (O_2001,N_24576,N_24841);
and UO_2002 (O_2002,N_24619,N_24771);
and UO_2003 (O_2003,N_24831,N_24535);
and UO_2004 (O_2004,N_24711,N_24955);
xor UO_2005 (O_2005,N_24923,N_24867);
or UO_2006 (O_2006,N_24705,N_24799);
nor UO_2007 (O_2007,N_24557,N_24875);
nand UO_2008 (O_2008,N_24976,N_24565);
and UO_2009 (O_2009,N_24819,N_24873);
and UO_2010 (O_2010,N_24773,N_24748);
nor UO_2011 (O_2011,N_24854,N_24671);
xnor UO_2012 (O_2012,N_24817,N_24901);
nand UO_2013 (O_2013,N_24800,N_24674);
nor UO_2014 (O_2014,N_24931,N_24559);
and UO_2015 (O_2015,N_24951,N_24618);
xnor UO_2016 (O_2016,N_24783,N_24546);
xor UO_2017 (O_2017,N_24556,N_24898);
xor UO_2018 (O_2018,N_24526,N_24979);
and UO_2019 (O_2019,N_24676,N_24555);
nor UO_2020 (O_2020,N_24640,N_24564);
nor UO_2021 (O_2021,N_24739,N_24978);
and UO_2022 (O_2022,N_24707,N_24591);
nor UO_2023 (O_2023,N_24705,N_24500);
or UO_2024 (O_2024,N_24739,N_24720);
and UO_2025 (O_2025,N_24814,N_24783);
or UO_2026 (O_2026,N_24928,N_24700);
nor UO_2027 (O_2027,N_24821,N_24797);
and UO_2028 (O_2028,N_24766,N_24643);
nor UO_2029 (O_2029,N_24934,N_24610);
nand UO_2030 (O_2030,N_24537,N_24772);
nand UO_2031 (O_2031,N_24671,N_24982);
nand UO_2032 (O_2032,N_24863,N_24990);
xnor UO_2033 (O_2033,N_24893,N_24921);
nand UO_2034 (O_2034,N_24755,N_24655);
and UO_2035 (O_2035,N_24937,N_24723);
or UO_2036 (O_2036,N_24648,N_24715);
and UO_2037 (O_2037,N_24565,N_24962);
xnor UO_2038 (O_2038,N_24552,N_24712);
and UO_2039 (O_2039,N_24547,N_24580);
nand UO_2040 (O_2040,N_24884,N_24506);
or UO_2041 (O_2041,N_24790,N_24510);
xnor UO_2042 (O_2042,N_24860,N_24676);
or UO_2043 (O_2043,N_24765,N_24506);
or UO_2044 (O_2044,N_24981,N_24958);
nor UO_2045 (O_2045,N_24882,N_24613);
nor UO_2046 (O_2046,N_24623,N_24746);
nor UO_2047 (O_2047,N_24997,N_24871);
xnor UO_2048 (O_2048,N_24871,N_24815);
nor UO_2049 (O_2049,N_24934,N_24518);
nand UO_2050 (O_2050,N_24567,N_24851);
or UO_2051 (O_2051,N_24892,N_24709);
nand UO_2052 (O_2052,N_24936,N_24763);
or UO_2053 (O_2053,N_24964,N_24579);
xnor UO_2054 (O_2054,N_24535,N_24598);
or UO_2055 (O_2055,N_24706,N_24769);
nand UO_2056 (O_2056,N_24649,N_24865);
or UO_2057 (O_2057,N_24547,N_24715);
or UO_2058 (O_2058,N_24988,N_24782);
xnor UO_2059 (O_2059,N_24574,N_24714);
nand UO_2060 (O_2060,N_24701,N_24872);
or UO_2061 (O_2061,N_24677,N_24806);
or UO_2062 (O_2062,N_24969,N_24940);
xnor UO_2063 (O_2063,N_24629,N_24514);
or UO_2064 (O_2064,N_24807,N_24760);
nor UO_2065 (O_2065,N_24668,N_24627);
or UO_2066 (O_2066,N_24837,N_24637);
nor UO_2067 (O_2067,N_24945,N_24599);
nand UO_2068 (O_2068,N_24606,N_24600);
nor UO_2069 (O_2069,N_24628,N_24721);
xor UO_2070 (O_2070,N_24821,N_24529);
nand UO_2071 (O_2071,N_24559,N_24760);
xor UO_2072 (O_2072,N_24893,N_24804);
and UO_2073 (O_2073,N_24839,N_24555);
or UO_2074 (O_2074,N_24674,N_24847);
nor UO_2075 (O_2075,N_24949,N_24896);
nor UO_2076 (O_2076,N_24548,N_24898);
nor UO_2077 (O_2077,N_24505,N_24547);
or UO_2078 (O_2078,N_24928,N_24605);
nand UO_2079 (O_2079,N_24634,N_24646);
nand UO_2080 (O_2080,N_24543,N_24800);
and UO_2081 (O_2081,N_24744,N_24841);
or UO_2082 (O_2082,N_24832,N_24998);
xor UO_2083 (O_2083,N_24528,N_24831);
or UO_2084 (O_2084,N_24777,N_24691);
or UO_2085 (O_2085,N_24586,N_24700);
nand UO_2086 (O_2086,N_24920,N_24996);
nand UO_2087 (O_2087,N_24797,N_24655);
or UO_2088 (O_2088,N_24738,N_24555);
nand UO_2089 (O_2089,N_24921,N_24742);
and UO_2090 (O_2090,N_24628,N_24855);
and UO_2091 (O_2091,N_24834,N_24982);
nor UO_2092 (O_2092,N_24699,N_24898);
or UO_2093 (O_2093,N_24639,N_24536);
or UO_2094 (O_2094,N_24906,N_24603);
nand UO_2095 (O_2095,N_24569,N_24855);
nand UO_2096 (O_2096,N_24940,N_24889);
and UO_2097 (O_2097,N_24916,N_24531);
xnor UO_2098 (O_2098,N_24760,N_24823);
xnor UO_2099 (O_2099,N_24770,N_24567);
and UO_2100 (O_2100,N_24817,N_24877);
or UO_2101 (O_2101,N_24997,N_24545);
and UO_2102 (O_2102,N_24756,N_24838);
nand UO_2103 (O_2103,N_24506,N_24671);
and UO_2104 (O_2104,N_24502,N_24836);
xnor UO_2105 (O_2105,N_24538,N_24572);
nor UO_2106 (O_2106,N_24873,N_24567);
xor UO_2107 (O_2107,N_24588,N_24565);
nor UO_2108 (O_2108,N_24970,N_24854);
xnor UO_2109 (O_2109,N_24931,N_24617);
xor UO_2110 (O_2110,N_24585,N_24553);
nor UO_2111 (O_2111,N_24761,N_24675);
and UO_2112 (O_2112,N_24545,N_24805);
xnor UO_2113 (O_2113,N_24855,N_24745);
nor UO_2114 (O_2114,N_24998,N_24638);
and UO_2115 (O_2115,N_24703,N_24891);
nor UO_2116 (O_2116,N_24562,N_24902);
nand UO_2117 (O_2117,N_24606,N_24645);
and UO_2118 (O_2118,N_24688,N_24572);
and UO_2119 (O_2119,N_24596,N_24563);
or UO_2120 (O_2120,N_24850,N_24664);
and UO_2121 (O_2121,N_24953,N_24906);
nor UO_2122 (O_2122,N_24948,N_24786);
or UO_2123 (O_2123,N_24636,N_24676);
nand UO_2124 (O_2124,N_24856,N_24572);
xor UO_2125 (O_2125,N_24687,N_24722);
and UO_2126 (O_2126,N_24875,N_24714);
or UO_2127 (O_2127,N_24819,N_24583);
or UO_2128 (O_2128,N_24646,N_24796);
or UO_2129 (O_2129,N_24519,N_24723);
and UO_2130 (O_2130,N_24860,N_24828);
or UO_2131 (O_2131,N_24554,N_24724);
nor UO_2132 (O_2132,N_24507,N_24531);
or UO_2133 (O_2133,N_24508,N_24804);
xor UO_2134 (O_2134,N_24901,N_24779);
xnor UO_2135 (O_2135,N_24711,N_24551);
and UO_2136 (O_2136,N_24586,N_24761);
xnor UO_2137 (O_2137,N_24805,N_24673);
nor UO_2138 (O_2138,N_24846,N_24728);
or UO_2139 (O_2139,N_24575,N_24503);
xnor UO_2140 (O_2140,N_24518,N_24994);
xnor UO_2141 (O_2141,N_24885,N_24981);
xor UO_2142 (O_2142,N_24990,N_24820);
nand UO_2143 (O_2143,N_24729,N_24565);
nor UO_2144 (O_2144,N_24510,N_24988);
xnor UO_2145 (O_2145,N_24604,N_24966);
nand UO_2146 (O_2146,N_24760,N_24577);
nor UO_2147 (O_2147,N_24922,N_24703);
and UO_2148 (O_2148,N_24612,N_24987);
nand UO_2149 (O_2149,N_24863,N_24582);
and UO_2150 (O_2150,N_24886,N_24818);
nand UO_2151 (O_2151,N_24664,N_24760);
nand UO_2152 (O_2152,N_24909,N_24963);
or UO_2153 (O_2153,N_24713,N_24622);
or UO_2154 (O_2154,N_24758,N_24968);
or UO_2155 (O_2155,N_24929,N_24645);
xor UO_2156 (O_2156,N_24532,N_24553);
nand UO_2157 (O_2157,N_24514,N_24933);
nor UO_2158 (O_2158,N_24951,N_24934);
xnor UO_2159 (O_2159,N_24883,N_24650);
xnor UO_2160 (O_2160,N_24626,N_24554);
nor UO_2161 (O_2161,N_24561,N_24741);
and UO_2162 (O_2162,N_24534,N_24976);
and UO_2163 (O_2163,N_24985,N_24545);
nor UO_2164 (O_2164,N_24924,N_24645);
nand UO_2165 (O_2165,N_24871,N_24690);
xor UO_2166 (O_2166,N_24593,N_24594);
xnor UO_2167 (O_2167,N_24694,N_24894);
and UO_2168 (O_2168,N_24729,N_24824);
xor UO_2169 (O_2169,N_24852,N_24977);
or UO_2170 (O_2170,N_24968,N_24637);
nor UO_2171 (O_2171,N_24674,N_24831);
or UO_2172 (O_2172,N_24814,N_24806);
xor UO_2173 (O_2173,N_24548,N_24574);
and UO_2174 (O_2174,N_24996,N_24932);
nand UO_2175 (O_2175,N_24627,N_24563);
xnor UO_2176 (O_2176,N_24748,N_24676);
nor UO_2177 (O_2177,N_24893,N_24503);
and UO_2178 (O_2178,N_24791,N_24597);
nor UO_2179 (O_2179,N_24702,N_24707);
and UO_2180 (O_2180,N_24509,N_24600);
xnor UO_2181 (O_2181,N_24767,N_24796);
and UO_2182 (O_2182,N_24594,N_24755);
nor UO_2183 (O_2183,N_24749,N_24892);
and UO_2184 (O_2184,N_24588,N_24880);
and UO_2185 (O_2185,N_24825,N_24743);
nand UO_2186 (O_2186,N_24663,N_24640);
or UO_2187 (O_2187,N_24576,N_24836);
and UO_2188 (O_2188,N_24938,N_24916);
nor UO_2189 (O_2189,N_24831,N_24612);
xnor UO_2190 (O_2190,N_24582,N_24850);
xnor UO_2191 (O_2191,N_24571,N_24970);
nor UO_2192 (O_2192,N_24899,N_24984);
or UO_2193 (O_2193,N_24694,N_24595);
xnor UO_2194 (O_2194,N_24714,N_24950);
xor UO_2195 (O_2195,N_24623,N_24646);
and UO_2196 (O_2196,N_24514,N_24511);
nor UO_2197 (O_2197,N_24809,N_24858);
nand UO_2198 (O_2198,N_24925,N_24610);
nor UO_2199 (O_2199,N_24598,N_24761);
and UO_2200 (O_2200,N_24648,N_24633);
xor UO_2201 (O_2201,N_24858,N_24846);
xor UO_2202 (O_2202,N_24927,N_24640);
nor UO_2203 (O_2203,N_24907,N_24770);
xnor UO_2204 (O_2204,N_24795,N_24844);
and UO_2205 (O_2205,N_24622,N_24847);
xor UO_2206 (O_2206,N_24765,N_24776);
or UO_2207 (O_2207,N_24678,N_24763);
and UO_2208 (O_2208,N_24890,N_24507);
and UO_2209 (O_2209,N_24940,N_24963);
or UO_2210 (O_2210,N_24530,N_24997);
nor UO_2211 (O_2211,N_24524,N_24938);
and UO_2212 (O_2212,N_24897,N_24669);
and UO_2213 (O_2213,N_24713,N_24844);
nor UO_2214 (O_2214,N_24546,N_24642);
and UO_2215 (O_2215,N_24828,N_24521);
xor UO_2216 (O_2216,N_24758,N_24979);
xnor UO_2217 (O_2217,N_24835,N_24721);
and UO_2218 (O_2218,N_24740,N_24580);
and UO_2219 (O_2219,N_24682,N_24997);
nor UO_2220 (O_2220,N_24587,N_24630);
nand UO_2221 (O_2221,N_24500,N_24981);
nand UO_2222 (O_2222,N_24990,N_24662);
nand UO_2223 (O_2223,N_24777,N_24841);
xor UO_2224 (O_2224,N_24758,N_24706);
nand UO_2225 (O_2225,N_24546,N_24927);
or UO_2226 (O_2226,N_24532,N_24934);
nor UO_2227 (O_2227,N_24985,N_24504);
nand UO_2228 (O_2228,N_24923,N_24974);
and UO_2229 (O_2229,N_24584,N_24520);
and UO_2230 (O_2230,N_24571,N_24560);
nand UO_2231 (O_2231,N_24701,N_24973);
nor UO_2232 (O_2232,N_24905,N_24879);
nand UO_2233 (O_2233,N_24660,N_24684);
and UO_2234 (O_2234,N_24851,N_24695);
or UO_2235 (O_2235,N_24570,N_24553);
or UO_2236 (O_2236,N_24608,N_24516);
nor UO_2237 (O_2237,N_24767,N_24693);
nand UO_2238 (O_2238,N_24855,N_24615);
nand UO_2239 (O_2239,N_24710,N_24980);
nand UO_2240 (O_2240,N_24819,N_24610);
xor UO_2241 (O_2241,N_24564,N_24778);
xor UO_2242 (O_2242,N_24506,N_24999);
nor UO_2243 (O_2243,N_24540,N_24771);
nand UO_2244 (O_2244,N_24961,N_24808);
nand UO_2245 (O_2245,N_24705,N_24700);
xor UO_2246 (O_2246,N_24978,N_24822);
nor UO_2247 (O_2247,N_24666,N_24899);
nor UO_2248 (O_2248,N_24855,N_24777);
nor UO_2249 (O_2249,N_24933,N_24500);
nor UO_2250 (O_2250,N_24756,N_24939);
xnor UO_2251 (O_2251,N_24581,N_24821);
or UO_2252 (O_2252,N_24574,N_24983);
nand UO_2253 (O_2253,N_24994,N_24727);
nor UO_2254 (O_2254,N_24709,N_24746);
nand UO_2255 (O_2255,N_24544,N_24671);
xor UO_2256 (O_2256,N_24696,N_24732);
nand UO_2257 (O_2257,N_24898,N_24983);
nand UO_2258 (O_2258,N_24962,N_24922);
and UO_2259 (O_2259,N_24546,N_24723);
xor UO_2260 (O_2260,N_24529,N_24715);
nor UO_2261 (O_2261,N_24671,N_24912);
nor UO_2262 (O_2262,N_24665,N_24774);
nand UO_2263 (O_2263,N_24563,N_24807);
nor UO_2264 (O_2264,N_24538,N_24738);
or UO_2265 (O_2265,N_24973,N_24774);
and UO_2266 (O_2266,N_24500,N_24655);
and UO_2267 (O_2267,N_24734,N_24565);
nor UO_2268 (O_2268,N_24559,N_24859);
or UO_2269 (O_2269,N_24568,N_24633);
or UO_2270 (O_2270,N_24917,N_24924);
and UO_2271 (O_2271,N_24667,N_24895);
nor UO_2272 (O_2272,N_24789,N_24794);
or UO_2273 (O_2273,N_24669,N_24532);
xor UO_2274 (O_2274,N_24693,N_24707);
and UO_2275 (O_2275,N_24576,N_24703);
and UO_2276 (O_2276,N_24864,N_24617);
or UO_2277 (O_2277,N_24553,N_24903);
nor UO_2278 (O_2278,N_24569,N_24891);
xnor UO_2279 (O_2279,N_24870,N_24958);
and UO_2280 (O_2280,N_24772,N_24981);
or UO_2281 (O_2281,N_24997,N_24954);
nor UO_2282 (O_2282,N_24739,N_24989);
nor UO_2283 (O_2283,N_24727,N_24834);
nor UO_2284 (O_2284,N_24788,N_24746);
or UO_2285 (O_2285,N_24788,N_24633);
xor UO_2286 (O_2286,N_24813,N_24555);
nor UO_2287 (O_2287,N_24932,N_24671);
nor UO_2288 (O_2288,N_24560,N_24739);
nor UO_2289 (O_2289,N_24523,N_24627);
nor UO_2290 (O_2290,N_24645,N_24720);
or UO_2291 (O_2291,N_24564,N_24541);
xnor UO_2292 (O_2292,N_24927,N_24589);
nand UO_2293 (O_2293,N_24635,N_24811);
nand UO_2294 (O_2294,N_24563,N_24511);
and UO_2295 (O_2295,N_24582,N_24729);
nor UO_2296 (O_2296,N_24542,N_24799);
nor UO_2297 (O_2297,N_24813,N_24702);
or UO_2298 (O_2298,N_24759,N_24864);
or UO_2299 (O_2299,N_24633,N_24771);
or UO_2300 (O_2300,N_24600,N_24876);
or UO_2301 (O_2301,N_24559,N_24937);
nor UO_2302 (O_2302,N_24899,N_24763);
nand UO_2303 (O_2303,N_24906,N_24910);
nand UO_2304 (O_2304,N_24895,N_24771);
or UO_2305 (O_2305,N_24883,N_24544);
or UO_2306 (O_2306,N_24977,N_24731);
nand UO_2307 (O_2307,N_24810,N_24753);
nor UO_2308 (O_2308,N_24877,N_24653);
nand UO_2309 (O_2309,N_24834,N_24702);
xor UO_2310 (O_2310,N_24621,N_24947);
or UO_2311 (O_2311,N_24570,N_24559);
xor UO_2312 (O_2312,N_24550,N_24958);
nand UO_2313 (O_2313,N_24684,N_24882);
nand UO_2314 (O_2314,N_24857,N_24523);
or UO_2315 (O_2315,N_24889,N_24917);
and UO_2316 (O_2316,N_24956,N_24816);
nand UO_2317 (O_2317,N_24709,N_24988);
xnor UO_2318 (O_2318,N_24990,N_24872);
nor UO_2319 (O_2319,N_24857,N_24685);
nor UO_2320 (O_2320,N_24798,N_24759);
nor UO_2321 (O_2321,N_24515,N_24804);
nand UO_2322 (O_2322,N_24942,N_24790);
and UO_2323 (O_2323,N_24594,N_24681);
nand UO_2324 (O_2324,N_24893,N_24848);
nor UO_2325 (O_2325,N_24527,N_24977);
nor UO_2326 (O_2326,N_24870,N_24751);
nand UO_2327 (O_2327,N_24874,N_24507);
nand UO_2328 (O_2328,N_24920,N_24743);
and UO_2329 (O_2329,N_24589,N_24934);
and UO_2330 (O_2330,N_24672,N_24745);
nor UO_2331 (O_2331,N_24826,N_24835);
nand UO_2332 (O_2332,N_24587,N_24706);
and UO_2333 (O_2333,N_24700,N_24783);
xnor UO_2334 (O_2334,N_24934,N_24566);
nand UO_2335 (O_2335,N_24685,N_24882);
and UO_2336 (O_2336,N_24791,N_24728);
nand UO_2337 (O_2337,N_24883,N_24995);
or UO_2338 (O_2338,N_24784,N_24629);
nor UO_2339 (O_2339,N_24946,N_24590);
nor UO_2340 (O_2340,N_24956,N_24754);
nor UO_2341 (O_2341,N_24956,N_24873);
and UO_2342 (O_2342,N_24733,N_24976);
nor UO_2343 (O_2343,N_24757,N_24674);
xor UO_2344 (O_2344,N_24733,N_24994);
nand UO_2345 (O_2345,N_24937,N_24540);
nand UO_2346 (O_2346,N_24521,N_24903);
or UO_2347 (O_2347,N_24544,N_24535);
nand UO_2348 (O_2348,N_24911,N_24898);
nand UO_2349 (O_2349,N_24987,N_24928);
or UO_2350 (O_2350,N_24551,N_24969);
nor UO_2351 (O_2351,N_24508,N_24519);
or UO_2352 (O_2352,N_24937,N_24519);
xnor UO_2353 (O_2353,N_24776,N_24740);
or UO_2354 (O_2354,N_24647,N_24612);
or UO_2355 (O_2355,N_24531,N_24528);
nor UO_2356 (O_2356,N_24933,N_24719);
or UO_2357 (O_2357,N_24534,N_24936);
and UO_2358 (O_2358,N_24855,N_24871);
nand UO_2359 (O_2359,N_24562,N_24610);
nor UO_2360 (O_2360,N_24899,N_24754);
or UO_2361 (O_2361,N_24916,N_24741);
xnor UO_2362 (O_2362,N_24548,N_24837);
xor UO_2363 (O_2363,N_24994,N_24508);
nor UO_2364 (O_2364,N_24604,N_24926);
xnor UO_2365 (O_2365,N_24870,N_24863);
nand UO_2366 (O_2366,N_24555,N_24683);
xor UO_2367 (O_2367,N_24936,N_24968);
nand UO_2368 (O_2368,N_24575,N_24820);
nand UO_2369 (O_2369,N_24793,N_24632);
xnor UO_2370 (O_2370,N_24860,N_24921);
nand UO_2371 (O_2371,N_24986,N_24529);
xnor UO_2372 (O_2372,N_24538,N_24600);
and UO_2373 (O_2373,N_24764,N_24763);
xor UO_2374 (O_2374,N_24902,N_24959);
xnor UO_2375 (O_2375,N_24518,N_24895);
xor UO_2376 (O_2376,N_24781,N_24767);
or UO_2377 (O_2377,N_24820,N_24727);
nor UO_2378 (O_2378,N_24690,N_24951);
nand UO_2379 (O_2379,N_24700,N_24744);
nand UO_2380 (O_2380,N_24915,N_24881);
and UO_2381 (O_2381,N_24527,N_24559);
xor UO_2382 (O_2382,N_24907,N_24929);
or UO_2383 (O_2383,N_24698,N_24656);
nor UO_2384 (O_2384,N_24942,N_24524);
nand UO_2385 (O_2385,N_24505,N_24728);
xor UO_2386 (O_2386,N_24864,N_24776);
nor UO_2387 (O_2387,N_24996,N_24633);
or UO_2388 (O_2388,N_24697,N_24579);
xnor UO_2389 (O_2389,N_24566,N_24836);
and UO_2390 (O_2390,N_24626,N_24852);
xor UO_2391 (O_2391,N_24614,N_24789);
xnor UO_2392 (O_2392,N_24566,N_24868);
and UO_2393 (O_2393,N_24535,N_24505);
and UO_2394 (O_2394,N_24879,N_24810);
xnor UO_2395 (O_2395,N_24981,N_24868);
nand UO_2396 (O_2396,N_24654,N_24623);
or UO_2397 (O_2397,N_24886,N_24608);
xnor UO_2398 (O_2398,N_24804,N_24778);
xor UO_2399 (O_2399,N_24892,N_24957);
or UO_2400 (O_2400,N_24921,N_24692);
nand UO_2401 (O_2401,N_24695,N_24926);
and UO_2402 (O_2402,N_24649,N_24709);
nand UO_2403 (O_2403,N_24820,N_24954);
nor UO_2404 (O_2404,N_24736,N_24537);
and UO_2405 (O_2405,N_24614,N_24781);
and UO_2406 (O_2406,N_24890,N_24502);
xor UO_2407 (O_2407,N_24612,N_24845);
nand UO_2408 (O_2408,N_24865,N_24502);
nand UO_2409 (O_2409,N_24941,N_24880);
nand UO_2410 (O_2410,N_24816,N_24973);
and UO_2411 (O_2411,N_24650,N_24709);
xnor UO_2412 (O_2412,N_24856,N_24749);
or UO_2413 (O_2413,N_24874,N_24803);
nand UO_2414 (O_2414,N_24520,N_24824);
nor UO_2415 (O_2415,N_24725,N_24924);
and UO_2416 (O_2416,N_24964,N_24900);
xnor UO_2417 (O_2417,N_24717,N_24582);
nor UO_2418 (O_2418,N_24700,N_24815);
nor UO_2419 (O_2419,N_24582,N_24712);
or UO_2420 (O_2420,N_24545,N_24717);
nor UO_2421 (O_2421,N_24787,N_24848);
nand UO_2422 (O_2422,N_24851,N_24513);
or UO_2423 (O_2423,N_24931,N_24514);
or UO_2424 (O_2424,N_24666,N_24513);
nor UO_2425 (O_2425,N_24642,N_24909);
or UO_2426 (O_2426,N_24974,N_24852);
xnor UO_2427 (O_2427,N_24713,N_24610);
or UO_2428 (O_2428,N_24888,N_24510);
xor UO_2429 (O_2429,N_24836,N_24700);
and UO_2430 (O_2430,N_24911,N_24692);
and UO_2431 (O_2431,N_24753,N_24697);
or UO_2432 (O_2432,N_24867,N_24984);
or UO_2433 (O_2433,N_24947,N_24824);
or UO_2434 (O_2434,N_24513,N_24919);
or UO_2435 (O_2435,N_24614,N_24725);
xnor UO_2436 (O_2436,N_24685,N_24702);
and UO_2437 (O_2437,N_24965,N_24921);
and UO_2438 (O_2438,N_24991,N_24839);
and UO_2439 (O_2439,N_24697,N_24859);
or UO_2440 (O_2440,N_24666,N_24735);
and UO_2441 (O_2441,N_24779,N_24702);
xor UO_2442 (O_2442,N_24591,N_24984);
nor UO_2443 (O_2443,N_24582,N_24666);
and UO_2444 (O_2444,N_24803,N_24905);
xnor UO_2445 (O_2445,N_24835,N_24740);
xnor UO_2446 (O_2446,N_24642,N_24978);
or UO_2447 (O_2447,N_24697,N_24632);
and UO_2448 (O_2448,N_24773,N_24949);
and UO_2449 (O_2449,N_24903,N_24853);
xor UO_2450 (O_2450,N_24990,N_24807);
or UO_2451 (O_2451,N_24681,N_24637);
or UO_2452 (O_2452,N_24549,N_24970);
nand UO_2453 (O_2453,N_24808,N_24535);
nand UO_2454 (O_2454,N_24879,N_24811);
and UO_2455 (O_2455,N_24511,N_24673);
xnor UO_2456 (O_2456,N_24876,N_24516);
xnor UO_2457 (O_2457,N_24578,N_24954);
and UO_2458 (O_2458,N_24665,N_24644);
nand UO_2459 (O_2459,N_24850,N_24775);
xnor UO_2460 (O_2460,N_24922,N_24894);
nor UO_2461 (O_2461,N_24628,N_24874);
or UO_2462 (O_2462,N_24701,N_24787);
xnor UO_2463 (O_2463,N_24865,N_24884);
nand UO_2464 (O_2464,N_24715,N_24967);
and UO_2465 (O_2465,N_24500,N_24536);
nand UO_2466 (O_2466,N_24901,N_24997);
nor UO_2467 (O_2467,N_24938,N_24838);
and UO_2468 (O_2468,N_24607,N_24687);
nor UO_2469 (O_2469,N_24792,N_24754);
nand UO_2470 (O_2470,N_24689,N_24574);
and UO_2471 (O_2471,N_24723,N_24712);
nor UO_2472 (O_2472,N_24989,N_24735);
xnor UO_2473 (O_2473,N_24888,N_24528);
xor UO_2474 (O_2474,N_24606,N_24817);
or UO_2475 (O_2475,N_24752,N_24846);
and UO_2476 (O_2476,N_24556,N_24924);
and UO_2477 (O_2477,N_24649,N_24640);
nor UO_2478 (O_2478,N_24686,N_24798);
nand UO_2479 (O_2479,N_24656,N_24748);
or UO_2480 (O_2480,N_24700,N_24608);
xnor UO_2481 (O_2481,N_24711,N_24641);
nand UO_2482 (O_2482,N_24685,N_24927);
xor UO_2483 (O_2483,N_24700,N_24871);
xor UO_2484 (O_2484,N_24771,N_24745);
nand UO_2485 (O_2485,N_24916,N_24935);
or UO_2486 (O_2486,N_24623,N_24717);
nor UO_2487 (O_2487,N_24653,N_24835);
xor UO_2488 (O_2488,N_24919,N_24967);
xor UO_2489 (O_2489,N_24574,N_24518);
nand UO_2490 (O_2490,N_24626,N_24647);
and UO_2491 (O_2491,N_24609,N_24631);
nand UO_2492 (O_2492,N_24859,N_24829);
nand UO_2493 (O_2493,N_24589,N_24876);
nand UO_2494 (O_2494,N_24527,N_24756);
xor UO_2495 (O_2495,N_24551,N_24895);
and UO_2496 (O_2496,N_24756,N_24721);
nand UO_2497 (O_2497,N_24568,N_24572);
nand UO_2498 (O_2498,N_24950,N_24975);
or UO_2499 (O_2499,N_24964,N_24655);
nor UO_2500 (O_2500,N_24894,N_24537);
xnor UO_2501 (O_2501,N_24937,N_24681);
or UO_2502 (O_2502,N_24872,N_24656);
nand UO_2503 (O_2503,N_24733,N_24980);
xor UO_2504 (O_2504,N_24801,N_24828);
nor UO_2505 (O_2505,N_24586,N_24772);
xnor UO_2506 (O_2506,N_24645,N_24554);
xor UO_2507 (O_2507,N_24715,N_24781);
or UO_2508 (O_2508,N_24976,N_24567);
xnor UO_2509 (O_2509,N_24840,N_24552);
nor UO_2510 (O_2510,N_24847,N_24607);
and UO_2511 (O_2511,N_24734,N_24891);
and UO_2512 (O_2512,N_24863,N_24611);
and UO_2513 (O_2513,N_24654,N_24766);
nor UO_2514 (O_2514,N_24699,N_24963);
and UO_2515 (O_2515,N_24968,N_24704);
and UO_2516 (O_2516,N_24549,N_24564);
nor UO_2517 (O_2517,N_24644,N_24746);
nor UO_2518 (O_2518,N_24886,N_24705);
and UO_2519 (O_2519,N_24721,N_24612);
nand UO_2520 (O_2520,N_24855,N_24993);
nand UO_2521 (O_2521,N_24750,N_24641);
nor UO_2522 (O_2522,N_24756,N_24525);
xnor UO_2523 (O_2523,N_24505,N_24760);
or UO_2524 (O_2524,N_24797,N_24887);
xnor UO_2525 (O_2525,N_24699,N_24879);
or UO_2526 (O_2526,N_24683,N_24830);
and UO_2527 (O_2527,N_24834,N_24654);
nor UO_2528 (O_2528,N_24547,N_24899);
or UO_2529 (O_2529,N_24660,N_24531);
xnor UO_2530 (O_2530,N_24883,N_24694);
and UO_2531 (O_2531,N_24586,N_24782);
or UO_2532 (O_2532,N_24530,N_24544);
xor UO_2533 (O_2533,N_24850,N_24567);
nand UO_2534 (O_2534,N_24978,N_24666);
or UO_2535 (O_2535,N_24914,N_24562);
nand UO_2536 (O_2536,N_24670,N_24737);
and UO_2537 (O_2537,N_24922,N_24648);
nor UO_2538 (O_2538,N_24908,N_24717);
xor UO_2539 (O_2539,N_24969,N_24541);
nor UO_2540 (O_2540,N_24622,N_24518);
or UO_2541 (O_2541,N_24776,N_24772);
or UO_2542 (O_2542,N_24868,N_24698);
nor UO_2543 (O_2543,N_24600,N_24813);
nand UO_2544 (O_2544,N_24822,N_24542);
nor UO_2545 (O_2545,N_24793,N_24845);
and UO_2546 (O_2546,N_24918,N_24856);
xor UO_2547 (O_2547,N_24848,N_24984);
xor UO_2548 (O_2548,N_24643,N_24938);
and UO_2549 (O_2549,N_24723,N_24625);
nor UO_2550 (O_2550,N_24835,N_24961);
or UO_2551 (O_2551,N_24593,N_24700);
or UO_2552 (O_2552,N_24763,N_24650);
and UO_2553 (O_2553,N_24803,N_24776);
or UO_2554 (O_2554,N_24917,N_24778);
nand UO_2555 (O_2555,N_24944,N_24844);
or UO_2556 (O_2556,N_24832,N_24516);
or UO_2557 (O_2557,N_24957,N_24918);
nand UO_2558 (O_2558,N_24549,N_24529);
or UO_2559 (O_2559,N_24994,N_24527);
nand UO_2560 (O_2560,N_24775,N_24926);
or UO_2561 (O_2561,N_24923,N_24841);
or UO_2562 (O_2562,N_24628,N_24842);
xor UO_2563 (O_2563,N_24714,N_24512);
and UO_2564 (O_2564,N_24565,N_24512);
xnor UO_2565 (O_2565,N_24595,N_24546);
xnor UO_2566 (O_2566,N_24841,N_24824);
or UO_2567 (O_2567,N_24819,N_24858);
xnor UO_2568 (O_2568,N_24936,N_24973);
or UO_2569 (O_2569,N_24857,N_24863);
and UO_2570 (O_2570,N_24717,N_24917);
or UO_2571 (O_2571,N_24930,N_24834);
xnor UO_2572 (O_2572,N_24988,N_24743);
nand UO_2573 (O_2573,N_24581,N_24985);
xnor UO_2574 (O_2574,N_24996,N_24692);
nand UO_2575 (O_2575,N_24973,N_24923);
or UO_2576 (O_2576,N_24592,N_24861);
or UO_2577 (O_2577,N_24783,N_24859);
and UO_2578 (O_2578,N_24958,N_24883);
or UO_2579 (O_2579,N_24580,N_24708);
nand UO_2580 (O_2580,N_24559,N_24676);
or UO_2581 (O_2581,N_24757,N_24864);
xnor UO_2582 (O_2582,N_24530,N_24548);
and UO_2583 (O_2583,N_24526,N_24909);
xor UO_2584 (O_2584,N_24552,N_24722);
xnor UO_2585 (O_2585,N_24526,N_24986);
nor UO_2586 (O_2586,N_24575,N_24621);
or UO_2587 (O_2587,N_24532,N_24998);
nand UO_2588 (O_2588,N_24649,N_24790);
or UO_2589 (O_2589,N_24637,N_24594);
nor UO_2590 (O_2590,N_24835,N_24831);
xor UO_2591 (O_2591,N_24738,N_24520);
and UO_2592 (O_2592,N_24999,N_24789);
or UO_2593 (O_2593,N_24514,N_24542);
and UO_2594 (O_2594,N_24942,N_24694);
nor UO_2595 (O_2595,N_24633,N_24906);
and UO_2596 (O_2596,N_24692,N_24769);
or UO_2597 (O_2597,N_24877,N_24587);
nor UO_2598 (O_2598,N_24817,N_24587);
xor UO_2599 (O_2599,N_24835,N_24706);
xnor UO_2600 (O_2600,N_24996,N_24599);
nand UO_2601 (O_2601,N_24931,N_24786);
xor UO_2602 (O_2602,N_24988,N_24857);
xor UO_2603 (O_2603,N_24840,N_24959);
xor UO_2604 (O_2604,N_24699,N_24952);
and UO_2605 (O_2605,N_24659,N_24812);
xor UO_2606 (O_2606,N_24993,N_24981);
and UO_2607 (O_2607,N_24659,N_24558);
or UO_2608 (O_2608,N_24641,N_24715);
xnor UO_2609 (O_2609,N_24974,N_24743);
and UO_2610 (O_2610,N_24610,N_24715);
nor UO_2611 (O_2611,N_24845,N_24969);
and UO_2612 (O_2612,N_24649,N_24750);
nand UO_2613 (O_2613,N_24574,N_24736);
nor UO_2614 (O_2614,N_24500,N_24772);
and UO_2615 (O_2615,N_24616,N_24538);
and UO_2616 (O_2616,N_24861,N_24660);
and UO_2617 (O_2617,N_24951,N_24733);
or UO_2618 (O_2618,N_24783,N_24772);
and UO_2619 (O_2619,N_24568,N_24761);
xnor UO_2620 (O_2620,N_24993,N_24951);
or UO_2621 (O_2621,N_24980,N_24779);
and UO_2622 (O_2622,N_24545,N_24599);
and UO_2623 (O_2623,N_24504,N_24782);
nor UO_2624 (O_2624,N_24761,N_24672);
and UO_2625 (O_2625,N_24913,N_24981);
xnor UO_2626 (O_2626,N_24885,N_24994);
nor UO_2627 (O_2627,N_24520,N_24618);
nor UO_2628 (O_2628,N_24955,N_24817);
xor UO_2629 (O_2629,N_24950,N_24751);
nand UO_2630 (O_2630,N_24853,N_24530);
xor UO_2631 (O_2631,N_24933,N_24930);
and UO_2632 (O_2632,N_24905,N_24862);
or UO_2633 (O_2633,N_24871,N_24751);
or UO_2634 (O_2634,N_24800,N_24656);
xnor UO_2635 (O_2635,N_24539,N_24912);
nor UO_2636 (O_2636,N_24712,N_24703);
and UO_2637 (O_2637,N_24892,N_24832);
or UO_2638 (O_2638,N_24958,N_24789);
xnor UO_2639 (O_2639,N_24577,N_24589);
or UO_2640 (O_2640,N_24671,N_24821);
or UO_2641 (O_2641,N_24808,N_24922);
xor UO_2642 (O_2642,N_24688,N_24759);
and UO_2643 (O_2643,N_24921,N_24537);
or UO_2644 (O_2644,N_24542,N_24805);
nand UO_2645 (O_2645,N_24644,N_24577);
and UO_2646 (O_2646,N_24713,N_24742);
nor UO_2647 (O_2647,N_24839,N_24762);
nand UO_2648 (O_2648,N_24772,N_24781);
nor UO_2649 (O_2649,N_24659,N_24819);
and UO_2650 (O_2650,N_24816,N_24571);
and UO_2651 (O_2651,N_24836,N_24708);
or UO_2652 (O_2652,N_24589,N_24630);
or UO_2653 (O_2653,N_24612,N_24627);
nor UO_2654 (O_2654,N_24656,N_24590);
or UO_2655 (O_2655,N_24648,N_24939);
or UO_2656 (O_2656,N_24984,N_24643);
xor UO_2657 (O_2657,N_24540,N_24866);
nor UO_2658 (O_2658,N_24939,N_24663);
and UO_2659 (O_2659,N_24990,N_24504);
nand UO_2660 (O_2660,N_24886,N_24989);
xor UO_2661 (O_2661,N_24656,N_24511);
nor UO_2662 (O_2662,N_24989,N_24823);
and UO_2663 (O_2663,N_24567,N_24685);
nand UO_2664 (O_2664,N_24820,N_24911);
nand UO_2665 (O_2665,N_24933,N_24647);
or UO_2666 (O_2666,N_24630,N_24516);
or UO_2667 (O_2667,N_24760,N_24937);
nand UO_2668 (O_2668,N_24690,N_24998);
nand UO_2669 (O_2669,N_24602,N_24988);
xnor UO_2670 (O_2670,N_24682,N_24514);
xnor UO_2671 (O_2671,N_24617,N_24854);
nor UO_2672 (O_2672,N_24889,N_24819);
or UO_2673 (O_2673,N_24631,N_24788);
nand UO_2674 (O_2674,N_24956,N_24675);
or UO_2675 (O_2675,N_24978,N_24515);
or UO_2676 (O_2676,N_24737,N_24746);
or UO_2677 (O_2677,N_24903,N_24518);
nor UO_2678 (O_2678,N_24854,N_24819);
nand UO_2679 (O_2679,N_24520,N_24869);
xor UO_2680 (O_2680,N_24774,N_24914);
and UO_2681 (O_2681,N_24973,N_24977);
nand UO_2682 (O_2682,N_24537,N_24673);
or UO_2683 (O_2683,N_24519,N_24715);
and UO_2684 (O_2684,N_24799,N_24683);
xnor UO_2685 (O_2685,N_24604,N_24977);
xor UO_2686 (O_2686,N_24680,N_24999);
and UO_2687 (O_2687,N_24866,N_24556);
nor UO_2688 (O_2688,N_24866,N_24941);
nor UO_2689 (O_2689,N_24777,N_24513);
nand UO_2690 (O_2690,N_24955,N_24868);
nand UO_2691 (O_2691,N_24511,N_24647);
nand UO_2692 (O_2692,N_24688,N_24859);
and UO_2693 (O_2693,N_24912,N_24852);
or UO_2694 (O_2694,N_24758,N_24914);
and UO_2695 (O_2695,N_24528,N_24501);
xor UO_2696 (O_2696,N_24552,N_24885);
nand UO_2697 (O_2697,N_24722,N_24810);
or UO_2698 (O_2698,N_24504,N_24760);
or UO_2699 (O_2699,N_24772,N_24660);
nand UO_2700 (O_2700,N_24737,N_24768);
nor UO_2701 (O_2701,N_24834,N_24801);
or UO_2702 (O_2702,N_24632,N_24932);
and UO_2703 (O_2703,N_24561,N_24961);
nand UO_2704 (O_2704,N_24986,N_24524);
xnor UO_2705 (O_2705,N_24929,N_24575);
and UO_2706 (O_2706,N_24764,N_24556);
xnor UO_2707 (O_2707,N_24995,N_24979);
nor UO_2708 (O_2708,N_24720,N_24911);
and UO_2709 (O_2709,N_24780,N_24573);
and UO_2710 (O_2710,N_24852,N_24796);
and UO_2711 (O_2711,N_24989,N_24717);
xor UO_2712 (O_2712,N_24875,N_24742);
and UO_2713 (O_2713,N_24774,N_24737);
xnor UO_2714 (O_2714,N_24519,N_24952);
or UO_2715 (O_2715,N_24797,N_24525);
or UO_2716 (O_2716,N_24735,N_24531);
nand UO_2717 (O_2717,N_24961,N_24965);
xor UO_2718 (O_2718,N_24929,N_24750);
nand UO_2719 (O_2719,N_24639,N_24501);
or UO_2720 (O_2720,N_24958,N_24709);
nand UO_2721 (O_2721,N_24805,N_24984);
and UO_2722 (O_2722,N_24767,N_24514);
nand UO_2723 (O_2723,N_24535,N_24523);
nor UO_2724 (O_2724,N_24634,N_24624);
and UO_2725 (O_2725,N_24780,N_24523);
or UO_2726 (O_2726,N_24521,N_24816);
nor UO_2727 (O_2727,N_24982,N_24616);
nand UO_2728 (O_2728,N_24688,N_24810);
and UO_2729 (O_2729,N_24986,N_24504);
and UO_2730 (O_2730,N_24696,N_24632);
nand UO_2731 (O_2731,N_24629,N_24796);
or UO_2732 (O_2732,N_24998,N_24579);
or UO_2733 (O_2733,N_24693,N_24689);
or UO_2734 (O_2734,N_24948,N_24530);
nor UO_2735 (O_2735,N_24863,N_24702);
xor UO_2736 (O_2736,N_24900,N_24674);
or UO_2737 (O_2737,N_24935,N_24563);
or UO_2738 (O_2738,N_24670,N_24880);
xor UO_2739 (O_2739,N_24903,N_24656);
nand UO_2740 (O_2740,N_24556,N_24643);
xnor UO_2741 (O_2741,N_24811,N_24977);
xor UO_2742 (O_2742,N_24549,N_24548);
nor UO_2743 (O_2743,N_24880,N_24630);
and UO_2744 (O_2744,N_24784,N_24547);
and UO_2745 (O_2745,N_24757,N_24692);
nor UO_2746 (O_2746,N_24655,N_24979);
xor UO_2747 (O_2747,N_24689,N_24768);
nand UO_2748 (O_2748,N_24814,N_24505);
nor UO_2749 (O_2749,N_24878,N_24635);
xnor UO_2750 (O_2750,N_24584,N_24566);
or UO_2751 (O_2751,N_24737,N_24862);
xor UO_2752 (O_2752,N_24549,N_24839);
nand UO_2753 (O_2753,N_24788,N_24881);
or UO_2754 (O_2754,N_24684,N_24780);
or UO_2755 (O_2755,N_24814,N_24629);
xnor UO_2756 (O_2756,N_24908,N_24904);
xor UO_2757 (O_2757,N_24959,N_24737);
nand UO_2758 (O_2758,N_24709,N_24945);
and UO_2759 (O_2759,N_24786,N_24542);
nand UO_2760 (O_2760,N_24722,N_24843);
nand UO_2761 (O_2761,N_24759,N_24768);
or UO_2762 (O_2762,N_24818,N_24970);
xor UO_2763 (O_2763,N_24972,N_24586);
or UO_2764 (O_2764,N_24563,N_24590);
nand UO_2765 (O_2765,N_24799,N_24647);
xnor UO_2766 (O_2766,N_24936,N_24778);
nor UO_2767 (O_2767,N_24899,N_24875);
nand UO_2768 (O_2768,N_24723,N_24575);
and UO_2769 (O_2769,N_24606,N_24599);
and UO_2770 (O_2770,N_24688,N_24745);
or UO_2771 (O_2771,N_24671,N_24709);
and UO_2772 (O_2772,N_24554,N_24564);
and UO_2773 (O_2773,N_24753,N_24899);
or UO_2774 (O_2774,N_24687,N_24791);
and UO_2775 (O_2775,N_24956,N_24688);
xnor UO_2776 (O_2776,N_24952,N_24715);
nand UO_2777 (O_2777,N_24599,N_24664);
nand UO_2778 (O_2778,N_24670,N_24573);
nand UO_2779 (O_2779,N_24959,N_24783);
or UO_2780 (O_2780,N_24598,N_24781);
nor UO_2781 (O_2781,N_24618,N_24683);
or UO_2782 (O_2782,N_24760,N_24576);
nand UO_2783 (O_2783,N_24700,N_24857);
and UO_2784 (O_2784,N_24667,N_24857);
xor UO_2785 (O_2785,N_24836,N_24841);
or UO_2786 (O_2786,N_24728,N_24838);
nand UO_2787 (O_2787,N_24997,N_24807);
nor UO_2788 (O_2788,N_24735,N_24833);
or UO_2789 (O_2789,N_24601,N_24880);
nand UO_2790 (O_2790,N_24758,N_24918);
or UO_2791 (O_2791,N_24686,N_24842);
nor UO_2792 (O_2792,N_24865,N_24772);
xor UO_2793 (O_2793,N_24703,N_24645);
nand UO_2794 (O_2794,N_24794,N_24684);
xor UO_2795 (O_2795,N_24612,N_24969);
or UO_2796 (O_2796,N_24810,N_24643);
nand UO_2797 (O_2797,N_24782,N_24790);
xor UO_2798 (O_2798,N_24995,N_24976);
and UO_2799 (O_2799,N_24888,N_24626);
or UO_2800 (O_2800,N_24788,N_24758);
xor UO_2801 (O_2801,N_24964,N_24971);
or UO_2802 (O_2802,N_24572,N_24699);
nor UO_2803 (O_2803,N_24788,N_24994);
nor UO_2804 (O_2804,N_24559,N_24890);
xor UO_2805 (O_2805,N_24678,N_24561);
and UO_2806 (O_2806,N_24673,N_24932);
xnor UO_2807 (O_2807,N_24750,N_24571);
nor UO_2808 (O_2808,N_24965,N_24588);
or UO_2809 (O_2809,N_24707,N_24521);
or UO_2810 (O_2810,N_24648,N_24927);
or UO_2811 (O_2811,N_24928,N_24576);
xor UO_2812 (O_2812,N_24602,N_24970);
or UO_2813 (O_2813,N_24521,N_24616);
or UO_2814 (O_2814,N_24704,N_24923);
or UO_2815 (O_2815,N_24804,N_24983);
xor UO_2816 (O_2816,N_24773,N_24714);
and UO_2817 (O_2817,N_24991,N_24763);
nor UO_2818 (O_2818,N_24678,N_24934);
or UO_2819 (O_2819,N_24731,N_24952);
or UO_2820 (O_2820,N_24682,N_24957);
and UO_2821 (O_2821,N_24534,N_24692);
xor UO_2822 (O_2822,N_24658,N_24920);
nor UO_2823 (O_2823,N_24738,N_24873);
nand UO_2824 (O_2824,N_24526,N_24723);
nor UO_2825 (O_2825,N_24839,N_24818);
or UO_2826 (O_2826,N_24943,N_24916);
nand UO_2827 (O_2827,N_24633,N_24703);
and UO_2828 (O_2828,N_24888,N_24925);
and UO_2829 (O_2829,N_24633,N_24512);
nor UO_2830 (O_2830,N_24882,N_24636);
nand UO_2831 (O_2831,N_24976,N_24709);
or UO_2832 (O_2832,N_24787,N_24938);
and UO_2833 (O_2833,N_24528,N_24685);
nand UO_2834 (O_2834,N_24780,N_24831);
and UO_2835 (O_2835,N_24983,N_24866);
and UO_2836 (O_2836,N_24577,N_24902);
or UO_2837 (O_2837,N_24736,N_24747);
nand UO_2838 (O_2838,N_24902,N_24762);
or UO_2839 (O_2839,N_24929,N_24849);
nor UO_2840 (O_2840,N_24838,N_24720);
xor UO_2841 (O_2841,N_24985,N_24713);
xor UO_2842 (O_2842,N_24562,N_24528);
xor UO_2843 (O_2843,N_24813,N_24567);
and UO_2844 (O_2844,N_24717,N_24811);
nand UO_2845 (O_2845,N_24825,N_24896);
nand UO_2846 (O_2846,N_24750,N_24879);
and UO_2847 (O_2847,N_24997,N_24960);
nand UO_2848 (O_2848,N_24994,N_24853);
and UO_2849 (O_2849,N_24731,N_24982);
nand UO_2850 (O_2850,N_24833,N_24806);
or UO_2851 (O_2851,N_24939,N_24912);
or UO_2852 (O_2852,N_24848,N_24776);
and UO_2853 (O_2853,N_24636,N_24779);
xor UO_2854 (O_2854,N_24950,N_24770);
nor UO_2855 (O_2855,N_24962,N_24910);
nor UO_2856 (O_2856,N_24552,N_24561);
nand UO_2857 (O_2857,N_24587,N_24662);
nor UO_2858 (O_2858,N_24567,N_24895);
or UO_2859 (O_2859,N_24513,N_24935);
and UO_2860 (O_2860,N_24503,N_24658);
xnor UO_2861 (O_2861,N_24545,N_24656);
xor UO_2862 (O_2862,N_24910,N_24864);
nand UO_2863 (O_2863,N_24687,N_24861);
nor UO_2864 (O_2864,N_24783,N_24623);
or UO_2865 (O_2865,N_24561,N_24702);
nand UO_2866 (O_2866,N_24885,N_24557);
nand UO_2867 (O_2867,N_24850,N_24809);
nor UO_2868 (O_2868,N_24860,N_24689);
nor UO_2869 (O_2869,N_24814,N_24895);
nor UO_2870 (O_2870,N_24971,N_24942);
and UO_2871 (O_2871,N_24538,N_24995);
nor UO_2872 (O_2872,N_24837,N_24511);
nor UO_2873 (O_2873,N_24846,N_24836);
nand UO_2874 (O_2874,N_24698,N_24730);
and UO_2875 (O_2875,N_24819,N_24698);
or UO_2876 (O_2876,N_24973,N_24932);
xnor UO_2877 (O_2877,N_24700,N_24982);
nand UO_2878 (O_2878,N_24754,N_24747);
xor UO_2879 (O_2879,N_24858,N_24501);
or UO_2880 (O_2880,N_24945,N_24766);
nor UO_2881 (O_2881,N_24722,N_24986);
nor UO_2882 (O_2882,N_24804,N_24884);
xnor UO_2883 (O_2883,N_24861,N_24887);
and UO_2884 (O_2884,N_24519,N_24861);
xnor UO_2885 (O_2885,N_24717,N_24904);
and UO_2886 (O_2886,N_24710,N_24861);
or UO_2887 (O_2887,N_24541,N_24586);
nor UO_2888 (O_2888,N_24677,N_24957);
nand UO_2889 (O_2889,N_24669,N_24998);
or UO_2890 (O_2890,N_24617,N_24778);
xnor UO_2891 (O_2891,N_24988,N_24909);
nor UO_2892 (O_2892,N_24821,N_24990);
nor UO_2893 (O_2893,N_24713,N_24797);
or UO_2894 (O_2894,N_24716,N_24721);
and UO_2895 (O_2895,N_24967,N_24687);
or UO_2896 (O_2896,N_24683,N_24518);
xor UO_2897 (O_2897,N_24668,N_24853);
xor UO_2898 (O_2898,N_24832,N_24893);
and UO_2899 (O_2899,N_24601,N_24805);
nand UO_2900 (O_2900,N_24729,N_24865);
nor UO_2901 (O_2901,N_24688,N_24561);
xor UO_2902 (O_2902,N_24864,N_24961);
or UO_2903 (O_2903,N_24950,N_24830);
nor UO_2904 (O_2904,N_24697,N_24733);
nor UO_2905 (O_2905,N_24664,N_24984);
nor UO_2906 (O_2906,N_24556,N_24564);
nand UO_2907 (O_2907,N_24685,N_24566);
xor UO_2908 (O_2908,N_24508,N_24895);
nand UO_2909 (O_2909,N_24904,N_24874);
nor UO_2910 (O_2910,N_24977,N_24575);
and UO_2911 (O_2911,N_24763,N_24504);
nor UO_2912 (O_2912,N_24825,N_24809);
or UO_2913 (O_2913,N_24690,N_24673);
and UO_2914 (O_2914,N_24986,N_24754);
or UO_2915 (O_2915,N_24501,N_24932);
xnor UO_2916 (O_2916,N_24758,N_24846);
nand UO_2917 (O_2917,N_24668,N_24788);
and UO_2918 (O_2918,N_24543,N_24982);
nand UO_2919 (O_2919,N_24653,N_24906);
nand UO_2920 (O_2920,N_24949,N_24910);
nor UO_2921 (O_2921,N_24894,N_24957);
or UO_2922 (O_2922,N_24587,N_24610);
nand UO_2923 (O_2923,N_24630,N_24934);
xor UO_2924 (O_2924,N_24948,N_24543);
xor UO_2925 (O_2925,N_24603,N_24899);
xnor UO_2926 (O_2926,N_24928,N_24552);
xnor UO_2927 (O_2927,N_24620,N_24989);
nor UO_2928 (O_2928,N_24908,N_24945);
nand UO_2929 (O_2929,N_24870,N_24664);
or UO_2930 (O_2930,N_24662,N_24845);
nand UO_2931 (O_2931,N_24719,N_24976);
nor UO_2932 (O_2932,N_24897,N_24916);
xor UO_2933 (O_2933,N_24881,N_24544);
and UO_2934 (O_2934,N_24789,N_24792);
nand UO_2935 (O_2935,N_24558,N_24792);
and UO_2936 (O_2936,N_24725,N_24884);
xor UO_2937 (O_2937,N_24627,N_24737);
and UO_2938 (O_2938,N_24661,N_24964);
or UO_2939 (O_2939,N_24769,N_24698);
nor UO_2940 (O_2940,N_24678,N_24597);
or UO_2941 (O_2941,N_24679,N_24737);
xor UO_2942 (O_2942,N_24944,N_24760);
and UO_2943 (O_2943,N_24753,N_24939);
or UO_2944 (O_2944,N_24643,N_24555);
and UO_2945 (O_2945,N_24961,N_24682);
nand UO_2946 (O_2946,N_24743,N_24734);
nor UO_2947 (O_2947,N_24685,N_24547);
nand UO_2948 (O_2948,N_24908,N_24512);
and UO_2949 (O_2949,N_24720,N_24694);
or UO_2950 (O_2950,N_24995,N_24830);
nand UO_2951 (O_2951,N_24836,N_24601);
nor UO_2952 (O_2952,N_24590,N_24648);
nand UO_2953 (O_2953,N_24734,N_24909);
nand UO_2954 (O_2954,N_24881,N_24566);
nand UO_2955 (O_2955,N_24936,N_24779);
nor UO_2956 (O_2956,N_24596,N_24837);
nor UO_2957 (O_2957,N_24742,N_24701);
nor UO_2958 (O_2958,N_24883,N_24892);
nor UO_2959 (O_2959,N_24954,N_24527);
nand UO_2960 (O_2960,N_24695,N_24523);
and UO_2961 (O_2961,N_24934,N_24643);
xor UO_2962 (O_2962,N_24754,N_24787);
nor UO_2963 (O_2963,N_24534,N_24616);
nand UO_2964 (O_2964,N_24991,N_24622);
or UO_2965 (O_2965,N_24944,N_24756);
or UO_2966 (O_2966,N_24855,N_24812);
xnor UO_2967 (O_2967,N_24984,N_24781);
xor UO_2968 (O_2968,N_24570,N_24950);
xor UO_2969 (O_2969,N_24826,N_24680);
or UO_2970 (O_2970,N_24505,N_24562);
nor UO_2971 (O_2971,N_24776,N_24799);
nand UO_2972 (O_2972,N_24799,N_24568);
xor UO_2973 (O_2973,N_24500,N_24645);
or UO_2974 (O_2974,N_24764,N_24869);
nand UO_2975 (O_2975,N_24645,N_24985);
xor UO_2976 (O_2976,N_24650,N_24974);
nor UO_2977 (O_2977,N_24941,N_24657);
nor UO_2978 (O_2978,N_24922,N_24707);
or UO_2979 (O_2979,N_24733,N_24598);
nor UO_2980 (O_2980,N_24772,N_24622);
nand UO_2981 (O_2981,N_24601,N_24513);
nand UO_2982 (O_2982,N_24578,N_24592);
and UO_2983 (O_2983,N_24715,N_24693);
xor UO_2984 (O_2984,N_24707,N_24611);
nor UO_2985 (O_2985,N_24659,N_24607);
or UO_2986 (O_2986,N_24622,N_24603);
xor UO_2987 (O_2987,N_24539,N_24861);
xnor UO_2988 (O_2988,N_24988,N_24947);
nand UO_2989 (O_2989,N_24772,N_24975);
nand UO_2990 (O_2990,N_24882,N_24550);
nand UO_2991 (O_2991,N_24605,N_24621);
nor UO_2992 (O_2992,N_24808,N_24749);
and UO_2993 (O_2993,N_24674,N_24958);
nand UO_2994 (O_2994,N_24624,N_24908);
and UO_2995 (O_2995,N_24761,N_24536);
nor UO_2996 (O_2996,N_24595,N_24927);
or UO_2997 (O_2997,N_24655,N_24696);
xnor UO_2998 (O_2998,N_24739,N_24541);
xor UO_2999 (O_2999,N_24647,N_24695);
endmodule