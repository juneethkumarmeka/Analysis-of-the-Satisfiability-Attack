module basic_2000_20000_2500_80_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nor U0 (N_0,In_367,In_77);
or U1 (N_1,In_1841,In_1173);
and U2 (N_2,In_1600,In_440);
nor U3 (N_3,In_1679,In_530);
and U4 (N_4,In_1967,In_342);
xor U5 (N_5,In_138,In_810);
nor U6 (N_6,In_581,In_1309);
xor U7 (N_7,In_1869,In_1867);
nand U8 (N_8,In_165,In_573);
and U9 (N_9,In_593,In_932);
xor U10 (N_10,In_826,In_1279);
nor U11 (N_11,In_1217,In_1810);
or U12 (N_12,In_1731,In_1260);
and U13 (N_13,In_527,In_1349);
nor U14 (N_14,In_546,In_1901);
nand U15 (N_15,In_1857,In_0);
nor U16 (N_16,In_1456,In_1278);
xor U17 (N_17,In_852,In_53);
and U18 (N_18,In_897,In_1678);
or U19 (N_19,In_849,In_148);
nor U20 (N_20,In_1608,In_1680);
nand U21 (N_21,In_1740,In_1108);
and U22 (N_22,In_778,In_1658);
nor U23 (N_23,In_1671,In_719);
xnor U24 (N_24,In_644,In_1845);
xnor U25 (N_25,In_1933,In_1317);
nand U26 (N_26,In_667,In_943);
and U27 (N_27,In_1590,In_443);
xor U28 (N_28,In_510,In_1313);
xnor U29 (N_29,In_1609,In_566);
or U30 (N_30,In_36,In_609);
nand U31 (N_31,In_18,In_1395);
nand U32 (N_32,In_1846,In_1368);
and U33 (N_33,In_463,In_405);
and U34 (N_34,In_1993,In_1668);
nor U35 (N_35,In_1814,In_758);
nor U36 (N_36,In_1128,In_812);
nand U37 (N_37,In_258,In_1992);
or U38 (N_38,In_290,In_717);
or U39 (N_39,In_15,In_819);
xor U40 (N_40,In_1233,In_74);
nand U41 (N_41,In_1136,In_677);
or U42 (N_42,In_974,In_1161);
or U43 (N_43,In_1374,In_1423);
and U44 (N_44,In_547,In_265);
and U45 (N_45,In_1406,In_537);
xnor U46 (N_46,In_212,In_531);
nand U47 (N_47,In_1965,In_1477);
and U48 (N_48,In_733,In_95);
nand U49 (N_49,In_1842,In_1460);
or U50 (N_50,In_1515,In_1811);
nor U51 (N_51,In_1102,In_818);
nor U52 (N_52,In_172,In_459);
and U53 (N_53,In_655,In_1468);
nor U54 (N_54,In_596,In_1734);
and U55 (N_55,In_1311,In_1411);
and U56 (N_56,In_1934,In_1733);
nand U57 (N_57,In_355,In_1489);
or U58 (N_58,In_35,In_1649);
or U59 (N_59,In_642,In_1427);
xor U60 (N_60,In_1225,In_1794);
or U61 (N_61,In_615,In_1451);
nand U62 (N_62,In_1617,In_279);
or U63 (N_63,In_1470,In_217);
and U64 (N_64,In_311,In_242);
xnor U65 (N_65,In_1069,In_629);
xor U66 (N_66,In_1327,In_397);
and U67 (N_67,In_1359,In_1135);
or U68 (N_68,In_208,In_1772);
and U69 (N_69,In_1726,In_626);
nand U70 (N_70,In_1826,In_574);
nor U71 (N_71,In_772,In_1791);
or U72 (N_72,In_814,In_1756);
and U73 (N_73,In_557,In_293);
xnor U74 (N_74,In_1381,In_792);
nand U75 (N_75,In_1516,In_425);
xor U76 (N_76,In_916,In_1224);
nand U77 (N_77,In_622,In_1818);
xor U78 (N_78,In_1727,In_395);
nand U79 (N_79,In_8,In_503);
xnor U80 (N_80,In_479,In_748);
or U81 (N_81,In_1090,In_214);
nand U82 (N_82,In_283,In_1693);
or U83 (N_83,In_825,In_1026);
nand U84 (N_84,In_183,In_1481);
xnor U85 (N_85,In_222,In_882);
nor U86 (N_86,In_1333,In_422);
nor U87 (N_87,In_1780,In_653);
nor U88 (N_88,In_82,In_1796);
xnor U89 (N_89,In_1616,In_1152);
or U90 (N_90,In_1252,In_550);
xnor U91 (N_91,In_1474,In_756);
nor U92 (N_92,In_590,In_432);
nand U93 (N_93,In_1521,In_1554);
and U94 (N_94,In_853,In_669);
and U95 (N_95,In_1035,In_1005);
xor U96 (N_96,In_1212,In_860);
xor U97 (N_97,In_1452,In_1930);
or U98 (N_98,In_374,In_1736);
nand U99 (N_99,In_845,In_1358);
and U100 (N_100,In_406,In_181);
nand U101 (N_101,In_1016,In_972);
and U102 (N_102,In_1566,In_1899);
nor U103 (N_103,In_1601,In_450);
nor U104 (N_104,In_1294,In_1614);
nand U105 (N_105,In_1774,In_1355);
nor U106 (N_106,In_1769,In_1206);
or U107 (N_107,In_1729,In_666);
xnor U108 (N_108,In_1235,In_1234);
nor U109 (N_109,In_238,In_1540);
nor U110 (N_110,In_175,In_1564);
xnor U111 (N_111,In_34,In_426);
nand U112 (N_112,In_816,In_461);
nor U113 (N_113,In_817,In_1438);
nand U114 (N_114,In_60,In_914);
and U115 (N_115,In_160,In_1512);
and U116 (N_116,In_610,In_1963);
or U117 (N_117,In_995,In_1393);
and U118 (N_118,In_384,In_501);
or U119 (N_119,In_1689,In_1275);
nand U120 (N_120,In_670,In_131);
or U121 (N_121,In_1433,In_1493);
and U122 (N_122,In_1085,In_378);
and U123 (N_123,In_1262,In_266);
or U124 (N_124,In_1413,In_1179);
xor U125 (N_125,In_1730,In_1246);
and U126 (N_126,In_182,In_1805);
or U127 (N_127,In_1284,In_705);
and U128 (N_128,In_1367,In_998);
nand U129 (N_129,In_1043,In_672);
nor U130 (N_130,In_1952,In_1110);
nand U131 (N_131,In_81,In_1691);
and U132 (N_132,In_194,In_1175);
and U133 (N_133,In_1118,In_1463);
xnor U134 (N_134,In_875,In_568);
nor U135 (N_135,In_1595,In_920);
nor U136 (N_136,In_1760,In_1315);
or U137 (N_137,In_723,In_1364);
xnor U138 (N_138,In_1449,In_399);
nor U139 (N_139,In_392,In_1299);
nor U140 (N_140,In_1401,In_713);
xor U141 (N_141,In_1209,In_725);
nand U142 (N_142,In_971,In_321);
nor U143 (N_143,In_1793,In_534);
xnor U144 (N_144,In_1897,In_901);
nor U145 (N_145,In_75,In_1008);
or U146 (N_146,In_977,In_1995);
or U147 (N_147,In_136,In_13);
xor U148 (N_148,In_331,In_1076);
and U149 (N_149,In_1428,In_1854);
xor U150 (N_150,In_1775,In_1486);
xnor U151 (N_151,In_701,In_368);
nor U152 (N_152,In_144,In_125);
or U153 (N_153,In_1404,In_1322);
or U154 (N_154,In_1018,In_641);
or U155 (N_155,In_200,In_303);
or U156 (N_156,In_322,In_1487);
and U157 (N_157,In_1412,In_379);
nand U158 (N_158,In_827,In_218);
xnor U159 (N_159,In_1635,In_366);
and U160 (N_160,In_444,In_1661);
nand U161 (N_161,In_1319,In_1431);
xnor U162 (N_162,In_798,In_1205);
xnor U163 (N_163,In_1753,In_714);
nor U164 (N_164,In_1720,In_1886);
xor U165 (N_165,In_300,In_1361);
and U166 (N_166,In_577,In_895);
nor U167 (N_167,In_1125,In_11);
nand U168 (N_168,In_885,In_1271);
nand U169 (N_169,In_1265,In_813);
and U170 (N_170,In_260,In_1316);
nor U171 (N_171,In_970,In_967);
nand U172 (N_172,In_690,In_616);
nor U173 (N_173,In_1778,In_741);
or U174 (N_174,In_722,In_1338);
or U175 (N_175,In_1346,In_1488);
or U176 (N_176,In_963,In_1045);
or U177 (N_177,In_337,In_204);
nand U178 (N_178,In_559,In_1162);
and U179 (N_179,In_1898,In_12);
or U180 (N_180,In_309,In_1560);
nand U181 (N_181,In_1010,In_1865);
nor U182 (N_182,In_1697,In_1858);
nand U183 (N_183,In_1674,In_1894);
nand U184 (N_184,In_1593,In_800);
nand U185 (N_185,In_519,In_447);
nand U186 (N_186,In_1094,In_1256);
and U187 (N_187,In_1931,In_1415);
nor U188 (N_188,In_1220,In_1801);
nand U189 (N_189,In_319,In_1804);
xnor U190 (N_190,In_1061,In_1844);
and U191 (N_191,In_1054,In_1107);
or U192 (N_192,In_973,In_1436);
or U193 (N_193,In_1721,In_928);
nand U194 (N_194,In_1066,In_1392);
and U195 (N_195,In_1621,In_877);
nor U196 (N_196,In_1182,In_494);
or U197 (N_197,In_1064,In_1859);
and U198 (N_198,In_565,In_1650);
or U199 (N_199,In_1944,In_649);
nand U200 (N_200,In_1940,In_1149);
nand U201 (N_201,In_454,In_835);
xor U202 (N_202,In_1557,In_1973);
xor U203 (N_203,In_1191,In_31);
nor U204 (N_204,In_323,In_370);
nor U205 (N_205,In_1341,In_162);
and U206 (N_206,In_1887,In_548);
xor U207 (N_207,In_1027,In_1354);
or U208 (N_208,In_46,In_52);
xor U209 (N_209,In_1945,In_1360);
or U210 (N_210,In_312,In_621);
xnor U211 (N_211,In_1222,In_1444);
nand U212 (N_212,In_1214,In_1519);
xnor U213 (N_213,In_1350,In_1227);
nor U214 (N_214,In_1188,In_1267);
and U215 (N_215,In_567,In_1855);
nor U216 (N_216,In_1631,In_1868);
and U217 (N_217,In_591,In_960);
or U218 (N_218,In_1573,In_1571);
nand U219 (N_219,In_270,In_292);
xor U220 (N_220,In_1105,In_360);
xnor U221 (N_221,In_157,In_297);
nor U222 (N_222,In_839,In_564);
or U223 (N_223,In_939,In_1623);
nor U224 (N_224,In_1690,In_1592);
nor U225 (N_225,In_190,In_146);
or U226 (N_226,In_837,In_1822);
and U227 (N_227,In_1919,In_1408);
xnor U228 (N_228,In_783,In_1870);
nor U229 (N_229,In_497,In_1509);
xor U230 (N_230,In_1484,In_199);
or U231 (N_231,In_1371,In_1913);
nor U232 (N_232,In_770,In_418);
xor U233 (N_233,In_632,In_1335);
or U234 (N_234,In_1074,In_561);
or U235 (N_235,In_703,In_23);
and U236 (N_236,In_1770,In_1639);
or U237 (N_237,In_1885,In_504);
or U238 (N_238,In_1240,In_668);
nand U239 (N_239,In_883,In_539);
or U240 (N_240,In_1356,In_1168);
xnor U241 (N_241,In_1292,In_761);
or U242 (N_242,In_1834,In_1031);
xor U243 (N_243,In_417,In_773);
and U244 (N_244,In_1856,In_1537);
nand U245 (N_245,In_1565,In_1158);
nor U246 (N_246,In_535,In_377);
or U247 (N_247,In_1662,In_502);
xor U248 (N_248,In_624,In_1059);
nand U249 (N_249,In_1203,In_1763);
and U250 (N_250,In_365,In_1975);
nor U251 (N_251,In_514,In_1765);
or U252 (N_252,In_506,In_254);
nor U253 (N_253,In_1825,In_933);
or U254 (N_254,In_987,In_1542);
and U255 (N_255,In_1496,In_1130);
nor U256 (N_256,In_161,In_876);
nand U257 (N_257,In_1790,In_1871);
nand U258 (N_258,In_873,N_122);
or U259 (N_259,In_728,In_2);
and U260 (N_260,In_1029,In_1155);
nand U261 (N_261,In_1528,In_153);
xnor U262 (N_262,In_1098,In_976);
xnor U263 (N_263,In_129,In_1387);
and U264 (N_264,In_1004,In_1669);
or U265 (N_265,In_1644,In_509);
nor U266 (N_266,N_183,N_194);
nor U267 (N_267,In_526,In_1799);
and U268 (N_268,In_1802,In_373);
or U269 (N_269,N_80,In_1507);
and U270 (N_270,In_1171,N_103);
nand U271 (N_271,In_915,In_1088);
nor U272 (N_272,In_315,In_455);
xnor U273 (N_273,In_1620,In_648);
or U274 (N_274,In_1847,In_562);
and U275 (N_275,In_888,In_1425);
xor U276 (N_276,In_1437,In_1738);
xor U277 (N_277,In_1950,In_1123);
nand U278 (N_278,In_269,In_147);
and U279 (N_279,In_1699,In_1003);
or U280 (N_280,In_991,In_1792);
nand U281 (N_281,In_874,N_10);
xnor U282 (N_282,In_1403,N_16);
nor U283 (N_283,In_727,In_28);
or U284 (N_284,In_475,In_119);
or U285 (N_285,In_286,N_90);
and U286 (N_286,In_1563,In_1875);
or U287 (N_287,In_103,In_344);
xor U288 (N_288,In_706,In_468);
nor U289 (N_289,In_1109,In_571);
xor U290 (N_290,In_1638,In_1385);
nor U291 (N_291,In_1439,In_675);
or U292 (N_292,In_1971,In_352);
nand U293 (N_293,N_230,In_665);
nor U294 (N_294,In_1189,In_679);
or U295 (N_295,In_1572,In_1862);
nand U296 (N_296,In_805,In_334);
xor U297 (N_297,In_879,In_1972);
and U298 (N_298,In_1028,In_1747);
or U299 (N_299,In_1737,In_477);
or U300 (N_300,In_1126,In_1999);
and U301 (N_301,In_291,In_1688);
and U302 (N_302,In_1194,In_117);
and U303 (N_303,In_1798,In_786);
or U304 (N_304,In_797,In_955);
nand U305 (N_305,In_1597,In_1277);
or U306 (N_306,In_1526,In_1302);
nor U307 (N_307,In_1071,In_295);
or U308 (N_308,In_168,In_333);
xnor U309 (N_309,In_1352,In_804);
or U310 (N_310,In_1337,In_1707);
or U311 (N_311,In_1742,In_1207);
and U312 (N_312,In_42,N_121);
nor U313 (N_313,In_881,In_742);
nand U314 (N_314,In_1213,In_1215);
nor U315 (N_315,In_364,In_544);
nor U316 (N_316,N_223,In_339);
or U317 (N_317,In_942,In_802);
nor U318 (N_318,In_1583,N_109);
nand U319 (N_319,In_1612,N_130);
nor U320 (N_320,In_209,In_349);
xnor U321 (N_321,In_1911,In_1848);
nor U322 (N_322,In_1282,N_124);
nor U323 (N_323,In_1419,In_661);
nor U324 (N_324,In_828,In_611);
or U325 (N_325,In_1459,N_186);
nor U326 (N_326,In_328,In_986);
xor U327 (N_327,In_1698,In_684);
nor U328 (N_328,N_70,In_1369);
or U329 (N_329,In_1711,In_558);
nor U330 (N_330,In_1049,In_515);
xor U331 (N_331,In_132,In_445);
nand U332 (N_332,In_850,N_61);
nand U333 (N_333,In_167,N_224);
and U334 (N_334,In_7,N_178);
nor U335 (N_335,N_206,In_1286);
nand U336 (N_336,N_220,In_1396);
nand U337 (N_337,In_1497,In_985);
nor U338 (N_338,In_1466,In_1938);
nor U339 (N_339,In_587,In_840);
or U340 (N_340,In_1786,In_435);
nor U341 (N_341,In_710,In_40);
and U342 (N_342,In_1946,In_1676);
xnor U343 (N_343,In_1659,In_32);
and U344 (N_344,In_480,In_1099);
or U345 (N_345,In_1866,In_724);
or U346 (N_346,In_983,In_249);
nor U347 (N_347,In_551,In_1714);
and U348 (N_348,In_886,In_1231);
or U349 (N_349,In_1712,In_1181);
and U350 (N_350,In_124,In_631);
nand U351 (N_351,In_1190,In_793);
nand U352 (N_352,In_1131,In_380);
or U353 (N_353,In_411,In_841);
xnor U354 (N_354,In_122,In_1087);
or U355 (N_355,In_1186,In_1684);
xor U356 (N_356,In_1482,In_1208);
xor U357 (N_357,In_486,N_107);
and U358 (N_358,In_1011,In_702);
and U359 (N_359,In_1450,N_131);
nand U360 (N_360,In_1771,In_754);
nand U361 (N_361,In_1843,In_996);
and U362 (N_362,In_193,N_69);
or U363 (N_363,N_15,In_1091);
or U364 (N_364,N_199,In_1062);
nor U365 (N_365,In_434,In_899);
and U366 (N_366,N_191,N_165);
or U367 (N_367,N_13,In_1757);
and U368 (N_368,In_21,In_1932);
xor U369 (N_369,In_1293,In_1832);
xor U370 (N_370,N_192,In_940);
nor U371 (N_371,In_536,N_174);
nor U372 (N_372,In_1079,In_1545);
or U373 (N_373,In_19,In_1046);
and U374 (N_374,In_674,In_1250);
or U375 (N_375,In_647,In_471);
xor U376 (N_376,In_1178,In_708);
xnor U377 (N_377,N_120,In_1892);
nor U378 (N_378,In_1785,In_887);
nor U379 (N_379,In_1243,In_1270);
or U380 (N_380,N_111,In_1830);
or U381 (N_381,N_135,In_428);
nand U382 (N_382,In_149,In_51);
xor U383 (N_383,In_1910,N_221);
and U384 (N_384,In_1543,In_1308);
nand U385 (N_385,In_583,N_172);
nand U386 (N_386,In_1637,In_1782);
nor U387 (N_387,In_1296,In_1550);
nand U388 (N_388,In_1642,In_739);
nor U389 (N_389,In_1127,In_1954);
nand U390 (N_390,N_217,In_1148);
nor U391 (N_391,In_580,In_313);
nor U392 (N_392,In_1274,In_211);
or U393 (N_393,In_634,In_599);
nand U394 (N_394,N_100,In_187);
nand U395 (N_395,In_401,In_1219);
nor U396 (N_396,In_1902,In_989);
and U397 (N_397,In_1210,In_469);
or U398 (N_398,In_90,In_650);
nor U399 (N_399,In_1514,In_1473);
nor U400 (N_400,In_906,In_811);
nor U401 (N_401,In_1112,In_1922);
nand U402 (N_402,In_362,In_969);
and U403 (N_403,N_247,In_738);
xor U404 (N_404,In_1159,N_83);
nor U405 (N_405,In_905,In_1295);
and U406 (N_406,In_700,N_36);
xor U407 (N_407,In_1229,N_118);
nor U408 (N_408,In_597,In_58);
xor U409 (N_409,In_934,In_1430);
xnor U410 (N_410,N_88,In_251);
and U411 (N_411,In_1465,In_1570);
and U412 (N_412,N_242,In_1618);
nand U413 (N_413,In_1000,In_1863);
or U414 (N_414,In_163,In_437);
and U415 (N_415,In_1912,N_38);
and U416 (N_416,In_1255,In_1705);
nor U417 (N_417,In_576,In_66);
nand U418 (N_418,In_902,In_1718);
nand U419 (N_419,In_1665,In_72);
nor U420 (N_420,In_1978,In_782);
or U421 (N_421,In_1204,In_169);
nand U422 (N_422,In_1551,In_436);
or U423 (N_423,In_575,In_1585);
xor U424 (N_424,In_1323,In_357);
or U425 (N_425,In_330,In_1837);
or U426 (N_426,In_603,In_284);
xnor U427 (N_427,In_1390,N_92);
or U428 (N_428,In_1926,In_809);
and U429 (N_429,In_711,In_171);
and U430 (N_430,In_1667,N_91);
and U431 (N_431,In_929,In_900);
and U432 (N_432,In_636,In_1629);
and U433 (N_433,In_1373,In_1084);
or U434 (N_434,In_1921,In_847);
nor U435 (N_435,In_1532,In_912);
xnor U436 (N_436,In_1339,In_277);
xnor U437 (N_437,N_60,In_78);
nand U438 (N_438,In_215,N_226);
xnor U439 (N_439,In_1056,N_175);
and U440 (N_440,In_186,In_1675);
nor U441 (N_441,In_1717,In_638);
nor U442 (N_442,N_51,N_33);
and U443 (N_443,In_1997,In_361);
and U444 (N_444,N_105,N_64);
xnor U445 (N_445,In_414,In_1372);
nor U446 (N_446,N_67,In_937);
nor U447 (N_447,In_413,N_167);
xor U448 (N_448,In_838,In_619);
xor U449 (N_449,In_1998,In_1510);
and U450 (N_450,In_25,In_359);
and U451 (N_451,In_1023,In_320);
and U452 (N_452,In_1682,In_855);
xnor U453 (N_453,In_388,In_1677);
nor U454 (N_454,In_1388,In_1695);
nor U455 (N_455,In_255,In_304);
nor U456 (N_456,N_23,In_263);
nand U457 (N_457,In_1024,N_189);
xnor U458 (N_458,In_1119,In_1523);
nor U459 (N_459,In_354,N_72);
or U460 (N_460,In_452,In_1336);
nand U461 (N_461,In_87,In_780);
or U462 (N_462,In_944,In_524);
nand U463 (N_463,In_1896,In_244);
nor U464 (N_464,N_238,In_472);
xor U465 (N_465,In_302,In_743);
and U466 (N_466,In_1363,In_1378);
nand U467 (N_467,In_549,In_498);
xor U468 (N_468,In_1139,In_1643);
xnor U469 (N_469,In_1903,In_842);
nor U470 (N_470,In_1582,In_822);
nand U471 (N_471,In_24,In_1351);
and U472 (N_472,In_981,In_438);
and U473 (N_473,In_1872,In_1513);
nand U474 (N_474,In_441,In_1710);
and U475 (N_475,In_820,In_219);
or U476 (N_476,In_1495,In_1983);
nand U477 (N_477,In_1610,In_521);
nor U478 (N_478,N_25,In_1535);
xnor U479 (N_479,In_488,N_54);
nor U480 (N_480,In_326,In_736);
nand U481 (N_481,In_1097,In_1143);
or U482 (N_482,In_821,In_1244);
and U483 (N_483,In_85,In_239);
nor U484 (N_484,In_846,In_715);
xnor U485 (N_485,In_1506,In_1657);
xor U486 (N_486,In_1957,In_1548);
nor U487 (N_487,In_63,In_33);
nor U488 (N_488,In_578,In_71);
or U489 (N_489,In_1701,N_89);
or U490 (N_490,In_1559,In_1732);
nor U491 (N_491,In_271,In_1176);
xnor U492 (N_492,In_262,In_1673);
nor U493 (N_493,N_26,In_478);
or U494 (N_494,In_628,In_779);
xnor U495 (N_495,In_1067,In_1305);
nand U496 (N_496,In_294,In_999);
xnor U497 (N_497,In_843,In_1254);
nor U498 (N_498,In_962,In_1281);
nor U499 (N_499,In_861,In_1929);
and U500 (N_500,In_1259,In_353);
and U501 (N_501,N_288,In_1410);
and U502 (N_502,N_257,In_1195);
and U503 (N_503,In_784,In_108);
and U504 (N_504,In_993,In_1539);
nor U505 (N_505,In_55,In_1121);
and U506 (N_506,In_99,In_716);
nand U507 (N_507,N_234,N_251);
and U508 (N_508,In_747,In_1201);
nand U509 (N_509,In_652,N_465);
nand U510 (N_510,N_438,In_1223);
or U511 (N_511,N_255,In_1956);
or U512 (N_512,In_1226,In_921);
xnor U513 (N_513,In_1604,N_293);
and U514 (N_514,N_56,In_1719);
and U515 (N_515,In_1266,In_1051);
nor U516 (N_516,In_1264,In_1402);
xor U517 (N_517,In_1587,In_253);
or U518 (N_518,In_685,N_126);
and U519 (N_519,In_823,In_495);
xor U520 (N_520,In_1095,N_466);
nor U521 (N_521,In_1883,N_346);
nor U522 (N_522,In_836,In_683);
nand U523 (N_523,In_423,In_662);
or U524 (N_524,In_155,N_281);
nand U525 (N_525,In_1146,In_1928);
nand U526 (N_526,In_1605,N_381);
nand U527 (N_527,In_130,N_96);
or U528 (N_528,In_296,In_340);
or U529 (N_529,In_1253,In_1328);
nand U530 (N_530,In_1672,In_1647);
or U531 (N_531,In_1384,In_1664);
nor U532 (N_532,In_1906,In_1248);
or U533 (N_533,In_1598,In_1777);
nor U534 (N_534,In_1479,In_1421);
and U535 (N_535,In_381,N_340);
nor U536 (N_536,N_98,In_1216);
nand U537 (N_537,In_1429,In_1300);
nor U538 (N_538,In_1820,In_1416);
nand U539 (N_539,In_1925,N_433);
and U540 (N_540,In_1398,In_595);
nor U541 (N_541,In_1947,In_1498);
xnor U542 (N_542,N_401,N_337);
or U543 (N_543,In_1636,N_68);
nand U544 (N_544,In_98,In_1426);
nor U545 (N_545,N_81,In_633);
nor U546 (N_546,In_17,In_1063);
or U547 (N_547,In_1133,In_348);
and U548 (N_548,In_493,In_1057);
nand U549 (N_549,In_1307,In_1376);
and U550 (N_550,In_966,In_734);
nor U551 (N_551,N_17,In_287);
nor U552 (N_552,In_1122,In_1891);
and U553 (N_553,N_269,In_604);
nand U554 (N_554,N_304,In_1918);
nand U555 (N_555,In_57,In_1407);
nor U556 (N_556,N_260,In_910);
nor U557 (N_557,In_1036,N_106);
and U558 (N_558,In_1042,In_1058);
nor U559 (N_559,N_338,In_1821);
or U560 (N_560,N_349,N_405);
nor U561 (N_561,In_1986,In_990);
nor U562 (N_562,In_630,N_59);
nor U563 (N_563,In_113,In_1283);
and U564 (N_564,N_378,In_1218);
nor U565 (N_565,In_660,N_457);
nand U566 (N_566,In_483,In_1602);
nor U567 (N_567,In_145,N_279);
nor U568 (N_568,In_1116,N_187);
or U569 (N_569,In_1704,In_29);
xnor U570 (N_570,In_317,In_120);
and U571 (N_571,In_372,N_400);
nand U572 (N_572,In_1312,N_404);
nor U573 (N_573,In_1574,In_485);
xor U574 (N_574,In_48,In_1709);
xnor U575 (N_575,N_263,In_941);
xnor U576 (N_576,In_729,In_848);
nor U577 (N_577,In_1124,In_1047);
xnor U578 (N_578,In_949,N_147);
or U579 (N_579,In_1494,In_500);
xnor U580 (N_580,N_45,In_431);
nor U581 (N_581,In_1746,In_1800);
or U582 (N_582,N_403,In_47);
nor U583 (N_583,In_1290,N_460);
nor U584 (N_584,In_1014,In_83);
xor U585 (N_585,In_1020,In_1624);
and U586 (N_586,In_1483,In_1441);
or U587 (N_587,N_355,In_97);
xnor U588 (N_588,In_1163,N_39);
or U589 (N_589,N_440,N_411);
nand U590 (N_590,In_476,N_275);
nor U591 (N_591,N_375,N_27);
and U592 (N_592,N_197,In_749);
nor U593 (N_593,In_1948,In_1784);
or U594 (N_594,In_1663,In_1819);
and U595 (N_595,In_600,In_791);
nand U596 (N_596,In_541,In_1078);
nor U597 (N_597,In_1435,In_1666);
and U598 (N_598,In_1228,In_1619);
nand U599 (N_599,In_1142,N_454);
and U600 (N_600,In_764,N_6);
nor U601 (N_601,In_1959,In_408);
nand U602 (N_602,In_1976,In_907);
and U603 (N_603,In_639,N_41);
nand U604 (N_604,N_373,N_452);
nor U605 (N_605,N_322,N_149);
nand U606 (N_606,N_262,In_612);
and U607 (N_607,In_865,In_245);
nand U608 (N_608,In_1382,In_1851);
or U609 (N_609,In_112,In_1007);
nor U610 (N_610,N_212,N_443);
or U611 (N_611,N_309,In_267);
xnor U612 (N_612,N_156,In_1237);
xnor U613 (N_613,In_489,In_273);
nor U614 (N_614,In_980,In_1331);
and U615 (N_615,In_1873,In_227);
or U616 (N_616,In_202,In_1626);
xor U617 (N_617,N_79,In_1797);
or U618 (N_618,In_1242,In_935);
xor U619 (N_619,In_195,In_682);
or U620 (N_620,In_673,In_737);
nor U621 (N_621,N_152,In_1996);
nor U622 (N_622,In_1092,In_698);
nor U623 (N_623,In_1968,In_115);
xor U624 (N_624,In_73,N_213);
nand U625 (N_625,In_419,In_688);
nor U626 (N_626,In_1781,In_257);
and U627 (N_627,In_803,N_362);
nand U628 (N_628,In_948,In_1198);
nand U629 (N_629,In_1471,In_1807);
xnor U630 (N_630,N_134,In_1457);
or U631 (N_631,In_170,In_1692);
or U632 (N_632,In_1916,In_1320);
nor U633 (N_633,N_424,In_329);
nor U634 (N_634,In_1878,In_275);
nor U635 (N_635,In_781,N_299);
nor U636 (N_636,In_1113,In_1594);
and U637 (N_637,In_529,In_868);
nor U638 (N_638,In_201,In_532);
xnor U639 (N_639,In_1951,In_50);
xnor U640 (N_640,In_243,In_65);
nor U641 (N_641,In_110,In_1081);
xnor U642 (N_642,N_436,In_1455);
or U643 (N_643,In_420,In_210);
and U644 (N_644,N_57,In_801);
xnor U645 (N_645,In_229,In_1655);
xnor U646 (N_646,N_426,N_65);
nor U647 (N_647,In_1890,In_191);
nand U648 (N_648,N_233,N_352);
and U649 (N_649,In_740,In_1779);
nor U650 (N_650,N_451,N_133);
xor U651 (N_651,N_188,In_1703);
or U652 (N_652,N_369,In_336);
nor U653 (N_653,In_299,N_480);
xor U654 (N_654,N_303,N_368);
and U655 (N_655,N_43,In_1030);
and U656 (N_656,In_520,In_393);
nand U657 (N_657,In_1860,In_686);
xor U658 (N_658,In_1467,In_1783);
xnor U659 (N_659,N_385,In_750);
and U660 (N_660,N_244,N_252);
nor U661 (N_661,In_1065,In_233);
nand U662 (N_662,In_1070,In_1882);
nand U663 (N_663,In_1584,N_473);
xnor U664 (N_664,In_1633,In_1909);
nor U665 (N_665,In_917,N_161);
nand U666 (N_666,In_1400,In_1157);
and U667 (N_667,In_1538,N_40);
and U668 (N_668,In_625,N_361);
nand U669 (N_669,In_453,In_281);
or U670 (N_670,In_1370,N_210);
nor U671 (N_671,N_332,In_256);
xnor U672 (N_672,In_56,In_1745);
nand U673 (N_673,N_432,N_289);
nand U674 (N_674,In_114,N_356);
nand U675 (N_675,N_231,In_1138);
and U676 (N_676,N_138,In_627);
nand U677 (N_677,N_391,In_1634);
and U678 (N_678,N_18,N_136);
nor U679 (N_679,In_456,N_225);
nor U680 (N_680,In_88,In_1174);
and U681 (N_681,In_704,In_1006);
nand U682 (N_682,In_982,In_1599);
or U683 (N_683,In_451,In_1586);
nor U684 (N_684,In_1681,In_1329);
nand U685 (N_685,In_369,N_487);
nand U686 (N_686,N_209,In_795);
and U687 (N_687,In_1491,N_296);
and U688 (N_688,In_556,N_498);
nand U689 (N_689,N_148,In_1589);
xnor U690 (N_690,In_936,In_45);
nand U691 (N_691,In_908,In_1485);
nor U692 (N_692,N_58,In_1838);
nand U693 (N_693,N_292,In_1504);
nor U694 (N_694,In_176,N_78);
nor U695 (N_695,In_975,N_229);
and U696 (N_696,In_104,In_261);
or U697 (N_697,In_552,In_1447);
nand U698 (N_698,N_19,N_484);
nand U699 (N_699,In_854,N_151);
and U700 (N_700,N_101,In_1200);
nor U701 (N_701,N_447,In_1257);
xnor U702 (N_702,In_984,In_755);
or U703 (N_703,N_1,N_259);
nand U704 (N_704,In_1015,In_1789);
nand U705 (N_705,N_497,N_265);
xor U706 (N_706,N_285,N_448);
xnor U707 (N_707,In_586,In_1375);
and U708 (N_708,In_1839,In_1552);
or U709 (N_709,N_222,In_1480);
xnor U710 (N_710,N_218,N_395);
and U711 (N_711,N_422,In_1330);
or U712 (N_712,In_1787,In_1141);
or U713 (N_713,In_1297,N_351);
nor U714 (N_714,In_232,In_1961);
xnor U715 (N_715,In_484,N_44);
and U716 (N_716,N_184,In_1713);
nor U717 (N_717,In_1432,In_1773);
nand U718 (N_718,In_1722,In_862);
or U719 (N_719,In_492,In_241);
nand U720 (N_720,In_988,N_55);
or U721 (N_721,In_449,N_308);
nand U722 (N_722,In_133,N_393);
nand U723 (N_723,In_893,In_1549);
nor U724 (N_724,N_14,In_1580);
and U725 (N_725,In_1478,N_287);
and U726 (N_726,N_494,In_1974);
nor U727 (N_727,N_52,N_48);
and U728 (N_728,N_328,In_1357);
or U729 (N_729,In_371,In_1652);
or U730 (N_730,In_487,In_1966);
or U731 (N_731,In_1759,N_358);
or U732 (N_732,In_387,In_508);
nor U733 (N_733,In_226,N_376);
nand U734 (N_734,In_152,N_345);
nor U735 (N_735,In_1039,In_325);
and U736 (N_736,In_1405,In_1247);
nor U737 (N_737,In_1117,In_102);
nand U738 (N_738,In_156,N_482);
and U739 (N_739,In_1353,In_1083);
xnor U740 (N_740,In_439,In_1280);
xnor U741 (N_741,In_718,In_1632);
nor U742 (N_742,In_579,N_250);
xor U743 (N_743,In_1980,N_301);
and U744 (N_744,N_267,In_1568);
or U745 (N_745,In_474,In_345);
nor U746 (N_746,In_1490,In_26);
or U747 (N_747,N_145,In_1531);
and U748 (N_748,In_856,N_62);
xor U749 (N_749,In_554,N_93);
nor U750 (N_750,N_413,In_16);
and U751 (N_751,N_291,N_402);
nand U752 (N_752,N_163,N_619);
and U753 (N_753,N_215,In_513);
xor U754 (N_754,N_294,N_414);
nor U755 (N_755,N_169,In_466);
or U756 (N_756,In_678,In_1755);
or U757 (N_757,In_694,N_560);
nor U758 (N_758,N_568,N_573);
nor U759 (N_759,In_1365,In_1272);
and U760 (N_760,N_672,In_1881);
and U761 (N_761,In_44,N_82);
nor U762 (N_762,N_331,N_286);
xnor U763 (N_763,In_909,In_752);
and U764 (N_764,In_385,In_282);
and U765 (N_765,N_665,N_495);
or U766 (N_766,N_599,N_656);
and U767 (N_767,In_1022,In_1383);
nand U768 (N_768,N_73,N_531);
and U769 (N_769,N_282,In_1879);
and U770 (N_770,In_618,In_871);
and U771 (N_771,In_1166,In_1055);
and U772 (N_772,In_391,In_1012);
or U773 (N_773,In_1628,In_1962);
nor U774 (N_774,In_116,N_581);
xor U775 (N_775,N_77,In_1749);
xor U776 (N_776,N_335,N_701);
nand U777 (N_777,N_9,In_1541);
or U778 (N_778,In_1261,In_1603);
xor U779 (N_779,In_1301,N_97);
nand U780 (N_780,N_412,N_99);
and U781 (N_781,N_445,In_1660);
nor U782 (N_782,In_957,In_1344);
or U783 (N_783,In_1106,In_1025);
nor U784 (N_784,N_84,In_400);
and U785 (N_785,In_775,N_205);
and U786 (N_786,In_1907,In_1500);
and U787 (N_787,N_601,N_663);
nor U788 (N_788,N_712,N_694);
nand U789 (N_789,In_1522,In_1380);
nor U790 (N_790,In_867,In_410);
and U791 (N_791,In_1314,In_851);
xnor U792 (N_792,N_614,N_745);
nor U793 (N_793,In_61,N_439);
and U794 (N_794,In_421,N_50);
nor U795 (N_795,In_1806,N_662);
and U796 (N_796,In_1446,In_196);
nor U797 (N_797,In_913,In_1132);
xor U798 (N_798,N_713,In_1391);
and U799 (N_799,In_1562,N_651);
or U800 (N_800,N_731,In_207);
and U801 (N_801,N_707,N_462);
nor U802 (N_802,In_1553,In_1183);
nor U803 (N_803,In_806,In_27);
nand U804 (N_804,N_579,N_566);
xnor U805 (N_805,In_1761,N_314);
or U806 (N_806,In_415,In_1192);
and U807 (N_807,N_668,In_992);
or U808 (N_808,N_645,In_206);
nand U809 (N_809,In_605,In_646);
nand U810 (N_810,N_699,In_216);
or U811 (N_811,In_496,In_252);
and U812 (N_812,In_796,In_1386);
and U813 (N_813,In_1040,N_114);
and U814 (N_814,In_1615,N_610);
or U815 (N_815,N_545,In_1288);
nor U816 (N_816,In_76,N_297);
and U817 (N_817,In_318,N_357);
xnor U818 (N_818,In_1795,N_730);
nor U819 (N_819,In_10,In_880);
or U820 (N_820,N_425,In_278);
xor U821 (N_821,In_952,In_903);
nand U822 (N_822,N_363,In_1418);
xor U823 (N_823,In_1185,In_1348);
or U824 (N_824,N_214,N_526);
xor U825 (N_825,In_1520,In_128);
and U826 (N_826,In_164,In_1741);
or U827 (N_827,In_613,In_869);
nor U828 (N_828,In_1694,N_453);
nand U829 (N_829,N_348,N_571);
nor U830 (N_830,In_904,N_446);
xor U831 (N_831,In_59,N_360);
or U832 (N_832,N_196,In_1829);
xor U833 (N_833,N_729,In_606);
or U834 (N_834,N_529,In_1808);
nand U835 (N_835,N_537,N_724);
nand U836 (N_836,In_68,In_1960);
or U837 (N_837,In_89,N_502);
xnor U838 (N_838,N_557,N_585);
xnor U839 (N_839,In_922,In_1145);
xnor U840 (N_840,N_638,In_1347);
xor U841 (N_841,In_664,In_1137);
nor U842 (N_842,In_830,N_697);
xor U843 (N_843,In_1101,N_632);
nor U844 (N_844,In_1861,N_146);
xnor U845 (N_845,In_1306,N_570);
and U846 (N_846,In_1706,N_3);
nor U847 (N_847,N_524,N_116);
or U848 (N_848,In_1342,N_559);
xor U849 (N_849,In_829,N_661);
nand U850 (N_850,N_598,In_687);
or U851 (N_851,In_1180,In_1230);
or U852 (N_852,In_1167,In_517);
and U853 (N_853,In_490,In_1424);
nor U854 (N_854,In_512,In_1461);
and U855 (N_855,In_891,N_544);
and U856 (N_856,N_696,N_266);
xnor U857 (N_857,In_223,In_753);
and U858 (N_858,N_491,In_1533);
nand U859 (N_859,N_475,In_1285);
xor U860 (N_860,N_676,In_220);
and U861 (N_861,N_474,In_777);
or U862 (N_862,N_682,N_505);
or U863 (N_863,In_1762,In_1394);
or U864 (N_864,In_767,In_1970);
or U865 (N_865,In_1249,In_166);
xor U866 (N_866,N_123,In_268);
nor U867 (N_867,In_997,In_280);
and U868 (N_868,N_164,N_660);
and U869 (N_869,In_1518,N_407);
xor U870 (N_870,In_978,N_507);
or U871 (N_871,N_132,In_1888);
nor U872 (N_872,N_622,In_884);
nor U873 (N_873,N_590,In_950);
nor U874 (N_874,N_323,In_91);
nor U875 (N_875,N_166,N_386);
or U876 (N_876,N_721,In_776);
or U877 (N_877,In_1754,In_1768);
nand U878 (N_878,N_549,N_155);
nor U879 (N_879,N_515,In_1434);
or U880 (N_880,N_374,N_305);
xor U881 (N_881,In_351,In_1588);
or U882 (N_882,In_1464,In_744);
and U883 (N_883,In_695,In_1915);
or U884 (N_884,In_1824,In_228);
nand U885 (N_885,In_308,N_12);
and U886 (N_886,N_236,In_1715);
nor U887 (N_887,In_964,N_653);
and U888 (N_888,N_539,N_483);
nand U889 (N_889,N_720,N_420);
nand U890 (N_890,In_205,N_290);
nand U891 (N_891,In_1752,In_246);
and U892 (N_892,N_596,In_457);
xnor U893 (N_893,In_335,In_1569);
nand U894 (N_894,N_567,N_383);
nand U895 (N_895,In_350,In_3);
and U896 (N_896,In_314,In_858);
nor U897 (N_897,In_1558,N_329);
nand U898 (N_898,N_141,In_726);
nor U899 (N_899,In_735,N_717);
and U900 (N_900,In_1544,In_106);
nor U901 (N_901,In_1263,N_158);
nor U902 (N_902,In_1082,N_584);
nand U903 (N_903,In_572,In_844);
xnor U904 (N_904,In_1268,N_688);
nor U905 (N_905,In_953,N_182);
nor U906 (N_906,In_123,In_1987);
nor U907 (N_907,N_399,In_1546);
nand U908 (N_908,In_358,N_464);
xnor U909 (N_909,In_1197,N_747);
or U910 (N_910,In_1900,In_745);
and U911 (N_911,In_1221,In_416);
xor U912 (N_912,In_225,In_184);
nor U913 (N_913,N_684,N_2);
nand U914 (N_914,In_1575,N_71);
nand U915 (N_915,In_403,N_419);
or U916 (N_916,N_42,In_1093);
or U917 (N_917,In_1077,In_394);
xor U918 (N_918,N_591,In_1303);
or U919 (N_919,In_306,In_1828);
or U920 (N_920,In_1,In_1454);
and U921 (N_921,In_589,In_1310);
nand U922 (N_922,N_655,In_1475);
nand U923 (N_923,N_207,N_551);
nand U924 (N_924,In_1239,In_994);
or U925 (N_925,In_555,In_1001);
nand U926 (N_926,In_1815,N_648);
nor U927 (N_927,In_896,In_307);
nor U928 (N_928,In_732,In_712);
nor U929 (N_929,N_102,N_430);
and U930 (N_930,In_866,N_434);
xnor U931 (N_931,In_1534,N_112);
or U932 (N_932,In_918,In_607);
nor U933 (N_933,N_623,In_41);
and U934 (N_934,N_37,N_738);
and U935 (N_935,N_637,In_1038);
nand U936 (N_936,In_1567,In_481);
xor U937 (N_937,N_703,In_465);
and U938 (N_938,In_327,N_298);
nor U939 (N_939,In_1577,N_396);
nand U940 (N_940,In_1269,N_521);
nor U941 (N_941,N_125,In_832);
nand U942 (N_942,In_1505,In_766);
and U943 (N_943,In_1687,N_193);
nand U944 (N_944,N_734,In_1927);
nor U945 (N_945,In_1080,N_737);
and U946 (N_946,N_216,In_62);
xor U947 (N_947,N_20,In_878);
and U948 (N_948,In_720,In_1321);
xor U949 (N_949,N_256,In_1529);
and U950 (N_950,In_1556,In_1591);
and U951 (N_951,N_75,In_189);
and U952 (N_952,In_1114,In_1625);
nand U953 (N_953,In_1153,N_504);
or U954 (N_954,In_142,In_926);
xnor U955 (N_955,In_769,N_24);
or U956 (N_956,In_954,In_1991);
or U957 (N_957,In_608,N_389);
nand U958 (N_958,In_1469,In_696);
nor U959 (N_959,N_540,N_277);
or U960 (N_960,In_1377,In_341);
nand U961 (N_961,In_127,In_923);
and U962 (N_962,In_1735,N_429);
and U963 (N_963,In_1723,N_284);
or U964 (N_964,N_364,In_1648);
or U965 (N_965,In_298,In_1273);
and U966 (N_966,In_137,In_588);
xor U967 (N_967,In_1724,N_21);
or U968 (N_968,N_576,N_550);
and U969 (N_969,In_301,N_527);
or U970 (N_970,In_1073,N_104);
or U971 (N_971,In_1803,In_1630);
and U972 (N_972,N_608,N_325);
nand U973 (N_973,N_488,N_273);
nand U974 (N_974,In_746,N_85);
nor U975 (N_975,In_788,In_158);
xor U976 (N_976,In_560,In_1696);
or U977 (N_977,In_1836,In_592);
xnor U978 (N_978,In_1096,In_1645);
xor U979 (N_979,N_652,N_667);
and U980 (N_980,N_586,N_461);
or U981 (N_981,In_389,N_377);
or U982 (N_982,N_245,N_654);
nor U983 (N_983,In_39,In_890);
and U984 (N_984,In_264,In_470);
and U985 (N_985,N_736,N_458);
and U986 (N_986,N_735,In_1686);
nand U987 (N_987,In_1202,In_141);
xnor U988 (N_988,In_1499,N_31);
and U989 (N_989,N_235,N_371);
xnor U990 (N_990,In_1060,In_1530);
xnor U991 (N_991,In_111,In_1670);
xnor U992 (N_992,N_716,N_536);
nor U993 (N_993,N_137,In_1864);
nand U994 (N_994,In_671,In_1935);
or U995 (N_995,N_392,In_958);
or U996 (N_996,In_429,In_1576);
or U997 (N_997,N_321,In_1611);
nor U998 (N_998,In_20,In_947);
or U999 (N_999,In_150,N_493);
nor U1000 (N_1000,In_709,In_1895);
and U1001 (N_1001,In_1750,In_951);
and U1002 (N_1002,In_1581,In_1017);
nor U1003 (N_1003,N_950,N_516);
and U1004 (N_1004,In_1748,N_949);
xnor U1005 (N_1005,In_347,In_1725);
or U1006 (N_1006,N_508,N_201);
xor U1007 (N_1007,N_844,N_5);
or U1008 (N_1008,In_857,In_1289);
nor U1009 (N_1009,In_96,In_424);
xnor U1010 (N_1010,N_975,In_1656);
or U1011 (N_1011,N_784,In_1251);
nand U1012 (N_1012,N_22,In_491);
xnor U1013 (N_1013,In_1536,N_477);
and U1014 (N_1014,N_316,N_562);
nand U1015 (N_1015,In_1527,N_63);
and U1016 (N_1016,In_1298,N_94);
or U1017 (N_1017,N_967,N_689);
nor U1018 (N_1018,N_558,N_589);
and U1019 (N_1019,N_799,N_302);
or U1020 (N_1020,N_489,N_517);
xor U1021 (N_1021,N_179,N_958);
or U1022 (N_1022,N_594,N_865);
nand U1023 (N_1023,N_326,In_831);
nor U1024 (N_1024,N_384,N_394);
xnor U1025 (N_1025,N_846,In_1032);
or U1026 (N_1026,In_221,N_832);
xor U1027 (N_1027,N_990,N_750);
or U1028 (N_1028,N_634,N_115);
xnor U1029 (N_1029,N_370,N_597);
or U1030 (N_1030,In_30,N_828);
and U1031 (N_1031,In_693,N_367);
nand U1032 (N_1032,N_319,N_441);
nand U1033 (N_1033,In_467,N_856);
nand U1034 (N_1034,N_850,N_605);
nor U1035 (N_1035,N_128,In_224);
nand U1036 (N_1036,In_965,N_630);
and U1037 (N_1037,N_911,N_624);
or U1038 (N_1038,N_867,N_897);
xor U1039 (N_1039,N_794,In_1276);
nand U1040 (N_1040,N_899,N_278);
nor U1041 (N_1041,N_757,In_248);
or U1042 (N_1042,N_556,In_505);
or U1043 (N_1043,N_449,In_105);
nor U1044 (N_1044,N_427,N_631);
and U1045 (N_1045,In_1685,N_330);
nor U1046 (N_1046,N_615,N_948);
nand U1047 (N_1047,In_1964,N_779);
xor U1048 (N_1048,In_1111,In_1445);
or U1049 (N_1049,In_623,In_1379);
nor U1050 (N_1050,N_324,N_765);
or U1051 (N_1051,N_692,N_117);
nor U1052 (N_1052,N_826,In_1876);
or U1053 (N_1053,N_613,N_200);
nor U1054 (N_1054,In_288,In_1075);
and U1055 (N_1055,N_592,N_753);
nand U1056 (N_1056,In_1409,N_988);
nand U1057 (N_1057,N_542,In_4);
and U1058 (N_1058,In_731,N_796);
nor U1059 (N_1059,N_778,In_404);
xnor U1060 (N_1060,N_719,N_243);
nand U1061 (N_1061,In_1984,In_1033);
nor U1062 (N_1062,N_317,N_479);
and U1063 (N_1063,N_686,N_874);
xnor U1064 (N_1064,In_433,N_944);
nor U1065 (N_1065,In_1103,In_659);
or U1066 (N_1066,N_842,In_1009);
nand U1067 (N_1067,N_961,N_627);
nand U1068 (N_1068,N_143,In_458);
nand U1069 (N_1069,N_353,N_463);
nor U1070 (N_1070,N_814,N_781);
and U1071 (N_1071,N_878,N_595);
xnor U1072 (N_1072,In_1044,N_241);
nand U1073 (N_1073,N_127,N_733);
nand U1074 (N_1074,In_699,N_968);
xnor U1075 (N_1075,In_1884,N_509);
nand U1076 (N_1076,N_860,N_973);
or U1077 (N_1077,N_270,N_759);
and U1078 (N_1078,N_941,In_188);
nor U1079 (N_1079,In_1052,N_872);
or U1080 (N_1080,In_1561,In_1555);
xnor U1081 (N_1081,In_553,In_1517);
nor U1082 (N_1082,N_687,N_803);
xor U1083 (N_1083,N_534,In_407);
and U1084 (N_1084,In_5,In_585);
or U1085 (N_1085,N_939,N_468);
and U1086 (N_1086,N_847,N_875);
xnor U1087 (N_1087,In_1193,In_892);
or U1088 (N_1088,N_980,In_1949);
xor U1089 (N_1089,N_641,N_239);
xor U1090 (N_1090,In_894,N_185);
xnor U1091 (N_1091,In_1607,N_620);
nor U1092 (N_1092,N_755,N_561);
and U1093 (N_1093,In_1654,In_324);
or U1094 (N_1094,N_914,N_885);
or U1095 (N_1095,In_635,In_247);
or U1096 (N_1096,N_989,In_1115);
or U1097 (N_1097,In_100,N_934);
xnor U1098 (N_1098,N_927,N_775);
nand U1099 (N_1099,N_723,In_346);
xnor U1100 (N_1100,In_1627,N_397);
and U1101 (N_1101,In_1129,In_1068);
xor U1102 (N_1102,In_197,N_806);
nor U1103 (N_1103,N_825,N_827);
or U1104 (N_1104,In_272,In_1985);
or U1105 (N_1105,N_372,N_456);
or U1106 (N_1106,N_29,In_1332);
or U1107 (N_1107,N_677,In_824);
and U1108 (N_1108,N_791,N_232);
nand U1109 (N_1109,In_730,N_963);
and U1110 (N_1110,N_691,In_198);
nor U1111 (N_1111,N_928,In_759);
nand U1112 (N_1112,N_154,In_1196);
nand U1113 (N_1113,N_833,N_771);
nand U1114 (N_1114,N_543,N_333);
or U1115 (N_1115,N_500,N_607);
or U1116 (N_1116,N_246,N_450);
or U1117 (N_1117,N_144,N_254);
nor U1118 (N_1118,N_722,In_1613);
and U1119 (N_1119,N_901,N_995);
nor U1120 (N_1120,In_898,In_1104);
or U1121 (N_1121,In_14,N_891);
or U1122 (N_1122,In_398,In_1840);
and U1123 (N_1123,In_1788,N_673);
and U1124 (N_1124,In_946,In_1462);
xor U1125 (N_1125,In_1547,N_336);
and U1126 (N_1126,N_129,N_679);
xor U1127 (N_1127,In_601,In_859);
and U1128 (N_1128,N_817,In_6);
nor U1129 (N_1129,N_929,N_931);
xnor U1130 (N_1130,In_135,In_768);
nor U1131 (N_1131,In_1920,N_782);
or U1132 (N_1132,N_644,N_108);
nor U1133 (N_1133,N_909,N_261);
nand U1134 (N_1134,N_683,In_234);
or U1135 (N_1135,N_892,In_178);
or U1136 (N_1136,N_919,In_570);
xnor U1137 (N_1137,N_160,In_310);
xnor U1138 (N_1138,N_767,N_957);
and U1139 (N_1139,N_258,N_808);
and U1140 (N_1140,N_643,N_514);
xnor U1141 (N_1141,N_87,In_637);
and U1142 (N_1142,N_887,N_635);
and U1143 (N_1143,In_1170,In_383);
nand U1144 (N_1144,In_1366,N_481);
xor U1145 (N_1145,In_1134,N_882);
nand U1146 (N_1146,N_908,In_563);
or U1147 (N_1147,N_583,N_444);
nand U1148 (N_1148,N_920,N_350);
nand U1149 (N_1149,N_924,N_587);
and U1150 (N_1150,In_945,In_979);
nor U1151 (N_1151,In_1853,In_1758);
nor U1152 (N_1152,In_1936,In_1034);
nand U1153 (N_1153,N_871,N_472);
nor U1154 (N_1154,N_831,N_492);
nand U1155 (N_1155,N_896,N_744);
nor U1156 (N_1156,N_881,In_79);
nand U1157 (N_1157,In_864,In_663);
and U1158 (N_1158,N_974,In_1002);
xor U1159 (N_1159,N_552,In_1977);
and U1160 (N_1160,N_816,N_625);
and U1161 (N_1161,N_569,N_649);
nand U1162 (N_1162,In_203,N_563);
nand U1163 (N_1163,N_204,N_520);
xnor U1164 (N_1164,N_773,N_912);
and U1165 (N_1165,In_22,N_611);
and U1166 (N_1166,N_203,In_180);
nand U1167 (N_1167,In_67,In_343);
nand U1168 (N_1168,In_134,N_709);
or U1169 (N_1169,N_227,In_1924);
nor U1170 (N_1170,N_925,In_1813);
nor U1171 (N_1171,In_1767,In_1982);
and U1172 (N_1172,N_830,In_236);
xnor U1173 (N_1173,In_338,N_838);
and U1174 (N_1174,In_1326,N_913);
xor U1175 (N_1175,N_418,N_0);
and U1176 (N_1176,In_154,N_538);
nor U1177 (N_1177,N_327,N_864);
nand U1178 (N_1178,N_150,N_960);
or U1179 (N_1179,In_1019,In_409);
xnor U1180 (N_1180,N_640,N_593);
xnor U1181 (N_1181,N_455,N_664);
and U1182 (N_1182,N_554,In_464);
xor U1183 (N_1183,N_470,In_602);
and U1184 (N_1184,N_932,In_1827);
nand U1185 (N_1185,N_862,N_906);
nand U1186 (N_1186,N_533,N_490);
nand U1187 (N_1187,N_942,In_1050);
nor U1188 (N_1188,N_666,N_818);
xor U1189 (N_1189,In_1041,N_889);
nand U1190 (N_1190,In_1941,N_442);
xnor U1191 (N_1191,N_718,N_763);
nor U1192 (N_1192,In_1739,In_1417);
nand U1193 (N_1193,In_1831,N_863);
xor U1194 (N_1194,N_280,N_626);
xnor U1195 (N_1195,In_528,N_813);
and U1196 (N_1196,In_617,N_519);
nand U1197 (N_1197,In_1578,N_930);
nor U1198 (N_1198,N_264,N_522);
nand U1199 (N_1199,In_1172,In_1304);
and U1200 (N_1200,In_697,N_202);
nor U1201 (N_1201,In_872,N_341);
or U1202 (N_1202,N_8,In_1874);
nand U1203 (N_1203,In_799,N_704);
xnor U1204 (N_1204,In_1908,N_153);
nand U1205 (N_1205,N_777,In_1852);
and U1206 (N_1206,N_905,N_849);
nand U1207 (N_1207,In_43,In_1164);
and U1208 (N_1208,In_1651,N_996);
xnor U1209 (N_1209,N_283,N_310);
xor U1210 (N_1210,N_943,N_976);
nand U1211 (N_1211,N_921,In_1817);
nand U1212 (N_1212,N_956,N_685);
nand U1213 (N_1213,N_760,N_698);
xnor U1214 (N_1214,N_32,In_1708);
or U1215 (N_1215,In_961,N_786);
and U1216 (N_1216,In_789,N_848);
or U1217 (N_1217,N_822,N_177);
or U1218 (N_1218,In_889,In_54);
xor U1219 (N_1219,In_1072,N_936);
or U1220 (N_1220,In_109,N_812);
and U1221 (N_1221,N_702,N_761);
or U1222 (N_1222,In_1943,In_1318);
nand U1223 (N_1223,In_1877,In_870);
nor U1224 (N_1224,N_74,N_706);
nand U1225 (N_1225,In_924,In_38);
and U1226 (N_1226,N_903,N_572);
and U1227 (N_1227,In_542,N_998);
xnor U1228 (N_1228,In_1751,In_681);
or U1229 (N_1229,In_1340,N_915);
or U1230 (N_1230,In_1641,In_1981);
and U1231 (N_1231,N_728,In_375);
or U1232 (N_1232,N_659,N_379);
nand U1233 (N_1233,In_1448,In_511);
and U1234 (N_1234,N_510,In_448);
nor U1235 (N_1235,In_1503,N_795);
xnor U1236 (N_1236,N_315,In_1120);
and U1237 (N_1237,In_1816,In_919);
and U1238 (N_1238,In_676,N_999);
nand U1239 (N_1239,N_801,In_1766);
and U1240 (N_1240,N_546,In_1606);
xnor U1241 (N_1241,N_926,N_532);
or U1242 (N_1242,In_1579,N_113);
or U1243 (N_1243,In_1325,N_983);
and U1244 (N_1244,N_437,N_170);
and U1245 (N_1245,In_1955,In_240);
xor U1246 (N_1246,N_528,N_553);
xnor U1247 (N_1247,N_334,N_923);
and U1248 (N_1248,N_708,In_179);
xor U1249 (N_1249,N_343,N_868);
and U1250 (N_1250,N_1192,In_657);
xnor U1251 (N_1251,N_1003,In_139);
nor U1252 (N_1252,N_119,N_904);
or U1253 (N_1253,N_947,In_545);
nand U1254 (N_1254,In_80,N_918);
or U1255 (N_1255,N_1099,N_774);
or U1256 (N_1256,N_884,In_1511);
and U1257 (N_1257,N_173,In_1904);
xor U1258 (N_1258,N_1004,In_1953);
nand U1259 (N_1259,N_541,In_1917);
xor U1260 (N_1260,In_620,N_1140);
nand U1261 (N_1261,N_1139,N_835);
and U1262 (N_1262,In_1420,N_1031);
and U1263 (N_1263,N_837,In_396);
or U1264 (N_1264,N_861,N_741);
nor U1265 (N_1265,N_1237,N_855);
and U1266 (N_1266,N_496,In_925);
nand U1267 (N_1267,In_173,In_1640);
or U1268 (N_1268,N_249,N_907);
nor U1269 (N_1269,N_1210,N_766);
nor U1270 (N_1270,In_462,N_1213);
and U1271 (N_1271,N_790,N_1134);
xnor U1272 (N_1272,N_1125,In_516);
and U1273 (N_1273,N_1204,N_501);
or U1274 (N_1274,N_606,N_311);
xnor U1275 (N_1275,In_1653,In_84);
and U1276 (N_1276,In_518,N_977);
and U1277 (N_1277,In_785,N_890);
xor U1278 (N_1278,N_1071,In_540);
nand U1279 (N_1279,N_959,N_1062);
xor U1280 (N_1280,N_535,N_1024);
or U1281 (N_1281,In_231,N_1047);
nand U1282 (N_1282,N_1053,N_1098);
xor U1283 (N_1283,In_446,N_982);
xor U1284 (N_1284,N_86,N_1015);
nand U1285 (N_1285,N_639,In_794);
nor U1286 (N_1286,N_1005,N_886);
nand U1287 (N_1287,In_151,In_1140);
xor U1288 (N_1288,N_1185,N_1067);
nand U1289 (N_1289,N_1208,N_476);
xor U1290 (N_1290,N_895,N_1249);
or U1291 (N_1291,In_1086,N_1211);
or U1292 (N_1292,N_917,N_756);
and U1293 (N_1293,N_1222,In_9);
xnor U1294 (N_1294,N_764,N_810);
nor U1295 (N_1295,In_1199,N_981);
xnor U1296 (N_1296,N_208,N_478);
or U1297 (N_1297,N_1243,N_751);
nor U1298 (N_1298,N_1058,N_1128);
nor U1299 (N_1299,N_1230,N_633);
nor U1300 (N_1300,N_1124,N_1034);
and U1301 (N_1301,N_780,N_1102);
xnor U1302 (N_1302,In_1238,In_1324);
and U1303 (N_1303,N_866,N_499);
nor U1304 (N_1304,In_1958,N_1158);
nor U1305 (N_1305,N_1127,N_388);
or U1306 (N_1306,N_577,N_693);
and U1307 (N_1307,In_569,N_787);
or U1308 (N_1308,N_798,N_1214);
and U1309 (N_1309,N_1085,N_1195);
nor U1310 (N_1310,In_305,In_1596);
xor U1311 (N_1311,N_1054,In_1937);
nor U1312 (N_1312,In_1362,In_1144);
or U1313 (N_1313,In_584,N_1059);
nand U1314 (N_1314,N_1025,N_181);
nand U1315 (N_1315,In_1893,In_582);
and U1316 (N_1316,N_840,N_176);
or U1317 (N_1317,N_409,In_1241);
and U1318 (N_1318,N_1007,N_382);
xor U1319 (N_1319,N_1151,In_1989);
xnor U1320 (N_1320,N_359,In_959);
and U1321 (N_1321,N_1044,N_1206);
and U1322 (N_1322,In_86,N_575);
and U1323 (N_1323,N_746,N_1164);
nor U1324 (N_1324,In_765,In_774);
or U1325 (N_1325,In_1156,N_344);
and U1326 (N_1326,N_1107,N_1184);
xor U1327 (N_1327,N_1154,N_617);
and U1328 (N_1328,N_1010,N_28);
nor U1329 (N_1329,N_602,N_110);
and U1330 (N_1330,N_1049,N_1233);
xor U1331 (N_1331,N_237,N_95);
nand U1332 (N_1332,In_1291,N_1104);
nand U1333 (N_1333,N_824,N_966);
nor U1334 (N_1334,In_460,N_1246);
nand U1335 (N_1335,In_316,N_916);
or U1336 (N_1336,N_858,N_1060);
and U1337 (N_1337,N_888,In_1988);
and U1338 (N_1338,N_839,N_1068);
nor U1339 (N_1339,N_1090,N_1247);
and U1340 (N_1340,N_820,In_1914);
nand U1341 (N_1341,N_428,In_1165);
nand U1342 (N_1342,N_675,N_159);
nand U1343 (N_1343,N_168,In_523);
or U1344 (N_1344,In_1994,In_931);
nor U1345 (N_1345,N_945,N_965);
xnor U1346 (N_1346,In_656,N_1144);
nand U1347 (N_1347,In_1236,N_984);
nor U1348 (N_1348,N_564,N_971);
xnor U1349 (N_1349,N_940,N_219);
or U1350 (N_1350,In_1211,N_1114);
or U1351 (N_1351,N_1150,N_1002);
xor U1352 (N_1352,N_47,In_1622);
xnor U1353 (N_1353,N_970,In_525);
and U1354 (N_1354,N_547,N_240);
xnor U1355 (N_1355,In_1728,N_1021);
nand U1356 (N_1356,In_1501,N_1033);
nand U1357 (N_1357,In_356,N_1178);
xnor U1358 (N_1358,In_1850,In_107);
xor U1359 (N_1359,N_962,N_681);
nand U1360 (N_1360,In_757,In_751);
nor U1361 (N_1361,In_499,N_35);
nand U1362 (N_1362,In_1812,N_900);
and U1363 (N_1363,N_1065,N_387);
nand U1364 (N_1364,In_834,N_1225);
nor U1365 (N_1365,In_1835,In_911);
nand U1366 (N_1366,In_213,In_285);
or U1367 (N_1367,N_139,N_616);
xor U1368 (N_1368,In_1397,N_991);
and U1369 (N_1369,N_1216,N_1095);
xnor U1370 (N_1370,In_37,N_894);
or U1371 (N_1371,N_1205,In_863);
nand U1372 (N_1372,N_1088,In_538);
nor U1373 (N_1373,In_402,N_211);
xnor U1374 (N_1374,N_1215,N_1212);
nor U1375 (N_1375,In_230,N_1038);
or U1376 (N_1376,N_823,N_1196);
nor U1377 (N_1377,In_1646,N_320);
nor U1378 (N_1378,N_754,N_1232);
nand U1379 (N_1379,N_1220,N_1012);
nand U1380 (N_1380,N_313,N_852);
nand U1381 (N_1381,N_1073,N_588);
and U1382 (N_1382,N_1110,N_805);
nor U1383 (N_1383,N_910,N_1087);
and U1384 (N_1384,N_762,In_1245);
or U1385 (N_1385,In_1492,N_1186);
and U1386 (N_1386,N_1175,N_678);
nand U1387 (N_1387,N_1086,N_1075);
or U1388 (N_1388,N_802,N_739);
nor U1389 (N_1389,In_651,In_807);
or U1390 (N_1390,N_354,In_140);
or U1391 (N_1391,N_1202,N_1041);
nand U1392 (N_1392,In_760,N_398);
nand U1393 (N_1393,N_1170,In_177);
xor U1394 (N_1394,N_1061,In_1472);
xnor U1395 (N_1395,N_636,N_1050);
xor U1396 (N_1396,In_289,In_1154);
nor U1397 (N_1397,In_1990,In_1150);
nor U1398 (N_1398,N_1245,In_259);
nor U1399 (N_1399,In_427,N_417);
nor U1400 (N_1400,N_1133,In_654);
or U1401 (N_1401,N_811,N_646);
nor U1402 (N_1402,N_1197,In_1389);
nand U1403 (N_1403,N_518,In_1524);
xor U1404 (N_1404,In_1232,In_412);
xnor U1405 (N_1405,N_312,N_1187);
nor U1406 (N_1406,N_157,N_1111);
xor U1407 (N_1407,N_380,In_1037);
or U1408 (N_1408,N_1117,N_1248);
nand U1409 (N_1409,N_506,In_70);
nor U1410 (N_1410,In_1979,N_421);
nand U1411 (N_1411,N_1069,N_1200);
and U1412 (N_1412,N_700,In_1969);
or U1413 (N_1413,In_1334,In_507);
and U1414 (N_1414,N_1239,N_416);
or U1415 (N_1415,N_669,N_600);
or U1416 (N_1416,N_1142,N_834);
or U1417 (N_1417,N_1063,N_793);
xor U1418 (N_1418,N_180,N_978);
nand U1419 (N_1419,N_804,N_1238);
nand U1420 (N_1420,N_274,N_1051);
nand U1421 (N_1421,N_140,N_715);
nand U1422 (N_1422,In_543,N_1076);
xor U1423 (N_1423,N_1019,N_1177);
xnor U1424 (N_1424,In_1184,N_870);
xor U1425 (N_1425,N_1166,N_1082);
xnor U1426 (N_1426,In_235,N_1236);
or U1427 (N_1427,In_658,N_1189);
nor U1428 (N_1428,N_1190,In_1716);
xnor U1429 (N_1429,N_671,N_815);
and U1430 (N_1430,N_1228,In_640);
nor U1431 (N_1431,N_1045,In_692);
nor U1432 (N_1432,N_1167,N_1103);
and U1433 (N_1433,N_972,N_809);
nor U1434 (N_1434,N_1056,In_1764);
or U1435 (N_1435,N_1101,N_992);
nand U1436 (N_1436,N_1244,N_190);
nor U1437 (N_1437,N_629,N_883);
xor U1438 (N_1438,N_1037,N_658);
nor U1439 (N_1439,In_386,In_598);
nor U1440 (N_1440,N_1057,N_618);
or U1441 (N_1441,N_1113,N_769);
nand U1442 (N_1442,In_833,N_1070);
nor U1443 (N_1443,N_628,In_1702);
and U1444 (N_1444,N_1152,N_1155);
nand U1445 (N_1445,N_271,N_670);
and U1446 (N_1446,N_857,N_390);
nor U1447 (N_1447,N_800,In_762);
nand U1448 (N_1448,N_1169,N_1163);
nand U1449 (N_1449,In_1809,In_1287);
nor U1450 (N_1450,N_1100,N_783);
nor U1451 (N_1451,N_770,N_1089);
xor U1452 (N_1452,N_1123,In_808);
or U1453 (N_1453,In_1021,N_295);
nor U1454 (N_1454,N_657,N_788);
nor U1455 (N_1455,N_34,N_272);
xor U1456 (N_1456,N_1149,N_1093);
xnor U1457 (N_1457,N_1027,N_1118);
and U1458 (N_1458,In_250,N_1129);
xnor U1459 (N_1459,In_815,In_1942);
nor U1460 (N_1460,N_727,N_469);
xnor U1461 (N_1461,N_1135,N_1028);
nand U1462 (N_1462,N_695,In_1458);
nand U1463 (N_1463,N_1201,N_307);
and U1464 (N_1464,N_1121,In_1160);
or U1465 (N_1465,In_1343,N_1116);
nand U1466 (N_1466,N_650,N_4);
and U1467 (N_1467,N_993,N_198);
or U1468 (N_1468,In_1476,N_582);
nor U1469 (N_1469,N_339,N_1168);
xnor U1470 (N_1470,N_1066,N_1043);
nor U1471 (N_1471,In_101,In_1053);
xnor U1472 (N_1472,In_69,N_711);
nor U1473 (N_1473,N_1091,N_318);
or U1474 (N_1474,N_609,N_162);
nor U1475 (N_1475,N_1209,N_1077);
nor U1476 (N_1476,N_1105,N_1112);
nor U1477 (N_1477,N_7,N_1126);
and U1478 (N_1478,N_612,In_1258);
xnor U1479 (N_1479,N_829,N_1193);
and U1480 (N_1480,N_893,N_937);
xor U1481 (N_1481,N_1055,In_1169);
or U1482 (N_1482,N_268,In_276);
nor U1483 (N_1483,N_853,N_621);
nand U1484 (N_1484,N_485,N_819);
nor U1485 (N_1485,N_1046,N_1180);
xnor U1486 (N_1486,In_763,N_1171);
xnor U1487 (N_1487,N_1188,In_92);
nand U1488 (N_1488,N_1020,In_1440);
xnor U1489 (N_1489,N_997,In_363);
nor U1490 (N_1490,N_1080,In_771);
nor U1491 (N_1491,N_933,N_985);
xor U1492 (N_1492,N_578,N_1153);
or U1493 (N_1493,In_1187,N_851);
or U1494 (N_1494,N_306,N_459);
nand U1495 (N_1495,N_1132,N_964);
xnor U1496 (N_1496,In_1889,N_1234);
xnor U1497 (N_1497,N_435,N_758);
and U1498 (N_1498,In_1443,N_1108);
nor U1499 (N_1499,N_1147,N_821);
or U1500 (N_1500,In_237,N_1064);
nand U1501 (N_1501,In_689,N_1405);
nor U1502 (N_1502,N_1263,N_1341);
xor U1503 (N_1503,N_1457,N_952);
and U1504 (N_1504,In_442,N_1137);
nor U1505 (N_1505,N_1282,In_614);
or U1506 (N_1506,N_776,In_174);
or U1507 (N_1507,In_790,N_1442);
nor U1508 (N_1508,N_1354,In_930);
or U1509 (N_1509,In_159,N_1323);
nand U1510 (N_1510,N_1487,N_1495);
nand U1511 (N_1511,In_1442,N_748);
xor U1512 (N_1512,In_1147,N_1298);
nor U1513 (N_1513,N_1026,N_1344);
xor U1514 (N_1514,In_968,N_1370);
and U1515 (N_1515,N_1436,N_1459);
xnor U1516 (N_1516,N_1444,N_1302);
and U1517 (N_1517,N_1250,N_486);
xnor U1518 (N_1518,N_1224,N_1468);
or U1519 (N_1519,In_376,N_732);
nor U1520 (N_1520,N_1431,N_898);
nor U1521 (N_1521,N_1252,N_1081);
or U1522 (N_1522,N_1030,N_1338);
xnor U1523 (N_1523,N_342,N_951);
and U1524 (N_1524,N_1219,N_1408);
nor U1525 (N_1525,In_927,N_1217);
and U1526 (N_1526,In_1923,N_1146);
or U1527 (N_1527,N_423,N_1411);
or U1528 (N_1528,N_1173,N_879);
nand U1529 (N_1529,N_1016,N_1381);
nand U1530 (N_1530,N_1242,N_1388);
nand U1531 (N_1531,In_533,N_471);
and U1532 (N_1532,N_1292,In_1151);
or U1533 (N_1533,N_1494,N_1039);
and U1534 (N_1534,N_1379,N_1227);
xor U1535 (N_1535,N_1413,N_1226);
nor U1536 (N_1536,N_772,In_1683);
xnor U1537 (N_1537,N_1321,N_1406);
and U1538 (N_1538,N_1359,N_841);
or U1539 (N_1539,N_877,In_1880);
xnor U1540 (N_1540,N_1083,N_1029);
xor U1541 (N_1541,N_1145,N_1465);
nor U1542 (N_1542,N_1429,N_1437);
and U1543 (N_1543,N_1262,N_276);
xor U1544 (N_1544,N_946,N_1013);
or U1545 (N_1545,N_1392,N_1430);
nand U1546 (N_1546,N_171,N_415);
and U1547 (N_1547,In_1502,N_513);
nand U1548 (N_1548,N_1376,N_1389);
nand U1549 (N_1549,N_740,N_1290);
nand U1550 (N_1550,N_1286,N_1276);
nand U1551 (N_1551,N_1275,N_1255);
xor U1552 (N_1552,N_1438,N_1412);
and U1553 (N_1553,N_1386,N_1448);
nor U1554 (N_1554,In_94,N_1447);
or U1555 (N_1555,N_725,N_1467);
nor U1556 (N_1556,N_680,N_1395);
xor U1557 (N_1557,N_253,N_1136);
nor U1558 (N_1558,N_1315,N_1254);
nor U1559 (N_1559,N_1475,N_1288);
nor U1560 (N_1560,In_1833,N_1426);
nand U1561 (N_1561,N_1308,N_836);
nand U1562 (N_1562,N_431,N_1156);
or U1563 (N_1563,N_1497,N_1331);
xor U1564 (N_1564,N_1048,In_482);
and U1565 (N_1565,In_1414,N_1294);
and U1566 (N_1566,N_792,N_1297);
nand U1567 (N_1567,In_332,N_1138);
xnor U1568 (N_1568,N_1489,N_1427);
and U1569 (N_1569,N_1466,N_1235);
nor U1570 (N_1570,In_1453,N_1040);
nand U1571 (N_1571,N_1306,N_1490);
nand U1572 (N_1572,N_1203,N_1143);
nor U1573 (N_1573,N_1273,N_76);
and U1574 (N_1574,N_1017,N_1074);
nor U1575 (N_1575,N_1218,N_1261);
or U1576 (N_1576,N_1317,N_1403);
xnor U1577 (N_1577,N_1314,N_1162);
and U1578 (N_1578,N_1410,N_1352);
and U1579 (N_1579,In_1177,N_565);
nor U1580 (N_1580,In_721,N_1305);
xnor U1581 (N_1581,N_807,N_603);
or U1582 (N_1582,N_1092,N_710);
xor U1583 (N_1583,In_1525,N_1499);
and U1584 (N_1584,N_1333,N_1482);
and U1585 (N_1585,N_1407,N_1373);
and U1586 (N_1586,N_1415,N_902);
and U1587 (N_1587,In_143,N_1366);
nor U1588 (N_1588,N_1384,N_1253);
and U1589 (N_1589,In_1399,N_922);
and U1590 (N_1590,In_185,N_1375);
nand U1591 (N_1591,N_1281,N_1347);
nor U1592 (N_1592,N_555,N_1471);
nor U1593 (N_1593,N_1148,In_430);
xnor U1594 (N_1594,N_674,N_1374);
or U1595 (N_1595,N_1367,In_1823);
nand U1596 (N_1596,N_1271,N_1364);
nand U1597 (N_1597,N_1318,N_1491);
nand U1598 (N_1598,N_1259,N_1371);
nand U1599 (N_1599,N_1327,N_1421);
nand U1600 (N_1600,N_1332,In_1744);
xnor U1601 (N_1601,N_1301,N_1141);
xnor U1602 (N_1602,N_1358,N_1032);
nand U1603 (N_1603,N_1404,N_53);
xor U1604 (N_1604,In_274,N_1397);
xor U1605 (N_1605,N_1369,N_1470);
and U1606 (N_1606,N_1401,In_645);
and U1607 (N_1607,N_1339,N_46);
nand U1608 (N_1608,N_1454,N_714);
or U1609 (N_1609,In_382,N_1312);
nor U1610 (N_1610,N_1336,N_410);
or U1611 (N_1611,N_1409,In_1939);
nor U1612 (N_1612,N_1283,N_548);
nand U1613 (N_1613,N_1334,N_955);
nand U1614 (N_1614,N_1455,N_705);
nor U1615 (N_1615,N_1439,N_1289);
nand U1616 (N_1616,N_1450,N_1097);
xor U1617 (N_1617,In_1100,In_707);
nor U1618 (N_1618,N_580,N_994);
nand U1619 (N_1619,N_1309,N_1131);
or U1620 (N_1620,N_953,N_1365);
nor U1621 (N_1621,N_1402,N_1313);
or U1622 (N_1622,N_248,N_1440);
or U1623 (N_1623,N_1052,N_1351);
xnor U1624 (N_1624,N_1417,N_1078);
nor U1625 (N_1625,N_1449,N_642);
and U1626 (N_1626,N_1009,N_1231);
nand U1627 (N_1627,In_121,N_752);
nand U1628 (N_1628,N_987,In_1345);
nand U1629 (N_1629,N_1320,N_1303);
and U1630 (N_1630,N_1194,N_1240);
xnor U1631 (N_1631,N_1355,N_1183);
nand U1632 (N_1632,N_1498,N_1399);
or U1633 (N_1633,N_1453,N_1496);
xnor U1634 (N_1634,In_192,N_1106);
and U1635 (N_1635,In_473,N_11);
xor U1636 (N_1636,In_956,N_1266);
or U1637 (N_1637,N_1435,N_873);
or U1638 (N_1638,N_1390,N_1361);
nor U1639 (N_1639,N_1461,In_938);
xor U1640 (N_1640,N_1036,N_406);
and U1641 (N_1641,N_785,N_797);
or U1642 (N_1642,N_1269,N_935);
or U1643 (N_1643,N_1277,N_1433);
nor U1644 (N_1644,N_1079,In_1743);
or U1645 (N_1645,N_845,N_1299);
xor U1646 (N_1646,N_1424,N_1042);
and U1647 (N_1647,In_680,N_1008);
xor U1648 (N_1648,N_1307,N_1265);
and U1649 (N_1649,N_1452,N_511);
and U1650 (N_1650,N_1441,N_1446);
or U1651 (N_1651,N_1159,N_1182);
xnor U1652 (N_1652,N_1418,N_1343);
nand U1653 (N_1653,In_93,N_1199);
and U1654 (N_1654,N_1472,N_1393);
and U1655 (N_1655,N_1368,N_1122);
nand U1656 (N_1656,N_1207,N_1325);
nor U1657 (N_1657,N_1300,N_523);
xnor U1658 (N_1658,N_1268,In_787);
or U1659 (N_1659,N_467,N_1014);
nor U1660 (N_1660,N_1251,In_1422);
or U1661 (N_1661,N_647,N_1161);
or U1662 (N_1662,N_1198,N_1394);
or U1663 (N_1663,N_1287,N_1348);
xnor U1664 (N_1664,N_1342,N_743);
or U1665 (N_1665,N_1414,N_1257);
and U1666 (N_1666,In_1089,N_512);
nor U1667 (N_1667,N_1425,N_408);
nand U1668 (N_1668,N_749,N_1432);
nand U1669 (N_1669,N_969,N_1130);
nand U1670 (N_1670,N_1492,N_1006);
and U1671 (N_1671,N_1383,N_1329);
and U1672 (N_1672,N_979,N_938);
or U1673 (N_1673,N_1120,N_1084);
nand U1674 (N_1674,N_1264,N_1241);
nor U1675 (N_1675,N_1396,N_1278);
nor U1676 (N_1676,N_1174,In_1776);
nand U1677 (N_1677,N_876,N_1462);
nand U1678 (N_1678,N_1221,N_1295);
xor U1679 (N_1679,N_1474,N_789);
nor U1680 (N_1680,N_1372,N_1291);
nor U1681 (N_1681,N_1000,N_530);
or U1682 (N_1682,N_1279,N_1023);
nor U1683 (N_1683,N_869,N_1445);
xor U1684 (N_1684,N_854,N_195);
nand U1685 (N_1685,In_1849,In_594);
or U1686 (N_1686,N_690,N_1420);
and U1687 (N_1687,N_1018,N_880);
and U1688 (N_1688,N_1094,N_1398);
xor U1689 (N_1689,N_1258,N_1362);
nand U1690 (N_1690,N_1304,N_1382);
or U1691 (N_1691,N_1416,N_1419);
xnor U1692 (N_1692,N_1363,In_1508);
nand U1693 (N_1693,N_1096,N_1479);
or U1694 (N_1694,N_1486,N_1328);
or U1695 (N_1695,N_1476,N_1280);
nand U1696 (N_1696,In_1905,N_1353);
and U1697 (N_1697,N_347,N_1346);
xor U1698 (N_1698,N_574,In_1048);
or U1699 (N_1699,N_1434,N_1345);
nand U1700 (N_1700,N_1310,N_1428);
and U1701 (N_1701,N_1349,In_522);
and U1702 (N_1702,N_30,N_726);
nand U1703 (N_1703,N_1483,N_1473);
nand U1704 (N_1704,N_1272,N_1378);
nor U1705 (N_1705,N_1001,In_691);
and U1706 (N_1706,N_1488,N_300);
nor U1707 (N_1707,N_1391,N_1322);
nand U1708 (N_1708,N_1458,N_1311);
xnor U1709 (N_1709,In_64,In_1700);
nor U1710 (N_1710,N_1022,N_1423);
or U1711 (N_1711,N_1456,N_1484);
and U1712 (N_1712,N_1072,N_1326);
or U1713 (N_1713,N_1493,N_1380);
nand U1714 (N_1714,N_1256,N_1478);
nand U1715 (N_1715,N_954,N_1469);
or U1716 (N_1716,N_843,N_1387);
nor U1717 (N_1717,N_1480,N_1335);
xor U1718 (N_1718,N_1229,N_1191);
xnor U1719 (N_1719,In_1013,N_365);
and U1720 (N_1720,N_1481,N_1285);
or U1721 (N_1721,N_1319,N_1316);
or U1722 (N_1722,N_1157,N_1451);
and U1723 (N_1723,N_1350,N_986);
and U1724 (N_1724,N_1340,In_118);
nor U1725 (N_1725,N_742,In_643);
and U1726 (N_1726,N_604,N_1400);
nand U1727 (N_1727,N_1119,N_859);
nand U1728 (N_1728,N_1115,N_1181);
nor U1729 (N_1729,N_1464,N_66);
nand U1730 (N_1730,N_1160,In_390);
or U1731 (N_1731,N_1223,N_1296);
nand U1732 (N_1732,N_1172,N_1293);
nor U1733 (N_1733,In_126,N_1011);
or U1734 (N_1734,N_1270,N_1260);
nor U1735 (N_1735,N_1274,N_1176);
nor U1736 (N_1736,N_1324,N_1356);
nor U1737 (N_1737,N_1377,N_1463);
or U1738 (N_1738,N_1422,N_1460);
nor U1739 (N_1739,In_49,N_1443);
or U1740 (N_1740,N_1485,N_1477);
xnor U1741 (N_1741,N_228,N_1284);
or U1742 (N_1742,N_1360,N_503);
nor U1743 (N_1743,N_1165,N_366);
xor U1744 (N_1744,N_49,N_1109);
xnor U1745 (N_1745,N_1385,N_1035);
nor U1746 (N_1746,N_1179,N_1357);
nand U1747 (N_1747,N_142,N_525);
xnor U1748 (N_1748,N_1337,N_1267);
or U1749 (N_1749,N_1330,N_768);
and U1750 (N_1750,N_1588,N_1545);
nor U1751 (N_1751,N_1745,N_1707);
nor U1752 (N_1752,N_1598,N_1694);
nand U1753 (N_1753,N_1739,N_1584);
nand U1754 (N_1754,N_1604,N_1563);
and U1755 (N_1755,N_1737,N_1668);
nand U1756 (N_1756,N_1705,N_1623);
xnor U1757 (N_1757,N_1519,N_1734);
or U1758 (N_1758,N_1695,N_1617);
nand U1759 (N_1759,N_1674,N_1503);
nor U1760 (N_1760,N_1552,N_1622);
or U1761 (N_1761,N_1501,N_1684);
and U1762 (N_1762,N_1644,N_1746);
and U1763 (N_1763,N_1649,N_1543);
xnor U1764 (N_1764,N_1675,N_1665);
nand U1765 (N_1765,N_1663,N_1693);
or U1766 (N_1766,N_1664,N_1625);
nor U1767 (N_1767,N_1553,N_1728);
xnor U1768 (N_1768,N_1560,N_1699);
and U1769 (N_1769,N_1690,N_1558);
nor U1770 (N_1770,N_1535,N_1578);
nor U1771 (N_1771,N_1506,N_1539);
or U1772 (N_1772,N_1743,N_1573);
and U1773 (N_1773,N_1517,N_1634);
xor U1774 (N_1774,N_1696,N_1609);
or U1775 (N_1775,N_1647,N_1606);
nor U1776 (N_1776,N_1616,N_1614);
nand U1777 (N_1777,N_1568,N_1706);
nor U1778 (N_1778,N_1725,N_1659);
nand U1779 (N_1779,N_1575,N_1631);
xnor U1780 (N_1780,N_1748,N_1718);
xor U1781 (N_1781,N_1580,N_1523);
nor U1782 (N_1782,N_1550,N_1505);
or U1783 (N_1783,N_1741,N_1642);
nand U1784 (N_1784,N_1708,N_1531);
and U1785 (N_1785,N_1522,N_1595);
or U1786 (N_1786,N_1747,N_1679);
and U1787 (N_1787,N_1726,N_1689);
and U1788 (N_1788,N_1507,N_1564);
and U1789 (N_1789,N_1658,N_1636);
or U1790 (N_1790,N_1525,N_1551);
or U1791 (N_1791,N_1597,N_1671);
and U1792 (N_1792,N_1736,N_1720);
and U1793 (N_1793,N_1530,N_1509);
xor U1794 (N_1794,N_1641,N_1585);
xor U1795 (N_1795,N_1610,N_1666);
and U1796 (N_1796,N_1715,N_1514);
nand U1797 (N_1797,N_1540,N_1735);
and U1798 (N_1798,N_1590,N_1562);
or U1799 (N_1799,N_1716,N_1630);
and U1800 (N_1800,N_1660,N_1600);
nand U1801 (N_1801,N_1723,N_1643);
nor U1802 (N_1802,N_1594,N_1678);
nand U1803 (N_1803,N_1592,N_1603);
xnor U1804 (N_1804,N_1656,N_1581);
nand U1805 (N_1805,N_1672,N_1730);
nand U1806 (N_1806,N_1516,N_1537);
and U1807 (N_1807,N_1719,N_1549);
xor U1808 (N_1808,N_1701,N_1653);
or U1809 (N_1809,N_1713,N_1591);
nor U1810 (N_1810,N_1686,N_1611);
and U1811 (N_1811,N_1621,N_1534);
nor U1812 (N_1812,N_1546,N_1577);
or U1813 (N_1813,N_1548,N_1740);
and U1814 (N_1814,N_1744,N_1638);
and U1815 (N_1815,N_1724,N_1650);
nor U1816 (N_1816,N_1742,N_1557);
nor U1817 (N_1817,N_1512,N_1566);
and U1818 (N_1818,N_1714,N_1619);
xor U1819 (N_1819,N_1618,N_1510);
or U1820 (N_1820,N_1710,N_1559);
nor U1821 (N_1821,N_1500,N_1700);
nand U1822 (N_1822,N_1587,N_1629);
or U1823 (N_1823,N_1536,N_1661);
xnor U1824 (N_1824,N_1593,N_1504);
nor U1825 (N_1825,N_1633,N_1555);
xor U1826 (N_1826,N_1627,N_1673);
or U1827 (N_1827,N_1607,N_1652);
or U1828 (N_1828,N_1583,N_1613);
nor U1829 (N_1829,N_1682,N_1569);
xnor U1830 (N_1830,N_1556,N_1691);
and U1831 (N_1831,N_1703,N_1579);
and U1832 (N_1832,N_1602,N_1651);
nor U1833 (N_1833,N_1632,N_1662);
xnor U1834 (N_1834,N_1729,N_1702);
nor U1835 (N_1835,N_1685,N_1738);
or U1836 (N_1836,N_1574,N_1692);
nor U1837 (N_1837,N_1677,N_1657);
nand U1838 (N_1838,N_1687,N_1608);
and U1839 (N_1839,N_1667,N_1518);
nor U1840 (N_1840,N_1711,N_1626);
nor U1841 (N_1841,N_1669,N_1646);
or U1842 (N_1842,N_1605,N_1565);
xor U1843 (N_1843,N_1533,N_1681);
or U1844 (N_1844,N_1547,N_1582);
and U1845 (N_1845,N_1640,N_1648);
nand U1846 (N_1846,N_1508,N_1628);
nor U1847 (N_1847,N_1521,N_1599);
xor U1848 (N_1848,N_1527,N_1567);
or U1849 (N_1849,N_1680,N_1697);
or U1850 (N_1850,N_1731,N_1727);
or U1851 (N_1851,N_1515,N_1502);
xnor U1852 (N_1852,N_1709,N_1698);
xor U1853 (N_1853,N_1645,N_1712);
and U1854 (N_1854,N_1529,N_1624);
or U1855 (N_1855,N_1637,N_1532);
nand U1856 (N_1856,N_1722,N_1670);
or U1857 (N_1857,N_1654,N_1511);
nand U1858 (N_1858,N_1576,N_1601);
nand U1859 (N_1859,N_1570,N_1717);
and U1860 (N_1860,N_1538,N_1571);
nor U1861 (N_1861,N_1596,N_1620);
nor U1862 (N_1862,N_1561,N_1554);
or U1863 (N_1863,N_1589,N_1524);
or U1864 (N_1864,N_1541,N_1572);
xnor U1865 (N_1865,N_1688,N_1676);
or U1866 (N_1866,N_1544,N_1612);
nand U1867 (N_1867,N_1721,N_1526);
or U1868 (N_1868,N_1615,N_1733);
nand U1869 (N_1869,N_1683,N_1639);
nor U1870 (N_1870,N_1542,N_1732);
nor U1871 (N_1871,N_1704,N_1513);
and U1872 (N_1872,N_1635,N_1528);
xor U1873 (N_1873,N_1520,N_1749);
and U1874 (N_1874,N_1655,N_1586);
and U1875 (N_1875,N_1714,N_1731);
nor U1876 (N_1876,N_1610,N_1639);
or U1877 (N_1877,N_1687,N_1708);
nor U1878 (N_1878,N_1658,N_1588);
or U1879 (N_1879,N_1742,N_1598);
or U1880 (N_1880,N_1744,N_1599);
nand U1881 (N_1881,N_1588,N_1645);
and U1882 (N_1882,N_1701,N_1610);
nor U1883 (N_1883,N_1626,N_1714);
xnor U1884 (N_1884,N_1556,N_1506);
nor U1885 (N_1885,N_1678,N_1584);
or U1886 (N_1886,N_1678,N_1506);
and U1887 (N_1887,N_1636,N_1560);
xor U1888 (N_1888,N_1536,N_1676);
and U1889 (N_1889,N_1730,N_1686);
xor U1890 (N_1890,N_1684,N_1547);
nand U1891 (N_1891,N_1644,N_1503);
or U1892 (N_1892,N_1642,N_1694);
nor U1893 (N_1893,N_1523,N_1561);
nor U1894 (N_1894,N_1525,N_1679);
xor U1895 (N_1895,N_1610,N_1650);
nor U1896 (N_1896,N_1519,N_1512);
nor U1897 (N_1897,N_1546,N_1557);
or U1898 (N_1898,N_1643,N_1599);
nand U1899 (N_1899,N_1638,N_1535);
xor U1900 (N_1900,N_1701,N_1659);
or U1901 (N_1901,N_1684,N_1714);
xor U1902 (N_1902,N_1705,N_1725);
and U1903 (N_1903,N_1639,N_1613);
xnor U1904 (N_1904,N_1565,N_1531);
nor U1905 (N_1905,N_1653,N_1535);
or U1906 (N_1906,N_1704,N_1531);
xnor U1907 (N_1907,N_1654,N_1723);
or U1908 (N_1908,N_1692,N_1550);
nor U1909 (N_1909,N_1601,N_1676);
and U1910 (N_1910,N_1691,N_1538);
nor U1911 (N_1911,N_1733,N_1536);
xnor U1912 (N_1912,N_1746,N_1583);
or U1913 (N_1913,N_1664,N_1694);
nand U1914 (N_1914,N_1561,N_1546);
xor U1915 (N_1915,N_1706,N_1585);
and U1916 (N_1916,N_1713,N_1562);
nor U1917 (N_1917,N_1625,N_1708);
and U1918 (N_1918,N_1728,N_1692);
xnor U1919 (N_1919,N_1543,N_1637);
nand U1920 (N_1920,N_1634,N_1514);
and U1921 (N_1921,N_1622,N_1688);
or U1922 (N_1922,N_1632,N_1626);
nor U1923 (N_1923,N_1731,N_1705);
or U1924 (N_1924,N_1503,N_1517);
and U1925 (N_1925,N_1561,N_1538);
nand U1926 (N_1926,N_1536,N_1541);
xnor U1927 (N_1927,N_1647,N_1605);
nand U1928 (N_1928,N_1689,N_1600);
or U1929 (N_1929,N_1548,N_1704);
or U1930 (N_1930,N_1663,N_1659);
xor U1931 (N_1931,N_1638,N_1704);
nand U1932 (N_1932,N_1515,N_1586);
and U1933 (N_1933,N_1708,N_1665);
xnor U1934 (N_1934,N_1518,N_1633);
xnor U1935 (N_1935,N_1722,N_1712);
or U1936 (N_1936,N_1557,N_1522);
or U1937 (N_1937,N_1639,N_1546);
and U1938 (N_1938,N_1636,N_1623);
nor U1939 (N_1939,N_1525,N_1523);
nor U1940 (N_1940,N_1709,N_1540);
nand U1941 (N_1941,N_1539,N_1573);
nand U1942 (N_1942,N_1634,N_1537);
nand U1943 (N_1943,N_1665,N_1558);
nand U1944 (N_1944,N_1500,N_1569);
nor U1945 (N_1945,N_1731,N_1553);
or U1946 (N_1946,N_1670,N_1505);
or U1947 (N_1947,N_1526,N_1728);
and U1948 (N_1948,N_1631,N_1692);
nand U1949 (N_1949,N_1620,N_1670);
xor U1950 (N_1950,N_1578,N_1597);
xor U1951 (N_1951,N_1540,N_1526);
and U1952 (N_1952,N_1533,N_1606);
nor U1953 (N_1953,N_1673,N_1507);
and U1954 (N_1954,N_1634,N_1687);
nor U1955 (N_1955,N_1640,N_1682);
xnor U1956 (N_1956,N_1537,N_1746);
and U1957 (N_1957,N_1519,N_1655);
nand U1958 (N_1958,N_1529,N_1630);
or U1959 (N_1959,N_1686,N_1618);
or U1960 (N_1960,N_1718,N_1671);
nor U1961 (N_1961,N_1729,N_1613);
nor U1962 (N_1962,N_1565,N_1582);
or U1963 (N_1963,N_1542,N_1703);
nand U1964 (N_1964,N_1570,N_1603);
nor U1965 (N_1965,N_1662,N_1690);
nand U1966 (N_1966,N_1517,N_1733);
and U1967 (N_1967,N_1670,N_1524);
and U1968 (N_1968,N_1549,N_1684);
xnor U1969 (N_1969,N_1583,N_1614);
nor U1970 (N_1970,N_1726,N_1642);
and U1971 (N_1971,N_1569,N_1712);
nand U1972 (N_1972,N_1553,N_1513);
nand U1973 (N_1973,N_1719,N_1746);
or U1974 (N_1974,N_1732,N_1591);
nor U1975 (N_1975,N_1514,N_1613);
nor U1976 (N_1976,N_1572,N_1688);
xor U1977 (N_1977,N_1565,N_1702);
nand U1978 (N_1978,N_1537,N_1563);
nand U1979 (N_1979,N_1742,N_1663);
xor U1980 (N_1980,N_1723,N_1661);
nand U1981 (N_1981,N_1515,N_1557);
nor U1982 (N_1982,N_1565,N_1594);
nand U1983 (N_1983,N_1641,N_1563);
nand U1984 (N_1984,N_1720,N_1731);
nand U1985 (N_1985,N_1663,N_1671);
nor U1986 (N_1986,N_1746,N_1533);
and U1987 (N_1987,N_1546,N_1646);
and U1988 (N_1988,N_1744,N_1511);
or U1989 (N_1989,N_1590,N_1702);
xnor U1990 (N_1990,N_1547,N_1530);
or U1991 (N_1991,N_1731,N_1686);
and U1992 (N_1992,N_1511,N_1526);
nor U1993 (N_1993,N_1551,N_1710);
nor U1994 (N_1994,N_1545,N_1625);
and U1995 (N_1995,N_1727,N_1598);
and U1996 (N_1996,N_1737,N_1639);
or U1997 (N_1997,N_1531,N_1620);
nor U1998 (N_1998,N_1504,N_1740);
nand U1999 (N_1999,N_1515,N_1638);
nand U2000 (N_2000,N_1980,N_1990);
nand U2001 (N_2001,N_1837,N_1935);
nand U2002 (N_2002,N_1945,N_1920);
nor U2003 (N_2003,N_1787,N_1893);
and U2004 (N_2004,N_1821,N_1951);
nor U2005 (N_2005,N_1810,N_1784);
or U2006 (N_2006,N_1939,N_1948);
xor U2007 (N_2007,N_1930,N_1831);
or U2008 (N_2008,N_1840,N_1823);
xor U2009 (N_2009,N_1923,N_1876);
nand U2010 (N_2010,N_1914,N_1752);
xnor U2011 (N_2011,N_1989,N_1828);
or U2012 (N_2012,N_1931,N_1934);
or U2013 (N_2013,N_1984,N_1834);
nand U2014 (N_2014,N_1909,N_1818);
xnor U2015 (N_2015,N_1897,N_1841);
xnor U2016 (N_2016,N_1906,N_1940);
nand U2017 (N_2017,N_1785,N_1757);
nor U2018 (N_2018,N_1864,N_1901);
nand U2019 (N_2019,N_1941,N_1777);
or U2020 (N_2020,N_1999,N_1965);
nand U2021 (N_2021,N_1826,N_1830);
and U2022 (N_2022,N_1822,N_1848);
nor U2023 (N_2023,N_1793,N_1960);
and U2024 (N_2024,N_1859,N_1884);
and U2025 (N_2025,N_1844,N_1987);
nand U2026 (N_2026,N_1946,N_1925);
nand U2027 (N_2027,N_1958,N_1872);
or U2028 (N_2028,N_1879,N_1938);
nor U2029 (N_2029,N_1781,N_1910);
or U2030 (N_2030,N_1776,N_1861);
and U2031 (N_2031,N_1800,N_1796);
and U2032 (N_2032,N_1877,N_1933);
and U2033 (N_2033,N_1887,N_1832);
nand U2034 (N_2034,N_1853,N_1790);
or U2035 (N_2035,N_1769,N_1838);
nor U2036 (N_2036,N_1806,N_1851);
nor U2037 (N_2037,N_1843,N_1847);
and U2038 (N_2038,N_1994,N_1928);
or U2039 (N_2039,N_1804,N_1882);
xor U2040 (N_2040,N_1802,N_1924);
xnor U2041 (N_2041,N_1981,N_1927);
or U2042 (N_2042,N_1978,N_1996);
or U2043 (N_2043,N_1943,N_1973);
and U2044 (N_2044,N_1795,N_1956);
or U2045 (N_2045,N_1904,N_1878);
xor U2046 (N_2046,N_1835,N_1805);
xor U2047 (N_2047,N_1783,N_1766);
nor U2048 (N_2048,N_1970,N_1916);
nand U2049 (N_2049,N_1883,N_1860);
or U2050 (N_2050,N_1949,N_1896);
or U2051 (N_2051,N_1880,N_1968);
nor U2052 (N_2052,N_1975,N_1858);
nand U2053 (N_2053,N_1891,N_1750);
or U2054 (N_2054,N_1812,N_1966);
xor U2055 (N_2055,N_1991,N_1993);
nor U2056 (N_2056,N_1971,N_1803);
nor U2057 (N_2057,N_1839,N_1873);
nor U2058 (N_2058,N_1936,N_1944);
xnor U2059 (N_2059,N_1801,N_1947);
nand U2060 (N_2060,N_1915,N_1833);
or U2061 (N_2061,N_1792,N_1767);
and U2062 (N_2062,N_1889,N_1842);
xnor U2063 (N_2063,N_1997,N_1798);
and U2064 (N_2064,N_1871,N_1808);
or U2065 (N_2065,N_1982,N_1825);
nand U2066 (N_2066,N_1778,N_1888);
and U2067 (N_2067,N_1772,N_1890);
nor U2068 (N_2068,N_1813,N_1942);
nor U2069 (N_2069,N_1881,N_1963);
xor U2070 (N_2070,N_1898,N_1952);
or U2071 (N_2071,N_1809,N_1751);
and U2072 (N_2072,N_1782,N_1850);
nor U2073 (N_2073,N_1870,N_1885);
xor U2074 (N_2074,N_1959,N_1950);
or U2075 (N_2075,N_1921,N_1900);
or U2076 (N_2076,N_1977,N_1829);
and U2077 (N_2077,N_1862,N_1845);
nor U2078 (N_2078,N_1854,N_1788);
or U2079 (N_2079,N_1976,N_1852);
and U2080 (N_2080,N_1824,N_1816);
xor U2081 (N_2081,N_1786,N_1998);
or U2082 (N_2082,N_1995,N_1986);
nand U2083 (N_2083,N_1929,N_1907);
nand U2084 (N_2084,N_1770,N_1985);
nor U2085 (N_2085,N_1819,N_1791);
or U2086 (N_2086,N_1857,N_1865);
and U2087 (N_2087,N_1836,N_1855);
and U2088 (N_2088,N_1773,N_1807);
nand U2089 (N_2089,N_1780,N_1955);
nor U2090 (N_2090,N_1756,N_1964);
or U2091 (N_2091,N_1972,N_1913);
nand U2092 (N_2092,N_1764,N_1820);
nor U2093 (N_2093,N_1875,N_1762);
nor U2094 (N_2094,N_1759,N_1911);
xnor U2095 (N_2095,N_1974,N_1918);
and U2096 (N_2096,N_1874,N_1919);
and U2097 (N_2097,N_1760,N_1753);
or U2098 (N_2098,N_1789,N_1917);
nand U2099 (N_2099,N_1869,N_1797);
xor U2100 (N_2100,N_1937,N_1758);
xnor U2101 (N_2101,N_1866,N_1932);
xnor U2102 (N_2102,N_1992,N_1892);
nor U2103 (N_2103,N_1794,N_1969);
xor U2104 (N_2104,N_1817,N_1761);
nand U2105 (N_2105,N_1908,N_1905);
nor U2106 (N_2106,N_1765,N_1988);
or U2107 (N_2107,N_1967,N_1926);
and U2108 (N_2108,N_1811,N_1867);
nand U2109 (N_2109,N_1895,N_1922);
nor U2110 (N_2110,N_1894,N_1983);
nor U2111 (N_2111,N_1763,N_1754);
xnor U2112 (N_2112,N_1954,N_1774);
nor U2113 (N_2113,N_1957,N_1856);
nand U2114 (N_2114,N_1755,N_1775);
nor U2115 (N_2115,N_1953,N_1779);
xor U2116 (N_2116,N_1799,N_1849);
nor U2117 (N_2117,N_1771,N_1768);
or U2118 (N_2118,N_1902,N_1979);
xnor U2119 (N_2119,N_1912,N_1899);
and U2120 (N_2120,N_1815,N_1886);
xnor U2121 (N_2121,N_1868,N_1962);
nand U2122 (N_2122,N_1814,N_1961);
or U2123 (N_2123,N_1846,N_1827);
nor U2124 (N_2124,N_1903,N_1863);
nand U2125 (N_2125,N_1804,N_1766);
nor U2126 (N_2126,N_1775,N_1798);
nand U2127 (N_2127,N_1877,N_1818);
nand U2128 (N_2128,N_1828,N_1859);
and U2129 (N_2129,N_1781,N_1922);
and U2130 (N_2130,N_1792,N_1794);
nor U2131 (N_2131,N_1805,N_1896);
nand U2132 (N_2132,N_1995,N_1921);
and U2133 (N_2133,N_1928,N_1975);
and U2134 (N_2134,N_1801,N_1779);
and U2135 (N_2135,N_1940,N_1981);
or U2136 (N_2136,N_1982,N_1818);
and U2137 (N_2137,N_1891,N_1910);
nor U2138 (N_2138,N_1898,N_1817);
nor U2139 (N_2139,N_1965,N_1766);
nor U2140 (N_2140,N_1980,N_1762);
nor U2141 (N_2141,N_1818,N_1898);
nor U2142 (N_2142,N_1843,N_1848);
xor U2143 (N_2143,N_1861,N_1820);
and U2144 (N_2144,N_1971,N_1838);
xnor U2145 (N_2145,N_1939,N_1996);
and U2146 (N_2146,N_1792,N_1865);
or U2147 (N_2147,N_1794,N_1966);
nand U2148 (N_2148,N_1782,N_1968);
or U2149 (N_2149,N_1757,N_1909);
xor U2150 (N_2150,N_1984,N_1843);
and U2151 (N_2151,N_1937,N_1901);
and U2152 (N_2152,N_1838,N_1786);
or U2153 (N_2153,N_1754,N_1838);
or U2154 (N_2154,N_1750,N_1795);
xor U2155 (N_2155,N_1950,N_1875);
or U2156 (N_2156,N_1991,N_1972);
nand U2157 (N_2157,N_1947,N_1998);
nor U2158 (N_2158,N_1841,N_1901);
and U2159 (N_2159,N_1810,N_1867);
nand U2160 (N_2160,N_1923,N_1990);
nor U2161 (N_2161,N_1926,N_1831);
nor U2162 (N_2162,N_1791,N_1938);
and U2163 (N_2163,N_1990,N_1941);
nand U2164 (N_2164,N_1814,N_1927);
and U2165 (N_2165,N_1851,N_1752);
or U2166 (N_2166,N_1813,N_1905);
nand U2167 (N_2167,N_1899,N_1791);
nor U2168 (N_2168,N_1798,N_1892);
nand U2169 (N_2169,N_1830,N_1849);
nand U2170 (N_2170,N_1791,N_1923);
and U2171 (N_2171,N_1872,N_1917);
or U2172 (N_2172,N_1806,N_1795);
xor U2173 (N_2173,N_1943,N_1926);
nand U2174 (N_2174,N_1817,N_1862);
nand U2175 (N_2175,N_1868,N_1988);
nand U2176 (N_2176,N_1893,N_1863);
xnor U2177 (N_2177,N_1779,N_1969);
nor U2178 (N_2178,N_1751,N_1783);
nor U2179 (N_2179,N_1975,N_1992);
xnor U2180 (N_2180,N_1865,N_1834);
or U2181 (N_2181,N_1953,N_1853);
nor U2182 (N_2182,N_1822,N_1926);
nand U2183 (N_2183,N_1840,N_1814);
xnor U2184 (N_2184,N_1859,N_1895);
xnor U2185 (N_2185,N_1835,N_1950);
and U2186 (N_2186,N_1944,N_1949);
xor U2187 (N_2187,N_1758,N_1987);
and U2188 (N_2188,N_1811,N_1896);
xor U2189 (N_2189,N_1761,N_1765);
xnor U2190 (N_2190,N_1822,N_1810);
nand U2191 (N_2191,N_1826,N_1861);
and U2192 (N_2192,N_1833,N_1923);
and U2193 (N_2193,N_1769,N_1857);
nor U2194 (N_2194,N_1833,N_1768);
xor U2195 (N_2195,N_1816,N_1843);
or U2196 (N_2196,N_1860,N_1829);
nor U2197 (N_2197,N_1774,N_1960);
nand U2198 (N_2198,N_1823,N_1986);
xnor U2199 (N_2199,N_1877,N_1858);
or U2200 (N_2200,N_1762,N_1977);
or U2201 (N_2201,N_1886,N_1767);
nand U2202 (N_2202,N_1793,N_1780);
xnor U2203 (N_2203,N_1901,N_1756);
or U2204 (N_2204,N_1863,N_1915);
xnor U2205 (N_2205,N_1990,N_1777);
xor U2206 (N_2206,N_1934,N_1866);
or U2207 (N_2207,N_1814,N_1934);
and U2208 (N_2208,N_1770,N_1794);
or U2209 (N_2209,N_1977,N_1795);
or U2210 (N_2210,N_1928,N_1757);
and U2211 (N_2211,N_1881,N_1789);
nor U2212 (N_2212,N_1803,N_1797);
and U2213 (N_2213,N_1889,N_1851);
or U2214 (N_2214,N_1852,N_1970);
or U2215 (N_2215,N_1898,N_1783);
and U2216 (N_2216,N_1871,N_1778);
nor U2217 (N_2217,N_1817,N_1927);
nand U2218 (N_2218,N_1998,N_1799);
nor U2219 (N_2219,N_1803,N_1857);
xor U2220 (N_2220,N_1963,N_1830);
nor U2221 (N_2221,N_1912,N_1987);
and U2222 (N_2222,N_1998,N_1845);
xor U2223 (N_2223,N_1800,N_1845);
or U2224 (N_2224,N_1953,N_1897);
xnor U2225 (N_2225,N_1798,N_1963);
nand U2226 (N_2226,N_1968,N_1862);
nand U2227 (N_2227,N_1938,N_1909);
nand U2228 (N_2228,N_1876,N_1791);
and U2229 (N_2229,N_1780,N_1771);
or U2230 (N_2230,N_1841,N_1755);
xor U2231 (N_2231,N_1945,N_1886);
nor U2232 (N_2232,N_1875,N_1781);
xnor U2233 (N_2233,N_1908,N_1991);
xnor U2234 (N_2234,N_1852,N_1908);
xnor U2235 (N_2235,N_1778,N_1782);
and U2236 (N_2236,N_1890,N_1847);
xnor U2237 (N_2237,N_1845,N_1969);
or U2238 (N_2238,N_1766,N_1827);
nand U2239 (N_2239,N_1859,N_1880);
nand U2240 (N_2240,N_1925,N_1989);
or U2241 (N_2241,N_1939,N_1883);
nand U2242 (N_2242,N_1810,N_1844);
or U2243 (N_2243,N_1986,N_1856);
or U2244 (N_2244,N_1919,N_1817);
or U2245 (N_2245,N_1934,N_1773);
xnor U2246 (N_2246,N_1799,N_1994);
and U2247 (N_2247,N_1830,N_1909);
nand U2248 (N_2248,N_1917,N_1869);
nand U2249 (N_2249,N_1938,N_1803);
and U2250 (N_2250,N_2072,N_2113);
and U2251 (N_2251,N_2187,N_2211);
or U2252 (N_2252,N_2112,N_2144);
nand U2253 (N_2253,N_2114,N_2058);
nand U2254 (N_2254,N_2078,N_2200);
and U2255 (N_2255,N_2123,N_2031);
or U2256 (N_2256,N_2015,N_2109);
and U2257 (N_2257,N_2244,N_2239);
nor U2258 (N_2258,N_2018,N_2236);
or U2259 (N_2259,N_2235,N_2183);
and U2260 (N_2260,N_2245,N_2080);
xor U2261 (N_2261,N_2110,N_2191);
nor U2262 (N_2262,N_2104,N_2141);
and U2263 (N_2263,N_2223,N_2051);
nand U2264 (N_2264,N_2026,N_2066);
nor U2265 (N_2265,N_2140,N_2180);
or U2266 (N_2266,N_2000,N_2093);
xor U2267 (N_2267,N_2130,N_2108);
and U2268 (N_2268,N_2238,N_2086);
and U2269 (N_2269,N_2192,N_2218);
nor U2270 (N_2270,N_2012,N_2036);
nand U2271 (N_2271,N_2160,N_2118);
nand U2272 (N_2272,N_2062,N_2069);
nand U2273 (N_2273,N_2045,N_2068);
or U2274 (N_2274,N_2161,N_2011);
nand U2275 (N_2275,N_2126,N_2122);
nor U2276 (N_2276,N_2025,N_2107);
or U2277 (N_2277,N_2179,N_2023);
nand U2278 (N_2278,N_2136,N_2052);
and U2279 (N_2279,N_2134,N_2013);
or U2280 (N_2280,N_2039,N_2171);
xnor U2281 (N_2281,N_2158,N_2081);
or U2282 (N_2282,N_2097,N_2247);
nand U2283 (N_2283,N_2102,N_2032);
xor U2284 (N_2284,N_2082,N_2129);
or U2285 (N_2285,N_2143,N_2040);
xor U2286 (N_2286,N_2079,N_2228);
nor U2287 (N_2287,N_2176,N_2221);
or U2288 (N_2288,N_2149,N_2248);
or U2289 (N_2289,N_2189,N_2207);
nor U2290 (N_2290,N_2215,N_2103);
or U2291 (N_2291,N_2226,N_2190);
nor U2292 (N_2292,N_2135,N_2150);
nand U2293 (N_2293,N_2001,N_2084);
nor U2294 (N_2294,N_2019,N_2137);
and U2295 (N_2295,N_2098,N_2153);
or U2296 (N_2296,N_2050,N_2243);
xnor U2297 (N_2297,N_2173,N_2185);
and U2298 (N_2298,N_2142,N_2182);
xor U2299 (N_2299,N_2155,N_2146);
and U2300 (N_2300,N_2085,N_2060);
nand U2301 (N_2301,N_2046,N_2196);
nor U2302 (N_2302,N_2044,N_2047);
nor U2303 (N_2303,N_2124,N_2101);
and U2304 (N_2304,N_2169,N_2120);
and U2305 (N_2305,N_2020,N_2198);
nor U2306 (N_2306,N_2028,N_2056);
nand U2307 (N_2307,N_2131,N_2194);
nand U2308 (N_2308,N_2111,N_2055);
or U2309 (N_2309,N_2145,N_2205);
xor U2310 (N_2310,N_2048,N_2174);
or U2311 (N_2311,N_2053,N_2240);
nand U2312 (N_2312,N_2208,N_2022);
or U2313 (N_2313,N_2237,N_2147);
or U2314 (N_2314,N_2202,N_2065);
nor U2315 (N_2315,N_2170,N_2159);
and U2316 (N_2316,N_2249,N_2116);
xnor U2317 (N_2317,N_2003,N_2059);
nor U2318 (N_2318,N_2178,N_2164);
nand U2319 (N_2319,N_2021,N_2231);
nand U2320 (N_2320,N_2076,N_2233);
and U2321 (N_2321,N_2214,N_2100);
and U2322 (N_2322,N_2206,N_2034);
nand U2323 (N_2323,N_2014,N_2027);
nand U2324 (N_2324,N_2168,N_2225);
and U2325 (N_2325,N_2105,N_2077);
nor U2326 (N_2326,N_2095,N_2106);
xnor U2327 (N_2327,N_2184,N_2212);
or U2328 (N_2328,N_2199,N_2125);
and U2329 (N_2329,N_2213,N_2156);
nor U2330 (N_2330,N_2121,N_2006);
and U2331 (N_2331,N_2075,N_2133);
and U2332 (N_2332,N_2004,N_2096);
and U2333 (N_2333,N_2167,N_2016);
nor U2334 (N_2334,N_2219,N_2089);
or U2335 (N_2335,N_2029,N_2151);
or U2336 (N_2336,N_2230,N_2242);
or U2337 (N_2337,N_2139,N_2210);
and U2338 (N_2338,N_2154,N_2073);
nor U2339 (N_2339,N_2119,N_2083);
nor U2340 (N_2340,N_2035,N_2224);
nand U2341 (N_2341,N_2157,N_2203);
xor U2342 (N_2342,N_2091,N_2177);
nand U2343 (N_2343,N_2024,N_2201);
nand U2344 (N_2344,N_2172,N_2094);
nor U2345 (N_2345,N_2054,N_2166);
or U2346 (N_2346,N_2043,N_2138);
nor U2347 (N_2347,N_2193,N_2049);
nand U2348 (N_2348,N_2186,N_2209);
nand U2349 (N_2349,N_2063,N_2002);
nor U2350 (N_2350,N_2216,N_2070);
nor U2351 (N_2351,N_2234,N_2127);
or U2352 (N_2352,N_2005,N_2181);
nor U2353 (N_2353,N_2099,N_2162);
or U2354 (N_2354,N_2064,N_2128);
nor U2355 (N_2355,N_2092,N_2175);
nor U2356 (N_2356,N_2009,N_2057);
xnor U2357 (N_2357,N_2115,N_2195);
or U2358 (N_2358,N_2061,N_2229);
nor U2359 (N_2359,N_2074,N_2041);
or U2360 (N_2360,N_2152,N_2090);
or U2361 (N_2361,N_2017,N_2030);
nand U2362 (N_2362,N_2132,N_2038);
or U2363 (N_2363,N_2067,N_2197);
nor U2364 (N_2364,N_2088,N_2165);
nor U2365 (N_2365,N_2246,N_2117);
nor U2366 (N_2366,N_2204,N_2010);
nor U2367 (N_2367,N_2232,N_2042);
and U2368 (N_2368,N_2222,N_2037);
nand U2369 (N_2369,N_2148,N_2033);
nand U2370 (N_2370,N_2188,N_2241);
or U2371 (N_2371,N_2217,N_2087);
and U2372 (N_2372,N_2008,N_2220);
nor U2373 (N_2373,N_2071,N_2163);
xnor U2374 (N_2374,N_2007,N_2227);
nand U2375 (N_2375,N_2093,N_2228);
or U2376 (N_2376,N_2159,N_2002);
nor U2377 (N_2377,N_2146,N_2136);
nand U2378 (N_2378,N_2013,N_2163);
and U2379 (N_2379,N_2207,N_2140);
or U2380 (N_2380,N_2238,N_2067);
nand U2381 (N_2381,N_2071,N_2016);
and U2382 (N_2382,N_2077,N_2159);
nand U2383 (N_2383,N_2205,N_2200);
nor U2384 (N_2384,N_2100,N_2006);
and U2385 (N_2385,N_2031,N_2205);
nor U2386 (N_2386,N_2182,N_2193);
nand U2387 (N_2387,N_2030,N_2181);
and U2388 (N_2388,N_2060,N_2225);
nand U2389 (N_2389,N_2041,N_2079);
nor U2390 (N_2390,N_2200,N_2068);
nor U2391 (N_2391,N_2065,N_2177);
and U2392 (N_2392,N_2107,N_2068);
xor U2393 (N_2393,N_2196,N_2049);
or U2394 (N_2394,N_2228,N_2009);
nand U2395 (N_2395,N_2071,N_2141);
nand U2396 (N_2396,N_2134,N_2021);
xor U2397 (N_2397,N_2110,N_2163);
or U2398 (N_2398,N_2060,N_2177);
nor U2399 (N_2399,N_2095,N_2104);
or U2400 (N_2400,N_2199,N_2196);
nor U2401 (N_2401,N_2042,N_2128);
xnor U2402 (N_2402,N_2141,N_2086);
xor U2403 (N_2403,N_2091,N_2102);
or U2404 (N_2404,N_2063,N_2113);
or U2405 (N_2405,N_2196,N_2142);
and U2406 (N_2406,N_2015,N_2196);
xnor U2407 (N_2407,N_2106,N_2236);
or U2408 (N_2408,N_2046,N_2049);
and U2409 (N_2409,N_2032,N_2183);
nand U2410 (N_2410,N_2141,N_2221);
and U2411 (N_2411,N_2239,N_2083);
xor U2412 (N_2412,N_2222,N_2080);
xnor U2413 (N_2413,N_2012,N_2086);
or U2414 (N_2414,N_2228,N_2158);
or U2415 (N_2415,N_2002,N_2160);
nor U2416 (N_2416,N_2245,N_2017);
nor U2417 (N_2417,N_2170,N_2198);
nand U2418 (N_2418,N_2126,N_2051);
nor U2419 (N_2419,N_2043,N_2115);
xor U2420 (N_2420,N_2064,N_2138);
nand U2421 (N_2421,N_2055,N_2227);
nand U2422 (N_2422,N_2054,N_2019);
nor U2423 (N_2423,N_2067,N_2236);
and U2424 (N_2424,N_2043,N_2226);
nor U2425 (N_2425,N_2005,N_2101);
nor U2426 (N_2426,N_2112,N_2217);
nand U2427 (N_2427,N_2227,N_2211);
nand U2428 (N_2428,N_2245,N_2244);
or U2429 (N_2429,N_2035,N_2181);
or U2430 (N_2430,N_2176,N_2244);
and U2431 (N_2431,N_2075,N_2046);
and U2432 (N_2432,N_2247,N_2143);
and U2433 (N_2433,N_2092,N_2143);
nor U2434 (N_2434,N_2139,N_2192);
or U2435 (N_2435,N_2249,N_2103);
and U2436 (N_2436,N_2076,N_2089);
nor U2437 (N_2437,N_2149,N_2193);
or U2438 (N_2438,N_2106,N_2052);
xnor U2439 (N_2439,N_2180,N_2012);
nand U2440 (N_2440,N_2082,N_2229);
nor U2441 (N_2441,N_2083,N_2069);
or U2442 (N_2442,N_2192,N_2163);
or U2443 (N_2443,N_2178,N_2135);
nor U2444 (N_2444,N_2203,N_2193);
nand U2445 (N_2445,N_2119,N_2106);
xnor U2446 (N_2446,N_2153,N_2034);
or U2447 (N_2447,N_2000,N_2102);
nand U2448 (N_2448,N_2193,N_2188);
xor U2449 (N_2449,N_2094,N_2081);
nand U2450 (N_2450,N_2106,N_2168);
and U2451 (N_2451,N_2237,N_2248);
nor U2452 (N_2452,N_2204,N_2086);
and U2453 (N_2453,N_2080,N_2158);
nor U2454 (N_2454,N_2007,N_2080);
or U2455 (N_2455,N_2248,N_2139);
or U2456 (N_2456,N_2156,N_2069);
nor U2457 (N_2457,N_2238,N_2188);
xnor U2458 (N_2458,N_2010,N_2006);
and U2459 (N_2459,N_2042,N_2040);
xnor U2460 (N_2460,N_2107,N_2026);
nand U2461 (N_2461,N_2195,N_2216);
or U2462 (N_2462,N_2193,N_2141);
nand U2463 (N_2463,N_2062,N_2040);
nand U2464 (N_2464,N_2225,N_2149);
or U2465 (N_2465,N_2108,N_2101);
nor U2466 (N_2466,N_2072,N_2184);
nand U2467 (N_2467,N_2197,N_2153);
nor U2468 (N_2468,N_2135,N_2239);
xnor U2469 (N_2469,N_2182,N_2223);
and U2470 (N_2470,N_2220,N_2178);
nor U2471 (N_2471,N_2040,N_2196);
or U2472 (N_2472,N_2106,N_2101);
nand U2473 (N_2473,N_2016,N_2039);
nand U2474 (N_2474,N_2067,N_2093);
and U2475 (N_2475,N_2247,N_2198);
nor U2476 (N_2476,N_2092,N_2068);
nor U2477 (N_2477,N_2238,N_2090);
and U2478 (N_2478,N_2205,N_2037);
nand U2479 (N_2479,N_2234,N_2197);
nor U2480 (N_2480,N_2165,N_2168);
and U2481 (N_2481,N_2125,N_2196);
and U2482 (N_2482,N_2056,N_2014);
xnor U2483 (N_2483,N_2118,N_2229);
nor U2484 (N_2484,N_2087,N_2133);
xor U2485 (N_2485,N_2053,N_2055);
nand U2486 (N_2486,N_2218,N_2025);
nor U2487 (N_2487,N_2094,N_2145);
xor U2488 (N_2488,N_2058,N_2122);
or U2489 (N_2489,N_2235,N_2229);
or U2490 (N_2490,N_2074,N_2114);
or U2491 (N_2491,N_2115,N_2098);
nand U2492 (N_2492,N_2126,N_2107);
or U2493 (N_2493,N_2181,N_2198);
xor U2494 (N_2494,N_2124,N_2118);
nand U2495 (N_2495,N_2093,N_2163);
or U2496 (N_2496,N_2041,N_2173);
xor U2497 (N_2497,N_2144,N_2132);
xnor U2498 (N_2498,N_2205,N_2156);
xor U2499 (N_2499,N_2029,N_2014);
nand U2500 (N_2500,N_2330,N_2472);
nor U2501 (N_2501,N_2413,N_2400);
and U2502 (N_2502,N_2433,N_2334);
or U2503 (N_2503,N_2403,N_2390);
and U2504 (N_2504,N_2349,N_2427);
and U2505 (N_2505,N_2291,N_2278);
or U2506 (N_2506,N_2262,N_2394);
nand U2507 (N_2507,N_2450,N_2387);
nand U2508 (N_2508,N_2339,N_2279);
xor U2509 (N_2509,N_2401,N_2492);
or U2510 (N_2510,N_2473,N_2280);
and U2511 (N_2511,N_2462,N_2360);
nand U2512 (N_2512,N_2455,N_2432);
nor U2513 (N_2513,N_2357,N_2377);
nor U2514 (N_2514,N_2251,N_2315);
nor U2515 (N_2515,N_2461,N_2420);
nor U2516 (N_2516,N_2428,N_2313);
nand U2517 (N_2517,N_2269,N_2454);
or U2518 (N_2518,N_2451,N_2437);
nand U2519 (N_2519,N_2407,N_2316);
nor U2520 (N_2520,N_2424,N_2258);
nand U2521 (N_2521,N_2396,N_2289);
nor U2522 (N_2522,N_2418,N_2345);
or U2523 (N_2523,N_2415,N_2267);
nand U2524 (N_2524,N_2331,N_2335);
or U2525 (N_2525,N_2302,N_2295);
and U2526 (N_2526,N_2355,N_2287);
nor U2527 (N_2527,N_2343,N_2449);
nor U2528 (N_2528,N_2388,N_2364);
or U2529 (N_2529,N_2479,N_2488);
or U2530 (N_2530,N_2442,N_2304);
xor U2531 (N_2531,N_2265,N_2435);
nor U2532 (N_2532,N_2333,N_2446);
and U2533 (N_2533,N_2310,N_2328);
or U2534 (N_2534,N_2372,N_2320);
or U2535 (N_2535,N_2478,N_2440);
xnor U2536 (N_2536,N_2294,N_2282);
nand U2537 (N_2537,N_2347,N_2392);
and U2538 (N_2538,N_2286,N_2417);
and U2539 (N_2539,N_2425,N_2452);
xnor U2540 (N_2540,N_2366,N_2476);
nor U2541 (N_2541,N_2419,N_2465);
or U2542 (N_2542,N_2380,N_2483);
or U2543 (N_2543,N_2374,N_2290);
xnor U2544 (N_2544,N_2429,N_2408);
or U2545 (N_2545,N_2378,N_2250);
nor U2546 (N_2546,N_2441,N_2395);
xnor U2547 (N_2547,N_2496,N_2327);
and U2548 (N_2548,N_2277,N_2490);
nor U2549 (N_2549,N_2404,N_2344);
and U2550 (N_2550,N_2480,N_2293);
nand U2551 (N_2551,N_2385,N_2272);
or U2552 (N_2552,N_2457,N_2351);
or U2553 (N_2553,N_2463,N_2296);
or U2554 (N_2554,N_2456,N_2324);
xor U2555 (N_2555,N_2284,N_2376);
nand U2556 (N_2556,N_2254,N_2382);
xnor U2557 (N_2557,N_2322,N_2271);
nor U2558 (N_2558,N_2439,N_2346);
and U2559 (N_2559,N_2270,N_2431);
xor U2560 (N_2560,N_2312,N_2308);
nor U2561 (N_2561,N_2484,N_2255);
or U2562 (N_2562,N_2356,N_2319);
nand U2563 (N_2563,N_2350,N_2253);
or U2564 (N_2564,N_2367,N_2363);
xnor U2565 (N_2565,N_2306,N_2336);
xor U2566 (N_2566,N_2263,N_2438);
nand U2567 (N_2567,N_2338,N_2281);
nand U2568 (N_2568,N_2353,N_2421);
nor U2569 (N_2569,N_2307,N_2303);
nand U2570 (N_2570,N_2311,N_2321);
nand U2571 (N_2571,N_2305,N_2361);
and U2572 (N_2572,N_2481,N_2423);
and U2573 (N_2573,N_2469,N_2383);
nor U2574 (N_2574,N_2292,N_2368);
or U2575 (N_2575,N_2399,N_2373);
xnor U2576 (N_2576,N_2371,N_2468);
xor U2577 (N_2577,N_2299,N_2348);
nand U2578 (N_2578,N_2358,N_2340);
nor U2579 (N_2579,N_2487,N_2416);
nor U2580 (N_2580,N_2430,N_2298);
nor U2581 (N_2581,N_2379,N_2436);
nor U2582 (N_2582,N_2393,N_2309);
or U2583 (N_2583,N_2409,N_2494);
nand U2584 (N_2584,N_2381,N_2273);
or U2585 (N_2585,N_2466,N_2285);
nand U2586 (N_2586,N_2475,N_2491);
or U2587 (N_2587,N_2410,N_2414);
nor U2588 (N_2588,N_2391,N_2362);
and U2589 (N_2589,N_2412,N_2314);
xnor U2590 (N_2590,N_2288,N_2489);
nor U2591 (N_2591,N_2365,N_2447);
or U2592 (N_2592,N_2317,N_2426);
and U2593 (N_2593,N_2467,N_2493);
xor U2594 (N_2594,N_2459,N_2359);
nor U2595 (N_2595,N_2337,N_2318);
or U2596 (N_2596,N_2325,N_2256);
and U2597 (N_2597,N_2464,N_2384);
nor U2598 (N_2598,N_2389,N_2386);
nor U2599 (N_2599,N_2444,N_2443);
nor U2600 (N_2600,N_2341,N_2261);
xnor U2601 (N_2601,N_2485,N_2252);
nor U2602 (N_2602,N_2445,N_2397);
and U2603 (N_2603,N_2274,N_2422);
and U2604 (N_2604,N_2474,N_2369);
nor U2605 (N_2605,N_2301,N_2411);
and U2606 (N_2606,N_2471,N_2497);
or U2607 (N_2607,N_2434,N_2352);
and U2608 (N_2608,N_2482,N_2375);
nor U2609 (N_2609,N_2264,N_2332);
or U2610 (N_2610,N_2266,N_2342);
and U2611 (N_2611,N_2297,N_2460);
nor U2612 (N_2612,N_2405,N_2275);
nand U2613 (N_2613,N_2370,N_2300);
or U2614 (N_2614,N_2495,N_2402);
or U2615 (N_2615,N_2486,N_2323);
or U2616 (N_2616,N_2276,N_2458);
and U2617 (N_2617,N_2477,N_2448);
xnor U2618 (N_2618,N_2326,N_2406);
xnor U2619 (N_2619,N_2257,N_2498);
nand U2620 (N_2620,N_2398,N_2453);
xor U2621 (N_2621,N_2354,N_2499);
and U2622 (N_2622,N_2283,N_2470);
xnor U2623 (N_2623,N_2259,N_2260);
nand U2624 (N_2624,N_2268,N_2329);
nor U2625 (N_2625,N_2309,N_2251);
xor U2626 (N_2626,N_2455,N_2420);
xor U2627 (N_2627,N_2432,N_2311);
xnor U2628 (N_2628,N_2475,N_2323);
xor U2629 (N_2629,N_2288,N_2266);
nand U2630 (N_2630,N_2387,N_2260);
or U2631 (N_2631,N_2275,N_2423);
or U2632 (N_2632,N_2280,N_2492);
nor U2633 (N_2633,N_2260,N_2453);
or U2634 (N_2634,N_2347,N_2308);
xor U2635 (N_2635,N_2474,N_2300);
or U2636 (N_2636,N_2289,N_2323);
or U2637 (N_2637,N_2452,N_2323);
or U2638 (N_2638,N_2291,N_2338);
nor U2639 (N_2639,N_2320,N_2387);
nor U2640 (N_2640,N_2367,N_2462);
nand U2641 (N_2641,N_2474,N_2269);
nand U2642 (N_2642,N_2493,N_2270);
xnor U2643 (N_2643,N_2400,N_2455);
nor U2644 (N_2644,N_2265,N_2273);
xor U2645 (N_2645,N_2302,N_2478);
nor U2646 (N_2646,N_2432,N_2274);
xnor U2647 (N_2647,N_2293,N_2302);
or U2648 (N_2648,N_2362,N_2498);
nand U2649 (N_2649,N_2319,N_2434);
nand U2650 (N_2650,N_2481,N_2388);
and U2651 (N_2651,N_2453,N_2320);
or U2652 (N_2652,N_2396,N_2349);
or U2653 (N_2653,N_2459,N_2416);
nor U2654 (N_2654,N_2489,N_2492);
xor U2655 (N_2655,N_2394,N_2275);
nand U2656 (N_2656,N_2495,N_2498);
and U2657 (N_2657,N_2431,N_2328);
nor U2658 (N_2658,N_2326,N_2380);
and U2659 (N_2659,N_2277,N_2458);
or U2660 (N_2660,N_2289,N_2338);
nor U2661 (N_2661,N_2385,N_2452);
and U2662 (N_2662,N_2385,N_2257);
or U2663 (N_2663,N_2272,N_2331);
nor U2664 (N_2664,N_2352,N_2386);
nor U2665 (N_2665,N_2452,N_2266);
xnor U2666 (N_2666,N_2439,N_2472);
nand U2667 (N_2667,N_2317,N_2439);
or U2668 (N_2668,N_2473,N_2452);
nor U2669 (N_2669,N_2310,N_2367);
nand U2670 (N_2670,N_2280,N_2406);
nor U2671 (N_2671,N_2457,N_2407);
or U2672 (N_2672,N_2306,N_2296);
or U2673 (N_2673,N_2402,N_2265);
or U2674 (N_2674,N_2313,N_2410);
nand U2675 (N_2675,N_2405,N_2378);
nand U2676 (N_2676,N_2422,N_2406);
or U2677 (N_2677,N_2323,N_2375);
nor U2678 (N_2678,N_2485,N_2323);
nand U2679 (N_2679,N_2348,N_2403);
and U2680 (N_2680,N_2291,N_2380);
nand U2681 (N_2681,N_2448,N_2499);
xor U2682 (N_2682,N_2421,N_2465);
or U2683 (N_2683,N_2341,N_2475);
nand U2684 (N_2684,N_2443,N_2260);
xor U2685 (N_2685,N_2309,N_2454);
nand U2686 (N_2686,N_2453,N_2362);
xnor U2687 (N_2687,N_2298,N_2316);
and U2688 (N_2688,N_2250,N_2497);
nor U2689 (N_2689,N_2429,N_2376);
and U2690 (N_2690,N_2319,N_2480);
and U2691 (N_2691,N_2482,N_2424);
or U2692 (N_2692,N_2309,N_2443);
and U2693 (N_2693,N_2453,N_2441);
xor U2694 (N_2694,N_2442,N_2386);
nor U2695 (N_2695,N_2492,N_2252);
or U2696 (N_2696,N_2375,N_2363);
xor U2697 (N_2697,N_2374,N_2364);
nand U2698 (N_2698,N_2459,N_2444);
or U2699 (N_2699,N_2275,N_2445);
xnor U2700 (N_2700,N_2292,N_2412);
xnor U2701 (N_2701,N_2264,N_2315);
and U2702 (N_2702,N_2471,N_2445);
nand U2703 (N_2703,N_2256,N_2479);
and U2704 (N_2704,N_2336,N_2450);
or U2705 (N_2705,N_2385,N_2307);
or U2706 (N_2706,N_2444,N_2397);
and U2707 (N_2707,N_2376,N_2324);
nor U2708 (N_2708,N_2348,N_2457);
and U2709 (N_2709,N_2446,N_2279);
xor U2710 (N_2710,N_2286,N_2496);
and U2711 (N_2711,N_2359,N_2312);
or U2712 (N_2712,N_2273,N_2484);
and U2713 (N_2713,N_2353,N_2322);
xor U2714 (N_2714,N_2487,N_2411);
and U2715 (N_2715,N_2256,N_2377);
and U2716 (N_2716,N_2468,N_2433);
nor U2717 (N_2717,N_2314,N_2486);
xnor U2718 (N_2718,N_2269,N_2310);
or U2719 (N_2719,N_2292,N_2350);
nor U2720 (N_2720,N_2428,N_2266);
nor U2721 (N_2721,N_2441,N_2278);
xnor U2722 (N_2722,N_2396,N_2254);
or U2723 (N_2723,N_2366,N_2297);
nor U2724 (N_2724,N_2306,N_2461);
or U2725 (N_2725,N_2471,N_2455);
and U2726 (N_2726,N_2296,N_2342);
nand U2727 (N_2727,N_2343,N_2365);
nor U2728 (N_2728,N_2370,N_2469);
nand U2729 (N_2729,N_2297,N_2353);
or U2730 (N_2730,N_2299,N_2393);
nor U2731 (N_2731,N_2499,N_2372);
and U2732 (N_2732,N_2260,N_2435);
or U2733 (N_2733,N_2417,N_2419);
or U2734 (N_2734,N_2273,N_2433);
xnor U2735 (N_2735,N_2356,N_2401);
nand U2736 (N_2736,N_2486,N_2319);
or U2737 (N_2737,N_2417,N_2482);
nor U2738 (N_2738,N_2335,N_2321);
nand U2739 (N_2739,N_2426,N_2306);
xnor U2740 (N_2740,N_2391,N_2319);
xor U2741 (N_2741,N_2435,N_2354);
nand U2742 (N_2742,N_2351,N_2269);
xor U2743 (N_2743,N_2399,N_2275);
nand U2744 (N_2744,N_2264,N_2380);
nor U2745 (N_2745,N_2356,N_2443);
xor U2746 (N_2746,N_2483,N_2481);
and U2747 (N_2747,N_2278,N_2415);
and U2748 (N_2748,N_2360,N_2265);
nor U2749 (N_2749,N_2476,N_2456);
or U2750 (N_2750,N_2740,N_2688);
and U2751 (N_2751,N_2746,N_2730);
and U2752 (N_2752,N_2630,N_2745);
and U2753 (N_2753,N_2723,N_2675);
and U2754 (N_2754,N_2742,N_2629);
or U2755 (N_2755,N_2601,N_2555);
and U2756 (N_2756,N_2574,N_2620);
or U2757 (N_2757,N_2591,N_2512);
and U2758 (N_2758,N_2611,N_2565);
or U2759 (N_2759,N_2505,N_2733);
xor U2760 (N_2760,N_2518,N_2508);
nor U2761 (N_2761,N_2524,N_2526);
nor U2762 (N_2762,N_2564,N_2588);
xnor U2763 (N_2763,N_2517,N_2682);
and U2764 (N_2764,N_2547,N_2576);
xor U2765 (N_2765,N_2624,N_2637);
xor U2766 (N_2766,N_2704,N_2737);
nor U2767 (N_2767,N_2627,N_2659);
and U2768 (N_2768,N_2600,N_2528);
nand U2769 (N_2769,N_2597,N_2502);
xor U2770 (N_2770,N_2748,N_2633);
nor U2771 (N_2771,N_2724,N_2676);
or U2772 (N_2772,N_2529,N_2587);
and U2773 (N_2773,N_2583,N_2510);
xor U2774 (N_2774,N_2527,N_2719);
xor U2775 (N_2775,N_2544,N_2613);
and U2776 (N_2776,N_2692,N_2551);
nor U2777 (N_2777,N_2718,N_2606);
and U2778 (N_2778,N_2603,N_2598);
or U2779 (N_2779,N_2680,N_2710);
or U2780 (N_2780,N_2739,N_2726);
nor U2781 (N_2781,N_2586,N_2647);
nor U2782 (N_2782,N_2521,N_2678);
and U2783 (N_2783,N_2605,N_2626);
xnor U2784 (N_2784,N_2595,N_2691);
and U2785 (N_2785,N_2687,N_2660);
nor U2786 (N_2786,N_2712,N_2674);
nand U2787 (N_2787,N_2522,N_2656);
nor U2788 (N_2788,N_2652,N_2609);
and U2789 (N_2789,N_2632,N_2649);
or U2790 (N_2790,N_2621,N_2658);
xor U2791 (N_2791,N_2725,N_2684);
or U2792 (N_2792,N_2590,N_2671);
nand U2793 (N_2793,N_2673,N_2594);
and U2794 (N_2794,N_2666,N_2523);
nor U2795 (N_2795,N_2728,N_2623);
or U2796 (N_2796,N_2501,N_2668);
nand U2797 (N_2797,N_2552,N_2511);
or U2798 (N_2798,N_2554,N_2634);
nand U2799 (N_2799,N_2667,N_2636);
nor U2800 (N_2800,N_2525,N_2734);
or U2801 (N_2801,N_2549,N_2604);
xor U2802 (N_2802,N_2639,N_2602);
or U2803 (N_2803,N_2542,N_2711);
and U2804 (N_2804,N_2701,N_2532);
xor U2805 (N_2805,N_2599,N_2727);
xor U2806 (N_2806,N_2720,N_2585);
nor U2807 (N_2807,N_2616,N_2628);
nor U2808 (N_2808,N_2622,N_2641);
and U2809 (N_2809,N_2507,N_2717);
or U2810 (N_2810,N_2556,N_2589);
nand U2811 (N_2811,N_2722,N_2643);
nand U2812 (N_2812,N_2703,N_2642);
nor U2813 (N_2813,N_2743,N_2625);
xor U2814 (N_2814,N_2580,N_2548);
xor U2815 (N_2815,N_2546,N_2545);
xnor U2816 (N_2816,N_2663,N_2566);
xor U2817 (N_2817,N_2608,N_2708);
xor U2818 (N_2818,N_2653,N_2563);
nand U2819 (N_2819,N_2694,N_2738);
and U2820 (N_2820,N_2533,N_2539);
xnor U2821 (N_2821,N_2593,N_2651);
or U2822 (N_2822,N_2749,N_2683);
nor U2823 (N_2823,N_2731,N_2655);
nand U2824 (N_2824,N_2575,N_2714);
nor U2825 (N_2825,N_2572,N_2614);
and U2826 (N_2826,N_2553,N_2541);
nor U2827 (N_2827,N_2699,N_2707);
nand U2828 (N_2828,N_2640,N_2540);
or U2829 (N_2829,N_2669,N_2509);
nand U2830 (N_2830,N_2741,N_2644);
nor U2831 (N_2831,N_2615,N_2581);
nand U2832 (N_2832,N_2662,N_2648);
and U2833 (N_2833,N_2559,N_2618);
xnor U2834 (N_2834,N_2698,N_2569);
nor U2835 (N_2835,N_2706,N_2700);
nand U2836 (N_2836,N_2535,N_2635);
or U2837 (N_2837,N_2513,N_2664);
and U2838 (N_2838,N_2685,N_2534);
nor U2839 (N_2839,N_2584,N_2530);
nand U2840 (N_2840,N_2577,N_2503);
and U2841 (N_2841,N_2672,N_2638);
nor U2842 (N_2842,N_2702,N_2619);
and U2843 (N_2843,N_2531,N_2665);
and U2844 (N_2844,N_2504,N_2557);
xor U2845 (N_2845,N_2661,N_2654);
or U2846 (N_2846,N_2650,N_2558);
or U2847 (N_2847,N_2744,N_2693);
xnor U2848 (N_2848,N_2568,N_2612);
nand U2849 (N_2849,N_2578,N_2582);
nand U2850 (N_2850,N_2721,N_2520);
xor U2851 (N_2851,N_2695,N_2696);
or U2852 (N_2852,N_2571,N_2506);
xnor U2853 (N_2853,N_2550,N_2536);
and U2854 (N_2854,N_2697,N_2689);
nor U2855 (N_2855,N_2579,N_2562);
nor U2856 (N_2856,N_2515,N_2514);
nand U2857 (N_2857,N_2716,N_2543);
xnor U2858 (N_2858,N_2500,N_2670);
xnor U2859 (N_2859,N_2610,N_2679);
or U2860 (N_2860,N_2537,N_2747);
or U2861 (N_2861,N_2690,N_2732);
or U2862 (N_2862,N_2645,N_2596);
nand U2863 (N_2863,N_2729,N_2631);
nand U2864 (N_2864,N_2715,N_2516);
xor U2865 (N_2865,N_2705,N_2686);
nor U2866 (N_2866,N_2538,N_2560);
and U2867 (N_2867,N_2573,N_2709);
xor U2868 (N_2868,N_2646,N_2570);
nand U2869 (N_2869,N_2677,N_2713);
and U2870 (N_2870,N_2607,N_2617);
xor U2871 (N_2871,N_2657,N_2592);
xnor U2872 (N_2872,N_2561,N_2519);
or U2873 (N_2873,N_2735,N_2736);
or U2874 (N_2874,N_2567,N_2681);
nand U2875 (N_2875,N_2701,N_2743);
nand U2876 (N_2876,N_2666,N_2638);
nand U2877 (N_2877,N_2623,N_2509);
xor U2878 (N_2878,N_2653,N_2685);
nand U2879 (N_2879,N_2546,N_2677);
nand U2880 (N_2880,N_2541,N_2643);
or U2881 (N_2881,N_2557,N_2704);
nand U2882 (N_2882,N_2632,N_2733);
nand U2883 (N_2883,N_2539,N_2574);
nand U2884 (N_2884,N_2727,N_2589);
or U2885 (N_2885,N_2748,N_2601);
xor U2886 (N_2886,N_2626,N_2677);
nor U2887 (N_2887,N_2615,N_2509);
nand U2888 (N_2888,N_2536,N_2590);
or U2889 (N_2889,N_2663,N_2522);
and U2890 (N_2890,N_2640,N_2624);
and U2891 (N_2891,N_2682,N_2588);
nand U2892 (N_2892,N_2612,N_2596);
nor U2893 (N_2893,N_2629,N_2565);
xnor U2894 (N_2894,N_2567,N_2682);
xor U2895 (N_2895,N_2536,N_2595);
or U2896 (N_2896,N_2520,N_2660);
nor U2897 (N_2897,N_2690,N_2611);
or U2898 (N_2898,N_2745,N_2722);
nand U2899 (N_2899,N_2628,N_2674);
or U2900 (N_2900,N_2743,N_2548);
nor U2901 (N_2901,N_2528,N_2523);
and U2902 (N_2902,N_2698,N_2593);
xor U2903 (N_2903,N_2739,N_2516);
nand U2904 (N_2904,N_2583,N_2527);
xor U2905 (N_2905,N_2555,N_2548);
nor U2906 (N_2906,N_2648,N_2564);
and U2907 (N_2907,N_2631,N_2566);
xnor U2908 (N_2908,N_2680,N_2667);
and U2909 (N_2909,N_2583,N_2544);
xor U2910 (N_2910,N_2723,N_2727);
xnor U2911 (N_2911,N_2654,N_2645);
xor U2912 (N_2912,N_2593,N_2655);
nor U2913 (N_2913,N_2705,N_2667);
nand U2914 (N_2914,N_2690,N_2555);
and U2915 (N_2915,N_2601,N_2572);
nand U2916 (N_2916,N_2683,N_2631);
and U2917 (N_2917,N_2528,N_2592);
nor U2918 (N_2918,N_2674,N_2688);
and U2919 (N_2919,N_2525,N_2624);
and U2920 (N_2920,N_2593,N_2680);
or U2921 (N_2921,N_2702,N_2627);
or U2922 (N_2922,N_2514,N_2564);
nor U2923 (N_2923,N_2724,N_2727);
and U2924 (N_2924,N_2507,N_2712);
and U2925 (N_2925,N_2522,N_2736);
or U2926 (N_2926,N_2571,N_2723);
nand U2927 (N_2927,N_2544,N_2512);
or U2928 (N_2928,N_2532,N_2534);
or U2929 (N_2929,N_2704,N_2609);
or U2930 (N_2930,N_2620,N_2526);
xnor U2931 (N_2931,N_2660,N_2581);
nand U2932 (N_2932,N_2634,N_2591);
xnor U2933 (N_2933,N_2694,N_2502);
nor U2934 (N_2934,N_2528,N_2580);
nand U2935 (N_2935,N_2540,N_2653);
nand U2936 (N_2936,N_2513,N_2503);
xnor U2937 (N_2937,N_2715,N_2587);
and U2938 (N_2938,N_2595,N_2569);
nor U2939 (N_2939,N_2632,N_2697);
nand U2940 (N_2940,N_2572,N_2637);
nand U2941 (N_2941,N_2628,N_2655);
nand U2942 (N_2942,N_2524,N_2606);
nand U2943 (N_2943,N_2619,N_2554);
nor U2944 (N_2944,N_2741,N_2703);
nor U2945 (N_2945,N_2576,N_2665);
and U2946 (N_2946,N_2631,N_2602);
nor U2947 (N_2947,N_2715,N_2691);
xnor U2948 (N_2948,N_2602,N_2555);
xnor U2949 (N_2949,N_2548,N_2602);
xnor U2950 (N_2950,N_2618,N_2629);
and U2951 (N_2951,N_2504,N_2626);
xnor U2952 (N_2952,N_2651,N_2553);
and U2953 (N_2953,N_2645,N_2629);
xor U2954 (N_2954,N_2734,N_2746);
nand U2955 (N_2955,N_2713,N_2616);
nor U2956 (N_2956,N_2508,N_2559);
xor U2957 (N_2957,N_2564,N_2666);
and U2958 (N_2958,N_2565,N_2583);
nor U2959 (N_2959,N_2722,N_2664);
or U2960 (N_2960,N_2578,N_2650);
and U2961 (N_2961,N_2582,N_2517);
and U2962 (N_2962,N_2633,N_2670);
nor U2963 (N_2963,N_2504,N_2558);
nor U2964 (N_2964,N_2572,N_2516);
xnor U2965 (N_2965,N_2705,N_2551);
and U2966 (N_2966,N_2686,N_2537);
nor U2967 (N_2967,N_2632,N_2702);
nor U2968 (N_2968,N_2701,N_2543);
xor U2969 (N_2969,N_2627,N_2680);
or U2970 (N_2970,N_2572,N_2699);
nand U2971 (N_2971,N_2585,N_2530);
nand U2972 (N_2972,N_2571,N_2533);
and U2973 (N_2973,N_2542,N_2604);
and U2974 (N_2974,N_2733,N_2529);
or U2975 (N_2975,N_2517,N_2569);
or U2976 (N_2976,N_2600,N_2504);
and U2977 (N_2977,N_2513,N_2658);
nand U2978 (N_2978,N_2504,N_2562);
nand U2979 (N_2979,N_2659,N_2708);
and U2980 (N_2980,N_2550,N_2574);
and U2981 (N_2981,N_2508,N_2723);
and U2982 (N_2982,N_2605,N_2708);
xor U2983 (N_2983,N_2673,N_2571);
nand U2984 (N_2984,N_2573,N_2670);
or U2985 (N_2985,N_2546,N_2638);
nor U2986 (N_2986,N_2649,N_2640);
or U2987 (N_2987,N_2504,N_2689);
nand U2988 (N_2988,N_2715,N_2537);
nand U2989 (N_2989,N_2552,N_2744);
and U2990 (N_2990,N_2738,N_2575);
and U2991 (N_2991,N_2570,N_2514);
xor U2992 (N_2992,N_2680,N_2517);
nor U2993 (N_2993,N_2521,N_2548);
nand U2994 (N_2994,N_2640,N_2742);
or U2995 (N_2995,N_2674,N_2597);
nor U2996 (N_2996,N_2596,N_2667);
xor U2997 (N_2997,N_2506,N_2624);
and U2998 (N_2998,N_2510,N_2632);
or U2999 (N_2999,N_2640,N_2564);
xnor U3000 (N_3000,N_2927,N_2821);
nor U3001 (N_3001,N_2878,N_2959);
or U3002 (N_3002,N_2920,N_2820);
or U3003 (N_3003,N_2816,N_2826);
nand U3004 (N_3004,N_2982,N_2795);
and U3005 (N_3005,N_2855,N_2757);
and U3006 (N_3006,N_2963,N_2922);
and U3007 (N_3007,N_2818,N_2781);
nand U3008 (N_3008,N_2997,N_2751);
xnor U3009 (N_3009,N_2805,N_2786);
and U3010 (N_3010,N_2951,N_2876);
nand U3011 (N_3011,N_2817,N_2775);
nor U3012 (N_3012,N_2886,N_2972);
nand U3013 (N_3013,N_2909,N_2849);
xnor U3014 (N_3014,N_2798,N_2938);
nor U3015 (N_3015,N_2806,N_2905);
nor U3016 (N_3016,N_2989,N_2772);
or U3017 (N_3017,N_2966,N_2801);
nor U3018 (N_3018,N_2888,N_2872);
xnor U3019 (N_3019,N_2840,N_2943);
xor U3020 (N_3020,N_2988,N_2904);
and U3021 (N_3021,N_2976,N_2809);
and U3022 (N_3022,N_2954,N_2933);
xor U3023 (N_3023,N_2811,N_2906);
or U3024 (N_3024,N_2918,N_2754);
nor U3025 (N_3025,N_2833,N_2823);
nor U3026 (N_3026,N_2994,N_2894);
nand U3027 (N_3027,N_2914,N_2908);
nor U3028 (N_3028,N_2926,N_2992);
xor U3029 (N_3029,N_2897,N_2893);
xor U3030 (N_3030,N_2907,N_2880);
nand U3031 (N_3031,N_2830,N_2971);
xor U3032 (N_3032,N_2841,N_2873);
nor U3033 (N_3033,N_2858,N_2766);
nand U3034 (N_3034,N_2862,N_2835);
xor U3035 (N_3035,N_2934,N_2783);
nor U3036 (N_3036,N_2881,N_2752);
or U3037 (N_3037,N_2928,N_2853);
nand U3038 (N_3038,N_2800,N_2923);
or U3039 (N_3039,N_2792,N_2990);
nand U3040 (N_3040,N_2902,N_2947);
nand U3041 (N_3041,N_2882,N_2856);
nand U3042 (N_3042,N_2812,N_2802);
xnor U3043 (N_3043,N_2970,N_2836);
or U3044 (N_3044,N_2919,N_2898);
and U3045 (N_3045,N_2998,N_2945);
and U3046 (N_3046,N_2771,N_2784);
nor U3047 (N_3047,N_2949,N_2819);
nand U3048 (N_3048,N_2760,N_2758);
xor U3049 (N_3049,N_2865,N_2985);
or U3050 (N_3050,N_2834,N_2861);
or U3051 (N_3051,N_2859,N_2790);
or U3052 (N_3052,N_2979,N_2965);
and U3053 (N_3053,N_2755,N_2848);
and U3054 (N_3054,N_2901,N_2750);
nor U3055 (N_3055,N_2968,N_2769);
nor U3056 (N_3056,N_2980,N_2846);
nand U3057 (N_3057,N_2774,N_2770);
or U3058 (N_3058,N_2753,N_2845);
or U3059 (N_3059,N_2764,N_2986);
nand U3060 (N_3060,N_2877,N_2955);
xor U3061 (N_3061,N_2891,N_2785);
nand U3062 (N_3062,N_2944,N_2956);
and U3063 (N_3063,N_2791,N_2779);
and U3064 (N_3064,N_2810,N_2782);
nor U3065 (N_3065,N_2883,N_2950);
xor U3066 (N_3066,N_2776,N_2958);
nand U3067 (N_3067,N_2870,N_2890);
xor U3068 (N_3068,N_2804,N_2767);
nand U3069 (N_3069,N_2860,N_2799);
or U3070 (N_3070,N_2829,N_2838);
nor U3071 (N_3071,N_2843,N_2763);
nor U3072 (N_3072,N_2924,N_2788);
nand U3073 (N_3073,N_2967,N_2863);
and U3074 (N_3074,N_2825,N_2837);
nor U3075 (N_3075,N_2868,N_2983);
and U3076 (N_3076,N_2822,N_2857);
nor U3077 (N_3077,N_2814,N_2889);
xnor U3078 (N_3078,N_2869,N_2773);
nand U3079 (N_3079,N_2975,N_2887);
nand U3080 (N_3080,N_2797,N_2991);
xnor U3081 (N_3081,N_2867,N_2948);
and U3082 (N_3082,N_2981,N_2900);
or U3083 (N_3083,N_2916,N_2871);
and U3084 (N_3084,N_2895,N_2842);
or U3085 (N_3085,N_2987,N_2864);
and U3086 (N_3086,N_2915,N_2999);
and U3087 (N_3087,N_2939,N_2852);
and U3088 (N_3088,N_2952,N_2778);
or U3089 (N_3089,N_2780,N_2953);
or U3090 (N_3090,N_2931,N_2828);
or U3091 (N_3091,N_2962,N_2996);
or U3092 (N_3092,N_2932,N_2941);
nand U3093 (N_3093,N_2929,N_2960);
nor U3094 (N_3094,N_2977,N_2844);
xor U3095 (N_3095,N_2875,N_2892);
and U3096 (N_3096,N_2815,N_2854);
xnor U3097 (N_3097,N_2974,N_2765);
and U3098 (N_3098,N_2759,N_2850);
and U3099 (N_3099,N_2995,N_2935);
and U3100 (N_3100,N_2813,N_2984);
nand U3101 (N_3101,N_2787,N_2957);
or U3102 (N_3102,N_2946,N_2827);
xor U3103 (N_3103,N_2993,N_2969);
or U3104 (N_3104,N_2807,N_2936);
and U3105 (N_3105,N_2910,N_2913);
or U3106 (N_3106,N_2911,N_2793);
and U3107 (N_3107,N_2899,N_2803);
or U3108 (N_3108,N_2832,N_2794);
or U3109 (N_3109,N_2937,N_2973);
and U3110 (N_3110,N_2874,N_2768);
nand U3111 (N_3111,N_2851,N_2879);
xnor U3112 (N_3112,N_2762,N_2866);
nor U3113 (N_3113,N_2831,N_2761);
and U3114 (N_3114,N_2917,N_2885);
nand U3115 (N_3115,N_2942,N_2789);
or U3116 (N_3116,N_2912,N_2796);
and U3117 (N_3117,N_2756,N_2940);
and U3118 (N_3118,N_2978,N_2839);
nand U3119 (N_3119,N_2896,N_2961);
and U3120 (N_3120,N_2777,N_2847);
nor U3121 (N_3121,N_2921,N_2824);
or U3122 (N_3122,N_2884,N_2930);
or U3123 (N_3123,N_2925,N_2964);
nand U3124 (N_3124,N_2808,N_2903);
nand U3125 (N_3125,N_2884,N_2944);
nor U3126 (N_3126,N_2838,N_2814);
nor U3127 (N_3127,N_2857,N_2814);
and U3128 (N_3128,N_2771,N_2897);
xor U3129 (N_3129,N_2875,N_2978);
xor U3130 (N_3130,N_2967,N_2861);
and U3131 (N_3131,N_2802,N_2818);
nand U3132 (N_3132,N_2903,N_2997);
nand U3133 (N_3133,N_2750,N_2885);
and U3134 (N_3134,N_2872,N_2848);
xor U3135 (N_3135,N_2835,N_2916);
xor U3136 (N_3136,N_2792,N_2874);
nand U3137 (N_3137,N_2799,N_2821);
xor U3138 (N_3138,N_2762,N_2882);
or U3139 (N_3139,N_2859,N_2757);
and U3140 (N_3140,N_2828,N_2934);
nand U3141 (N_3141,N_2956,N_2821);
and U3142 (N_3142,N_2892,N_2964);
and U3143 (N_3143,N_2907,N_2764);
or U3144 (N_3144,N_2825,N_2937);
nor U3145 (N_3145,N_2786,N_2961);
nand U3146 (N_3146,N_2879,N_2957);
nor U3147 (N_3147,N_2951,N_2843);
nand U3148 (N_3148,N_2783,N_2948);
xor U3149 (N_3149,N_2934,N_2887);
nand U3150 (N_3150,N_2909,N_2895);
nor U3151 (N_3151,N_2860,N_2918);
and U3152 (N_3152,N_2937,N_2965);
or U3153 (N_3153,N_2867,N_2802);
nor U3154 (N_3154,N_2965,N_2885);
or U3155 (N_3155,N_2867,N_2836);
nand U3156 (N_3156,N_2857,N_2839);
and U3157 (N_3157,N_2918,N_2804);
xor U3158 (N_3158,N_2926,N_2795);
xor U3159 (N_3159,N_2852,N_2987);
xor U3160 (N_3160,N_2804,N_2835);
nor U3161 (N_3161,N_2797,N_2798);
nor U3162 (N_3162,N_2903,N_2990);
nor U3163 (N_3163,N_2805,N_2956);
nand U3164 (N_3164,N_2956,N_2830);
or U3165 (N_3165,N_2960,N_2796);
nand U3166 (N_3166,N_2919,N_2980);
and U3167 (N_3167,N_2905,N_2920);
xnor U3168 (N_3168,N_2800,N_2852);
nor U3169 (N_3169,N_2830,N_2898);
or U3170 (N_3170,N_2962,N_2862);
and U3171 (N_3171,N_2962,N_2865);
and U3172 (N_3172,N_2859,N_2983);
and U3173 (N_3173,N_2776,N_2953);
and U3174 (N_3174,N_2929,N_2824);
nand U3175 (N_3175,N_2753,N_2798);
nand U3176 (N_3176,N_2756,N_2920);
xor U3177 (N_3177,N_2826,N_2812);
or U3178 (N_3178,N_2796,N_2821);
xor U3179 (N_3179,N_2910,N_2873);
and U3180 (N_3180,N_2960,N_2984);
nor U3181 (N_3181,N_2944,N_2964);
nor U3182 (N_3182,N_2893,N_2784);
and U3183 (N_3183,N_2879,N_2870);
or U3184 (N_3184,N_2873,N_2760);
xor U3185 (N_3185,N_2757,N_2785);
and U3186 (N_3186,N_2767,N_2966);
nor U3187 (N_3187,N_2892,N_2942);
xor U3188 (N_3188,N_2986,N_2979);
xor U3189 (N_3189,N_2991,N_2860);
xor U3190 (N_3190,N_2983,N_2957);
nor U3191 (N_3191,N_2762,N_2954);
nor U3192 (N_3192,N_2948,N_2990);
xor U3193 (N_3193,N_2991,N_2965);
nand U3194 (N_3194,N_2835,N_2788);
and U3195 (N_3195,N_2787,N_2757);
or U3196 (N_3196,N_2818,N_2864);
or U3197 (N_3197,N_2939,N_2980);
or U3198 (N_3198,N_2764,N_2762);
xor U3199 (N_3199,N_2862,N_2905);
and U3200 (N_3200,N_2960,N_2765);
and U3201 (N_3201,N_2763,N_2781);
nor U3202 (N_3202,N_2944,N_2762);
xnor U3203 (N_3203,N_2771,N_2887);
nor U3204 (N_3204,N_2873,N_2918);
and U3205 (N_3205,N_2908,N_2962);
nor U3206 (N_3206,N_2976,N_2797);
xor U3207 (N_3207,N_2870,N_2974);
or U3208 (N_3208,N_2828,N_2825);
nand U3209 (N_3209,N_2801,N_2844);
xor U3210 (N_3210,N_2885,N_2944);
and U3211 (N_3211,N_2764,N_2824);
and U3212 (N_3212,N_2855,N_2890);
and U3213 (N_3213,N_2891,N_2855);
or U3214 (N_3214,N_2808,N_2960);
xnor U3215 (N_3215,N_2895,N_2808);
and U3216 (N_3216,N_2785,N_2934);
xnor U3217 (N_3217,N_2796,N_2901);
nor U3218 (N_3218,N_2872,N_2785);
nor U3219 (N_3219,N_2758,N_2886);
xnor U3220 (N_3220,N_2926,N_2816);
and U3221 (N_3221,N_2996,N_2966);
nor U3222 (N_3222,N_2913,N_2836);
nand U3223 (N_3223,N_2947,N_2869);
nor U3224 (N_3224,N_2953,N_2889);
nand U3225 (N_3225,N_2840,N_2787);
xnor U3226 (N_3226,N_2959,N_2898);
and U3227 (N_3227,N_2910,N_2823);
and U3228 (N_3228,N_2995,N_2780);
xor U3229 (N_3229,N_2966,N_2938);
nand U3230 (N_3230,N_2930,N_2916);
and U3231 (N_3231,N_2751,N_2855);
nor U3232 (N_3232,N_2975,N_2953);
xor U3233 (N_3233,N_2867,N_2940);
xnor U3234 (N_3234,N_2872,N_2890);
or U3235 (N_3235,N_2971,N_2770);
nor U3236 (N_3236,N_2957,N_2883);
and U3237 (N_3237,N_2872,N_2924);
xnor U3238 (N_3238,N_2890,N_2918);
nand U3239 (N_3239,N_2960,N_2881);
or U3240 (N_3240,N_2792,N_2982);
and U3241 (N_3241,N_2826,N_2785);
and U3242 (N_3242,N_2869,N_2780);
nor U3243 (N_3243,N_2826,N_2833);
and U3244 (N_3244,N_2806,N_2790);
nor U3245 (N_3245,N_2923,N_2954);
and U3246 (N_3246,N_2907,N_2962);
nor U3247 (N_3247,N_2986,N_2772);
nor U3248 (N_3248,N_2829,N_2912);
and U3249 (N_3249,N_2807,N_2783);
xor U3250 (N_3250,N_3191,N_3061);
and U3251 (N_3251,N_3068,N_3145);
nand U3252 (N_3252,N_3077,N_3097);
nand U3253 (N_3253,N_3238,N_3092);
nor U3254 (N_3254,N_3067,N_3165);
nand U3255 (N_3255,N_3190,N_3080);
nand U3256 (N_3256,N_3195,N_3128);
xnor U3257 (N_3257,N_3249,N_3139);
or U3258 (N_3258,N_3159,N_3149);
xor U3259 (N_3259,N_3166,N_3236);
and U3260 (N_3260,N_3079,N_3181);
nor U3261 (N_3261,N_3132,N_3086);
xor U3262 (N_3262,N_3216,N_3221);
nor U3263 (N_3263,N_3019,N_3242);
nor U3264 (N_3264,N_3057,N_3107);
xnor U3265 (N_3265,N_3028,N_3151);
and U3266 (N_3266,N_3228,N_3150);
nand U3267 (N_3267,N_3235,N_3192);
xnor U3268 (N_3268,N_3202,N_3185);
or U3269 (N_3269,N_3072,N_3026);
or U3270 (N_3270,N_3143,N_3188);
and U3271 (N_3271,N_3046,N_3146);
nor U3272 (N_3272,N_3002,N_3135);
or U3273 (N_3273,N_3214,N_3137);
nand U3274 (N_3274,N_3204,N_3099);
nor U3275 (N_3275,N_3194,N_3048);
xor U3276 (N_3276,N_3127,N_3016);
and U3277 (N_3277,N_3123,N_3144);
and U3278 (N_3278,N_3167,N_3164);
and U3279 (N_3279,N_3121,N_3248);
nor U3280 (N_3280,N_3170,N_3119);
nor U3281 (N_3281,N_3113,N_3125);
or U3282 (N_3282,N_3233,N_3075);
nor U3283 (N_3283,N_3005,N_3102);
nor U3284 (N_3284,N_3162,N_3037);
nor U3285 (N_3285,N_3074,N_3219);
nand U3286 (N_3286,N_3062,N_3239);
or U3287 (N_3287,N_3206,N_3241);
nor U3288 (N_3288,N_3025,N_3215);
nor U3289 (N_3289,N_3234,N_3232);
nor U3290 (N_3290,N_3040,N_3160);
or U3291 (N_3291,N_3171,N_3010);
xor U3292 (N_3292,N_3060,N_3231);
or U3293 (N_3293,N_3182,N_3017);
xnor U3294 (N_3294,N_3087,N_3096);
or U3295 (N_3295,N_3014,N_3110);
and U3296 (N_3296,N_3155,N_3180);
nand U3297 (N_3297,N_3131,N_3209);
nor U3298 (N_3298,N_3029,N_3038);
nand U3299 (N_3299,N_3174,N_3198);
xnor U3300 (N_3300,N_3020,N_3201);
and U3301 (N_3301,N_3199,N_3063);
nand U3302 (N_3302,N_3176,N_3184);
or U3303 (N_3303,N_3100,N_3012);
nor U3304 (N_3304,N_3032,N_3120);
and U3305 (N_3305,N_3189,N_3015);
nor U3306 (N_3306,N_3051,N_3006);
nand U3307 (N_3307,N_3187,N_3147);
and U3308 (N_3308,N_3141,N_3197);
nor U3309 (N_3309,N_3076,N_3045);
nand U3310 (N_3310,N_3001,N_3211);
nor U3311 (N_3311,N_3161,N_3000);
xor U3312 (N_3312,N_3085,N_3126);
nor U3313 (N_3313,N_3196,N_3049);
xnor U3314 (N_3314,N_3091,N_3244);
nand U3315 (N_3315,N_3183,N_3065);
xnor U3316 (N_3316,N_3039,N_3089);
or U3317 (N_3317,N_3226,N_3245);
or U3318 (N_3318,N_3033,N_3008);
and U3319 (N_3319,N_3152,N_3179);
nand U3320 (N_3320,N_3052,N_3193);
nand U3321 (N_3321,N_3059,N_3203);
nand U3322 (N_3322,N_3237,N_3210);
xor U3323 (N_3323,N_3083,N_3178);
xor U3324 (N_3324,N_3212,N_3043);
and U3325 (N_3325,N_3070,N_3047);
and U3326 (N_3326,N_3229,N_3240);
or U3327 (N_3327,N_3230,N_3243);
or U3328 (N_3328,N_3106,N_3117);
and U3329 (N_3329,N_3218,N_3208);
and U3330 (N_3330,N_3118,N_3066);
and U3331 (N_3331,N_3090,N_3207);
xnor U3332 (N_3332,N_3018,N_3227);
nand U3333 (N_3333,N_3173,N_3078);
nor U3334 (N_3334,N_3129,N_3115);
or U3335 (N_3335,N_3222,N_3154);
nor U3336 (N_3336,N_3130,N_3247);
xor U3337 (N_3337,N_3133,N_3036);
or U3338 (N_3338,N_3158,N_3163);
or U3339 (N_3339,N_3084,N_3224);
nor U3340 (N_3340,N_3024,N_3069);
nand U3341 (N_3341,N_3175,N_3004);
or U3342 (N_3342,N_3071,N_3109);
and U3343 (N_3343,N_3042,N_3082);
nor U3344 (N_3344,N_3058,N_3142);
xnor U3345 (N_3345,N_3056,N_3007);
and U3346 (N_3346,N_3093,N_3035);
and U3347 (N_3347,N_3021,N_3169);
nand U3348 (N_3348,N_3200,N_3044);
or U3349 (N_3349,N_3138,N_3140);
nor U3350 (N_3350,N_3055,N_3054);
nand U3351 (N_3351,N_3034,N_3011);
xnor U3352 (N_3352,N_3116,N_3022);
xnor U3353 (N_3353,N_3156,N_3220);
or U3354 (N_3354,N_3064,N_3114);
xor U3355 (N_3355,N_3186,N_3041);
or U3356 (N_3356,N_3095,N_3223);
xor U3357 (N_3357,N_3088,N_3030);
nor U3358 (N_3358,N_3023,N_3136);
nor U3359 (N_3359,N_3104,N_3153);
xor U3360 (N_3360,N_3105,N_3217);
and U3361 (N_3361,N_3027,N_3134);
and U3362 (N_3362,N_3111,N_3050);
nor U3363 (N_3363,N_3177,N_3124);
xnor U3364 (N_3364,N_3168,N_3213);
or U3365 (N_3365,N_3053,N_3108);
nand U3366 (N_3366,N_3225,N_3101);
nand U3367 (N_3367,N_3013,N_3172);
or U3368 (N_3368,N_3081,N_3103);
nand U3369 (N_3369,N_3098,N_3157);
xnor U3370 (N_3370,N_3031,N_3009);
xnor U3371 (N_3371,N_3094,N_3122);
and U3372 (N_3372,N_3205,N_3112);
xnor U3373 (N_3373,N_3148,N_3246);
nand U3374 (N_3374,N_3003,N_3073);
xor U3375 (N_3375,N_3233,N_3188);
or U3376 (N_3376,N_3132,N_3072);
and U3377 (N_3377,N_3036,N_3247);
nand U3378 (N_3378,N_3133,N_3193);
nand U3379 (N_3379,N_3036,N_3013);
nand U3380 (N_3380,N_3074,N_3209);
nand U3381 (N_3381,N_3146,N_3044);
nand U3382 (N_3382,N_3039,N_3042);
nor U3383 (N_3383,N_3144,N_3075);
xor U3384 (N_3384,N_3120,N_3179);
xnor U3385 (N_3385,N_3174,N_3123);
and U3386 (N_3386,N_3041,N_3119);
nor U3387 (N_3387,N_3135,N_3028);
xor U3388 (N_3388,N_3220,N_3029);
nor U3389 (N_3389,N_3073,N_3039);
nand U3390 (N_3390,N_3001,N_3233);
nor U3391 (N_3391,N_3180,N_3194);
xnor U3392 (N_3392,N_3224,N_3242);
or U3393 (N_3393,N_3059,N_3174);
and U3394 (N_3394,N_3041,N_3203);
and U3395 (N_3395,N_3088,N_3000);
or U3396 (N_3396,N_3248,N_3241);
or U3397 (N_3397,N_3172,N_3195);
and U3398 (N_3398,N_3144,N_3016);
and U3399 (N_3399,N_3130,N_3086);
xor U3400 (N_3400,N_3155,N_3156);
xnor U3401 (N_3401,N_3077,N_3221);
nand U3402 (N_3402,N_3243,N_3245);
nand U3403 (N_3403,N_3236,N_3123);
nor U3404 (N_3404,N_3168,N_3167);
nor U3405 (N_3405,N_3163,N_3127);
nor U3406 (N_3406,N_3105,N_3082);
nor U3407 (N_3407,N_3107,N_3041);
nor U3408 (N_3408,N_3194,N_3181);
nand U3409 (N_3409,N_3196,N_3179);
nand U3410 (N_3410,N_3148,N_3173);
xnor U3411 (N_3411,N_3059,N_3222);
nor U3412 (N_3412,N_3235,N_3034);
and U3413 (N_3413,N_3161,N_3182);
xor U3414 (N_3414,N_3223,N_3249);
nor U3415 (N_3415,N_3199,N_3235);
nand U3416 (N_3416,N_3185,N_3193);
xor U3417 (N_3417,N_3227,N_3086);
nand U3418 (N_3418,N_3079,N_3001);
or U3419 (N_3419,N_3153,N_3070);
nor U3420 (N_3420,N_3113,N_3115);
xnor U3421 (N_3421,N_3191,N_3038);
and U3422 (N_3422,N_3064,N_3247);
and U3423 (N_3423,N_3118,N_3091);
xnor U3424 (N_3424,N_3036,N_3205);
nand U3425 (N_3425,N_3123,N_3213);
xor U3426 (N_3426,N_3150,N_3121);
xor U3427 (N_3427,N_3062,N_3078);
or U3428 (N_3428,N_3050,N_3006);
xnor U3429 (N_3429,N_3148,N_3114);
and U3430 (N_3430,N_3158,N_3114);
xnor U3431 (N_3431,N_3170,N_3063);
nor U3432 (N_3432,N_3185,N_3090);
xor U3433 (N_3433,N_3001,N_3104);
nor U3434 (N_3434,N_3128,N_3113);
nand U3435 (N_3435,N_3202,N_3074);
nand U3436 (N_3436,N_3002,N_3133);
nor U3437 (N_3437,N_3106,N_3115);
nand U3438 (N_3438,N_3132,N_3158);
nand U3439 (N_3439,N_3161,N_3014);
or U3440 (N_3440,N_3047,N_3247);
nand U3441 (N_3441,N_3219,N_3137);
xor U3442 (N_3442,N_3083,N_3044);
nor U3443 (N_3443,N_3182,N_3239);
and U3444 (N_3444,N_3231,N_3185);
and U3445 (N_3445,N_3154,N_3115);
nand U3446 (N_3446,N_3132,N_3065);
or U3447 (N_3447,N_3064,N_3096);
nand U3448 (N_3448,N_3139,N_3166);
or U3449 (N_3449,N_3034,N_3071);
nor U3450 (N_3450,N_3000,N_3206);
nor U3451 (N_3451,N_3012,N_3074);
nor U3452 (N_3452,N_3092,N_3063);
or U3453 (N_3453,N_3072,N_3060);
and U3454 (N_3454,N_3195,N_3227);
xor U3455 (N_3455,N_3050,N_3192);
xnor U3456 (N_3456,N_3071,N_3065);
or U3457 (N_3457,N_3073,N_3214);
or U3458 (N_3458,N_3060,N_3221);
xnor U3459 (N_3459,N_3237,N_3218);
nand U3460 (N_3460,N_3128,N_3001);
xor U3461 (N_3461,N_3165,N_3120);
and U3462 (N_3462,N_3017,N_3115);
and U3463 (N_3463,N_3197,N_3129);
or U3464 (N_3464,N_3200,N_3107);
xor U3465 (N_3465,N_3079,N_3058);
or U3466 (N_3466,N_3150,N_3243);
or U3467 (N_3467,N_3020,N_3144);
or U3468 (N_3468,N_3128,N_3175);
nor U3469 (N_3469,N_3076,N_3100);
nor U3470 (N_3470,N_3030,N_3071);
or U3471 (N_3471,N_3216,N_3069);
or U3472 (N_3472,N_3193,N_3215);
or U3473 (N_3473,N_3029,N_3060);
nor U3474 (N_3474,N_3155,N_3223);
xnor U3475 (N_3475,N_3037,N_3080);
nor U3476 (N_3476,N_3221,N_3039);
nor U3477 (N_3477,N_3125,N_3118);
or U3478 (N_3478,N_3027,N_3025);
xnor U3479 (N_3479,N_3196,N_3147);
and U3480 (N_3480,N_3221,N_3122);
or U3481 (N_3481,N_3129,N_3097);
or U3482 (N_3482,N_3035,N_3044);
and U3483 (N_3483,N_3029,N_3076);
and U3484 (N_3484,N_3015,N_3050);
nor U3485 (N_3485,N_3160,N_3072);
nand U3486 (N_3486,N_3020,N_3143);
and U3487 (N_3487,N_3153,N_3182);
nor U3488 (N_3488,N_3028,N_3142);
xor U3489 (N_3489,N_3145,N_3221);
and U3490 (N_3490,N_3194,N_3187);
xor U3491 (N_3491,N_3216,N_3086);
nor U3492 (N_3492,N_3221,N_3231);
nand U3493 (N_3493,N_3221,N_3123);
nand U3494 (N_3494,N_3033,N_3038);
xnor U3495 (N_3495,N_3154,N_3237);
xor U3496 (N_3496,N_3145,N_3176);
and U3497 (N_3497,N_3079,N_3135);
nor U3498 (N_3498,N_3247,N_3054);
nor U3499 (N_3499,N_3134,N_3126);
or U3500 (N_3500,N_3458,N_3393);
nand U3501 (N_3501,N_3308,N_3442);
or U3502 (N_3502,N_3432,N_3498);
nor U3503 (N_3503,N_3348,N_3364);
xor U3504 (N_3504,N_3335,N_3401);
or U3505 (N_3505,N_3396,N_3254);
nand U3506 (N_3506,N_3324,N_3457);
nand U3507 (N_3507,N_3384,N_3270);
nor U3508 (N_3508,N_3456,N_3399);
and U3509 (N_3509,N_3259,N_3444);
nor U3510 (N_3510,N_3321,N_3279);
xor U3511 (N_3511,N_3451,N_3311);
nor U3512 (N_3512,N_3306,N_3433);
xor U3513 (N_3513,N_3405,N_3356);
nor U3514 (N_3514,N_3411,N_3302);
nor U3515 (N_3515,N_3459,N_3377);
xnor U3516 (N_3516,N_3414,N_3470);
xnor U3517 (N_3517,N_3445,N_3272);
and U3518 (N_3518,N_3469,N_3395);
nand U3519 (N_3519,N_3253,N_3331);
xnor U3520 (N_3520,N_3305,N_3391);
nand U3521 (N_3521,N_3298,N_3278);
and U3522 (N_3522,N_3256,N_3418);
and U3523 (N_3523,N_3425,N_3483);
nand U3524 (N_3524,N_3275,N_3338);
and U3525 (N_3525,N_3413,N_3334);
nand U3526 (N_3526,N_3251,N_3443);
or U3527 (N_3527,N_3441,N_3368);
nor U3528 (N_3528,N_3255,N_3388);
xnor U3529 (N_3529,N_3427,N_3492);
or U3530 (N_3530,N_3477,N_3261);
nor U3531 (N_3531,N_3467,N_3271);
or U3532 (N_3532,N_3354,N_3472);
xor U3533 (N_3533,N_3361,N_3428);
xor U3534 (N_3534,N_3318,N_3314);
nand U3535 (N_3535,N_3316,N_3408);
nor U3536 (N_3536,N_3385,N_3468);
xor U3537 (N_3537,N_3336,N_3479);
nand U3538 (N_3538,N_3297,N_3339);
or U3539 (N_3539,N_3319,N_3486);
and U3540 (N_3540,N_3285,N_3389);
nor U3541 (N_3541,N_3283,N_3482);
nand U3542 (N_3542,N_3478,N_3287);
nor U3543 (N_3543,N_3375,N_3410);
or U3544 (N_3544,N_3351,N_3474);
or U3545 (N_3545,N_3415,N_3439);
nor U3546 (N_3546,N_3344,N_3370);
nor U3547 (N_3547,N_3400,N_3371);
and U3548 (N_3548,N_3485,N_3455);
nand U3549 (N_3549,N_3258,N_3326);
xor U3550 (N_3550,N_3440,N_3394);
nor U3551 (N_3551,N_3471,N_3496);
or U3552 (N_3552,N_3277,N_3494);
or U3553 (N_3553,N_3299,N_3480);
or U3554 (N_3554,N_3355,N_3269);
and U3555 (N_3555,N_3390,N_3363);
or U3556 (N_3556,N_3295,N_3490);
nand U3557 (N_3557,N_3450,N_3296);
nand U3558 (N_3558,N_3429,N_3322);
nor U3559 (N_3559,N_3362,N_3290);
xor U3560 (N_3560,N_3497,N_3487);
and U3561 (N_3561,N_3262,N_3381);
xnor U3562 (N_3562,N_3421,N_3300);
and U3563 (N_3563,N_3293,N_3280);
or U3564 (N_3564,N_3309,N_3317);
or U3565 (N_3565,N_3406,N_3260);
xor U3566 (N_3566,N_3378,N_3423);
nand U3567 (N_3567,N_3284,N_3349);
nand U3568 (N_3568,N_3347,N_3386);
xor U3569 (N_3569,N_3464,N_3301);
nand U3570 (N_3570,N_3449,N_3426);
xnor U3571 (N_3571,N_3397,N_3422);
or U3572 (N_3572,N_3430,N_3304);
xor U3573 (N_3573,N_3447,N_3332);
nor U3574 (N_3574,N_3346,N_3343);
and U3575 (N_3575,N_3453,N_3294);
or U3576 (N_3576,N_3446,N_3327);
or U3577 (N_3577,N_3436,N_3267);
nand U3578 (N_3578,N_3281,N_3465);
xor U3579 (N_3579,N_3367,N_3360);
nor U3580 (N_3580,N_3357,N_3376);
and U3581 (N_3581,N_3374,N_3372);
xor U3582 (N_3582,N_3424,N_3268);
nand U3583 (N_3583,N_3475,N_3291);
nand U3584 (N_3584,N_3263,N_3412);
xor U3585 (N_3585,N_3489,N_3387);
nor U3586 (N_3586,N_3476,N_3491);
nor U3587 (N_3587,N_3473,N_3448);
and U3588 (N_3588,N_3392,N_3416);
and U3589 (N_3589,N_3274,N_3438);
or U3590 (N_3590,N_3452,N_3265);
or U3591 (N_3591,N_3481,N_3409);
nor U3592 (N_3592,N_3312,N_3325);
or U3593 (N_3593,N_3350,N_3454);
nand U3594 (N_3594,N_3328,N_3461);
nor U3595 (N_3595,N_3419,N_3329);
and U3596 (N_3596,N_3403,N_3365);
and U3597 (N_3597,N_3286,N_3330);
and U3598 (N_3598,N_3323,N_3250);
nor U3599 (N_3599,N_3417,N_3257);
nand U3600 (N_3600,N_3358,N_3380);
nand U3601 (N_3601,N_3379,N_3431);
or U3602 (N_3602,N_3266,N_3289);
nor U3603 (N_3603,N_3398,N_3288);
nor U3604 (N_3604,N_3462,N_3282);
or U3605 (N_3605,N_3342,N_3320);
nand U3606 (N_3606,N_3313,N_3407);
xnor U3607 (N_3607,N_3359,N_3495);
and U3608 (N_3608,N_3273,N_3337);
or U3609 (N_3609,N_3276,N_3420);
nor U3610 (N_3610,N_3310,N_3466);
and U3611 (N_3611,N_3434,N_3383);
nor U3612 (N_3612,N_3369,N_3402);
or U3613 (N_3613,N_3382,N_3352);
or U3614 (N_3614,N_3264,N_3315);
and U3615 (N_3615,N_3345,N_3252);
xor U3616 (N_3616,N_3366,N_3303);
nand U3617 (N_3617,N_3340,N_3488);
nand U3618 (N_3618,N_3292,N_3484);
xnor U3619 (N_3619,N_3404,N_3437);
nor U3620 (N_3620,N_3341,N_3353);
nand U3621 (N_3621,N_3499,N_3333);
nor U3622 (N_3622,N_3435,N_3493);
nor U3623 (N_3623,N_3463,N_3373);
or U3624 (N_3624,N_3460,N_3307);
or U3625 (N_3625,N_3275,N_3281);
and U3626 (N_3626,N_3488,N_3404);
nor U3627 (N_3627,N_3353,N_3478);
nand U3628 (N_3628,N_3402,N_3394);
nor U3629 (N_3629,N_3393,N_3344);
or U3630 (N_3630,N_3364,N_3436);
and U3631 (N_3631,N_3499,N_3267);
or U3632 (N_3632,N_3370,N_3419);
and U3633 (N_3633,N_3458,N_3386);
and U3634 (N_3634,N_3364,N_3310);
or U3635 (N_3635,N_3360,N_3481);
and U3636 (N_3636,N_3373,N_3488);
and U3637 (N_3637,N_3352,N_3475);
nand U3638 (N_3638,N_3488,N_3280);
nand U3639 (N_3639,N_3310,N_3330);
nor U3640 (N_3640,N_3390,N_3282);
xnor U3641 (N_3641,N_3293,N_3276);
nand U3642 (N_3642,N_3427,N_3482);
and U3643 (N_3643,N_3281,N_3295);
nor U3644 (N_3644,N_3368,N_3334);
and U3645 (N_3645,N_3312,N_3341);
nor U3646 (N_3646,N_3303,N_3318);
nor U3647 (N_3647,N_3262,N_3430);
nand U3648 (N_3648,N_3452,N_3420);
or U3649 (N_3649,N_3491,N_3464);
nand U3650 (N_3650,N_3422,N_3393);
nand U3651 (N_3651,N_3325,N_3336);
nand U3652 (N_3652,N_3446,N_3465);
or U3653 (N_3653,N_3373,N_3450);
xor U3654 (N_3654,N_3314,N_3361);
and U3655 (N_3655,N_3269,N_3486);
and U3656 (N_3656,N_3337,N_3351);
and U3657 (N_3657,N_3353,N_3321);
xor U3658 (N_3658,N_3441,N_3331);
nand U3659 (N_3659,N_3496,N_3460);
and U3660 (N_3660,N_3366,N_3309);
and U3661 (N_3661,N_3341,N_3383);
and U3662 (N_3662,N_3357,N_3434);
and U3663 (N_3663,N_3425,N_3342);
nand U3664 (N_3664,N_3287,N_3415);
nor U3665 (N_3665,N_3449,N_3268);
nand U3666 (N_3666,N_3478,N_3260);
nand U3667 (N_3667,N_3456,N_3448);
nor U3668 (N_3668,N_3284,N_3490);
nand U3669 (N_3669,N_3384,N_3484);
or U3670 (N_3670,N_3453,N_3319);
nor U3671 (N_3671,N_3269,N_3348);
and U3672 (N_3672,N_3372,N_3381);
and U3673 (N_3673,N_3442,N_3343);
and U3674 (N_3674,N_3401,N_3293);
xnor U3675 (N_3675,N_3496,N_3383);
nor U3676 (N_3676,N_3313,N_3269);
and U3677 (N_3677,N_3477,N_3499);
nor U3678 (N_3678,N_3321,N_3299);
nor U3679 (N_3679,N_3365,N_3489);
or U3680 (N_3680,N_3450,N_3477);
xnor U3681 (N_3681,N_3482,N_3478);
and U3682 (N_3682,N_3347,N_3266);
nand U3683 (N_3683,N_3342,N_3436);
nand U3684 (N_3684,N_3358,N_3283);
or U3685 (N_3685,N_3341,N_3339);
nand U3686 (N_3686,N_3387,N_3439);
nand U3687 (N_3687,N_3408,N_3403);
xor U3688 (N_3688,N_3431,N_3270);
nor U3689 (N_3689,N_3461,N_3434);
xnor U3690 (N_3690,N_3284,N_3369);
xnor U3691 (N_3691,N_3385,N_3487);
nand U3692 (N_3692,N_3346,N_3442);
and U3693 (N_3693,N_3438,N_3339);
nor U3694 (N_3694,N_3428,N_3332);
xnor U3695 (N_3695,N_3363,N_3326);
nand U3696 (N_3696,N_3405,N_3443);
xnor U3697 (N_3697,N_3373,N_3425);
xor U3698 (N_3698,N_3457,N_3468);
nand U3699 (N_3699,N_3446,N_3279);
nand U3700 (N_3700,N_3260,N_3407);
xor U3701 (N_3701,N_3345,N_3358);
xnor U3702 (N_3702,N_3314,N_3279);
nor U3703 (N_3703,N_3386,N_3402);
or U3704 (N_3704,N_3379,N_3473);
and U3705 (N_3705,N_3327,N_3299);
and U3706 (N_3706,N_3391,N_3395);
nand U3707 (N_3707,N_3358,N_3315);
and U3708 (N_3708,N_3390,N_3456);
nand U3709 (N_3709,N_3361,N_3393);
and U3710 (N_3710,N_3476,N_3380);
and U3711 (N_3711,N_3417,N_3433);
nor U3712 (N_3712,N_3455,N_3467);
nand U3713 (N_3713,N_3398,N_3424);
or U3714 (N_3714,N_3441,N_3256);
and U3715 (N_3715,N_3372,N_3308);
nor U3716 (N_3716,N_3416,N_3383);
or U3717 (N_3717,N_3322,N_3358);
nand U3718 (N_3718,N_3418,N_3380);
or U3719 (N_3719,N_3290,N_3395);
or U3720 (N_3720,N_3311,N_3487);
or U3721 (N_3721,N_3358,N_3485);
or U3722 (N_3722,N_3387,N_3391);
and U3723 (N_3723,N_3343,N_3347);
and U3724 (N_3724,N_3433,N_3492);
xnor U3725 (N_3725,N_3458,N_3434);
or U3726 (N_3726,N_3438,N_3385);
and U3727 (N_3727,N_3382,N_3480);
nor U3728 (N_3728,N_3307,N_3293);
nand U3729 (N_3729,N_3364,N_3373);
nand U3730 (N_3730,N_3304,N_3382);
xnor U3731 (N_3731,N_3354,N_3370);
or U3732 (N_3732,N_3289,N_3409);
or U3733 (N_3733,N_3495,N_3387);
nand U3734 (N_3734,N_3430,N_3475);
and U3735 (N_3735,N_3305,N_3339);
nand U3736 (N_3736,N_3438,N_3288);
or U3737 (N_3737,N_3336,N_3328);
or U3738 (N_3738,N_3456,N_3468);
nor U3739 (N_3739,N_3426,N_3295);
nand U3740 (N_3740,N_3400,N_3450);
nor U3741 (N_3741,N_3430,N_3259);
nor U3742 (N_3742,N_3430,N_3251);
and U3743 (N_3743,N_3376,N_3406);
and U3744 (N_3744,N_3256,N_3314);
and U3745 (N_3745,N_3421,N_3396);
nand U3746 (N_3746,N_3440,N_3447);
and U3747 (N_3747,N_3355,N_3421);
and U3748 (N_3748,N_3261,N_3367);
nor U3749 (N_3749,N_3267,N_3402);
or U3750 (N_3750,N_3680,N_3734);
nor U3751 (N_3751,N_3511,N_3719);
nor U3752 (N_3752,N_3577,N_3560);
and U3753 (N_3753,N_3733,N_3564);
nand U3754 (N_3754,N_3662,N_3715);
and U3755 (N_3755,N_3697,N_3693);
and U3756 (N_3756,N_3723,N_3724);
xor U3757 (N_3757,N_3614,N_3544);
or U3758 (N_3758,N_3574,N_3519);
and U3759 (N_3759,N_3710,N_3507);
and U3760 (N_3760,N_3513,N_3626);
nor U3761 (N_3761,N_3656,N_3539);
nor U3762 (N_3762,N_3637,N_3592);
nand U3763 (N_3763,N_3565,N_3527);
or U3764 (N_3764,N_3669,N_3631);
xor U3765 (N_3765,N_3543,N_3714);
or U3766 (N_3766,N_3546,N_3573);
xor U3767 (N_3767,N_3562,N_3506);
or U3768 (N_3768,N_3602,N_3595);
xor U3769 (N_3769,N_3738,N_3736);
nand U3770 (N_3770,N_3533,N_3709);
or U3771 (N_3771,N_3745,N_3650);
or U3772 (N_3772,N_3705,N_3643);
and U3773 (N_3773,N_3532,N_3717);
xnor U3774 (N_3774,N_3557,N_3561);
or U3775 (N_3775,N_3605,N_3747);
xnor U3776 (N_3776,N_3629,N_3538);
or U3777 (N_3777,N_3608,N_3508);
and U3778 (N_3778,N_3676,N_3694);
xor U3779 (N_3779,N_3516,N_3699);
xor U3780 (N_3780,N_3526,N_3661);
nor U3781 (N_3781,N_3563,N_3684);
or U3782 (N_3782,N_3665,N_3703);
nor U3783 (N_3783,N_3593,N_3590);
xor U3784 (N_3784,N_3581,N_3702);
and U3785 (N_3785,N_3673,N_3691);
xor U3786 (N_3786,N_3728,N_3525);
and U3787 (N_3787,N_3512,N_3580);
or U3788 (N_3788,N_3555,N_3554);
xor U3789 (N_3789,N_3542,N_3531);
and U3790 (N_3790,N_3737,N_3571);
and U3791 (N_3791,N_3594,N_3576);
or U3792 (N_3792,N_3514,N_3686);
nor U3793 (N_3793,N_3541,N_3657);
and U3794 (N_3794,N_3628,N_3748);
xor U3795 (N_3795,N_3741,N_3729);
and U3796 (N_3796,N_3722,N_3569);
or U3797 (N_3797,N_3718,N_3599);
and U3798 (N_3798,N_3647,N_3721);
and U3799 (N_3799,N_3547,N_3585);
nand U3800 (N_3800,N_3621,N_3671);
nor U3801 (N_3801,N_3720,N_3652);
nand U3802 (N_3802,N_3708,N_3627);
xor U3803 (N_3803,N_3730,N_3640);
nor U3804 (N_3804,N_3536,N_3530);
or U3805 (N_3805,N_3504,N_3632);
nor U3806 (N_3806,N_3505,N_3591);
nor U3807 (N_3807,N_3666,N_3653);
and U3808 (N_3808,N_3683,N_3655);
and U3809 (N_3809,N_3687,N_3500);
nand U3810 (N_3810,N_3534,N_3634);
or U3811 (N_3811,N_3617,N_3510);
or U3812 (N_3812,N_3735,N_3550);
nand U3813 (N_3813,N_3528,N_3559);
or U3814 (N_3814,N_3537,N_3623);
xnor U3815 (N_3815,N_3579,N_3688);
and U3816 (N_3816,N_3556,N_3636);
and U3817 (N_3817,N_3586,N_3567);
nor U3818 (N_3818,N_3551,N_3578);
xor U3819 (N_3819,N_3520,N_3712);
nand U3820 (N_3820,N_3695,N_3746);
or U3821 (N_3821,N_3700,N_3558);
or U3822 (N_3822,N_3611,N_3535);
or U3823 (N_3823,N_3641,N_3707);
nand U3824 (N_3824,N_3690,N_3692);
or U3825 (N_3825,N_3596,N_3587);
nor U3826 (N_3826,N_3615,N_3501);
and U3827 (N_3827,N_3570,N_3610);
or U3828 (N_3828,N_3606,N_3743);
or U3829 (N_3829,N_3624,N_3619);
xor U3830 (N_3830,N_3604,N_3646);
and U3831 (N_3831,N_3659,N_3701);
nand U3832 (N_3832,N_3706,N_3716);
nor U3833 (N_3833,N_3622,N_3568);
xor U3834 (N_3834,N_3613,N_3521);
nor U3835 (N_3835,N_3553,N_3612);
nor U3836 (N_3836,N_3545,N_3658);
nor U3837 (N_3837,N_3725,N_3618);
and U3838 (N_3838,N_3654,N_3698);
nand U3839 (N_3839,N_3682,N_3502);
and U3840 (N_3840,N_3667,N_3552);
nor U3841 (N_3841,N_3515,N_3549);
and U3842 (N_3842,N_3645,N_3696);
or U3843 (N_3843,N_3675,N_3677);
and U3844 (N_3844,N_3727,N_3749);
and U3845 (N_3845,N_3517,N_3670);
nand U3846 (N_3846,N_3739,N_3660);
and U3847 (N_3847,N_3704,N_3731);
and U3848 (N_3848,N_3523,N_3664);
or U3849 (N_3849,N_3548,N_3678);
nor U3850 (N_3850,N_3651,N_3620);
nor U3851 (N_3851,N_3522,N_3589);
nand U3852 (N_3852,N_3597,N_3588);
nor U3853 (N_3853,N_3524,N_3607);
xor U3854 (N_3854,N_3679,N_3726);
nand U3855 (N_3855,N_3711,N_3638);
nand U3856 (N_3856,N_3649,N_3601);
and U3857 (N_3857,N_3732,N_3648);
or U3858 (N_3858,N_3572,N_3616);
or U3859 (N_3859,N_3598,N_3509);
nor U3860 (N_3860,N_3740,N_3529);
nand U3861 (N_3861,N_3644,N_3540);
and U3862 (N_3862,N_3630,N_3635);
nor U3863 (N_3863,N_3503,N_3583);
or U3864 (N_3864,N_3674,N_3609);
xnor U3865 (N_3865,N_3582,N_3663);
xor U3866 (N_3866,N_3685,N_3742);
or U3867 (N_3867,N_3713,N_3625);
and U3868 (N_3868,N_3689,N_3633);
nor U3869 (N_3869,N_3668,N_3575);
nor U3870 (N_3870,N_3518,N_3744);
xnor U3871 (N_3871,N_3603,N_3566);
nand U3872 (N_3872,N_3600,N_3584);
and U3873 (N_3873,N_3639,N_3681);
nor U3874 (N_3874,N_3642,N_3672);
and U3875 (N_3875,N_3549,N_3635);
and U3876 (N_3876,N_3605,N_3722);
nor U3877 (N_3877,N_3592,N_3588);
or U3878 (N_3878,N_3730,N_3552);
nand U3879 (N_3879,N_3692,N_3720);
xor U3880 (N_3880,N_3574,N_3658);
and U3881 (N_3881,N_3655,N_3552);
xor U3882 (N_3882,N_3687,N_3688);
nand U3883 (N_3883,N_3530,N_3574);
nand U3884 (N_3884,N_3681,N_3631);
and U3885 (N_3885,N_3656,N_3658);
xnor U3886 (N_3886,N_3534,N_3730);
nor U3887 (N_3887,N_3723,N_3504);
and U3888 (N_3888,N_3653,N_3734);
xor U3889 (N_3889,N_3654,N_3549);
and U3890 (N_3890,N_3545,N_3523);
or U3891 (N_3891,N_3638,N_3561);
xnor U3892 (N_3892,N_3608,N_3720);
or U3893 (N_3893,N_3696,N_3639);
and U3894 (N_3894,N_3608,N_3685);
and U3895 (N_3895,N_3588,N_3603);
xnor U3896 (N_3896,N_3534,N_3722);
and U3897 (N_3897,N_3747,N_3536);
xnor U3898 (N_3898,N_3715,N_3670);
nand U3899 (N_3899,N_3715,N_3569);
and U3900 (N_3900,N_3573,N_3704);
xnor U3901 (N_3901,N_3592,N_3583);
and U3902 (N_3902,N_3682,N_3619);
and U3903 (N_3903,N_3734,N_3541);
or U3904 (N_3904,N_3634,N_3590);
nor U3905 (N_3905,N_3642,N_3671);
nand U3906 (N_3906,N_3632,N_3712);
and U3907 (N_3907,N_3534,N_3512);
and U3908 (N_3908,N_3505,N_3595);
xnor U3909 (N_3909,N_3675,N_3682);
and U3910 (N_3910,N_3604,N_3644);
xnor U3911 (N_3911,N_3658,N_3635);
xor U3912 (N_3912,N_3549,N_3556);
and U3913 (N_3913,N_3672,N_3502);
nand U3914 (N_3914,N_3663,N_3542);
and U3915 (N_3915,N_3721,N_3644);
or U3916 (N_3916,N_3668,N_3521);
and U3917 (N_3917,N_3735,N_3541);
xor U3918 (N_3918,N_3575,N_3652);
nor U3919 (N_3919,N_3602,N_3633);
nor U3920 (N_3920,N_3537,N_3654);
and U3921 (N_3921,N_3684,N_3673);
xnor U3922 (N_3922,N_3592,N_3691);
xnor U3923 (N_3923,N_3744,N_3678);
and U3924 (N_3924,N_3706,N_3590);
nand U3925 (N_3925,N_3648,N_3613);
nand U3926 (N_3926,N_3649,N_3515);
and U3927 (N_3927,N_3693,N_3592);
nor U3928 (N_3928,N_3707,N_3573);
or U3929 (N_3929,N_3600,N_3599);
xor U3930 (N_3930,N_3650,N_3713);
and U3931 (N_3931,N_3503,N_3617);
and U3932 (N_3932,N_3611,N_3681);
or U3933 (N_3933,N_3746,N_3522);
nor U3934 (N_3934,N_3576,N_3527);
xor U3935 (N_3935,N_3728,N_3748);
nor U3936 (N_3936,N_3671,N_3726);
or U3937 (N_3937,N_3563,N_3528);
xnor U3938 (N_3938,N_3540,N_3515);
and U3939 (N_3939,N_3625,N_3673);
xnor U3940 (N_3940,N_3736,N_3673);
nand U3941 (N_3941,N_3744,N_3680);
and U3942 (N_3942,N_3748,N_3734);
nor U3943 (N_3943,N_3654,N_3509);
nor U3944 (N_3944,N_3642,N_3670);
and U3945 (N_3945,N_3513,N_3540);
and U3946 (N_3946,N_3691,N_3711);
nor U3947 (N_3947,N_3640,N_3581);
or U3948 (N_3948,N_3516,N_3578);
xor U3949 (N_3949,N_3508,N_3602);
nand U3950 (N_3950,N_3734,N_3698);
xnor U3951 (N_3951,N_3743,N_3529);
nor U3952 (N_3952,N_3625,N_3526);
or U3953 (N_3953,N_3698,N_3677);
or U3954 (N_3954,N_3641,N_3566);
nand U3955 (N_3955,N_3535,N_3536);
xor U3956 (N_3956,N_3642,N_3680);
and U3957 (N_3957,N_3565,N_3520);
nand U3958 (N_3958,N_3732,N_3610);
nor U3959 (N_3959,N_3582,N_3681);
or U3960 (N_3960,N_3644,N_3646);
xnor U3961 (N_3961,N_3638,N_3587);
xor U3962 (N_3962,N_3724,N_3656);
or U3963 (N_3963,N_3557,N_3520);
nor U3964 (N_3964,N_3636,N_3709);
nor U3965 (N_3965,N_3713,N_3608);
and U3966 (N_3966,N_3735,N_3671);
nand U3967 (N_3967,N_3679,N_3544);
xor U3968 (N_3968,N_3579,N_3712);
nand U3969 (N_3969,N_3622,N_3726);
nand U3970 (N_3970,N_3517,N_3746);
or U3971 (N_3971,N_3541,N_3717);
xor U3972 (N_3972,N_3503,N_3680);
or U3973 (N_3973,N_3571,N_3725);
nand U3974 (N_3974,N_3674,N_3657);
and U3975 (N_3975,N_3663,N_3507);
nor U3976 (N_3976,N_3576,N_3672);
nand U3977 (N_3977,N_3509,N_3581);
and U3978 (N_3978,N_3655,N_3719);
and U3979 (N_3979,N_3681,N_3703);
or U3980 (N_3980,N_3508,N_3572);
nand U3981 (N_3981,N_3572,N_3520);
nor U3982 (N_3982,N_3630,N_3732);
xor U3983 (N_3983,N_3511,N_3510);
xor U3984 (N_3984,N_3624,N_3512);
or U3985 (N_3985,N_3535,N_3504);
and U3986 (N_3986,N_3529,N_3670);
nand U3987 (N_3987,N_3716,N_3516);
nand U3988 (N_3988,N_3551,N_3532);
or U3989 (N_3989,N_3523,N_3726);
or U3990 (N_3990,N_3633,N_3501);
and U3991 (N_3991,N_3681,N_3744);
xor U3992 (N_3992,N_3696,N_3728);
nand U3993 (N_3993,N_3636,N_3747);
nand U3994 (N_3994,N_3603,N_3695);
or U3995 (N_3995,N_3694,N_3602);
or U3996 (N_3996,N_3717,N_3697);
nand U3997 (N_3997,N_3651,N_3598);
and U3998 (N_3998,N_3701,N_3520);
or U3999 (N_3999,N_3673,N_3592);
nand U4000 (N_4000,N_3802,N_3994);
xnor U4001 (N_4001,N_3837,N_3942);
and U4002 (N_4002,N_3763,N_3900);
and U4003 (N_4003,N_3933,N_3958);
nand U4004 (N_4004,N_3969,N_3953);
or U4005 (N_4005,N_3948,N_3776);
xor U4006 (N_4006,N_3854,N_3916);
or U4007 (N_4007,N_3975,N_3937);
nor U4008 (N_4008,N_3944,N_3805);
nor U4009 (N_4009,N_3964,N_3811);
or U4010 (N_4010,N_3984,N_3795);
xor U4011 (N_4011,N_3810,N_3853);
and U4012 (N_4012,N_3947,N_3989);
nand U4013 (N_4013,N_3777,N_3824);
nor U4014 (N_4014,N_3796,N_3949);
nand U4015 (N_4015,N_3981,N_3825);
or U4016 (N_4016,N_3803,N_3954);
nand U4017 (N_4017,N_3915,N_3914);
nor U4018 (N_4018,N_3771,N_3974);
xnor U4019 (N_4019,N_3875,N_3952);
xnor U4020 (N_4020,N_3898,N_3750);
or U4021 (N_4021,N_3759,N_3813);
xor U4022 (N_4022,N_3926,N_3993);
xor U4023 (N_4023,N_3892,N_3986);
and U4024 (N_4024,N_3979,N_3876);
or U4025 (N_4025,N_3788,N_3864);
or U4026 (N_4026,N_3768,N_3767);
nor U4027 (N_4027,N_3903,N_3826);
or U4028 (N_4028,N_3922,N_3846);
nand U4029 (N_4029,N_3930,N_3770);
nand U4030 (N_4030,N_3762,N_3961);
nor U4031 (N_4031,N_3843,N_3867);
xor U4032 (N_4032,N_3963,N_3834);
or U4033 (N_4033,N_3976,N_3809);
and U4034 (N_4034,N_3753,N_3880);
and U4035 (N_4035,N_3780,N_3857);
xnor U4036 (N_4036,N_3863,N_3800);
nor U4037 (N_4037,N_3869,N_3957);
nand U4038 (N_4038,N_3886,N_3760);
nand U4039 (N_4039,N_3887,N_3983);
and U4040 (N_4040,N_3939,N_3852);
nand U4041 (N_4041,N_3789,N_3787);
xnor U4042 (N_4042,N_3962,N_3924);
and U4043 (N_4043,N_3784,N_3971);
nand U4044 (N_4044,N_3814,N_3917);
xor U4045 (N_4045,N_3932,N_3778);
and U4046 (N_4046,N_3978,N_3833);
or U4047 (N_4047,N_3883,N_3848);
or U4048 (N_4048,N_3782,N_3808);
nor U4049 (N_4049,N_3877,N_3908);
nand U4050 (N_4050,N_3797,N_3791);
or U4051 (N_4051,N_3938,N_3910);
nand U4052 (N_4052,N_3968,N_3835);
xnor U4053 (N_4053,N_3923,N_3856);
and U4054 (N_4054,N_3890,N_3905);
nor U4055 (N_4055,N_3828,N_3827);
and U4056 (N_4056,N_3865,N_3911);
xnor U4057 (N_4057,N_3861,N_3992);
or U4058 (N_4058,N_3966,N_3836);
nand U4059 (N_4059,N_3891,N_3906);
xnor U4060 (N_4060,N_3881,N_3941);
nor U4061 (N_4061,N_3781,N_3985);
or U4062 (N_4062,N_3965,N_3940);
xnor U4063 (N_4063,N_3844,N_3831);
xnor U4064 (N_4064,N_3988,N_3859);
nor U4065 (N_4065,N_3858,N_3847);
or U4066 (N_4066,N_3996,N_3899);
xnor U4067 (N_4067,N_3879,N_3998);
nor U4068 (N_4068,N_3765,N_3956);
or U4069 (N_4069,N_3775,N_3756);
nand U4070 (N_4070,N_3896,N_3871);
and U4071 (N_4071,N_3991,N_3872);
or U4072 (N_4072,N_3866,N_3786);
nor U4073 (N_4073,N_3913,N_3884);
or U4074 (N_4074,N_3918,N_3766);
and U4075 (N_4075,N_3959,N_3987);
or U4076 (N_4076,N_3970,N_3849);
nand U4077 (N_4077,N_3841,N_3845);
or U4078 (N_4078,N_3895,N_3819);
or U4079 (N_4079,N_3928,N_3785);
nand U4080 (N_4080,N_3838,N_3855);
nor U4081 (N_4081,N_3773,N_3794);
nand U4082 (N_4082,N_3874,N_3769);
or U4083 (N_4083,N_3839,N_3904);
xnor U4084 (N_4084,N_3931,N_3820);
xnor U4085 (N_4085,N_3792,N_3885);
or U4086 (N_4086,N_3980,N_3946);
nand U4087 (N_4087,N_3889,N_3882);
nand U4088 (N_4088,N_3967,N_3764);
and U4089 (N_4089,N_3943,N_3868);
nor U4090 (N_4090,N_3757,N_3909);
or U4091 (N_4091,N_3929,N_3862);
nand U4092 (N_4092,N_3888,N_3783);
nor U4093 (N_4093,N_3925,N_3893);
or U4094 (N_4094,N_3793,N_3945);
nand U4095 (N_4095,N_3997,N_3897);
nand U4096 (N_4096,N_3999,N_3935);
and U4097 (N_4097,N_3822,N_3951);
nor U4098 (N_4098,N_3829,N_3818);
xor U4099 (N_4099,N_3921,N_3752);
nor U4100 (N_4100,N_3815,N_3790);
nor U4101 (N_4101,N_3761,N_3842);
or U4102 (N_4102,N_3955,N_3801);
nand U4103 (N_4103,N_3850,N_3798);
nand U4104 (N_4104,N_3973,N_3840);
and U4105 (N_4105,N_3873,N_3817);
or U4106 (N_4106,N_3936,N_3927);
nor U4107 (N_4107,N_3821,N_3812);
and U4108 (N_4108,N_3830,N_3823);
nand U4109 (N_4109,N_3755,N_3754);
and U4110 (N_4110,N_3779,N_3878);
and U4111 (N_4111,N_3774,N_3851);
nor U4112 (N_4112,N_3772,N_3758);
xnor U4113 (N_4113,N_3832,N_3960);
and U4114 (N_4114,N_3870,N_3950);
xnor U4115 (N_4115,N_3799,N_3816);
and U4116 (N_4116,N_3902,N_3990);
and U4117 (N_4117,N_3807,N_3907);
and U4118 (N_4118,N_3751,N_3894);
xor U4119 (N_4119,N_3995,N_3977);
xnor U4120 (N_4120,N_3806,N_3901);
or U4121 (N_4121,N_3920,N_3982);
nor U4122 (N_4122,N_3934,N_3912);
nand U4123 (N_4123,N_3804,N_3860);
xor U4124 (N_4124,N_3972,N_3919);
xnor U4125 (N_4125,N_3861,N_3765);
and U4126 (N_4126,N_3788,N_3750);
or U4127 (N_4127,N_3800,N_3965);
xnor U4128 (N_4128,N_3962,N_3956);
or U4129 (N_4129,N_3997,N_3837);
or U4130 (N_4130,N_3863,N_3972);
nand U4131 (N_4131,N_3790,N_3844);
xor U4132 (N_4132,N_3913,N_3996);
nor U4133 (N_4133,N_3771,N_3798);
xnor U4134 (N_4134,N_3944,N_3854);
xnor U4135 (N_4135,N_3873,N_3981);
or U4136 (N_4136,N_3830,N_3947);
or U4137 (N_4137,N_3995,N_3800);
nor U4138 (N_4138,N_3980,N_3926);
or U4139 (N_4139,N_3976,N_3912);
nand U4140 (N_4140,N_3828,N_3782);
nor U4141 (N_4141,N_3897,N_3829);
or U4142 (N_4142,N_3980,N_3809);
and U4143 (N_4143,N_3798,N_3979);
nand U4144 (N_4144,N_3795,N_3889);
and U4145 (N_4145,N_3762,N_3987);
nand U4146 (N_4146,N_3950,N_3895);
nor U4147 (N_4147,N_3918,N_3945);
nand U4148 (N_4148,N_3910,N_3936);
or U4149 (N_4149,N_3982,N_3768);
and U4150 (N_4150,N_3915,N_3846);
nand U4151 (N_4151,N_3793,N_3960);
nand U4152 (N_4152,N_3820,N_3787);
or U4153 (N_4153,N_3759,N_3809);
nand U4154 (N_4154,N_3884,N_3781);
xnor U4155 (N_4155,N_3958,N_3961);
nand U4156 (N_4156,N_3975,N_3795);
nand U4157 (N_4157,N_3769,N_3774);
xnor U4158 (N_4158,N_3847,N_3888);
or U4159 (N_4159,N_3949,N_3804);
xnor U4160 (N_4160,N_3755,N_3872);
and U4161 (N_4161,N_3901,N_3841);
xnor U4162 (N_4162,N_3899,N_3915);
xnor U4163 (N_4163,N_3936,N_3990);
nor U4164 (N_4164,N_3801,N_3759);
nand U4165 (N_4165,N_3928,N_3966);
nand U4166 (N_4166,N_3867,N_3990);
nor U4167 (N_4167,N_3840,N_3896);
xor U4168 (N_4168,N_3923,N_3933);
nor U4169 (N_4169,N_3764,N_3875);
or U4170 (N_4170,N_3978,N_3754);
nor U4171 (N_4171,N_3759,N_3957);
nor U4172 (N_4172,N_3921,N_3881);
nand U4173 (N_4173,N_3849,N_3958);
and U4174 (N_4174,N_3999,N_3754);
nor U4175 (N_4175,N_3847,N_3950);
and U4176 (N_4176,N_3999,N_3937);
or U4177 (N_4177,N_3814,N_3780);
nor U4178 (N_4178,N_3997,N_3828);
or U4179 (N_4179,N_3876,N_3948);
and U4180 (N_4180,N_3900,N_3786);
nor U4181 (N_4181,N_3905,N_3931);
and U4182 (N_4182,N_3974,N_3996);
nor U4183 (N_4183,N_3947,N_3752);
and U4184 (N_4184,N_3994,N_3828);
or U4185 (N_4185,N_3776,N_3829);
nand U4186 (N_4186,N_3910,N_3980);
or U4187 (N_4187,N_3948,N_3763);
and U4188 (N_4188,N_3776,N_3931);
nor U4189 (N_4189,N_3917,N_3773);
xor U4190 (N_4190,N_3925,N_3869);
or U4191 (N_4191,N_3813,N_3928);
nand U4192 (N_4192,N_3768,N_3998);
xor U4193 (N_4193,N_3934,N_3936);
or U4194 (N_4194,N_3975,N_3768);
and U4195 (N_4195,N_3794,N_3802);
nor U4196 (N_4196,N_3873,N_3833);
nor U4197 (N_4197,N_3806,N_3766);
or U4198 (N_4198,N_3860,N_3956);
nand U4199 (N_4199,N_3789,N_3927);
xnor U4200 (N_4200,N_3777,N_3998);
xnor U4201 (N_4201,N_3914,N_3752);
or U4202 (N_4202,N_3755,N_3831);
xor U4203 (N_4203,N_3911,N_3966);
nand U4204 (N_4204,N_3878,N_3868);
nor U4205 (N_4205,N_3844,N_3981);
or U4206 (N_4206,N_3998,N_3953);
nand U4207 (N_4207,N_3972,N_3865);
xnor U4208 (N_4208,N_3822,N_3757);
nor U4209 (N_4209,N_3929,N_3889);
and U4210 (N_4210,N_3902,N_3823);
xor U4211 (N_4211,N_3793,N_3947);
and U4212 (N_4212,N_3825,N_3856);
or U4213 (N_4213,N_3763,N_3939);
nand U4214 (N_4214,N_3868,N_3866);
xor U4215 (N_4215,N_3818,N_3763);
and U4216 (N_4216,N_3847,N_3874);
xnor U4217 (N_4217,N_3854,N_3819);
xor U4218 (N_4218,N_3963,N_3754);
xnor U4219 (N_4219,N_3769,N_3981);
or U4220 (N_4220,N_3821,N_3877);
or U4221 (N_4221,N_3934,N_3900);
or U4222 (N_4222,N_3876,N_3830);
and U4223 (N_4223,N_3974,N_3825);
and U4224 (N_4224,N_3771,N_3821);
and U4225 (N_4225,N_3840,N_3757);
nor U4226 (N_4226,N_3766,N_3838);
xnor U4227 (N_4227,N_3945,N_3928);
nand U4228 (N_4228,N_3913,N_3968);
or U4229 (N_4229,N_3767,N_3950);
or U4230 (N_4230,N_3889,N_3839);
xnor U4231 (N_4231,N_3991,N_3817);
and U4232 (N_4232,N_3878,N_3879);
nor U4233 (N_4233,N_3971,N_3927);
nor U4234 (N_4234,N_3861,N_3842);
or U4235 (N_4235,N_3820,N_3877);
nand U4236 (N_4236,N_3868,N_3885);
nand U4237 (N_4237,N_3925,N_3983);
nand U4238 (N_4238,N_3966,N_3925);
nor U4239 (N_4239,N_3938,N_3838);
nand U4240 (N_4240,N_3999,N_3871);
or U4241 (N_4241,N_3790,N_3836);
nor U4242 (N_4242,N_3829,N_3884);
nand U4243 (N_4243,N_3867,N_3758);
xnor U4244 (N_4244,N_3983,N_3997);
and U4245 (N_4245,N_3762,N_3935);
xnor U4246 (N_4246,N_3913,N_3870);
nand U4247 (N_4247,N_3952,N_3864);
xnor U4248 (N_4248,N_3847,N_3791);
xnor U4249 (N_4249,N_3798,N_3949);
xor U4250 (N_4250,N_4185,N_4046);
xnor U4251 (N_4251,N_4172,N_4019);
nor U4252 (N_4252,N_4175,N_4101);
and U4253 (N_4253,N_4063,N_4065);
xor U4254 (N_4254,N_4029,N_4064);
and U4255 (N_4255,N_4199,N_4060);
nor U4256 (N_4256,N_4201,N_4118);
nand U4257 (N_4257,N_4051,N_4194);
or U4258 (N_4258,N_4009,N_4216);
xnor U4259 (N_4259,N_4163,N_4197);
nor U4260 (N_4260,N_4139,N_4129);
nand U4261 (N_4261,N_4239,N_4031);
and U4262 (N_4262,N_4195,N_4234);
or U4263 (N_4263,N_4189,N_4224);
and U4264 (N_4264,N_4020,N_4231);
or U4265 (N_4265,N_4081,N_4002);
xnor U4266 (N_4266,N_4115,N_4169);
or U4267 (N_4267,N_4208,N_4240);
or U4268 (N_4268,N_4110,N_4220);
xor U4269 (N_4269,N_4232,N_4067);
nor U4270 (N_4270,N_4157,N_4187);
or U4271 (N_4271,N_4089,N_4132);
xor U4272 (N_4272,N_4047,N_4249);
and U4273 (N_4273,N_4092,N_4087);
or U4274 (N_4274,N_4083,N_4088);
and U4275 (N_4275,N_4230,N_4135);
xor U4276 (N_4276,N_4015,N_4096);
xor U4277 (N_4277,N_4095,N_4026);
xor U4278 (N_4278,N_4117,N_4145);
nor U4279 (N_4279,N_4165,N_4179);
xor U4280 (N_4280,N_4209,N_4138);
and U4281 (N_4281,N_4071,N_4143);
nor U4282 (N_4282,N_4061,N_4114);
xnor U4283 (N_4283,N_4121,N_4207);
xnor U4284 (N_4284,N_4038,N_4164);
nand U4285 (N_4285,N_4133,N_4093);
nand U4286 (N_4286,N_4192,N_4235);
xnor U4287 (N_4287,N_4109,N_4069);
xnor U4288 (N_4288,N_4237,N_4200);
nand U4289 (N_4289,N_4097,N_4106);
and U4290 (N_4290,N_4146,N_4098);
xnor U4291 (N_4291,N_4050,N_4241);
xor U4292 (N_4292,N_4198,N_4018);
and U4293 (N_4293,N_4193,N_4040);
or U4294 (N_4294,N_4105,N_4225);
nor U4295 (N_4295,N_4131,N_4032);
and U4296 (N_4296,N_4127,N_4104);
xnor U4297 (N_4297,N_4119,N_4034);
and U4298 (N_4298,N_4123,N_4148);
and U4299 (N_4299,N_4149,N_4073);
or U4300 (N_4300,N_4217,N_4013);
nor U4301 (N_4301,N_4111,N_4141);
or U4302 (N_4302,N_4022,N_4228);
nor U4303 (N_4303,N_4017,N_4108);
nand U4304 (N_4304,N_4044,N_4025);
xor U4305 (N_4305,N_4007,N_4014);
nor U4306 (N_4306,N_4184,N_4153);
xor U4307 (N_4307,N_4024,N_4159);
and U4308 (N_4308,N_4052,N_4102);
xor U4309 (N_4309,N_4057,N_4113);
xnor U4310 (N_4310,N_4030,N_4103);
nand U4311 (N_4311,N_4245,N_4076);
nor U4312 (N_4312,N_4016,N_4037);
or U4313 (N_4313,N_4176,N_4028);
or U4314 (N_4314,N_4190,N_4130);
xnor U4315 (N_4315,N_4134,N_4191);
and U4316 (N_4316,N_4229,N_4086);
or U4317 (N_4317,N_4116,N_4162);
nor U4318 (N_4318,N_4221,N_4167);
and U4319 (N_4319,N_4154,N_4211);
and U4320 (N_4320,N_4010,N_4171);
or U4321 (N_4321,N_4210,N_4074);
xor U4322 (N_4322,N_4178,N_4120);
and U4323 (N_4323,N_4222,N_4036);
xor U4324 (N_4324,N_4170,N_4203);
xor U4325 (N_4325,N_4227,N_4005);
nor U4326 (N_4326,N_4001,N_4023);
or U4327 (N_4327,N_4219,N_4125);
or U4328 (N_4328,N_4011,N_4054);
nor U4329 (N_4329,N_4147,N_4226);
nor U4330 (N_4330,N_4246,N_4077);
nor U4331 (N_4331,N_4158,N_4248);
or U4332 (N_4332,N_4155,N_4173);
nand U4333 (N_4333,N_4055,N_4218);
and U4334 (N_4334,N_4233,N_4039);
nand U4335 (N_4335,N_4004,N_4186);
nand U4336 (N_4336,N_4181,N_4128);
nand U4337 (N_4337,N_4042,N_4160);
and U4338 (N_4338,N_4150,N_4003);
and U4339 (N_4339,N_4033,N_4021);
and U4340 (N_4340,N_4045,N_4070);
and U4341 (N_4341,N_4080,N_4094);
and U4342 (N_4342,N_4084,N_4124);
or U4343 (N_4343,N_4078,N_4215);
and U4344 (N_4344,N_4056,N_4238);
nor U4345 (N_4345,N_4053,N_4188);
nor U4346 (N_4346,N_4242,N_4223);
nor U4347 (N_4347,N_4059,N_4099);
nand U4348 (N_4348,N_4214,N_4100);
or U4349 (N_4349,N_4043,N_4152);
xnor U4350 (N_4350,N_4072,N_4174);
nand U4351 (N_4351,N_4137,N_4068);
nor U4352 (N_4352,N_4085,N_4107);
nand U4353 (N_4353,N_4041,N_4244);
or U4354 (N_4354,N_4183,N_4062);
and U4355 (N_4355,N_4166,N_4142);
nor U4356 (N_4356,N_4136,N_4202);
and U4357 (N_4357,N_4140,N_4205);
nand U4358 (N_4358,N_4243,N_4161);
and U4359 (N_4359,N_4247,N_4182);
xor U4360 (N_4360,N_4012,N_4212);
nand U4361 (N_4361,N_4049,N_4079);
and U4362 (N_4362,N_4168,N_4122);
xnor U4363 (N_4363,N_4090,N_4177);
and U4364 (N_4364,N_4000,N_4048);
nor U4365 (N_4365,N_4196,N_4058);
and U4366 (N_4366,N_4066,N_4156);
nor U4367 (N_4367,N_4006,N_4091);
nand U4368 (N_4368,N_4236,N_4204);
and U4369 (N_4369,N_4082,N_4027);
nand U4370 (N_4370,N_4213,N_4008);
and U4371 (N_4371,N_4180,N_4112);
or U4372 (N_4372,N_4151,N_4144);
nand U4373 (N_4373,N_4126,N_4206);
nor U4374 (N_4374,N_4075,N_4035);
xor U4375 (N_4375,N_4114,N_4170);
and U4376 (N_4376,N_4015,N_4239);
nor U4377 (N_4377,N_4226,N_4199);
nand U4378 (N_4378,N_4146,N_4142);
xnor U4379 (N_4379,N_4156,N_4177);
xor U4380 (N_4380,N_4090,N_4082);
nor U4381 (N_4381,N_4249,N_4104);
nand U4382 (N_4382,N_4185,N_4108);
nor U4383 (N_4383,N_4241,N_4055);
xor U4384 (N_4384,N_4062,N_4090);
nand U4385 (N_4385,N_4048,N_4235);
nor U4386 (N_4386,N_4249,N_4019);
or U4387 (N_4387,N_4143,N_4036);
or U4388 (N_4388,N_4249,N_4151);
nor U4389 (N_4389,N_4096,N_4188);
and U4390 (N_4390,N_4122,N_4215);
and U4391 (N_4391,N_4096,N_4186);
xor U4392 (N_4392,N_4222,N_4216);
nor U4393 (N_4393,N_4226,N_4071);
or U4394 (N_4394,N_4224,N_4167);
nor U4395 (N_4395,N_4213,N_4039);
and U4396 (N_4396,N_4083,N_4239);
nor U4397 (N_4397,N_4205,N_4167);
or U4398 (N_4398,N_4036,N_4203);
nor U4399 (N_4399,N_4203,N_4222);
xor U4400 (N_4400,N_4009,N_4000);
and U4401 (N_4401,N_4071,N_4037);
xor U4402 (N_4402,N_4126,N_4044);
nand U4403 (N_4403,N_4144,N_4227);
nand U4404 (N_4404,N_4055,N_4163);
nand U4405 (N_4405,N_4070,N_4225);
nor U4406 (N_4406,N_4105,N_4064);
xor U4407 (N_4407,N_4104,N_4170);
xnor U4408 (N_4408,N_4172,N_4157);
nand U4409 (N_4409,N_4036,N_4054);
or U4410 (N_4410,N_4197,N_4001);
or U4411 (N_4411,N_4013,N_4073);
nor U4412 (N_4412,N_4012,N_4213);
xor U4413 (N_4413,N_4043,N_4022);
nor U4414 (N_4414,N_4061,N_4159);
or U4415 (N_4415,N_4005,N_4168);
nand U4416 (N_4416,N_4087,N_4177);
or U4417 (N_4417,N_4045,N_4176);
and U4418 (N_4418,N_4016,N_4070);
or U4419 (N_4419,N_4152,N_4052);
xnor U4420 (N_4420,N_4076,N_4080);
or U4421 (N_4421,N_4187,N_4245);
or U4422 (N_4422,N_4122,N_4220);
nand U4423 (N_4423,N_4204,N_4213);
nand U4424 (N_4424,N_4150,N_4172);
xnor U4425 (N_4425,N_4138,N_4204);
nand U4426 (N_4426,N_4129,N_4180);
or U4427 (N_4427,N_4186,N_4231);
or U4428 (N_4428,N_4026,N_4098);
nand U4429 (N_4429,N_4124,N_4106);
nand U4430 (N_4430,N_4116,N_4055);
xnor U4431 (N_4431,N_4224,N_4198);
xnor U4432 (N_4432,N_4186,N_4052);
nor U4433 (N_4433,N_4078,N_4172);
nor U4434 (N_4434,N_4063,N_4001);
and U4435 (N_4435,N_4151,N_4235);
or U4436 (N_4436,N_4181,N_4217);
nor U4437 (N_4437,N_4193,N_4097);
or U4438 (N_4438,N_4176,N_4181);
and U4439 (N_4439,N_4021,N_4113);
or U4440 (N_4440,N_4128,N_4082);
nand U4441 (N_4441,N_4133,N_4088);
nor U4442 (N_4442,N_4179,N_4145);
nand U4443 (N_4443,N_4079,N_4076);
and U4444 (N_4444,N_4051,N_4015);
xor U4445 (N_4445,N_4099,N_4094);
nand U4446 (N_4446,N_4120,N_4180);
and U4447 (N_4447,N_4236,N_4122);
or U4448 (N_4448,N_4166,N_4165);
nor U4449 (N_4449,N_4157,N_4160);
nor U4450 (N_4450,N_4011,N_4038);
nor U4451 (N_4451,N_4197,N_4101);
and U4452 (N_4452,N_4134,N_4128);
nor U4453 (N_4453,N_4015,N_4236);
or U4454 (N_4454,N_4105,N_4130);
nand U4455 (N_4455,N_4045,N_4034);
xor U4456 (N_4456,N_4046,N_4189);
and U4457 (N_4457,N_4098,N_4010);
nor U4458 (N_4458,N_4034,N_4038);
and U4459 (N_4459,N_4158,N_4231);
or U4460 (N_4460,N_4249,N_4057);
or U4461 (N_4461,N_4214,N_4213);
nor U4462 (N_4462,N_4070,N_4048);
and U4463 (N_4463,N_4210,N_4118);
and U4464 (N_4464,N_4223,N_4001);
nor U4465 (N_4465,N_4088,N_4192);
nand U4466 (N_4466,N_4222,N_4052);
and U4467 (N_4467,N_4080,N_4083);
nand U4468 (N_4468,N_4247,N_4243);
nand U4469 (N_4469,N_4118,N_4054);
or U4470 (N_4470,N_4009,N_4037);
and U4471 (N_4471,N_4232,N_4109);
xor U4472 (N_4472,N_4141,N_4034);
nand U4473 (N_4473,N_4022,N_4007);
xor U4474 (N_4474,N_4038,N_4081);
nand U4475 (N_4475,N_4174,N_4207);
nor U4476 (N_4476,N_4023,N_4142);
xnor U4477 (N_4477,N_4047,N_4207);
nor U4478 (N_4478,N_4039,N_4138);
or U4479 (N_4479,N_4015,N_4016);
xnor U4480 (N_4480,N_4042,N_4219);
nor U4481 (N_4481,N_4078,N_4079);
nor U4482 (N_4482,N_4043,N_4075);
nand U4483 (N_4483,N_4248,N_4055);
nor U4484 (N_4484,N_4136,N_4013);
nand U4485 (N_4485,N_4051,N_4088);
and U4486 (N_4486,N_4205,N_4029);
and U4487 (N_4487,N_4039,N_4095);
or U4488 (N_4488,N_4180,N_4140);
and U4489 (N_4489,N_4036,N_4020);
xnor U4490 (N_4490,N_4168,N_4081);
and U4491 (N_4491,N_4208,N_4207);
nand U4492 (N_4492,N_4034,N_4143);
nor U4493 (N_4493,N_4102,N_4083);
xor U4494 (N_4494,N_4008,N_4232);
and U4495 (N_4495,N_4093,N_4149);
and U4496 (N_4496,N_4125,N_4156);
nand U4497 (N_4497,N_4114,N_4194);
xnor U4498 (N_4498,N_4086,N_4235);
and U4499 (N_4499,N_4178,N_4034);
and U4500 (N_4500,N_4483,N_4397);
or U4501 (N_4501,N_4305,N_4330);
nand U4502 (N_4502,N_4302,N_4316);
or U4503 (N_4503,N_4400,N_4338);
and U4504 (N_4504,N_4441,N_4474);
nand U4505 (N_4505,N_4287,N_4383);
and U4506 (N_4506,N_4456,N_4303);
nor U4507 (N_4507,N_4380,N_4429);
nor U4508 (N_4508,N_4356,N_4258);
xnor U4509 (N_4509,N_4279,N_4496);
nand U4510 (N_4510,N_4486,N_4365);
and U4511 (N_4511,N_4490,N_4373);
xor U4512 (N_4512,N_4253,N_4299);
xor U4513 (N_4513,N_4321,N_4339);
or U4514 (N_4514,N_4276,N_4291);
xnor U4515 (N_4515,N_4307,N_4317);
xnor U4516 (N_4516,N_4460,N_4322);
and U4517 (N_4517,N_4323,N_4327);
and U4518 (N_4518,N_4359,N_4379);
and U4519 (N_4519,N_4271,N_4407);
xor U4520 (N_4520,N_4479,N_4416);
nand U4521 (N_4521,N_4455,N_4284);
nand U4522 (N_4522,N_4403,N_4375);
and U4523 (N_4523,N_4275,N_4300);
nor U4524 (N_4524,N_4434,N_4467);
nand U4525 (N_4525,N_4289,N_4354);
or U4526 (N_4526,N_4454,N_4470);
and U4527 (N_4527,N_4415,N_4335);
nor U4528 (N_4528,N_4462,N_4360);
nor U4529 (N_4529,N_4385,N_4402);
and U4530 (N_4530,N_4315,N_4469);
and U4531 (N_4531,N_4278,N_4311);
xor U4532 (N_4532,N_4286,N_4256);
nor U4533 (N_4533,N_4353,N_4346);
xor U4534 (N_4534,N_4386,N_4266);
xnor U4535 (N_4535,N_4304,N_4450);
nor U4536 (N_4536,N_4267,N_4314);
nand U4537 (N_4537,N_4263,N_4370);
nand U4538 (N_4538,N_4398,N_4423);
or U4539 (N_4539,N_4259,N_4369);
nand U4540 (N_4540,N_4274,N_4343);
xor U4541 (N_4541,N_4439,N_4306);
nand U4542 (N_4542,N_4412,N_4301);
or U4543 (N_4543,N_4366,N_4282);
xor U4544 (N_4544,N_4324,N_4340);
or U4545 (N_4545,N_4485,N_4308);
or U4546 (N_4546,N_4355,N_4482);
xor U4547 (N_4547,N_4499,N_4288);
and U4548 (N_4548,N_4442,N_4494);
nand U4549 (N_4549,N_4408,N_4443);
or U4550 (N_4550,N_4336,N_4491);
or U4551 (N_4551,N_4477,N_4458);
xor U4552 (N_4552,N_4478,N_4390);
xor U4553 (N_4553,N_4328,N_4362);
or U4554 (N_4554,N_4350,N_4440);
nor U4555 (N_4555,N_4252,N_4413);
and U4556 (N_4556,N_4420,N_4272);
nand U4557 (N_4557,N_4424,N_4293);
or U4558 (N_4558,N_4466,N_4384);
nand U4559 (N_4559,N_4295,N_4254);
nand U4560 (N_4560,N_4364,N_4472);
and U4561 (N_4561,N_4399,N_4351);
nand U4562 (N_4562,N_4417,N_4461);
nand U4563 (N_4563,N_4435,N_4358);
nand U4564 (N_4564,N_4325,N_4463);
nor U4565 (N_4565,N_4487,N_4476);
and U4566 (N_4566,N_4337,N_4387);
nor U4567 (N_4567,N_4404,N_4382);
and U4568 (N_4568,N_4427,N_4392);
nand U4569 (N_4569,N_4492,N_4372);
nand U4570 (N_4570,N_4395,N_4331);
nor U4571 (N_4571,N_4446,N_4270);
xor U4572 (N_4572,N_4347,N_4459);
xor U4573 (N_4573,N_4401,N_4457);
nor U4574 (N_4574,N_4444,N_4333);
xnor U4575 (N_4575,N_4394,N_4448);
xnor U4576 (N_4576,N_4409,N_4464);
xor U4577 (N_4577,N_4332,N_4363);
nand U4578 (N_4578,N_4264,N_4273);
nand U4579 (N_4579,N_4422,N_4312);
or U4580 (N_4580,N_4309,N_4344);
nand U4581 (N_4581,N_4349,N_4447);
and U4582 (N_4582,N_4433,N_4378);
xor U4583 (N_4583,N_4481,N_4342);
nor U4584 (N_4584,N_4292,N_4453);
and U4585 (N_4585,N_4357,N_4445);
and U4586 (N_4586,N_4431,N_4393);
xnor U4587 (N_4587,N_4451,N_4320);
or U4588 (N_4588,N_4277,N_4341);
or U4589 (N_4589,N_4497,N_4352);
and U4590 (N_4590,N_4260,N_4449);
and U4591 (N_4591,N_4294,N_4495);
xor U4592 (N_4592,N_4438,N_4334);
nor U4593 (N_4593,N_4419,N_4269);
or U4594 (N_4594,N_4488,N_4255);
or U4595 (N_4595,N_4452,N_4391);
nor U4596 (N_4596,N_4489,N_4329);
nand U4597 (N_4597,N_4414,N_4290);
nand U4598 (N_4598,N_4406,N_4426);
nor U4599 (N_4599,N_4265,N_4436);
nand U4600 (N_4600,N_4425,N_4471);
xnor U4601 (N_4601,N_4468,N_4310);
and U4602 (N_4602,N_4367,N_4410);
xnor U4603 (N_4603,N_4377,N_4418);
xnor U4604 (N_4604,N_4251,N_4493);
and U4605 (N_4605,N_4250,N_4318);
nand U4606 (N_4606,N_4428,N_4368);
or U4607 (N_4607,N_4296,N_4381);
or U4608 (N_4608,N_4345,N_4297);
or U4609 (N_4609,N_4298,N_4374);
and U4610 (N_4610,N_4432,N_4326);
nor U4611 (N_4611,N_4376,N_4396);
and U4612 (N_4612,N_4484,N_4421);
nor U4613 (N_4613,N_4348,N_4480);
xnor U4614 (N_4614,N_4411,N_4389);
xor U4615 (N_4615,N_4257,N_4430);
xor U4616 (N_4616,N_4313,N_4283);
nor U4617 (N_4617,N_4405,N_4465);
or U4618 (N_4618,N_4281,N_4498);
xnor U4619 (N_4619,N_4361,N_4262);
or U4620 (N_4620,N_4473,N_4280);
nor U4621 (N_4621,N_4268,N_4261);
or U4622 (N_4622,N_4475,N_4285);
or U4623 (N_4623,N_4388,N_4437);
or U4624 (N_4624,N_4371,N_4319);
nor U4625 (N_4625,N_4479,N_4443);
nand U4626 (N_4626,N_4497,N_4407);
and U4627 (N_4627,N_4473,N_4448);
xor U4628 (N_4628,N_4308,N_4323);
xor U4629 (N_4629,N_4351,N_4279);
nor U4630 (N_4630,N_4407,N_4428);
nand U4631 (N_4631,N_4360,N_4415);
and U4632 (N_4632,N_4422,N_4387);
nand U4633 (N_4633,N_4427,N_4487);
or U4634 (N_4634,N_4428,N_4482);
nor U4635 (N_4635,N_4293,N_4473);
nor U4636 (N_4636,N_4371,N_4464);
nand U4637 (N_4637,N_4495,N_4262);
or U4638 (N_4638,N_4258,N_4336);
nand U4639 (N_4639,N_4355,N_4464);
nand U4640 (N_4640,N_4256,N_4484);
nor U4641 (N_4641,N_4471,N_4466);
nor U4642 (N_4642,N_4290,N_4318);
nand U4643 (N_4643,N_4315,N_4253);
xor U4644 (N_4644,N_4291,N_4325);
nand U4645 (N_4645,N_4451,N_4331);
or U4646 (N_4646,N_4475,N_4427);
xnor U4647 (N_4647,N_4455,N_4447);
and U4648 (N_4648,N_4400,N_4468);
nor U4649 (N_4649,N_4281,N_4465);
and U4650 (N_4650,N_4386,N_4490);
and U4651 (N_4651,N_4473,N_4356);
and U4652 (N_4652,N_4345,N_4403);
xnor U4653 (N_4653,N_4467,N_4363);
or U4654 (N_4654,N_4350,N_4474);
nand U4655 (N_4655,N_4383,N_4498);
nor U4656 (N_4656,N_4469,N_4368);
nor U4657 (N_4657,N_4277,N_4458);
nand U4658 (N_4658,N_4403,N_4274);
and U4659 (N_4659,N_4299,N_4303);
nand U4660 (N_4660,N_4296,N_4407);
xnor U4661 (N_4661,N_4322,N_4482);
nand U4662 (N_4662,N_4330,N_4444);
or U4663 (N_4663,N_4268,N_4424);
nor U4664 (N_4664,N_4366,N_4435);
nand U4665 (N_4665,N_4338,N_4349);
nor U4666 (N_4666,N_4345,N_4333);
nand U4667 (N_4667,N_4334,N_4471);
and U4668 (N_4668,N_4408,N_4316);
xor U4669 (N_4669,N_4388,N_4382);
or U4670 (N_4670,N_4397,N_4314);
xnor U4671 (N_4671,N_4422,N_4339);
and U4672 (N_4672,N_4475,N_4400);
nand U4673 (N_4673,N_4280,N_4315);
and U4674 (N_4674,N_4382,N_4286);
or U4675 (N_4675,N_4490,N_4378);
and U4676 (N_4676,N_4490,N_4420);
or U4677 (N_4677,N_4393,N_4432);
nand U4678 (N_4678,N_4293,N_4264);
xnor U4679 (N_4679,N_4451,N_4371);
nor U4680 (N_4680,N_4415,N_4268);
and U4681 (N_4681,N_4285,N_4399);
or U4682 (N_4682,N_4456,N_4419);
nor U4683 (N_4683,N_4349,N_4401);
or U4684 (N_4684,N_4356,N_4470);
nor U4685 (N_4685,N_4378,N_4318);
and U4686 (N_4686,N_4399,N_4467);
or U4687 (N_4687,N_4433,N_4383);
xor U4688 (N_4688,N_4330,N_4285);
or U4689 (N_4689,N_4365,N_4324);
nor U4690 (N_4690,N_4434,N_4341);
nand U4691 (N_4691,N_4358,N_4479);
and U4692 (N_4692,N_4337,N_4310);
or U4693 (N_4693,N_4471,N_4373);
or U4694 (N_4694,N_4279,N_4407);
nand U4695 (N_4695,N_4302,N_4377);
nand U4696 (N_4696,N_4268,N_4353);
or U4697 (N_4697,N_4305,N_4297);
or U4698 (N_4698,N_4489,N_4478);
nor U4699 (N_4699,N_4408,N_4281);
xnor U4700 (N_4700,N_4365,N_4295);
or U4701 (N_4701,N_4375,N_4486);
xor U4702 (N_4702,N_4293,N_4253);
nand U4703 (N_4703,N_4277,N_4313);
xor U4704 (N_4704,N_4311,N_4423);
nor U4705 (N_4705,N_4258,N_4370);
xnor U4706 (N_4706,N_4274,N_4456);
and U4707 (N_4707,N_4338,N_4335);
or U4708 (N_4708,N_4373,N_4429);
nor U4709 (N_4709,N_4316,N_4447);
xor U4710 (N_4710,N_4360,N_4305);
xnor U4711 (N_4711,N_4471,N_4310);
xor U4712 (N_4712,N_4310,N_4371);
and U4713 (N_4713,N_4436,N_4455);
xor U4714 (N_4714,N_4494,N_4287);
and U4715 (N_4715,N_4322,N_4378);
and U4716 (N_4716,N_4356,N_4330);
and U4717 (N_4717,N_4421,N_4420);
nand U4718 (N_4718,N_4254,N_4296);
xor U4719 (N_4719,N_4404,N_4417);
or U4720 (N_4720,N_4425,N_4261);
xnor U4721 (N_4721,N_4461,N_4429);
nand U4722 (N_4722,N_4290,N_4374);
nand U4723 (N_4723,N_4396,N_4344);
nand U4724 (N_4724,N_4461,N_4289);
or U4725 (N_4725,N_4253,N_4440);
or U4726 (N_4726,N_4480,N_4284);
or U4727 (N_4727,N_4342,N_4271);
xnor U4728 (N_4728,N_4403,N_4395);
nand U4729 (N_4729,N_4355,N_4292);
nor U4730 (N_4730,N_4397,N_4496);
nor U4731 (N_4731,N_4475,N_4394);
or U4732 (N_4732,N_4404,N_4321);
nor U4733 (N_4733,N_4267,N_4391);
nand U4734 (N_4734,N_4292,N_4255);
nor U4735 (N_4735,N_4443,N_4378);
nand U4736 (N_4736,N_4253,N_4270);
nor U4737 (N_4737,N_4302,N_4361);
nand U4738 (N_4738,N_4286,N_4491);
nand U4739 (N_4739,N_4429,N_4281);
nor U4740 (N_4740,N_4485,N_4439);
or U4741 (N_4741,N_4365,N_4316);
xor U4742 (N_4742,N_4360,N_4483);
or U4743 (N_4743,N_4340,N_4298);
nand U4744 (N_4744,N_4382,N_4480);
nand U4745 (N_4745,N_4456,N_4354);
or U4746 (N_4746,N_4353,N_4422);
xnor U4747 (N_4747,N_4303,N_4489);
and U4748 (N_4748,N_4358,N_4398);
nor U4749 (N_4749,N_4253,N_4493);
or U4750 (N_4750,N_4545,N_4537);
xnor U4751 (N_4751,N_4523,N_4525);
xor U4752 (N_4752,N_4544,N_4747);
or U4753 (N_4753,N_4699,N_4739);
or U4754 (N_4754,N_4737,N_4532);
nor U4755 (N_4755,N_4654,N_4612);
nand U4756 (N_4756,N_4711,N_4517);
or U4757 (N_4757,N_4571,N_4568);
nor U4758 (N_4758,N_4666,N_4633);
xnor U4759 (N_4759,N_4604,N_4681);
nor U4760 (N_4760,N_4621,N_4719);
xnor U4761 (N_4761,N_4581,N_4565);
xor U4762 (N_4762,N_4520,N_4600);
and U4763 (N_4763,N_4589,N_4697);
nand U4764 (N_4764,N_4569,N_4730);
and U4765 (N_4765,N_4631,N_4695);
xnor U4766 (N_4766,N_4658,N_4587);
nand U4767 (N_4767,N_4614,N_4682);
nor U4768 (N_4768,N_4701,N_4536);
or U4769 (N_4769,N_4669,N_4686);
nand U4770 (N_4770,N_4570,N_4659);
or U4771 (N_4771,N_4744,N_4736);
nand U4772 (N_4772,N_4519,N_4579);
or U4773 (N_4773,N_4512,N_4567);
and U4774 (N_4774,N_4628,N_4749);
and U4775 (N_4775,N_4732,N_4691);
nand U4776 (N_4776,N_4647,N_4574);
and U4777 (N_4777,N_4746,N_4690);
xnor U4778 (N_4778,N_4521,N_4615);
and U4779 (N_4779,N_4726,N_4649);
or U4780 (N_4780,N_4653,N_4529);
or U4781 (N_4781,N_4616,N_4680);
nor U4782 (N_4782,N_4675,N_4602);
and U4783 (N_4783,N_4625,N_4601);
and U4784 (N_4784,N_4588,N_4668);
nor U4785 (N_4785,N_4578,N_4594);
nand U4786 (N_4786,N_4677,N_4640);
and U4787 (N_4787,N_4643,N_4582);
nand U4788 (N_4788,N_4700,N_4651);
and U4789 (N_4789,N_4524,N_4598);
nor U4790 (N_4790,N_4539,N_4636);
nand U4791 (N_4791,N_4703,N_4549);
xnor U4792 (N_4792,N_4663,N_4577);
or U4793 (N_4793,N_4721,N_4678);
nand U4794 (N_4794,N_4531,N_4500);
nor U4795 (N_4795,N_4627,N_4731);
nand U4796 (N_4796,N_4620,N_4717);
nand U4797 (N_4797,N_4554,N_4684);
and U4798 (N_4798,N_4683,N_4644);
xnor U4799 (N_4799,N_4559,N_4667);
and U4800 (N_4800,N_4630,N_4502);
nor U4801 (N_4801,N_4557,N_4650);
or U4802 (N_4802,N_4605,N_4655);
or U4803 (N_4803,N_4685,N_4505);
nor U4804 (N_4804,N_4706,N_4560);
or U4805 (N_4805,N_4634,N_4573);
or U4806 (N_4806,N_4696,N_4635);
or U4807 (N_4807,N_4617,N_4725);
or U4808 (N_4808,N_4507,N_4506);
nor U4809 (N_4809,N_4641,N_4508);
and U4810 (N_4810,N_4530,N_4714);
nand U4811 (N_4811,N_4606,N_4608);
or U4812 (N_4812,N_4564,N_4660);
and U4813 (N_4813,N_4548,N_4671);
nand U4814 (N_4814,N_4694,N_4503);
nor U4815 (N_4815,N_4563,N_4556);
or U4816 (N_4816,N_4592,N_4709);
and U4817 (N_4817,N_4527,N_4713);
nand U4818 (N_4818,N_4585,N_4642);
and U4819 (N_4819,N_4638,N_4715);
and U4820 (N_4820,N_4716,N_4613);
or U4821 (N_4821,N_4551,N_4522);
nand U4822 (N_4822,N_4722,N_4727);
and U4823 (N_4823,N_4610,N_4619);
nor U4824 (N_4824,N_4637,N_4710);
or U4825 (N_4825,N_4692,N_4679);
or U4826 (N_4826,N_4618,N_4657);
or U4827 (N_4827,N_4504,N_4550);
or U4828 (N_4828,N_4639,N_4704);
xor U4829 (N_4829,N_4552,N_4586);
xor U4830 (N_4830,N_4595,N_4541);
or U4831 (N_4831,N_4665,N_4661);
and U4832 (N_4832,N_4599,N_4702);
nor U4833 (N_4833,N_4543,N_4729);
nor U4834 (N_4834,N_4741,N_4624);
nand U4835 (N_4835,N_4590,N_4623);
xnor U4836 (N_4836,N_4591,N_4670);
nor U4837 (N_4837,N_4745,N_4566);
or U4838 (N_4838,N_4648,N_4705);
nand U4839 (N_4839,N_4738,N_4733);
and U4840 (N_4840,N_4707,N_4611);
or U4841 (N_4841,N_4740,N_4513);
or U4842 (N_4842,N_4646,N_4580);
nand U4843 (N_4843,N_4672,N_4533);
nor U4844 (N_4844,N_4673,N_4547);
nor U4845 (N_4845,N_4526,N_4742);
nand U4846 (N_4846,N_4662,N_4652);
nand U4847 (N_4847,N_4597,N_4510);
nand U4848 (N_4848,N_4555,N_4688);
nand U4849 (N_4849,N_4734,N_4632);
nand U4850 (N_4850,N_4708,N_4553);
and U4851 (N_4851,N_4622,N_4596);
xor U4852 (N_4852,N_4584,N_4674);
or U4853 (N_4853,N_4576,N_4514);
and U4854 (N_4854,N_4515,N_4693);
or U4855 (N_4855,N_4575,N_4712);
xor U4856 (N_4856,N_4593,N_4562);
or U4857 (N_4857,N_4542,N_4609);
xnor U4858 (N_4858,N_4528,N_4720);
or U4859 (N_4859,N_4511,N_4735);
xnor U4860 (N_4860,N_4534,N_4558);
nor U4861 (N_4861,N_4629,N_4518);
xor U4862 (N_4862,N_4509,N_4656);
or U4863 (N_4863,N_4698,N_4546);
and U4864 (N_4864,N_4626,N_4748);
xnor U4865 (N_4865,N_4724,N_4561);
xor U4866 (N_4866,N_4689,N_4501);
nand U4867 (N_4867,N_4728,N_4516);
nor U4868 (N_4868,N_4743,N_4538);
nor U4869 (N_4869,N_4723,N_4540);
xor U4870 (N_4870,N_4583,N_4645);
or U4871 (N_4871,N_4687,N_4676);
or U4872 (N_4872,N_4572,N_4607);
or U4873 (N_4873,N_4664,N_4603);
nand U4874 (N_4874,N_4535,N_4718);
xor U4875 (N_4875,N_4738,N_4577);
xor U4876 (N_4876,N_4620,N_4685);
xor U4877 (N_4877,N_4651,N_4689);
and U4878 (N_4878,N_4684,N_4658);
nand U4879 (N_4879,N_4633,N_4722);
nor U4880 (N_4880,N_4514,N_4550);
and U4881 (N_4881,N_4702,N_4678);
xor U4882 (N_4882,N_4682,N_4749);
or U4883 (N_4883,N_4660,N_4507);
nor U4884 (N_4884,N_4620,N_4548);
or U4885 (N_4885,N_4717,N_4733);
nand U4886 (N_4886,N_4629,N_4638);
or U4887 (N_4887,N_4652,N_4620);
or U4888 (N_4888,N_4587,N_4727);
nand U4889 (N_4889,N_4592,N_4575);
nand U4890 (N_4890,N_4582,N_4501);
and U4891 (N_4891,N_4503,N_4664);
and U4892 (N_4892,N_4706,N_4531);
nor U4893 (N_4893,N_4677,N_4671);
xor U4894 (N_4894,N_4614,N_4545);
nand U4895 (N_4895,N_4673,N_4711);
and U4896 (N_4896,N_4664,N_4629);
nor U4897 (N_4897,N_4699,N_4582);
nand U4898 (N_4898,N_4646,N_4711);
or U4899 (N_4899,N_4591,N_4630);
or U4900 (N_4900,N_4693,N_4609);
nor U4901 (N_4901,N_4722,N_4698);
or U4902 (N_4902,N_4548,N_4690);
xor U4903 (N_4903,N_4618,N_4692);
nor U4904 (N_4904,N_4749,N_4655);
xnor U4905 (N_4905,N_4597,N_4613);
and U4906 (N_4906,N_4748,N_4525);
and U4907 (N_4907,N_4587,N_4693);
xor U4908 (N_4908,N_4588,N_4550);
and U4909 (N_4909,N_4591,N_4502);
xnor U4910 (N_4910,N_4630,N_4660);
or U4911 (N_4911,N_4712,N_4651);
xor U4912 (N_4912,N_4571,N_4508);
or U4913 (N_4913,N_4681,N_4533);
nand U4914 (N_4914,N_4504,N_4699);
and U4915 (N_4915,N_4556,N_4673);
or U4916 (N_4916,N_4664,N_4607);
and U4917 (N_4917,N_4729,N_4645);
and U4918 (N_4918,N_4666,N_4651);
and U4919 (N_4919,N_4718,N_4707);
nor U4920 (N_4920,N_4601,N_4623);
and U4921 (N_4921,N_4602,N_4705);
xnor U4922 (N_4922,N_4531,N_4574);
nor U4923 (N_4923,N_4634,N_4584);
nor U4924 (N_4924,N_4676,N_4680);
nor U4925 (N_4925,N_4642,N_4714);
nor U4926 (N_4926,N_4538,N_4568);
and U4927 (N_4927,N_4514,N_4635);
nor U4928 (N_4928,N_4708,N_4734);
nand U4929 (N_4929,N_4614,N_4559);
or U4930 (N_4930,N_4565,N_4553);
nand U4931 (N_4931,N_4571,N_4611);
or U4932 (N_4932,N_4728,N_4708);
and U4933 (N_4933,N_4629,N_4721);
xnor U4934 (N_4934,N_4694,N_4691);
xor U4935 (N_4935,N_4573,N_4744);
nor U4936 (N_4936,N_4571,N_4553);
and U4937 (N_4937,N_4674,N_4582);
nor U4938 (N_4938,N_4707,N_4658);
nand U4939 (N_4939,N_4623,N_4616);
nand U4940 (N_4940,N_4632,N_4732);
xnor U4941 (N_4941,N_4625,N_4670);
nor U4942 (N_4942,N_4540,N_4582);
nor U4943 (N_4943,N_4645,N_4559);
and U4944 (N_4944,N_4574,N_4567);
nor U4945 (N_4945,N_4616,N_4556);
nor U4946 (N_4946,N_4727,N_4719);
or U4947 (N_4947,N_4557,N_4659);
nor U4948 (N_4948,N_4605,N_4628);
or U4949 (N_4949,N_4677,N_4735);
xnor U4950 (N_4950,N_4613,N_4696);
or U4951 (N_4951,N_4684,N_4641);
nand U4952 (N_4952,N_4595,N_4514);
xnor U4953 (N_4953,N_4558,N_4736);
nand U4954 (N_4954,N_4610,N_4682);
nand U4955 (N_4955,N_4525,N_4611);
xnor U4956 (N_4956,N_4743,N_4745);
xnor U4957 (N_4957,N_4582,N_4655);
and U4958 (N_4958,N_4534,N_4500);
or U4959 (N_4959,N_4659,N_4634);
and U4960 (N_4960,N_4621,N_4629);
and U4961 (N_4961,N_4592,N_4515);
nand U4962 (N_4962,N_4652,N_4732);
nand U4963 (N_4963,N_4591,N_4507);
nor U4964 (N_4964,N_4527,N_4711);
xor U4965 (N_4965,N_4520,N_4586);
or U4966 (N_4966,N_4596,N_4711);
nor U4967 (N_4967,N_4658,N_4669);
nor U4968 (N_4968,N_4709,N_4729);
nand U4969 (N_4969,N_4619,N_4504);
or U4970 (N_4970,N_4611,N_4568);
and U4971 (N_4971,N_4534,N_4637);
nor U4972 (N_4972,N_4623,N_4724);
nand U4973 (N_4973,N_4569,N_4740);
or U4974 (N_4974,N_4539,N_4717);
nor U4975 (N_4975,N_4567,N_4681);
xnor U4976 (N_4976,N_4749,N_4677);
xor U4977 (N_4977,N_4701,N_4741);
or U4978 (N_4978,N_4675,N_4706);
or U4979 (N_4979,N_4681,N_4693);
xor U4980 (N_4980,N_4665,N_4690);
nand U4981 (N_4981,N_4689,N_4724);
nor U4982 (N_4982,N_4585,N_4666);
xnor U4983 (N_4983,N_4664,N_4702);
nor U4984 (N_4984,N_4720,N_4518);
and U4985 (N_4985,N_4595,N_4603);
and U4986 (N_4986,N_4586,N_4533);
and U4987 (N_4987,N_4507,N_4543);
or U4988 (N_4988,N_4690,N_4677);
and U4989 (N_4989,N_4649,N_4535);
xnor U4990 (N_4990,N_4607,N_4548);
and U4991 (N_4991,N_4664,N_4517);
or U4992 (N_4992,N_4546,N_4642);
or U4993 (N_4993,N_4570,N_4728);
xor U4994 (N_4994,N_4632,N_4717);
nand U4995 (N_4995,N_4746,N_4644);
nand U4996 (N_4996,N_4636,N_4725);
and U4997 (N_4997,N_4561,N_4594);
nand U4998 (N_4998,N_4510,N_4504);
nor U4999 (N_4999,N_4559,N_4656);
and U5000 (N_5000,N_4950,N_4990);
nor U5001 (N_5001,N_4857,N_4947);
or U5002 (N_5002,N_4877,N_4953);
or U5003 (N_5003,N_4822,N_4848);
and U5004 (N_5004,N_4915,N_4799);
or U5005 (N_5005,N_4780,N_4881);
nand U5006 (N_5006,N_4942,N_4756);
and U5007 (N_5007,N_4791,N_4826);
nand U5008 (N_5008,N_4927,N_4931);
nor U5009 (N_5009,N_4824,N_4963);
nor U5010 (N_5010,N_4911,N_4803);
nand U5011 (N_5011,N_4818,N_4933);
and U5012 (N_5012,N_4750,N_4984);
and U5013 (N_5013,N_4979,N_4789);
or U5014 (N_5014,N_4825,N_4980);
or U5015 (N_5015,N_4934,N_4919);
and U5016 (N_5016,N_4775,N_4971);
and U5017 (N_5017,N_4921,N_4782);
xor U5018 (N_5018,N_4974,N_4955);
and U5019 (N_5019,N_4809,N_4916);
nand U5020 (N_5020,N_4752,N_4753);
or U5021 (N_5021,N_4948,N_4998);
nand U5022 (N_5022,N_4935,N_4802);
xor U5023 (N_5023,N_4972,N_4843);
or U5024 (N_5024,N_4801,N_4983);
or U5025 (N_5025,N_4944,N_4964);
or U5026 (N_5026,N_4829,N_4781);
xor U5027 (N_5027,N_4783,N_4952);
nand U5028 (N_5028,N_4771,N_4913);
nand U5029 (N_5029,N_4899,N_4855);
nor U5030 (N_5030,N_4999,N_4924);
and U5031 (N_5031,N_4943,N_4859);
nor U5032 (N_5032,N_4914,N_4954);
nand U5033 (N_5033,N_4978,N_4922);
and U5034 (N_5034,N_4897,N_4965);
or U5035 (N_5035,N_4985,N_4865);
xnor U5036 (N_5036,N_4957,N_4808);
xor U5037 (N_5037,N_4800,N_4806);
nor U5038 (N_5038,N_4977,N_4768);
and U5039 (N_5039,N_4997,N_4937);
nor U5040 (N_5040,N_4787,N_4844);
and U5041 (N_5041,N_4784,N_4797);
or U5042 (N_5042,N_4755,N_4982);
nor U5043 (N_5043,N_4760,N_4839);
nor U5044 (N_5044,N_4941,N_4907);
nand U5045 (N_5045,N_4976,N_4830);
and U5046 (N_5046,N_4866,N_4932);
nand U5047 (N_5047,N_4975,N_4905);
nor U5048 (N_5048,N_4902,N_4879);
and U5049 (N_5049,N_4908,N_4923);
and U5050 (N_5050,N_4906,N_4946);
and U5051 (N_5051,N_4793,N_4969);
or U5052 (N_5052,N_4772,N_4838);
nand U5053 (N_5053,N_4798,N_4956);
or U5054 (N_5054,N_4811,N_4821);
and U5055 (N_5055,N_4837,N_4917);
nand U5056 (N_5056,N_4867,N_4961);
and U5057 (N_5057,N_4892,N_4765);
and U5058 (N_5058,N_4850,N_4873);
xor U5059 (N_5059,N_4926,N_4849);
and U5060 (N_5060,N_4847,N_4841);
and U5061 (N_5061,N_4757,N_4883);
nand U5062 (N_5062,N_4819,N_4846);
xnor U5063 (N_5063,N_4949,N_4898);
or U5064 (N_5064,N_4903,N_4761);
nand U5065 (N_5065,N_4938,N_4823);
xnor U5066 (N_5066,N_4989,N_4900);
or U5067 (N_5067,N_4889,N_4875);
nand U5068 (N_5068,N_4835,N_4868);
and U5069 (N_5069,N_4777,N_4778);
nor U5070 (N_5070,N_4754,N_4786);
or U5071 (N_5071,N_4992,N_4884);
or U5072 (N_5072,N_4779,N_4805);
and U5073 (N_5073,N_4790,N_4895);
and U5074 (N_5074,N_4770,N_4886);
and U5075 (N_5075,N_4810,N_4795);
or U5076 (N_5076,N_4861,N_4885);
xnor U5077 (N_5077,N_4813,N_4968);
nor U5078 (N_5078,N_4834,N_4842);
nor U5079 (N_5079,N_4967,N_4958);
xnor U5080 (N_5080,N_4820,N_4758);
and U5081 (N_5081,N_4788,N_4854);
or U5082 (N_5082,N_4759,N_4893);
nor U5083 (N_5083,N_4827,N_4909);
xnor U5084 (N_5084,N_4774,N_4880);
or U5085 (N_5085,N_4945,N_4993);
nor U5086 (N_5086,N_4876,N_4872);
nand U5087 (N_5087,N_4767,N_4988);
or U5088 (N_5088,N_4891,N_4904);
nor U5089 (N_5089,N_4856,N_4970);
nor U5090 (N_5090,N_4888,N_4792);
xnor U5091 (N_5091,N_4870,N_4852);
or U5092 (N_5092,N_4858,N_4940);
or U5093 (N_5093,N_4910,N_4878);
and U5094 (N_5094,N_4832,N_4807);
or U5095 (N_5095,N_4814,N_4966);
or U5096 (N_5096,N_4831,N_4929);
and U5097 (N_5097,N_4763,N_4986);
and U5098 (N_5098,N_4833,N_4882);
nand U5099 (N_5099,N_4794,N_4901);
xnor U5100 (N_5100,N_4816,N_4815);
xor U5101 (N_5101,N_4766,N_4951);
xor U5102 (N_5102,N_4896,N_4804);
nand U5103 (N_5103,N_4751,N_4887);
xnor U5104 (N_5104,N_4862,N_4840);
or U5105 (N_5105,N_4796,N_4764);
nor U5106 (N_5106,N_4962,N_4845);
nor U5107 (N_5107,N_4853,N_4762);
and U5108 (N_5108,N_4851,N_4871);
nor U5109 (N_5109,N_4936,N_4995);
nor U5110 (N_5110,N_4817,N_4769);
or U5111 (N_5111,N_4920,N_4785);
nor U5112 (N_5112,N_4939,N_4912);
xor U5113 (N_5113,N_4890,N_4869);
xor U5114 (N_5114,N_4930,N_4987);
nor U5115 (N_5115,N_4860,N_4864);
nand U5116 (N_5116,N_4812,N_4996);
and U5117 (N_5117,N_4863,N_4874);
xor U5118 (N_5118,N_4918,N_4994);
nand U5119 (N_5119,N_4991,N_4981);
and U5120 (N_5120,N_4836,N_4973);
or U5121 (N_5121,N_4828,N_4773);
nor U5122 (N_5122,N_4960,N_4894);
or U5123 (N_5123,N_4959,N_4776);
nor U5124 (N_5124,N_4925,N_4928);
and U5125 (N_5125,N_4835,N_4966);
nor U5126 (N_5126,N_4923,N_4899);
nand U5127 (N_5127,N_4955,N_4952);
xnor U5128 (N_5128,N_4994,N_4887);
and U5129 (N_5129,N_4858,N_4771);
nand U5130 (N_5130,N_4803,N_4902);
xnor U5131 (N_5131,N_4769,N_4783);
and U5132 (N_5132,N_4890,N_4881);
or U5133 (N_5133,N_4805,N_4976);
nand U5134 (N_5134,N_4917,N_4781);
and U5135 (N_5135,N_4907,N_4999);
nor U5136 (N_5136,N_4825,N_4842);
and U5137 (N_5137,N_4775,N_4931);
xor U5138 (N_5138,N_4852,N_4931);
nand U5139 (N_5139,N_4881,N_4850);
and U5140 (N_5140,N_4856,N_4990);
xnor U5141 (N_5141,N_4956,N_4994);
and U5142 (N_5142,N_4973,N_4838);
nor U5143 (N_5143,N_4769,N_4892);
nor U5144 (N_5144,N_4776,N_4950);
nor U5145 (N_5145,N_4760,N_4864);
nor U5146 (N_5146,N_4988,N_4832);
or U5147 (N_5147,N_4863,N_4929);
nand U5148 (N_5148,N_4809,N_4898);
nand U5149 (N_5149,N_4844,N_4882);
nor U5150 (N_5150,N_4991,N_4872);
nand U5151 (N_5151,N_4929,N_4835);
and U5152 (N_5152,N_4938,N_4872);
nand U5153 (N_5153,N_4788,N_4779);
xnor U5154 (N_5154,N_4800,N_4860);
or U5155 (N_5155,N_4857,N_4890);
xnor U5156 (N_5156,N_4866,N_4799);
and U5157 (N_5157,N_4915,N_4838);
and U5158 (N_5158,N_4924,N_4912);
nand U5159 (N_5159,N_4823,N_4880);
and U5160 (N_5160,N_4996,N_4976);
and U5161 (N_5161,N_4877,N_4832);
nand U5162 (N_5162,N_4784,N_4974);
or U5163 (N_5163,N_4969,N_4849);
nor U5164 (N_5164,N_4861,N_4849);
and U5165 (N_5165,N_4873,N_4967);
nor U5166 (N_5166,N_4883,N_4824);
or U5167 (N_5167,N_4847,N_4873);
and U5168 (N_5168,N_4760,N_4876);
xnor U5169 (N_5169,N_4906,N_4871);
nand U5170 (N_5170,N_4845,N_4931);
nor U5171 (N_5171,N_4890,N_4936);
xor U5172 (N_5172,N_4840,N_4960);
or U5173 (N_5173,N_4829,N_4971);
and U5174 (N_5174,N_4842,N_4807);
nor U5175 (N_5175,N_4999,N_4925);
and U5176 (N_5176,N_4934,N_4806);
nor U5177 (N_5177,N_4986,N_4888);
xnor U5178 (N_5178,N_4890,N_4776);
and U5179 (N_5179,N_4850,N_4750);
nand U5180 (N_5180,N_4958,N_4841);
and U5181 (N_5181,N_4987,N_4909);
and U5182 (N_5182,N_4828,N_4791);
xor U5183 (N_5183,N_4854,N_4856);
nor U5184 (N_5184,N_4921,N_4978);
nand U5185 (N_5185,N_4777,N_4997);
nor U5186 (N_5186,N_4890,N_4866);
and U5187 (N_5187,N_4810,N_4954);
xnor U5188 (N_5188,N_4937,N_4897);
xnor U5189 (N_5189,N_4835,N_4811);
nor U5190 (N_5190,N_4978,N_4941);
nand U5191 (N_5191,N_4870,N_4925);
or U5192 (N_5192,N_4928,N_4858);
nand U5193 (N_5193,N_4978,N_4917);
nor U5194 (N_5194,N_4990,N_4772);
xor U5195 (N_5195,N_4785,N_4970);
nand U5196 (N_5196,N_4984,N_4902);
nand U5197 (N_5197,N_4797,N_4862);
nor U5198 (N_5198,N_4894,N_4751);
xnor U5199 (N_5199,N_4798,N_4852);
or U5200 (N_5200,N_4787,N_4958);
or U5201 (N_5201,N_4899,N_4859);
nand U5202 (N_5202,N_4975,N_4983);
nand U5203 (N_5203,N_4971,N_4842);
or U5204 (N_5204,N_4887,N_4883);
or U5205 (N_5205,N_4917,N_4770);
xor U5206 (N_5206,N_4946,N_4838);
nor U5207 (N_5207,N_4813,N_4871);
xnor U5208 (N_5208,N_4808,N_4896);
and U5209 (N_5209,N_4966,N_4906);
xnor U5210 (N_5210,N_4956,N_4812);
nand U5211 (N_5211,N_4771,N_4856);
and U5212 (N_5212,N_4817,N_4985);
and U5213 (N_5213,N_4800,N_4813);
nand U5214 (N_5214,N_4970,N_4843);
nand U5215 (N_5215,N_4904,N_4883);
nand U5216 (N_5216,N_4780,N_4932);
xnor U5217 (N_5217,N_4772,N_4959);
nand U5218 (N_5218,N_4809,N_4867);
xnor U5219 (N_5219,N_4836,N_4805);
nor U5220 (N_5220,N_4796,N_4789);
and U5221 (N_5221,N_4898,N_4782);
nand U5222 (N_5222,N_4776,N_4783);
and U5223 (N_5223,N_4823,N_4789);
nor U5224 (N_5224,N_4802,N_4966);
nor U5225 (N_5225,N_4830,N_4877);
and U5226 (N_5226,N_4988,N_4804);
or U5227 (N_5227,N_4937,N_4847);
xnor U5228 (N_5228,N_4856,N_4781);
nor U5229 (N_5229,N_4811,N_4885);
xnor U5230 (N_5230,N_4845,N_4821);
xor U5231 (N_5231,N_4912,N_4848);
nor U5232 (N_5232,N_4912,N_4791);
and U5233 (N_5233,N_4857,N_4923);
xnor U5234 (N_5234,N_4939,N_4975);
nor U5235 (N_5235,N_4819,N_4993);
or U5236 (N_5236,N_4955,N_4971);
nor U5237 (N_5237,N_4778,N_4898);
xor U5238 (N_5238,N_4778,N_4772);
and U5239 (N_5239,N_4894,N_4903);
and U5240 (N_5240,N_4987,N_4897);
xor U5241 (N_5241,N_4764,N_4865);
nor U5242 (N_5242,N_4807,N_4865);
nor U5243 (N_5243,N_4794,N_4954);
xor U5244 (N_5244,N_4911,N_4953);
and U5245 (N_5245,N_4803,N_4872);
xnor U5246 (N_5246,N_4920,N_4876);
and U5247 (N_5247,N_4880,N_4897);
and U5248 (N_5248,N_4954,N_4799);
nand U5249 (N_5249,N_4788,N_4767);
and U5250 (N_5250,N_5052,N_5049);
nand U5251 (N_5251,N_5096,N_5097);
nand U5252 (N_5252,N_5171,N_5087);
xnor U5253 (N_5253,N_5142,N_5086);
nor U5254 (N_5254,N_5125,N_5148);
or U5255 (N_5255,N_5071,N_5139);
xnor U5256 (N_5256,N_5136,N_5245);
nor U5257 (N_5257,N_5181,N_5176);
and U5258 (N_5258,N_5029,N_5064);
and U5259 (N_5259,N_5130,N_5199);
nand U5260 (N_5260,N_5046,N_5188);
or U5261 (N_5261,N_5144,N_5015);
xor U5262 (N_5262,N_5031,N_5111);
and U5263 (N_5263,N_5002,N_5212);
xor U5264 (N_5264,N_5109,N_5075);
or U5265 (N_5265,N_5247,N_5126);
nand U5266 (N_5266,N_5184,N_5113);
nor U5267 (N_5267,N_5070,N_5037);
nor U5268 (N_5268,N_5135,N_5214);
and U5269 (N_5269,N_5057,N_5025);
or U5270 (N_5270,N_5063,N_5090);
nor U5271 (N_5271,N_5106,N_5107);
nor U5272 (N_5272,N_5044,N_5244);
or U5273 (N_5273,N_5116,N_5165);
or U5274 (N_5274,N_5082,N_5124);
or U5275 (N_5275,N_5041,N_5159);
or U5276 (N_5276,N_5168,N_5152);
nand U5277 (N_5277,N_5003,N_5218);
and U5278 (N_5278,N_5153,N_5236);
nand U5279 (N_5279,N_5009,N_5054);
xnor U5280 (N_5280,N_5164,N_5093);
or U5281 (N_5281,N_5206,N_5155);
and U5282 (N_5282,N_5065,N_5095);
or U5283 (N_5283,N_5027,N_5233);
or U5284 (N_5284,N_5022,N_5040);
nand U5285 (N_5285,N_5205,N_5223);
and U5286 (N_5286,N_5024,N_5129);
nand U5287 (N_5287,N_5076,N_5196);
nor U5288 (N_5288,N_5104,N_5201);
xor U5289 (N_5289,N_5230,N_5014);
and U5290 (N_5290,N_5195,N_5121);
and U5291 (N_5291,N_5013,N_5032);
nand U5292 (N_5292,N_5007,N_5043);
xor U5293 (N_5293,N_5157,N_5221);
nand U5294 (N_5294,N_5162,N_5010);
or U5295 (N_5295,N_5118,N_5177);
nand U5296 (N_5296,N_5140,N_5156);
nand U5297 (N_5297,N_5045,N_5098);
xnor U5298 (N_5298,N_5068,N_5114);
and U5299 (N_5299,N_5160,N_5217);
xnor U5300 (N_5300,N_5239,N_5048);
and U5301 (N_5301,N_5018,N_5133);
or U5302 (N_5302,N_5078,N_5035);
nand U5303 (N_5303,N_5163,N_5122);
nand U5304 (N_5304,N_5067,N_5237);
and U5305 (N_5305,N_5209,N_5210);
and U5306 (N_5306,N_5026,N_5175);
or U5307 (N_5307,N_5141,N_5213);
or U5308 (N_5308,N_5241,N_5147);
nand U5309 (N_5309,N_5150,N_5050);
xor U5310 (N_5310,N_5186,N_5085);
nor U5311 (N_5311,N_5169,N_5115);
xnor U5312 (N_5312,N_5231,N_5202);
or U5313 (N_5313,N_5059,N_5038);
nand U5314 (N_5314,N_5047,N_5058);
nand U5315 (N_5315,N_5081,N_5033);
and U5316 (N_5316,N_5051,N_5146);
nor U5317 (N_5317,N_5088,N_5108);
or U5318 (N_5318,N_5017,N_5226);
xor U5319 (N_5319,N_5193,N_5123);
or U5320 (N_5320,N_5006,N_5072);
or U5321 (N_5321,N_5149,N_5232);
and U5322 (N_5322,N_5204,N_5132);
and U5323 (N_5323,N_5220,N_5216);
nor U5324 (N_5324,N_5178,N_5222);
xnor U5325 (N_5325,N_5170,N_5229);
and U5326 (N_5326,N_5119,N_5080);
nor U5327 (N_5327,N_5180,N_5151);
and U5328 (N_5328,N_5145,N_5042);
and U5329 (N_5329,N_5053,N_5174);
and U5330 (N_5330,N_5074,N_5039);
or U5331 (N_5331,N_5127,N_5189);
or U5332 (N_5332,N_5143,N_5099);
xor U5333 (N_5333,N_5154,N_5187);
or U5334 (N_5334,N_5005,N_5228);
xor U5335 (N_5335,N_5182,N_5028);
nand U5336 (N_5336,N_5138,N_5137);
or U5337 (N_5337,N_5083,N_5172);
nor U5338 (N_5338,N_5240,N_5084);
and U5339 (N_5339,N_5060,N_5224);
xnor U5340 (N_5340,N_5248,N_5036);
nand U5341 (N_5341,N_5055,N_5101);
or U5342 (N_5342,N_5077,N_5243);
xnor U5343 (N_5343,N_5012,N_5225);
xor U5344 (N_5344,N_5079,N_5167);
nand U5345 (N_5345,N_5249,N_5004);
and U5346 (N_5346,N_5001,N_5191);
or U5347 (N_5347,N_5134,N_5238);
and U5348 (N_5348,N_5030,N_5219);
xnor U5349 (N_5349,N_5000,N_5131);
nor U5350 (N_5350,N_5117,N_5102);
nand U5351 (N_5351,N_5066,N_5056);
and U5352 (N_5352,N_5161,N_5211);
and U5353 (N_5353,N_5197,N_5179);
nand U5354 (N_5354,N_5194,N_5166);
and U5355 (N_5355,N_5069,N_5192);
or U5356 (N_5356,N_5020,N_5246);
or U5357 (N_5357,N_5235,N_5110);
and U5358 (N_5358,N_5120,N_5208);
nor U5359 (N_5359,N_5021,N_5016);
xnor U5360 (N_5360,N_5011,N_5062);
xor U5361 (N_5361,N_5190,N_5112);
nor U5362 (N_5362,N_5128,N_5094);
xnor U5363 (N_5363,N_5198,N_5091);
xnor U5364 (N_5364,N_5092,N_5242);
nand U5365 (N_5365,N_5061,N_5203);
nor U5366 (N_5366,N_5105,N_5023);
or U5367 (N_5367,N_5185,N_5183);
and U5368 (N_5368,N_5100,N_5227);
nand U5369 (N_5369,N_5008,N_5103);
nor U5370 (N_5370,N_5034,N_5019);
nand U5371 (N_5371,N_5173,N_5207);
or U5372 (N_5372,N_5073,N_5158);
and U5373 (N_5373,N_5089,N_5200);
and U5374 (N_5374,N_5234,N_5215);
and U5375 (N_5375,N_5097,N_5128);
nor U5376 (N_5376,N_5017,N_5199);
nor U5377 (N_5377,N_5111,N_5206);
and U5378 (N_5378,N_5168,N_5085);
and U5379 (N_5379,N_5217,N_5172);
nand U5380 (N_5380,N_5150,N_5156);
nand U5381 (N_5381,N_5175,N_5228);
nor U5382 (N_5382,N_5129,N_5171);
and U5383 (N_5383,N_5056,N_5203);
nor U5384 (N_5384,N_5120,N_5217);
nor U5385 (N_5385,N_5199,N_5160);
xnor U5386 (N_5386,N_5016,N_5034);
and U5387 (N_5387,N_5099,N_5044);
and U5388 (N_5388,N_5100,N_5111);
xor U5389 (N_5389,N_5161,N_5026);
nor U5390 (N_5390,N_5035,N_5058);
nor U5391 (N_5391,N_5014,N_5006);
xor U5392 (N_5392,N_5249,N_5138);
and U5393 (N_5393,N_5151,N_5201);
or U5394 (N_5394,N_5036,N_5129);
nand U5395 (N_5395,N_5208,N_5198);
or U5396 (N_5396,N_5211,N_5129);
and U5397 (N_5397,N_5015,N_5009);
nor U5398 (N_5398,N_5161,N_5077);
nand U5399 (N_5399,N_5055,N_5078);
nand U5400 (N_5400,N_5029,N_5231);
and U5401 (N_5401,N_5211,N_5188);
xor U5402 (N_5402,N_5151,N_5183);
or U5403 (N_5403,N_5006,N_5146);
and U5404 (N_5404,N_5175,N_5064);
xnor U5405 (N_5405,N_5003,N_5104);
xnor U5406 (N_5406,N_5027,N_5202);
nand U5407 (N_5407,N_5004,N_5121);
nand U5408 (N_5408,N_5152,N_5203);
nand U5409 (N_5409,N_5022,N_5041);
nand U5410 (N_5410,N_5242,N_5081);
and U5411 (N_5411,N_5075,N_5190);
or U5412 (N_5412,N_5067,N_5128);
xnor U5413 (N_5413,N_5076,N_5152);
and U5414 (N_5414,N_5089,N_5230);
or U5415 (N_5415,N_5240,N_5088);
nand U5416 (N_5416,N_5009,N_5095);
xor U5417 (N_5417,N_5098,N_5082);
nand U5418 (N_5418,N_5149,N_5212);
and U5419 (N_5419,N_5110,N_5225);
nor U5420 (N_5420,N_5138,N_5169);
nor U5421 (N_5421,N_5093,N_5014);
nor U5422 (N_5422,N_5167,N_5029);
xor U5423 (N_5423,N_5090,N_5082);
or U5424 (N_5424,N_5240,N_5030);
and U5425 (N_5425,N_5212,N_5091);
or U5426 (N_5426,N_5176,N_5213);
nand U5427 (N_5427,N_5056,N_5147);
xor U5428 (N_5428,N_5168,N_5230);
or U5429 (N_5429,N_5045,N_5044);
or U5430 (N_5430,N_5002,N_5192);
or U5431 (N_5431,N_5205,N_5092);
nor U5432 (N_5432,N_5141,N_5028);
xnor U5433 (N_5433,N_5197,N_5146);
xnor U5434 (N_5434,N_5133,N_5121);
xnor U5435 (N_5435,N_5249,N_5136);
and U5436 (N_5436,N_5060,N_5088);
xor U5437 (N_5437,N_5177,N_5046);
xor U5438 (N_5438,N_5185,N_5107);
nand U5439 (N_5439,N_5090,N_5003);
and U5440 (N_5440,N_5080,N_5143);
or U5441 (N_5441,N_5141,N_5187);
xnor U5442 (N_5442,N_5077,N_5064);
xnor U5443 (N_5443,N_5210,N_5100);
and U5444 (N_5444,N_5079,N_5110);
xnor U5445 (N_5445,N_5112,N_5024);
nor U5446 (N_5446,N_5041,N_5194);
nand U5447 (N_5447,N_5160,N_5016);
nor U5448 (N_5448,N_5018,N_5121);
and U5449 (N_5449,N_5171,N_5227);
and U5450 (N_5450,N_5105,N_5010);
nand U5451 (N_5451,N_5017,N_5086);
or U5452 (N_5452,N_5203,N_5025);
or U5453 (N_5453,N_5152,N_5079);
xnor U5454 (N_5454,N_5059,N_5144);
nand U5455 (N_5455,N_5029,N_5143);
and U5456 (N_5456,N_5194,N_5096);
nor U5457 (N_5457,N_5124,N_5050);
and U5458 (N_5458,N_5205,N_5200);
xor U5459 (N_5459,N_5155,N_5082);
or U5460 (N_5460,N_5246,N_5184);
nor U5461 (N_5461,N_5005,N_5011);
or U5462 (N_5462,N_5219,N_5142);
and U5463 (N_5463,N_5110,N_5135);
nor U5464 (N_5464,N_5236,N_5045);
nor U5465 (N_5465,N_5112,N_5162);
or U5466 (N_5466,N_5246,N_5239);
and U5467 (N_5467,N_5152,N_5177);
xor U5468 (N_5468,N_5156,N_5137);
nand U5469 (N_5469,N_5133,N_5230);
xor U5470 (N_5470,N_5014,N_5097);
nand U5471 (N_5471,N_5009,N_5057);
nand U5472 (N_5472,N_5098,N_5213);
nand U5473 (N_5473,N_5013,N_5014);
nand U5474 (N_5474,N_5005,N_5208);
and U5475 (N_5475,N_5007,N_5002);
xor U5476 (N_5476,N_5016,N_5085);
nor U5477 (N_5477,N_5090,N_5120);
xor U5478 (N_5478,N_5015,N_5246);
nor U5479 (N_5479,N_5127,N_5187);
xor U5480 (N_5480,N_5065,N_5119);
nor U5481 (N_5481,N_5077,N_5215);
xor U5482 (N_5482,N_5004,N_5149);
or U5483 (N_5483,N_5102,N_5189);
and U5484 (N_5484,N_5089,N_5105);
and U5485 (N_5485,N_5031,N_5104);
or U5486 (N_5486,N_5113,N_5033);
nand U5487 (N_5487,N_5108,N_5118);
and U5488 (N_5488,N_5147,N_5009);
and U5489 (N_5489,N_5052,N_5059);
nand U5490 (N_5490,N_5156,N_5081);
or U5491 (N_5491,N_5228,N_5018);
or U5492 (N_5492,N_5194,N_5032);
nand U5493 (N_5493,N_5183,N_5115);
xnor U5494 (N_5494,N_5078,N_5219);
and U5495 (N_5495,N_5147,N_5214);
and U5496 (N_5496,N_5027,N_5119);
xor U5497 (N_5497,N_5006,N_5118);
nand U5498 (N_5498,N_5244,N_5226);
xor U5499 (N_5499,N_5127,N_5140);
nor U5500 (N_5500,N_5405,N_5425);
xor U5501 (N_5501,N_5428,N_5438);
nor U5502 (N_5502,N_5416,N_5431);
nor U5503 (N_5503,N_5479,N_5474);
nor U5504 (N_5504,N_5483,N_5486);
xnor U5505 (N_5505,N_5429,N_5415);
nand U5506 (N_5506,N_5304,N_5426);
nor U5507 (N_5507,N_5446,N_5331);
and U5508 (N_5508,N_5396,N_5255);
xnor U5509 (N_5509,N_5273,N_5381);
nand U5510 (N_5510,N_5358,N_5252);
or U5511 (N_5511,N_5349,N_5364);
and U5512 (N_5512,N_5351,N_5263);
nand U5513 (N_5513,N_5414,N_5285);
nand U5514 (N_5514,N_5402,N_5420);
nor U5515 (N_5515,N_5280,N_5475);
nor U5516 (N_5516,N_5250,N_5413);
or U5517 (N_5517,N_5251,N_5366);
and U5518 (N_5518,N_5393,N_5461);
nor U5519 (N_5519,N_5254,N_5394);
and U5520 (N_5520,N_5336,N_5308);
xor U5521 (N_5521,N_5400,N_5344);
nand U5522 (N_5522,N_5452,N_5312);
nand U5523 (N_5523,N_5283,N_5380);
and U5524 (N_5524,N_5318,N_5301);
nor U5525 (N_5525,N_5311,N_5407);
and U5526 (N_5526,N_5499,N_5332);
nor U5527 (N_5527,N_5403,N_5490);
or U5528 (N_5528,N_5302,N_5383);
nand U5529 (N_5529,N_5333,N_5287);
nand U5530 (N_5530,N_5343,N_5496);
or U5531 (N_5531,N_5478,N_5354);
xnor U5532 (N_5532,N_5278,N_5362);
xnor U5533 (N_5533,N_5340,N_5265);
xnor U5534 (N_5534,N_5262,N_5458);
nand U5535 (N_5535,N_5266,N_5307);
nor U5536 (N_5536,N_5495,N_5348);
xnor U5537 (N_5537,N_5445,N_5370);
nor U5538 (N_5538,N_5309,N_5295);
nand U5539 (N_5539,N_5320,N_5417);
nand U5540 (N_5540,N_5433,N_5453);
nand U5541 (N_5541,N_5327,N_5256);
xor U5542 (N_5542,N_5324,N_5338);
nor U5543 (N_5543,N_5377,N_5481);
and U5544 (N_5544,N_5465,N_5471);
xnor U5545 (N_5545,N_5470,N_5390);
and U5546 (N_5546,N_5282,N_5469);
nor U5547 (N_5547,N_5284,N_5401);
or U5548 (N_5548,N_5296,N_5382);
or U5549 (N_5549,N_5257,N_5317);
nand U5550 (N_5550,N_5253,N_5337);
nor U5551 (N_5551,N_5356,N_5488);
nor U5552 (N_5552,N_5480,N_5306);
xnor U5553 (N_5553,N_5374,N_5409);
and U5554 (N_5554,N_5298,N_5325);
xnor U5555 (N_5555,N_5494,N_5436);
xnor U5556 (N_5556,N_5310,N_5261);
or U5557 (N_5557,N_5323,N_5267);
and U5558 (N_5558,N_5321,N_5427);
xor U5559 (N_5559,N_5388,N_5360);
nor U5560 (N_5560,N_5326,N_5449);
nand U5561 (N_5561,N_5375,N_5467);
or U5562 (N_5562,N_5484,N_5447);
or U5563 (N_5563,N_5432,N_5270);
xnor U5564 (N_5564,N_5423,N_5455);
nor U5565 (N_5565,N_5271,N_5493);
xor U5566 (N_5566,N_5339,N_5466);
xnor U5567 (N_5567,N_5411,N_5492);
nor U5568 (N_5568,N_5424,N_5442);
nor U5569 (N_5569,N_5459,N_5286);
xnor U5570 (N_5570,N_5292,N_5462);
or U5571 (N_5571,N_5372,N_5485);
xnor U5572 (N_5572,N_5316,N_5378);
and U5573 (N_5573,N_5443,N_5464);
nand U5574 (N_5574,N_5448,N_5361);
xor U5575 (N_5575,N_5384,N_5305);
xor U5576 (N_5576,N_5497,N_5363);
nand U5577 (N_5577,N_5487,N_5352);
or U5578 (N_5578,N_5389,N_5303);
nand U5579 (N_5579,N_5347,N_5260);
or U5580 (N_5580,N_5258,N_5444);
nand U5581 (N_5581,N_5476,N_5328);
nand U5582 (N_5582,N_5274,N_5440);
and U5583 (N_5583,N_5468,N_5367);
and U5584 (N_5584,N_5281,N_5322);
nor U5585 (N_5585,N_5272,N_5300);
nor U5586 (N_5586,N_5365,N_5435);
xnor U5587 (N_5587,N_5353,N_5451);
and U5588 (N_5588,N_5439,N_5368);
xnor U5589 (N_5589,N_5294,N_5350);
or U5590 (N_5590,N_5376,N_5355);
and U5591 (N_5591,N_5288,N_5450);
and U5592 (N_5592,N_5460,N_5391);
or U5593 (N_5593,N_5290,N_5463);
xnor U5594 (N_5594,N_5275,N_5441);
nor U5595 (N_5595,N_5430,N_5269);
xnor U5596 (N_5596,N_5408,N_5335);
nand U5597 (N_5597,N_5359,N_5264);
nand U5598 (N_5598,N_5419,N_5345);
xor U5599 (N_5599,N_5277,N_5418);
or U5600 (N_5600,N_5434,N_5299);
nand U5601 (N_5601,N_5397,N_5456);
nor U5602 (N_5602,N_5489,N_5385);
or U5603 (N_5603,N_5293,N_5315);
xnor U5604 (N_5604,N_5371,N_5342);
and U5605 (N_5605,N_5373,N_5482);
or U5606 (N_5606,N_5437,N_5457);
xor U5607 (N_5607,N_5491,N_5392);
nor U5608 (N_5608,N_5379,N_5334);
nor U5609 (N_5609,N_5386,N_5279);
xnor U5610 (N_5610,N_5404,N_5395);
or U5611 (N_5611,N_5341,N_5289);
xnor U5612 (N_5612,N_5329,N_5313);
xnor U5613 (N_5613,N_5346,N_5477);
nand U5614 (N_5614,N_5421,N_5410);
xnor U5615 (N_5615,N_5454,N_5473);
xnor U5616 (N_5616,N_5387,N_5422);
xnor U5617 (N_5617,N_5268,N_5399);
xor U5618 (N_5618,N_5319,N_5314);
and U5619 (N_5619,N_5297,N_5276);
xnor U5620 (N_5620,N_5330,N_5498);
nor U5621 (N_5621,N_5406,N_5357);
nor U5622 (N_5622,N_5472,N_5291);
xor U5623 (N_5623,N_5259,N_5369);
and U5624 (N_5624,N_5412,N_5398);
or U5625 (N_5625,N_5318,N_5337);
nor U5626 (N_5626,N_5464,N_5372);
or U5627 (N_5627,N_5356,N_5484);
nor U5628 (N_5628,N_5410,N_5378);
or U5629 (N_5629,N_5262,N_5272);
xnor U5630 (N_5630,N_5343,N_5268);
and U5631 (N_5631,N_5468,N_5321);
and U5632 (N_5632,N_5289,N_5301);
or U5633 (N_5633,N_5349,N_5325);
and U5634 (N_5634,N_5311,N_5375);
nand U5635 (N_5635,N_5460,N_5372);
nor U5636 (N_5636,N_5371,N_5298);
and U5637 (N_5637,N_5264,N_5440);
and U5638 (N_5638,N_5251,N_5422);
xnor U5639 (N_5639,N_5414,N_5367);
xnor U5640 (N_5640,N_5495,N_5313);
and U5641 (N_5641,N_5403,N_5496);
and U5642 (N_5642,N_5422,N_5398);
nor U5643 (N_5643,N_5260,N_5481);
and U5644 (N_5644,N_5343,N_5398);
nand U5645 (N_5645,N_5289,N_5440);
nor U5646 (N_5646,N_5483,N_5359);
xor U5647 (N_5647,N_5389,N_5345);
nor U5648 (N_5648,N_5357,N_5250);
or U5649 (N_5649,N_5369,N_5364);
or U5650 (N_5650,N_5350,N_5385);
xor U5651 (N_5651,N_5350,N_5459);
nand U5652 (N_5652,N_5415,N_5373);
xnor U5653 (N_5653,N_5399,N_5441);
nor U5654 (N_5654,N_5458,N_5334);
and U5655 (N_5655,N_5358,N_5315);
nand U5656 (N_5656,N_5370,N_5317);
xnor U5657 (N_5657,N_5436,N_5439);
nand U5658 (N_5658,N_5446,N_5460);
and U5659 (N_5659,N_5285,N_5438);
and U5660 (N_5660,N_5482,N_5382);
or U5661 (N_5661,N_5320,N_5363);
and U5662 (N_5662,N_5470,N_5322);
or U5663 (N_5663,N_5335,N_5331);
nand U5664 (N_5664,N_5366,N_5261);
or U5665 (N_5665,N_5263,N_5481);
or U5666 (N_5666,N_5376,N_5328);
xnor U5667 (N_5667,N_5470,N_5356);
nor U5668 (N_5668,N_5437,N_5292);
and U5669 (N_5669,N_5263,N_5486);
and U5670 (N_5670,N_5289,N_5472);
and U5671 (N_5671,N_5307,N_5328);
and U5672 (N_5672,N_5392,N_5383);
nor U5673 (N_5673,N_5253,N_5254);
and U5674 (N_5674,N_5440,N_5462);
or U5675 (N_5675,N_5361,N_5347);
nand U5676 (N_5676,N_5492,N_5495);
xor U5677 (N_5677,N_5411,N_5351);
nand U5678 (N_5678,N_5285,N_5344);
xor U5679 (N_5679,N_5433,N_5480);
or U5680 (N_5680,N_5437,N_5495);
xor U5681 (N_5681,N_5302,N_5459);
nor U5682 (N_5682,N_5413,N_5464);
xor U5683 (N_5683,N_5264,N_5352);
or U5684 (N_5684,N_5442,N_5465);
nor U5685 (N_5685,N_5299,N_5279);
xnor U5686 (N_5686,N_5388,N_5468);
and U5687 (N_5687,N_5307,N_5353);
and U5688 (N_5688,N_5299,N_5480);
or U5689 (N_5689,N_5271,N_5374);
or U5690 (N_5690,N_5252,N_5489);
nand U5691 (N_5691,N_5489,N_5390);
nor U5692 (N_5692,N_5386,N_5310);
and U5693 (N_5693,N_5327,N_5369);
nor U5694 (N_5694,N_5290,N_5427);
nand U5695 (N_5695,N_5278,N_5391);
nand U5696 (N_5696,N_5287,N_5293);
nor U5697 (N_5697,N_5413,N_5438);
xor U5698 (N_5698,N_5431,N_5432);
xnor U5699 (N_5699,N_5272,N_5305);
and U5700 (N_5700,N_5326,N_5412);
nand U5701 (N_5701,N_5491,N_5431);
and U5702 (N_5702,N_5478,N_5443);
nand U5703 (N_5703,N_5362,N_5354);
nand U5704 (N_5704,N_5436,N_5413);
xnor U5705 (N_5705,N_5375,N_5465);
xor U5706 (N_5706,N_5399,N_5431);
xnor U5707 (N_5707,N_5391,N_5365);
and U5708 (N_5708,N_5476,N_5423);
nor U5709 (N_5709,N_5419,N_5333);
nand U5710 (N_5710,N_5419,N_5344);
xnor U5711 (N_5711,N_5326,N_5269);
nand U5712 (N_5712,N_5271,N_5335);
nand U5713 (N_5713,N_5441,N_5434);
xnor U5714 (N_5714,N_5308,N_5292);
or U5715 (N_5715,N_5393,N_5433);
and U5716 (N_5716,N_5469,N_5495);
nand U5717 (N_5717,N_5317,N_5482);
nor U5718 (N_5718,N_5260,N_5360);
nand U5719 (N_5719,N_5471,N_5317);
and U5720 (N_5720,N_5448,N_5446);
and U5721 (N_5721,N_5425,N_5452);
and U5722 (N_5722,N_5494,N_5482);
nor U5723 (N_5723,N_5300,N_5264);
xnor U5724 (N_5724,N_5324,N_5418);
or U5725 (N_5725,N_5301,N_5258);
and U5726 (N_5726,N_5277,N_5426);
nor U5727 (N_5727,N_5359,N_5398);
and U5728 (N_5728,N_5415,N_5264);
or U5729 (N_5729,N_5296,N_5338);
and U5730 (N_5730,N_5330,N_5286);
and U5731 (N_5731,N_5441,N_5365);
nand U5732 (N_5732,N_5341,N_5402);
nand U5733 (N_5733,N_5346,N_5374);
or U5734 (N_5734,N_5487,N_5400);
xnor U5735 (N_5735,N_5380,N_5453);
nand U5736 (N_5736,N_5267,N_5489);
nor U5737 (N_5737,N_5411,N_5467);
and U5738 (N_5738,N_5398,N_5402);
or U5739 (N_5739,N_5381,N_5340);
or U5740 (N_5740,N_5441,N_5290);
and U5741 (N_5741,N_5470,N_5430);
nor U5742 (N_5742,N_5440,N_5308);
or U5743 (N_5743,N_5412,N_5361);
and U5744 (N_5744,N_5377,N_5358);
nand U5745 (N_5745,N_5462,N_5302);
and U5746 (N_5746,N_5292,N_5457);
nand U5747 (N_5747,N_5310,N_5273);
nand U5748 (N_5748,N_5416,N_5255);
or U5749 (N_5749,N_5323,N_5414);
or U5750 (N_5750,N_5569,N_5656);
xnor U5751 (N_5751,N_5588,N_5559);
xnor U5752 (N_5752,N_5722,N_5721);
and U5753 (N_5753,N_5577,N_5583);
nor U5754 (N_5754,N_5552,N_5600);
or U5755 (N_5755,N_5503,N_5648);
and U5756 (N_5756,N_5706,N_5595);
xor U5757 (N_5757,N_5695,N_5718);
nand U5758 (N_5758,N_5670,N_5726);
nand U5759 (N_5759,N_5679,N_5635);
nor U5760 (N_5760,N_5568,N_5561);
and U5761 (N_5761,N_5744,N_5547);
xor U5762 (N_5762,N_5748,N_5589);
nand U5763 (N_5763,N_5614,N_5615);
nand U5764 (N_5764,N_5644,N_5541);
xnor U5765 (N_5765,N_5564,N_5729);
nand U5766 (N_5766,N_5657,N_5502);
nor U5767 (N_5767,N_5551,N_5566);
nand U5768 (N_5768,N_5544,N_5620);
nand U5769 (N_5769,N_5654,N_5522);
nand U5770 (N_5770,N_5639,N_5542);
nor U5771 (N_5771,N_5616,N_5701);
or U5772 (N_5772,N_5591,N_5719);
nand U5773 (N_5773,N_5525,N_5578);
and U5774 (N_5774,N_5501,N_5678);
nand U5775 (N_5775,N_5733,N_5675);
nor U5776 (N_5776,N_5709,N_5628);
or U5777 (N_5777,N_5693,N_5734);
nor U5778 (N_5778,N_5554,N_5596);
nand U5779 (N_5779,N_5608,N_5643);
nor U5780 (N_5780,N_5540,N_5563);
xnor U5781 (N_5781,N_5690,N_5747);
or U5782 (N_5782,N_5609,N_5698);
xor U5783 (N_5783,N_5584,N_5691);
nand U5784 (N_5784,N_5619,N_5672);
and U5785 (N_5785,N_5586,N_5731);
nand U5786 (N_5786,N_5611,N_5587);
nand U5787 (N_5787,N_5703,N_5618);
or U5788 (N_5788,N_5562,N_5732);
xor U5789 (N_5789,N_5601,N_5515);
xor U5790 (N_5790,N_5686,N_5711);
or U5791 (N_5791,N_5650,N_5712);
xnor U5792 (N_5792,N_5571,N_5716);
and U5793 (N_5793,N_5521,N_5694);
nor U5794 (N_5794,N_5702,N_5500);
nor U5795 (N_5795,N_5543,N_5518);
nor U5796 (N_5796,N_5524,N_5555);
xnor U5797 (N_5797,N_5574,N_5558);
nand U5798 (N_5798,N_5653,N_5730);
nand U5799 (N_5799,N_5580,N_5681);
and U5800 (N_5800,N_5603,N_5594);
and U5801 (N_5801,N_5667,N_5550);
nand U5802 (N_5802,N_5669,N_5642);
xor U5803 (N_5803,N_5623,N_5740);
nand U5804 (N_5804,N_5590,N_5556);
xnor U5805 (N_5805,N_5570,N_5510);
and U5806 (N_5806,N_5683,N_5560);
nor U5807 (N_5807,N_5508,N_5526);
xnor U5808 (N_5808,N_5607,N_5705);
and U5809 (N_5809,N_5606,N_5724);
nand U5810 (N_5810,N_5743,N_5717);
xnor U5811 (N_5811,N_5520,N_5576);
nor U5812 (N_5812,N_5592,N_5506);
nor U5813 (N_5813,N_5685,N_5626);
xnor U5814 (N_5814,N_5739,N_5687);
and U5815 (N_5815,N_5688,N_5512);
or U5816 (N_5816,N_5636,N_5677);
nand U5817 (N_5817,N_5742,N_5700);
xor U5818 (N_5818,N_5696,N_5599);
or U5819 (N_5819,N_5519,N_5646);
nor U5820 (N_5820,N_5538,N_5523);
nor U5821 (N_5821,N_5707,N_5581);
and U5822 (N_5822,N_5533,N_5708);
and U5823 (N_5823,N_5664,N_5692);
xnor U5824 (N_5824,N_5689,N_5680);
or U5825 (N_5825,N_5668,N_5527);
nand U5826 (N_5826,N_5567,N_5638);
nand U5827 (N_5827,N_5504,N_5684);
or U5828 (N_5828,N_5736,N_5610);
xnor U5829 (N_5829,N_5652,N_5660);
xor U5830 (N_5830,N_5545,N_5661);
and U5831 (N_5831,N_5715,N_5713);
xnor U5832 (N_5832,N_5665,N_5617);
xor U5833 (N_5833,N_5651,N_5659);
and U5834 (N_5834,N_5728,N_5516);
nor U5835 (N_5835,N_5671,N_5676);
nor U5836 (N_5836,N_5629,N_5507);
xnor U5837 (N_5837,N_5714,N_5546);
nor U5838 (N_5838,N_5735,N_5621);
or U5839 (N_5839,N_5674,N_5710);
or U5840 (N_5840,N_5631,N_5645);
nor U5841 (N_5841,N_5604,N_5530);
or U5842 (N_5842,N_5682,N_5622);
and U5843 (N_5843,N_5737,N_5511);
and U5844 (N_5844,N_5597,N_5613);
and U5845 (N_5845,N_5598,N_5579);
xor U5846 (N_5846,N_5529,N_5513);
nor U5847 (N_5847,N_5602,N_5633);
nor U5848 (N_5848,N_5514,N_5535);
or U5849 (N_5849,N_5634,N_5699);
nand U5850 (N_5850,N_5627,N_5572);
nor U5851 (N_5851,N_5557,N_5624);
nor U5852 (N_5852,N_5632,N_5582);
xnor U5853 (N_5853,N_5704,N_5749);
nand U5854 (N_5854,N_5727,N_5528);
nand U5855 (N_5855,N_5630,N_5534);
or U5856 (N_5856,N_5509,N_5658);
or U5857 (N_5857,N_5723,N_5746);
nor U5858 (N_5858,N_5517,N_5738);
or U5859 (N_5859,N_5548,N_5662);
xnor U5860 (N_5860,N_5605,N_5649);
nand U5861 (N_5861,N_5741,N_5593);
and U5862 (N_5862,N_5655,N_5531);
nor U5863 (N_5863,N_5539,N_5666);
xor U5864 (N_5864,N_5537,N_5725);
xor U5865 (N_5865,N_5637,N_5647);
and U5866 (N_5866,N_5536,N_5697);
or U5867 (N_5867,N_5585,N_5720);
nand U5868 (N_5868,N_5673,N_5663);
and U5869 (N_5869,N_5565,N_5573);
or U5870 (N_5870,N_5575,N_5549);
or U5871 (N_5871,N_5625,N_5553);
or U5872 (N_5872,N_5505,N_5745);
or U5873 (N_5873,N_5640,N_5532);
or U5874 (N_5874,N_5641,N_5612);
or U5875 (N_5875,N_5605,N_5629);
or U5876 (N_5876,N_5586,N_5687);
or U5877 (N_5877,N_5615,N_5729);
nor U5878 (N_5878,N_5651,N_5681);
nor U5879 (N_5879,N_5743,N_5537);
nand U5880 (N_5880,N_5734,N_5533);
and U5881 (N_5881,N_5734,N_5686);
or U5882 (N_5882,N_5736,N_5697);
or U5883 (N_5883,N_5694,N_5560);
or U5884 (N_5884,N_5639,N_5628);
or U5885 (N_5885,N_5619,N_5541);
or U5886 (N_5886,N_5733,N_5666);
nor U5887 (N_5887,N_5640,N_5595);
nor U5888 (N_5888,N_5537,N_5509);
xnor U5889 (N_5889,N_5596,N_5591);
nand U5890 (N_5890,N_5604,N_5734);
nand U5891 (N_5891,N_5541,N_5670);
xnor U5892 (N_5892,N_5509,N_5679);
nand U5893 (N_5893,N_5588,N_5528);
xnor U5894 (N_5894,N_5547,N_5628);
xnor U5895 (N_5895,N_5646,N_5645);
nor U5896 (N_5896,N_5747,N_5645);
nor U5897 (N_5897,N_5532,N_5524);
or U5898 (N_5898,N_5551,N_5717);
and U5899 (N_5899,N_5686,N_5581);
nor U5900 (N_5900,N_5731,N_5537);
xnor U5901 (N_5901,N_5708,N_5748);
nand U5902 (N_5902,N_5582,N_5665);
and U5903 (N_5903,N_5610,N_5714);
nor U5904 (N_5904,N_5732,N_5696);
nand U5905 (N_5905,N_5603,N_5625);
or U5906 (N_5906,N_5649,N_5576);
nand U5907 (N_5907,N_5649,N_5503);
xor U5908 (N_5908,N_5735,N_5692);
and U5909 (N_5909,N_5673,N_5722);
xor U5910 (N_5910,N_5652,N_5515);
nand U5911 (N_5911,N_5532,N_5651);
or U5912 (N_5912,N_5535,N_5654);
xnor U5913 (N_5913,N_5673,N_5706);
and U5914 (N_5914,N_5684,N_5710);
nand U5915 (N_5915,N_5677,N_5625);
and U5916 (N_5916,N_5725,N_5727);
xnor U5917 (N_5917,N_5520,N_5600);
nand U5918 (N_5918,N_5655,N_5532);
nand U5919 (N_5919,N_5531,N_5665);
nor U5920 (N_5920,N_5723,N_5558);
nor U5921 (N_5921,N_5607,N_5722);
or U5922 (N_5922,N_5714,N_5547);
and U5923 (N_5923,N_5707,N_5597);
nand U5924 (N_5924,N_5715,N_5644);
nor U5925 (N_5925,N_5650,N_5611);
or U5926 (N_5926,N_5508,N_5728);
or U5927 (N_5927,N_5539,N_5668);
and U5928 (N_5928,N_5565,N_5625);
nand U5929 (N_5929,N_5687,N_5695);
and U5930 (N_5930,N_5689,N_5743);
and U5931 (N_5931,N_5668,N_5643);
nor U5932 (N_5932,N_5562,N_5544);
nor U5933 (N_5933,N_5733,N_5659);
xor U5934 (N_5934,N_5569,N_5564);
nor U5935 (N_5935,N_5684,N_5729);
nor U5936 (N_5936,N_5654,N_5544);
nand U5937 (N_5937,N_5586,N_5743);
nand U5938 (N_5938,N_5559,N_5563);
nor U5939 (N_5939,N_5635,N_5580);
xnor U5940 (N_5940,N_5555,N_5525);
nor U5941 (N_5941,N_5712,N_5540);
xnor U5942 (N_5942,N_5647,N_5654);
nor U5943 (N_5943,N_5701,N_5698);
xor U5944 (N_5944,N_5742,N_5713);
nand U5945 (N_5945,N_5732,N_5643);
xor U5946 (N_5946,N_5502,N_5745);
and U5947 (N_5947,N_5676,N_5737);
xor U5948 (N_5948,N_5632,N_5703);
nand U5949 (N_5949,N_5624,N_5500);
xnor U5950 (N_5950,N_5743,N_5723);
nor U5951 (N_5951,N_5535,N_5569);
or U5952 (N_5952,N_5627,N_5611);
or U5953 (N_5953,N_5602,N_5622);
xnor U5954 (N_5954,N_5593,N_5575);
or U5955 (N_5955,N_5617,N_5735);
and U5956 (N_5956,N_5661,N_5634);
or U5957 (N_5957,N_5634,N_5610);
xor U5958 (N_5958,N_5573,N_5528);
or U5959 (N_5959,N_5737,N_5574);
and U5960 (N_5960,N_5553,N_5685);
nand U5961 (N_5961,N_5622,N_5533);
nand U5962 (N_5962,N_5634,N_5612);
or U5963 (N_5963,N_5630,N_5564);
xnor U5964 (N_5964,N_5641,N_5712);
or U5965 (N_5965,N_5588,N_5687);
xnor U5966 (N_5966,N_5545,N_5599);
and U5967 (N_5967,N_5712,N_5589);
or U5968 (N_5968,N_5512,N_5525);
nor U5969 (N_5969,N_5594,N_5693);
and U5970 (N_5970,N_5621,N_5521);
nand U5971 (N_5971,N_5726,N_5607);
nor U5972 (N_5972,N_5575,N_5557);
xor U5973 (N_5973,N_5553,N_5690);
or U5974 (N_5974,N_5513,N_5506);
nand U5975 (N_5975,N_5617,N_5652);
or U5976 (N_5976,N_5656,N_5747);
nand U5977 (N_5977,N_5688,N_5718);
nor U5978 (N_5978,N_5568,N_5554);
nor U5979 (N_5979,N_5585,N_5642);
nor U5980 (N_5980,N_5743,N_5600);
nand U5981 (N_5981,N_5697,N_5619);
nor U5982 (N_5982,N_5713,N_5505);
nor U5983 (N_5983,N_5668,N_5602);
or U5984 (N_5984,N_5664,N_5661);
or U5985 (N_5985,N_5611,N_5686);
nor U5986 (N_5986,N_5637,N_5563);
nand U5987 (N_5987,N_5627,N_5628);
and U5988 (N_5988,N_5561,N_5538);
and U5989 (N_5989,N_5640,N_5565);
nor U5990 (N_5990,N_5644,N_5531);
xnor U5991 (N_5991,N_5679,N_5567);
and U5992 (N_5992,N_5665,N_5716);
or U5993 (N_5993,N_5540,N_5509);
nand U5994 (N_5994,N_5604,N_5699);
nor U5995 (N_5995,N_5608,N_5653);
and U5996 (N_5996,N_5666,N_5738);
xnor U5997 (N_5997,N_5664,N_5543);
nand U5998 (N_5998,N_5667,N_5739);
and U5999 (N_5999,N_5731,N_5509);
nor U6000 (N_6000,N_5766,N_5893);
nor U6001 (N_6001,N_5953,N_5907);
or U6002 (N_6002,N_5920,N_5877);
xnor U6003 (N_6003,N_5971,N_5935);
nor U6004 (N_6004,N_5934,N_5960);
or U6005 (N_6005,N_5992,N_5933);
xnor U6006 (N_6006,N_5777,N_5886);
nor U6007 (N_6007,N_5758,N_5950);
and U6008 (N_6008,N_5962,N_5987);
and U6009 (N_6009,N_5847,N_5880);
xnor U6010 (N_6010,N_5804,N_5810);
or U6011 (N_6011,N_5913,N_5900);
nor U6012 (N_6012,N_5854,N_5999);
xor U6013 (N_6013,N_5863,N_5883);
and U6014 (N_6014,N_5795,N_5946);
and U6015 (N_6015,N_5957,N_5760);
xnor U6016 (N_6016,N_5836,N_5849);
or U6017 (N_6017,N_5914,N_5927);
nand U6018 (N_6018,N_5846,N_5816);
nor U6019 (N_6019,N_5947,N_5918);
nor U6020 (N_6020,N_5764,N_5970);
or U6021 (N_6021,N_5983,N_5806);
and U6022 (N_6022,N_5955,N_5991);
or U6023 (N_6023,N_5928,N_5945);
nand U6024 (N_6024,N_5871,N_5903);
and U6025 (N_6025,N_5808,N_5974);
nor U6026 (N_6026,N_5936,N_5911);
nor U6027 (N_6027,N_5762,N_5770);
and U6028 (N_6028,N_5985,N_5839);
xnor U6029 (N_6029,N_5790,N_5842);
xor U6030 (N_6030,N_5941,N_5771);
nand U6031 (N_6031,N_5819,N_5862);
xor U6032 (N_6032,N_5759,N_5830);
xor U6033 (N_6033,N_5767,N_5832);
xnor U6034 (N_6034,N_5834,N_5932);
nor U6035 (N_6035,N_5889,N_5856);
nor U6036 (N_6036,N_5898,N_5929);
nand U6037 (N_6037,N_5781,N_5807);
nor U6038 (N_6038,N_5984,N_5772);
and U6039 (N_6039,N_5905,N_5964);
nor U6040 (N_6040,N_5761,N_5969);
nand U6041 (N_6041,N_5958,N_5919);
nand U6042 (N_6042,N_5835,N_5851);
or U6043 (N_6043,N_5861,N_5915);
or U6044 (N_6044,N_5943,N_5850);
nand U6045 (N_6045,N_5848,N_5845);
xnor U6046 (N_6046,N_5809,N_5961);
xnor U6047 (N_6047,N_5859,N_5876);
or U6048 (N_6048,N_5838,N_5949);
or U6049 (N_6049,N_5799,N_5890);
nand U6050 (N_6050,N_5860,N_5986);
or U6051 (N_6051,N_5888,N_5784);
nor U6052 (N_6052,N_5930,N_5908);
nand U6053 (N_6053,N_5925,N_5972);
nor U6054 (N_6054,N_5896,N_5820);
and U6055 (N_6055,N_5973,N_5829);
and U6056 (N_6056,N_5875,N_5811);
xnor U6057 (N_6057,N_5996,N_5786);
xor U6058 (N_6058,N_5872,N_5873);
xor U6059 (N_6059,N_5793,N_5787);
nand U6060 (N_6060,N_5768,N_5754);
nand U6061 (N_6061,N_5874,N_5756);
or U6062 (N_6062,N_5977,N_5884);
nand U6063 (N_6063,N_5942,N_5965);
xnor U6064 (N_6064,N_5878,N_5813);
nand U6065 (N_6065,N_5844,N_5822);
xnor U6066 (N_6066,N_5833,N_5885);
and U6067 (N_6067,N_5881,N_5774);
xnor U6068 (N_6068,N_5892,N_5831);
nand U6069 (N_6069,N_5792,N_5975);
nor U6070 (N_6070,N_5750,N_5870);
or U6071 (N_6071,N_5765,N_5923);
and U6072 (N_6072,N_5773,N_5843);
or U6073 (N_6073,N_5779,N_5828);
or U6074 (N_6074,N_5904,N_5789);
xor U6075 (N_6075,N_5865,N_5858);
xnor U6076 (N_6076,N_5780,N_5864);
and U6077 (N_6077,N_5994,N_5818);
or U6078 (N_6078,N_5823,N_5753);
xor U6079 (N_6079,N_5967,N_5948);
xnor U6080 (N_6080,N_5752,N_5853);
nand U6081 (N_6081,N_5939,N_5866);
xnor U6082 (N_6082,N_5924,N_5937);
xnor U6083 (N_6083,N_5812,N_5827);
nand U6084 (N_6084,N_5794,N_5815);
nor U6085 (N_6085,N_5966,N_5954);
xnor U6086 (N_6086,N_5921,N_5901);
nor U6087 (N_6087,N_5998,N_5990);
nand U6088 (N_6088,N_5887,N_5791);
nand U6089 (N_6089,N_5869,N_5995);
or U6090 (N_6090,N_5951,N_5852);
nand U6091 (N_6091,N_5803,N_5788);
xor U6092 (N_6092,N_5797,N_5963);
or U6093 (N_6093,N_5931,N_5800);
nand U6094 (N_6094,N_5968,N_5897);
nand U6095 (N_6095,N_5769,N_5825);
nor U6096 (N_6096,N_5902,N_5899);
nor U6097 (N_6097,N_5926,N_5978);
or U6098 (N_6098,N_5895,N_5959);
or U6099 (N_6099,N_5805,N_5802);
xor U6100 (N_6100,N_5785,N_5755);
xor U6101 (N_6101,N_5882,N_5976);
and U6102 (N_6102,N_5922,N_5891);
nand U6103 (N_6103,N_5916,N_5940);
and U6104 (N_6104,N_5775,N_5814);
xor U6105 (N_6105,N_5980,N_5956);
xnor U6106 (N_6106,N_5867,N_5824);
and U6107 (N_6107,N_5912,N_5917);
nor U6108 (N_6108,N_5841,N_5840);
and U6109 (N_6109,N_5894,N_5989);
xnor U6110 (N_6110,N_5821,N_5988);
nor U6111 (N_6111,N_5801,N_5944);
xor U6112 (N_6112,N_5763,N_5778);
or U6113 (N_6113,N_5776,N_5981);
xor U6114 (N_6114,N_5783,N_5782);
xor U6115 (N_6115,N_5817,N_5982);
or U6116 (N_6116,N_5938,N_5906);
or U6117 (N_6117,N_5751,N_5952);
xnor U6118 (N_6118,N_5993,N_5909);
and U6119 (N_6119,N_5798,N_5857);
nand U6120 (N_6120,N_5868,N_5997);
or U6121 (N_6121,N_5757,N_5826);
xor U6122 (N_6122,N_5855,N_5910);
nor U6123 (N_6123,N_5979,N_5796);
nor U6124 (N_6124,N_5837,N_5879);
or U6125 (N_6125,N_5850,N_5800);
xor U6126 (N_6126,N_5823,N_5888);
nand U6127 (N_6127,N_5810,N_5924);
or U6128 (N_6128,N_5910,N_5995);
or U6129 (N_6129,N_5939,N_5779);
nor U6130 (N_6130,N_5800,N_5768);
and U6131 (N_6131,N_5885,N_5967);
xnor U6132 (N_6132,N_5941,N_5908);
and U6133 (N_6133,N_5956,N_5997);
nand U6134 (N_6134,N_5840,N_5948);
and U6135 (N_6135,N_5932,N_5777);
xnor U6136 (N_6136,N_5822,N_5931);
xnor U6137 (N_6137,N_5764,N_5757);
xor U6138 (N_6138,N_5940,N_5906);
xor U6139 (N_6139,N_5886,N_5926);
nor U6140 (N_6140,N_5993,N_5930);
xnor U6141 (N_6141,N_5757,N_5906);
nand U6142 (N_6142,N_5943,N_5815);
xor U6143 (N_6143,N_5862,N_5872);
nand U6144 (N_6144,N_5883,N_5796);
nand U6145 (N_6145,N_5921,N_5853);
nor U6146 (N_6146,N_5950,N_5905);
nand U6147 (N_6147,N_5824,N_5806);
nand U6148 (N_6148,N_5906,N_5814);
nand U6149 (N_6149,N_5836,N_5905);
or U6150 (N_6150,N_5776,N_5923);
nor U6151 (N_6151,N_5794,N_5765);
nor U6152 (N_6152,N_5917,N_5787);
xnor U6153 (N_6153,N_5870,N_5918);
and U6154 (N_6154,N_5819,N_5923);
xnor U6155 (N_6155,N_5804,N_5812);
or U6156 (N_6156,N_5911,N_5974);
and U6157 (N_6157,N_5870,N_5777);
xor U6158 (N_6158,N_5883,N_5845);
nand U6159 (N_6159,N_5771,N_5751);
nor U6160 (N_6160,N_5878,N_5786);
or U6161 (N_6161,N_5778,N_5962);
nor U6162 (N_6162,N_5870,N_5786);
nor U6163 (N_6163,N_5800,N_5919);
xnor U6164 (N_6164,N_5856,N_5969);
and U6165 (N_6165,N_5931,N_5951);
or U6166 (N_6166,N_5828,N_5931);
nand U6167 (N_6167,N_5976,N_5954);
xor U6168 (N_6168,N_5773,N_5798);
nor U6169 (N_6169,N_5862,N_5929);
or U6170 (N_6170,N_5959,N_5992);
nor U6171 (N_6171,N_5972,N_5975);
nand U6172 (N_6172,N_5919,N_5848);
and U6173 (N_6173,N_5894,N_5996);
xnor U6174 (N_6174,N_5840,N_5867);
and U6175 (N_6175,N_5785,N_5992);
and U6176 (N_6176,N_5927,N_5959);
or U6177 (N_6177,N_5782,N_5943);
or U6178 (N_6178,N_5836,N_5873);
nor U6179 (N_6179,N_5786,N_5909);
xnor U6180 (N_6180,N_5952,N_5916);
nand U6181 (N_6181,N_5830,N_5899);
nor U6182 (N_6182,N_5868,N_5822);
or U6183 (N_6183,N_5859,N_5940);
xor U6184 (N_6184,N_5772,N_5831);
nand U6185 (N_6185,N_5983,N_5955);
nor U6186 (N_6186,N_5952,N_5974);
nand U6187 (N_6187,N_5940,N_5976);
xor U6188 (N_6188,N_5875,N_5796);
xnor U6189 (N_6189,N_5996,N_5854);
nor U6190 (N_6190,N_5912,N_5973);
xor U6191 (N_6191,N_5818,N_5897);
xor U6192 (N_6192,N_5991,N_5916);
xnor U6193 (N_6193,N_5918,N_5972);
or U6194 (N_6194,N_5928,N_5979);
and U6195 (N_6195,N_5822,N_5836);
nand U6196 (N_6196,N_5989,N_5893);
and U6197 (N_6197,N_5832,N_5840);
and U6198 (N_6198,N_5837,N_5924);
xnor U6199 (N_6199,N_5877,N_5861);
nand U6200 (N_6200,N_5960,N_5820);
xnor U6201 (N_6201,N_5926,N_5913);
nor U6202 (N_6202,N_5777,N_5785);
nand U6203 (N_6203,N_5760,N_5861);
and U6204 (N_6204,N_5750,N_5863);
nor U6205 (N_6205,N_5847,N_5935);
xor U6206 (N_6206,N_5898,N_5893);
xnor U6207 (N_6207,N_5938,N_5799);
nand U6208 (N_6208,N_5825,N_5818);
xor U6209 (N_6209,N_5751,N_5972);
nor U6210 (N_6210,N_5774,N_5889);
and U6211 (N_6211,N_5959,N_5930);
nand U6212 (N_6212,N_5844,N_5974);
and U6213 (N_6213,N_5901,N_5899);
nand U6214 (N_6214,N_5885,N_5753);
nand U6215 (N_6215,N_5983,N_5892);
nor U6216 (N_6216,N_5994,N_5915);
nand U6217 (N_6217,N_5756,N_5837);
or U6218 (N_6218,N_5918,N_5801);
nor U6219 (N_6219,N_5900,N_5826);
and U6220 (N_6220,N_5755,N_5987);
or U6221 (N_6221,N_5887,N_5920);
xor U6222 (N_6222,N_5789,N_5953);
nand U6223 (N_6223,N_5878,N_5869);
or U6224 (N_6224,N_5907,N_5891);
and U6225 (N_6225,N_5801,N_5842);
nor U6226 (N_6226,N_5856,N_5992);
xnor U6227 (N_6227,N_5909,N_5992);
nand U6228 (N_6228,N_5982,N_5839);
nand U6229 (N_6229,N_5771,N_5802);
nand U6230 (N_6230,N_5970,N_5770);
or U6231 (N_6231,N_5841,N_5767);
nand U6232 (N_6232,N_5895,N_5807);
or U6233 (N_6233,N_5998,N_5788);
xor U6234 (N_6234,N_5874,N_5909);
nand U6235 (N_6235,N_5957,N_5965);
or U6236 (N_6236,N_5754,N_5897);
and U6237 (N_6237,N_5877,N_5976);
xor U6238 (N_6238,N_5808,N_5868);
nand U6239 (N_6239,N_5980,N_5874);
nor U6240 (N_6240,N_5913,N_5853);
or U6241 (N_6241,N_5985,N_5811);
xor U6242 (N_6242,N_5970,N_5983);
and U6243 (N_6243,N_5885,N_5978);
nand U6244 (N_6244,N_5974,N_5813);
or U6245 (N_6245,N_5913,N_5994);
nor U6246 (N_6246,N_5761,N_5882);
or U6247 (N_6247,N_5772,N_5970);
nand U6248 (N_6248,N_5995,N_5863);
xnor U6249 (N_6249,N_5936,N_5800);
nor U6250 (N_6250,N_6096,N_6233);
nand U6251 (N_6251,N_6224,N_6151);
and U6252 (N_6252,N_6026,N_6176);
and U6253 (N_6253,N_6015,N_6013);
xor U6254 (N_6254,N_6077,N_6180);
or U6255 (N_6255,N_6241,N_6119);
nand U6256 (N_6256,N_6101,N_6040);
or U6257 (N_6257,N_6060,N_6097);
or U6258 (N_6258,N_6192,N_6243);
and U6259 (N_6259,N_6211,N_6073);
xnor U6260 (N_6260,N_6194,N_6091);
and U6261 (N_6261,N_6152,N_6029);
xnor U6262 (N_6262,N_6126,N_6054);
or U6263 (N_6263,N_6174,N_6093);
xnor U6264 (N_6264,N_6167,N_6076);
nor U6265 (N_6265,N_6129,N_6206);
xor U6266 (N_6266,N_6062,N_6057);
xnor U6267 (N_6267,N_6090,N_6199);
or U6268 (N_6268,N_6136,N_6201);
or U6269 (N_6269,N_6216,N_6186);
xor U6270 (N_6270,N_6113,N_6042);
nand U6271 (N_6271,N_6037,N_6231);
nand U6272 (N_6272,N_6149,N_6132);
or U6273 (N_6273,N_6031,N_6095);
xnor U6274 (N_6274,N_6162,N_6035);
xor U6275 (N_6275,N_6058,N_6014);
nand U6276 (N_6276,N_6247,N_6171);
nand U6277 (N_6277,N_6049,N_6155);
xnor U6278 (N_6278,N_6086,N_6087);
nand U6279 (N_6279,N_6102,N_6160);
xor U6280 (N_6280,N_6238,N_6010);
nand U6281 (N_6281,N_6080,N_6056);
nand U6282 (N_6282,N_6130,N_6222);
xnor U6283 (N_6283,N_6033,N_6084);
or U6284 (N_6284,N_6217,N_6225);
nor U6285 (N_6285,N_6154,N_6190);
nor U6286 (N_6286,N_6147,N_6043);
nor U6287 (N_6287,N_6214,N_6012);
nor U6288 (N_6288,N_6131,N_6107);
or U6289 (N_6289,N_6146,N_6242);
xnor U6290 (N_6290,N_6011,N_6221);
nor U6291 (N_6291,N_6111,N_6127);
nor U6292 (N_6292,N_6065,N_6023);
nor U6293 (N_6293,N_6038,N_6025);
xor U6294 (N_6294,N_6144,N_6178);
and U6295 (N_6295,N_6182,N_6083);
or U6296 (N_6296,N_6220,N_6067);
nor U6297 (N_6297,N_6046,N_6019);
xnor U6298 (N_6298,N_6244,N_6110);
xor U6299 (N_6299,N_6141,N_6226);
xor U6300 (N_6300,N_6179,N_6237);
nand U6301 (N_6301,N_6016,N_6165);
nor U6302 (N_6302,N_6034,N_6169);
nor U6303 (N_6303,N_6064,N_6123);
nand U6304 (N_6304,N_6196,N_6005);
and U6305 (N_6305,N_6234,N_6209);
or U6306 (N_6306,N_6120,N_6175);
nand U6307 (N_6307,N_6204,N_6114);
and U6308 (N_6308,N_6183,N_6134);
and U6309 (N_6309,N_6230,N_6082);
and U6310 (N_6310,N_6198,N_6089);
nand U6311 (N_6311,N_6055,N_6170);
and U6312 (N_6312,N_6164,N_6189);
or U6313 (N_6313,N_6008,N_6195);
and U6314 (N_6314,N_6024,N_6156);
and U6315 (N_6315,N_6092,N_6177);
and U6316 (N_6316,N_6163,N_6105);
nor U6317 (N_6317,N_6103,N_6161);
and U6318 (N_6318,N_6187,N_6041);
or U6319 (N_6319,N_6068,N_6115);
nor U6320 (N_6320,N_6227,N_6124);
nand U6321 (N_6321,N_6071,N_6246);
xnor U6322 (N_6322,N_6248,N_6223);
nor U6323 (N_6323,N_6094,N_6003);
or U6324 (N_6324,N_6061,N_6063);
and U6325 (N_6325,N_6205,N_6020);
nand U6326 (N_6326,N_6050,N_6081);
nor U6327 (N_6327,N_6159,N_6116);
and U6328 (N_6328,N_6240,N_6215);
or U6329 (N_6329,N_6053,N_6036);
or U6330 (N_6330,N_6207,N_6059);
or U6331 (N_6331,N_6000,N_6006);
xnor U6332 (N_6332,N_6007,N_6184);
nor U6333 (N_6333,N_6004,N_6173);
or U6334 (N_6334,N_6001,N_6188);
nor U6335 (N_6335,N_6203,N_6099);
nand U6336 (N_6336,N_6219,N_6021);
or U6337 (N_6337,N_6172,N_6212);
or U6338 (N_6338,N_6200,N_6245);
nor U6339 (N_6339,N_6143,N_6249);
nand U6340 (N_6340,N_6157,N_6229);
or U6341 (N_6341,N_6051,N_6117);
and U6342 (N_6342,N_6139,N_6193);
xnor U6343 (N_6343,N_6191,N_6137);
and U6344 (N_6344,N_6135,N_6032);
nand U6345 (N_6345,N_6133,N_6128);
and U6346 (N_6346,N_6202,N_6145);
nand U6347 (N_6347,N_6079,N_6109);
nand U6348 (N_6348,N_6168,N_6236);
nor U6349 (N_6349,N_6052,N_6108);
nand U6350 (N_6350,N_6045,N_6075);
and U6351 (N_6351,N_6158,N_6085);
nand U6352 (N_6352,N_6166,N_6197);
and U6353 (N_6353,N_6030,N_6150);
nor U6354 (N_6354,N_6148,N_6066);
or U6355 (N_6355,N_6118,N_6140);
and U6356 (N_6356,N_6017,N_6106);
nand U6357 (N_6357,N_6208,N_6122);
xor U6358 (N_6358,N_6112,N_6239);
xor U6359 (N_6359,N_6009,N_6098);
nor U6360 (N_6360,N_6181,N_6125);
or U6361 (N_6361,N_6210,N_6142);
nor U6362 (N_6362,N_6022,N_6185);
xnor U6363 (N_6363,N_6044,N_6002);
or U6364 (N_6364,N_6039,N_6028);
nand U6365 (N_6365,N_6232,N_6100);
xnor U6366 (N_6366,N_6228,N_6027);
xnor U6367 (N_6367,N_6153,N_6074);
nor U6368 (N_6368,N_6218,N_6088);
xor U6369 (N_6369,N_6121,N_6104);
or U6370 (N_6370,N_6047,N_6213);
or U6371 (N_6371,N_6018,N_6078);
xnor U6372 (N_6372,N_6069,N_6138);
xnor U6373 (N_6373,N_6235,N_6048);
xor U6374 (N_6374,N_6072,N_6070);
and U6375 (N_6375,N_6151,N_6050);
or U6376 (N_6376,N_6028,N_6061);
and U6377 (N_6377,N_6030,N_6078);
nand U6378 (N_6378,N_6020,N_6083);
xor U6379 (N_6379,N_6196,N_6009);
or U6380 (N_6380,N_6091,N_6080);
and U6381 (N_6381,N_6165,N_6241);
nor U6382 (N_6382,N_6205,N_6051);
and U6383 (N_6383,N_6186,N_6077);
nand U6384 (N_6384,N_6047,N_6179);
nor U6385 (N_6385,N_6033,N_6191);
or U6386 (N_6386,N_6040,N_6108);
xor U6387 (N_6387,N_6193,N_6060);
xor U6388 (N_6388,N_6117,N_6046);
and U6389 (N_6389,N_6249,N_6149);
xor U6390 (N_6390,N_6211,N_6147);
nand U6391 (N_6391,N_6078,N_6043);
xnor U6392 (N_6392,N_6082,N_6031);
and U6393 (N_6393,N_6060,N_6042);
or U6394 (N_6394,N_6136,N_6112);
xnor U6395 (N_6395,N_6131,N_6196);
or U6396 (N_6396,N_6232,N_6243);
nor U6397 (N_6397,N_6194,N_6017);
xnor U6398 (N_6398,N_6116,N_6163);
xor U6399 (N_6399,N_6168,N_6091);
or U6400 (N_6400,N_6232,N_6114);
nand U6401 (N_6401,N_6096,N_6095);
and U6402 (N_6402,N_6005,N_6024);
xnor U6403 (N_6403,N_6198,N_6162);
xor U6404 (N_6404,N_6117,N_6023);
nand U6405 (N_6405,N_6228,N_6068);
and U6406 (N_6406,N_6065,N_6246);
xor U6407 (N_6407,N_6232,N_6109);
and U6408 (N_6408,N_6215,N_6066);
and U6409 (N_6409,N_6151,N_6149);
and U6410 (N_6410,N_6113,N_6032);
or U6411 (N_6411,N_6053,N_6091);
xnor U6412 (N_6412,N_6161,N_6125);
nor U6413 (N_6413,N_6004,N_6053);
nand U6414 (N_6414,N_6130,N_6003);
nand U6415 (N_6415,N_6243,N_6112);
and U6416 (N_6416,N_6095,N_6214);
and U6417 (N_6417,N_6083,N_6242);
nor U6418 (N_6418,N_6000,N_6123);
nor U6419 (N_6419,N_6022,N_6214);
nor U6420 (N_6420,N_6168,N_6112);
nor U6421 (N_6421,N_6217,N_6162);
xor U6422 (N_6422,N_6165,N_6114);
and U6423 (N_6423,N_6102,N_6174);
and U6424 (N_6424,N_6079,N_6104);
and U6425 (N_6425,N_6183,N_6035);
xnor U6426 (N_6426,N_6136,N_6022);
or U6427 (N_6427,N_6099,N_6003);
nor U6428 (N_6428,N_6054,N_6075);
nor U6429 (N_6429,N_6022,N_6060);
and U6430 (N_6430,N_6246,N_6038);
or U6431 (N_6431,N_6049,N_6081);
and U6432 (N_6432,N_6055,N_6228);
and U6433 (N_6433,N_6080,N_6140);
or U6434 (N_6434,N_6147,N_6032);
nor U6435 (N_6435,N_6048,N_6136);
nor U6436 (N_6436,N_6034,N_6036);
or U6437 (N_6437,N_6001,N_6127);
and U6438 (N_6438,N_6190,N_6085);
nand U6439 (N_6439,N_6241,N_6028);
and U6440 (N_6440,N_6055,N_6123);
nor U6441 (N_6441,N_6026,N_6168);
nand U6442 (N_6442,N_6084,N_6073);
or U6443 (N_6443,N_6140,N_6247);
xnor U6444 (N_6444,N_6170,N_6026);
nor U6445 (N_6445,N_6203,N_6131);
nand U6446 (N_6446,N_6138,N_6214);
and U6447 (N_6447,N_6087,N_6157);
nand U6448 (N_6448,N_6207,N_6061);
xnor U6449 (N_6449,N_6053,N_6139);
or U6450 (N_6450,N_6149,N_6230);
nor U6451 (N_6451,N_6087,N_6057);
nor U6452 (N_6452,N_6214,N_6114);
and U6453 (N_6453,N_6091,N_6106);
nand U6454 (N_6454,N_6240,N_6196);
xnor U6455 (N_6455,N_6028,N_6187);
and U6456 (N_6456,N_6196,N_6059);
nor U6457 (N_6457,N_6105,N_6180);
nand U6458 (N_6458,N_6123,N_6233);
nand U6459 (N_6459,N_6094,N_6045);
nor U6460 (N_6460,N_6123,N_6212);
xnor U6461 (N_6461,N_6177,N_6116);
nor U6462 (N_6462,N_6212,N_6014);
or U6463 (N_6463,N_6097,N_6220);
nor U6464 (N_6464,N_6087,N_6011);
or U6465 (N_6465,N_6088,N_6132);
nand U6466 (N_6466,N_6152,N_6158);
or U6467 (N_6467,N_6096,N_6069);
xnor U6468 (N_6468,N_6172,N_6127);
nor U6469 (N_6469,N_6180,N_6207);
nor U6470 (N_6470,N_6029,N_6168);
nor U6471 (N_6471,N_6124,N_6137);
xnor U6472 (N_6472,N_6089,N_6108);
or U6473 (N_6473,N_6227,N_6186);
nand U6474 (N_6474,N_6083,N_6221);
or U6475 (N_6475,N_6200,N_6166);
and U6476 (N_6476,N_6072,N_6019);
xor U6477 (N_6477,N_6113,N_6014);
xor U6478 (N_6478,N_6200,N_6095);
nand U6479 (N_6479,N_6131,N_6174);
and U6480 (N_6480,N_6240,N_6113);
xor U6481 (N_6481,N_6062,N_6195);
xor U6482 (N_6482,N_6122,N_6124);
and U6483 (N_6483,N_6039,N_6210);
or U6484 (N_6484,N_6246,N_6025);
or U6485 (N_6485,N_6092,N_6228);
or U6486 (N_6486,N_6225,N_6156);
or U6487 (N_6487,N_6109,N_6243);
nor U6488 (N_6488,N_6235,N_6140);
and U6489 (N_6489,N_6093,N_6005);
nand U6490 (N_6490,N_6058,N_6140);
nand U6491 (N_6491,N_6172,N_6091);
or U6492 (N_6492,N_6069,N_6132);
nand U6493 (N_6493,N_6197,N_6082);
nand U6494 (N_6494,N_6021,N_6243);
and U6495 (N_6495,N_6144,N_6026);
xor U6496 (N_6496,N_6011,N_6191);
xnor U6497 (N_6497,N_6242,N_6085);
xor U6498 (N_6498,N_6218,N_6081);
or U6499 (N_6499,N_6171,N_6086);
and U6500 (N_6500,N_6283,N_6481);
xor U6501 (N_6501,N_6330,N_6315);
nor U6502 (N_6502,N_6418,N_6294);
nand U6503 (N_6503,N_6341,N_6395);
xnor U6504 (N_6504,N_6498,N_6253);
nand U6505 (N_6505,N_6484,N_6331);
and U6506 (N_6506,N_6466,N_6348);
xnor U6507 (N_6507,N_6364,N_6404);
nor U6508 (N_6508,N_6363,N_6372);
nor U6509 (N_6509,N_6281,N_6293);
nand U6510 (N_6510,N_6478,N_6270);
xor U6511 (N_6511,N_6384,N_6425);
or U6512 (N_6512,N_6413,N_6426);
nor U6513 (N_6513,N_6491,N_6254);
nor U6514 (N_6514,N_6431,N_6467);
xnor U6515 (N_6515,N_6310,N_6290);
or U6516 (N_6516,N_6366,N_6287);
or U6517 (N_6517,N_6276,N_6439);
xnor U6518 (N_6518,N_6397,N_6311);
or U6519 (N_6519,N_6403,N_6494);
nor U6520 (N_6520,N_6453,N_6409);
and U6521 (N_6521,N_6321,N_6358);
or U6522 (N_6522,N_6252,N_6250);
nand U6523 (N_6523,N_6463,N_6346);
xor U6524 (N_6524,N_6441,N_6393);
nand U6525 (N_6525,N_6324,N_6490);
or U6526 (N_6526,N_6256,N_6492);
nand U6527 (N_6527,N_6452,N_6415);
nor U6528 (N_6528,N_6405,N_6299);
or U6529 (N_6529,N_6303,N_6265);
or U6530 (N_6530,N_6268,N_6308);
nor U6531 (N_6531,N_6455,N_6370);
nand U6532 (N_6532,N_6474,N_6314);
nand U6533 (N_6533,N_6319,N_6318);
nor U6534 (N_6534,N_6386,N_6304);
nand U6535 (N_6535,N_6255,N_6489);
nand U6536 (N_6536,N_6445,N_6416);
and U6537 (N_6537,N_6412,N_6473);
nor U6538 (N_6538,N_6482,N_6266);
nand U6539 (N_6539,N_6450,N_6335);
or U6540 (N_6540,N_6385,N_6406);
xnor U6541 (N_6541,N_6496,N_6329);
nand U6542 (N_6542,N_6320,N_6284);
xnor U6543 (N_6543,N_6343,N_6381);
nor U6544 (N_6544,N_6390,N_6388);
and U6545 (N_6545,N_6355,N_6440);
nor U6546 (N_6546,N_6428,N_6408);
or U6547 (N_6547,N_6407,N_6307);
or U6548 (N_6548,N_6394,N_6485);
or U6549 (N_6549,N_6359,N_6251);
nor U6550 (N_6550,N_6344,N_6471);
and U6551 (N_6551,N_6362,N_6323);
nand U6552 (N_6552,N_6487,N_6479);
and U6553 (N_6553,N_6483,N_6443);
and U6554 (N_6554,N_6387,N_6476);
or U6555 (N_6555,N_6258,N_6295);
and U6556 (N_6556,N_6423,N_6462);
or U6557 (N_6557,N_6279,N_6257);
nor U6558 (N_6558,N_6277,N_6398);
and U6559 (N_6559,N_6396,N_6309);
and U6560 (N_6560,N_6470,N_6419);
nor U6561 (N_6561,N_6264,N_6472);
and U6562 (N_6562,N_6435,N_6437);
nand U6563 (N_6563,N_6424,N_6429);
nand U6564 (N_6564,N_6449,N_6371);
xnor U6565 (N_6565,N_6298,N_6444);
xnor U6566 (N_6566,N_6322,N_6480);
nor U6567 (N_6567,N_6430,N_6414);
nand U6568 (N_6568,N_6340,N_6338);
or U6569 (N_6569,N_6282,N_6300);
xnor U6570 (N_6570,N_6327,N_6325);
xor U6571 (N_6571,N_6417,N_6306);
nor U6572 (N_6572,N_6497,N_6336);
nand U6573 (N_6573,N_6438,N_6273);
nand U6574 (N_6574,N_6392,N_6361);
xor U6575 (N_6575,N_6486,N_6302);
nor U6576 (N_6576,N_6442,N_6349);
xor U6577 (N_6577,N_6451,N_6259);
or U6578 (N_6578,N_6468,N_6456);
and U6579 (N_6579,N_6495,N_6339);
nand U6580 (N_6580,N_6465,N_6305);
nand U6581 (N_6581,N_6289,N_6278);
or U6582 (N_6582,N_6488,N_6313);
or U6583 (N_6583,N_6375,N_6378);
and U6584 (N_6584,N_6368,N_6382);
and U6585 (N_6585,N_6458,N_6334);
nand U6586 (N_6586,N_6499,N_6410);
or U6587 (N_6587,N_6272,N_6354);
or U6588 (N_6588,N_6326,N_6271);
xor U6589 (N_6589,N_6291,N_6317);
nand U6590 (N_6590,N_6475,N_6427);
xnor U6591 (N_6591,N_6493,N_6373);
nand U6592 (N_6592,N_6269,N_6274);
xor U6593 (N_6593,N_6345,N_6275);
nor U6594 (N_6594,N_6477,N_6267);
and U6595 (N_6595,N_6448,N_6433);
nor U6596 (N_6596,N_6360,N_6342);
or U6597 (N_6597,N_6454,N_6389);
nand U6598 (N_6598,N_6337,N_6377);
and U6599 (N_6599,N_6301,N_6263);
or U6600 (N_6600,N_6280,N_6401);
nand U6601 (N_6601,N_6447,N_6333);
and U6602 (N_6602,N_6262,N_6402);
nand U6603 (N_6603,N_6421,N_6446);
nand U6604 (N_6604,N_6461,N_6459);
nor U6605 (N_6605,N_6391,N_6347);
xor U6606 (N_6606,N_6436,N_6420);
xor U6607 (N_6607,N_6399,N_6369);
or U6608 (N_6608,N_6296,N_6357);
nand U6609 (N_6609,N_6261,N_6353);
nand U6610 (N_6610,N_6411,N_6376);
xor U6611 (N_6611,N_6365,N_6286);
xor U6612 (N_6612,N_6383,N_6356);
nand U6613 (N_6613,N_6352,N_6328);
nor U6614 (N_6614,N_6469,N_6460);
nand U6615 (N_6615,N_6422,N_6350);
nand U6616 (N_6616,N_6332,N_6297);
or U6617 (N_6617,N_6457,N_6379);
xnor U6618 (N_6618,N_6464,N_6312);
nor U6619 (N_6619,N_6288,N_6292);
xor U6620 (N_6620,N_6432,N_6380);
and U6621 (N_6621,N_6285,N_6367);
or U6622 (N_6622,N_6351,N_6434);
nor U6623 (N_6623,N_6316,N_6260);
nand U6624 (N_6624,N_6374,N_6400);
nand U6625 (N_6625,N_6260,N_6409);
or U6626 (N_6626,N_6402,N_6466);
or U6627 (N_6627,N_6258,N_6463);
xor U6628 (N_6628,N_6493,N_6332);
nand U6629 (N_6629,N_6344,N_6293);
nand U6630 (N_6630,N_6367,N_6336);
or U6631 (N_6631,N_6453,N_6437);
or U6632 (N_6632,N_6363,N_6485);
nor U6633 (N_6633,N_6297,N_6268);
or U6634 (N_6634,N_6292,N_6300);
nor U6635 (N_6635,N_6360,N_6290);
nand U6636 (N_6636,N_6254,N_6333);
or U6637 (N_6637,N_6364,N_6314);
xnor U6638 (N_6638,N_6476,N_6262);
or U6639 (N_6639,N_6312,N_6452);
and U6640 (N_6640,N_6339,N_6277);
nor U6641 (N_6641,N_6292,N_6439);
xnor U6642 (N_6642,N_6490,N_6323);
or U6643 (N_6643,N_6371,N_6415);
and U6644 (N_6644,N_6492,N_6418);
xor U6645 (N_6645,N_6439,N_6299);
nand U6646 (N_6646,N_6471,N_6437);
and U6647 (N_6647,N_6284,N_6295);
nand U6648 (N_6648,N_6419,N_6382);
nand U6649 (N_6649,N_6303,N_6254);
or U6650 (N_6650,N_6253,N_6481);
xnor U6651 (N_6651,N_6470,N_6398);
nand U6652 (N_6652,N_6454,N_6429);
nor U6653 (N_6653,N_6493,N_6347);
and U6654 (N_6654,N_6392,N_6462);
and U6655 (N_6655,N_6290,N_6485);
or U6656 (N_6656,N_6340,N_6397);
nor U6657 (N_6657,N_6403,N_6365);
nand U6658 (N_6658,N_6253,N_6493);
and U6659 (N_6659,N_6282,N_6345);
and U6660 (N_6660,N_6374,N_6464);
or U6661 (N_6661,N_6476,N_6404);
nor U6662 (N_6662,N_6272,N_6415);
nand U6663 (N_6663,N_6450,N_6418);
nand U6664 (N_6664,N_6268,N_6301);
xnor U6665 (N_6665,N_6406,N_6310);
nand U6666 (N_6666,N_6498,N_6323);
nor U6667 (N_6667,N_6456,N_6439);
nand U6668 (N_6668,N_6387,N_6345);
xnor U6669 (N_6669,N_6390,N_6414);
nand U6670 (N_6670,N_6458,N_6362);
xor U6671 (N_6671,N_6457,N_6341);
and U6672 (N_6672,N_6363,N_6354);
nor U6673 (N_6673,N_6466,N_6305);
and U6674 (N_6674,N_6326,N_6300);
nor U6675 (N_6675,N_6270,N_6373);
nand U6676 (N_6676,N_6465,N_6297);
nor U6677 (N_6677,N_6493,N_6431);
nor U6678 (N_6678,N_6311,N_6483);
nand U6679 (N_6679,N_6431,N_6428);
xnor U6680 (N_6680,N_6271,N_6396);
nand U6681 (N_6681,N_6354,N_6273);
nand U6682 (N_6682,N_6408,N_6285);
or U6683 (N_6683,N_6326,N_6357);
xnor U6684 (N_6684,N_6340,N_6374);
nor U6685 (N_6685,N_6462,N_6261);
nand U6686 (N_6686,N_6464,N_6376);
nand U6687 (N_6687,N_6259,N_6470);
and U6688 (N_6688,N_6431,N_6276);
nor U6689 (N_6689,N_6419,N_6324);
nand U6690 (N_6690,N_6261,N_6278);
xnor U6691 (N_6691,N_6302,N_6392);
nor U6692 (N_6692,N_6480,N_6427);
xnor U6693 (N_6693,N_6462,N_6273);
nor U6694 (N_6694,N_6449,N_6469);
nor U6695 (N_6695,N_6465,N_6403);
and U6696 (N_6696,N_6428,N_6425);
nand U6697 (N_6697,N_6399,N_6401);
nand U6698 (N_6698,N_6363,N_6489);
nor U6699 (N_6699,N_6339,N_6293);
nand U6700 (N_6700,N_6493,N_6370);
xor U6701 (N_6701,N_6367,N_6308);
or U6702 (N_6702,N_6410,N_6398);
xor U6703 (N_6703,N_6274,N_6363);
or U6704 (N_6704,N_6462,N_6257);
nor U6705 (N_6705,N_6389,N_6284);
or U6706 (N_6706,N_6386,N_6427);
xnor U6707 (N_6707,N_6267,N_6431);
and U6708 (N_6708,N_6452,N_6375);
xnor U6709 (N_6709,N_6323,N_6456);
nor U6710 (N_6710,N_6278,N_6379);
or U6711 (N_6711,N_6370,N_6454);
xor U6712 (N_6712,N_6494,N_6364);
xnor U6713 (N_6713,N_6292,N_6374);
or U6714 (N_6714,N_6369,N_6279);
nand U6715 (N_6715,N_6405,N_6273);
xor U6716 (N_6716,N_6371,N_6467);
nand U6717 (N_6717,N_6356,N_6351);
and U6718 (N_6718,N_6284,N_6451);
and U6719 (N_6719,N_6483,N_6269);
nand U6720 (N_6720,N_6290,N_6467);
or U6721 (N_6721,N_6403,N_6473);
nor U6722 (N_6722,N_6385,N_6461);
nand U6723 (N_6723,N_6365,N_6436);
nor U6724 (N_6724,N_6253,N_6279);
xnor U6725 (N_6725,N_6399,N_6312);
nor U6726 (N_6726,N_6297,N_6346);
nor U6727 (N_6727,N_6496,N_6327);
nor U6728 (N_6728,N_6261,N_6494);
nor U6729 (N_6729,N_6480,N_6309);
nand U6730 (N_6730,N_6302,N_6398);
nor U6731 (N_6731,N_6449,N_6297);
and U6732 (N_6732,N_6263,N_6415);
and U6733 (N_6733,N_6274,N_6360);
nand U6734 (N_6734,N_6288,N_6418);
nand U6735 (N_6735,N_6425,N_6335);
and U6736 (N_6736,N_6383,N_6378);
and U6737 (N_6737,N_6488,N_6398);
xnor U6738 (N_6738,N_6252,N_6291);
nor U6739 (N_6739,N_6332,N_6490);
xnor U6740 (N_6740,N_6440,N_6463);
and U6741 (N_6741,N_6482,N_6412);
nor U6742 (N_6742,N_6355,N_6336);
and U6743 (N_6743,N_6333,N_6400);
and U6744 (N_6744,N_6291,N_6413);
and U6745 (N_6745,N_6434,N_6475);
nand U6746 (N_6746,N_6267,N_6352);
and U6747 (N_6747,N_6452,N_6462);
nand U6748 (N_6748,N_6345,N_6465);
nand U6749 (N_6749,N_6350,N_6334);
or U6750 (N_6750,N_6734,N_6631);
nand U6751 (N_6751,N_6725,N_6538);
xnor U6752 (N_6752,N_6690,N_6544);
or U6753 (N_6753,N_6622,N_6739);
or U6754 (N_6754,N_6576,N_6749);
nor U6755 (N_6755,N_6722,N_6558);
or U6756 (N_6756,N_6712,N_6530);
nor U6757 (N_6757,N_6503,N_6587);
and U6758 (N_6758,N_6557,N_6602);
nor U6759 (N_6759,N_6528,N_6523);
nor U6760 (N_6760,N_6646,N_6672);
nor U6761 (N_6761,N_6628,N_6603);
nor U6762 (N_6762,N_6569,N_6556);
nor U6763 (N_6763,N_6651,N_6644);
or U6764 (N_6764,N_6552,N_6521);
and U6765 (N_6765,N_6508,N_6661);
and U6766 (N_6766,N_6529,N_6565);
and U6767 (N_6767,N_6550,N_6667);
and U6768 (N_6768,N_6720,N_6709);
or U6769 (N_6769,N_6633,N_6677);
nand U6770 (N_6770,N_6581,N_6694);
or U6771 (N_6771,N_6669,N_6618);
or U6772 (N_6772,N_6533,N_6572);
nand U6773 (N_6773,N_6684,N_6516);
nand U6774 (N_6774,N_6708,N_6645);
and U6775 (N_6775,N_6500,N_6687);
and U6776 (N_6776,N_6578,N_6619);
nor U6777 (N_6777,N_6674,N_6657);
nand U6778 (N_6778,N_6737,N_6517);
nand U6779 (N_6779,N_6607,N_6616);
xor U6780 (N_6780,N_6600,N_6729);
xor U6781 (N_6781,N_6601,N_6654);
nand U6782 (N_6782,N_6647,N_6553);
xor U6783 (N_6783,N_6717,N_6609);
nor U6784 (N_6784,N_6745,N_6641);
nand U6785 (N_6785,N_6548,N_6649);
nor U6786 (N_6786,N_6748,N_6540);
nor U6787 (N_6787,N_6582,N_6597);
xor U6788 (N_6788,N_6642,N_6696);
xnor U6789 (N_6789,N_6727,N_6704);
or U6790 (N_6790,N_6588,N_6590);
or U6791 (N_6791,N_6698,N_6534);
nor U6792 (N_6792,N_6509,N_6626);
nand U6793 (N_6793,N_6630,N_6728);
nand U6794 (N_6794,N_6736,N_6726);
nand U6795 (N_6795,N_6671,N_6604);
nand U6796 (N_6796,N_6542,N_6716);
nor U6797 (N_6797,N_6697,N_6639);
nand U6798 (N_6798,N_6643,N_6502);
and U6799 (N_6799,N_6514,N_6636);
and U6800 (N_6800,N_6658,N_6732);
xor U6801 (N_6801,N_6614,N_6714);
xor U6802 (N_6802,N_6606,N_6623);
or U6803 (N_6803,N_6613,N_6547);
nor U6804 (N_6804,N_6605,N_6589);
or U6805 (N_6805,N_6515,N_6598);
nand U6806 (N_6806,N_6611,N_6634);
or U6807 (N_6807,N_6585,N_6580);
or U6808 (N_6808,N_6546,N_6656);
nand U6809 (N_6809,N_6568,N_6573);
nand U6810 (N_6810,N_6504,N_6561);
nor U6811 (N_6811,N_6664,N_6525);
xnor U6812 (N_6812,N_6742,N_6705);
or U6813 (N_6813,N_6537,N_6668);
or U6814 (N_6814,N_6678,N_6659);
and U6815 (N_6815,N_6507,N_6543);
nand U6816 (N_6816,N_6738,N_6526);
nor U6817 (N_6817,N_6570,N_6615);
xnor U6818 (N_6818,N_6591,N_6563);
nand U6819 (N_6819,N_6686,N_6715);
nor U6820 (N_6820,N_6711,N_6685);
nor U6821 (N_6821,N_6571,N_6740);
and U6822 (N_6822,N_6741,N_6520);
xor U6823 (N_6823,N_6730,N_6594);
xor U6824 (N_6824,N_6747,N_6662);
xnor U6825 (N_6825,N_6673,N_6701);
and U6826 (N_6826,N_6640,N_6617);
and U6827 (N_6827,N_6596,N_6566);
and U6828 (N_6828,N_6743,N_6718);
and U6829 (N_6829,N_6505,N_6536);
or U6830 (N_6830,N_6638,N_6660);
nor U6831 (N_6831,N_6665,N_6562);
nor U6832 (N_6832,N_6652,N_6692);
nand U6833 (N_6833,N_6612,N_6555);
nor U6834 (N_6834,N_6621,N_6532);
nand U6835 (N_6835,N_6522,N_6731);
nor U6836 (N_6836,N_6527,N_6511);
nand U6837 (N_6837,N_6599,N_6695);
and U6838 (N_6838,N_6567,N_6702);
nand U6839 (N_6839,N_6531,N_6512);
and U6840 (N_6840,N_6577,N_6635);
xnor U6841 (N_6841,N_6524,N_6501);
nand U6842 (N_6842,N_6584,N_6625);
nor U6843 (N_6843,N_6549,N_6683);
or U6844 (N_6844,N_6650,N_6719);
or U6845 (N_6845,N_6608,N_6575);
nor U6846 (N_6846,N_6551,N_6666);
or U6847 (N_6847,N_6682,N_6535);
nor U6848 (N_6848,N_6691,N_6513);
and U6849 (N_6849,N_6627,N_6703);
nand U6850 (N_6850,N_6632,N_6541);
and U6851 (N_6851,N_6653,N_6699);
nand U6852 (N_6852,N_6545,N_6539);
or U6853 (N_6853,N_6680,N_6560);
nand U6854 (N_6854,N_6721,N_6554);
nand U6855 (N_6855,N_6746,N_6663);
or U6856 (N_6856,N_6655,N_6620);
and U6857 (N_6857,N_6564,N_6610);
or U6858 (N_6858,N_6592,N_6579);
or U6859 (N_6859,N_6689,N_6724);
nand U6860 (N_6860,N_6723,N_6629);
nor U6861 (N_6861,N_6681,N_6583);
nand U6862 (N_6862,N_6733,N_6676);
nor U6863 (N_6863,N_6679,N_6707);
nand U6864 (N_6864,N_6675,N_6735);
and U6865 (N_6865,N_6710,N_6586);
xor U6866 (N_6866,N_6637,N_6559);
or U6867 (N_6867,N_6706,N_6593);
xnor U6868 (N_6868,N_6693,N_6510);
nand U6869 (N_6869,N_6518,N_6700);
and U6870 (N_6870,N_6519,N_6648);
nor U6871 (N_6871,N_6688,N_6506);
nor U6872 (N_6872,N_6624,N_6574);
and U6873 (N_6873,N_6670,N_6713);
or U6874 (N_6874,N_6744,N_6595);
xor U6875 (N_6875,N_6520,N_6603);
and U6876 (N_6876,N_6527,N_6719);
nand U6877 (N_6877,N_6689,N_6649);
nand U6878 (N_6878,N_6733,N_6553);
xor U6879 (N_6879,N_6636,N_6571);
xor U6880 (N_6880,N_6521,N_6722);
xor U6881 (N_6881,N_6673,N_6730);
nor U6882 (N_6882,N_6576,N_6500);
nand U6883 (N_6883,N_6707,N_6723);
nor U6884 (N_6884,N_6720,N_6673);
nor U6885 (N_6885,N_6678,N_6696);
xnor U6886 (N_6886,N_6615,N_6565);
and U6887 (N_6887,N_6507,N_6684);
nand U6888 (N_6888,N_6674,N_6654);
nand U6889 (N_6889,N_6632,N_6740);
nand U6890 (N_6890,N_6628,N_6608);
and U6891 (N_6891,N_6547,N_6509);
nor U6892 (N_6892,N_6573,N_6686);
nand U6893 (N_6893,N_6727,N_6522);
nand U6894 (N_6894,N_6524,N_6602);
nand U6895 (N_6895,N_6735,N_6558);
nand U6896 (N_6896,N_6649,N_6703);
nor U6897 (N_6897,N_6735,N_6622);
nand U6898 (N_6898,N_6665,N_6533);
xnor U6899 (N_6899,N_6743,N_6687);
nor U6900 (N_6900,N_6557,N_6567);
nand U6901 (N_6901,N_6624,N_6507);
nor U6902 (N_6902,N_6591,N_6666);
xor U6903 (N_6903,N_6536,N_6530);
xnor U6904 (N_6904,N_6548,N_6521);
nand U6905 (N_6905,N_6703,N_6607);
or U6906 (N_6906,N_6714,N_6549);
or U6907 (N_6907,N_6556,N_6692);
and U6908 (N_6908,N_6679,N_6543);
or U6909 (N_6909,N_6561,N_6582);
xor U6910 (N_6910,N_6639,N_6626);
xor U6911 (N_6911,N_6554,N_6526);
nor U6912 (N_6912,N_6611,N_6737);
nand U6913 (N_6913,N_6651,N_6670);
or U6914 (N_6914,N_6695,N_6509);
or U6915 (N_6915,N_6542,N_6647);
or U6916 (N_6916,N_6610,N_6615);
or U6917 (N_6917,N_6577,N_6542);
nand U6918 (N_6918,N_6699,N_6570);
nand U6919 (N_6919,N_6618,N_6523);
and U6920 (N_6920,N_6559,N_6519);
or U6921 (N_6921,N_6562,N_6689);
xnor U6922 (N_6922,N_6695,N_6536);
nor U6923 (N_6923,N_6738,N_6605);
nand U6924 (N_6924,N_6742,N_6745);
nand U6925 (N_6925,N_6625,N_6717);
or U6926 (N_6926,N_6717,N_6641);
and U6927 (N_6927,N_6640,N_6747);
or U6928 (N_6928,N_6642,N_6520);
xnor U6929 (N_6929,N_6712,N_6567);
and U6930 (N_6930,N_6743,N_6616);
xnor U6931 (N_6931,N_6593,N_6644);
nor U6932 (N_6932,N_6667,N_6595);
or U6933 (N_6933,N_6619,N_6541);
or U6934 (N_6934,N_6609,N_6650);
nor U6935 (N_6935,N_6503,N_6694);
nor U6936 (N_6936,N_6609,N_6543);
nor U6937 (N_6937,N_6515,N_6724);
or U6938 (N_6938,N_6648,N_6507);
or U6939 (N_6939,N_6636,N_6643);
nand U6940 (N_6940,N_6737,N_6572);
xor U6941 (N_6941,N_6523,N_6558);
xor U6942 (N_6942,N_6631,N_6549);
nor U6943 (N_6943,N_6633,N_6585);
xnor U6944 (N_6944,N_6511,N_6504);
nor U6945 (N_6945,N_6620,N_6631);
and U6946 (N_6946,N_6714,N_6648);
nor U6947 (N_6947,N_6697,N_6538);
and U6948 (N_6948,N_6509,N_6740);
nand U6949 (N_6949,N_6520,N_6513);
and U6950 (N_6950,N_6540,N_6714);
and U6951 (N_6951,N_6530,N_6612);
and U6952 (N_6952,N_6604,N_6597);
or U6953 (N_6953,N_6716,N_6719);
or U6954 (N_6954,N_6528,N_6734);
nor U6955 (N_6955,N_6592,N_6544);
and U6956 (N_6956,N_6582,N_6599);
nor U6957 (N_6957,N_6724,N_6695);
nand U6958 (N_6958,N_6685,N_6501);
or U6959 (N_6959,N_6725,N_6721);
nand U6960 (N_6960,N_6716,N_6599);
xor U6961 (N_6961,N_6610,N_6541);
xor U6962 (N_6962,N_6591,N_6536);
xor U6963 (N_6963,N_6507,N_6506);
and U6964 (N_6964,N_6543,N_6567);
nand U6965 (N_6965,N_6648,N_6667);
or U6966 (N_6966,N_6651,N_6603);
and U6967 (N_6967,N_6546,N_6627);
nor U6968 (N_6968,N_6702,N_6727);
nand U6969 (N_6969,N_6634,N_6683);
or U6970 (N_6970,N_6510,N_6582);
xnor U6971 (N_6971,N_6536,N_6576);
and U6972 (N_6972,N_6651,N_6664);
or U6973 (N_6973,N_6577,N_6591);
or U6974 (N_6974,N_6555,N_6643);
xor U6975 (N_6975,N_6564,N_6693);
xnor U6976 (N_6976,N_6721,N_6635);
or U6977 (N_6977,N_6680,N_6519);
or U6978 (N_6978,N_6735,N_6639);
nor U6979 (N_6979,N_6553,N_6666);
xor U6980 (N_6980,N_6732,N_6700);
xor U6981 (N_6981,N_6643,N_6501);
and U6982 (N_6982,N_6731,N_6626);
or U6983 (N_6983,N_6696,N_6554);
xnor U6984 (N_6984,N_6697,N_6562);
xnor U6985 (N_6985,N_6612,N_6709);
and U6986 (N_6986,N_6742,N_6522);
and U6987 (N_6987,N_6729,N_6593);
nor U6988 (N_6988,N_6730,N_6704);
nor U6989 (N_6989,N_6589,N_6633);
nor U6990 (N_6990,N_6624,N_6522);
and U6991 (N_6991,N_6744,N_6742);
nand U6992 (N_6992,N_6743,N_6543);
xnor U6993 (N_6993,N_6546,N_6745);
nor U6994 (N_6994,N_6724,N_6567);
nand U6995 (N_6995,N_6662,N_6564);
and U6996 (N_6996,N_6695,N_6614);
or U6997 (N_6997,N_6733,N_6582);
or U6998 (N_6998,N_6560,N_6729);
and U6999 (N_6999,N_6633,N_6548);
or U7000 (N_7000,N_6912,N_6908);
xnor U7001 (N_7001,N_6941,N_6835);
nand U7002 (N_7002,N_6988,N_6878);
nand U7003 (N_7003,N_6994,N_6825);
xnor U7004 (N_7004,N_6942,N_6961);
nand U7005 (N_7005,N_6872,N_6924);
nor U7006 (N_7006,N_6809,N_6867);
nand U7007 (N_7007,N_6896,N_6863);
and U7008 (N_7008,N_6767,N_6976);
xnor U7009 (N_7009,N_6894,N_6783);
xnor U7010 (N_7010,N_6773,N_6937);
xor U7011 (N_7011,N_6965,N_6876);
nand U7012 (N_7012,N_6926,N_6819);
xor U7013 (N_7013,N_6887,N_6800);
xor U7014 (N_7014,N_6815,N_6838);
and U7015 (N_7015,N_6962,N_6877);
nand U7016 (N_7016,N_6852,N_6890);
or U7017 (N_7017,N_6788,N_6799);
and U7018 (N_7018,N_6834,N_6824);
xnor U7019 (N_7019,N_6957,N_6880);
nand U7020 (N_7020,N_6810,N_6861);
xnor U7021 (N_7021,N_6911,N_6780);
or U7022 (N_7022,N_6946,N_6998);
nand U7023 (N_7023,N_6982,N_6794);
xor U7024 (N_7024,N_6903,N_6768);
nor U7025 (N_7025,N_6847,N_6980);
and U7026 (N_7026,N_6811,N_6820);
nand U7027 (N_7027,N_6906,N_6918);
or U7028 (N_7028,N_6923,N_6921);
and U7029 (N_7029,N_6754,N_6977);
and U7030 (N_7030,N_6840,N_6856);
nand U7031 (N_7031,N_6904,N_6944);
xnor U7032 (N_7032,N_6983,N_6750);
xor U7033 (N_7033,N_6868,N_6936);
and U7034 (N_7034,N_6857,N_6789);
nand U7035 (N_7035,N_6764,N_6949);
and U7036 (N_7036,N_6828,N_6855);
and U7037 (N_7037,N_6902,N_6948);
nor U7038 (N_7038,N_6973,N_6837);
xor U7039 (N_7039,N_6844,N_6755);
and U7040 (N_7040,N_6845,N_6774);
or U7041 (N_7041,N_6785,N_6969);
or U7042 (N_7042,N_6787,N_6757);
and U7043 (N_7043,N_6939,N_6829);
nand U7044 (N_7044,N_6790,N_6843);
nand U7045 (N_7045,N_6899,N_6934);
xnor U7046 (N_7046,N_6905,N_6882);
and U7047 (N_7047,N_6895,N_6752);
nand U7048 (N_7048,N_6920,N_6771);
nor U7049 (N_7049,N_6953,N_6897);
xor U7050 (N_7050,N_6805,N_6816);
or U7051 (N_7051,N_6830,N_6913);
or U7052 (N_7052,N_6874,N_6889);
nand U7053 (N_7053,N_6821,N_6968);
or U7054 (N_7054,N_6818,N_6963);
nand U7055 (N_7055,N_6823,N_6893);
xor U7056 (N_7056,N_6802,N_6775);
nor U7057 (N_7057,N_6925,N_6986);
or U7058 (N_7058,N_6971,N_6884);
or U7059 (N_7059,N_6756,N_6807);
nor U7060 (N_7060,N_6778,N_6827);
nand U7061 (N_7061,N_6916,N_6769);
nor U7062 (N_7062,N_6833,N_6964);
xnor U7063 (N_7063,N_6770,N_6801);
and U7064 (N_7064,N_6883,N_6761);
and U7065 (N_7065,N_6786,N_6766);
nor U7066 (N_7066,N_6808,N_6832);
nand U7067 (N_7067,N_6960,N_6974);
nand U7068 (N_7068,N_6952,N_6929);
or U7069 (N_7069,N_6814,N_6782);
or U7070 (N_7070,N_6922,N_6991);
or U7071 (N_7071,N_6781,N_6993);
or U7072 (N_7072,N_6853,N_6812);
or U7073 (N_7073,N_6917,N_6846);
xor U7074 (N_7074,N_6898,N_6792);
nand U7075 (N_7075,N_6772,N_6915);
xor U7076 (N_7076,N_6959,N_6866);
nand U7077 (N_7077,N_6854,N_6839);
xnor U7078 (N_7078,N_6901,N_6940);
xnor U7079 (N_7079,N_6813,N_6870);
nor U7080 (N_7080,N_6871,N_6975);
xor U7081 (N_7081,N_6989,N_6806);
and U7082 (N_7082,N_6900,N_6945);
and U7083 (N_7083,N_6987,N_6979);
nor U7084 (N_7084,N_6981,N_6763);
and U7085 (N_7085,N_6933,N_6803);
and U7086 (N_7086,N_6985,N_6875);
xnor U7087 (N_7087,N_6888,N_6795);
or U7088 (N_7088,N_6762,N_6892);
and U7089 (N_7089,N_6950,N_6848);
or U7090 (N_7090,N_6841,N_6784);
and U7091 (N_7091,N_6927,N_6751);
xor U7092 (N_7092,N_6885,N_6955);
and U7093 (N_7093,N_6958,N_6860);
and U7094 (N_7094,N_6760,N_6966);
and U7095 (N_7095,N_6836,N_6817);
nor U7096 (N_7096,N_6851,N_6858);
nor U7097 (N_7097,N_6753,N_6992);
or U7098 (N_7098,N_6869,N_6997);
nand U7099 (N_7099,N_6797,N_6777);
nand U7100 (N_7100,N_6930,N_6990);
xor U7101 (N_7101,N_6938,N_6842);
xnor U7102 (N_7102,N_6910,N_6970);
or U7103 (N_7103,N_6779,N_6931);
nand U7104 (N_7104,N_6865,N_6956);
nand U7105 (N_7105,N_6864,N_6859);
or U7106 (N_7106,N_6862,N_6996);
and U7107 (N_7107,N_6873,N_6850);
nor U7108 (N_7108,N_6849,N_6914);
xnor U7109 (N_7109,N_6793,N_6891);
or U7110 (N_7110,N_6984,N_6967);
nand U7111 (N_7111,N_6826,N_6954);
nand U7112 (N_7112,N_6995,N_6879);
nor U7113 (N_7113,N_6791,N_6798);
and U7114 (N_7114,N_6907,N_6928);
xor U7115 (N_7115,N_6765,N_6759);
xor U7116 (N_7116,N_6999,N_6935);
xor U7117 (N_7117,N_6831,N_6804);
nor U7118 (N_7118,N_6932,N_6919);
nor U7119 (N_7119,N_6881,N_6947);
xor U7120 (N_7120,N_6909,N_6796);
nand U7121 (N_7121,N_6972,N_6758);
or U7122 (N_7122,N_6822,N_6776);
nor U7123 (N_7123,N_6951,N_6886);
xnor U7124 (N_7124,N_6943,N_6978);
xnor U7125 (N_7125,N_6969,N_6872);
nor U7126 (N_7126,N_6811,N_6995);
nand U7127 (N_7127,N_6863,N_6819);
xnor U7128 (N_7128,N_6802,N_6816);
nand U7129 (N_7129,N_6913,N_6768);
or U7130 (N_7130,N_6794,N_6987);
xor U7131 (N_7131,N_6942,N_6999);
nor U7132 (N_7132,N_6773,N_6766);
nand U7133 (N_7133,N_6773,N_6844);
nand U7134 (N_7134,N_6925,N_6984);
xor U7135 (N_7135,N_6965,N_6993);
xor U7136 (N_7136,N_6771,N_6767);
and U7137 (N_7137,N_6843,N_6802);
nor U7138 (N_7138,N_6975,N_6831);
xnor U7139 (N_7139,N_6854,N_6893);
nor U7140 (N_7140,N_6993,N_6783);
nor U7141 (N_7141,N_6808,N_6868);
and U7142 (N_7142,N_6934,N_6956);
nor U7143 (N_7143,N_6872,N_6807);
or U7144 (N_7144,N_6773,N_6936);
nand U7145 (N_7145,N_6783,N_6964);
and U7146 (N_7146,N_6810,N_6823);
or U7147 (N_7147,N_6857,N_6932);
or U7148 (N_7148,N_6764,N_6994);
nand U7149 (N_7149,N_6990,N_6897);
nand U7150 (N_7150,N_6990,N_6767);
nor U7151 (N_7151,N_6917,N_6897);
nor U7152 (N_7152,N_6998,N_6872);
nand U7153 (N_7153,N_6880,N_6864);
nand U7154 (N_7154,N_6923,N_6942);
or U7155 (N_7155,N_6759,N_6807);
and U7156 (N_7156,N_6976,N_6811);
and U7157 (N_7157,N_6979,N_6898);
or U7158 (N_7158,N_6909,N_6752);
xnor U7159 (N_7159,N_6801,N_6755);
or U7160 (N_7160,N_6987,N_6972);
nor U7161 (N_7161,N_6971,N_6817);
or U7162 (N_7162,N_6831,N_6933);
xor U7163 (N_7163,N_6889,N_6818);
nor U7164 (N_7164,N_6879,N_6967);
nor U7165 (N_7165,N_6859,N_6946);
nand U7166 (N_7166,N_6805,N_6772);
or U7167 (N_7167,N_6760,N_6807);
and U7168 (N_7168,N_6931,N_6941);
and U7169 (N_7169,N_6762,N_6956);
or U7170 (N_7170,N_6983,N_6842);
xor U7171 (N_7171,N_6869,N_6815);
and U7172 (N_7172,N_6995,N_6812);
nand U7173 (N_7173,N_6925,N_6950);
or U7174 (N_7174,N_6958,N_6985);
nor U7175 (N_7175,N_6792,N_6885);
nand U7176 (N_7176,N_6774,N_6825);
xor U7177 (N_7177,N_6814,N_6932);
nand U7178 (N_7178,N_6812,N_6750);
nor U7179 (N_7179,N_6946,N_6851);
xnor U7180 (N_7180,N_6997,N_6842);
xnor U7181 (N_7181,N_6881,N_6959);
and U7182 (N_7182,N_6948,N_6931);
nand U7183 (N_7183,N_6796,N_6764);
xor U7184 (N_7184,N_6859,N_6987);
nand U7185 (N_7185,N_6833,N_6985);
or U7186 (N_7186,N_6794,N_6923);
and U7187 (N_7187,N_6908,N_6902);
nand U7188 (N_7188,N_6836,N_6952);
or U7189 (N_7189,N_6789,N_6996);
nand U7190 (N_7190,N_6762,N_6931);
xnor U7191 (N_7191,N_6800,N_6805);
nor U7192 (N_7192,N_6960,N_6946);
nor U7193 (N_7193,N_6928,N_6992);
xnor U7194 (N_7194,N_6970,N_6852);
and U7195 (N_7195,N_6760,N_6887);
xnor U7196 (N_7196,N_6967,N_6823);
or U7197 (N_7197,N_6992,N_6752);
nor U7198 (N_7198,N_6999,N_6837);
xor U7199 (N_7199,N_6984,N_6894);
or U7200 (N_7200,N_6808,N_6912);
and U7201 (N_7201,N_6788,N_6751);
nand U7202 (N_7202,N_6895,N_6891);
xnor U7203 (N_7203,N_6993,N_6827);
or U7204 (N_7204,N_6756,N_6776);
nor U7205 (N_7205,N_6807,N_6980);
and U7206 (N_7206,N_6961,N_6762);
nor U7207 (N_7207,N_6935,N_6986);
and U7208 (N_7208,N_6971,N_6949);
or U7209 (N_7209,N_6845,N_6968);
nand U7210 (N_7210,N_6886,N_6797);
and U7211 (N_7211,N_6853,N_6919);
xor U7212 (N_7212,N_6781,N_6978);
nor U7213 (N_7213,N_6936,N_6889);
xnor U7214 (N_7214,N_6879,N_6890);
or U7215 (N_7215,N_6888,N_6953);
nand U7216 (N_7216,N_6895,N_6866);
and U7217 (N_7217,N_6942,N_6758);
nor U7218 (N_7218,N_6818,N_6980);
or U7219 (N_7219,N_6869,N_6878);
or U7220 (N_7220,N_6851,N_6771);
xnor U7221 (N_7221,N_6862,N_6761);
xor U7222 (N_7222,N_6762,N_6932);
or U7223 (N_7223,N_6915,N_6896);
or U7224 (N_7224,N_6939,N_6770);
nor U7225 (N_7225,N_6904,N_6826);
or U7226 (N_7226,N_6901,N_6778);
nor U7227 (N_7227,N_6989,N_6910);
or U7228 (N_7228,N_6765,N_6931);
or U7229 (N_7229,N_6948,N_6953);
nor U7230 (N_7230,N_6847,N_6990);
nand U7231 (N_7231,N_6785,N_6949);
nand U7232 (N_7232,N_6946,N_6918);
or U7233 (N_7233,N_6832,N_6847);
and U7234 (N_7234,N_6814,N_6921);
nor U7235 (N_7235,N_6943,N_6938);
nand U7236 (N_7236,N_6908,N_6879);
nand U7237 (N_7237,N_6920,N_6890);
and U7238 (N_7238,N_6916,N_6799);
nand U7239 (N_7239,N_6780,N_6944);
nand U7240 (N_7240,N_6901,N_6897);
and U7241 (N_7241,N_6866,N_6756);
and U7242 (N_7242,N_6885,N_6950);
nand U7243 (N_7243,N_6863,N_6795);
and U7244 (N_7244,N_6825,N_6861);
nand U7245 (N_7245,N_6790,N_6987);
nor U7246 (N_7246,N_6927,N_6979);
and U7247 (N_7247,N_6887,N_6764);
nand U7248 (N_7248,N_6788,N_6899);
nor U7249 (N_7249,N_6791,N_6903);
or U7250 (N_7250,N_7028,N_7019);
or U7251 (N_7251,N_7031,N_7163);
and U7252 (N_7252,N_7158,N_7212);
and U7253 (N_7253,N_7110,N_7011);
xnor U7254 (N_7254,N_7085,N_7190);
nand U7255 (N_7255,N_7153,N_7173);
xor U7256 (N_7256,N_7225,N_7146);
xnor U7257 (N_7257,N_7125,N_7160);
and U7258 (N_7258,N_7023,N_7042);
xnor U7259 (N_7259,N_7230,N_7072);
nor U7260 (N_7260,N_7005,N_7202);
and U7261 (N_7261,N_7029,N_7026);
xor U7262 (N_7262,N_7104,N_7142);
xnor U7263 (N_7263,N_7210,N_7245);
nor U7264 (N_7264,N_7004,N_7180);
xnor U7265 (N_7265,N_7059,N_7036);
nor U7266 (N_7266,N_7095,N_7074);
and U7267 (N_7267,N_7209,N_7183);
xnor U7268 (N_7268,N_7115,N_7079);
and U7269 (N_7269,N_7047,N_7108);
xor U7270 (N_7270,N_7052,N_7081);
or U7271 (N_7271,N_7088,N_7194);
nand U7272 (N_7272,N_7000,N_7168);
or U7273 (N_7273,N_7053,N_7109);
and U7274 (N_7274,N_7188,N_7126);
nor U7275 (N_7275,N_7143,N_7178);
or U7276 (N_7276,N_7101,N_7227);
or U7277 (N_7277,N_7239,N_7224);
nor U7278 (N_7278,N_7169,N_7097);
or U7279 (N_7279,N_7119,N_7164);
xnor U7280 (N_7280,N_7181,N_7165);
xor U7281 (N_7281,N_7204,N_7135);
nand U7282 (N_7282,N_7128,N_7046);
nor U7283 (N_7283,N_7054,N_7175);
or U7284 (N_7284,N_7069,N_7035);
and U7285 (N_7285,N_7151,N_7201);
and U7286 (N_7286,N_7091,N_7080);
or U7287 (N_7287,N_7191,N_7131);
and U7288 (N_7288,N_7056,N_7040);
and U7289 (N_7289,N_7130,N_7243);
xor U7290 (N_7290,N_7099,N_7211);
nand U7291 (N_7291,N_7187,N_7015);
nand U7292 (N_7292,N_7002,N_7145);
xnor U7293 (N_7293,N_7103,N_7177);
or U7294 (N_7294,N_7122,N_7231);
xnor U7295 (N_7295,N_7228,N_7112);
nor U7296 (N_7296,N_7203,N_7063);
and U7297 (N_7297,N_7123,N_7086);
or U7298 (N_7298,N_7102,N_7010);
xor U7299 (N_7299,N_7066,N_7033);
and U7300 (N_7300,N_7197,N_7229);
or U7301 (N_7301,N_7248,N_7235);
xnor U7302 (N_7302,N_7120,N_7226);
nor U7303 (N_7303,N_7106,N_7043);
nand U7304 (N_7304,N_7208,N_7022);
xnor U7305 (N_7305,N_7207,N_7223);
nor U7306 (N_7306,N_7077,N_7111);
and U7307 (N_7307,N_7214,N_7013);
or U7308 (N_7308,N_7113,N_7138);
and U7309 (N_7309,N_7057,N_7121);
xnor U7310 (N_7310,N_7070,N_7075);
or U7311 (N_7311,N_7117,N_7009);
nand U7312 (N_7312,N_7141,N_7156);
xor U7313 (N_7313,N_7242,N_7105);
xnor U7314 (N_7314,N_7246,N_7039);
nand U7315 (N_7315,N_7144,N_7100);
xnor U7316 (N_7316,N_7003,N_7071);
xnor U7317 (N_7317,N_7132,N_7060);
or U7318 (N_7318,N_7024,N_7020);
nand U7319 (N_7319,N_7233,N_7032);
nor U7320 (N_7320,N_7068,N_7176);
nor U7321 (N_7321,N_7152,N_7195);
and U7322 (N_7322,N_7082,N_7084);
or U7323 (N_7323,N_7041,N_7236);
xnor U7324 (N_7324,N_7206,N_7014);
xor U7325 (N_7325,N_7192,N_7205);
nand U7326 (N_7326,N_7037,N_7237);
xor U7327 (N_7327,N_7167,N_7007);
xor U7328 (N_7328,N_7027,N_7172);
or U7329 (N_7329,N_7221,N_7137);
xnor U7330 (N_7330,N_7018,N_7185);
nor U7331 (N_7331,N_7073,N_7162);
nand U7332 (N_7332,N_7008,N_7218);
and U7333 (N_7333,N_7133,N_7124);
nor U7334 (N_7334,N_7189,N_7220);
nand U7335 (N_7335,N_7170,N_7179);
or U7336 (N_7336,N_7136,N_7062);
nand U7337 (N_7337,N_7050,N_7051);
or U7338 (N_7338,N_7148,N_7098);
and U7339 (N_7339,N_7198,N_7078);
or U7340 (N_7340,N_7200,N_7017);
nor U7341 (N_7341,N_7038,N_7067);
nand U7342 (N_7342,N_7092,N_7030);
and U7343 (N_7343,N_7161,N_7215);
or U7344 (N_7344,N_7249,N_7149);
and U7345 (N_7345,N_7016,N_7107);
or U7346 (N_7346,N_7001,N_7193);
nand U7347 (N_7347,N_7150,N_7147);
and U7348 (N_7348,N_7093,N_7058);
or U7349 (N_7349,N_7241,N_7222);
nor U7350 (N_7350,N_7089,N_7114);
nand U7351 (N_7351,N_7234,N_7213);
nor U7352 (N_7352,N_7116,N_7154);
or U7353 (N_7353,N_7064,N_7157);
xor U7354 (N_7354,N_7184,N_7083);
or U7355 (N_7355,N_7021,N_7166);
nand U7356 (N_7356,N_7127,N_7090);
nor U7357 (N_7357,N_7140,N_7134);
xnor U7358 (N_7358,N_7044,N_7247);
xor U7359 (N_7359,N_7076,N_7055);
xnor U7360 (N_7360,N_7129,N_7238);
and U7361 (N_7361,N_7216,N_7186);
nor U7362 (N_7362,N_7196,N_7045);
and U7363 (N_7363,N_7219,N_7012);
nand U7364 (N_7364,N_7159,N_7006);
xor U7365 (N_7365,N_7025,N_7232);
or U7366 (N_7366,N_7061,N_7155);
or U7367 (N_7367,N_7049,N_7217);
and U7368 (N_7368,N_7094,N_7096);
nand U7369 (N_7369,N_7244,N_7118);
nand U7370 (N_7370,N_7034,N_7048);
nand U7371 (N_7371,N_7139,N_7199);
or U7372 (N_7372,N_7182,N_7087);
nand U7373 (N_7373,N_7174,N_7240);
xor U7374 (N_7374,N_7065,N_7171);
nand U7375 (N_7375,N_7021,N_7188);
xor U7376 (N_7376,N_7194,N_7167);
xor U7377 (N_7377,N_7092,N_7127);
nor U7378 (N_7378,N_7112,N_7160);
nor U7379 (N_7379,N_7240,N_7188);
xnor U7380 (N_7380,N_7082,N_7192);
or U7381 (N_7381,N_7141,N_7079);
xnor U7382 (N_7382,N_7052,N_7158);
nor U7383 (N_7383,N_7136,N_7202);
and U7384 (N_7384,N_7148,N_7149);
xnor U7385 (N_7385,N_7122,N_7133);
and U7386 (N_7386,N_7221,N_7145);
nor U7387 (N_7387,N_7110,N_7167);
nor U7388 (N_7388,N_7118,N_7246);
xor U7389 (N_7389,N_7069,N_7029);
nand U7390 (N_7390,N_7151,N_7239);
nor U7391 (N_7391,N_7175,N_7060);
or U7392 (N_7392,N_7158,N_7151);
nor U7393 (N_7393,N_7163,N_7159);
xnor U7394 (N_7394,N_7136,N_7058);
nor U7395 (N_7395,N_7095,N_7130);
or U7396 (N_7396,N_7104,N_7190);
or U7397 (N_7397,N_7171,N_7099);
or U7398 (N_7398,N_7233,N_7248);
nor U7399 (N_7399,N_7153,N_7187);
nor U7400 (N_7400,N_7191,N_7174);
nor U7401 (N_7401,N_7231,N_7228);
xnor U7402 (N_7402,N_7000,N_7107);
and U7403 (N_7403,N_7049,N_7199);
and U7404 (N_7404,N_7129,N_7011);
nand U7405 (N_7405,N_7085,N_7098);
and U7406 (N_7406,N_7153,N_7133);
nor U7407 (N_7407,N_7218,N_7042);
nand U7408 (N_7408,N_7084,N_7034);
nand U7409 (N_7409,N_7217,N_7170);
or U7410 (N_7410,N_7113,N_7070);
nand U7411 (N_7411,N_7113,N_7034);
nor U7412 (N_7412,N_7177,N_7176);
nand U7413 (N_7413,N_7027,N_7077);
xnor U7414 (N_7414,N_7051,N_7198);
and U7415 (N_7415,N_7229,N_7224);
xor U7416 (N_7416,N_7199,N_7064);
and U7417 (N_7417,N_7136,N_7047);
nor U7418 (N_7418,N_7064,N_7059);
nand U7419 (N_7419,N_7195,N_7122);
and U7420 (N_7420,N_7238,N_7157);
nand U7421 (N_7421,N_7236,N_7046);
or U7422 (N_7422,N_7223,N_7225);
xnor U7423 (N_7423,N_7164,N_7129);
and U7424 (N_7424,N_7189,N_7232);
nor U7425 (N_7425,N_7087,N_7051);
xnor U7426 (N_7426,N_7086,N_7102);
or U7427 (N_7427,N_7171,N_7105);
and U7428 (N_7428,N_7186,N_7159);
or U7429 (N_7429,N_7145,N_7118);
and U7430 (N_7430,N_7051,N_7249);
or U7431 (N_7431,N_7234,N_7151);
nor U7432 (N_7432,N_7072,N_7079);
nand U7433 (N_7433,N_7127,N_7183);
or U7434 (N_7434,N_7041,N_7162);
xor U7435 (N_7435,N_7186,N_7228);
xnor U7436 (N_7436,N_7165,N_7076);
or U7437 (N_7437,N_7006,N_7146);
xnor U7438 (N_7438,N_7176,N_7118);
xnor U7439 (N_7439,N_7012,N_7024);
nand U7440 (N_7440,N_7092,N_7124);
or U7441 (N_7441,N_7045,N_7147);
or U7442 (N_7442,N_7039,N_7078);
nand U7443 (N_7443,N_7049,N_7117);
xor U7444 (N_7444,N_7050,N_7110);
nor U7445 (N_7445,N_7168,N_7169);
nor U7446 (N_7446,N_7196,N_7158);
or U7447 (N_7447,N_7210,N_7244);
and U7448 (N_7448,N_7047,N_7035);
nor U7449 (N_7449,N_7054,N_7111);
xnor U7450 (N_7450,N_7112,N_7185);
nand U7451 (N_7451,N_7028,N_7005);
nand U7452 (N_7452,N_7035,N_7008);
xor U7453 (N_7453,N_7213,N_7027);
nand U7454 (N_7454,N_7030,N_7191);
xor U7455 (N_7455,N_7192,N_7167);
nand U7456 (N_7456,N_7096,N_7157);
nand U7457 (N_7457,N_7149,N_7207);
or U7458 (N_7458,N_7098,N_7150);
xnor U7459 (N_7459,N_7007,N_7218);
and U7460 (N_7460,N_7174,N_7248);
nand U7461 (N_7461,N_7005,N_7088);
xnor U7462 (N_7462,N_7186,N_7122);
and U7463 (N_7463,N_7192,N_7097);
or U7464 (N_7464,N_7162,N_7168);
nand U7465 (N_7465,N_7203,N_7236);
nor U7466 (N_7466,N_7193,N_7158);
nand U7467 (N_7467,N_7162,N_7167);
xor U7468 (N_7468,N_7055,N_7105);
nor U7469 (N_7469,N_7196,N_7185);
nor U7470 (N_7470,N_7185,N_7059);
nor U7471 (N_7471,N_7058,N_7170);
xor U7472 (N_7472,N_7242,N_7211);
nor U7473 (N_7473,N_7206,N_7221);
or U7474 (N_7474,N_7085,N_7246);
xor U7475 (N_7475,N_7025,N_7175);
and U7476 (N_7476,N_7084,N_7119);
or U7477 (N_7477,N_7077,N_7154);
nor U7478 (N_7478,N_7099,N_7208);
xor U7479 (N_7479,N_7002,N_7160);
nand U7480 (N_7480,N_7158,N_7060);
nor U7481 (N_7481,N_7140,N_7235);
xnor U7482 (N_7482,N_7216,N_7239);
nand U7483 (N_7483,N_7217,N_7056);
nor U7484 (N_7484,N_7138,N_7054);
nand U7485 (N_7485,N_7193,N_7012);
nand U7486 (N_7486,N_7190,N_7103);
or U7487 (N_7487,N_7210,N_7067);
and U7488 (N_7488,N_7009,N_7164);
nor U7489 (N_7489,N_7054,N_7062);
nor U7490 (N_7490,N_7039,N_7047);
xor U7491 (N_7491,N_7121,N_7056);
or U7492 (N_7492,N_7240,N_7040);
nor U7493 (N_7493,N_7124,N_7042);
nand U7494 (N_7494,N_7206,N_7195);
nand U7495 (N_7495,N_7075,N_7094);
or U7496 (N_7496,N_7012,N_7111);
xor U7497 (N_7497,N_7108,N_7137);
nor U7498 (N_7498,N_7232,N_7134);
xnor U7499 (N_7499,N_7050,N_7236);
nand U7500 (N_7500,N_7323,N_7448);
or U7501 (N_7501,N_7281,N_7381);
nand U7502 (N_7502,N_7359,N_7445);
xor U7503 (N_7503,N_7416,N_7284);
or U7504 (N_7504,N_7317,N_7333);
nor U7505 (N_7505,N_7392,N_7278);
nor U7506 (N_7506,N_7482,N_7374);
or U7507 (N_7507,N_7465,N_7340);
nand U7508 (N_7508,N_7300,N_7262);
xor U7509 (N_7509,N_7270,N_7382);
or U7510 (N_7510,N_7490,N_7437);
and U7511 (N_7511,N_7475,N_7439);
nor U7512 (N_7512,N_7354,N_7388);
nor U7513 (N_7513,N_7295,N_7302);
nor U7514 (N_7514,N_7287,N_7318);
and U7515 (N_7515,N_7307,N_7251);
nand U7516 (N_7516,N_7476,N_7413);
or U7517 (N_7517,N_7479,N_7393);
xnor U7518 (N_7518,N_7467,N_7419);
xnor U7519 (N_7519,N_7297,N_7498);
nand U7520 (N_7520,N_7310,N_7320);
and U7521 (N_7521,N_7435,N_7442);
nor U7522 (N_7522,N_7337,N_7463);
nor U7523 (N_7523,N_7377,N_7254);
xnor U7524 (N_7524,N_7384,N_7412);
or U7525 (N_7525,N_7368,N_7394);
and U7526 (N_7526,N_7361,N_7369);
or U7527 (N_7527,N_7461,N_7426);
and U7528 (N_7528,N_7325,N_7378);
and U7529 (N_7529,N_7473,N_7275);
nand U7530 (N_7530,N_7294,N_7343);
nand U7531 (N_7531,N_7492,N_7316);
or U7532 (N_7532,N_7370,N_7304);
and U7533 (N_7533,N_7446,N_7334);
and U7534 (N_7534,N_7298,N_7272);
and U7535 (N_7535,N_7288,N_7391);
xor U7536 (N_7536,N_7415,N_7466);
nor U7537 (N_7537,N_7422,N_7495);
and U7538 (N_7538,N_7265,N_7366);
nor U7539 (N_7539,N_7268,N_7313);
nor U7540 (N_7540,N_7328,N_7273);
nor U7541 (N_7541,N_7408,N_7371);
or U7542 (N_7542,N_7331,N_7289);
or U7543 (N_7543,N_7380,N_7450);
nor U7544 (N_7544,N_7303,N_7497);
nand U7545 (N_7545,N_7383,N_7329);
xor U7546 (N_7546,N_7430,N_7395);
or U7547 (N_7547,N_7271,N_7396);
nand U7548 (N_7548,N_7356,N_7459);
nor U7549 (N_7549,N_7363,N_7264);
nand U7550 (N_7550,N_7259,N_7364);
and U7551 (N_7551,N_7314,N_7403);
or U7552 (N_7552,N_7376,N_7496);
nor U7553 (N_7553,N_7420,N_7398);
or U7554 (N_7554,N_7493,N_7326);
nand U7555 (N_7555,N_7260,N_7404);
xor U7556 (N_7556,N_7283,N_7353);
nand U7557 (N_7557,N_7425,N_7282);
and U7558 (N_7558,N_7432,N_7362);
or U7559 (N_7559,N_7311,N_7332);
nor U7560 (N_7560,N_7464,N_7436);
nor U7561 (N_7561,N_7296,N_7458);
xor U7562 (N_7562,N_7279,N_7274);
and U7563 (N_7563,N_7453,N_7256);
and U7564 (N_7564,N_7253,N_7276);
and U7565 (N_7565,N_7489,N_7421);
or U7566 (N_7566,N_7306,N_7335);
xor U7567 (N_7567,N_7385,N_7389);
nor U7568 (N_7568,N_7454,N_7358);
nand U7569 (N_7569,N_7327,N_7299);
or U7570 (N_7570,N_7485,N_7372);
nand U7571 (N_7571,N_7417,N_7348);
xnor U7572 (N_7572,N_7427,N_7250);
nor U7573 (N_7573,N_7347,N_7301);
nand U7574 (N_7574,N_7373,N_7367);
xor U7575 (N_7575,N_7305,N_7434);
or U7576 (N_7576,N_7257,N_7474);
or U7577 (N_7577,N_7488,N_7407);
nand U7578 (N_7578,N_7471,N_7267);
xnor U7579 (N_7579,N_7266,N_7263);
or U7580 (N_7580,N_7286,N_7338);
or U7581 (N_7581,N_7410,N_7478);
and U7582 (N_7582,N_7440,N_7285);
and U7583 (N_7583,N_7441,N_7357);
and U7584 (N_7584,N_7345,N_7428);
xnor U7585 (N_7585,N_7386,N_7405);
nand U7586 (N_7586,N_7312,N_7477);
nor U7587 (N_7587,N_7423,N_7486);
or U7588 (N_7588,N_7433,N_7292);
xor U7589 (N_7589,N_7402,N_7469);
nor U7590 (N_7590,N_7290,N_7462);
xor U7591 (N_7591,N_7349,N_7470);
nor U7592 (N_7592,N_7344,N_7293);
nor U7593 (N_7593,N_7411,N_7447);
nor U7594 (N_7594,N_7261,N_7255);
or U7595 (N_7595,N_7499,N_7319);
or U7596 (N_7596,N_7258,N_7438);
xor U7597 (N_7597,N_7429,N_7444);
or U7598 (N_7598,N_7321,N_7365);
nand U7599 (N_7599,N_7387,N_7456);
xor U7600 (N_7600,N_7280,N_7457);
or U7601 (N_7601,N_7355,N_7487);
nand U7602 (N_7602,N_7390,N_7401);
nand U7603 (N_7603,N_7397,N_7460);
or U7604 (N_7604,N_7481,N_7269);
xor U7605 (N_7605,N_7342,N_7379);
xnor U7606 (N_7606,N_7350,N_7443);
nor U7607 (N_7607,N_7418,N_7360);
nor U7608 (N_7608,N_7336,N_7483);
or U7609 (N_7609,N_7309,N_7330);
and U7610 (N_7610,N_7322,N_7494);
and U7611 (N_7611,N_7424,N_7277);
xnor U7612 (N_7612,N_7455,N_7291);
xor U7613 (N_7613,N_7472,N_7324);
or U7614 (N_7614,N_7341,N_7431);
or U7615 (N_7615,N_7484,N_7452);
xor U7616 (N_7616,N_7414,N_7451);
or U7617 (N_7617,N_7315,N_7468);
or U7618 (N_7618,N_7375,N_7409);
nor U7619 (N_7619,N_7308,N_7406);
xor U7620 (N_7620,N_7339,N_7252);
or U7621 (N_7621,N_7480,N_7449);
nor U7622 (N_7622,N_7352,N_7399);
nor U7623 (N_7623,N_7400,N_7491);
xor U7624 (N_7624,N_7351,N_7346);
nor U7625 (N_7625,N_7472,N_7312);
nor U7626 (N_7626,N_7418,N_7410);
nor U7627 (N_7627,N_7293,N_7250);
nor U7628 (N_7628,N_7266,N_7451);
nand U7629 (N_7629,N_7481,N_7372);
and U7630 (N_7630,N_7417,N_7266);
or U7631 (N_7631,N_7381,N_7319);
and U7632 (N_7632,N_7313,N_7423);
nor U7633 (N_7633,N_7363,N_7494);
and U7634 (N_7634,N_7409,N_7301);
nor U7635 (N_7635,N_7321,N_7460);
or U7636 (N_7636,N_7387,N_7410);
xnor U7637 (N_7637,N_7442,N_7390);
nor U7638 (N_7638,N_7360,N_7287);
xnor U7639 (N_7639,N_7472,N_7416);
nand U7640 (N_7640,N_7423,N_7288);
and U7641 (N_7641,N_7341,N_7421);
nand U7642 (N_7642,N_7475,N_7410);
nor U7643 (N_7643,N_7256,N_7450);
or U7644 (N_7644,N_7253,N_7446);
nand U7645 (N_7645,N_7403,N_7454);
and U7646 (N_7646,N_7476,N_7409);
nand U7647 (N_7647,N_7358,N_7384);
or U7648 (N_7648,N_7410,N_7305);
nor U7649 (N_7649,N_7262,N_7307);
nor U7650 (N_7650,N_7395,N_7467);
and U7651 (N_7651,N_7280,N_7353);
nor U7652 (N_7652,N_7269,N_7403);
nor U7653 (N_7653,N_7486,N_7418);
and U7654 (N_7654,N_7340,N_7484);
nor U7655 (N_7655,N_7403,N_7417);
nand U7656 (N_7656,N_7386,N_7316);
or U7657 (N_7657,N_7378,N_7340);
or U7658 (N_7658,N_7445,N_7340);
or U7659 (N_7659,N_7353,N_7378);
and U7660 (N_7660,N_7337,N_7382);
xnor U7661 (N_7661,N_7406,N_7478);
or U7662 (N_7662,N_7435,N_7461);
or U7663 (N_7663,N_7330,N_7264);
or U7664 (N_7664,N_7365,N_7470);
or U7665 (N_7665,N_7386,N_7499);
nand U7666 (N_7666,N_7496,N_7444);
or U7667 (N_7667,N_7473,N_7321);
and U7668 (N_7668,N_7265,N_7394);
nor U7669 (N_7669,N_7267,N_7343);
nor U7670 (N_7670,N_7418,N_7308);
or U7671 (N_7671,N_7361,N_7484);
and U7672 (N_7672,N_7340,N_7284);
nand U7673 (N_7673,N_7321,N_7296);
xor U7674 (N_7674,N_7322,N_7263);
nand U7675 (N_7675,N_7406,N_7294);
and U7676 (N_7676,N_7426,N_7463);
nand U7677 (N_7677,N_7289,N_7464);
and U7678 (N_7678,N_7383,N_7389);
xnor U7679 (N_7679,N_7475,N_7445);
or U7680 (N_7680,N_7487,N_7257);
and U7681 (N_7681,N_7480,N_7440);
or U7682 (N_7682,N_7269,N_7300);
nor U7683 (N_7683,N_7439,N_7461);
nor U7684 (N_7684,N_7477,N_7393);
nor U7685 (N_7685,N_7391,N_7350);
xor U7686 (N_7686,N_7369,N_7419);
or U7687 (N_7687,N_7493,N_7347);
xnor U7688 (N_7688,N_7487,N_7395);
nand U7689 (N_7689,N_7403,N_7296);
nor U7690 (N_7690,N_7317,N_7338);
and U7691 (N_7691,N_7498,N_7467);
and U7692 (N_7692,N_7415,N_7444);
xnor U7693 (N_7693,N_7429,N_7318);
or U7694 (N_7694,N_7384,N_7392);
nand U7695 (N_7695,N_7353,N_7335);
nand U7696 (N_7696,N_7450,N_7302);
xor U7697 (N_7697,N_7465,N_7413);
xnor U7698 (N_7698,N_7279,N_7255);
xnor U7699 (N_7699,N_7275,N_7436);
or U7700 (N_7700,N_7476,N_7408);
or U7701 (N_7701,N_7335,N_7439);
or U7702 (N_7702,N_7460,N_7370);
xnor U7703 (N_7703,N_7466,N_7305);
or U7704 (N_7704,N_7271,N_7472);
nor U7705 (N_7705,N_7325,N_7496);
xnor U7706 (N_7706,N_7277,N_7497);
xnor U7707 (N_7707,N_7363,N_7339);
or U7708 (N_7708,N_7454,N_7434);
xor U7709 (N_7709,N_7396,N_7490);
nand U7710 (N_7710,N_7359,N_7398);
nand U7711 (N_7711,N_7301,N_7401);
nor U7712 (N_7712,N_7252,N_7288);
nor U7713 (N_7713,N_7318,N_7373);
or U7714 (N_7714,N_7470,N_7485);
nand U7715 (N_7715,N_7370,N_7468);
and U7716 (N_7716,N_7472,N_7415);
and U7717 (N_7717,N_7300,N_7302);
nand U7718 (N_7718,N_7422,N_7413);
and U7719 (N_7719,N_7370,N_7303);
nor U7720 (N_7720,N_7437,N_7441);
and U7721 (N_7721,N_7288,N_7474);
xnor U7722 (N_7722,N_7382,N_7277);
and U7723 (N_7723,N_7388,N_7435);
xor U7724 (N_7724,N_7259,N_7288);
nor U7725 (N_7725,N_7281,N_7461);
or U7726 (N_7726,N_7422,N_7305);
nor U7727 (N_7727,N_7278,N_7280);
xnor U7728 (N_7728,N_7442,N_7413);
and U7729 (N_7729,N_7313,N_7294);
and U7730 (N_7730,N_7261,N_7456);
and U7731 (N_7731,N_7254,N_7275);
nand U7732 (N_7732,N_7399,N_7423);
and U7733 (N_7733,N_7419,N_7425);
and U7734 (N_7734,N_7495,N_7427);
nand U7735 (N_7735,N_7267,N_7319);
and U7736 (N_7736,N_7369,N_7323);
nor U7737 (N_7737,N_7434,N_7457);
nand U7738 (N_7738,N_7277,N_7489);
xnor U7739 (N_7739,N_7311,N_7323);
or U7740 (N_7740,N_7283,N_7306);
xnor U7741 (N_7741,N_7469,N_7480);
xnor U7742 (N_7742,N_7391,N_7333);
xor U7743 (N_7743,N_7282,N_7407);
nor U7744 (N_7744,N_7491,N_7479);
or U7745 (N_7745,N_7476,N_7335);
and U7746 (N_7746,N_7476,N_7435);
nor U7747 (N_7747,N_7309,N_7448);
xnor U7748 (N_7748,N_7351,N_7362);
nor U7749 (N_7749,N_7288,N_7406);
nor U7750 (N_7750,N_7600,N_7535);
and U7751 (N_7751,N_7520,N_7567);
and U7752 (N_7752,N_7516,N_7598);
and U7753 (N_7753,N_7710,N_7503);
nand U7754 (N_7754,N_7713,N_7500);
nand U7755 (N_7755,N_7612,N_7748);
and U7756 (N_7756,N_7607,N_7708);
or U7757 (N_7757,N_7678,N_7568);
nand U7758 (N_7758,N_7539,N_7694);
xnor U7759 (N_7759,N_7665,N_7709);
nor U7760 (N_7760,N_7714,N_7613);
nand U7761 (N_7761,N_7614,N_7590);
nor U7762 (N_7762,N_7589,N_7533);
nand U7763 (N_7763,N_7625,N_7513);
or U7764 (N_7764,N_7749,N_7517);
nor U7765 (N_7765,N_7674,N_7543);
nand U7766 (N_7766,N_7574,N_7644);
nand U7767 (N_7767,N_7556,N_7615);
and U7768 (N_7768,N_7702,N_7744);
nand U7769 (N_7769,N_7681,N_7599);
or U7770 (N_7770,N_7652,N_7634);
xnor U7771 (N_7771,N_7668,N_7645);
nor U7772 (N_7772,N_7696,N_7701);
nor U7773 (N_7773,N_7659,N_7584);
nand U7774 (N_7774,N_7742,N_7730);
nand U7775 (N_7775,N_7686,N_7655);
xnor U7776 (N_7776,N_7711,N_7571);
and U7777 (N_7777,N_7538,N_7546);
nand U7778 (N_7778,N_7586,N_7580);
or U7779 (N_7779,N_7728,N_7509);
and U7780 (N_7780,N_7675,N_7627);
and U7781 (N_7781,N_7527,N_7582);
xor U7782 (N_7782,N_7657,N_7530);
nor U7783 (N_7783,N_7667,N_7680);
and U7784 (N_7784,N_7604,N_7606);
and U7785 (N_7785,N_7723,N_7510);
or U7786 (N_7786,N_7691,N_7725);
xnor U7787 (N_7787,N_7676,N_7561);
xor U7788 (N_7788,N_7554,N_7529);
or U7789 (N_7789,N_7724,N_7643);
xor U7790 (N_7790,N_7630,N_7650);
xor U7791 (N_7791,N_7553,N_7649);
or U7792 (N_7792,N_7640,N_7642);
and U7793 (N_7793,N_7578,N_7617);
nand U7794 (N_7794,N_7564,N_7536);
xnor U7795 (N_7795,N_7526,N_7658);
and U7796 (N_7796,N_7569,N_7514);
nor U7797 (N_7797,N_7523,N_7718);
xor U7798 (N_7798,N_7560,N_7693);
xnor U7799 (N_7799,N_7706,N_7544);
and U7800 (N_7800,N_7712,N_7648);
and U7801 (N_7801,N_7684,N_7591);
and U7802 (N_7802,N_7559,N_7651);
or U7803 (N_7803,N_7747,N_7647);
nand U7804 (N_7804,N_7522,N_7532);
nor U7805 (N_7805,N_7682,N_7661);
xnor U7806 (N_7806,N_7610,N_7666);
nand U7807 (N_7807,N_7733,N_7566);
nand U7808 (N_7808,N_7623,N_7621);
nor U7809 (N_7809,N_7572,N_7729);
or U7810 (N_7810,N_7528,N_7739);
and U7811 (N_7811,N_7700,N_7732);
xor U7812 (N_7812,N_7511,N_7707);
and U7813 (N_7813,N_7631,N_7746);
xor U7814 (N_7814,N_7552,N_7542);
and U7815 (N_7815,N_7641,N_7705);
nand U7816 (N_7816,N_7620,N_7638);
nand U7817 (N_7817,N_7534,N_7558);
or U7818 (N_7818,N_7646,N_7562);
or U7819 (N_7819,N_7577,N_7601);
or U7820 (N_7820,N_7618,N_7603);
nor U7821 (N_7821,N_7579,N_7632);
and U7822 (N_7822,N_7507,N_7690);
and U7823 (N_7823,N_7619,N_7508);
nor U7824 (N_7824,N_7537,N_7743);
nor U7825 (N_7825,N_7502,N_7721);
or U7826 (N_7826,N_7611,N_7695);
or U7827 (N_7827,N_7518,N_7626);
or U7828 (N_7828,N_7677,N_7519);
and U7829 (N_7829,N_7672,N_7704);
nand U7830 (N_7830,N_7637,N_7673);
and U7831 (N_7831,N_7588,N_7573);
nor U7832 (N_7832,N_7585,N_7524);
nand U7833 (N_7833,N_7740,N_7549);
and U7834 (N_7834,N_7576,N_7551);
or U7835 (N_7835,N_7583,N_7570);
and U7836 (N_7836,N_7587,N_7512);
and U7837 (N_7837,N_7745,N_7656);
nor U7838 (N_7838,N_7506,N_7715);
nor U7839 (N_7839,N_7602,N_7505);
xor U7840 (N_7840,N_7624,N_7545);
and U7841 (N_7841,N_7628,N_7596);
or U7842 (N_7842,N_7679,N_7515);
nor U7843 (N_7843,N_7697,N_7605);
xnor U7844 (N_7844,N_7720,N_7689);
and U7845 (N_7845,N_7670,N_7563);
and U7846 (N_7846,N_7662,N_7734);
xor U7847 (N_7847,N_7504,N_7633);
xor U7848 (N_7848,N_7687,N_7736);
or U7849 (N_7849,N_7699,N_7727);
and U7850 (N_7850,N_7692,N_7575);
nand U7851 (N_7851,N_7629,N_7550);
nor U7852 (N_7852,N_7547,N_7635);
xnor U7853 (N_7853,N_7669,N_7608);
xnor U7854 (N_7854,N_7717,N_7592);
and U7855 (N_7855,N_7521,N_7609);
nor U7856 (N_7856,N_7703,N_7741);
xor U7857 (N_7857,N_7719,N_7663);
nand U7858 (N_7858,N_7636,N_7671);
nor U7859 (N_7859,N_7557,N_7735);
nand U7860 (N_7860,N_7555,N_7716);
xor U7861 (N_7861,N_7595,N_7593);
nor U7862 (N_7862,N_7597,N_7685);
and U7863 (N_7863,N_7548,N_7737);
xor U7864 (N_7864,N_7683,N_7660);
nand U7865 (N_7865,N_7501,N_7731);
and U7866 (N_7866,N_7653,N_7722);
or U7867 (N_7867,N_7540,N_7654);
xnor U7868 (N_7868,N_7565,N_7541);
nor U7869 (N_7869,N_7616,N_7726);
and U7870 (N_7870,N_7622,N_7531);
and U7871 (N_7871,N_7525,N_7664);
and U7872 (N_7872,N_7698,N_7581);
or U7873 (N_7873,N_7688,N_7594);
nor U7874 (N_7874,N_7639,N_7738);
and U7875 (N_7875,N_7526,N_7513);
and U7876 (N_7876,N_7655,N_7515);
xor U7877 (N_7877,N_7670,N_7677);
or U7878 (N_7878,N_7653,N_7683);
or U7879 (N_7879,N_7683,N_7716);
nor U7880 (N_7880,N_7503,N_7555);
nand U7881 (N_7881,N_7661,N_7547);
xnor U7882 (N_7882,N_7660,N_7608);
nand U7883 (N_7883,N_7532,N_7705);
and U7884 (N_7884,N_7566,N_7716);
xnor U7885 (N_7885,N_7687,N_7698);
nand U7886 (N_7886,N_7579,N_7501);
or U7887 (N_7887,N_7708,N_7514);
nor U7888 (N_7888,N_7703,N_7557);
and U7889 (N_7889,N_7605,N_7675);
xor U7890 (N_7890,N_7706,N_7552);
xor U7891 (N_7891,N_7506,N_7559);
xnor U7892 (N_7892,N_7600,N_7633);
nor U7893 (N_7893,N_7566,N_7644);
and U7894 (N_7894,N_7530,N_7579);
and U7895 (N_7895,N_7640,N_7617);
or U7896 (N_7896,N_7568,N_7509);
or U7897 (N_7897,N_7714,N_7554);
nand U7898 (N_7898,N_7693,N_7710);
nand U7899 (N_7899,N_7556,N_7655);
xnor U7900 (N_7900,N_7568,N_7716);
or U7901 (N_7901,N_7669,N_7718);
and U7902 (N_7902,N_7565,N_7665);
nand U7903 (N_7903,N_7606,N_7501);
nand U7904 (N_7904,N_7696,N_7748);
and U7905 (N_7905,N_7711,N_7625);
or U7906 (N_7906,N_7638,N_7674);
or U7907 (N_7907,N_7749,N_7688);
nor U7908 (N_7908,N_7552,N_7616);
or U7909 (N_7909,N_7700,N_7530);
and U7910 (N_7910,N_7715,N_7618);
nor U7911 (N_7911,N_7579,N_7741);
nor U7912 (N_7912,N_7712,N_7500);
nor U7913 (N_7913,N_7619,N_7598);
nor U7914 (N_7914,N_7732,N_7632);
nor U7915 (N_7915,N_7506,N_7684);
and U7916 (N_7916,N_7636,N_7568);
nor U7917 (N_7917,N_7592,N_7638);
nand U7918 (N_7918,N_7638,N_7545);
xor U7919 (N_7919,N_7555,N_7663);
nand U7920 (N_7920,N_7585,N_7697);
and U7921 (N_7921,N_7638,N_7736);
nor U7922 (N_7922,N_7730,N_7735);
and U7923 (N_7923,N_7647,N_7642);
nor U7924 (N_7924,N_7581,N_7542);
and U7925 (N_7925,N_7674,N_7676);
nor U7926 (N_7926,N_7731,N_7730);
nand U7927 (N_7927,N_7510,N_7623);
nand U7928 (N_7928,N_7746,N_7547);
xnor U7929 (N_7929,N_7740,N_7702);
nor U7930 (N_7930,N_7675,N_7528);
and U7931 (N_7931,N_7737,N_7549);
xnor U7932 (N_7932,N_7521,N_7719);
nand U7933 (N_7933,N_7733,N_7721);
and U7934 (N_7934,N_7697,N_7508);
xor U7935 (N_7935,N_7747,N_7506);
nor U7936 (N_7936,N_7602,N_7563);
or U7937 (N_7937,N_7638,N_7737);
nor U7938 (N_7938,N_7550,N_7527);
xor U7939 (N_7939,N_7703,N_7634);
xor U7940 (N_7940,N_7715,N_7531);
or U7941 (N_7941,N_7557,N_7545);
xnor U7942 (N_7942,N_7747,N_7534);
or U7943 (N_7943,N_7718,N_7528);
nand U7944 (N_7944,N_7718,N_7703);
or U7945 (N_7945,N_7544,N_7671);
and U7946 (N_7946,N_7681,N_7627);
or U7947 (N_7947,N_7551,N_7682);
nand U7948 (N_7948,N_7516,N_7608);
nor U7949 (N_7949,N_7564,N_7614);
xor U7950 (N_7950,N_7654,N_7544);
or U7951 (N_7951,N_7665,N_7652);
nor U7952 (N_7952,N_7722,N_7541);
nand U7953 (N_7953,N_7565,N_7509);
or U7954 (N_7954,N_7704,N_7601);
nand U7955 (N_7955,N_7669,N_7605);
nor U7956 (N_7956,N_7522,N_7742);
or U7957 (N_7957,N_7578,N_7575);
or U7958 (N_7958,N_7715,N_7649);
nand U7959 (N_7959,N_7571,N_7689);
and U7960 (N_7960,N_7588,N_7595);
nand U7961 (N_7961,N_7732,N_7748);
nand U7962 (N_7962,N_7691,N_7658);
nor U7963 (N_7963,N_7733,N_7676);
or U7964 (N_7964,N_7705,N_7638);
xor U7965 (N_7965,N_7528,N_7527);
nand U7966 (N_7966,N_7604,N_7698);
nand U7967 (N_7967,N_7500,N_7741);
and U7968 (N_7968,N_7515,N_7620);
nor U7969 (N_7969,N_7705,N_7735);
xor U7970 (N_7970,N_7643,N_7644);
or U7971 (N_7971,N_7508,N_7591);
and U7972 (N_7972,N_7536,N_7643);
nor U7973 (N_7973,N_7533,N_7709);
or U7974 (N_7974,N_7659,N_7608);
and U7975 (N_7975,N_7607,N_7687);
nand U7976 (N_7976,N_7736,N_7545);
nand U7977 (N_7977,N_7564,N_7590);
nor U7978 (N_7978,N_7603,N_7520);
and U7979 (N_7979,N_7584,N_7618);
nand U7980 (N_7980,N_7710,N_7708);
nor U7981 (N_7981,N_7602,N_7567);
xnor U7982 (N_7982,N_7681,N_7699);
or U7983 (N_7983,N_7575,N_7511);
nand U7984 (N_7984,N_7731,N_7736);
nand U7985 (N_7985,N_7550,N_7727);
nor U7986 (N_7986,N_7624,N_7532);
nand U7987 (N_7987,N_7599,N_7526);
or U7988 (N_7988,N_7663,N_7695);
and U7989 (N_7989,N_7654,N_7680);
nand U7990 (N_7990,N_7504,N_7685);
or U7991 (N_7991,N_7706,N_7727);
nand U7992 (N_7992,N_7670,N_7668);
and U7993 (N_7993,N_7656,N_7662);
nand U7994 (N_7994,N_7715,N_7643);
or U7995 (N_7995,N_7697,N_7717);
or U7996 (N_7996,N_7650,N_7507);
nand U7997 (N_7997,N_7708,N_7501);
xor U7998 (N_7998,N_7679,N_7536);
nor U7999 (N_7999,N_7554,N_7682);
or U8000 (N_8000,N_7823,N_7941);
and U8001 (N_8001,N_7841,N_7842);
xnor U8002 (N_8002,N_7825,N_7959);
nor U8003 (N_8003,N_7937,N_7915);
nor U8004 (N_8004,N_7783,N_7866);
nand U8005 (N_8005,N_7900,N_7913);
or U8006 (N_8006,N_7813,N_7805);
nand U8007 (N_8007,N_7831,N_7898);
or U8008 (N_8008,N_7750,N_7756);
xnor U8009 (N_8009,N_7869,N_7821);
and U8010 (N_8010,N_7888,N_7882);
nor U8011 (N_8011,N_7980,N_7987);
or U8012 (N_8012,N_7757,N_7901);
nand U8013 (N_8013,N_7801,N_7972);
nor U8014 (N_8014,N_7799,N_7778);
or U8015 (N_8015,N_7928,N_7846);
nand U8016 (N_8016,N_7909,N_7920);
and U8017 (N_8017,N_7818,N_7874);
nor U8018 (N_8018,N_7808,N_7763);
and U8019 (N_8019,N_7963,N_7964);
xor U8020 (N_8020,N_7923,N_7760);
and U8021 (N_8021,N_7833,N_7766);
nand U8022 (N_8022,N_7781,N_7809);
and U8023 (N_8023,N_7988,N_7970);
nand U8024 (N_8024,N_7896,N_7895);
nand U8025 (N_8025,N_7777,N_7989);
or U8026 (N_8026,N_7932,N_7780);
or U8027 (N_8027,N_7782,N_7857);
or U8028 (N_8028,N_7954,N_7776);
xor U8029 (N_8029,N_7795,N_7877);
or U8030 (N_8030,N_7908,N_7811);
nand U8031 (N_8031,N_7761,N_7971);
and U8032 (N_8032,N_7824,N_7998);
and U8033 (N_8033,N_7802,N_7925);
xnor U8034 (N_8034,N_7765,N_7837);
nor U8035 (N_8035,N_7981,N_7992);
xor U8036 (N_8036,N_7960,N_7976);
or U8037 (N_8037,N_7899,N_7863);
and U8038 (N_8038,N_7804,N_7844);
xnor U8039 (N_8039,N_7800,N_7919);
and U8040 (N_8040,N_7807,N_7843);
nand U8041 (N_8041,N_7878,N_7851);
or U8042 (N_8042,N_7864,N_7940);
nor U8043 (N_8043,N_7885,N_7769);
and U8044 (N_8044,N_7814,N_7754);
xor U8045 (N_8045,N_7906,N_7930);
and U8046 (N_8046,N_7984,N_7789);
xor U8047 (N_8047,N_7770,N_7768);
xnor U8048 (N_8048,N_7839,N_7966);
nor U8049 (N_8049,N_7952,N_7994);
and U8050 (N_8050,N_7829,N_7806);
and U8051 (N_8051,N_7921,N_7929);
xor U8052 (N_8052,N_7907,N_7872);
and U8053 (N_8053,N_7859,N_7995);
nand U8054 (N_8054,N_7944,N_7867);
xor U8055 (N_8055,N_7847,N_7845);
nor U8056 (N_8056,N_7934,N_7978);
or U8057 (N_8057,N_7911,N_7973);
or U8058 (N_8058,N_7986,N_7794);
nor U8059 (N_8059,N_7969,N_7835);
nand U8060 (N_8060,N_7828,N_7751);
nor U8061 (N_8061,N_7817,N_7979);
xor U8062 (N_8062,N_7860,N_7945);
or U8063 (N_8063,N_7965,N_7939);
and U8064 (N_8064,N_7875,N_7893);
xor U8065 (N_8065,N_7894,N_7834);
xor U8066 (N_8066,N_7759,N_7942);
xnor U8067 (N_8067,N_7933,N_7922);
nor U8068 (N_8068,N_7950,N_7957);
nor U8069 (N_8069,N_7916,N_7832);
and U8070 (N_8070,N_7883,N_7822);
or U8071 (N_8071,N_7853,N_7927);
or U8072 (N_8072,N_7924,N_7861);
and U8073 (N_8073,N_7891,N_7996);
xor U8074 (N_8074,N_7938,N_7762);
nor U8075 (N_8075,N_7880,N_7955);
nand U8076 (N_8076,N_7773,N_7786);
nand U8077 (N_8077,N_7926,N_7931);
nand U8078 (N_8078,N_7812,N_7943);
and U8079 (N_8079,N_7870,N_7862);
and U8080 (N_8080,N_7910,N_7764);
nand U8081 (N_8081,N_7949,N_7858);
or U8082 (N_8082,N_7767,N_7962);
and U8083 (N_8083,N_7752,N_7903);
nor U8084 (N_8084,N_7849,N_7784);
nor U8085 (N_8085,N_7999,N_7755);
nor U8086 (N_8086,N_7886,N_7753);
nand U8087 (N_8087,N_7868,N_7826);
xor U8088 (N_8088,N_7793,N_7772);
nand U8089 (N_8089,N_7904,N_7865);
nor U8090 (N_8090,N_7990,N_7889);
and U8091 (N_8091,N_7820,N_7958);
nor U8092 (N_8092,N_7819,N_7947);
nor U8093 (N_8093,N_7897,N_7991);
nor U8094 (N_8094,N_7997,N_7977);
nand U8095 (N_8095,N_7774,N_7758);
or U8096 (N_8096,N_7902,N_7850);
xor U8097 (N_8097,N_7974,N_7840);
nor U8098 (N_8098,N_7797,N_7836);
or U8099 (N_8099,N_7790,N_7838);
xnor U8100 (N_8100,N_7953,N_7935);
or U8101 (N_8101,N_7787,N_7982);
or U8102 (N_8102,N_7914,N_7879);
nand U8103 (N_8103,N_7803,N_7855);
or U8104 (N_8104,N_7873,N_7775);
and U8105 (N_8105,N_7948,N_7961);
xnor U8106 (N_8106,N_7798,N_7785);
xnor U8107 (N_8107,N_7968,N_7884);
nand U8108 (N_8108,N_7771,N_7912);
nand U8109 (N_8109,N_7946,N_7993);
and U8110 (N_8110,N_7983,N_7876);
xor U8111 (N_8111,N_7810,N_7936);
xnor U8112 (N_8112,N_7852,N_7985);
xor U8113 (N_8113,N_7975,N_7856);
nor U8114 (N_8114,N_7815,N_7788);
or U8115 (N_8115,N_7881,N_7871);
or U8116 (N_8116,N_7917,N_7892);
nor U8117 (N_8117,N_7830,N_7796);
xnor U8118 (N_8118,N_7779,N_7792);
and U8119 (N_8119,N_7918,N_7890);
nand U8120 (N_8120,N_7967,N_7956);
or U8121 (N_8121,N_7905,N_7951);
or U8122 (N_8122,N_7848,N_7816);
or U8123 (N_8123,N_7887,N_7827);
nand U8124 (N_8124,N_7791,N_7854);
nor U8125 (N_8125,N_7766,N_7755);
xnor U8126 (N_8126,N_7908,N_7870);
nor U8127 (N_8127,N_7753,N_7907);
and U8128 (N_8128,N_7789,N_7931);
xnor U8129 (N_8129,N_7873,N_7790);
nand U8130 (N_8130,N_7919,N_7918);
xor U8131 (N_8131,N_7972,N_7995);
and U8132 (N_8132,N_7850,N_7761);
nor U8133 (N_8133,N_7790,N_7783);
xor U8134 (N_8134,N_7763,N_7995);
nor U8135 (N_8135,N_7864,N_7938);
xnor U8136 (N_8136,N_7938,N_7870);
or U8137 (N_8137,N_7761,N_7987);
nor U8138 (N_8138,N_7863,N_7841);
nor U8139 (N_8139,N_7936,N_7791);
nor U8140 (N_8140,N_7920,N_7936);
and U8141 (N_8141,N_7923,N_7964);
and U8142 (N_8142,N_7997,N_7911);
xnor U8143 (N_8143,N_7784,N_7787);
or U8144 (N_8144,N_7972,N_7784);
or U8145 (N_8145,N_7905,N_7844);
and U8146 (N_8146,N_7861,N_7811);
or U8147 (N_8147,N_7757,N_7887);
and U8148 (N_8148,N_7778,N_7995);
nand U8149 (N_8149,N_7760,N_7838);
xor U8150 (N_8150,N_7882,N_7827);
and U8151 (N_8151,N_7880,N_7841);
nor U8152 (N_8152,N_7954,N_7947);
and U8153 (N_8153,N_7939,N_7798);
nor U8154 (N_8154,N_7822,N_7870);
or U8155 (N_8155,N_7816,N_7786);
xor U8156 (N_8156,N_7768,N_7802);
xor U8157 (N_8157,N_7777,N_7792);
xnor U8158 (N_8158,N_7795,N_7957);
xnor U8159 (N_8159,N_7983,N_7766);
and U8160 (N_8160,N_7853,N_7919);
nand U8161 (N_8161,N_7836,N_7915);
xnor U8162 (N_8162,N_7828,N_7851);
nor U8163 (N_8163,N_7889,N_7802);
nor U8164 (N_8164,N_7858,N_7923);
or U8165 (N_8165,N_7906,N_7807);
and U8166 (N_8166,N_7969,N_7852);
xnor U8167 (N_8167,N_7757,N_7750);
nand U8168 (N_8168,N_7896,N_7974);
nand U8169 (N_8169,N_7780,N_7950);
or U8170 (N_8170,N_7903,N_7889);
and U8171 (N_8171,N_7893,N_7766);
nand U8172 (N_8172,N_7952,N_7948);
nor U8173 (N_8173,N_7898,N_7971);
xnor U8174 (N_8174,N_7764,N_7882);
xnor U8175 (N_8175,N_7844,N_7797);
or U8176 (N_8176,N_7961,N_7864);
xor U8177 (N_8177,N_7780,N_7885);
nand U8178 (N_8178,N_7836,N_7779);
nand U8179 (N_8179,N_7954,N_7857);
nand U8180 (N_8180,N_7979,N_7953);
or U8181 (N_8181,N_7990,N_7959);
nand U8182 (N_8182,N_7777,N_7830);
xnor U8183 (N_8183,N_7877,N_7885);
or U8184 (N_8184,N_7987,N_7774);
and U8185 (N_8185,N_7840,N_7969);
and U8186 (N_8186,N_7754,N_7902);
xor U8187 (N_8187,N_7997,N_7995);
xnor U8188 (N_8188,N_7972,N_7842);
nand U8189 (N_8189,N_7833,N_7855);
nor U8190 (N_8190,N_7937,N_7941);
nor U8191 (N_8191,N_7993,N_7909);
nor U8192 (N_8192,N_7955,N_7900);
xor U8193 (N_8193,N_7940,N_7862);
nand U8194 (N_8194,N_7824,N_7850);
nand U8195 (N_8195,N_7993,N_7855);
nand U8196 (N_8196,N_7883,N_7829);
nor U8197 (N_8197,N_7927,N_7814);
and U8198 (N_8198,N_7769,N_7789);
and U8199 (N_8199,N_7840,N_7821);
nor U8200 (N_8200,N_7870,N_7784);
nand U8201 (N_8201,N_7775,N_7952);
nand U8202 (N_8202,N_7896,N_7767);
nand U8203 (N_8203,N_7875,N_7983);
or U8204 (N_8204,N_7801,N_7894);
xnor U8205 (N_8205,N_7880,N_7911);
nor U8206 (N_8206,N_7812,N_7799);
nand U8207 (N_8207,N_7982,N_7899);
and U8208 (N_8208,N_7852,N_7811);
xor U8209 (N_8209,N_7847,N_7887);
xor U8210 (N_8210,N_7934,N_7756);
nand U8211 (N_8211,N_7917,N_7985);
nor U8212 (N_8212,N_7804,N_7873);
and U8213 (N_8213,N_7877,N_7993);
nand U8214 (N_8214,N_7971,N_7999);
nor U8215 (N_8215,N_7999,N_7883);
or U8216 (N_8216,N_7960,N_7896);
xnor U8217 (N_8217,N_7782,N_7877);
or U8218 (N_8218,N_7850,N_7770);
or U8219 (N_8219,N_7774,N_7868);
xor U8220 (N_8220,N_7889,N_7983);
xnor U8221 (N_8221,N_7825,N_7807);
or U8222 (N_8222,N_7910,N_7757);
or U8223 (N_8223,N_7871,N_7992);
nand U8224 (N_8224,N_7924,N_7833);
nor U8225 (N_8225,N_7753,N_7936);
or U8226 (N_8226,N_7914,N_7856);
nor U8227 (N_8227,N_7921,N_7961);
xor U8228 (N_8228,N_7901,N_7953);
nand U8229 (N_8229,N_7836,N_7946);
nor U8230 (N_8230,N_7887,N_7851);
nand U8231 (N_8231,N_7989,N_7810);
and U8232 (N_8232,N_7818,N_7893);
xor U8233 (N_8233,N_7824,N_7801);
xor U8234 (N_8234,N_7780,N_7978);
xor U8235 (N_8235,N_7825,N_7900);
or U8236 (N_8236,N_7975,N_7986);
nand U8237 (N_8237,N_7769,N_7977);
and U8238 (N_8238,N_7960,N_7920);
or U8239 (N_8239,N_7974,N_7972);
nand U8240 (N_8240,N_7770,N_7760);
or U8241 (N_8241,N_7843,N_7963);
nor U8242 (N_8242,N_7863,N_7950);
and U8243 (N_8243,N_7941,N_7873);
xor U8244 (N_8244,N_7892,N_7882);
xnor U8245 (N_8245,N_7847,N_7901);
nand U8246 (N_8246,N_7816,N_7916);
xor U8247 (N_8247,N_7810,N_7981);
nor U8248 (N_8248,N_7864,N_7773);
or U8249 (N_8249,N_7807,N_7834);
nor U8250 (N_8250,N_8021,N_8211);
or U8251 (N_8251,N_8036,N_8203);
nand U8252 (N_8252,N_8209,N_8137);
and U8253 (N_8253,N_8073,N_8236);
and U8254 (N_8254,N_8007,N_8132);
and U8255 (N_8255,N_8048,N_8078);
nor U8256 (N_8256,N_8076,N_8186);
and U8257 (N_8257,N_8090,N_8049);
nand U8258 (N_8258,N_8027,N_8217);
or U8259 (N_8259,N_8020,N_8115);
nor U8260 (N_8260,N_8063,N_8181);
nor U8261 (N_8261,N_8199,N_8180);
xnor U8262 (N_8262,N_8219,N_8026);
or U8263 (N_8263,N_8127,N_8111);
xor U8264 (N_8264,N_8239,N_8023);
nand U8265 (N_8265,N_8192,N_8099);
nor U8266 (N_8266,N_8013,N_8001);
nand U8267 (N_8267,N_8054,N_8247);
or U8268 (N_8268,N_8113,N_8228);
nand U8269 (N_8269,N_8109,N_8240);
nand U8270 (N_8270,N_8174,N_8101);
xnor U8271 (N_8271,N_8002,N_8167);
xor U8272 (N_8272,N_8053,N_8159);
xor U8273 (N_8273,N_8231,N_8162);
xor U8274 (N_8274,N_8237,N_8194);
xnor U8275 (N_8275,N_8056,N_8197);
xor U8276 (N_8276,N_8178,N_8171);
and U8277 (N_8277,N_8226,N_8069);
nor U8278 (N_8278,N_8123,N_8031);
nor U8279 (N_8279,N_8096,N_8082);
nand U8280 (N_8280,N_8151,N_8080);
xnor U8281 (N_8281,N_8064,N_8147);
nand U8282 (N_8282,N_8223,N_8238);
or U8283 (N_8283,N_8097,N_8037);
and U8284 (N_8284,N_8157,N_8105);
xnor U8285 (N_8285,N_8138,N_8195);
and U8286 (N_8286,N_8177,N_8148);
and U8287 (N_8287,N_8065,N_8163);
nand U8288 (N_8288,N_8179,N_8193);
xnor U8289 (N_8289,N_8019,N_8100);
nor U8290 (N_8290,N_8050,N_8225);
nand U8291 (N_8291,N_8154,N_8224);
or U8292 (N_8292,N_8057,N_8006);
nor U8293 (N_8293,N_8112,N_8214);
nand U8294 (N_8294,N_8246,N_8029);
and U8295 (N_8295,N_8158,N_8213);
nand U8296 (N_8296,N_8117,N_8183);
nor U8297 (N_8297,N_8169,N_8046);
and U8298 (N_8298,N_8206,N_8120);
or U8299 (N_8299,N_8155,N_8009);
and U8300 (N_8300,N_8124,N_8201);
xor U8301 (N_8301,N_8134,N_8204);
xnor U8302 (N_8302,N_8081,N_8133);
or U8303 (N_8303,N_8191,N_8200);
nor U8304 (N_8304,N_8074,N_8220);
or U8305 (N_8305,N_8098,N_8070);
nand U8306 (N_8306,N_8173,N_8085);
and U8307 (N_8307,N_8165,N_8114);
and U8308 (N_8308,N_8005,N_8059);
or U8309 (N_8309,N_8212,N_8035);
xnor U8310 (N_8310,N_8129,N_8189);
nor U8311 (N_8311,N_8218,N_8150);
xor U8312 (N_8312,N_8235,N_8018);
nor U8313 (N_8313,N_8093,N_8043);
or U8314 (N_8314,N_8108,N_8122);
xor U8315 (N_8315,N_8175,N_8116);
xnor U8316 (N_8316,N_8092,N_8041);
and U8317 (N_8317,N_8000,N_8216);
nor U8318 (N_8318,N_8075,N_8079);
or U8319 (N_8319,N_8089,N_8118);
or U8320 (N_8320,N_8103,N_8243);
or U8321 (N_8321,N_8038,N_8003);
nand U8322 (N_8322,N_8095,N_8012);
or U8323 (N_8323,N_8060,N_8010);
or U8324 (N_8324,N_8153,N_8034);
nor U8325 (N_8325,N_8128,N_8051);
or U8326 (N_8326,N_8182,N_8143);
nor U8327 (N_8327,N_8131,N_8024);
and U8328 (N_8328,N_8160,N_8068);
xor U8329 (N_8329,N_8210,N_8135);
nor U8330 (N_8330,N_8110,N_8086);
nand U8331 (N_8331,N_8176,N_8198);
nor U8332 (N_8332,N_8166,N_8229);
nand U8333 (N_8333,N_8126,N_8071);
and U8334 (N_8334,N_8072,N_8011);
nand U8335 (N_8335,N_8106,N_8025);
xor U8336 (N_8336,N_8244,N_8017);
or U8337 (N_8337,N_8205,N_8088);
xor U8338 (N_8338,N_8139,N_8202);
or U8339 (N_8339,N_8145,N_8091);
nor U8340 (N_8340,N_8102,N_8022);
nand U8341 (N_8341,N_8121,N_8187);
nand U8342 (N_8342,N_8125,N_8140);
xor U8343 (N_8343,N_8185,N_8241);
xnor U8344 (N_8344,N_8146,N_8077);
nand U8345 (N_8345,N_8156,N_8084);
nand U8346 (N_8346,N_8230,N_8055);
and U8347 (N_8347,N_8033,N_8149);
and U8348 (N_8348,N_8196,N_8242);
nor U8349 (N_8349,N_8188,N_8014);
and U8350 (N_8350,N_8142,N_8130);
or U8351 (N_8351,N_8058,N_8016);
xnor U8352 (N_8352,N_8215,N_8141);
nor U8353 (N_8353,N_8066,N_8040);
or U8354 (N_8354,N_8104,N_8045);
and U8355 (N_8355,N_8062,N_8168);
nand U8356 (N_8356,N_8249,N_8208);
or U8357 (N_8357,N_8030,N_8136);
or U8358 (N_8358,N_8061,N_8190);
nand U8359 (N_8359,N_8008,N_8044);
nand U8360 (N_8360,N_8047,N_8164);
nand U8361 (N_8361,N_8227,N_8232);
and U8362 (N_8362,N_8233,N_8172);
or U8363 (N_8363,N_8184,N_8245);
nor U8364 (N_8364,N_8119,N_8170);
xor U8365 (N_8365,N_8248,N_8094);
xnor U8366 (N_8366,N_8207,N_8152);
and U8367 (N_8367,N_8083,N_8234);
and U8368 (N_8368,N_8144,N_8032);
nand U8369 (N_8369,N_8052,N_8067);
and U8370 (N_8370,N_8161,N_8015);
xnor U8371 (N_8371,N_8028,N_8004);
or U8372 (N_8372,N_8221,N_8222);
and U8373 (N_8373,N_8039,N_8087);
nor U8374 (N_8374,N_8107,N_8042);
nor U8375 (N_8375,N_8238,N_8240);
nor U8376 (N_8376,N_8187,N_8010);
and U8377 (N_8377,N_8029,N_8244);
xor U8378 (N_8378,N_8056,N_8022);
nor U8379 (N_8379,N_8059,N_8126);
nand U8380 (N_8380,N_8131,N_8092);
and U8381 (N_8381,N_8028,N_8179);
nand U8382 (N_8382,N_8217,N_8091);
nor U8383 (N_8383,N_8222,N_8101);
or U8384 (N_8384,N_8227,N_8082);
or U8385 (N_8385,N_8052,N_8062);
xnor U8386 (N_8386,N_8106,N_8100);
and U8387 (N_8387,N_8015,N_8147);
nor U8388 (N_8388,N_8110,N_8019);
xor U8389 (N_8389,N_8246,N_8048);
nor U8390 (N_8390,N_8031,N_8171);
xor U8391 (N_8391,N_8010,N_8043);
xnor U8392 (N_8392,N_8204,N_8195);
nand U8393 (N_8393,N_8050,N_8005);
and U8394 (N_8394,N_8087,N_8219);
nor U8395 (N_8395,N_8094,N_8081);
nor U8396 (N_8396,N_8051,N_8184);
nor U8397 (N_8397,N_8041,N_8147);
nor U8398 (N_8398,N_8016,N_8040);
and U8399 (N_8399,N_8200,N_8181);
and U8400 (N_8400,N_8044,N_8065);
xnor U8401 (N_8401,N_8150,N_8183);
or U8402 (N_8402,N_8224,N_8038);
or U8403 (N_8403,N_8069,N_8149);
xor U8404 (N_8404,N_8151,N_8139);
nand U8405 (N_8405,N_8082,N_8223);
or U8406 (N_8406,N_8225,N_8047);
nand U8407 (N_8407,N_8210,N_8226);
nand U8408 (N_8408,N_8122,N_8012);
and U8409 (N_8409,N_8173,N_8094);
xnor U8410 (N_8410,N_8164,N_8053);
xor U8411 (N_8411,N_8117,N_8228);
nand U8412 (N_8412,N_8069,N_8193);
nor U8413 (N_8413,N_8154,N_8064);
nand U8414 (N_8414,N_8014,N_8099);
nor U8415 (N_8415,N_8204,N_8123);
or U8416 (N_8416,N_8152,N_8094);
nor U8417 (N_8417,N_8067,N_8226);
or U8418 (N_8418,N_8002,N_8219);
and U8419 (N_8419,N_8158,N_8045);
nand U8420 (N_8420,N_8158,N_8202);
nand U8421 (N_8421,N_8021,N_8001);
nand U8422 (N_8422,N_8109,N_8066);
nand U8423 (N_8423,N_8243,N_8007);
nor U8424 (N_8424,N_8010,N_8240);
and U8425 (N_8425,N_8206,N_8091);
and U8426 (N_8426,N_8005,N_8249);
and U8427 (N_8427,N_8090,N_8232);
or U8428 (N_8428,N_8139,N_8135);
nor U8429 (N_8429,N_8085,N_8161);
and U8430 (N_8430,N_8192,N_8016);
and U8431 (N_8431,N_8128,N_8127);
nand U8432 (N_8432,N_8044,N_8060);
nor U8433 (N_8433,N_8182,N_8098);
and U8434 (N_8434,N_8079,N_8076);
nand U8435 (N_8435,N_8193,N_8167);
or U8436 (N_8436,N_8163,N_8106);
nand U8437 (N_8437,N_8203,N_8012);
nand U8438 (N_8438,N_8170,N_8060);
nand U8439 (N_8439,N_8211,N_8166);
nor U8440 (N_8440,N_8072,N_8060);
xor U8441 (N_8441,N_8227,N_8173);
and U8442 (N_8442,N_8238,N_8113);
nor U8443 (N_8443,N_8138,N_8187);
nor U8444 (N_8444,N_8217,N_8025);
xor U8445 (N_8445,N_8207,N_8195);
or U8446 (N_8446,N_8070,N_8168);
or U8447 (N_8447,N_8118,N_8153);
and U8448 (N_8448,N_8229,N_8148);
nand U8449 (N_8449,N_8109,N_8046);
xnor U8450 (N_8450,N_8057,N_8238);
nand U8451 (N_8451,N_8078,N_8003);
nand U8452 (N_8452,N_8086,N_8008);
nor U8453 (N_8453,N_8220,N_8141);
xor U8454 (N_8454,N_8155,N_8040);
xor U8455 (N_8455,N_8149,N_8035);
nor U8456 (N_8456,N_8215,N_8028);
nand U8457 (N_8457,N_8137,N_8100);
nand U8458 (N_8458,N_8052,N_8148);
nand U8459 (N_8459,N_8239,N_8161);
and U8460 (N_8460,N_8136,N_8163);
or U8461 (N_8461,N_8041,N_8076);
xnor U8462 (N_8462,N_8197,N_8237);
xnor U8463 (N_8463,N_8193,N_8176);
nand U8464 (N_8464,N_8093,N_8203);
and U8465 (N_8465,N_8202,N_8124);
or U8466 (N_8466,N_8135,N_8088);
nor U8467 (N_8467,N_8082,N_8191);
and U8468 (N_8468,N_8106,N_8241);
xor U8469 (N_8469,N_8085,N_8232);
nand U8470 (N_8470,N_8042,N_8059);
xnor U8471 (N_8471,N_8074,N_8060);
or U8472 (N_8472,N_8222,N_8127);
nor U8473 (N_8473,N_8216,N_8126);
nor U8474 (N_8474,N_8040,N_8050);
or U8475 (N_8475,N_8020,N_8043);
nand U8476 (N_8476,N_8000,N_8017);
xor U8477 (N_8477,N_8006,N_8165);
and U8478 (N_8478,N_8213,N_8062);
nor U8479 (N_8479,N_8099,N_8216);
nor U8480 (N_8480,N_8019,N_8234);
or U8481 (N_8481,N_8233,N_8108);
xor U8482 (N_8482,N_8069,N_8176);
or U8483 (N_8483,N_8160,N_8175);
and U8484 (N_8484,N_8040,N_8033);
nor U8485 (N_8485,N_8064,N_8091);
and U8486 (N_8486,N_8053,N_8117);
or U8487 (N_8487,N_8021,N_8046);
or U8488 (N_8488,N_8145,N_8034);
and U8489 (N_8489,N_8178,N_8072);
or U8490 (N_8490,N_8204,N_8119);
or U8491 (N_8491,N_8116,N_8149);
xor U8492 (N_8492,N_8014,N_8185);
nor U8493 (N_8493,N_8037,N_8127);
nor U8494 (N_8494,N_8244,N_8150);
nor U8495 (N_8495,N_8220,N_8018);
nand U8496 (N_8496,N_8047,N_8220);
or U8497 (N_8497,N_8006,N_8022);
xor U8498 (N_8498,N_8028,N_8073);
nand U8499 (N_8499,N_8129,N_8124);
nor U8500 (N_8500,N_8466,N_8281);
xor U8501 (N_8501,N_8334,N_8475);
nand U8502 (N_8502,N_8458,N_8438);
and U8503 (N_8503,N_8273,N_8384);
or U8504 (N_8504,N_8369,N_8288);
nor U8505 (N_8505,N_8477,N_8425);
or U8506 (N_8506,N_8390,N_8305);
or U8507 (N_8507,N_8387,N_8381);
nand U8508 (N_8508,N_8331,N_8484);
xnor U8509 (N_8509,N_8278,N_8328);
nor U8510 (N_8510,N_8299,N_8327);
or U8511 (N_8511,N_8271,N_8440);
nor U8512 (N_8512,N_8364,N_8285);
nand U8513 (N_8513,N_8252,N_8471);
xnor U8514 (N_8514,N_8362,N_8416);
or U8515 (N_8515,N_8361,N_8374);
and U8516 (N_8516,N_8332,N_8368);
and U8517 (N_8517,N_8419,N_8437);
nor U8518 (N_8518,N_8307,N_8447);
nand U8519 (N_8519,N_8263,N_8279);
nor U8520 (N_8520,N_8375,N_8460);
xnor U8521 (N_8521,N_8376,N_8396);
xor U8522 (N_8522,N_8456,N_8256);
nand U8523 (N_8523,N_8359,N_8311);
xnor U8524 (N_8524,N_8424,N_8257);
and U8525 (N_8525,N_8428,N_8323);
nand U8526 (N_8526,N_8302,N_8457);
nand U8527 (N_8527,N_8345,N_8344);
or U8528 (N_8528,N_8270,N_8267);
nor U8529 (N_8529,N_8338,N_8451);
and U8530 (N_8530,N_8349,N_8325);
nand U8531 (N_8531,N_8414,N_8371);
xnor U8532 (N_8532,N_8322,N_8446);
and U8533 (N_8533,N_8467,N_8356);
or U8534 (N_8534,N_8335,N_8410);
xnor U8535 (N_8535,N_8498,N_8272);
or U8536 (N_8536,N_8319,N_8391);
and U8537 (N_8537,N_8315,N_8493);
nor U8538 (N_8538,N_8499,N_8340);
nand U8539 (N_8539,N_8432,N_8380);
or U8540 (N_8540,N_8337,N_8261);
nand U8541 (N_8541,N_8353,N_8379);
or U8542 (N_8542,N_8405,N_8312);
nor U8543 (N_8543,N_8304,N_8255);
and U8544 (N_8544,N_8491,N_8295);
nand U8545 (N_8545,N_8439,N_8420);
and U8546 (N_8546,N_8465,N_8486);
nand U8547 (N_8547,N_8348,N_8321);
or U8548 (N_8548,N_8277,N_8297);
nand U8549 (N_8549,N_8452,N_8352);
or U8550 (N_8550,N_8407,N_8434);
nand U8551 (N_8551,N_8365,N_8427);
or U8552 (N_8552,N_8430,N_8265);
xnor U8553 (N_8553,N_8284,N_8413);
or U8554 (N_8554,N_8314,N_8382);
and U8555 (N_8555,N_8462,N_8399);
nor U8556 (N_8556,N_8274,N_8421);
or U8557 (N_8557,N_8301,N_8294);
xnor U8558 (N_8558,N_8268,N_8494);
nand U8559 (N_8559,N_8287,N_8495);
or U8560 (N_8560,N_8351,N_8482);
nor U8561 (N_8561,N_8318,N_8378);
nor U8562 (N_8562,N_8431,N_8300);
nand U8563 (N_8563,N_8269,N_8476);
nor U8564 (N_8564,N_8443,N_8490);
and U8565 (N_8565,N_8330,N_8259);
nor U8566 (N_8566,N_8343,N_8426);
and U8567 (N_8567,N_8481,N_8472);
nor U8568 (N_8568,N_8292,N_8479);
or U8569 (N_8569,N_8409,N_8354);
nor U8570 (N_8570,N_8441,N_8290);
nor U8571 (N_8571,N_8324,N_8463);
and U8572 (N_8572,N_8346,N_8429);
nand U8573 (N_8573,N_8286,N_8289);
nand U8574 (N_8574,N_8342,N_8393);
nand U8575 (N_8575,N_8400,N_8389);
xnor U8576 (N_8576,N_8464,N_8291);
nor U8577 (N_8577,N_8316,N_8398);
and U8578 (N_8578,N_8411,N_8461);
or U8579 (N_8579,N_8282,N_8310);
nor U8580 (N_8580,N_8402,N_8296);
nor U8581 (N_8581,N_8436,N_8308);
nor U8582 (N_8582,N_8469,N_8317);
nand U8583 (N_8583,N_8473,N_8320);
or U8584 (N_8584,N_8459,N_8341);
and U8585 (N_8585,N_8485,N_8404);
nand U8586 (N_8586,N_8403,N_8417);
and U8587 (N_8587,N_8406,N_8388);
or U8588 (N_8588,N_8448,N_8276);
xnor U8589 (N_8589,N_8250,N_8360);
or U8590 (N_8590,N_8253,N_8468);
nand U8591 (N_8591,N_8373,N_8370);
nor U8592 (N_8592,N_8264,N_8313);
nor U8593 (N_8593,N_8363,N_8497);
and U8594 (N_8594,N_8366,N_8260);
nand U8595 (N_8595,N_8350,N_8336);
and U8596 (N_8596,N_8347,N_8455);
xnor U8597 (N_8597,N_8266,N_8445);
nand U8598 (N_8598,N_8254,N_8258);
nand U8599 (N_8599,N_8478,N_8358);
or U8600 (N_8600,N_8262,N_8422);
nand U8601 (N_8601,N_8280,N_8454);
nand U8602 (N_8602,N_8453,N_8283);
nand U8603 (N_8603,N_8418,N_8377);
nor U8604 (N_8604,N_8395,N_8385);
and U8605 (N_8605,N_8480,N_8397);
or U8606 (N_8606,N_8383,N_8483);
xnor U8607 (N_8607,N_8412,N_8372);
and U8608 (N_8608,N_8309,N_8386);
or U8609 (N_8609,N_8492,N_8487);
or U8610 (N_8610,N_8298,N_8326);
or U8611 (N_8611,N_8306,N_8496);
nor U8612 (N_8612,N_8329,N_8394);
xnor U8613 (N_8613,N_8433,N_8367);
nand U8614 (N_8614,N_8357,N_8449);
or U8615 (N_8615,N_8435,N_8275);
nor U8616 (N_8616,N_8423,N_8489);
and U8617 (N_8617,N_8392,N_8401);
nand U8618 (N_8618,N_8339,N_8470);
or U8619 (N_8619,N_8450,N_8474);
or U8620 (N_8620,N_8442,N_8415);
and U8621 (N_8621,N_8293,N_8408);
and U8622 (N_8622,N_8333,N_8251);
nand U8623 (N_8623,N_8303,N_8355);
and U8624 (N_8624,N_8444,N_8488);
nand U8625 (N_8625,N_8415,N_8424);
xnor U8626 (N_8626,N_8357,N_8252);
xnor U8627 (N_8627,N_8381,N_8489);
nand U8628 (N_8628,N_8463,N_8485);
nand U8629 (N_8629,N_8265,N_8392);
xnor U8630 (N_8630,N_8438,N_8374);
and U8631 (N_8631,N_8349,N_8425);
xor U8632 (N_8632,N_8491,N_8499);
nand U8633 (N_8633,N_8432,N_8456);
xor U8634 (N_8634,N_8404,N_8336);
nand U8635 (N_8635,N_8417,N_8256);
and U8636 (N_8636,N_8384,N_8371);
nor U8637 (N_8637,N_8387,N_8446);
or U8638 (N_8638,N_8275,N_8259);
and U8639 (N_8639,N_8318,N_8443);
xor U8640 (N_8640,N_8488,N_8337);
nor U8641 (N_8641,N_8300,N_8264);
or U8642 (N_8642,N_8484,N_8458);
nand U8643 (N_8643,N_8463,N_8446);
and U8644 (N_8644,N_8262,N_8406);
nor U8645 (N_8645,N_8451,N_8381);
and U8646 (N_8646,N_8272,N_8474);
nor U8647 (N_8647,N_8310,N_8308);
nand U8648 (N_8648,N_8373,N_8421);
xnor U8649 (N_8649,N_8457,N_8313);
and U8650 (N_8650,N_8353,N_8344);
nor U8651 (N_8651,N_8499,N_8377);
and U8652 (N_8652,N_8303,N_8343);
xor U8653 (N_8653,N_8447,N_8422);
nor U8654 (N_8654,N_8396,N_8412);
xor U8655 (N_8655,N_8432,N_8383);
nor U8656 (N_8656,N_8284,N_8429);
xnor U8657 (N_8657,N_8286,N_8363);
nor U8658 (N_8658,N_8409,N_8312);
and U8659 (N_8659,N_8343,N_8286);
xor U8660 (N_8660,N_8326,N_8297);
nand U8661 (N_8661,N_8399,N_8473);
or U8662 (N_8662,N_8294,N_8495);
nor U8663 (N_8663,N_8480,N_8380);
nor U8664 (N_8664,N_8442,N_8432);
nor U8665 (N_8665,N_8378,N_8316);
nor U8666 (N_8666,N_8350,N_8289);
nand U8667 (N_8667,N_8482,N_8491);
nor U8668 (N_8668,N_8301,N_8313);
xor U8669 (N_8669,N_8290,N_8312);
nand U8670 (N_8670,N_8349,N_8391);
nor U8671 (N_8671,N_8422,N_8295);
or U8672 (N_8672,N_8408,N_8346);
or U8673 (N_8673,N_8324,N_8486);
xnor U8674 (N_8674,N_8445,N_8476);
and U8675 (N_8675,N_8482,N_8410);
xor U8676 (N_8676,N_8264,N_8478);
and U8677 (N_8677,N_8368,N_8379);
xor U8678 (N_8678,N_8260,N_8438);
nand U8679 (N_8679,N_8483,N_8470);
nor U8680 (N_8680,N_8406,N_8315);
nor U8681 (N_8681,N_8458,N_8399);
or U8682 (N_8682,N_8334,N_8338);
and U8683 (N_8683,N_8420,N_8423);
and U8684 (N_8684,N_8283,N_8254);
or U8685 (N_8685,N_8460,N_8419);
or U8686 (N_8686,N_8448,N_8433);
and U8687 (N_8687,N_8476,N_8357);
nand U8688 (N_8688,N_8263,N_8384);
and U8689 (N_8689,N_8398,N_8497);
xor U8690 (N_8690,N_8478,N_8317);
or U8691 (N_8691,N_8361,N_8264);
and U8692 (N_8692,N_8323,N_8424);
nor U8693 (N_8693,N_8315,N_8474);
nand U8694 (N_8694,N_8457,N_8371);
nor U8695 (N_8695,N_8430,N_8422);
nand U8696 (N_8696,N_8291,N_8443);
or U8697 (N_8697,N_8317,N_8382);
and U8698 (N_8698,N_8311,N_8472);
nor U8699 (N_8699,N_8336,N_8424);
and U8700 (N_8700,N_8354,N_8267);
xor U8701 (N_8701,N_8283,N_8389);
or U8702 (N_8702,N_8312,N_8302);
and U8703 (N_8703,N_8327,N_8279);
and U8704 (N_8704,N_8304,N_8302);
or U8705 (N_8705,N_8328,N_8450);
xnor U8706 (N_8706,N_8455,N_8453);
or U8707 (N_8707,N_8369,N_8485);
xor U8708 (N_8708,N_8380,N_8451);
nand U8709 (N_8709,N_8292,N_8266);
nor U8710 (N_8710,N_8387,N_8391);
nand U8711 (N_8711,N_8467,N_8443);
xor U8712 (N_8712,N_8310,N_8448);
xnor U8713 (N_8713,N_8352,N_8253);
nand U8714 (N_8714,N_8401,N_8496);
and U8715 (N_8715,N_8361,N_8350);
nand U8716 (N_8716,N_8297,N_8273);
nor U8717 (N_8717,N_8370,N_8344);
xor U8718 (N_8718,N_8420,N_8267);
or U8719 (N_8719,N_8266,N_8389);
nor U8720 (N_8720,N_8290,N_8389);
xnor U8721 (N_8721,N_8470,N_8365);
or U8722 (N_8722,N_8265,N_8375);
or U8723 (N_8723,N_8495,N_8404);
xnor U8724 (N_8724,N_8266,N_8388);
nand U8725 (N_8725,N_8397,N_8294);
nand U8726 (N_8726,N_8468,N_8309);
nor U8727 (N_8727,N_8423,N_8306);
nor U8728 (N_8728,N_8425,N_8306);
nand U8729 (N_8729,N_8298,N_8458);
and U8730 (N_8730,N_8455,N_8372);
xor U8731 (N_8731,N_8350,N_8465);
and U8732 (N_8732,N_8280,N_8477);
or U8733 (N_8733,N_8303,N_8350);
nand U8734 (N_8734,N_8413,N_8448);
or U8735 (N_8735,N_8475,N_8451);
nor U8736 (N_8736,N_8368,N_8418);
nand U8737 (N_8737,N_8476,N_8365);
nor U8738 (N_8738,N_8349,N_8424);
nor U8739 (N_8739,N_8481,N_8424);
nor U8740 (N_8740,N_8481,N_8251);
nand U8741 (N_8741,N_8336,N_8453);
xor U8742 (N_8742,N_8465,N_8409);
and U8743 (N_8743,N_8379,N_8460);
nand U8744 (N_8744,N_8429,N_8475);
nand U8745 (N_8745,N_8449,N_8397);
nand U8746 (N_8746,N_8453,N_8304);
nor U8747 (N_8747,N_8487,N_8394);
nor U8748 (N_8748,N_8476,N_8372);
nand U8749 (N_8749,N_8254,N_8318);
xor U8750 (N_8750,N_8730,N_8574);
nand U8751 (N_8751,N_8700,N_8654);
nor U8752 (N_8752,N_8674,N_8668);
nand U8753 (N_8753,N_8504,N_8536);
and U8754 (N_8754,N_8633,N_8659);
and U8755 (N_8755,N_8617,N_8718);
nor U8756 (N_8756,N_8732,N_8639);
nand U8757 (N_8757,N_8747,N_8699);
nor U8758 (N_8758,N_8685,N_8527);
nand U8759 (N_8759,N_8612,N_8728);
or U8760 (N_8760,N_8604,N_8535);
nand U8761 (N_8761,N_8680,N_8634);
nand U8762 (N_8762,N_8560,N_8585);
nor U8763 (N_8763,N_8610,N_8726);
or U8764 (N_8764,N_8652,N_8598);
xor U8765 (N_8765,N_8614,N_8505);
or U8766 (N_8766,N_8664,N_8520);
and U8767 (N_8767,N_8740,N_8651);
or U8768 (N_8768,N_8736,N_8507);
nand U8769 (N_8769,N_8596,N_8570);
xnor U8770 (N_8770,N_8569,N_8717);
nand U8771 (N_8771,N_8551,N_8526);
nor U8772 (N_8772,N_8653,N_8546);
nand U8773 (N_8773,N_8545,N_8713);
and U8774 (N_8774,N_8741,N_8684);
xor U8775 (N_8775,N_8648,N_8589);
nor U8776 (N_8776,N_8539,N_8559);
or U8777 (N_8777,N_8580,N_8622);
nand U8778 (N_8778,N_8739,N_8603);
and U8779 (N_8779,N_8588,N_8661);
xnor U8780 (N_8780,N_8655,N_8723);
and U8781 (N_8781,N_8675,N_8558);
xnor U8782 (N_8782,N_8537,N_8609);
and U8783 (N_8783,N_8660,N_8522);
xor U8784 (N_8784,N_8693,N_8708);
and U8785 (N_8785,N_8694,N_8669);
nor U8786 (N_8786,N_8646,N_8529);
and U8787 (N_8787,N_8666,N_8600);
nor U8788 (N_8788,N_8679,N_8689);
and U8789 (N_8789,N_8583,N_8641);
nand U8790 (N_8790,N_8613,N_8615);
nand U8791 (N_8791,N_8688,N_8626);
xnor U8792 (N_8792,N_8709,N_8592);
and U8793 (N_8793,N_8575,N_8550);
nand U8794 (N_8794,N_8698,N_8725);
and U8795 (N_8795,N_8638,N_8673);
or U8796 (N_8796,N_8542,N_8636);
xor U8797 (N_8797,N_8548,N_8735);
xnor U8798 (N_8798,N_8722,N_8543);
nor U8799 (N_8799,N_8538,N_8681);
nand U8800 (N_8800,N_8662,N_8625);
nand U8801 (N_8801,N_8595,N_8720);
nor U8802 (N_8802,N_8564,N_8519);
nor U8803 (N_8803,N_8534,N_8606);
and U8804 (N_8804,N_8555,N_8593);
nor U8805 (N_8805,N_8678,N_8733);
and U8806 (N_8806,N_8657,N_8640);
or U8807 (N_8807,N_8599,N_8523);
nor U8808 (N_8808,N_8517,N_8530);
nand U8809 (N_8809,N_8509,N_8690);
nand U8810 (N_8810,N_8682,N_8686);
nor U8811 (N_8811,N_8586,N_8511);
nor U8812 (N_8812,N_8642,N_8544);
nor U8813 (N_8813,N_8576,N_8621);
and U8814 (N_8814,N_8581,N_8587);
nor U8815 (N_8815,N_8671,N_8670);
and U8816 (N_8816,N_8711,N_8712);
and U8817 (N_8817,N_8676,N_8532);
xor U8818 (N_8818,N_8578,N_8719);
and U8819 (N_8819,N_8518,N_8649);
xnor U8820 (N_8820,N_8553,N_8746);
nand U8821 (N_8821,N_8724,N_8687);
and U8822 (N_8822,N_8540,N_8703);
xor U8823 (N_8823,N_8714,N_8742);
nor U8824 (N_8824,N_8658,N_8528);
and U8825 (N_8825,N_8514,N_8738);
or U8826 (N_8826,N_8557,N_8696);
xor U8827 (N_8827,N_8629,N_8510);
nand U8828 (N_8828,N_8608,N_8620);
and U8829 (N_8829,N_8635,N_8547);
or U8830 (N_8830,N_8607,N_8549);
nand U8831 (N_8831,N_8566,N_8710);
xnor U8832 (N_8832,N_8631,N_8748);
nand U8833 (N_8833,N_8737,N_8573);
nor U8834 (N_8834,N_8695,N_8565);
nand U8835 (N_8835,N_8582,N_8691);
and U8836 (N_8836,N_8508,N_8734);
and U8837 (N_8837,N_8590,N_8597);
xor U8838 (N_8838,N_8561,N_8513);
nand U8839 (N_8839,N_8647,N_8749);
and U8840 (N_8840,N_8643,N_8524);
and U8841 (N_8841,N_8611,N_8656);
and U8842 (N_8842,N_8562,N_8502);
xnor U8843 (N_8843,N_8637,N_8706);
xnor U8844 (N_8844,N_8619,N_8672);
nand U8845 (N_8845,N_8716,N_8533);
nor U8846 (N_8846,N_8503,N_8515);
or U8847 (N_8847,N_8697,N_8572);
or U8848 (N_8848,N_8624,N_8650);
nand U8849 (N_8849,N_8506,N_8705);
and U8850 (N_8850,N_8628,N_8601);
xor U8851 (N_8851,N_8584,N_8721);
nor U8852 (N_8852,N_8579,N_8727);
and U8853 (N_8853,N_8556,N_8577);
or U8854 (N_8854,N_8704,N_8541);
or U8855 (N_8855,N_8512,N_8667);
or U8856 (N_8856,N_8644,N_8677);
xnor U8857 (N_8857,N_8632,N_8745);
or U8858 (N_8858,N_8521,N_8525);
xor U8859 (N_8859,N_8707,N_8605);
and U8860 (N_8860,N_8630,N_8531);
xor U8861 (N_8861,N_8500,N_8594);
or U8862 (N_8862,N_8702,N_8616);
or U8863 (N_8863,N_8563,N_8729);
and U8864 (N_8864,N_8731,N_8568);
xor U8865 (N_8865,N_8602,N_8663);
xor U8866 (N_8866,N_8591,N_8665);
nand U8867 (N_8867,N_8715,N_8645);
xor U8868 (N_8868,N_8501,N_8683);
and U8869 (N_8869,N_8623,N_8744);
xor U8870 (N_8870,N_8692,N_8627);
or U8871 (N_8871,N_8567,N_8618);
or U8872 (N_8872,N_8743,N_8701);
nor U8873 (N_8873,N_8571,N_8552);
or U8874 (N_8874,N_8516,N_8554);
or U8875 (N_8875,N_8638,N_8517);
nor U8876 (N_8876,N_8509,N_8714);
nor U8877 (N_8877,N_8725,N_8580);
nand U8878 (N_8878,N_8637,N_8719);
and U8879 (N_8879,N_8720,N_8645);
nand U8880 (N_8880,N_8514,N_8689);
and U8881 (N_8881,N_8640,N_8500);
or U8882 (N_8882,N_8576,N_8528);
nand U8883 (N_8883,N_8525,N_8642);
nand U8884 (N_8884,N_8526,N_8537);
nor U8885 (N_8885,N_8514,N_8688);
and U8886 (N_8886,N_8666,N_8717);
nand U8887 (N_8887,N_8561,N_8518);
nor U8888 (N_8888,N_8533,N_8665);
or U8889 (N_8889,N_8520,N_8675);
and U8890 (N_8890,N_8698,N_8703);
nand U8891 (N_8891,N_8744,N_8676);
and U8892 (N_8892,N_8619,N_8624);
nor U8893 (N_8893,N_8557,N_8595);
nand U8894 (N_8894,N_8505,N_8613);
nand U8895 (N_8895,N_8571,N_8721);
xnor U8896 (N_8896,N_8593,N_8573);
xnor U8897 (N_8897,N_8509,N_8534);
xor U8898 (N_8898,N_8693,N_8661);
or U8899 (N_8899,N_8565,N_8562);
nor U8900 (N_8900,N_8635,N_8622);
xnor U8901 (N_8901,N_8682,N_8557);
nand U8902 (N_8902,N_8703,N_8710);
xor U8903 (N_8903,N_8615,N_8552);
nor U8904 (N_8904,N_8506,N_8680);
xnor U8905 (N_8905,N_8627,N_8610);
and U8906 (N_8906,N_8699,N_8510);
nor U8907 (N_8907,N_8550,N_8669);
xnor U8908 (N_8908,N_8694,N_8554);
nand U8909 (N_8909,N_8548,N_8528);
nand U8910 (N_8910,N_8707,N_8649);
xnor U8911 (N_8911,N_8535,N_8566);
or U8912 (N_8912,N_8700,N_8605);
and U8913 (N_8913,N_8648,N_8666);
or U8914 (N_8914,N_8556,N_8655);
xnor U8915 (N_8915,N_8530,N_8716);
nor U8916 (N_8916,N_8721,N_8574);
nand U8917 (N_8917,N_8736,N_8617);
nand U8918 (N_8918,N_8725,N_8621);
nand U8919 (N_8919,N_8672,N_8725);
or U8920 (N_8920,N_8557,N_8649);
or U8921 (N_8921,N_8550,N_8651);
nand U8922 (N_8922,N_8631,N_8532);
or U8923 (N_8923,N_8624,N_8622);
nand U8924 (N_8924,N_8633,N_8613);
xor U8925 (N_8925,N_8662,N_8545);
and U8926 (N_8926,N_8699,N_8646);
or U8927 (N_8927,N_8505,N_8741);
nor U8928 (N_8928,N_8557,N_8628);
and U8929 (N_8929,N_8531,N_8617);
or U8930 (N_8930,N_8709,N_8563);
nor U8931 (N_8931,N_8621,N_8720);
xnor U8932 (N_8932,N_8527,N_8691);
xnor U8933 (N_8933,N_8506,N_8509);
xor U8934 (N_8934,N_8596,N_8531);
xor U8935 (N_8935,N_8585,N_8584);
xnor U8936 (N_8936,N_8570,N_8562);
xnor U8937 (N_8937,N_8561,N_8673);
and U8938 (N_8938,N_8714,N_8689);
and U8939 (N_8939,N_8572,N_8684);
nand U8940 (N_8940,N_8599,N_8666);
and U8941 (N_8941,N_8541,N_8672);
and U8942 (N_8942,N_8639,N_8574);
or U8943 (N_8943,N_8573,N_8509);
xor U8944 (N_8944,N_8741,N_8546);
xnor U8945 (N_8945,N_8635,N_8587);
xor U8946 (N_8946,N_8616,N_8690);
nor U8947 (N_8947,N_8645,N_8524);
and U8948 (N_8948,N_8641,N_8553);
xor U8949 (N_8949,N_8574,N_8630);
and U8950 (N_8950,N_8644,N_8502);
xnor U8951 (N_8951,N_8713,N_8668);
xor U8952 (N_8952,N_8545,N_8583);
and U8953 (N_8953,N_8555,N_8702);
nor U8954 (N_8954,N_8504,N_8528);
xor U8955 (N_8955,N_8590,N_8662);
and U8956 (N_8956,N_8745,N_8524);
xnor U8957 (N_8957,N_8703,N_8735);
or U8958 (N_8958,N_8575,N_8723);
or U8959 (N_8959,N_8565,N_8635);
and U8960 (N_8960,N_8527,N_8584);
or U8961 (N_8961,N_8574,N_8579);
or U8962 (N_8962,N_8743,N_8657);
or U8963 (N_8963,N_8740,N_8655);
nand U8964 (N_8964,N_8558,N_8705);
and U8965 (N_8965,N_8566,N_8552);
nand U8966 (N_8966,N_8666,N_8553);
or U8967 (N_8967,N_8745,N_8611);
nand U8968 (N_8968,N_8583,N_8721);
or U8969 (N_8969,N_8645,N_8567);
xor U8970 (N_8970,N_8725,N_8687);
nor U8971 (N_8971,N_8644,N_8512);
nand U8972 (N_8972,N_8599,N_8543);
nand U8973 (N_8973,N_8748,N_8647);
xnor U8974 (N_8974,N_8607,N_8686);
and U8975 (N_8975,N_8742,N_8505);
xor U8976 (N_8976,N_8549,N_8588);
and U8977 (N_8977,N_8639,N_8683);
xor U8978 (N_8978,N_8656,N_8735);
and U8979 (N_8979,N_8532,N_8557);
xnor U8980 (N_8980,N_8529,N_8544);
nand U8981 (N_8981,N_8716,N_8630);
nor U8982 (N_8982,N_8727,N_8647);
nand U8983 (N_8983,N_8632,N_8637);
and U8984 (N_8984,N_8585,N_8520);
xnor U8985 (N_8985,N_8579,N_8728);
and U8986 (N_8986,N_8646,N_8675);
or U8987 (N_8987,N_8734,N_8703);
xnor U8988 (N_8988,N_8663,N_8617);
nor U8989 (N_8989,N_8527,N_8534);
xor U8990 (N_8990,N_8528,N_8697);
or U8991 (N_8991,N_8520,N_8622);
nor U8992 (N_8992,N_8575,N_8656);
or U8993 (N_8993,N_8564,N_8672);
and U8994 (N_8994,N_8717,N_8641);
or U8995 (N_8995,N_8740,N_8578);
nor U8996 (N_8996,N_8596,N_8671);
and U8997 (N_8997,N_8677,N_8715);
or U8998 (N_8998,N_8745,N_8739);
nor U8999 (N_8999,N_8632,N_8735);
nor U9000 (N_9000,N_8907,N_8976);
nand U9001 (N_9001,N_8784,N_8862);
and U9002 (N_9002,N_8810,N_8765);
or U9003 (N_9003,N_8776,N_8966);
nor U9004 (N_9004,N_8970,N_8787);
nor U9005 (N_9005,N_8897,N_8918);
xnor U9006 (N_9006,N_8969,N_8890);
and U9007 (N_9007,N_8985,N_8769);
nor U9008 (N_9008,N_8874,N_8791);
nand U9009 (N_9009,N_8829,N_8799);
and U9010 (N_9010,N_8886,N_8980);
xnor U9011 (N_9011,N_8906,N_8992);
nand U9012 (N_9012,N_8910,N_8831);
and U9013 (N_9013,N_8993,N_8943);
xor U9014 (N_9014,N_8837,N_8783);
nor U9015 (N_9015,N_8861,N_8770);
nand U9016 (N_9016,N_8940,N_8815);
and U9017 (N_9017,N_8841,N_8795);
and U9018 (N_9018,N_8979,N_8871);
nand U9019 (N_9019,N_8800,N_8796);
nand U9020 (N_9020,N_8935,N_8928);
xnor U9021 (N_9021,N_8982,N_8905);
or U9022 (N_9022,N_8998,N_8900);
or U9023 (N_9023,N_8822,N_8768);
and U9024 (N_9024,N_8760,N_8779);
or U9025 (N_9025,N_8830,N_8858);
xnor U9026 (N_9026,N_8855,N_8938);
or U9027 (N_9027,N_8798,N_8794);
xnor U9028 (N_9028,N_8773,N_8898);
xnor U9029 (N_9029,N_8946,N_8869);
and U9030 (N_9030,N_8961,N_8952);
nand U9031 (N_9031,N_8836,N_8911);
and U9032 (N_9032,N_8756,N_8925);
and U9033 (N_9033,N_8967,N_8842);
nor U9034 (N_9034,N_8843,N_8932);
and U9035 (N_9035,N_8885,N_8939);
xor U9036 (N_9036,N_8949,N_8922);
nor U9037 (N_9037,N_8959,N_8806);
xnor U9038 (N_9038,N_8936,N_8927);
xnor U9039 (N_9039,N_8920,N_8973);
xnor U9040 (N_9040,N_8751,N_8995);
nor U9041 (N_9041,N_8947,N_8767);
xor U9042 (N_9042,N_8872,N_8945);
or U9043 (N_9043,N_8817,N_8917);
or U9044 (N_9044,N_8934,N_8974);
or U9045 (N_9045,N_8875,N_8848);
xor U9046 (N_9046,N_8963,N_8852);
nor U9047 (N_9047,N_8893,N_8811);
nand U9048 (N_9048,N_8851,N_8924);
xnor U9049 (N_9049,N_8792,N_8833);
and U9050 (N_9050,N_8816,N_8987);
and U9051 (N_9051,N_8790,N_8864);
and U9052 (N_9052,N_8990,N_8901);
or U9053 (N_9053,N_8954,N_8996);
or U9054 (N_9054,N_8902,N_8785);
and U9055 (N_9055,N_8919,N_8950);
nor U9056 (N_9056,N_8797,N_8951);
and U9057 (N_9057,N_8754,N_8884);
and U9058 (N_9058,N_8860,N_8827);
and U9059 (N_9059,N_8908,N_8834);
nand U9060 (N_9060,N_8809,N_8888);
nor U9061 (N_9061,N_8866,N_8962);
and U9062 (N_9062,N_8999,N_8757);
or U9063 (N_9063,N_8899,N_8802);
nand U9064 (N_9064,N_8981,N_8929);
nand U9065 (N_9065,N_8984,N_8820);
or U9066 (N_9066,N_8892,N_8804);
or U9067 (N_9067,N_8873,N_8994);
nor U9068 (N_9068,N_8965,N_8821);
or U9069 (N_9069,N_8989,N_8953);
xnor U9070 (N_9070,N_8759,N_8904);
or U9071 (N_9071,N_8882,N_8846);
nand U9072 (N_9072,N_8930,N_8788);
xor U9073 (N_9073,N_8891,N_8778);
or U9074 (N_9074,N_8896,N_8828);
nand U9075 (N_9075,N_8941,N_8983);
or U9076 (N_9076,N_8801,N_8844);
or U9077 (N_9077,N_8845,N_8823);
nor U9078 (N_9078,N_8877,N_8880);
or U9079 (N_9079,N_8789,N_8913);
or U9080 (N_9080,N_8782,N_8781);
nand U9081 (N_9081,N_8771,N_8761);
and U9082 (N_9082,N_8857,N_8988);
nand U9083 (N_9083,N_8755,N_8964);
and U9084 (N_9084,N_8840,N_8942);
nor U9085 (N_9085,N_8955,N_8876);
or U9086 (N_9086,N_8838,N_8889);
and U9087 (N_9087,N_8859,N_8752);
and U9088 (N_9088,N_8786,N_8793);
and U9089 (N_9089,N_8933,N_8839);
nand U9090 (N_9090,N_8774,N_8826);
nand U9091 (N_9091,N_8997,N_8926);
or U9092 (N_9092,N_8832,N_8975);
xnor U9093 (N_9093,N_8780,N_8854);
xnor U9094 (N_9094,N_8931,N_8956);
nor U9095 (N_9095,N_8763,N_8764);
nor U9096 (N_9096,N_8968,N_8818);
nand U9097 (N_9097,N_8895,N_8819);
nand U9098 (N_9098,N_8775,N_8958);
or U9099 (N_9099,N_8803,N_8825);
nor U9100 (N_9100,N_8868,N_8903);
nor U9101 (N_9101,N_8863,N_8808);
nand U9102 (N_9102,N_8865,N_8847);
nor U9103 (N_9103,N_8813,N_8960);
nor U9104 (N_9104,N_8881,N_8753);
xor U9105 (N_9105,N_8909,N_8957);
xor U9106 (N_9106,N_8777,N_8883);
nor U9107 (N_9107,N_8766,N_8758);
nand U9108 (N_9108,N_8879,N_8812);
and U9109 (N_9109,N_8750,N_8887);
nor U9110 (N_9110,N_8894,N_8867);
nor U9111 (N_9111,N_8835,N_8824);
and U9112 (N_9112,N_8986,N_8916);
nor U9113 (N_9113,N_8991,N_8849);
xor U9114 (N_9114,N_8805,N_8914);
xor U9115 (N_9115,N_8853,N_8870);
and U9116 (N_9116,N_8814,N_8948);
xnor U9117 (N_9117,N_8972,N_8762);
or U9118 (N_9118,N_8944,N_8807);
and U9119 (N_9119,N_8923,N_8772);
xor U9120 (N_9120,N_8937,N_8912);
or U9121 (N_9121,N_8856,N_8915);
nor U9122 (N_9122,N_8850,N_8921);
and U9123 (N_9123,N_8978,N_8878);
and U9124 (N_9124,N_8977,N_8971);
or U9125 (N_9125,N_8939,N_8914);
or U9126 (N_9126,N_8860,N_8971);
nor U9127 (N_9127,N_8846,N_8945);
nand U9128 (N_9128,N_8919,N_8862);
and U9129 (N_9129,N_8878,N_8844);
xor U9130 (N_9130,N_8756,N_8806);
nor U9131 (N_9131,N_8882,N_8934);
xor U9132 (N_9132,N_8867,N_8880);
nand U9133 (N_9133,N_8781,N_8904);
nand U9134 (N_9134,N_8844,N_8756);
and U9135 (N_9135,N_8890,N_8955);
nor U9136 (N_9136,N_8953,N_8899);
nor U9137 (N_9137,N_8897,N_8961);
nand U9138 (N_9138,N_8856,N_8879);
xor U9139 (N_9139,N_8805,N_8960);
nand U9140 (N_9140,N_8851,N_8921);
xnor U9141 (N_9141,N_8965,N_8914);
xor U9142 (N_9142,N_8999,N_8847);
or U9143 (N_9143,N_8892,N_8963);
nand U9144 (N_9144,N_8831,N_8841);
nor U9145 (N_9145,N_8921,N_8830);
or U9146 (N_9146,N_8936,N_8793);
nor U9147 (N_9147,N_8991,N_8932);
xnor U9148 (N_9148,N_8800,N_8909);
nor U9149 (N_9149,N_8750,N_8949);
xor U9150 (N_9150,N_8782,N_8864);
xor U9151 (N_9151,N_8874,N_8916);
or U9152 (N_9152,N_8843,N_8946);
xor U9153 (N_9153,N_8798,N_8872);
nand U9154 (N_9154,N_8962,N_8984);
nor U9155 (N_9155,N_8964,N_8880);
or U9156 (N_9156,N_8842,N_8799);
nor U9157 (N_9157,N_8862,N_8927);
nand U9158 (N_9158,N_8979,N_8923);
xor U9159 (N_9159,N_8998,N_8771);
nor U9160 (N_9160,N_8937,N_8996);
and U9161 (N_9161,N_8799,N_8935);
and U9162 (N_9162,N_8782,N_8804);
or U9163 (N_9163,N_8945,N_8860);
or U9164 (N_9164,N_8788,N_8932);
or U9165 (N_9165,N_8814,N_8956);
nand U9166 (N_9166,N_8835,N_8945);
or U9167 (N_9167,N_8785,N_8865);
xnor U9168 (N_9168,N_8791,N_8816);
nand U9169 (N_9169,N_8982,N_8891);
or U9170 (N_9170,N_8897,N_8847);
or U9171 (N_9171,N_8901,N_8774);
nand U9172 (N_9172,N_8883,N_8829);
and U9173 (N_9173,N_8892,N_8877);
and U9174 (N_9174,N_8858,N_8825);
xor U9175 (N_9175,N_8878,N_8772);
nand U9176 (N_9176,N_8872,N_8764);
xor U9177 (N_9177,N_8890,N_8802);
nand U9178 (N_9178,N_8937,N_8762);
xnor U9179 (N_9179,N_8753,N_8990);
nor U9180 (N_9180,N_8839,N_8898);
and U9181 (N_9181,N_8771,N_8975);
xnor U9182 (N_9182,N_8769,N_8949);
xnor U9183 (N_9183,N_8919,N_8986);
nand U9184 (N_9184,N_8852,N_8928);
or U9185 (N_9185,N_8759,N_8825);
and U9186 (N_9186,N_8980,N_8876);
xor U9187 (N_9187,N_8964,N_8851);
or U9188 (N_9188,N_8830,N_8833);
nor U9189 (N_9189,N_8847,N_8772);
or U9190 (N_9190,N_8946,N_8815);
nand U9191 (N_9191,N_8860,N_8778);
or U9192 (N_9192,N_8792,N_8821);
or U9193 (N_9193,N_8827,N_8911);
and U9194 (N_9194,N_8976,N_8774);
xnor U9195 (N_9195,N_8794,N_8774);
xor U9196 (N_9196,N_8781,N_8750);
xnor U9197 (N_9197,N_8857,N_8820);
xnor U9198 (N_9198,N_8854,N_8962);
and U9199 (N_9199,N_8978,N_8778);
or U9200 (N_9200,N_8913,N_8942);
nand U9201 (N_9201,N_8814,N_8908);
or U9202 (N_9202,N_8841,N_8981);
and U9203 (N_9203,N_8978,N_8996);
or U9204 (N_9204,N_8821,N_8901);
nand U9205 (N_9205,N_8949,N_8789);
and U9206 (N_9206,N_8757,N_8853);
or U9207 (N_9207,N_8774,N_8930);
nor U9208 (N_9208,N_8752,N_8751);
and U9209 (N_9209,N_8881,N_8821);
xnor U9210 (N_9210,N_8811,N_8955);
or U9211 (N_9211,N_8921,N_8764);
xnor U9212 (N_9212,N_8784,N_8811);
xor U9213 (N_9213,N_8896,N_8832);
nand U9214 (N_9214,N_8835,N_8998);
and U9215 (N_9215,N_8855,N_8800);
or U9216 (N_9216,N_8752,N_8812);
xnor U9217 (N_9217,N_8871,N_8861);
nor U9218 (N_9218,N_8784,N_8826);
nor U9219 (N_9219,N_8836,N_8885);
or U9220 (N_9220,N_8917,N_8776);
nor U9221 (N_9221,N_8910,N_8752);
nand U9222 (N_9222,N_8762,N_8814);
or U9223 (N_9223,N_8956,N_8795);
nor U9224 (N_9224,N_8807,N_8977);
nand U9225 (N_9225,N_8812,N_8891);
and U9226 (N_9226,N_8824,N_8855);
and U9227 (N_9227,N_8839,N_8982);
or U9228 (N_9228,N_8868,N_8844);
and U9229 (N_9229,N_8752,N_8918);
and U9230 (N_9230,N_8873,N_8924);
and U9231 (N_9231,N_8873,N_8909);
or U9232 (N_9232,N_8800,N_8987);
or U9233 (N_9233,N_8986,N_8834);
xnor U9234 (N_9234,N_8942,N_8862);
nor U9235 (N_9235,N_8937,N_8834);
nor U9236 (N_9236,N_8882,N_8754);
and U9237 (N_9237,N_8837,N_8804);
nand U9238 (N_9238,N_8940,N_8929);
or U9239 (N_9239,N_8861,N_8777);
and U9240 (N_9240,N_8940,N_8941);
nor U9241 (N_9241,N_8906,N_8819);
xor U9242 (N_9242,N_8905,N_8953);
nand U9243 (N_9243,N_8783,N_8811);
nand U9244 (N_9244,N_8856,N_8796);
and U9245 (N_9245,N_8903,N_8994);
or U9246 (N_9246,N_8828,N_8802);
xnor U9247 (N_9247,N_8875,N_8874);
and U9248 (N_9248,N_8886,N_8942);
nand U9249 (N_9249,N_8965,N_8977);
nand U9250 (N_9250,N_9165,N_9120);
and U9251 (N_9251,N_9024,N_9012);
nand U9252 (N_9252,N_9002,N_9137);
nand U9253 (N_9253,N_9074,N_9243);
nor U9254 (N_9254,N_9086,N_9046);
or U9255 (N_9255,N_9192,N_9108);
nor U9256 (N_9256,N_9173,N_9064);
or U9257 (N_9257,N_9031,N_9244);
xnor U9258 (N_9258,N_9090,N_9197);
and U9259 (N_9259,N_9205,N_9220);
nor U9260 (N_9260,N_9154,N_9195);
nand U9261 (N_9261,N_9021,N_9101);
nor U9262 (N_9262,N_9214,N_9081);
nor U9263 (N_9263,N_9163,N_9223);
nor U9264 (N_9264,N_9034,N_9210);
or U9265 (N_9265,N_9056,N_9040);
or U9266 (N_9266,N_9150,N_9116);
nor U9267 (N_9267,N_9060,N_9174);
nand U9268 (N_9268,N_9077,N_9201);
and U9269 (N_9269,N_9067,N_9114);
nand U9270 (N_9270,N_9122,N_9038);
or U9271 (N_9271,N_9198,N_9117);
xor U9272 (N_9272,N_9048,N_9093);
xor U9273 (N_9273,N_9027,N_9143);
nand U9274 (N_9274,N_9176,N_9148);
nor U9275 (N_9275,N_9115,N_9153);
nand U9276 (N_9276,N_9014,N_9099);
xor U9277 (N_9277,N_9129,N_9005);
nand U9278 (N_9278,N_9080,N_9149);
and U9279 (N_9279,N_9042,N_9218);
or U9280 (N_9280,N_9190,N_9248);
nand U9281 (N_9281,N_9249,N_9051);
and U9282 (N_9282,N_9194,N_9052);
or U9283 (N_9283,N_9206,N_9239);
xnor U9284 (N_9284,N_9202,N_9241);
nand U9285 (N_9285,N_9008,N_9219);
nor U9286 (N_9286,N_9082,N_9016);
nor U9287 (N_9287,N_9083,N_9096);
and U9288 (N_9288,N_9144,N_9097);
or U9289 (N_9289,N_9215,N_9134);
and U9290 (N_9290,N_9030,N_9025);
or U9291 (N_9291,N_9098,N_9123);
or U9292 (N_9292,N_9217,N_9212);
xor U9293 (N_9293,N_9170,N_9085);
and U9294 (N_9294,N_9103,N_9004);
xor U9295 (N_9295,N_9247,N_9124);
and U9296 (N_9296,N_9141,N_9213);
nor U9297 (N_9297,N_9135,N_9053);
nand U9298 (N_9298,N_9169,N_9235);
xor U9299 (N_9299,N_9015,N_9232);
xor U9300 (N_9300,N_9068,N_9199);
nor U9301 (N_9301,N_9032,N_9111);
nor U9302 (N_9302,N_9233,N_9185);
nand U9303 (N_9303,N_9036,N_9062);
or U9304 (N_9304,N_9230,N_9227);
nand U9305 (N_9305,N_9009,N_9125);
xor U9306 (N_9306,N_9196,N_9171);
and U9307 (N_9307,N_9087,N_9224);
nand U9308 (N_9308,N_9152,N_9079);
nand U9309 (N_9309,N_9119,N_9059);
nor U9310 (N_9310,N_9172,N_9006);
nand U9311 (N_9311,N_9045,N_9229);
nand U9312 (N_9312,N_9022,N_9092);
or U9313 (N_9313,N_9130,N_9066);
or U9314 (N_9314,N_9164,N_9076);
xnor U9315 (N_9315,N_9069,N_9179);
nand U9316 (N_9316,N_9140,N_9033);
or U9317 (N_9317,N_9007,N_9011);
nor U9318 (N_9318,N_9017,N_9238);
and U9319 (N_9319,N_9072,N_9216);
or U9320 (N_9320,N_9094,N_9175);
nor U9321 (N_9321,N_9246,N_9181);
and U9322 (N_9322,N_9095,N_9049);
xor U9323 (N_9323,N_9146,N_9110);
nand U9324 (N_9324,N_9157,N_9139);
or U9325 (N_9325,N_9001,N_9167);
xnor U9326 (N_9326,N_9209,N_9204);
nor U9327 (N_9327,N_9073,N_9102);
or U9328 (N_9328,N_9188,N_9028);
or U9329 (N_9329,N_9100,N_9225);
and U9330 (N_9330,N_9180,N_9003);
xor U9331 (N_9331,N_9211,N_9142);
nand U9332 (N_9332,N_9193,N_9065);
or U9333 (N_9333,N_9156,N_9055);
nor U9334 (N_9334,N_9236,N_9020);
xor U9335 (N_9335,N_9151,N_9105);
nand U9336 (N_9336,N_9104,N_9078);
nand U9337 (N_9337,N_9183,N_9121);
or U9338 (N_9338,N_9231,N_9161);
and U9339 (N_9339,N_9162,N_9043);
and U9340 (N_9340,N_9226,N_9178);
xnor U9341 (N_9341,N_9088,N_9228);
and U9342 (N_9342,N_9189,N_9184);
xnor U9343 (N_9343,N_9132,N_9245);
xnor U9344 (N_9344,N_9159,N_9013);
nand U9345 (N_9345,N_9061,N_9010);
or U9346 (N_9346,N_9138,N_9145);
xor U9347 (N_9347,N_9208,N_9063);
or U9348 (N_9348,N_9221,N_9133);
xnor U9349 (N_9349,N_9041,N_9158);
or U9350 (N_9350,N_9075,N_9019);
xor U9351 (N_9351,N_9037,N_9187);
xor U9352 (N_9352,N_9029,N_9240);
nand U9353 (N_9353,N_9191,N_9054);
and U9354 (N_9354,N_9109,N_9106);
nor U9355 (N_9355,N_9147,N_9160);
nor U9356 (N_9356,N_9018,N_9237);
xnor U9357 (N_9357,N_9182,N_9177);
xor U9358 (N_9358,N_9186,N_9155);
nand U9359 (N_9359,N_9071,N_9070);
xor U9360 (N_9360,N_9131,N_9089);
and U9361 (N_9361,N_9136,N_9127);
xnor U9362 (N_9362,N_9057,N_9222);
xor U9363 (N_9363,N_9242,N_9026);
nand U9364 (N_9364,N_9168,N_9050);
and U9365 (N_9365,N_9112,N_9091);
xnor U9366 (N_9366,N_9126,N_9044);
or U9367 (N_9367,N_9113,N_9207);
xor U9368 (N_9368,N_9039,N_9084);
nor U9369 (N_9369,N_9234,N_9023);
nand U9370 (N_9370,N_9000,N_9107);
and U9371 (N_9371,N_9203,N_9118);
xor U9372 (N_9372,N_9058,N_9128);
xnor U9373 (N_9373,N_9035,N_9166);
nand U9374 (N_9374,N_9200,N_9047);
or U9375 (N_9375,N_9119,N_9184);
nand U9376 (N_9376,N_9027,N_9185);
or U9377 (N_9377,N_9227,N_9115);
nand U9378 (N_9378,N_9249,N_9176);
nand U9379 (N_9379,N_9191,N_9100);
xor U9380 (N_9380,N_9120,N_9056);
or U9381 (N_9381,N_9082,N_9067);
nand U9382 (N_9382,N_9148,N_9023);
or U9383 (N_9383,N_9188,N_9150);
nand U9384 (N_9384,N_9239,N_9114);
or U9385 (N_9385,N_9171,N_9018);
xnor U9386 (N_9386,N_9015,N_9034);
xnor U9387 (N_9387,N_9085,N_9078);
nand U9388 (N_9388,N_9083,N_9221);
xnor U9389 (N_9389,N_9187,N_9046);
nand U9390 (N_9390,N_9220,N_9248);
nor U9391 (N_9391,N_9246,N_9045);
and U9392 (N_9392,N_9083,N_9077);
and U9393 (N_9393,N_9190,N_9160);
or U9394 (N_9394,N_9069,N_9086);
nand U9395 (N_9395,N_9196,N_9080);
xor U9396 (N_9396,N_9110,N_9013);
nor U9397 (N_9397,N_9161,N_9214);
nor U9398 (N_9398,N_9003,N_9054);
and U9399 (N_9399,N_9104,N_9145);
xnor U9400 (N_9400,N_9223,N_9249);
nor U9401 (N_9401,N_9195,N_9059);
xor U9402 (N_9402,N_9080,N_9110);
nand U9403 (N_9403,N_9027,N_9125);
and U9404 (N_9404,N_9090,N_9005);
or U9405 (N_9405,N_9102,N_9192);
nand U9406 (N_9406,N_9233,N_9119);
and U9407 (N_9407,N_9024,N_9098);
nor U9408 (N_9408,N_9054,N_9098);
nor U9409 (N_9409,N_9139,N_9085);
or U9410 (N_9410,N_9128,N_9169);
nor U9411 (N_9411,N_9146,N_9142);
nor U9412 (N_9412,N_9118,N_9003);
xnor U9413 (N_9413,N_9209,N_9229);
nand U9414 (N_9414,N_9128,N_9122);
xor U9415 (N_9415,N_9208,N_9045);
and U9416 (N_9416,N_9049,N_9176);
nor U9417 (N_9417,N_9026,N_9128);
xor U9418 (N_9418,N_9101,N_9019);
or U9419 (N_9419,N_9104,N_9138);
and U9420 (N_9420,N_9038,N_9156);
and U9421 (N_9421,N_9204,N_9171);
nor U9422 (N_9422,N_9172,N_9228);
nand U9423 (N_9423,N_9082,N_9050);
xnor U9424 (N_9424,N_9003,N_9213);
nor U9425 (N_9425,N_9050,N_9034);
nand U9426 (N_9426,N_9065,N_9123);
xnor U9427 (N_9427,N_9052,N_9201);
nor U9428 (N_9428,N_9247,N_9021);
nor U9429 (N_9429,N_9104,N_9214);
and U9430 (N_9430,N_9163,N_9184);
nor U9431 (N_9431,N_9005,N_9052);
nand U9432 (N_9432,N_9148,N_9242);
xor U9433 (N_9433,N_9014,N_9131);
nor U9434 (N_9434,N_9095,N_9118);
or U9435 (N_9435,N_9132,N_9045);
nand U9436 (N_9436,N_9210,N_9187);
nand U9437 (N_9437,N_9226,N_9030);
nand U9438 (N_9438,N_9066,N_9194);
xor U9439 (N_9439,N_9010,N_9200);
nor U9440 (N_9440,N_9069,N_9243);
and U9441 (N_9441,N_9108,N_9121);
xnor U9442 (N_9442,N_9198,N_9214);
nand U9443 (N_9443,N_9200,N_9224);
or U9444 (N_9444,N_9203,N_9208);
nand U9445 (N_9445,N_9178,N_9026);
and U9446 (N_9446,N_9103,N_9215);
or U9447 (N_9447,N_9142,N_9220);
nand U9448 (N_9448,N_9008,N_9203);
xnor U9449 (N_9449,N_9040,N_9110);
xnor U9450 (N_9450,N_9249,N_9239);
nand U9451 (N_9451,N_9042,N_9099);
and U9452 (N_9452,N_9099,N_9194);
nor U9453 (N_9453,N_9208,N_9151);
xor U9454 (N_9454,N_9085,N_9233);
xor U9455 (N_9455,N_9120,N_9051);
or U9456 (N_9456,N_9219,N_9016);
xor U9457 (N_9457,N_9209,N_9041);
xnor U9458 (N_9458,N_9175,N_9079);
nand U9459 (N_9459,N_9131,N_9174);
and U9460 (N_9460,N_9162,N_9207);
xnor U9461 (N_9461,N_9155,N_9249);
or U9462 (N_9462,N_9069,N_9195);
and U9463 (N_9463,N_9208,N_9011);
and U9464 (N_9464,N_9015,N_9027);
and U9465 (N_9465,N_9154,N_9124);
or U9466 (N_9466,N_9092,N_9103);
nand U9467 (N_9467,N_9214,N_9190);
nand U9468 (N_9468,N_9024,N_9185);
nor U9469 (N_9469,N_9181,N_9051);
nand U9470 (N_9470,N_9030,N_9176);
xor U9471 (N_9471,N_9211,N_9205);
or U9472 (N_9472,N_9083,N_9049);
and U9473 (N_9473,N_9000,N_9184);
or U9474 (N_9474,N_9065,N_9196);
xnor U9475 (N_9475,N_9103,N_9245);
or U9476 (N_9476,N_9117,N_9109);
or U9477 (N_9477,N_9116,N_9065);
nor U9478 (N_9478,N_9028,N_9238);
xor U9479 (N_9479,N_9136,N_9173);
or U9480 (N_9480,N_9050,N_9183);
and U9481 (N_9481,N_9055,N_9033);
xnor U9482 (N_9482,N_9158,N_9148);
nand U9483 (N_9483,N_9160,N_9181);
xnor U9484 (N_9484,N_9198,N_9226);
nor U9485 (N_9485,N_9081,N_9161);
nor U9486 (N_9486,N_9016,N_9065);
and U9487 (N_9487,N_9243,N_9137);
or U9488 (N_9488,N_9027,N_9074);
nand U9489 (N_9489,N_9183,N_9082);
nand U9490 (N_9490,N_9232,N_9217);
nand U9491 (N_9491,N_9141,N_9102);
or U9492 (N_9492,N_9038,N_9213);
and U9493 (N_9493,N_9199,N_9094);
nor U9494 (N_9494,N_9034,N_9012);
xor U9495 (N_9495,N_9183,N_9163);
xor U9496 (N_9496,N_9119,N_9081);
and U9497 (N_9497,N_9225,N_9126);
or U9498 (N_9498,N_9249,N_9010);
xor U9499 (N_9499,N_9205,N_9005);
nand U9500 (N_9500,N_9286,N_9491);
or U9501 (N_9501,N_9282,N_9316);
nand U9502 (N_9502,N_9329,N_9368);
and U9503 (N_9503,N_9362,N_9303);
nand U9504 (N_9504,N_9292,N_9348);
xor U9505 (N_9505,N_9455,N_9261);
nand U9506 (N_9506,N_9379,N_9407);
nor U9507 (N_9507,N_9410,N_9294);
nor U9508 (N_9508,N_9440,N_9394);
or U9509 (N_9509,N_9464,N_9287);
nand U9510 (N_9510,N_9473,N_9417);
or U9511 (N_9511,N_9443,N_9357);
and U9512 (N_9512,N_9398,N_9382);
nand U9513 (N_9513,N_9301,N_9263);
or U9514 (N_9514,N_9408,N_9343);
nand U9515 (N_9515,N_9428,N_9274);
or U9516 (N_9516,N_9460,N_9389);
and U9517 (N_9517,N_9290,N_9265);
nand U9518 (N_9518,N_9314,N_9465);
or U9519 (N_9519,N_9461,N_9317);
or U9520 (N_9520,N_9497,N_9436);
xor U9521 (N_9521,N_9418,N_9441);
nand U9522 (N_9522,N_9421,N_9453);
and U9523 (N_9523,N_9470,N_9479);
or U9524 (N_9524,N_9431,N_9383);
or U9525 (N_9525,N_9325,N_9323);
or U9526 (N_9526,N_9445,N_9340);
nor U9527 (N_9527,N_9385,N_9254);
and U9528 (N_9528,N_9486,N_9406);
nand U9529 (N_9529,N_9264,N_9331);
or U9530 (N_9530,N_9482,N_9356);
xor U9531 (N_9531,N_9283,N_9289);
nor U9532 (N_9532,N_9487,N_9285);
nor U9533 (N_9533,N_9377,N_9442);
or U9534 (N_9534,N_9412,N_9402);
or U9535 (N_9535,N_9277,N_9432);
or U9536 (N_9536,N_9485,N_9349);
nand U9537 (N_9537,N_9475,N_9496);
xor U9538 (N_9538,N_9457,N_9435);
nor U9539 (N_9539,N_9478,N_9392);
nand U9540 (N_9540,N_9257,N_9424);
nand U9541 (N_9541,N_9373,N_9448);
and U9542 (N_9542,N_9269,N_9336);
xor U9543 (N_9543,N_9481,N_9313);
and U9544 (N_9544,N_9419,N_9439);
xnor U9545 (N_9545,N_9327,N_9293);
or U9546 (N_9546,N_9492,N_9366);
or U9547 (N_9547,N_9409,N_9344);
and U9548 (N_9548,N_9321,N_9312);
and U9549 (N_9549,N_9401,N_9476);
nand U9550 (N_9550,N_9469,N_9472);
or U9551 (N_9551,N_9271,N_9291);
xor U9552 (N_9552,N_9498,N_9463);
xor U9553 (N_9553,N_9365,N_9395);
and U9554 (N_9554,N_9280,N_9420);
and U9555 (N_9555,N_9466,N_9422);
nand U9556 (N_9556,N_9459,N_9309);
nand U9557 (N_9557,N_9360,N_9388);
nor U9558 (N_9558,N_9296,N_9376);
xnor U9559 (N_9559,N_9295,N_9468);
xor U9560 (N_9560,N_9370,N_9405);
or U9561 (N_9561,N_9251,N_9335);
xnor U9562 (N_9562,N_9495,N_9477);
or U9563 (N_9563,N_9452,N_9353);
xor U9564 (N_9564,N_9429,N_9415);
and U9565 (N_9565,N_9299,N_9446);
or U9566 (N_9566,N_9259,N_9404);
nor U9567 (N_9567,N_9350,N_9328);
or U9568 (N_9568,N_9427,N_9268);
nor U9569 (N_9569,N_9381,N_9437);
and U9570 (N_9570,N_9260,N_9449);
nand U9571 (N_9571,N_9266,N_9267);
or U9572 (N_9572,N_9480,N_9341);
nor U9573 (N_9573,N_9387,N_9414);
and U9574 (N_9574,N_9272,N_9494);
and U9575 (N_9575,N_9255,N_9337);
or U9576 (N_9576,N_9275,N_9338);
xnor U9577 (N_9577,N_9430,N_9311);
nand U9578 (N_9578,N_9345,N_9324);
or U9579 (N_9579,N_9330,N_9273);
nor U9580 (N_9580,N_9456,N_9433);
nand U9581 (N_9581,N_9367,N_9450);
xor U9582 (N_9582,N_9444,N_9484);
and U9583 (N_9583,N_9396,N_9393);
nor U9584 (N_9584,N_9426,N_9397);
and U9585 (N_9585,N_9333,N_9258);
nand U9586 (N_9586,N_9454,N_9281);
or U9587 (N_9587,N_9342,N_9315);
xnor U9588 (N_9588,N_9352,N_9298);
nand U9589 (N_9589,N_9326,N_9347);
nor U9590 (N_9590,N_9320,N_9451);
xor U9591 (N_9591,N_9363,N_9369);
nand U9592 (N_9592,N_9302,N_9332);
nor U9593 (N_9593,N_9447,N_9334);
nor U9594 (N_9594,N_9305,N_9413);
nand U9595 (N_9595,N_9284,N_9391);
nor U9596 (N_9596,N_9471,N_9270);
xnor U9597 (N_9597,N_9493,N_9416);
nand U9598 (N_9598,N_9399,N_9288);
or U9599 (N_9599,N_9310,N_9339);
or U9600 (N_9600,N_9386,N_9278);
nor U9601 (N_9601,N_9364,N_9488);
and U9602 (N_9602,N_9279,N_9355);
and U9603 (N_9603,N_9374,N_9318);
xor U9604 (N_9604,N_9483,N_9262);
or U9605 (N_9605,N_9423,N_9308);
nand U9606 (N_9606,N_9384,N_9400);
or U9607 (N_9607,N_9375,N_9489);
xor U9608 (N_9608,N_9306,N_9276);
or U9609 (N_9609,N_9256,N_9462);
nand U9610 (N_9610,N_9354,N_9297);
nor U9611 (N_9611,N_9300,N_9474);
nand U9612 (N_9612,N_9378,N_9351);
and U9613 (N_9613,N_9411,N_9490);
and U9614 (N_9614,N_9458,N_9346);
xor U9615 (N_9615,N_9319,N_9434);
and U9616 (N_9616,N_9403,N_9372);
xor U9617 (N_9617,N_9425,N_9371);
nand U9618 (N_9618,N_9438,N_9380);
nand U9619 (N_9619,N_9499,N_9250);
nand U9620 (N_9620,N_9467,N_9304);
and U9621 (N_9621,N_9361,N_9358);
or U9622 (N_9622,N_9359,N_9390);
or U9623 (N_9623,N_9322,N_9253);
nand U9624 (N_9624,N_9307,N_9252);
or U9625 (N_9625,N_9286,N_9327);
xnor U9626 (N_9626,N_9362,N_9250);
xor U9627 (N_9627,N_9304,N_9431);
nand U9628 (N_9628,N_9436,N_9454);
nor U9629 (N_9629,N_9317,N_9365);
or U9630 (N_9630,N_9397,N_9399);
nor U9631 (N_9631,N_9416,N_9376);
xnor U9632 (N_9632,N_9266,N_9311);
and U9633 (N_9633,N_9297,N_9430);
and U9634 (N_9634,N_9440,N_9391);
and U9635 (N_9635,N_9321,N_9287);
or U9636 (N_9636,N_9406,N_9366);
nand U9637 (N_9637,N_9391,N_9304);
and U9638 (N_9638,N_9298,N_9465);
nand U9639 (N_9639,N_9324,N_9461);
nor U9640 (N_9640,N_9365,N_9335);
xnor U9641 (N_9641,N_9496,N_9368);
or U9642 (N_9642,N_9270,N_9305);
and U9643 (N_9643,N_9440,N_9251);
or U9644 (N_9644,N_9303,N_9493);
and U9645 (N_9645,N_9281,N_9437);
nand U9646 (N_9646,N_9433,N_9255);
nand U9647 (N_9647,N_9323,N_9400);
or U9648 (N_9648,N_9473,N_9343);
nor U9649 (N_9649,N_9267,N_9362);
nand U9650 (N_9650,N_9261,N_9259);
and U9651 (N_9651,N_9468,N_9449);
xnor U9652 (N_9652,N_9318,N_9416);
and U9653 (N_9653,N_9316,N_9371);
nor U9654 (N_9654,N_9296,N_9335);
xnor U9655 (N_9655,N_9331,N_9454);
xnor U9656 (N_9656,N_9414,N_9484);
or U9657 (N_9657,N_9487,N_9261);
nor U9658 (N_9658,N_9430,N_9355);
xor U9659 (N_9659,N_9406,N_9271);
xor U9660 (N_9660,N_9338,N_9323);
nand U9661 (N_9661,N_9253,N_9442);
nand U9662 (N_9662,N_9495,N_9266);
nand U9663 (N_9663,N_9288,N_9440);
nand U9664 (N_9664,N_9419,N_9361);
nand U9665 (N_9665,N_9368,N_9487);
nor U9666 (N_9666,N_9256,N_9421);
and U9667 (N_9667,N_9426,N_9412);
and U9668 (N_9668,N_9290,N_9316);
nor U9669 (N_9669,N_9370,N_9254);
nor U9670 (N_9670,N_9261,N_9266);
or U9671 (N_9671,N_9366,N_9465);
xnor U9672 (N_9672,N_9427,N_9482);
nand U9673 (N_9673,N_9292,N_9428);
xnor U9674 (N_9674,N_9334,N_9422);
and U9675 (N_9675,N_9281,N_9410);
xnor U9676 (N_9676,N_9495,N_9268);
or U9677 (N_9677,N_9373,N_9314);
or U9678 (N_9678,N_9429,N_9266);
xnor U9679 (N_9679,N_9424,N_9322);
xor U9680 (N_9680,N_9332,N_9494);
nor U9681 (N_9681,N_9331,N_9312);
xnor U9682 (N_9682,N_9385,N_9456);
nand U9683 (N_9683,N_9456,N_9333);
or U9684 (N_9684,N_9252,N_9387);
nand U9685 (N_9685,N_9251,N_9272);
xnor U9686 (N_9686,N_9346,N_9284);
and U9687 (N_9687,N_9258,N_9283);
nand U9688 (N_9688,N_9467,N_9374);
and U9689 (N_9689,N_9450,N_9374);
and U9690 (N_9690,N_9269,N_9353);
or U9691 (N_9691,N_9262,N_9390);
and U9692 (N_9692,N_9315,N_9458);
nand U9693 (N_9693,N_9260,N_9372);
nor U9694 (N_9694,N_9269,N_9251);
or U9695 (N_9695,N_9404,N_9330);
and U9696 (N_9696,N_9257,N_9413);
xor U9697 (N_9697,N_9395,N_9337);
nand U9698 (N_9698,N_9381,N_9408);
or U9699 (N_9699,N_9448,N_9377);
nor U9700 (N_9700,N_9444,N_9273);
xnor U9701 (N_9701,N_9495,N_9436);
nor U9702 (N_9702,N_9326,N_9382);
and U9703 (N_9703,N_9300,N_9483);
nor U9704 (N_9704,N_9357,N_9430);
and U9705 (N_9705,N_9278,N_9413);
xor U9706 (N_9706,N_9281,N_9418);
xor U9707 (N_9707,N_9297,N_9285);
xnor U9708 (N_9708,N_9361,N_9372);
nand U9709 (N_9709,N_9456,N_9254);
nor U9710 (N_9710,N_9365,N_9349);
xnor U9711 (N_9711,N_9362,N_9456);
nand U9712 (N_9712,N_9495,N_9311);
or U9713 (N_9713,N_9427,N_9344);
and U9714 (N_9714,N_9299,N_9383);
nand U9715 (N_9715,N_9455,N_9309);
or U9716 (N_9716,N_9305,N_9299);
xnor U9717 (N_9717,N_9273,N_9437);
nor U9718 (N_9718,N_9259,N_9445);
nand U9719 (N_9719,N_9394,N_9396);
xnor U9720 (N_9720,N_9493,N_9300);
and U9721 (N_9721,N_9479,N_9414);
xnor U9722 (N_9722,N_9380,N_9461);
or U9723 (N_9723,N_9402,N_9293);
nand U9724 (N_9724,N_9455,N_9454);
and U9725 (N_9725,N_9302,N_9445);
and U9726 (N_9726,N_9494,N_9486);
and U9727 (N_9727,N_9286,N_9268);
or U9728 (N_9728,N_9468,N_9338);
xor U9729 (N_9729,N_9360,N_9400);
nor U9730 (N_9730,N_9484,N_9261);
nand U9731 (N_9731,N_9353,N_9492);
nor U9732 (N_9732,N_9359,N_9314);
and U9733 (N_9733,N_9364,N_9415);
nand U9734 (N_9734,N_9432,N_9420);
nor U9735 (N_9735,N_9431,N_9305);
and U9736 (N_9736,N_9386,N_9289);
and U9737 (N_9737,N_9252,N_9346);
and U9738 (N_9738,N_9418,N_9268);
or U9739 (N_9739,N_9316,N_9254);
or U9740 (N_9740,N_9299,N_9314);
or U9741 (N_9741,N_9282,N_9367);
and U9742 (N_9742,N_9293,N_9480);
xnor U9743 (N_9743,N_9491,N_9399);
nor U9744 (N_9744,N_9263,N_9322);
nand U9745 (N_9745,N_9326,N_9427);
or U9746 (N_9746,N_9284,N_9339);
and U9747 (N_9747,N_9379,N_9413);
nand U9748 (N_9748,N_9416,N_9362);
nor U9749 (N_9749,N_9380,N_9354);
xor U9750 (N_9750,N_9737,N_9500);
nand U9751 (N_9751,N_9725,N_9708);
nor U9752 (N_9752,N_9698,N_9501);
nor U9753 (N_9753,N_9513,N_9676);
nor U9754 (N_9754,N_9514,N_9535);
and U9755 (N_9755,N_9591,N_9522);
xnor U9756 (N_9756,N_9570,N_9610);
xor U9757 (N_9757,N_9504,N_9686);
xor U9758 (N_9758,N_9672,N_9696);
nand U9759 (N_9759,N_9553,N_9651);
xor U9760 (N_9760,N_9619,N_9697);
nor U9761 (N_9761,N_9705,N_9604);
nor U9762 (N_9762,N_9681,N_9679);
and U9763 (N_9763,N_9709,N_9730);
nand U9764 (N_9764,N_9509,N_9541);
and U9765 (N_9765,N_9726,N_9638);
nand U9766 (N_9766,N_9569,N_9673);
nor U9767 (N_9767,N_9559,N_9617);
or U9768 (N_9768,N_9586,N_9719);
and U9769 (N_9769,N_9689,N_9624);
or U9770 (N_9770,N_9675,N_9585);
nor U9771 (N_9771,N_9680,N_9615);
nand U9772 (N_9772,N_9685,N_9526);
nand U9773 (N_9773,N_9718,N_9732);
or U9774 (N_9774,N_9688,N_9506);
nand U9775 (N_9775,N_9613,N_9543);
nor U9776 (N_9776,N_9712,N_9614);
nor U9777 (N_9777,N_9592,N_9601);
nor U9778 (N_9778,N_9656,N_9555);
or U9779 (N_9779,N_9580,N_9652);
xor U9780 (N_9780,N_9665,N_9744);
xnor U9781 (N_9781,N_9561,N_9520);
or U9782 (N_9782,N_9551,N_9505);
nor U9783 (N_9783,N_9529,N_9578);
and U9784 (N_9784,N_9663,N_9702);
and U9785 (N_9785,N_9516,N_9723);
xor U9786 (N_9786,N_9627,N_9538);
nand U9787 (N_9787,N_9695,N_9508);
nor U9788 (N_9788,N_9557,N_9722);
xor U9789 (N_9789,N_9565,N_9525);
nand U9790 (N_9790,N_9710,N_9666);
or U9791 (N_9791,N_9518,N_9727);
nand U9792 (N_9792,N_9671,N_9734);
or U9793 (N_9793,N_9667,N_9622);
and U9794 (N_9794,N_9691,N_9662);
nand U9795 (N_9795,N_9632,N_9593);
and U9796 (N_9796,N_9620,N_9634);
xor U9797 (N_9797,N_9560,N_9558);
xnor U9798 (N_9798,N_9524,N_9531);
xnor U9799 (N_9799,N_9660,N_9661);
and U9800 (N_9800,N_9637,N_9678);
xnor U9801 (N_9801,N_9556,N_9720);
nand U9802 (N_9802,N_9628,N_9519);
nor U9803 (N_9803,N_9684,N_9621);
and U9804 (N_9804,N_9567,N_9715);
nor U9805 (N_9805,N_9546,N_9608);
nor U9806 (N_9806,N_9612,N_9707);
nor U9807 (N_9807,N_9742,N_9544);
or U9808 (N_9808,N_9502,N_9731);
or U9809 (N_9809,N_9640,N_9577);
xor U9810 (N_9810,N_9631,N_9598);
or U9811 (N_9811,N_9517,N_9587);
or U9812 (N_9812,N_9701,N_9668);
nand U9813 (N_9813,N_9515,N_9534);
or U9814 (N_9814,N_9528,N_9674);
xnor U9815 (N_9815,N_9590,N_9741);
nand U9816 (N_9816,N_9735,N_9657);
xnor U9817 (N_9817,N_9611,N_9653);
or U9818 (N_9818,N_9639,N_9711);
or U9819 (N_9819,N_9699,N_9523);
xnor U9820 (N_9820,N_9575,N_9713);
nand U9821 (N_9821,N_9717,N_9700);
nor U9822 (N_9822,N_9616,N_9690);
and U9823 (N_9823,N_9600,N_9602);
nor U9824 (N_9824,N_9564,N_9716);
xnor U9825 (N_9825,N_9747,N_9636);
or U9826 (N_9826,N_9669,N_9582);
nand U9827 (N_9827,N_9579,N_9589);
or U9828 (N_9828,N_9736,N_9644);
xnor U9829 (N_9829,N_9659,N_9706);
or U9830 (N_9830,N_9596,N_9588);
nor U9831 (N_9831,N_9670,N_9568);
or U9832 (N_9832,N_9658,N_9549);
or U9833 (N_9833,N_9703,N_9626);
xor U9834 (N_9834,N_9542,N_9547);
and U9835 (N_9835,N_9566,N_9682);
or U9836 (N_9836,N_9563,N_9635);
nand U9837 (N_9837,N_9704,N_9724);
nor U9838 (N_9838,N_9599,N_9643);
nand U9839 (N_9839,N_9692,N_9654);
nor U9840 (N_9840,N_9650,N_9574);
xor U9841 (N_9841,N_9694,N_9625);
or U9842 (N_9842,N_9687,N_9645);
nor U9843 (N_9843,N_9641,N_9721);
or U9844 (N_9844,N_9739,N_9603);
nor U9845 (N_9845,N_9609,N_9664);
nor U9846 (N_9846,N_9597,N_9746);
nor U9847 (N_9847,N_9536,N_9554);
or U9848 (N_9848,N_9745,N_9594);
xor U9849 (N_9849,N_9507,N_9738);
and U9850 (N_9850,N_9521,N_9527);
and U9851 (N_9851,N_9595,N_9649);
or U9852 (N_9852,N_9552,N_9512);
nor U9853 (N_9853,N_9539,N_9548);
nor U9854 (N_9854,N_9532,N_9729);
or U9855 (N_9855,N_9629,N_9607);
nand U9856 (N_9856,N_9540,N_9584);
nand U9857 (N_9857,N_9573,N_9633);
or U9858 (N_9858,N_9623,N_9683);
nand U9859 (N_9859,N_9605,N_9655);
and U9860 (N_9860,N_9583,N_9503);
nand U9861 (N_9861,N_9572,N_9642);
or U9862 (N_9862,N_9646,N_9545);
or U9863 (N_9863,N_9606,N_9728);
and U9864 (N_9864,N_9714,N_9733);
or U9865 (N_9865,N_9571,N_9562);
or U9866 (N_9866,N_9740,N_9743);
xnor U9867 (N_9867,N_9530,N_9618);
nand U9868 (N_9868,N_9537,N_9647);
nor U9869 (N_9869,N_9748,N_9510);
nor U9870 (N_9870,N_9550,N_9581);
nand U9871 (N_9871,N_9677,N_9511);
nor U9872 (N_9872,N_9648,N_9749);
xor U9873 (N_9873,N_9576,N_9533);
and U9874 (N_9874,N_9630,N_9693);
nand U9875 (N_9875,N_9652,N_9658);
or U9876 (N_9876,N_9626,N_9746);
xnor U9877 (N_9877,N_9562,N_9523);
nand U9878 (N_9878,N_9648,N_9633);
and U9879 (N_9879,N_9548,N_9702);
xnor U9880 (N_9880,N_9569,N_9711);
xor U9881 (N_9881,N_9730,N_9714);
xor U9882 (N_9882,N_9655,N_9595);
xor U9883 (N_9883,N_9621,N_9577);
nor U9884 (N_9884,N_9720,N_9508);
nor U9885 (N_9885,N_9591,N_9607);
and U9886 (N_9886,N_9715,N_9686);
nand U9887 (N_9887,N_9628,N_9556);
nor U9888 (N_9888,N_9536,N_9715);
or U9889 (N_9889,N_9705,N_9622);
nand U9890 (N_9890,N_9673,N_9576);
and U9891 (N_9891,N_9540,N_9537);
xnor U9892 (N_9892,N_9570,N_9672);
nor U9893 (N_9893,N_9545,N_9732);
xnor U9894 (N_9894,N_9560,N_9649);
or U9895 (N_9895,N_9722,N_9702);
or U9896 (N_9896,N_9700,N_9723);
nor U9897 (N_9897,N_9708,N_9647);
or U9898 (N_9898,N_9593,N_9609);
xnor U9899 (N_9899,N_9596,N_9592);
or U9900 (N_9900,N_9597,N_9598);
xnor U9901 (N_9901,N_9610,N_9635);
and U9902 (N_9902,N_9727,N_9689);
nor U9903 (N_9903,N_9655,N_9715);
nor U9904 (N_9904,N_9599,N_9684);
or U9905 (N_9905,N_9505,N_9576);
nor U9906 (N_9906,N_9595,N_9722);
nor U9907 (N_9907,N_9674,N_9613);
or U9908 (N_9908,N_9604,N_9653);
nand U9909 (N_9909,N_9721,N_9741);
or U9910 (N_9910,N_9615,N_9579);
nand U9911 (N_9911,N_9699,N_9721);
xor U9912 (N_9912,N_9610,N_9676);
and U9913 (N_9913,N_9652,N_9615);
and U9914 (N_9914,N_9707,N_9611);
nand U9915 (N_9915,N_9700,N_9650);
xor U9916 (N_9916,N_9663,N_9717);
or U9917 (N_9917,N_9743,N_9745);
nand U9918 (N_9918,N_9562,N_9660);
or U9919 (N_9919,N_9597,N_9678);
nand U9920 (N_9920,N_9685,N_9566);
xnor U9921 (N_9921,N_9625,N_9510);
xnor U9922 (N_9922,N_9721,N_9636);
nand U9923 (N_9923,N_9706,N_9630);
and U9924 (N_9924,N_9593,N_9560);
nand U9925 (N_9925,N_9577,N_9582);
xnor U9926 (N_9926,N_9696,N_9523);
and U9927 (N_9927,N_9598,N_9626);
and U9928 (N_9928,N_9594,N_9542);
nor U9929 (N_9929,N_9657,N_9608);
nand U9930 (N_9930,N_9594,N_9695);
or U9931 (N_9931,N_9621,N_9636);
nor U9932 (N_9932,N_9675,N_9740);
nand U9933 (N_9933,N_9698,N_9592);
nor U9934 (N_9934,N_9550,N_9513);
and U9935 (N_9935,N_9633,N_9651);
or U9936 (N_9936,N_9617,N_9664);
nor U9937 (N_9937,N_9721,N_9737);
nand U9938 (N_9938,N_9644,N_9721);
nor U9939 (N_9939,N_9568,N_9504);
xnor U9940 (N_9940,N_9701,N_9732);
nor U9941 (N_9941,N_9600,N_9503);
nor U9942 (N_9942,N_9580,N_9655);
and U9943 (N_9943,N_9574,N_9577);
and U9944 (N_9944,N_9518,N_9602);
nand U9945 (N_9945,N_9700,N_9571);
nand U9946 (N_9946,N_9642,N_9621);
or U9947 (N_9947,N_9604,N_9605);
or U9948 (N_9948,N_9600,N_9530);
xor U9949 (N_9949,N_9723,N_9535);
nand U9950 (N_9950,N_9586,N_9521);
nor U9951 (N_9951,N_9557,N_9686);
nor U9952 (N_9952,N_9633,N_9660);
or U9953 (N_9953,N_9619,N_9659);
nand U9954 (N_9954,N_9555,N_9652);
nor U9955 (N_9955,N_9584,N_9552);
and U9956 (N_9956,N_9617,N_9745);
and U9957 (N_9957,N_9745,N_9555);
xor U9958 (N_9958,N_9680,N_9670);
and U9959 (N_9959,N_9506,N_9687);
nand U9960 (N_9960,N_9688,N_9541);
or U9961 (N_9961,N_9666,N_9500);
nand U9962 (N_9962,N_9728,N_9642);
nor U9963 (N_9963,N_9675,N_9699);
nand U9964 (N_9964,N_9568,N_9596);
and U9965 (N_9965,N_9595,N_9624);
or U9966 (N_9966,N_9644,N_9620);
nand U9967 (N_9967,N_9572,N_9511);
nor U9968 (N_9968,N_9560,N_9706);
or U9969 (N_9969,N_9582,N_9683);
or U9970 (N_9970,N_9732,N_9680);
and U9971 (N_9971,N_9683,N_9692);
and U9972 (N_9972,N_9723,N_9671);
nor U9973 (N_9973,N_9693,N_9662);
xor U9974 (N_9974,N_9653,N_9721);
and U9975 (N_9975,N_9559,N_9557);
and U9976 (N_9976,N_9659,N_9558);
or U9977 (N_9977,N_9630,N_9738);
and U9978 (N_9978,N_9669,N_9506);
and U9979 (N_9979,N_9584,N_9728);
nor U9980 (N_9980,N_9550,N_9520);
nor U9981 (N_9981,N_9596,N_9590);
or U9982 (N_9982,N_9554,N_9516);
nor U9983 (N_9983,N_9606,N_9556);
or U9984 (N_9984,N_9720,N_9524);
or U9985 (N_9985,N_9564,N_9569);
or U9986 (N_9986,N_9559,N_9589);
and U9987 (N_9987,N_9691,N_9685);
and U9988 (N_9988,N_9530,N_9610);
xor U9989 (N_9989,N_9586,N_9532);
and U9990 (N_9990,N_9651,N_9625);
xor U9991 (N_9991,N_9650,N_9596);
and U9992 (N_9992,N_9721,N_9521);
and U9993 (N_9993,N_9609,N_9728);
and U9994 (N_9994,N_9733,N_9665);
nand U9995 (N_9995,N_9630,N_9502);
nand U9996 (N_9996,N_9715,N_9530);
nand U9997 (N_9997,N_9614,N_9647);
xnor U9998 (N_9998,N_9620,N_9648);
or U9999 (N_9999,N_9606,N_9729);
nor U10000 (N_10000,N_9855,N_9984);
xnor U10001 (N_10001,N_9861,N_9840);
nor U10002 (N_10002,N_9970,N_9874);
nor U10003 (N_10003,N_9974,N_9815);
or U10004 (N_10004,N_9752,N_9863);
or U10005 (N_10005,N_9981,N_9826);
xor U10006 (N_10006,N_9779,N_9844);
nand U10007 (N_10007,N_9813,N_9839);
or U10008 (N_10008,N_9838,N_9817);
nand U10009 (N_10009,N_9912,N_9938);
xor U10010 (N_10010,N_9973,N_9896);
or U10011 (N_10011,N_9765,N_9927);
xor U10012 (N_10012,N_9999,N_9976);
and U10013 (N_10013,N_9866,N_9825);
nand U10014 (N_10014,N_9908,N_9794);
xnor U10015 (N_10015,N_9954,N_9800);
nor U10016 (N_10016,N_9963,N_9919);
xnor U10017 (N_10017,N_9862,N_9795);
and U10018 (N_10018,N_9947,N_9818);
nand U10019 (N_10019,N_9835,N_9906);
and U10020 (N_10020,N_9848,N_9966);
nand U10021 (N_10021,N_9824,N_9916);
and U10022 (N_10022,N_9873,N_9870);
nand U10023 (N_10023,N_9780,N_9771);
or U10024 (N_10024,N_9995,N_9933);
nor U10025 (N_10025,N_9790,N_9997);
nand U10026 (N_10026,N_9860,N_9936);
xnor U10027 (N_10027,N_9992,N_9769);
nor U10028 (N_10028,N_9775,N_9998);
nor U10029 (N_10029,N_9994,N_9853);
nand U10030 (N_10030,N_9903,N_9847);
or U10031 (N_10031,N_9834,N_9975);
or U10032 (N_10032,N_9943,N_9968);
xor U10033 (N_10033,N_9778,N_9909);
or U10034 (N_10034,N_9956,N_9964);
nand U10035 (N_10035,N_9923,N_9996);
and U10036 (N_10036,N_9821,N_9899);
xnor U10037 (N_10037,N_9932,N_9805);
and U10038 (N_10038,N_9878,N_9756);
nand U10039 (N_10039,N_9910,N_9799);
and U10040 (N_10040,N_9952,N_9955);
xor U10041 (N_10041,N_9785,N_9843);
or U10042 (N_10042,N_9776,N_9883);
or U10043 (N_10043,N_9930,N_9961);
xor U10044 (N_10044,N_9922,N_9812);
or U10045 (N_10045,N_9986,N_9935);
nand U10046 (N_10046,N_9792,N_9946);
nand U10047 (N_10047,N_9757,N_9987);
or U10048 (N_10048,N_9833,N_9991);
or U10049 (N_10049,N_9880,N_9753);
xor U10050 (N_10050,N_9877,N_9884);
xnor U10051 (N_10051,N_9811,N_9879);
or U10052 (N_10052,N_9993,N_9772);
nand U10053 (N_10053,N_9828,N_9979);
xnor U10054 (N_10054,N_9900,N_9761);
nor U10055 (N_10055,N_9786,N_9965);
nand U10056 (N_10056,N_9854,N_9888);
and U10057 (N_10057,N_9798,N_9985);
nand U10058 (N_10058,N_9876,N_9777);
and U10059 (N_10059,N_9967,N_9842);
and U10060 (N_10060,N_9750,N_9960);
nor U10061 (N_10061,N_9832,N_9885);
xnor U10062 (N_10062,N_9829,N_9886);
xor U10063 (N_10063,N_9977,N_9934);
nand U10064 (N_10064,N_9945,N_9980);
nand U10065 (N_10065,N_9806,N_9949);
xnor U10066 (N_10066,N_9751,N_9897);
nor U10067 (N_10067,N_9762,N_9841);
nand U10068 (N_10068,N_9783,N_9989);
xor U10069 (N_10069,N_9898,N_9972);
nand U10070 (N_10070,N_9808,N_9809);
xnor U10071 (N_10071,N_9937,N_9957);
xnor U10072 (N_10072,N_9836,N_9882);
nor U10073 (N_10073,N_9755,N_9814);
xnor U10074 (N_10074,N_9871,N_9969);
nor U10075 (N_10075,N_9971,N_9768);
xor U10076 (N_10076,N_9858,N_9929);
nor U10077 (N_10077,N_9770,N_9950);
nor U10078 (N_10078,N_9948,N_9856);
xnor U10079 (N_10079,N_9905,N_9881);
nand U10080 (N_10080,N_9962,N_9774);
xnor U10081 (N_10081,N_9754,N_9941);
nor U10082 (N_10082,N_9924,N_9990);
xor U10083 (N_10083,N_9865,N_9801);
xnor U10084 (N_10084,N_9827,N_9864);
xor U10085 (N_10085,N_9823,N_9958);
nor U10086 (N_10086,N_9837,N_9820);
or U10087 (N_10087,N_9917,N_9891);
nand U10088 (N_10088,N_9890,N_9816);
or U10089 (N_10089,N_9907,N_9920);
or U10090 (N_10090,N_9928,N_9789);
and U10091 (N_10091,N_9849,N_9831);
or U10092 (N_10092,N_9782,N_9819);
nor U10093 (N_10093,N_9781,N_9944);
nor U10094 (N_10094,N_9913,N_9931);
nand U10095 (N_10095,N_9788,N_9807);
nor U10096 (N_10096,N_9857,N_9796);
or U10097 (N_10097,N_9894,N_9988);
and U10098 (N_10098,N_9868,N_9804);
and U10099 (N_10099,N_9982,N_9759);
xor U10100 (N_10100,N_9959,N_9791);
or U10101 (N_10101,N_9850,N_9851);
nand U10102 (N_10102,N_9983,N_9926);
nand U10103 (N_10103,N_9940,N_9915);
or U10104 (N_10104,N_9758,N_9852);
xor U10105 (N_10105,N_9911,N_9803);
nand U10106 (N_10106,N_9869,N_9793);
nand U10107 (N_10107,N_9822,N_9889);
xor U10108 (N_10108,N_9953,N_9978);
xnor U10109 (N_10109,N_9846,N_9810);
xnor U10110 (N_10110,N_9921,N_9887);
or U10111 (N_10111,N_9893,N_9892);
or U10112 (N_10112,N_9859,N_9802);
xnor U10113 (N_10113,N_9875,N_9787);
xor U10114 (N_10114,N_9942,N_9901);
xnor U10115 (N_10115,N_9760,N_9867);
or U10116 (N_10116,N_9914,N_9904);
nand U10117 (N_10117,N_9784,N_9872);
nand U10118 (N_10118,N_9939,N_9918);
and U10119 (N_10119,N_9797,N_9773);
or U10120 (N_10120,N_9767,N_9951);
nor U10121 (N_10121,N_9830,N_9895);
nor U10122 (N_10122,N_9766,N_9764);
xnor U10123 (N_10123,N_9902,N_9845);
nand U10124 (N_10124,N_9925,N_9763);
xnor U10125 (N_10125,N_9965,N_9828);
nor U10126 (N_10126,N_9912,N_9967);
or U10127 (N_10127,N_9923,N_9779);
and U10128 (N_10128,N_9896,N_9800);
nor U10129 (N_10129,N_9955,N_9772);
nand U10130 (N_10130,N_9929,N_9773);
and U10131 (N_10131,N_9846,N_9929);
nand U10132 (N_10132,N_9834,N_9824);
and U10133 (N_10133,N_9769,N_9987);
nor U10134 (N_10134,N_9811,N_9828);
or U10135 (N_10135,N_9908,N_9961);
xnor U10136 (N_10136,N_9924,N_9875);
or U10137 (N_10137,N_9946,N_9843);
nand U10138 (N_10138,N_9906,N_9773);
nand U10139 (N_10139,N_9990,N_9923);
nand U10140 (N_10140,N_9936,N_9996);
and U10141 (N_10141,N_9898,N_9823);
and U10142 (N_10142,N_9916,N_9818);
or U10143 (N_10143,N_9846,N_9849);
xnor U10144 (N_10144,N_9803,N_9750);
or U10145 (N_10145,N_9866,N_9828);
xor U10146 (N_10146,N_9803,N_9753);
nor U10147 (N_10147,N_9895,N_9855);
nand U10148 (N_10148,N_9839,N_9811);
and U10149 (N_10149,N_9810,N_9842);
or U10150 (N_10150,N_9891,N_9953);
or U10151 (N_10151,N_9920,N_9934);
and U10152 (N_10152,N_9963,N_9975);
or U10153 (N_10153,N_9782,N_9901);
nand U10154 (N_10154,N_9845,N_9834);
and U10155 (N_10155,N_9766,N_9928);
nor U10156 (N_10156,N_9858,N_9831);
nor U10157 (N_10157,N_9891,N_9920);
nor U10158 (N_10158,N_9904,N_9910);
and U10159 (N_10159,N_9799,N_9899);
or U10160 (N_10160,N_9817,N_9965);
and U10161 (N_10161,N_9923,N_9934);
nor U10162 (N_10162,N_9752,N_9941);
nor U10163 (N_10163,N_9776,N_9876);
xnor U10164 (N_10164,N_9992,N_9790);
nor U10165 (N_10165,N_9778,N_9884);
or U10166 (N_10166,N_9855,N_9887);
or U10167 (N_10167,N_9893,N_9975);
nand U10168 (N_10168,N_9790,N_9802);
or U10169 (N_10169,N_9912,N_9892);
nor U10170 (N_10170,N_9822,N_9956);
and U10171 (N_10171,N_9990,N_9993);
and U10172 (N_10172,N_9755,N_9820);
nor U10173 (N_10173,N_9818,N_9905);
nand U10174 (N_10174,N_9957,N_9852);
nand U10175 (N_10175,N_9903,N_9785);
and U10176 (N_10176,N_9871,N_9897);
and U10177 (N_10177,N_9953,N_9811);
nor U10178 (N_10178,N_9776,N_9919);
xnor U10179 (N_10179,N_9802,N_9867);
and U10180 (N_10180,N_9899,N_9813);
nand U10181 (N_10181,N_9984,N_9828);
or U10182 (N_10182,N_9988,N_9782);
and U10183 (N_10183,N_9875,N_9911);
or U10184 (N_10184,N_9901,N_9786);
nor U10185 (N_10185,N_9790,N_9814);
and U10186 (N_10186,N_9862,N_9807);
and U10187 (N_10187,N_9824,N_9765);
xnor U10188 (N_10188,N_9923,N_9824);
nor U10189 (N_10189,N_9876,N_9989);
and U10190 (N_10190,N_9812,N_9860);
nor U10191 (N_10191,N_9786,N_9921);
xor U10192 (N_10192,N_9862,N_9819);
nor U10193 (N_10193,N_9781,N_9841);
nor U10194 (N_10194,N_9807,N_9838);
xnor U10195 (N_10195,N_9856,N_9813);
or U10196 (N_10196,N_9791,N_9965);
or U10197 (N_10197,N_9986,N_9857);
nor U10198 (N_10198,N_9815,N_9828);
xnor U10199 (N_10199,N_9840,N_9988);
and U10200 (N_10200,N_9907,N_9755);
nand U10201 (N_10201,N_9962,N_9753);
or U10202 (N_10202,N_9950,N_9941);
nand U10203 (N_10203,N_9805,N_9829);
or U10204 (N_10204,N_9799,N_9940);
or U10205 (N_10205,N_9894,N_9853);
and U10206 (N_10206,N_9872,N_9877);
nor U10207 (N_10207,N_9776,N_9816);
and U10208 (N_10208,N_9913,N_9929);
and U10209 (N_10209,N_9894,N_9847);
xor U10210 (N_10210,N_9987,N_9954);
nor U10211 (N_10211,N_9788,N_9822);
xor U10212 (N_10212,N_9952,N_9916);
nand U10213 (N_10213,N_9985,N_9970);
nand U10214 (N_10214,N_9954,N_9898);
xnor U10215 (N_10215,N_9829,N_9831);
nor U10216 (N_10216,N_9871,N_9901);
nor U10217 (N_10217,N_9765,N_9834);
or U10218 (N_10218,N_9989,N_9937);
xor U10219 (N_10219,N_9935,N_9924);
or U10220 (N_10220,N_9757,N_9863);
and U10221 (N_10221,N_9771,N_9904);
nand U10222 (N_10222,N_9945,N_9920);
xor U10223 (N_10223,N_9968,N_9898);
nor U10224 (N_10224,N_9823,N_9977);
nand U10225 (N_10225,N_9916,N_9898);
nand U10226 (N_10226,N_9904,N_9764);
nand U10227 (N_10227,N_9766,N_9778);
nand U10228 (N_10228,N_9757,N_9808);
nand U10229 (N_10229,N_9778,N_9788);
nand U10230 (N_10230,N_9780,N_9994);
or U10231 (N_10231,N_9938,N_9916);
nor U10232 (N_10232,N_9761,N_9786);
nor U10233 (N_10233,N_9780,N_9986);
xor U10234 (N_10234,N_9987,N_9751);
xnor U10235 (N_10235,N_9967,N_9931);
and U10236 (N_10236,N_9905,N_9847);
xor U10237 (N_10237,N_9899,N_9837);
or U10238 (N_10238,N_9800,N_9964);
nor U10239 (N_10239,N_9944,N_9850);
nor U10240 (N_10240,N_9944,N_9774);
xor U10241 (N_10241,N_9867,N_9821);
or U10242 (N_10242,N_9901,N_9852);
nand U10243 (N_10243,N_9766,N_9946);
nand U10244 (N_10244,N_9892,N_9763);
or U10245 (N_10245,N_9773,N_9852);
and U10246 (N_10246,N_9945,N_9998);
or U10247 (N_10247,N_9804,N_9992);
nor U10248 (N_10248,N_9833,N_9882);
or U10249 (N_10249,N_9931,N_9917);
nand U10250 (N_10250,N_10144,N_10136);
or U10251 (N_10251,N_10199,N_10226);
xor U10252 (N_10252,N_10039,N_10228);
and U10253 (N_10253,N_10145,N_10003);
nor U10254 (N_10254,N_10059,N_10132);
and U10255 (N_10255,N_10211,N_10128);
nor U10256 (N_10256,N_10115,N_10159);
and U10257 (N_10257,N_10109,N_10125);
nor U10258 (N_10258,N_10241,N_10095);
and U10259 (N_10259,N_10158,N_10223);
xor U10260 (N_10260,N_10013,N_10033);
nand U10261 (N_10261,N_10209,N_10058);
xor U10262 (N_10262,N_10204,N_10085);
or U10263 (N_10263,N_10126,N_10134);
nand U10264 (N_10264,N_10164,N_10161);
xor U10265 (N_10265,N_10081,N_10171);
and U10266 (N_10266,N_10230,N_10071);
or U10267 (N_10267,N_10110,N_10190);
and U10268 (N_10268,N_10246,N_10045);
nand U10269 (N_10269,N_10076,N_10247);
and U10270 (N_10270,N_10111,N_10043);
or U10271 (N_10271,N_10133,N_10102);
nor U10272 (N_10272,N_10060,N_10070);
xor U10273 (N_10273,N_10140,N_10001);
nand U10274 (N_10274,N_10052,N_10152);
nor U10275 (N_10275,N_10112,N_10201);
nor U10276 (N_10276,N_10107,N_10062);
nor U10277 (N_10277,N_10038,N_10127);
or U10278 (N_10278,N_10005,N_10222);
and U10279 (N_10279,N_10116,N_10180);
nor U10280 (N_10280,N_10200,N_10146);
xnor U10281 (N_10281,N_10175,N_10177);
nor U10282 (N_10282,N_10023,N_10216);
and U10283 (N_10283,N_10179,N_10196);
and U10284 (N_10284,N_10061,N_10153);
or U10285 (N_10285,N_10031,N_10097);
or U10286 (N_10286,N_10151,N_10220);
nor U10287 (N_10287,N_10096,N_10008);
and U10288 (N_10288,N_10022,N_10026);
or U10289 (N_10289,N_10217,N_10067);
or U10290 (N_10290,N_10227,N_10093);
nand U10291 (N_10291,N_10002,N_10210);
nor U10292 (N_10292,N_10129,N_10068);
xnor U10293 (N_10293,N_10169,N_10162);
and U10294 (N_10294,N_10014,N_10044);
nand U10295 (N_10295,N_10009,N_10206);
nand U10296 (N_10296,N_10123,N_10142);
and U10297 (N_10297,N_10188,N_10057);
and U10298 (N_10298,N_10156,N_10098);
and U10299 (N_10299,N_10173,N_10154);
nor U10300 (N_10300,N_10212,N_10150);
or U10301 (N_10301,N_10007,N_10141);
and U10302 (N_10302,N_10114,N_10147);
nor U10303 (N_10303,N_10019,N_10036);
xor U10304 (N_10304,N_10056,N_10198);
nand U10305 (N_10305,N_10028,N_10080);
or U10306 (N_10306,N_10089,N_10054);
nor U10307 (N_10307,N_10225,N_10163);
nand U10308 (N_10308,N_10103,N_10077);
nor U10309 (N_10309,N_10202,N_10037);
nor U10310 (N_10310,N_10138,N_10051);
and U10311 (N_10311,N_10193,N_10040);
nor U10312 (N_10312,N_10047,N_10078);
and U10313 (N_10313,N_10083,N_10224);
nand U10314 (N_10314,N_10029,N_10063);
xnor U10315 (N_10315,N_10178,N_10122);
or U10316 (N_10316,N_10205,N_10189);
nor U10317 (N_10317,N_10119,N_10203);
or U10318 (N_10318,N_10139,N_10155);
and U10319 (N_10319,N_10035,N_10042);
or U10320 (N_10320,N_10087,N_10207);
nand U10321 (N_10321,N_10243,N_10242);
and U10322 (N_10322,N_10094,N_10011);
nor U10323 (N_10323,N_10176,N_10240);
or U10324 (N_10324,N_10099,N_10239);
or U10325 (N_10325,N_10075,N_10181);
nor U10326 (N_10326,N_10167,N_10249);
and U10327 (N_10327,N_10105,N_10090);
and U10328 (N_10328,N_10234,N_10064);
or U10329 (N_10329,N_10182,N_10018);
nand U10330 (N_10330,N_10048,N_10172);
or U10331 (N_10331,N_10229,N_10106);
nand U10332 (N_10332,N_10012,N_10030);
xor U10333 (N_10333,N_10006,N_10010);
xnor U10334 (N_10334,N_10025,N_10174);
nor U10335 (N_10335,N_10066,N_10192);
nor U10336 (N_10336,N_10084,N_10118);
xor U10337 (N_10337,N_10124,N_10074);
xor U10338 (N_10338,N_10232,N_10131);
and U10339 (N_10339,N_10072,N_10237);
nand U10340 (N_10340,N_10135,N_10184);
xor U10341 (N_10341,N_10000,N_10130);
or U10342 (N_10342,N_10218,N_10065);
and U10343 (N_10343,N_10233,N_10149);
xor U10344 (N_10344,N_10004,N_10166);
xor U10345 (N_10345,N_10137,N_10143);
or U10346 (N_10346,N_10215,N_10214);
and U10347 (N_10347,N_10231,N_10245);
nor U10348 (N_10348,N_10015,N_10027);
and U10349 (N_10349,N_10020,N_10238);
nor U10350 (N_10350,N_10108,N_10055);
nand U10351 (N_10351,N_10236,N_10186);
or U10352 (N_10352,N_10244,N_10016);
xor U10353 (N_10353,N_10092,N_10221);
or U10354 (N_10354,N_10213,N_10165);
nor U10355 (N_10355,N_10121,N_10017);
nor U10356 (N_10356,N_10248,N_10049);
nand U10357 (N_10357,N_10073,N_10160);
xor U10358 (N_10358,N_10148,N_10120);
nor U10359 (N_10359,N_10168,N_10187);
and U10360 (N_10360,N_10091,N_10021);
nor U10361 (N_10361,N_10235,N_10082);
nand U10362 (N_10362,N_10197,N_10104);
nand U10363 (N_10363,N_10069,N_10041);
or U10364 (N_10364,N_10046,N_10113);
and U10365 (N_10365,N_10157,N_10183);
xor U10366 (N_10366,N_10086,N_10024);
nand U10367 (N_10367,N_10208,N_10195);
and U10368 (N_10368,N_10053,N_10032);
xnor U10369 (N_10369,N_10219,N_10050);
or U10370 (N_10370,N_10079,N_10088);
nor U10371 (N_10371,N_10117,N_10185);
nand U10372 (N_10372,N_10034,N_10170);
nor U10373 (N_10373,N_10194,N_10191);
nor U10374 (N_10374,N_10101,N_10100);
xnor U10375 (N_10375,N_10129,N_10028);
and U10376 (N_10376,N_10153,N_10137);
nor U10377 (N_10377,N_10130,N_10115);
nand U10378 (N_10378,N_10080,N_10022);
and U10379 (N_10379,N_10101,N_10099);
or U10380 (N_10380,N_10052,N_10078);
and U10381 (N_10381,N_10018,N_10100);
nand U10382 (N_10382,N_10247,N_10175);
or U10383 (N_10383,N_10094,N_10237);
and U10384 (N_10384,N_10239,N_10166);
nor U10385 (N_10385,N_10226,N_10182);
nor U10386 (N_10386,N_10192,N_10127);
and U10387 (N_10387,N_10112,N_10089);
nor U10388 (N_10388,N_10173,N_10181);
xnor U10389 (N_10389,N_10216,N_10178);
or U10390 (N_10390,N_10171,N_10178);
xor U10391 (N_10391,N_10073,N_10214);
and U10392 (N_10392,N_10235,N_10204);
nand U10393 (N_10393,N_10156,N_10219);
or U10394 (N_10394,N_10175,N_10020);
nand U10395 (N_10395,N_10117,N_10198);
and U10396 (N_10396,N_10002,N_10242);
nand U10397 (N_10397,N_10068,N_10012);
nor U10398 (N_10398,N_10015,N_10110);
and U10399 (N_10399,N_10154,N_10097);
xnor U10400 (N_10400,N_10210,N_10206);
and U10401 (N_10401,N_10024,N_10011);
xor U10402 (N_10402,N_10127,N_10175);
nor U10403 (N_10403,N_10154,N_10011);
nor U10404 (N_10404,N_10246,N_10207);
or U10405 (N_10405,N_10111,N_10205);
nand U10406 (N_10406,N_10151,N_10065);
or U10407 (N_10407,N_10207,N_10076);
xor U10408 (N_10408,N_10105,N_10087);
xor U10409 (N_10409,N_10082,N_10150);
nand U10410 (N_10410,N_10197,N_10023);
or U10411 (N_10411,N_10176,N_10114);
nand U10412 (N_10412,N_10085,N_10039);
nor U10413 (N_10413,N_10038,N_10062);
nand U10414 (N_10414,N_10071,N_10099);
xor U10415 (N_10415,N_10010,N_10114);
nand U10416 (N_10416,N_10005,N_10212);
nand U10417 (N_10417,N_10011,N_10127);
nand U10418 (N_10418,N_10092,N_10074);
or U10419 (N_10419,N_10159,N_10203);
xnor U10420 (N_10420,N_10077,N_10087);
xnor U10421 (N_10421,N_10200,N_10046);
or U10422 (N_10422,N_10079,N_10127);
nand U10423 (N_10423,N_10178,N_10192);
nor U10424 (N_10424,N_10092,N_10089);
nand U10425 (N_10425,N_10130,N_10179);
or U10426 (N_10426,N_10031,N_10054);
nand U10427 (N_10427,N_10058,N_10141);
nor U10428 (N_10428,N_10199,N_10086);
and U10429 (N_10429,N_10147,N_10044);
nand U10430 (N_10430,N_10165,N_10173);
nor U10431 (N_10431,N_10091,N_10121);
nand U10432 (N_10432,N_10159,N_10125);
xor U10433 (N_10433,N_10014,N_10176);
and U10434 (N_10434,N_10233,N_10005);
xor U10435 (N_10435,N_10241,N_10215);
and U10436 (N_10436,N_10143,N_10152);
or U10437 (N_10437,N_10004,N_10170);
xor U10438 (N_10438,N_10243,N_10122);
nor U10439 (N_10439,N_10019,N_10214);
xor U10440 (N_10440,N_10017,N_10108);
nor U10441 (N_10441,N_10154,N_10167);
nor U10442 (N_10442,N_10166,N_10076);
xnor U10443 (N_10443,N_10004,N_10068);
nor U10444 (N_10444,N_10157,N_10172);
and U10445 (N_10445,N_10057,N_10155);
nor U10446 (N_10446,N_10072,N_10222);
nand U10447 (N_10447,N_10132,N_10192);
xor U10448 (N_10448,N_10039,N_10023);
nand U10449 (N_10449,N_10041,N_10159);
or U10450 (N_10450,N_10164,N_10141);
nor U10451 (N_10451,N_10188,N_10161);
nor U10452 (N_10452,N_10101,N_10160);
nor U10453 (N_10453,N_10075,N_10023);
xor U10454 (N_10454,N_10182,N_10107);
or U10455 (N_10455,N_10223,N_10047);
or U10456 (N_10456,N_10212,N_10030);
nor U10457 (N_10457,N_10085,N_10249);
xor U10458 (N_10458,N_10098,N_10001);
nor U10459 (N_10459,N_10127,N_10126);
nand U10460 (N_10460,N_10030,N_10215);
or U10461 (N_10461,N_10174,N_10052);
or U10462 (N_10462,N_10134,N_10211);
nand U10463 (N_10463,N_10220,N_10245);
nor U10464 (N_10464,N_10086,N_10068);
nand U10465 (N_10465,N_10118,N_10124);
and U10466 (N_10466,N_10110,N_10204);
xor U10467 (N_10467,N_10089,N_10166);
nand U10468 (N_10468,N_10198,N_10018);
nor U10469 (N_10469,N_10227,N_10210);
xnor U10470 (N_10470,N_10035,N_10244);
and U10471 (N_10471,N_10097,N_10000);
or U10472 (N_10472,N_10104,N_10169);
or U10473 (N_10473,N_10207,N_10012);
nand U10474 (N_10474,N_10180,N_10027);
and U10475 (N_10475,N_10124,N_10206);
or U10476 (N_10476,N_10177,N_10036);
or U10477 (N_10477,N_10047,N_10236);
nor U10478 (N_10478,N_10022,N_10110);
and U10479 (N_10479,N_10124,N_10014);
nand U10480 (N_10480,N_10006,N_10083);
xor U10481 (N_10481,N_10090,N_10222);
nor U10482 (N_10482,N_10124,N_10121);
nand U10483 (N_10483,N_10222,N_10118);
or U10484 (N_10484,N_10008,N_10047);
or U10485 (N_10485,N_10228,N_10052);
nor U10486 (N_10486,N_10101,N_10102);
or U10487 (N_10487,N_10128,N_10206);
or U10488 (N_10488,N_10070,N_10108);
or U10489 (N_10489,N_10189,N_10217);
and U10490 (N_10490,N_10110,N_10138);
xnor U10491 (N_10491,N_10185,N_10068);
or U10492 (N_10492,N_10022,N_10139);
nor U10493 (N_10493,N_10235,N_10158);
nand U10494 (N_10494,N_10147,N_10182);
nor U10495 (N_10495,N_10156,N_10229);
xor U10496 (N_10496,N_10192,N_10068);
or U10497 (N_10497,N_10103,N_10070);
nor U10498 (N_10498,N_10105,N_10167);
nor U10499 (N_10499,N_10117,N_10029);
nand U10500 (N_10500,N_10422,N_10331);
or U10501 (N_10501,N_10303,N_10277);
or U10502 (N_10502,N_10358,N_10292);
and U10503 (N_10503,N_10425,N_10278);
nand U10504 (N_10504,N_10411,N_10275);
xor U10505 (N_10505,N_10271,N_10360);
nor U10506 (N_10506,N_10469,N_10431);
xnor U10507 (N_10507,N_10429,N_10433);
or U10508 (N_10508,N_10324,N_10366);
or U10509 (N_10509,N_10492,N_10305);
nor U10510 (N_10510,N_10444,N_10397);
or U10511 (N_10511,N_10385,N_10461);
or U10512 (N_10512,N_10262,N_10452);
or U10513 (N_10513,N_10339,N_10463);
and U10514 (N_10514,N_10441,N_10494);
or U10515 (N_10515,N_10352,N_10491);
nand U10516 (N_10516,N_10322,N_10318);
and U10517 (N_10517,N_10270,N_10384);
nor U10518 (N_10518,N_10474,N_10319);
xnor U10519 (N_10519,N_10282,N_10398);
xor U10520 (N_10520,N_10298,N_10455);
nand U10521 (N_10521,N_10269,N_10458);
nor U10522 (N_10522,N_10481,N_10294);
nand U10523 (N_10523,N_10283,N_10403);
and U10524 (N_10524,N_10432,N_10436);
and U10525 (N_10525,N_10389,N_10295);
or U10526 (N_10526,N_10465,N_10453);
nand U10527 (N_10527,N_10310,N_10409);
nor U10528 (N_10528,N_10430,N_10258);
nand U10529 (N_10529,N_10382,N_10467);
and U10530 (N_10530,N_10479,N_10497);
or U10531 (N_10531,N_10256,N_10364);
xnor U10532 (N_10532,N_10290,N_10427);
nor U10533 (N_10533,N_10407,N_10288);
and U10534 (N_10534,N_10377,N_10372);
xnor U10535 (N_10535,N_10468,N_10350);
xnor U10536 (N_10536,N_10406,N_10442);
and U10537 (N_10537,N_10268,N_10466);
nand U10538 (N_10538,N_10284,N_10253);
or U10539 (N_10539,N_10287,N_10296);
nand U10540 (N_10540,N_10289,N_10402);
nor U10541 (N_10541,N_10304,N_10456);
and U10542 (N_10542,N_10381,N_10336);
xor U10543 (N_10543,N_10308,N_10399);
nor U10544 (N_10544,N_10485,N_10250);
nor U10545 (N_10545,N_10482,N_10415);
nand U10546 (N_10546,N_10274,N_10487);
nand U10547 (N_10547,N_10301,N_10311);
or U10548 (N_10548,N_10499,N_10363);
nor U10549 (N_10549,N_10367,N_10255);
or U10550 (N_10550,N_10328,N_10323);
nor U10551 (N_10551,N_10405,N_10483);
nand U10552 (N_10552,N_10417,N_10327);
xor U10553 (N_10553,N_10261,N_10299);
nor U10554 (N_10554,N_10267,N_10314);
and U10555 (N_10555,N_10393,N_10378);
xor U10556 (N_10556,N_10484,N_10471);
and U10557 (N_10557,N_10281,N_10330);
nand U10558 (N_10558,N_10306,N_10419);
and U10559 (N_10559,N_10280,N_10451);
and U10560 (N_10560,N_10259,N_10357);
or U10561 (N_10561,N_10450,N_10349);
or U10562 (N_10562,N_10416,N_10495);
and U10563 (N_10563,N_10401,N_10344);
xor U10564 (N_10564,N_10439,N_10476);
xnor U10565 (N_10565,N_10293,N_10437);
nor U10566 (N_10566,N_10320,N_10337);
nand U10567 (N_10567,N_10462,N_10365);
nor U10568 (N_10568,N_10457,N_10414);
nand U10569 (N_10569,N_10470,N_10346);
xor U10570 (N_10570,N_10252,N_10276);
or U10571 (N_10571,N_10359,N_10257);
and U10572 (N_10572,N_10446,N_10376);
and U10573 (N_10573,N_10345,N_10477);
or U10574 (N_10574,N_10395,N_10263);
nor U10575 (N_10575,N_10353,N_10307);
or U10576 (N_10576,N_10373,N_10408);
or U10577 (N_10577,N_10434,N_10272);
nor U10578 (N_10578,N_10354,N_10392);
xnor U10579 (N_10579,N_10266,N_10420);
and U10580 (N_10580,N_10454,N_10410);
or U10581 (N_10581,N_10371,N_10412);
or U10582 (N_10582,N_10370,N_10480);
xnor U10583 (N_10583,N_10300,N_10362);
and U10584 (N_10584,N_10369,N_10251);
nor U10585 (N_10585,N_10291,N_10348);
xnor U10586 (N_10586,N_10356,N_10326);
or U10587 (N_10587,N_10460,N_10341);
nor U10588 (N_10588,N_10343,N_10285);
nor U10589 (N_10589,N_10390,N_10347);
and U10590 (N_10590,N_10321,N_10418);
or U10591 (N_10591,N_10498,N_10489);
xor U10592 (N_10592,N_10400,N_10421);
xnor U10593 (N_10593,N_10375,N_10368);
xnor U10594 (N_10594,N_10380,N_10329);
or U10595 (N_10595,N_10279,N_10309);
nor U10596 (N_10596,N_10426,N_10254);
nor U10597 (N_10597,N_10448,N_10404);
or U10598 (N_10598,N_10312,N_10286);
or U10599 (N_10599,N_10447,N_10313);
or U10600 (N_10600,N_10334,N_10265);
or U10601 (N_10601,N_10413,N_10332);
and U10602 (N_10602,N_10342,N_10388);
and U10603 (N_10603,N_10374,N_10325);
nor U10604 (N_10604,N_10361,N_10493);
xor U10605 (N_10605,N_10440,N_10264);
and U10606 (N_10606,N_10387,N_10475);
or U10607 (N_10607,N_10317,N_10449);
nor U10608 (N_10608,N_10379,N_10355);
xor U10609 (N_10609,N_10488,N_10391);
xor U10610 (N_10610,N_10424,N_10472);
nor U10611 (N_10611,N_10435,N_10490);
and U10612 (N_10612,N_10333,N_10459);
and U10613 (N_10613,N_10496,N_10486);
nor U10614 (N_10614,N_10260,N_10315);
xor U10615 (N_10615,N_10464,N_10297);
xnor U10616 (N_10616,N_10445,N_10473);
or U10617 (N_10617,N_10338,N_10340);
nor U10618 (N_10618,N_10396,N_10351);
and U10619 (N_10619,N_10316,N_10386);
or U10620 (N_10620,N_10423,N_10443);
nor U10621 (N_10621,N_10335,N_10394);
or U10622 (N_10622,N_10438,N_10428);
and U10623 (N_10623,N_10273,N_10383);
or U10624 (N_10624,N_10478,N_10302);
nand U10625 (N_10625,N_10329,N_10368);
nand U10626 (N_10626,N_10255,N_10424);
nor U10627 (N_10627,N_10455,N_10428);
and U10628 (N_10628,N_10296,N_10453);
and U10629 (N_10629,N_10422,N_10499);
and U10630 (N_10630,N_10336,N_10499);
and U10631 (N_10631,N_10277,N_10339);
and U10632 (N_10632,N_10461,N_10474);
nand U10633 (N_10633,N_10250,N_10391);
or U10634 (N_10634,N_10258,N_10451);
or U10635 (N_10635,N_10456,N_10377);
and U10636 (N_10636,N_10256,N_10332);
xor U10637 (N_10637,N_10287,N_10282);
nand U10638 (N_10638,N_10381,N_10431);
or U10639 (N_10639,N_10351,N_10262);
or U10640 (N_10640,N_10457,N_10318);
and U10641 (N_10641,N_10436,N_10409);
nand U10642 (N_10642,N_10483,N_10289);
and U10643 (N_10643,N_10464,N_10402);
nand U10644 (N_10644,N_10358,N_10373);
or U10645 (N_10645,N_10266,N_10271);
or U10646 (N_10646,N_10457,N_10278);
nand U10647 (N_10647,N_10397,N_10395);
nand U10648 (N_10648,N_10360,N_10459);
and U10649 (N_10649,N_10256,N_10430);
nor U10650 (N_10650,N_10341,N_10494);
or U10651 (N_10651,N_10288,N_10426);
or U10652 (N_10652,N_10449,N_10338);
nor U10653 (N_10653,N_10447,N_10276);
nand U10654 (N_10654,N_10485,N_10397);
or U10655 (N_10655,N_10319,N_10350);
or U10656 (N_10656,N_10497,N_10372);
and U10657 (N_10657,N_10345,N_10380);
nand U10658 (N_10658,N_10493,N_10354);
nand U10659 (N_10659,N_10351,N_10488);
nor U10660 (N_10660,N_10264,N_10419);
or U10661 (N_10661,N_10475,N_10283);
or U10662 (N_10662,N_10464,N_10271);
xor U10663 (N_10663,N_10432,N_10380);
and U10664 (N_10664,N_10408,N_10462);
xnor U10665 (N_10665,N_10275,N_10378);
or U10666 (N_10666,N_10329,N_10280);
xnor U10667 (N_10667,N_10374,N_10429);
and U10668 (N_10668,N_10397,N_10353);
or U10669 (N_10669,N_10300,N_10449);
and U10670 (N_10670,N_10288,N_10422);
nand U10671 (N_10671,N_10313,N_10295);
nand U10672 (N_10672,N_10456,N_10347);
or U10673 (N_10673,N_10389,N_10401);
or U10674 (N_10674,N_10324,N_10314);
or U10675 (N_10675,N_10398,N_10402);
nor U10676 (N_10676,N_10257,N_10313);
or U10677 (N_10677,N_10310,N_10384);
and U10678 (N_10678,N_10359,N_10260);
xor U10679 (N_10679,N_10350,N_10388);
xor U10680 (N_10680,N_10378,N_10370);
or U10681 (N_10681,N_10400,N_10276);
and U10682 (N_10682,N_10471,N_10340);
or U10683 (N_10683,N_10387,N_10351);
or U10684 (N_10684,N_10294,N_10316);
xor U10685 (N_10685,N_10361,N_10274);
nor U10686 (N_10686,N_10357,N_10291);
and U10687 (N_10687,N_10276,N_10312);
nor U10688 (N_10688,N_10287,N_10475);
or U10689 (N_10689,N_10410,N_10419);
nand U10690 (N_10690,N_10271,N_10297);
and U10691 (N_10691,N_10259,N_10468);
nor U10692 (N_10692,N_10413,N_10365);
and U10693 (N_10693,N_10463,N_10444);
xnor U10694 (N_10694,N_10392,N_10280);
and U10695 (N_10695,N_10380,N_10438);
nor U10696 (N_10696,N_10489,N_10402);
nor U10697 (N_10697,N_10300,N_10417);
and U10698 (N_10698,N_10493,N_10369);
or U10699 (N_10699,N_10482,N_10492);
xnor U10700 (N_10700,N_10360,N_10320);
or U10701 (N_10701,N_10256,N_10354);
xnor U10702 (N_10702,N_10281,N_10473);
nand U10703 (N_10703,N_10442,N_10421);
or U10704 (N_10704,N_10430,N_10428);
nor U10705 (N_10705,N_10379,N_10490);
nor U10706 (N_10706,N_10439,N_10413);
and U10707 (N_10707,N_10341,N_10466);
nor U10708 (N_10708,N_10437,N_10374);
nor U10709 (N_10709,N_10284,N_10433);
and U10710 (N_10710,N_10255,N_10465);
and U10711 (N_10711,N_10364,N_10268);
nor U10712 (N_10712,N_10477,N_10462);
nor U10713 (N_10713,N_10391,N_10398);
and U10714 (N_10714,N_10331,N_10426);
or U10715 (N_10715,N_10488,N_10331);
nor U10716 (N_10716,N_10473,N_10477);
or U10717 (N_10717,N_10391,N_10491);
nand U10718 (N_10718,N_10387,N_10256);
and U10719 (N_10719,N_10358,N_10345);
or U10720 (N_10720,N_10485,N_10259);
or U10721 (N_10721,N_10305,N_10268);
nor U10722 (N_10722,N_10456,N_10276);
nor U10723 (N_10723,N_10424,N_10293);
and U10724 (N_10724,N_10372,N_10411);
xnor U10725 (N_10725,N_10464,N_10448);
and U10726 (N_10726,N_10413,N_10361);
nand U10727 (N_10727,N_10350,N_10324);
nor U10728 (N_10728,N_10419,N_10409);
nor U10729 (N_10729,N_10386,N_10421);
nand U10730 (N_10730,N_10263,N_10442);
and U10731 (N_10731,N_10390,N_10315);
nor U10732 (N_10732,N_10289,N_10370);
nand U10733 (N_10733,N_10458,N_10482);
nor U10734 (N_10734,N_10379,N_10328);
xnor U10735 (N_10735,N_10491,N_10301);
xnor U10736 (N_10736,N_10258,N_10305);
nor U10737 (N_10737,N_10307,N_10289);
or U10738 (N_10738,N_10254,N_10440);
nor U10739 (N_10739,N_10454,N_10381);
nand U10740 (N_10740,N_10326,N_10312);
or U10741 (N_10741,N_10261,N_10307);
and U10742 (N_10742,N_10385,N_10375);
and U10743 (N_10743,N_10476,N_10261);
nand U10744 (N_10744,N_10446,N_10437);
nor U10745 (N_10745,N_10479,N_10319);
xor U10746 (N_10746,N_10308,N_10434);
nor U10747 (N_10747,N_10273,N_10495);
nand U10748 (N_10748,N_10471,N_10433);
nand U10749 (N_10749,N_10285,N_10383);
and U10750 (N_10750,N_10506,N_10605);
or U10751 (N_10751,N_10632,N_10732);
and U10752 (N_10752,N_10642,N_10600);
nand U10753 (N_10753,N_10628,N_10552);
nand U10754 (N_10754,N_10741,N_10652);
xnor U10755 (N_10755,N_10687,N_10596);
nor U10756 (N_10756,N_10518,N_10546);
nor U10757 (N_10757,N_10705,N_10556);
nand U10758 (N_10758,N_10611,N_10661);
xor U10759 (N_10759,N_10582,N_10640);
or U10760 (N_10760,N_10578,N_10604);
nand U10761 (N_10761,N_10625,N_10509);
xor U10762 (N_10762,N_10638,N_10601);
nand U10763 (N_10763,N_10514,N_10505);
nor U10764 (N_10764,N_10579,N_10629);
nor U10765 (N_10765,N_10694,N_10635);
xnor U10766 (N_10766,N_10621,N_10570);
nand U10767 (N_10767,N_10550,N_10738);
or U10768 (N_10768,N_10670,N_10520);
nand U10769 (N_10769,N_10606,N_10698);
or U10770 (N_10770,N_10585,N_10569);
nand U10771 (N_10771,N_10526,N_10697);
xnor U10772 (N_10772,N_10691,N_10744);
nor U10773 (N_10773,N_10549,N_10648);
xor U10774 (N_10774,N_10508,N_10676);
and U10775 (N_10775,N_10567,N_10589);
nor U10776 (N_10776,N_10731,N_10673);
nand U10777 (N_10777,N_10564,N_10710);
and U10778 (N_10778,N_10669,N_10735);
nor U10779 (N_10779,N_10725,N_10533);
nand U10780 (N_10780,N_10630,N_10713);
nor U10781 (N_10781,N_10516,N_10610);
xnor U10782 (N_10782,N_10507,N_10523);
nand U10783 (N_10783,N_10666,N_10541);
nor U10784 (N_10784,N_10667,N_10620);
or U10785 (N_10785,N_10672,N_10534);
nand U10786 (N_10786,N_10524,N_10536);
nor U10787 (N_10787,N_10597,N_10679);
or U10788 (N_10788,N_10531,N_10709);
and U10789 (N_10789,N_10733,N_10558);
nand U10790 (N_10790,N_10522,N_10609);
nor U10791 (N_10791,N_10535,N_10528);
nand U10792 (N_10792,N_10702,N_10581);
or U10793 (N_10793,N_10723,N_10721);
and U10794 (N_10794,N_10665,N_10686);
xor U10795 (N_10795,N_10651,N_10706);
nor U10796 (N_10796,N_10746,N_10650);
xor U10797 (N_10797,N_10500,N_10511);
nand U10798 (N_10798,N_10704,N_10748);
and U10799 (N_10799,N_10594,N_10515);
and U10800 (N_10800,N_10747,N_10510);
and U10801 (N_10801,N_10561,N_10649);
nand U10802 (N_10802,N_10657,N_10599);
xnor U10803 (N_10803,N_10583,N_10623);
and U10804 (N_10804,N_10565,N_10719);
nor U10805 (N_10805,N_10654,N_10695);
nand U10806 (N_10806,N_10587,N_10519);
nand U10807 (N_10807,N_10591,N_10512);
or U10808 (N_10808,N_10634,N_10503);
nand U10809 (N_10809,N_10707,N_10544);
nand U10810 (N_10810,N_10712,N_10745);
nor U10811 (N_10811,N_10660,N_10580);
nor U10812 (N_10812,N_10714,N_10532);
xnor U10813 (N_10813,N_10685,N_10645);
and U10814 (N_10814,N_10680,N_10668);
xor U10815 (N_10815,N_10681,N_10644);
xnor U10816 (N_10816,N_10543,N_10734);
xnor U10817 (N_10817,N_10622,N_10577);
or U10818 (N_10818,N_10529,N_10548);
xor U10819 (N_10819,N_10737,N_10742);
xor U10820 (N_10820,N_10607,N_10688);
and U10821 (N_10821,N_10658,N_10643);
nor U10822 (N_10822,N_10545,N_10720);
or U10823 (N_10823,N_10722,N_10554);
nand U10824 (N_10824,N_10568,N_10527);
xnor U10825 (N_10825,N_10726,N_10525);
or U10826 (N_10826,N_10690,N_10730);
nor U10827 (N_10827,N_10663,N_10555);
or U10828 (N_10828,N_10617,N_10728);
nand U10829 (N_10829,N_10736,N_10504);
or U10830 (N_10830,N_10674,N_10675);
nor U10831 (N_10831,N_10696,N_10739);
xnor U10832 (N_10832,N_10647,N_10557);
xor U10833 (N_10833,N_10530,N_10573);
xor U10834 (N_10834,N_10717,N_10624);
xor U10835 (N_10835,N_10590,N_10566);
or U10836 (N_10836,N_10592,N_10718);
nand U10837 (N_10837,N_10615,N_10641);
xor U10838 (N_10838,N_10683,N_10614);
and U10839 (N_10839,N_10700,N_10693);
nand U10840 (N_10840,N_10659,N_10631);
nand U10841 (N_10841,N_10501,N_10633);
and U10842 (N_10842,N_10560,N_10586);
or U10843 (N_10843,N_10551,N_10646);
nand U10844 (N_10844,N_10729,N_10538);
nor U10845 (N_10845,N_10584,N_10572);
nor U10846 (N_10846,N_10656,N_10689);
or U10847 (N_10847,N_10616,N_10517);
and U10848 (N_10848,N_10711,N_10575);
or U10849 (N_10849,N_10636,N_10684);
xnor U10850 (N_10850,N_10671,N_10574);
nor U10851 (N_10851,N_10540,N_10602);
nor U10852 (N_10852,N_10655,N_10502);
nand U10853 (N_10853,N_10724,N_10598);
nand U10854 (N_10854,N_10562,N_10639);
or U10855 (N_10855,N_10715,N_10576);
nand U10856 (N_10856,N_10703,N_10618);
nand U10857 (N_10857,N_10627,N_10662);
or U10858 (N_10858,N_10603,N_10595);
nand U10859 (N_10859,N_10613,N_10699);
nand U10860 (N_10860,N_10677,N_10521);
nor U10861 (N_10861,N_10542,N_10537);
xor U10862 (N_10862,N_10619,N_10664);
or U10863 (N_10863,N_10553,N_10727);
or U10864 (N_10864,N_10692,N_10637);
and U10865 (N_10865,N_10716,N_10563);
and U10866 (N_10866,N_10653,N_10708);
nor U10867 (N_10867,N_10593,N_10539);
and U10868 (N_10868,N_10608,N_10626);
xnor U10869 (N_10869,N_10588,N_10559);
or U10870 (N_10870,N_10701,N_10749);
or U10871 (N_10871,N_10740,N_10612);
xor U10872 (N_10872,N_10743,N_10513);
and U10873 (N_10873,N_10571,N_10547);
or U10874 (N_10874,N_10682,N_10678);
xnor U10875 (N_10875,N_10655,N_10690);
xor U10876 (N_10876,N_10615,N_10733);
nor U10877 (N_10877,N_10587,N_10723);
nor U10878 (N_10878,N_10695,N_10679);
and U10879 (N_10879,N_10633,N_10644);
or U10880 (N_10880,N_10535,N_10641);
or U10881 (N_10881,N_10515,N_10589);
and U10882 (N_10882,N_10668,N_10682);
and U10883 (N_10883,N_10512,N_10635);
nor U10884 (N_10884,N_10692,N_10595);
nand U10885 (N_10885,N_10510,N_10556);
nor U10886 (N_10886,N_10580,N_10625);
and U10887 (N_10887,N_10537,N_10651);
nor U10888 (N_10888,N_10603,N_10511);
nor U10889 (N_10889,N_10522,N_10532);
or U10890 (N_10890,N_10539,N_10644);
nand U10891 (N_10891,N_10656,N_10657);
and U10892 (N_10892,N_10683,N_10539);
and U10893 (N_10893,N_10610,N_10727);
or U10894 (N_10894,N_10702,N_10624);
xor U10895 (N_10895,N_10744,N_10567);
nand U10896 (N_10896,N_10623,N_10671);
nor U10897 (N_10897,N_10561,N_10667);
xnor U10898 (N_10898,N_10641,N_10589);
and U10899 (N_10899,N_10586,N_10675);
xor U10900 (N_10900,N_10704,N_10603);
and U10901 (N_10901,N_10594,N_10605);
or U10902 (N_10902,N_10698,N_10510);
and U10903 (N_10903,N_10745,N_10738);
xor U10904 (N_10904,N_10619,N_10515);
nand U10905 (N_10905,N_10728,N_10541);
nor U10906 (N_10906,N_10540,N_10715);
and U10907 (N_10907,N_10553,N_10541);
nor U10908 (N_10908,N_10661,N_10592);
xor U10909 (N_10909,N_10718,N_10584);
nor U10910 (N_10910,N_10500,N_10632);
nand U10911 (N_10911,N_10649,N_10526);
nor U10912 (N_10912,N_10516,N_10645);
or U10913 (N_10913,N_10654,N_10680);
or U10914 (N_10914,N_10700,N_10505);
nor U10915 (N_10915,N_10512,N_10648);
xor U10916 (N_10916,N_10742,N_10663);
nand U10917 (N_10917,N_10728,N_10527);
nand U10918 (N_10918,N_10613,N_10629);
nand U10919 (N_10919,N_10602,N_10680);
xnor U10920 (N_10920,N_10662,N_10532);
or U10921 (N_10921,N_10512,N_10531);
or U10922 (N_10922,N_10542,N_10635);
nand U10923 (N_10923,N_10565,N_10652);
nor U10924 (N_10924,N_10547,N_10544);
and U10925 (N_10925,N_10604,N_10694);
xnor U10926 (N_10926,N_10549,N_10525);
and U10927 (N_10927,N_10722,N_10657);
nand U10928 (N_10928,N_10723,N_10555);
and U10929 (N_10929,N_10614,N_10531);
nand U10930 (N_10930,N_10606,N_10683);
nor U10931 (N_10931,N_10711,N_10653);
nor U10932 (N_10932,N_10551,N_10579);
and U10933 (N_10933,N_10672,N_10595);
nand U10934 (N_10934,N_10727,N_10584);
or U10935 (N_10935,N_10729,N_10591);
xor U10936 (N_10936,N_10660,N_10690);
or U10937 (N_10937,N_10573,N_10512);
xor U10938 (N_10938,N_10574,N_10573);
nand U10939 (N_10939,N_10715,N_10563);
and U10940 (N_10940,N_10634,N_10554);
nand U10941 (N_10941,N_10681,N_10655);
nand U10942 (N_10942,N_10529,N_10558);
or U10943 (N_10943,N_10640,N_10721);
nor U10944 (N_10944,N_10505,N_10693);
nand U10945 (N_10945,N_10666,N_10729);
or U10946 (N_10946,N_10651,N_10608);
xor U10947 (N_10947,N_10652,N_10705);
nand U10948 (N_10948,N_10574,N_10524);
nor U10949 (N_10949,N_10747,N_10718);
or U10950 (N_10950,N_10585,N_10680);
and U10951 (N_10951,N_10500,N_10609);
xnor U10952 (N_10952,N_10523,N_10622);
nand U10953 (N_10953,N_10554,N_10713);
xnor U10954 (N_10954,N_10570,N_10568);
nand U10955 (N_10955,N_10719,N_10720);
nor U10956 (N_10956,N_10692,N_10585);
xnor U10957 (N_10957,N_10678,N_10500);
nor U10958 (N_10958,N_10603,N_10609);
nor U10959 (N_10959,N_10615,N_10734);
and U10960 (N_10960,N_10502,N_10615);
nand U10961 (N_10961,N_10721,N_10672);
and U10962 (N_10962,N_10685,N_10541);
or U10963 (N_10963,N_10714,N_10551);
nor U10964 (N_10964,N_10596,N_10645);
and U10965 (N_10965,N_10547,N_10651);
or U10966 (N_10966,N_10587,N_10505);
and U10967 (N_10967,N_10597,N_10528);
nand U10968 (N_10968,N_10581,N_10531);
nand U10969 (N_10969,N_10737,N_10556);
nand U10970 (N_10970,N_10626,N_10524);
nand U10971 (N_10971,N_10562,N_10553);
and U10972 (N_10972,N_10703,N_10711);
and U10973 (N_10973,N_10731,N_10695);
nand U10974 (N_10974,N_10540,N_10685);
or U10975 (N_10975,N_10626,N_10643);
and U10976 (N_10976,N_10726,N_10695);
or U10977 (N_10977,N_10608,N_10568);
or U10978 (N_10978,N_10720,N_10678);
nand U10979 (N_10979,N_10619,N_10656);
or U10980 (N_10980,N_10614,N_10621);
or U10981 (N_10981,N_10703,N_10715);
nand U10982 (N_10982,N_10646,N_10745);
and U10983 (N_10983,N_10689,N_10513);
nor U10984 (N_10984,N_10659,N_10620);
nor U10985 (N_10985,N_10563,N_10649);
and U10986 (N_10986,N_10676,N_10560);
nor U10987 (N_10987,N_10514,N_10650);
nand U10988 (N_10988,N_10725,N_10694);
nand U10989 (N_10989,N_10729,N_10595);
xor U10990 (N_10990,N_10549,N_10611);
nor U10991 (N_10991,N_10627,N_10529);
xor U10992 (N_10992,N_10642,N_10721);
and U10993 (N_10993,N_10716,N_10709);
and U10994 (N_10994,N_10628,N_10534);
nor U10995 (N_10995,N_10556,N_10617);
nand U10996 (N_10996,N_10563,N_10502);
nor U10997 (N_10997,N_10539,N_10731);
and U10998 (N_10998,N_10601,N_10529);
nand U10999 (N_10999,N_10573,N_10678);
nor U11000 (N_11000,N_10896,N_10809);
nand U11001 (N_11001,N_10788,N_10959);
xnor U11002 (N_11002,N_10843,N_10785);
or U11003 (N_11003,N_10957,N_10958);
nand U11004 (N_11004,N_10772,N_10903);
or U11005 (N_11005,N_10755,N_10965);
nand U11006 (N_11006,N_10986,N_10987);
nand U11007 (N_11007,N_10806,N_10997);
nand U11008 (N_11008,N_10906,N_10895);
nor U11009 (N_11009,N_10966,N_10898);
nand U11010 (N_11010,N_10830,N_10792);
and U11011 (N_11011,N_10962,N_10796);
nor U11012 (N_11012,N_10905,N_10827);
nor U11013 (N_11013,N_10841,N_10797);
and U11014 (N_11014,N_10976,N_10812);
nand U11015 (N_11015,N_10984,N_10920);
or U11016 (N_11016,N_10818,N_10932);
nor U11017 (N_11017,N_10759,N_10771);
nand U11018 (N_11018,N_10767,N_10793);
or U11019 (N_11019,N_10828,N_10996);
xnor U11020 (N_11020,N_10878,N_10963);
nor U11021 (N_11021,N_10825,N_10840);
xnor U11022 (N_11022,N_10938,N_10935);
nor U11023 (N_11023,N_10844,N_10801);
nand U11024 (N_11024,N_10946,N_10979);
and U11025 (N_11025,N_10995,N_10776);
xor U11026 (N_11026,N_10831,N_10846);
nand U11027 (N_11027,N_10972,N_10768);
and U11028 (N_11028,N_10899,N_10832);
and U11029 (N_11029,N_10873,N_10800);
xor U11030 (N_11030,N_10872,N_10975);
nand U11031 (N_11031,N_10762,N_10819);
and U11032 (N_11032,N_10813,N_10769);
nor U11033 (N_11033,N_10940,N_10973);
nand U11034 (N_11034,N_10980,N_10934);
or U11035 (N_11035,N_10784,N_10835);
and U11036 (N_11036,N_10950,N_10875);
xnor U11037 (N_11037,N_10939,N_10971);
or U11038 (N_11038,N_10910,N_10886);
nor U11039 (N_11039,N_10765,N_10829);
or U11040 (N_11040,N_10804,N_10894);
or U11041 (N_11041,N_10777,N_10968);
xor U11042 (N_11042,N_10851,N_10954);
or U11043 (N_11043,N_10833,N_10794);
nand U11044 (N_11044,N_10955,N_10807);
nand U11045 (N_11045,N_10871,N_10775);
and U11046 (N_11046,N_10856,N_10853);
xnor U11047 (N_11047,N_10754,N_10823);
xnor U11048 (N_11048,N_10960,N_10988);
and U11049 (N_11049,N_10751,N_10931);
nand U11050 (N_11050,N_10956,N_10845);
and U11051 (N_11051,N_10786,N_10921);
or U11052 (N_11052,N_10991,N_10880);
and U11053 (N_11053,N_10925,N_10834);
and U11054 (N_11054,N_10820,N_10847);
nand U11055 (N_11055,N_10757,N_10821);
nand U11056 (N_11056,N_10884,N_10752);
nor U11057 (N_11057,N_10766,N_10928);
xor U11058 (N_11058,N_10782,N_10941);
nand U11059 (N_11059,N_10808,N_10817);
xor U11060 (N_11060,N_10937,N_10814);
nand U11061 (N_11061,N_10867,N_10791);
nor U11062 (N_11062,N_10964,N_10949);
nor U11063 (N_11063,N_10866,N_10837);
and U11064 (N_11064,N_10913,N_10909);
nor U11065 (N_11065,N_10985,N_10865);
or U11066 (N_11066,N_10876,N_10907);
nand U11067 (N_11067,N_10815,N_10978);
and U11068 (N_11068,N_10904,N_10858);
or U11069 (N_11069,N_10838,N_10998);
and U11070 (N_11070,N_10773,N_10803);
nand U11071 (N_11071,N_10753,N_10936);
nor U11072 (N_11072,N_10994,N_10779);
or U11073 (N_11073,N_10961,N_10929);
and U11074 (N_11074,N_10848,N_10862);
nor U11075 (N_11075,N_10864,N_10982);
nor U11076 (N_11076,N_10914,N_10992);
nor U11077 (N_11077,N_10863,N_10850);
xnor U11078 (N_11078,N_10981,N_10882);
xor U11079 (N_11079,N_10854,N_10933);
and U11080 (N_11080,N_10842,N_10883);
nand U11081 (N_11081,N_10888,N_10974);
nor U11082 (N_11082,N_10917,N_10892);
nor U11083 (N_11083,N_10923,N_10967);
nand U11084 (N_11084,N_10802,N_10778);
nand U11085 (N_11085,N_10983,N_10868);
xnor U11086 (N_11086,N_10805,N_10897);
or U11087 (N_11087,N_10889,N_10943);
nor U11088 (N_11088,N_10893,N_10911);
or U11089 (N_11089,N_10953,N_10912);
nand U11090 (N_11090,N_10795,N_10926);
nand U11091 (N_11091,N_10874,N_10787);
nor U11092 (N_11092,N_10919,N_10774);
nand U11093 (N_11093,N_10869,N_10836);
or U11094 (N_11094,N_10790,N_10924);
xor U11095 (N_11095,N_10877,N_10902);
and U11096 (N_11096,N_10870,N_10761);
or U11097 (N_11097,N_10900,N_10879);
nand U11098 (N_11098,N_10945,N_10849);
nor U11099 (N_11099,N_10763,N_10799);
nand U11100 (N_11100,N_10780,N_10970);
or U11101 (N_11101,N_10750,N_10908);
and U11102 (N_11102,N_10891,N_10839);
xor U11103 (N_11103,N_10989,N_10859);
or U11104 (N_11104,N_10824,N_10810);
xor U11105 (N_11105,N_10764,N_10756);
nand U11106 (N_11106,N_10918,N_10999);
nand U11107 (N_11107,N_10952,N_10855);
nand U11108 (N_11108,N_10922,N_10760);
nand U11109 (N_11109,N_10885,N_10781);
or U11110 (N_11110,N_10948,N_10816);
or U11111 (N_11111,N_10890,N_10758);
xor U11112 (N_11112,N_10927,N_10783);
nor U11113 (N_11113,N_10887,N_10993);
nand U11114 (N_11114,N_10990,N_10852);
nor U11115 (N_11115,N_10969,N_10947);
nand U11116 (N_11116,N_10951,N_10977);
and U11117 (N_11117,N_10915,N_10916);
nand U11118 (N_11118,N_10930,N_10881);
nand U11119 (N_11119,N_10826,N_10944);
or U11120 (N_11120,N_10861,N_10860);
or U11121 (N_11121,N_10811,N_10798);
xnor U11122 (N_11122,N_10857,N_10942);
or U11123 (N_11123,N_10770,N_10901);
nor U11124 (N_11124,N_10822,N_10789);
or U11125 (N_11125,N_10784,N_10960);
nor U11126 (N_11126,N_10773,N_10771);
xnor U11127 (N_11127,N_10884,N_10774);
or U11128 (N_11128,N_10943,N_10888);
nor U11129 (N_11129,N_10971,N_10825);
and U11130 (N_11130,N_10906,N_10845);
xnor U11131 (N_11131,N_10821,N_10752);
nand U11132 (N_11132,N_10775,N_10854);
nor U11133 (N_11133,N_10927,N_10842);
and U11134 (N_11134,N_10752,N_10956);
or U11135 (N_11135,N_10788,N_10834);
and U11136 (N_11136,N_10869,N_10981);
and U11137 (N_11137,N_10819,N_10853);
or U11138 (N_11138,N_10941,N_10751);
xor U11139 (N_11139,N_10821,N_10996);
nor U11140 (N_11140,N_10951,N_10773);
nand U11141 (N_11141,N_10837,N_10778);
nand U11142 (N_11142,N_10823,N_10848);
nand U11143 (N_11143,N_10974,N_10851);
nor U11144 (N_11144,N_10984,N_10939);
nor U11145 (N_11145,N_10777,N_10841);
or U11146 (N_11146,N_10885,N_10970);
or U11147 (N_11147,N_10984,N_10990);
and U11148 (N_11148,N_10891,N_10755);
nand U11149 (N_11149,N_10913,N_10967);
nor U11150 (N_11150,N_10980,N_10782);
nor U11151 (N_11151,N_10981,N_10885);
or U11152 (N_11152,N_10767,N_10860);
nand U11153 (N_11153,N_10920,N_10996);
nor U11154 (N_11154,N_10846,N_10906);
nand U11155 (N_11155,N_10846,N_10886);
xnor U11156 (N_11156,N_10792,N_10775);
and U11157 (N_11157,N_10897,N_10942);
nand U11158 (N_11158,N_10834,N_10913);
xor U11159 (N_11159,N_10960,N_10821);
nand U11160 (N_11160,N_10906,N_10924);
nor U11161 (N_11161,N_10912,N_10825);
nand U11162 (N_11162,N_10768,N_10836);
nor U11163 (N_11163,N_10969,N_10941);
nor U11164 (N_11164,N_10936,N_10911);
nand U11165 (N_11165,N_10852,N_10770);
and U11166 (N_11166,N_10912,N_10918);
or U11167 (N_11167,N_10785,N_10775);
nor U11168 (N_11168,N_10857,N_10848);
nor U11169 (N_11169,N_10753,N_10779);
or U11170 (N_11170,N_10831,N_10911);
xor U11171 (N_11171,N_10961,N_10809);
xor U11172 (N_11172,N_10943,N_10752);
or U11173 (N_11173,N_10920,N_10819);
nand U11174 (N_11174,N_10826,N_10905);
nor U11175 (N_11175,N_10849,N_10786);
nand U11176 (N_11176,N_10866,N_10894);
nor U11177 (N_11177,N_10969,N_10942);
xnor U11178 (N_11178,N_10829,N_10974);
xor U11179 (N_11179,N_10923,N_10986);
xnor U11180 (N_11180,N_10881,N_10762);
nand U11181 (N_11181,N_10804,N_10783);
nor U11182 (N_11182,N_10971,N_10873);
and U11183 (N_11183,N_10772,N_10870);
or U11184 (N_11184,N_10848,N_10942);
or U11185 (N_11185,N_10812,N_10855);
or U11186 (N_11186,N_10890,N_10762);
or U11187 (N_11187,N_10796,N_10854);
or U11188 (N_11188,N_10877,N_10751);
nand U11189 (N_11189,N_10792,N_10754);
and U11190 (N_11190,N_10835,N_10966);
nand U11191 (N_11191,N_10843,N_10824);
xnor U11192 (N_11192,N_10886,N_10979);
nor U11193 (N_11193,N_10925,N_10927);
nor U11194 (N_11194,N_10942,N_10953);
and U11195 (N_11195,N_10922,N_10761);
and U11196 (N_11196,N_10873,N_10815);
nor U11197 (N_11197,N_10926,N_10904);
nand U11198 (N_11198,N_10964,N_10756);
or U11199 (N_11199,N_10904,N_10836);
nand U11200 (N_11200,N_10904,N_10865);
or U11201 (N_11201,N_10973,N_10900);
nand U11202 (N_11202,N_10856,N_10963);
or U11203 (N_11203,N_10830,N_10832);
nand U11204 (N_11204,N_10886,N_10800);
xnor U11205 (N_11205,N_10779,N_10990);
or U11206 (N_11206,N_10960,N_10762);
nor U11207 (N_11207,N_10836,N_10929);
and U11208 (N_11208,N_10985,N_10842);
nand U11209 (N_11209,N_10871,N_10955);
nand U11210 (N_11210,N_10853,N_10915);
nor U11211 (N_11211,N_10871,N_10828);
nor U11212 (N_11212,N_10923,N_10810);
nor U11213 (N_11213,N_10832,N_10934);
xor U11214 (N_11214,N_10842,N_10808);
nand U11215 (N_11215,N_10970,N_10969);
or U11216 (N_11216,N_10804,N_10983);
xnor U11217 (N_11217,N_10870,N_10900);
and U11218 (N_11218,N_10928,N_10780);
nand U11219 (N_11219,N_10927,N_10851);
and U11220 (N_11220,N_10795,N_10885);
nand U11221 (N_11221,N_10988,N_10763);
and U11222 (N_11222,N_10956,N_10959);
nand U11223 (N_11223,N_10961,N_10834);
xor U11224 (N_11224,N_10890,N_10862);
nand U11225 (N_11225,N_10893,N_10760);
and U11226 (N_11226,N_10972,N_10965);
nand U11227 (N_11227,N_10957,N_10995);
or U11228 (N_11228,N_10906,N_10884);
and U11229 (N_11229,N_10795,N_10755);
nand U11230 (N_11230,N_10960,N_10993);
nor U11231 (N_11231,N_10891,N_10781);
and U11232 (N_11232,N_10857,N_10958);
nand U11233 (N_11233,N_10822,N_10921);
nor U11234 (N_11234,N_10930,N_10914);
nand U11235 (N_11235,N_10908,N_10955);
nand U11236 (N_11236,N_10964,N_10893);
nand U11237 (N_11237,N_10868,N_10970);
or U11238 (N_11238,N_10875,N_10997);
or U11239 (N_11239,N_10909,N_10926);
or U11240 (N_11240,N_10826,N_10917);
xor U11241 (N_11241,N_10839,N_10755);
xnor U11242 (N_11242,N_10768,N_10787);
nor U11243 (N_11243,N_10935,N_10983);
xnor U11244 (N_11244,N_10789,N_10964);
nor U11245 (N_11245,N_10908,N_10895);
nor U11246 (N_11246,N_10906,N_10965);
nor U11247 (N_11247,N_10974,N_10787);
and U11248 (N_11248,N_10910,N_10836);
or U11249 (N_11249,N_10809,N_10759);
or U11250 (N_11250,N_11014,N_11139);
and U11251 (N_11251,N_11120,N_11114);
nor U11252 (N_11252,N_11186,N_11245);
nor U11253 (N_11253,N_11191,N_11220);
or U11254 (N_11254,N_11082,N_11215);
nand U11255 (N_11255,N_11075,N_11153);
nor U11256 (N_11256,N_11063,N_11171);
and U11257 (N_11257,N_11002,N_11109);
nor U11258 (N_11258,N_11174,N_11098);
nor U11259 (N_11259,N_11047,N_11104);
nand U11260 (N_11260,N_11119,N_11126);
nor U11261 (N_11261,N_11091,N_11200);
xor U11262 (N_11262,N_11168,N_11132);
nand U11263 (N_11263,N_11165,N_11240);
xor U11264 (N_11264,N_11013,N_11164);
or U11265 (N_11265,N_11198,N_11003);
xor U11266 (N_11266,N_11090,N_11100);
nand U11267 (N_11267,N_11026,N_11084);
nor U11268 (N_11268,N_11166,N_11218);
nor U11269 (N_11269,N_11085,N_11017);
nand U11270 (N_11270,N_11000,N_11124);
or U11271 (N_11271,N_11073,N_11018);
nand U11272 (N_11272,N_11185,N_11057);
or U11273 (N_11273,N_11233,N_11049);
or U11274 (N_11274,N_11123,N_11155);
and U11275 (N_11275,N_11223,N_11181);
and U11276 (N_11276,N_11176,N_11169);
nand U11277 (N_11277,N_11024,N_11077);
and U11278 (N_11278,N_11056,N_11137);
nand U11279 (N_11279,N_11053,N_11162);
nor U11280 (N_11280,N_11127,N_11228);
nor U11281 (N_11281,N_11148,N_11236);
or U11282 (N_11282,N_11193,N_11217);
xor U11283 (N_11283,N_11212,N_11242);
or U11284 (N_11284,N_11029,N_11197);
and U11285 (N_11285,N_11161,N_11052);
nand U11286 (N_11286,N_11247,N_11042);
or U11287 (N_11287,N_11081,N_11149);
nor U11288 (N_11288,N_11087,N_11136);
and U11289 (N_11289,N_11115,N_11088);
xor U11290 (N_11290,N_11234,N_11008);
or U11291 (N_11291,N_11158,N_11130);
xnor U11292 (N_11292,N_11069,N_11179);
or U11293 (N_11293,N_11203,N_11140);
nand U11294 (N_11294,N_11107,N_11142);
xnor U11295 (N_11295,N_11070,N_11235);
and U11296 (N_11296,N_11188,N_11071);
or U11297 (N_11297,N_11205,N_11011);
and U11298 (N_11298,N_11201,N_11040);
and U11299 (N_11299,N_11210,N_11116);
or U11300 (N_11300,N_11159,N_11046);
nor U11301 (N_11301,N_11020,N_11044);
nand U11302 (N_11302,N_11241,N_11065);
or U11303 (N_11303,N_11041,N_11019);
or U11304 (N_11304,N_11204,N_11054);
and U11305 (N_11305,N_11001,N_11093);
xor U11306 (N_11306,N_11134,N_11055);
nand U11307 (N_11307,N_11195,N_11227);
xnor U11308 (N_11308,N_11086,N_11199);
nand U11309 (N_11309,N_11023,N_11007);
xnor U11310 (N_11310,N_11202,N_11089);
or U11311 (N_11311,N_11170,N_11010);
xor U11312 (N_11312,N_11180,N_11105);
or U11313 (N_11313,N_11156,N_11160);
nand U11314 (N_11314,N_11244,N_11133);
xor U11315 (N_11315,N_11110,N_11005);
and U11316 (N_11316,N_11028,N_11224);
or U11317 (N_11317,N_11230,N_11232);
and U11318 (N_11318,N_11059,N_11106);
or U11319 (N_11319,N_11015,N_11045);
or U11320 (N_11320,N_11012,N_11048);
and U11321 (N_11321,N_11184,N_11113);
nor U11322 (N_11322,N_11222,N_11187);
and U11323 (N_11323,N_11214,N_11211);
nand U11324 (N_11324,N_11138,N_11035);
or U11325 (N_11325,N_11238,N_11150);
nand U11326 (N_11326,N_11226,N_11025);
or U11327 (N_11327,N_11021,N_11072);
or U11328 (N_11328,N_11190,N_11237);
xor U11329 (N_11329,N_11039,N_11213);
or U11330 (N_11330,N_11067,N_11079);
or U11331 (N_11331,N_11208,N_11248);
nor U11332 (N_11332,N_11207,N_11101);
nor U11333 (N_11333,N_11051,N_11239);
xnor U11334 (N_11334,N_11177,N_11050);
xnor U11335 (N_11335,N_11145,N_11102);
or U11336 (N_11336,N_11225,N_11016);
or U11337 (N_11337,N_11030,N_11032);
nor U11338 (N_11338,N_11246,N_11221);
nor U11339 (N_11339,N_11099,N_11129);
and U11340 (N_11340,N_11229,N_11112);
xor U11341 (N_11341,N_11022,N_11206);
or U11342 (N_11342,N_11034,N_11183);
nand U11343 (N_11343,N_11108,N_11122);
nand U11344 (N_11344,N_11173,N_11094);
xnor U11345 (N_11345,N_11058,N_11249);
nor U11346 (N_11346,N_11121,N_11095);
and U11347 (N_11347,N_11163,N_11076);
nor U11348 (N_11348,N_11189,N_11080);
nand U11349 (N_11349,N_11209,N_11178);
or U11350 (N_11350,N_11066,N_11037);
xor U11351 (N_11351,N_11143,N_11092);
nor U11352 (N_11352,N_11118,N_11146);
and U11353 (N_11353,N_11231,N_11078);
xor U11354 (N_11354,N_11167,N_11196);
or U11355 (N_11355,N_11064,N_11194);
nand U11356 (N_11356,N_11157,N_11243);
nand U11357 (N_11357,N_11111,N_11062);
nand U11358 (N_11358,N_11038,N_11036);
nor U11359 (N_11359,N_11009,N_11125);
or U11360 (N_11360,N_11043,N_11141);
nand U11361 (N_11361,N_11033,N_11097);
nand U11362 (N_11362,N_11074,N_11151);
nor U11363 (N_11363,N_11027,N_11061);
xnor U11364 (N_11364,N_11144,N_11216);
nor U11365 (N_11365,N_11096,N_11083);
and U11366 (N_11366,N_11152,N_11128);
and U11367 (N_11367,N_11192,N_11006);
nor U11368 (N_11368,N_11103,N_11031);
or U11369 (N_11369,N_11154,N_11131);
xor U11370 (N_11370,N_11117,N_11060);
and U11371 (N_11371,N_11219,N_11147);
nand U11372 (N_11372,N_11135,N_11175);
and U11373 (N_11373,N_11004,N_11068);
nor U11374 (N_11374,N_11182,N_11172);
nand U11375 (N_11375,N_11085,N_11090);
or U11376 (N_11376,N_11188,N_11042);
nand U11377 (N_11377,N_11065,N_11050);
and U11378 (N_11378,N_11190,N_11014);
xor U11379 (N_11379,N_11087,N_11173);
nand U11380 (N_11380,N_11144,N_11132);
nand U11381 (N_11381,N_11096,N_11128);
or U11382 (N_11382,N_11170,N_11014);
nor U11383 (N_11383,N_11133,N_11109);
xnor U11384 (N_11384,N_11042,N_11065);
nand U11385 (N_11385,N_11191,N_11245);
nand U11386 (N_11386,N_11203,N_11048);
xor U11387 (N_11387,N_11057,N_11157);
xnor U11388 (N_11388,N_11035,N_11129);
nand U11389 (N_11389,N_11021,N_11027);
or U11390 (N_11390,N_11170,N_11029);
nand U11391 (N_11391,N_11092,N_11222);
nand U11392 (N_11392,N_11102,N_11118);
nor U11393 (N_11393,N_11100,N_11161);
or U11394 (N_11394,N_11074,N_11144);
and U11395 (N_11395,N_11211,N_11055);
nand U11396 (N_11396,N_11186,N_11055);
nor U11397 (N_11397,N_11160,N_11180);
and U11398 (N_11398,N_11102,N_11066);
nand U11399 (N_11399,N_11036,N_11172);
xor U11400 (N_11400,N_11047,N_11203);
xor U11401 (N_11401,N_11123,N_11009);
or U11402 (N_11402,N_11185,N_11032);
nor U11403 (N_11403,N_11071,N_11069);
nor U11404 (N_11404,N_11091,N_11106);
xor U11405 (N_11405,N_11243,N_11094);
xnor U11406 (N_11406,N_11002,N_11037);
nor U11407 (N_11407,N_11218,N_11232);
and U11408 (N_11408,N_11144,N_11089);
and U11409 (N_11409,N_11235,N_11230);
nor U11410 (N_11410,N_11010,N_11054);
nor U11411 (N_11411,N_11071,N_11095);
nor U11412 (N_11412,N_11137,N_11185);
nor U11413 (N_11413,N_11047,N_11046);
and U11414 (N_11414,N_11136,N_11100);
or U11415 (N_11415,N_11249,N_11088);
nor U11416 (N_11416,N_11145,N_11014);
nor U11417 (N_11417,N_11113,N_11246);
nor U11418 (N_11418,N_11142,N_11144);
nor U11419 (N_11419,N_11092,N_11239);
or U11420 (N_11420,N_11192,N_11083);
and U11421 (N_11421,N_11054,N_11182);
nor U11422 (N_11422,N_11129,N_11222);
nand U11423 (N_11423,N_11236,N_11085);
nor U11424 (N_11424,N_11036,N_11188);
xor U11425 (N_11425,N_11163,N_11095);
or U11426 (N_11426,N_11229,N_11160);
and U11427 (N_11427,N_11117,N_11037);
and U11428 (N_11428,N_11051,N_11021);
or U11429 (N_11429,N_11110,N_11065);
or U11430 (N_11430,N_11129,N_11029);
nor U11431 (N_11431,N_11193,N_11123);
xor U11432 (N_11432,N_11159,N_11216);
nor U11433 (N_11433,N_11005,N_11167);
nand U11434 (N_11434,N_11012,N_11042);
and U11435 (N_11435,N_11230,N_11140);
nor U11436 (N_11436,N_11033,N_11026);
and U11437 (N_11437,N_11233,N_11186);
nand U11438 (N_11438,N_11144,N_11210);
xor U11439 (N_11439,N_11248,N_11242);
xor U11440 (N_11440,N_11023,N_11216);
nand U11441 (N_11441,N_11113,N_11045);
nand U11442 (N_11442,N_11188,N_11037);
and U11443 (N_11443,N_11038,N_11125);
nand U11444 (N_11444,N_11236,N_11126);
nand U11445 (N_11445,N_11133,N_11163);
or U11446 (N_11446,N_11096,N_11195);
or U11447 (N_11447,N_11189,N_11095);
nand U11448 (N_11448,N_11110,N_11248);
xnor U11449 (N_11449,N_11072,N_11004);
or U11450 (N_11450,N_11239,N_11065);
nand U11451 (N_11451,N_11138,N_11230);
and U11452 (N_11452,N_11225,N_11067);
and U11453 (N_11453,N_11195,N_11119);
xor U11454 (N_11454,N_11216,N_11219);
nand U11455 (N_11455,N_11049,N_11223);
xnor U11456 (N_11456,N_11094,N_11111);
and U11457 (N_11457,N_11116,N_11022);
nand U11458 (N_11458,N_11180,N_11239);
or U11459 (N_11459,N_11068,N_11223);
nor U11460 (N_11460,N_11008,N_11028);
nor U11461 (N_11461,N_11046,N_11144);
xnor U11462 (N_11462,N_11214,N_11037);
or U11463 (N_11463,N_11185,N_11144);
or U11464 (N_11464,N_11035,N_11201);
or U11465 (N_11465,N_11113,N_11061);
xnor U11466 (N_11466,N_11058,N_11220);
nand U11467 (N_11467,N_11223,N_11184);
or U11468 (N_11468,N_11245,N_11181);
and U11469 (N_11469,N_11123,N_11045);
or U11470 (N_11470,N_11221,N_11073);
or U11471 (N_11471,N_11019,N_11028);
and U11472 (N_11472,N_11193,N_11002);
and U11473 (N_11473,N_11222,N_11130);
xnor U11474 (N_11474,N_11224,N_11111);
xor U11475 (N_11475,N_11179,N_11209);
xnor U11476 (N_11476,N_11030,N_11141);
nor U11477 (N_11477,N_11016,N_11187);
nor U11478 (N_11478,N_11182,N_11018);
and U11479 (N_11479,N_11095,N_11103);
and U11480 (N_11480,N_11168,N_11072);
xor U11481 (N_11481,N_11162,N_11128);
nor U11482 (N_11482,N_11034,N_11057);
or U11483 (N_11483,N_11117,N_11122);
or U11484 (N_11484,N_11191,N_11057);
xnor U11485 (N_11485,N_11224,N_11193);
and U11486 (N_11486,N_11241,N_11007);
or U11487 (N_11487,N_11121,N_11177);
and U11488 (N_11488,N_11051,N_11157);
nor U11489 (N_11489,N_11193,N_11000);
and U11490 (N_11490,N_11079,N_11148);
nor U11491 (N_11491,N_11053,N_11166);
nor U11492 (N_11492,N_11153,N_11009);
xnor U11493 (N_11493,N_11246,N_11022);
nor U11494 (N_11494,N_11070,N_11162);
xor U11495 (N_11495,N_11044,N_11027);
and U11496 (N_11496,N_11073,N_11196);
nand U11497 (N_11497,N_11121,N_11126);
or U11498 (N_11498,N_11102,N_11211);
xor U11499 (N_11499,N_11220,N_11222);
and U11500 (N_11500,N_11278,N_11365);
xnor U11501 (N_11501,N_11378,N_11271);
nand U11502 (N_11502,N_11440,N_11451);
or U11503 (N_11503,N_11461,N_11374);
xnor U11504 (N_11504,N_11474,N_11464);
and U11505 (N_11505,N_11277,N_11429);
or U11506 (N_11506,N_11299,N_11309);
and U11507 (N_11507,N_11251,N_11263);
and U11508 (N_11508,N_11274,N_11485);
and U11509 (N_11509,N_11488,N_11421);
xor U11510 (N_11510,N_11487,N_11325);
xnor U11511 (N_11511,N_11326,N_11492);
nand U11512 (N_11512,N_11304,N_11286);
nor U11513 (N_11513,N_11352,N_11457);
nor U11514 (N_11514,N_11285,N_11341);
xnor U11515 (N_11515,N_11496,N_11427);
nand U11516 (N_11516,N_11256,N_11489);
nor U11517 (N_11517,N_11327,N_11302);
xor U11518 (N_11518,N_11337,N_11253);
xor U11519 (N_11519,N_11361,N_11407);
xor U11520 (N_11520,N_11476,N_11279);
or U11521 (N_11521,N_11390,N_11426);
or U11522 (N_11522,N_11284,N_11323);
nor U11523 (N_11523,N_11296,N_11291);
or U11524 (N_11524,N_11450,N_11437);
or U11525 (N_11525,N_11298,N_11436);
nand U11526 (N_11526,N_11287,N_11475);
or U11527 (N_11527,N_11481,N_11452);
nand U11528 (N_11528,N_11313,N_11369);
or U11529 (N_11529,N_11359,N_11430);
and U11530 (N_11530,N_11267,N_11435);
or U11531 (N_11531,N_11354,N_11269);
nor U11532 (N_11532,N_11310,N_11493);
xnor U11533 (N_11533,N_11389,N_11420);
or U11534 (N_11534,N_11348,N_11388);
xor U11535 (N_11535,N_11342,N_11293);
and U11536 (N_11536,N_11446,N_11273);
and U11537 (N_11537,N_11433,N_11300);
nor U11538 (N_11538,N_11467,N_11394);
and U11539 (N_11539,N_11470,N_11259);
or U11540 (N_11540,N_11473,N_11281);
or U11541 (N_11541,N_11479,N_11412);
xnor U11542 (N_11542,N_11490,N_11372);
nand U11543 (N_11543,N_11356,N_11398);
xnor U11544 (N_11544,N_11422,N_11431);
nor U11545 (N_11545,N_11424,N_11379);
or U11546 (N_11546,N_11373,N_11401);
nor U11547 (N_11547,N_11497,N_11261);
xor U11548 (N_11548,N_11494,N_11397);
or U11549 (N_11549,N_11305,N_11468);
xnor U11550 (N_11550,N_11417,N_11384);
or U11551 (N_11551,N_11297,N_11366);
nor U11552 (N_11552,N_11317,N_11283);
xor U11553 (N_11553,N_11498,N_11322);
and U11554 (N_11554,N_11402,N_11458);
nor U11555 (N_11555,N_11466,N_11355);
or U11556 (N_11556,N_11264,N_11331);
or U11557 (N_11557,N_11288,N_11295);
nand U11558 (N_11558,N_11328,N_11252);
nor U11559 (N_11559,N_11292,N_11339);
nor U11560 (N_11560,N_11371,N_11347);
nand U11561 (N_11561,N_11442,N_11350);
and U11562 (N_11562,N_11301,N_11334);
nor U11563 (N_11563,N_11255,N_11336);
and U11564 (N_11564,N_11363,N_11453);
nor U11565 (N_11565,N_11351,N_11260);
and U11566 (N_11566,N_11258,N_11425);
and U11567 (N_11567,N_11290,N_11480);
nand U11568 (N_11568,N_11439,N_11270);
or U11569 (N_11569,N_11445,N_11340);
or U11570 (N_11570,N_11266,N_11408);
nand U11571 (N_11571,N_11262,N_11399);
and U11572 (N_11572,N_11469,N_11478);
nand U11573 (N_11573,N_11448,N_11306);
nor U11574 (N_11574,N_11268,N_11393);
nor U11575 (N_11575,N_11491,N_11432);
or U11576 (N_11576,N_11319,N_11353);
or U11577 (N_11577,N_11345,N_11376);
xnor U11578 (N_11578,N_11343,N_11403);
and U11579 (N_11579,N_11472,N_11416);
xor U11580 (N_11580,N_11250,N_11276);
nand U11581 (N_11581,N_11335,N_11409);
and U11582 (N_11582,N_11438,N_11465);
and U11583 (N_11583,N_11392,N_11308);
or U11584 (N_11584,N_11303,N_11411);
and U11585 (N_11585,N_11375,N_11330);
nand U11586 (N_11586,N_11349,N_11362);
nor U11587 (N_11587,N_11484,N_11315);
xor U11588 (N_11588,N_11456,N_11368);
and U11589 (N_11589,N_11333,N_11383);
nand U11590 (N_11590,N_11385,N_11396);
xnor U11591 (N_11591,N_11294,N_11454);
xor U11592 (N_11592,N_11357,N_11386);
or U11593 (N_11593,N_11406,N_11377);
and U11594 (N_11594,N_11275,N_11367);
nor U11595 (N_11595,N_11444,N_11332);
xnor U11596 (N_11596,N_11364,N_11360);
nor U11597 (N_11597,N_11370,N_11410);
nor U11598 (N_11598,N_11471,N_11460);
xnor U11599 (N_11599,N_11346,N_11455);
xnor U11600 (N_11600,N_11344,N_11312);
xnor U11601 (N_11601,N_11314,N_11381);
or U11602 (N_11602,N_11358,N_11423);
xnor U11603 (N_11603,N_11324,N_11320);
and U11604 (N_11604,N_11414,N_11282);
nand U11605 (N_11605,N_11404,N_11318);
nor U11606 (N_11606,N_11486,N_11499);
and U11607 (N_11607,N_11495,N_11462);
and U11608 (N_11608,N_11311,N_11483);
nand U11609 (N_11609,N_11419,N_11447);
xnor U11610 (N_11610,N_11428,N_11280);
or U11611 (N_11611,N_11395,N_11272);
or U11612 (N_11612,N_11265,N_11434);
nor U11613 (N_11613,N_11380,N_11463);
nor U11614 (N_11614,N_11316,N_11257);
xnor U11615 (N_11615,N_11391,N_11387);
and U11616 (N_11616,N_11382,N_11289);
and U11617 (N_11617,N_11441,N_11415);
nand U11618 (N_11618,N_11405,N_11449);
nand U11619 (N_11619,N_11329,N_11307);
xor U11620 (N_11620,N_11482,N_11413);
or U11621 (N_11621,N_11443,N_11338);
or U11622 (N_11622,N_11418,N_11477);
xnor U11623 (N_11623,N_11321,N_11459);
xor U11624 (N_11624,N_11400,N_11254);
and U11625 (N_11625,N_11341,N_11299);
nor U11626 (N_11626,N_11310,N_11336);
nor U11627 (N_11627,N_11274,N_11452);
xor U11628 (N_11628,N_11392,N_11347);
xnor U11629 (N_11629,N_11365,N_11290);
xor U11630 (N_11630,N_11345,N_11470);
or U11631 (N_11631,N_11255,N_11411);
xnor U11632 (N_11632,N_11449,N_11311);
nor U11633 (N_11633,N_11366,N_11413);
xnor U11634 (N_11634,N_11499,N_11460);
and U11635 (N_11635,N_11442,N_11452);
nor U11636 (N_11636,N_11466,N_11490);
nand U11637 (N_11637,N_11423,N_11450);
nor U11638 (N_11638,N_11438,N_11450);
nand U11639 (N_11639,N_11414,N_11431);
nor U11640 (N_11640,N_11307,N_11374);
xor U11641 (N_11641,N_11454,N_11311);
or U11642 (N_11642,N_11327,N_11282);
nor U11643 (N_11643,N_11252,N_11382);
and U11644 (N_11644,N_11300,N_11328);
or U11645 (N_11645,N_11421,N_11487);
and U11646 (N_11646,N_11277,N_11403);
nor U11647 (N_11647,N_11261,N_11392);
and U11648 (N_11648,N_11267,N_11478);
nand U11649 (N_11649,N_11382,N_11277);
and U11650 (N_11650,N_11319,N_11378);
nor U11651 (N_11651,N_11480,N_11343);
and U11652 (N_11652,N_11326,N_11410);
nor U11653 (N_11653,N_11309,N_11313);
or U11654 (N_11654,N_11264,N_11420);
or U11655 (N_11655,N_11425,N_11335);
xnor U11656 (N_11656,N_11405,N_11365);
nand U11657 (N_11657,N_11440,N_11351);
nand U11658 (N_11658,N_11344,N_11303);
or U11659 (N_11659,N_11253,N_11367);
nand U11660 (N_11660,N_11371,N_11379);
nand U11661 (N_11661,N_11349,N_11251);
nor U11662 (N_11662,N_11350,N_11386);
or U11663 (N_11663,N_11398,N_11437);
or U11664 (N_11664,N_11250,N_11336);
nor U11665 (N_11665,N_11350,N_11347);
or U11666 (N_11666,N_11468,N_11279);
nor U11667 (N_11667,N_11468,N_11407);
xnor U11668 (N_11668,N_11298,N_11349);
xor U11669 (N_11669,N_11269,N_11465);
and U11670 (N_11670,N_11316,N_11357);
or U11671 (N_11671,N_11455,N_11347);
and U11672 (N_11672,N_11408,N_11299);
and U11673 (N_11673,N_11337,N_11498);
and U11674 (N_11674,N_11408,N_11480);
or U11675 (N_11675,N_11327,N_11445);
and U11676 (N_11676,N_11334,N_11374);
and U11677 (N_11677,N_11370,N_11459);
and U11678 (N_11678,N_11282,N_11393);
or U11679 (N_11679,N_11270,N_11430);
nand U11680 (N_11680,N_11265,N_11448);
or U11681 (N_11681,N_11474,N_11270);
xor U11682 (N_11682,N_11346,N_11410);
nand U11683 (N_11683,N_11296,N_11499);
xnor U11684 (N_11684,N_11260,N_11477);
nor U11685 (N_11685,N_11397,N_11436);
nor U11686 (N_11686,N_11280,N_11360);
xor U11687 (N_11687,N_11251,N_11393);
or U11688 (N_11688,N_11441,N_11307);
or U11689 (N_11689,N_11403,N_11485);
xnor U11690 (N_11690,N_11387,N_11397);
nor U11691 (N_11691,N_11455,N_11426);
nand U11692 (N_11692,N_11309,N_11404);
nor U11693 (N_11693,N_11457,N_11337);
nand U11694 (N_11694,N_11414,N_11310);
and U11695 (N_11695,N_11374,N_11345);
nand U11696 (N_11696,N_11361,N_11423);
xnor U11697 (N_11697,N_11411,N_11351);
nand U11698 (N_11698,N_11361,N_11278);
or U11699 (N_11699,N_11442,N_11261);
and U11700 (N_11700,N_11274,N_11310);
xnor U11701 (N_11701,N_11355,N_11359);
nor U11702 (N_11702,N_11466,N_11486);
or U11703 (N_11703,N_11317,N_11273);
nor U11704 (N_11704,N_11478,N_11361);
xor U11705 (N_11705,N_11495,N_11411);
and U11706 (N_11706,N_11498,N_11464);
xor U11707 (N_11707,N_11419,N_11312);
nand U11708 (N_11708,N_11445,N_11286);
nor U11709 (N_11709,N_11472,N_11377);
and U11710 (N_11710,N_11407,N_11388);
nand U11711 (N_11711,N_11474,N_11338);
or U11712 (N_11712,N_11410,N_11289);
xnor U11713 (N_11713,N_11268,N_11440);
xor U11714 (N_11714,N_11300,N_11410);
xor U11715 (N_11715,N_11461,N_11389);
nand U11716 (N_11716,N_11329,N_11374);
or U11717 (N_11717,N_11395,N_11399);
nor U11718 (N_11718,N_11349,N_11411);
nand U11719 (N_11719,N_11341,N_11434);
nand U11720 (N_11720,N_11432,N_11330);
and U11721 (N_11721,N_11440,N_11383);
nand U11722 (N_11722,N_11305,N_11434);
nor U11723 (N_11723,N_11274,N_11453);
or U11724 (N_11724,N_11328,N_11485);
nor U11725 (N_11725,N_11479,N_11422);
or U11726 (N_11726,N_11259,N_11285);
nor U11727 (N_11727,N_11266,N_11372);
xor U11728 (N_11728,N_11346,N_11300);
xor U11729 (N_11729,N_11383,N_11349);
and U11730 (N_11730,N_11368,N_11438);
nand U11731 (N_11731,N_11404,N_11360);
or U11732 (N_11732,N_11321,N_11277);
nor U11733 (N_11733,N_11451,N_11415);
and U11734 (N_11734,N_11328,N_11306);
or U11735 (N_11735,N_11443,N_11360);
nor U11736 (N_11736,N_11419,N_11418);
xor U11737 (N_11737,N_11423,N_11471);
nor U11738 (N_11738,N_11329,N_11335);
and U11739 (N_11739,N_11409,N_11285);
and U11740 (N_11740,N_11460,N_11347);
nor U11741 (N_11741,N_11423,N_11413);
xnor U11742 (N_11742,N_11427,N_11400);
nand U11743 (N_11743,N_11278,N_11426);
nor U11744 (N_11744,N_11297,N_11407);
and U11745 (N_11745,N_11433,N_11425);
nor U11746 (N_11746,N_11268,N_11333);
nand U11747 (N_11747,N_11411,N_11392);
nand U11748 (N_11748,N_11260,N_11290);
xnor U11749 (N_11749,N_11365,N_11323);
nor U11750 (N_11750,N_11733,N_11539);
or U11751 (N_11751,N_11723,N_11640);
and U11752 (N_11752,N_11701,N_11556);
and U11753 (N_11753,N_11529,N_11703);
and U11754 (N_11754,N_11522,N_11536);
nor U11755 (N_11755,N_11661,N_11714);
and U11756 (N_11756,N_11745,N_11528);
nand U11757 (N_11757,N_11666,N_11742);
xnor U11758 (N_11758,N_11644,N_11656);
nand U11759 (N_11759,N_11577,N_11713);
nand U11760 (N_11760,N_11515,N_11610);
and U11761 (N_11761,N_11537,N_11696);
nor U11762 (N_11762,N_11524,N_11594);
or U11763 (N_11763,N_11639,N_11500);
nand U11764 (N_11764,N_11591,N_11698);
and U11765 (N_11765,N_11635,N_11676);
nor U11766 (N_11766,N_11562,N_11715);
or U11767 (N_11767,N_11711,N_11568);
or U11768 (N_11768,N_11580,N_11626);
or U11769 (N_11769,N_11535,N_11619);
or U11770 (N_11770,N_11633,N_11622);
xor U11771 (N_11771,N_11743,N_11514);
xor U11772 (N_11772,N_11678,N_11718);
nor U11773 (N_11773,N_11726,N_11706);
xnor U11774 (N_11774,N_11675,N_11617);
nand U11775 (N_11775,N_11531,N_11663);
nand U11776 (N_11776,N_11566,N_11513);
or U11777 (N_11777,N_11729,N_11605);
nand U11778 (N_11778,N_11658,N_11637);
xnor U11779 (N_11779,N_11673,N_11560);
nor U11780 (N_11780,N_11542,N_11685);
and U11781 (N_11781,N_11692,N_11590);
nand U11782 (N_11782,N_11611,N_11749);
nor U11783 (N_11783,N_11693,N_11501);
and U11784 (N_11784,N_11550,N_11554);
xor U11785 (N_11785,N_11563,N_11732);
or U11786 (N_11786,N_11683,N_11695);
or U11787 (N_11787,N_11652,N_11547);
xnor U11788 (N_11788,N_11670,N_11662);
xnor U11789 (N_11789,N_11541,N_11603);
and U11790 (N_11790,N_11565,N_11721);
xnor U11791 (N_11791,N_11601,N_11735);
or U11792 (N_11792,N_11671,N_11588);
and U11793 (N_11793,N_11686,N_11578);
nor U11794 (N_11794,N_11651,N_11579);
nand U11795 (N_11795,N_11621,N_11697);
or U11796 (N_11796,N_11570,N_11704);
xor U11797 (N_11797,N_11629,N_11689);
and U11798 (N_11798,N_11725,N_11564);
xnor U11799 (N_11799,N_11506,N_11625);
and U11800 (N_11800,N_11600,N_11700);
nand U11801 (N_11801,N_11719,N_11624);
nand U11802 (N_11802,N_11608,N_11727);
or U11803 (N_11803,N_11618,N_11614);
or U11804 (N_11804,N_11572,N_11620);
or U11805 (N_11805,N_11731,N_11709);
and U11806 (N_11806,N_11592,N_11609);
nor U11807 (N_11807,N_11660,N_11634);
nand U11808 (N_11808,N_11687,N_11615);
nand U11809 (N_11809,N_11505,N_11523);
xnor U11810 (N_11810,N_11654,N_11544);
nor U11811 (N_11811,N_11606,N_11672);
and U11812 (N_11812,N_11641,N_11737);
xor U11813 (N_11813,N_11503,N_11589);
or U11814 (N_11814,N_11728,N_11583);
xor U11815 (N_11815,N_11741,N_11525);
or U11816 (N_11816,N_11538,N_11584);
and U11817 (N_11817,N_11680,N_11585);
nor U11818 (N_11818,N_11543,N_11534);
and U11819 (N_11819,N_11631,N_11712);
nor U11820 (N_11820,N_11736,N_11521);
xnor U11821 (N_11821,N_11630,N_11677);
and U11822 (N_11822,N_11738,N_11667);
and U11823 (N_11823,N_11645,N_11682);
or U11824 (N_11824,N_11558,N_11596);
nor U11825 (N_11825,N_11607,N_11730);
xor U11826 (N_11826,N_11613,N_11582);
xnor U11827 (N_11827,N_11679,N_11587);
nor U11828 (N_11828,N_11746,N_11520);
or U11829 (N_11829,N_11708,N_11688);
xnor U11830 (N_11830,N_11722,N_11648);
nand U11831 (N_11831,N_11517,N_11552);
nand U11832 (N_11832,N_11502,N_11616);
and U11833 (N_11833,N_11623,N_11567);
xnor U11834 (N_11834,N_11694,N_11668);
nand U11835 (N_11835,N_11657,N_11724);
and U11836 (N_11836,N_11548,N_11598);
xnor U11837 (N_11837,N_11576,N_11530);
nand U11838 (N_11838,N_11553,N_11581);
or U11839 (N_11839,N_11707,N_11551);
nor U11840 (N_11840,N_11511,N_11504);
xor U11841 (N_11841,N_11717,N_11734);
nor U11842 (N_11842,N_11740,N_11512);
nand U11843 (N_11843,N_11612,N_11699);
nor U11844 (N_11844,N_11602,N_11540);
nand U11845 (N_11845,N_11595,N_11664);
nand U11846 (N_11846,N_11569,N_11638);
nand U11847 (N_11847,N_11628,N_11518);
nor U11848 (N_11848,N_11650,N_11561);
or U11849 (N_11849,N_11527,N_11681);
nand U11850 (N_11850,N_11716,N_11636);
or U11851 (N_11851,N_11507,N_11586);
and U11852 (N_11852,N_11647,N_11649);
and U11853 (N_11853,N_11546,N_11627);
and U11854 (N_11854,N_11747,N_11557);
xor U11855 (N_11855,N_11549,N_11599);
or U11856 (N_11856,N_11559,N_11533);
nor U11857 (N_11857,N_11690,N_11720);
nand U11858 (N_11858,N_11702,N_11508);
nor U11859 (N_11859,N_11643,N_11575);
and U11860 (N_11860,N_11509,N_11574);
and U11861 (N_11861,N_11519,N_11555);
and U11862 (N_11862,N_11516,N_11545);
or U11863 (N_11863,N_11705,N_11684);
nor U11864 (N_11864,N_11710,N_11655);
or U11865 (N_11865,N_11739,N_11593);
nand U11866 (N_11866,N_11573,N_11642);
and U11867 (N_11867,N_11510,N_11646);
xor U11868 (N_11868,N_11674,N_11632);
xnor U11869 (N_11869,N_11597,N_11659);
nor U11870 (N_11870,N_11526,N_11665);
nor U11871 (N_11871,N_11532,N_11653);
xor U11872 (N_11872,N_11748,N_11571);
nor U11873 (N_11873,N_11691,N_11604);
xor U11874 (N_11874,N_11744,N_11669);
xor U11875 (N_11875,N_11719,N_11610);
nand U11876 (N_11876,N_11693,N_11527);
nand U11877 (N_11877,N_11559,N_11640);
and U11878 (N_11878,N_11599,N_11593);
nand U11879 (N_11879,N_11708,N_11675);
or U11880 (N_11880,N_11646,N_11740);
nor U11881 (N_11881,N_11585,N_11545);
or U11882 (N_11882,N_11715,N_11548);
and U11883 (N_11883,N_11714,N_11615);
and U11884 (N_11884,N_11677,N_11687);
xor U11885 (N_11885,N_11657,N_11602);
or U11886 (N_11886,N_11638,N_11530);
nor U11887 (N_11887,N_11522,N_11668);
nand U11888 (N_11888,N_11696,N_11647);
xor U11889 (N_11889,N_11529,N_11526);
xor U11890 (N_11890,N_11570,N_11697);
and U11891 (N_11891,N_11684,N_11679);
nor U11892 (N_11892,N_11606,N_11577);
nor U11893 (N_11893,N_11562,N_11675);
nand U11894 (N_11894,N_11552,N_11562);
and U11895 (N_11895,N_11651,N_11543);
or U11896 (N_11896,N_11679,N_11729);
xnor U11897 (N_11897,N_11669,N_11576);
or U11898 (N_11898,N_11506,N_11694);
nor U11899 (N_11899,N_11570,N_11718);
nand U11900 (N_11900,N_11525,N_11717);
nand U11901 (N_11901,N_11602,N_11678);
nor U11902 (N_11902,N_11526,N_11663);
xnor U11903 (N_11903,N_11662,N_11591);
and U11904 (N_11904,N_11514,N_11626);
nor U11905 (N_11905,N_11684,N_11632);
nand U11906 (N_11906,N_11540,N_11588);
and U11907 (N_11907,N_11587,N_11667);
nand U11908 (N_11908,N_11629,N_11503);
or U11909 (N_11909,N_11566,N_11643);
or U11910 (N_11910,N_11740,N_11663);
xnor U11911 (N_11911,N_11711,N_11525);
nand U11912 (N_11912,N_11639,N_11654);
or U11913 (N_11913,N_11583,N_11698);
nand U11914 (N_11914,N_11544,N_11640);
nor U11915 (N_11915,N_11511,N_11623);
or U11916 (N_11916,N_11542,N_11513);
and U11917 (N_11917,N_11504,N_11660);
xor U11918 (N_11918,N_11525,N_11746);
nand U11919 (N_11919,N_11557,N_11734);
nand U11920 (N_11920,N_11668,N_11535);
xnor U11921 (N_11921,N_11524,N_11677);
xor U11922 (N_11922,N_11549,N_11626);
nor U11923 (N_11923,N_11505,N_11710);
nor U11924 (N_11924,N_11607,N_11589);
xnor U11925 (N_11925,N_11556,N_11652);
nand U11926 (N_11926,N_11653,N_11572);
nand U11927 (N_11927,N_11606,N_11584);
xnor U11928 (N_11928,N_11717,N_11588);
or U11929 (N_11929,N_11578,N_11647);
or U11930 (N_11930,N_11732,N_11608);
xnor U11931 (N_11931,N_11597,N_11714);
and U11932 (N_11932,N_11585,N_11669);
xnor U11933 (N_11933,N_11575,N_11621);
or U11934 (N_11934,N_11542,N_11586);
xnor U11935 (N_11935,N_11710,N_11672);
nor U11936 (N_11936,N_11716,N_11558);
nor U11937 (N_11937,N_11695,N_11540);
nand U11938 (N_11938,N_11616,N_11643);
and U11939 (N_11939,N_11710,N_11571);
or U11940 (N_11940,N_11509,N_11633);
or U11941 (N_11941,N_11697,N_11686);
and U11942 (N_11942,N_11713,N_11723);
and U11943 (N_11943,N_11719,N_11513);
or U11944 (N_11944,N_11739,N_11546);
nand U11945 (N_11945,N_11564,N_11601);
or U11946 (N_11946,N_11539,N_11697);
nand U11947 (N_11947,N_11612,N_11654);
and U11948 (N_11948,N_11548,N_11697);
and U11949 (N_11949,N_11665,N_11678);
or U11950 (N_11950,N_11632,N_11548);
nor U11951 (N_11951,N_11529,N_11702);
nand U11952 (N_11952,N_11563,N_11504);
or U11953 (N_11953,N_11709,N_11645);
or U11954 (N_11954,N_11593,N_11559);
nand U11955 (N_11955,N_11642,N_11594);
nand U11956 (N_11956,N_11544,N_11664);
nor U11957 (N_11957,N_11681,N_11514);
xnor U11958 (N_11958,N_11658,N_11728);
xnor U11959 (N_11959,N_11571,N_11736);
xnor U11960 (N_11960,N_11710,N_11536);
nor U11961 (N_11961,N_11718,N_11688);
xnor U11962 (N_11962,N_11608,N_11690);
xor U11963 (N_11963,N_11540,N_11542);
or U11964 (N_11964,N_11535,N_11642);
nand U11965 (N_11965,N_11577,N_11620);
or U11966 (N_11966,N_11607,N_11725);
nand U11967 (N_11967,N_11668,N_11602);
or U11968 (N_11968,N_11718,N_11691);
and U11969 (N_11969,N_11670,N_11722);
or U11970 (N_11970,N_11545,N_11608);
nor U11971 (N_11971,N_11566,N_11515);
nand U11972 (N_11972,N_11721,N_11580);
xor U11973 (N_11973,N_11637,N_11722);
nor U11974 (N_11974,N_11732,N_11513);
xnor U11975 (N_11975,N_11622,N_11728);
and U11976 (N_11976,N_11600,N_11630);
nand U11977 (N_11977,N_11668,N_11532);
xor U11978 (N_11978,N_11521,N_11748);
nand U11979 (N_11979,N_11667,N_11559);
nand U11980 (N_11980,N_11670,N_11543);
or U11981 (N_11981,N_11683,N_11613);
and U11982 (N_11982,N_11614,N_11638);
nor U11983 (N_11983,N_11697,N_11600);
xnor U11984 (N_11984,N_11743,N_11635);
xor U11985 (N_11985,N_11614,N_11641);
or U11986 (N_11986,N_11576,N_11676);
nand U11987 (N_11987,N_11555,N_11634);
or U11988 (N_11988,N_11586,N_11659);
or U11989 (N_11989,N_11619,N_11735);
nor U11990 (N_11990,N_11542,N_11729);
nand U11991 (N_11991,N_11651,N_11585);
or U11992 (N_11992,N_11651,N_11638);
nand U11993 (N_11993,N_11747,N_11578);
nor U11994 (N_11994,N_11666,N_11647);
nor U11995 (N_11995,N_11625,N_11633);
or U11996 (N_11996,N_11723,N_11627);
nand U11997 (N_11997,N_11599,N_11545);
or U11998 (N_11998,N_11500,N_11592);
nand U11999 (N_11999,N_11681,N_11512);
nor U12000 (N_12000,N_11912,N_11996);
xor U12001 (N_12001,N_11998,N_11786);
nand U12002 (N_12002,N_11922,N_11958);
and U12003 (N_12003,N_11900,N_11992);
nand U12004 (N_12004,N_11853,N_11827);
nand U12005 (N_12005,N_11888,N_11797);
or U12006 (N_12006,N_11999,N_11779);
xor U12007 (N_12007,N_11793,N_11944);
or U12008 (N_12008,N_11753,N_11765);
or U12009 (N_12009,N_11927,N_11831);
and U12010 (N_12010,N_11948,N_11868);
and U12011 (N_12011,N_11795,N_11955);
and U12012 (N_12012,N_11775,N_11890);
and U12013 (N_12013,N_11805,N_11990);
xor U12014 (N_12014,N_11938,N_11787);
and U12015 (N_12015,N_11752,N_11925);
or U12016 (N_12016,N_11909,N_11821);
or U12017 (N_12017,N_11979,N_11920);
xor U12018 (N_12018,N_11977,N_11761);
nor U12019 (N_12019,N_11806,N_11984);
nand U12020 (N_12020,N_11875,N_11928);
or U12021 (N_12021,N_11834,N_11844);
or U12022 (N_12022,N_11758,N_11874);
nor U12023 (N_12023,N_11790,N_11937);
nor U12024 (N_12024,N_11845,N_11864);
and U12025 (N_12025,N_11921,N_11974);
nand U12026 (N_12026,N_11870,N_11902);
nand U12027 (N_12027,N_11987,N_11785);
xnor U12028 (N_12028,N_11898,N_11896);
or U12029 (N_12029,N_11822,N_11768);
or U12030 (N_12030,N_11796,N_11802);
and U12031 (N_12031,N_11771,N_11947);
nor U12032 (N_12032,N_11774,N_11965);
nand U12033 (N_12033,N_11970,N_11887);
nand U12034 (N_12034,N_11762,N_11910);
nor U12035 (N_12035,N_11757,N_11832);
nor U12036 (N_12036,N_11976,N_11781);
xor U12037 (N_12037,N_11972,N_11931);
nand U12038 (N_12038,N_11830,N_11945);
nand U12039 (N_12039,N_11892,N_11897);
xnor U12040 (N_12040,N_11751,N_11985);
nor U12041 (N_12041,N_11895,N_11867);
xor U12042 (N_12042,N_11962,N_11828);
xor U12043 (N_12043,N_11759,N_11951);
and U12044 (N_12044,N_11993,N_11840);
nor U12045 (N_12045,N_11924,N_11764);
nor U12046 (N_12046,N_11926,N_11846);
and U12047 (N_12047,N_11772,N_11923);
nand U12048 (N_12048,N_11776,N_11847);
and U12049 (N_12049,N_11963,N_11769);
and U12050 (N_12050,N_11916,N_11906);
xnor U12051 (N_12051,N_11811,N_11754);
nor U12052 (N_12052,N_11756,N_11825);
nand U12053 (N_12053,N_11881,N_11879);
and U12054 (N_12054,N_11959,N_11953);
nand U12055 (N_12055,N_11939,N_11943);
xnor U12056 (N_12056,N_11843,N_11873);
or U12057 (N_12057,N_11978,N_11966);
and U12058 (N_12058,N_11901,N_11782);
or U12059 (N_12059,N_11982,N_11994);
or U12060 (N_12060,N_11824,N_11935);
nand U12061 (N_12061,N_11933,N_11871);
or U12062 (N_12062,N_11940,N_11904);
nand U12063 (N_12063,N_11755,N_11856);
and U12064 (N_12064,N_11889,N_11784);
or U12065 (N_12065,N_11988,N_11918);
nor U12066 (N_12066,N_11878,N_11778);
and U12067 (N_12067,N_11913,N_11882);
xor U12068 (N_12068,N_11810,N_11852);
nand U12069 (N_12069,N_11961,N_11934);
xor U12070 (N_12070,N_11876,N_11971);
and U12071 (N_12071,N_11919,N_11780);
nor U12072 (N_12072,N_11995,N_11957);
and U12073 (N_12073,N_11858,N_11863);
nand U12074 (N_12074,N_11880,N_11964);
nand U12075 (N_12075,N_11997,N_11777);
or U12076 (N_12076,N_11766,N_11866);
xnor U12077 (N_12077,N_11883,N_11798);
and U12078 (N_12078,N_11808,N_11989);
nor U12079 (N_12079,N_11980,N_11930);
xnor U12080 (N_12080,N_11815,N_11773);
nand U12081 (N_12081,N_11891,N_11829);
nand U12082 (N_12082,N_11855,N_11849);
nand U12083 (N_12083,N_11929,N_11817);
nand U12084 (N_12084,N_11915,N_11884);
xnor U12085 (N_12085,N_11767,N_11869);
and U12086 (N_12086,N_11789,N_11813);
and U12087 (N_12087,N_11981,N_11804);
or U12088 (N_12088,N_11986,N_11942);
nand U12089 (N_12089,N_11872,N_11914);
nand U12090 (N_12090,N_11812,N_11905);
or U12091 (N_12091,N_11837,N_11949);
xnor U12092 (N_12092,N_11911,N_11960);
and U12093 (N_12093,N_11886,N_11835);
xor U12094 (N_12094,N_11973,N_11818);
nor U12095 (N_12095,N_11791,N_11783);
xor U12096 (N_12096,N_11975,N_11952);
nand U12097 (N_12097,N_11799,N_11857);
nor U12098 (N_12098,N_11851,N_11842);
and U12099 (N_12099,N_11760,N_11809);
and U12100 (N_12100,N_11792,N_11946);
nor U12101 (N_12101,N_11859,N_11936);
or U12102 (N_12102,N_11820,N_11861);
nand U12103 (N_12103,N_11750,N_11801);
nor U12104 (N_12104,N_11763,N_11794);
nor U12105 (N_12105,N_11854,N_11803);
or U12106 (N_12106,N_11932,N_11956);
or U12107 (N_12107,N_11823,N_11899);
nand U12108 (N_12108,N_11841,N_11903);
nor U12109 (N_12109,N_11807,N_11967);
and U12110 (N_12110,N_11950,N_11848);
nor U12111 (N_12111,N_11991,N_11839);
nand U12112 (N_12112,N_11838,N_11907);
nand U12113 (N_12113,N_11814,N_11908);
nand U12114 (N_12114,N_11800,N_11862);
or U12115 (N_12115,N_11877,N_11917);
xor U12116 (N_12116,N_11833,N_11816);
or U12117 (N_12117,N_11941,N_11819);
or U12118 (N_12118,N_11770,N_11983);
and U12119 (N_12119,N_11893,N_11850);
and U12120 (N_12120,N_11894,N_11836);
xnor U12121 (N_12121,N_11865,N_11969);
and U12122 (N_12122,N_11826,N_11788);
or U12123 (N_12123,N_11954,N_11885);
and U12124 (N_12124,N_11860,N_11968);
nand U12125 (N_12125,N_11829,N_11811);
nor U12126 (N_12126,N_11934,N_11968);
or U12127 (N_12127,N_11773,N_11951);
and U12128 (N_12128,N_11817,N_11883);
and U12129 (N_12129,N_11867,N_11863);
or U12130 (N_12130,N_11846,N_11925);
nand U12131 (N_12131,N_11898,N_11928);
or U12132 (N_12132,N_11803,N_11810);
or U12133 (N_12133,N_11796,N_11887);
or U12134 (N_12134,N_11904,N_11926);
xnor U12135 (N_12135,N_11945,N_11813);
or U12136 (N_12136,N_11946,N_11862);
and U12137 (N_12137,N_11800,N_11826);
or U12138 (N_12138,N_11761,N_11959);
or U12139 (N_12139,N_11963,N_11960);
or U12140 (N_12140,N_11935,N_11855);
nand U12141 (N_12141,N_11930,N_11883);
nor U12142 (N_12142,N_11863,N_11913);
xnor U12143 (N_12143,N_11813,N_11977);
xnor U12144 (N_12144,N_11965,N_11901);
xor U12145 (N_12145,N_11912,N_11971);
nand U12146 (N_12146,N_11874,N_11994);
nand U12147 (N_12147,N_11827,N_11793);
nand U12148 (N_12148,N_11877,N_11817);
nor U12149 (N_12149,N_11776,N_11851);
xor U12150 (N_12150,N_11809,N_11785);
nand U12151 (N_12151,N_11835,N_11848);
or U12152 (N_12152,N_11771,N_11871);
nor U12153 (N_12153,N_11754,N_11994);
and U12154 (N_12154,N_11983,N_11968);
nand U12155 (N_12155,N_11968,N_11781);
or U12156 (N_12156,N_11858,N_11845);
and U12157 (N_12157,N_11797,N_11781);
nand U12158 (N_12158,N_11812,N_11847);
and U12159 (N_12159,N_11814,N_11844);
nand U12160 (N_12160,N_11965,N_11998);
or U12161 (N_12161,N_11791,N_11829);
xnor U12162 (N_12162,N_11770,N_11961);
or U12163 (N_12163,N_11952,N_11918);
xnor U12164 (N_12164,N_11761,N_11931);
or U12165 (N_12165,N_11997,N_11788);
xor U12166 (N_12166,N_11988,N_11769);
nand U12167 (N_12167,N_11926,N_11772);
nor U12168 (N_12168,N_11998,N_11906);
or U12169 (N_12169,N_11894,N_11777);
nand U12170 (N_12170,N_11867,N_11916);
xor U12171 (N_12171,N_11861,N_11765);
nand U12172 (N_12172,N_11990,N_11932);
nor U12173 (N_12173,N_11915,N_11786);
or U12174 (N_12174,N_11959,N_11937);
xnor U12175 (N_12175,N_11798,N_11996);
nand U12176 (N_12176,N_11980,N_11835);
and U12177 (N_12177,N_11935,N_11998);
nand U12178 (N_12178,N_11973,N_11849);
nand U12179 (N_12179,N_11882,N_11757);
or U12180 (N_12180,N_11958,N_11942);
nor U12181 (N_12181,N_11905,N_11864);
or U12182 (N_12182,N_11794,N_11860);
nor U12183 (N_12183,N_11807,N_11908);
or U12184 (N_12184,N_11913,N_11801);
and U12185 (N_12185,N_11753,N_11884);
xnor U12186 (N_12186,N_11796,N_11834);
nor U12187 (N_12187,N_11972,N_11819);
or U12188 (N_12188,N_11763,N_11877);
nor U12189 (N_12189,N_11867,N_11800);
or U12190 (N_12190,N_11758,N_11995);
and U12191 (N_12191,N_11841,N_11853);
nand U12192 (N_12192,N_11949,N_11805);
or U12193 (N_12193,N_11993,N_11990);
nor U12194 (N_12194,N_11852,N_11811);
nor U12195 (N_12195,N_11877,N_11822);
nor U12196 (N_12196,N_11919,N_11807);
and U12197 (N_12197,N_11944,N_11917);
or U12198 (N_12198,N_11937,N_11800);
nand U12199 (N_12199,N_11970,N_11847);
xor U12200 (N_12200,N_11812,N_11924);
and U12201 (N_12201,N_11998,N_11899);
nor U12202 (N_12202,N_11763,N_11809);
nor U12203 (N_12203,N_11930,N_11770);
or U12204 (N_12204,N_11852,N_11848);
or U12205 (N_12205,N_11869,N_11852);
nor U12206 (N_12206,N_11788,N_11862);
nand U12207 (N_12207,N_11909,N_11788);
nand U12208 (N_12208,N_11885,N_11997);
nand U12209 (N_12209,N_11874,N_11973);
nor U12210 (N_12210,N_11923,N_11751);
and U12211 (N_12211,N_11953,N_11873);
nand U12212 (N_12212,N_11807,N_11864);
nor U12213 (N_12213,N_11952,N_11900);
and U12214 (N_12214,N_11892,N_11833);
and U12215 (N_12215,N_11799,N_11755);
and U12216 (N_12216,N_11959,N_11978);
and U12217 (N_12217,N_11863,N_11902);
nand U12218 (N_12218,N_11803,N_11999);
and U12219 (N_12219,N_11817,N_11825);
or U12220 (N_12220,N_11943,N_11974);
xnor U12221 (N_12221,N_11861,N_11753);
nand U12222 (N_12222,N_11915,N_11956);
nand U12223 (N_12223,N_11927,N_11839);
xor U12224 (N_12224,N_11752,N_11899);
or U12225 (N_12225,N_11790,N_11970);
and U12226 (N_12226,N_11759,N_11791);
xnor U12227 (N_12227,N_11755,N_11823);
xnor U12228 (N_12228,N_11761,N_11784);
nor U12229 (N_12229,N_11787,N_11753);
or U12230 (N_12230,N_11873,N_11878);
and U12231 (N_12231,N_11914,N_11827);
and U12232 (N_12232,N_11921,N_11813);
nor U12233 (N_12233,N_11782,N_11828);
or U12234 (N_12234,N_11882,N_11784);
and U12235 (N_12235,N_11841,N_11805);
and U12236 (N_12236,N_11790,N_11811);
or U12237 (N_12237,N_11815,N_11843);
xor U12238 (N_12238,N_11798,N_11791);
and U12239 (N_12239,N_11959,N_11770);
or U12240 (N_12240,N_11907,N_11808);
or U12241 (N_12241,N_11787,N_11834);
xnor U12242 (N_12242,N_11925,N_11958);
xnor U12243 (N_12243,N_11812,N_11987);
nand U12244 (N_12244,N_11853,N_11938);
nand U12245 (N_12245,N_11761,N_11895);
nand U12246 (N_12246,N_11914,N_11845);
and U12247 (N_12247,N_11774,N_11932);
nand U12248 (N_12248,N_11770,N_11971);
or U12249 (N_12249,N_11798,N_11818);
nor U12250 (N_12250,N_12145,N_12138);
nor U12251 (N_12251,N_12037,N_12116);
nor U12252 (N_12252,N_12157,N_12014);
nand U12253 (N_12253,N_12063,N_12081);
nor U12254 (N_12254,N_12148,N_12082);
and U12255 (N_12255,N_12098,N_12072);
nor U12256 (N_12256,N_12057,N_12182);
nand U12257 (N_12257,N_12217,N_12067);
nand U12258 (N_12258,N_12084,N_12033);
and U12259 (N_12259,N_12097,N_12127);
nand U12260 (N_12260,N_12078,N_12123);
nand U12261 (N_12261,N_12109,N_12134);
and U12262 (N_12262,N_12003,N_12144);
xnor U12263 (N_12263,N_12112,N_12178);
or U12264 (N_12264,N_12215,N_12017);
xor U12265 (N_12265,N_12120,N_12086);
or U12266 (N_12266,N_12149,N_12042);
and U12267 (N_12267,N_12228,N_12136);
or U12268 (N_12268,N_12154,N_12010);
nand U12269 (N_12269,N_12040,N_12066);
and U12270 (N_12270,N_12119,N_12226);
nand U12271 (N_12271,N_12247,N_12176);
nand U12272 (N_12272,N_12019,N_12183);
nor U12273 (N_12273,N_12096,N_12065);
nor U12274 (N_12274,N_12049,N_12043);
nand U12275 (N_12275,N_12093,N_12091);
or U12276 (N_12276,N_12195,N_12077);
nor U12277 (N_12277,N_12175,N_12216);
xor U12278 (N_12278,N_12179,N_12237);
nor U12279 (N_12279,N_12155,N_12076);
or U12280 (N_12280,N_12204,N_12191);
nor U12281 (N_12281,N_12012,N_12186);
xor U12282 (N_12282,N_12064,N_12054);
xor U12283 (N_12283,N_12160,N_12130);
xnor U12284 (N_12284,N_12075,N_12180);
or U12285 (N_12285,N_12169,N_12047);
nand U12286 (N_12286,N_12241,N_12151);
nand U12287 (N_12287,N_12087,N_12202);
nand U12288 (N_12288,N_12126,N_12041);
xnor U12289 (N_12289,N_12245,N_12106);
nor U12290 (N_12290,N_12188,N_12122);
and U12291 (N_12291,N_12060,N_12194);
or U12292 (N_12292,N_12015,N_12227);
xnor U12293 (N_12293,N_12142,N_12146);
or U12294 (N_12294,N_12115,N_12048);
or U12295 (N_12295,N_12059,N_12213);
or U12296 (N_12296,N_12212,N_12234);
and U12297 (N_12297,N_12132,N_12099);
and U12298 (N_12298,N_12107,N_12210);
nor U12299 (N_12299,N_12231,N_12219);
nor U12300 (N_12300,N_12249,N_12208);
nor U12301 (N_12301,N_12211,N_12069);
and U12302 (N_12302,N_12030,N_12052);
and U12303 (N_12303,N_12135,N_12239);
xor U12304 (N_12304,N_12036,N_12139);
xnor U12305 (N_12305,N_12095,N_12173);
nor U12306 (N_12306,N_12187,N_12000);
nor U12307 (N_12307,N_12198,N_12094);
or U12308 (N_12308,N_12235,N_12008);
xor U12309 (N_12309,N_12232,N_12053);
xnor U12310 (N_12310,N_12248,N_12080);
nor U12311 (N_12311,N_12246,N_12058);
nand U12312 (N_12312,N_12102,N_12056);
nor U12313 (N_12313,N_12035,N_12137);
nand U12314 (N_12314,N_12150,N_12143);
nand U12315 (N_12315,N_12090,N_12029);
or U12316 (N_12316,N_12197,N_12177);
xor U12317 (N_12317,N_12161,N_12006);
and U12318 (N_12318,N_12238,N_12214);
nor U12319 (N_12319,N_12171,N_12181);
or U12320 (N_12320,N_12156,N_12224);
nand U12321 (N_12321,N_12159,N_12152);
and U12322 (N_12322,N_12113,N_12070);
nand U12323 (N_12323,N_12103,N_12189);
or U12324 (N_12324,N_12051,N_12021);
xnor U12325 (N_12325,N_12168,N_12147);
nor U12326 (N_12326,N_12218,N_12034);
nor U12327 (N_12327,N_12024,N_12193);
or U12328 (N_12328,N_12223,N_12167);
or U12329 (N_12329,N_12092,N_12174);
and U12330 (N_12330,N_12044,N_12050);
nand U12331 (N_12331,N_12089,N_12068);
nand U12332 (N_12332,N_12240,N_12242);
or U12333 (N_12333,N_12170,N_12158);
nor U12334 (N_12334,N_12205,N_12125);
and U12335 (N_12335,N_12011,N_12206);
xor U12336 (N_12336,N_12140,N_12018);
xor U12337 (N_12337,N_12105,N_12083);
nand U12338 (N_12338,N_12166,N_12209);
or U12339 (N_12339,N_12162,N_12163);
nor U12340 (N_12340,N_12071,N_12200);
and U12341 (N_12341,N_12009,N_12185);
and U12342 (N_12342,N_12124,N_12201);
nand U12343 (N_12343,N_12062,N_12244);
nand U12344 (N_12344,N_12016,N_12079);
or U12345 (N_12345,N_12153,N_12131);
nand U12346 (N_12346,N_12165,N_12046);
and U12347 (N_12347,N_12172,N_12028);
and U12348 (N_12348,N_12164,N_12236);
nor U12349 (N_12349,N_12243,N_12111);
xor U12350 (N_12350,N_12196,N_12184);
nor U12351 (N_12351,N_12027,N_12007);
nor U12352 (N_12352,N_12203,N_12207);
nor U12353 (N_12353,N_12073,N_12026);
nor U12354 (N_12354,N_12141,N_12117);
nor U12355 (N_12355,N_12133,N_12230);
xor U12356 (N_12356,N_12055,N_12101);
nand U12357 (N_12357,N_12104,N_12199);
and U12358 (N_12358,N_12225,N_12061);
nand U12359 (N_12359,N_12025,N_12233);
xor U12360 (N_12360,N_12129,N_12100);
or U12361 (N_12361,N_12128,N_12013);
xor U12362 (N_12362,N_12121,N_12004);
and U12363 (N_12363,N_12001,N_12045);
xor U12364 (N_12364,N_12039,N_12114);
and U12365 (N_12365,N_12220,N_12222);
xnor U12366 (N_12366,N_12085,N_12031);
xnor U12367 (N_12367,N_12108,N_12088);
xor U12368 (N_12368,N_12038,N_12118);
and U12369 (N_12369,N_12005,N_12023);
and U12370 (N_12370,N_12020,N_12002);
nand U12371 (N_12371,N_12022,N_12074);
nand U12372 (N_12372,N_12190,N_12032);
and U12373 (N_12373,N_12110,N_12192);
xnor U12374 (N_12374,N_12221,N_12229);
nor U12375 (N_12375,N_12202,N_12105);
nor U12376 (N_12376,N_12039,N_12246);
and U12377 (N_12377,N_12186,N_12171);
or U12378 (N_12378,N_12041,N_12047);
and U12379 (N_12379,N_12030,N_12039);
and U12380 (N_12380,N_12129,N_12103);
or U12381 (N_12381,N_12004,N_12212);
nor U12382 (N_12382,N_12207,N_12212);
xor U12383 (N_12383,N_12052,N_12004);
nand U12384 (N_12384,N_12171,N_12094);
nand U12385 (N_12385,N_12159,N_12087);
nor U12386 (N_12386,N_12112,N_12218);
xor U12387 (N_12387,N_12064,N_12012);
nor U12388 (N_12388,N_12153,N_12217);
and U12389 (N_12389,N_12175,N_12172);
nor U12390 (N_12390,N_12069,N_12056);
or U12391 (N_12391,N_12218,N_12053);
nand U12392 (N_12392,N_12136,N_12014);
nor U12393 (N_12393,N_12183,N_12078);
nand U12394 (N_12394,N_12164,N_12245);
nor U12395 (N_12395,N_12006,N_12188);
nand U12396 (N_12396,N_12043,N_12192);
or U12397 (N_12397,N_12040,N_12111);
xor U12398 (N_12398,N_12000,N_12114);
nor U12399 (N_12399,N_12041,N_12028);
nor U12400 (N_12400,N_12227,N_12105);
and U12401 (N_12401,N_12017,N_12003);
nor U12402 (N_12402,N_12103,N_12019);
nand U12403 (N_12403,N_12224,N_12139);
and U12404 (N_12404,N_12039,N_12043);
or U12405 (N_12405,N_12124,N_12100);
xnor U12406 (N_12406,N_12205,N_12028);
xor U12407 (N_12407,N_12097,N_12139);
and U12408 (N_12408,N_12126,N_12238);
or U12409 (N_12409,N_12168,N_12127);
or U12410 (N_12410,N_12162,N_12175);
or U12411 (N_12411,N_12077,N_12166);
nor U12412 (N_12412,N_12035,N_12232);
nand U12413 (N_12413,N_12209,N_12033);
nand U12414 (N_12414,N_12173,N_12003);
and U12415 (N_12415,N_12057,N_12179);
xor U12416 (N_12416,N_12099,N_12013);
nand U12417 (N_12417,N_12027,N_12054);
xor U12418 (N_12418,N_12159,N_12070);
or U12419 (N_12419,N_12177,N_12077);
nor U12420 (N_12420,N_12108,N_12134);
xnor U12421 (N_12421,N_12143,N_12154);
and U12422 (N_12422,N_12245,N_12219);
nor U12423 (N_12423,N_12037,N_12023);
or U12424 (N_12424,N_12087,N_12018);
xor U12425 (N_12425,N_12171,N_12041);
nor U12426 (N_12426,N_12197,N_12207);
xnor U12427 (N_12427,N_12181,N_12175);
xnor U12428 (N_12428,N_12177,N_12081);
nor U12429 (N_12429,N_12029,N_12008);
xnor U12430 (N_12430,N_12055,N_12176);
and U12431 (N_12431,N_12029,N_12139);
and U12432 (N_12432,N_12234,N_12060);
nand U12433 (N_12433,N_12229,N_12246);
nand U12434 (N_12434,N_12137,N_12015);
and U12435 (N_12435,N_12003,N_12134);
nand U12436 (N_12436,N_12153,N_12006);
and U12437 (N_12437,N_12229,N_12213);
nor U12438 (N_12438,N_12095,N_12207);
or U12439 (N_12439,N_12063,N_12031);
nor U12440 (N_12440,N_12052,N_12186);
nand U12441 (N_12441,N_12140,N_12153);
and U12442 (N_12442,N_12180,N_12097);
and U12443 (N_12443,N_12048,N_12104);
nor U12444 (N_12444,N_12108,N_12017);
and U12445 (N_12445,N_12248,N_12059);
nand U12446 (N_12446,N_12166,N_12126);
nand U12447 (N_12447,N_12235,N_12139);
nand U12448 (N_12448,N_12192,N_12199);
xor U12449 (N_12449,N_12122,N_12003);
and U12450 (N_12450,N_12179,N_12130);
and U12451 (N_12451,N_12160,N_12079);
nand U12452 (N_12452,N_12217,N_12117);
or U12453 (N_12453,N_12159,N_12104);
xnor U12454 (N_12454,N_12083,N_12122);
nor U12455 (N_12455,N_12019,N_12241);
or U12456 (N_12456,N_12001,N_12069);
and U12457 (N_12457,N_12240,N_12038);
xor U12458 (N_12458,N_12092,N_12068);
and U12459 (N_12459,N_12025,N_12032);
and U12460 (N_12460,N_12097,N_12151);
nor U12461 (N_12461,N_12017,N_12076);
xor U12462 (N_12462,N_12144,N_12020);
xor U12463 (N_12463,N_12138,N_12202);
nor U12464 (N_12464,N_12047,N_12029);
xor U12465 (N_12465,N_12002,N_12081);
nand U12466 (N_12466,N_12116,N_12215);
and U12467 (N_12467,N_12145,N_12142);
and U12468 (N_12468,N_12122,N_12017);
or U12469 (N_12469,N_12085,N_12194);
or U12470 (N_12470,N_12224,N_12061);
and U12471 (N_12471,N_12248,N_12206);
or U12472 (N_12472,N_12054,N_12047);
nor U12473 (N_12473,N_12225,N_12083);
or U12474 (N_12474,N_12061,N_12116);
or U12475 (N_12475,N_12130,N_12076);
xnor U12476 (N_12476,N_12101,N_12119);
nand U12477 (N_12477,N_12221,N_12076);
nand U12478 (N_12478,N_12139,N_12108);
and U12479 (N_12479,N_12043,N_12102);
xnor U12480 (N_12480,N_12234,N_12030);
and U12481 (N_12481,N_12090,N_12031);
nor U12482 (N_12482,N_12024,N_12079);
xor U12483 (N_12483,N_12052,N_12120);
and U12484 (N_12484,N_12074,N_12092);
nand U12485 (N_12485,N_12123,N_12164);
and U12486 (N_12486,N_12071,N_12057);
xnor U12487 (N_12487,N_12019,N_12021);
nand U12488 (N_12488,N_12216,N_12034);
xor U12489 (N_12489,N_12199,N_12066);
nand U12490 (N_12490,N_12067,N_12009);
and U12491 (N_12491,N_12059,N_12086);
and U12492 (N_12492,N_12217,N_12114);
nand U12493 (N_12493,N_12110,N_12060);
or U12494 (N_12494,N_12048,N_12200);
xor U12495 (N_12495,N_12173,N_12140);
or U12496 (N_12496,N_12155,N_12082);
nand U12497 (N_12497,N_12060,N_12103);
or U12498 (N_12498,N_12213,N_12045);
xnor U12499 (N_12499,N_12229,N_12222);
or U12500 (N_12500,N_12360,N_12326);
nor U12501 (N_12501,N_12310,N_12458);
nor U12502 (N_12502,N_12298,N_12390);
nand U12503 (N_12503,N_12357,N_12328);
xor U12504 (N_12504,N_12494,N_12422);
xnor U12505 (N_12505,N_12352,N_12374);
xor U12506 (N_12506,N_12448,N_12256);
nor U12507 (N_12507,N_12491,N_12294);
nand U12508 (N_12508,N_12366,N_12351);
and U12509 (N_12509,N_12464,N_12460);
or U12510 (N_12510,N_12307,N_12492);
xor U12511 (N_12511,N_12417,N_12465);
nor U12512 (N_12512,N_12312,N_12274);
and U12513 (N_12513,N_12336,N_12385);
or U12514 (N_12514,N_12322,N_12441);
nor U12515 (N_12515,N_12395,N_12305);
xor U12516 (N_12516,N_12479,N_12313);
nor U12517 (N_12517,N_12444,N_12271);
and U12518 (N_12518,N_12462,N_12414);
or U12519 (N_12519,N_12445,N_12497);
nor U12520 (N_12520,N_12436,N_12283);
xnor U12521 (N_12521,N_12498,N_12412);
xnor U12522 (N_12522,N_12253,N_12499);
nand U12523 (N_12523,N_12365,N_12387);
or U12524 (N_12524,N_12413,N_12478);
and U12525 (N_12525,N_12306,N_12471);
nor U12526 (N_12526,N_12435,N_12375);
xnor U12527 (N_12527,N_12254,N_12321);
nor U12528 (N_12528,N_12451,N_12275);
or U12529 (N_12529,N_12350,N_12411);
and U12530 (N_12530,N_12324,N_12457);
or U12531 (N_12531,N_12403,N_12373);
nand U12532 (N_12532,N_12269,N_12439);
xor U12533 (N_12533,N_12370,N_12355);
nor U12534 (N_12534,N_12386,N_12371);
nand U12535 (N_12535,N_12258,N_12361);
or U12536 (N_12536,N_12347,N_12308);
nand U12537 (N_12537,N_12282,N_12391);
and U12538 (N_12538,N_12354,N_12250);
xor U12539 (N_12539,N_12482,N_12261);
nand U12540 (N_12540,N_12267,N_12300);
nand U12541 (N_12541,N_12486,N_12472);
nor U12542 (N_12542,N_12466,N_12331);
nor U12543 (N_12543,N_12348,N_12335);
xnor U12544 (N_12544,N_12393,N_12264);
xor U12545 (N_12545,N_12311,N_12286);
and U12546 (N_12546,N_12406,N_12323);
nand U12547 (N_12547,N_12430,N_12255);
xnor U12548 (N_12548,N_12447,N_12424);
xor U12549 (N_12549,N_12303,N_12293);
nor U12550 (N_12550,N_12442,N_12450);
and U12551 (N_12551,N_12349,N_12296);
or U12552 (N_12552,N_12470,N_12426);
and U12553 (N_12553,N_12287,N_12405);
nor U12554 (N_12554,N_12290,N_12474);
or U12555 (N_12555,N_12333,N_12408);
xor U12556 (N_12556,N_12358,N_12364);
xor U12557 (N_12557,N_12420,N_12493);
xnor U12558 (N_12558,N_12401,N_12456);
nand U12559 (N_12559,N_12398,N_12276);
or U12560 (N_12560,N_12257,N_12388);
nand U12561 (N_12561,N_12315,N_12475);
nand U12562 (N_12562,N_12377,N_12483);
nor U12563 (N_12563,N_12265,N_12372);
and U12564 (N_12564,N_12489,N_12297);
and U12565 (N_12565,N_12278,N_12356);
nand U12566 (N_12566,N_12400,N_12433);
and U12567 (N_12567,N_12416,N_12337);
and U12568 (N_12568,N_12484,N_12363);
nand U12569 (N_12569,N_12446,N_12485);
xnor U12570 (N_12570,N_12302,N_12318);
or U12571 (N_12571,N_12284,N_12251);
nand U12572 (N_12572,N_12359,N_12459);
and U12573 (N_12573,N_12266,N_12380);
and U12574 (N_12574,N_12353,N_12378);
or U12575 (N_12575,N_12299,N_12453);
xnor U12576 (N_12576,N_12394,N_12399);
and U12577 (N_12577,N_12367,N_12467);
nand U12578 (N_12578,N_12440,N_12423);
or U12579 (N_12579,N_12427,N_12341);
nor U12580 (N_12580,N_12437,N_12443);
xnor U12581 (N_12581,N_12309,N_12425);
and U12582 (N_12582,N_12454,N_12468);
nor U12583 (N_12583,N_12476,N_12382);
xnor U12584 (N_12584,N_12273,N_12396);
xnor U12585 (N_12585,N_12407,N_12272);
nor U12586 (N_12586,N_12327,N_12340);
and U12587 (N_12587,N_12379,N_12344);
xor U12588 (N_12588,N_12421,N_12432);
nand U12589 (N_12589,N_12330,N_12263);
and U12590 (N_12590,N_12376,N_12292);
xnor U12591 (N_12591,N_12496,N_12277);
nand U12592 (N_12592,N_12281,N_12259);
or U12593 (N_12593,N_12304,N_12270);
or U12594 (N_12594,N_12301,N_12342);
or U12595 (N_12595,N_12452,N_12383);
or U12596 (N_12596,N_12487,N_12316);
or U12597 (N_12597,N_12280,N_12488);
nor U12598 (N_12598,N_12345,N_12317);
or U12599 (N_12599,N_12314,N_12339);
or U12600 (N_12600,N_12402,N_12455);
or U12601 (N_12601,N_12419,N_12279);
xnor U12602 (N_12602,N_12343,N_12404);
nand U12603 (N_12603,N_12288,N_12295);
nand U12604 (N_12604,N_12481,N_12428);
or U12605 (N_12605,N_12415,N_12431);
nor U12606 (N_12606,N_12260,N_12473);
and U12607 (N_12607,N_12495,N_12434);
xnor U12608 (N_12608,N_12469,N_12477);
xor U12609 (N_12609,N_12397,N_12320);
nand U12610 (N_12610,N_12252,N_12429);
nor U12611 (N_12611,N_12490,N_12389);
or U12612 (N_12612,N_12480,N_12289);
and U12613 (N_12613,N_12461,N_12369);
and U12614 (N_12614,N_12463,N_12392);
or U12615 (N_12615,N_12325,N_12334);
and U12616 (N_12616,N_12291,N_12285);
and U12617 (N_12617,N_12418,N_12346);
nand U12618 (N_12618,N_12319,N_12332);
or U12619 (N_12619,N_12410,N_12409);
nand U12620 (N_12620,N_12384,N_12329);
nor U12621 (N_12621,N_12438,N_12268);
xor U12622 (N_12622,N_12368,N_12362);
and U12623 (N_12623,N_12338,N_12381);
nor U12624 (N_12624,N_12262,N_12449);
xnor U12625 (N_12625,N_12259,N_12264);
nand U12626 (N_12626,N_12269,N_12442);
nand U12627 (N_12627,N_12426,N_12471);
nor U12628 (N_12628,N_12284,N_12420);
nand U12629 (N_12629,N_12433,N_12414);
or U12630 (N_12630,N_12288,N_12270);
nand U12631 (N_12631,N_12433,N_12370);
and U12632 (N_12632,N_12435,N_12453);
or U12633 (N_12633,N_12254,N_12450);
and U12634 (N_12634,N_12470,N_12284);
nor U12635 (N_12635,N_12399,N_12423);
or U12636 (N_12636,N_12293,N_12451);
nor U12637 (N_12637,N_12351,N_12288);
or U12638 (N_12638,N_12453,N_12305);
nor U12639 (N_12639,N_12385,N_12270);
or U12640 (N_12640,N_12401,N_12452);
nor U12641 (N_12641,N_12499,N_12378);
xor U12642 (N_12642,N_12390,N_12352);
and U12643 (N_12643,N_12312,N_12262);
and U12644 (N_12644,N_12315,N_12478);
nand U12645 (N_12645,N_12491,N_12378);
nand U12646 (N_12646,N_12254,N_12462);
or U12647 (N_12647,N_12313,N_12263);
nor U12648 (N_12648,N_12374,N_12365);
or U12649 (N_12649,N_12488,N_12414);
and U12650 (N_12650,N_12431,N_12492);
xnor U12651 (N_12651,N_12325,N_12464);
xor U12652 (N_12652,N_12304,N_12280);
or U12653 (N_12653,N_12269,N_12410);
nand U12654 (N_12654,N_12388,N_12392);
nand U12655 (N_12655,N_12418,N_12445);
xnor U12656 (N_12656,N_12374,N_12495);
and U12657 (N_12657,N_12413,N_12387);
nand U12658 (N_12658,N_12356,N_12307);
nand U12659 (N_12659,N_12476,N_12456);
nand U12660 (N_12660,N_12287,N_12416);
nor U12661 (N_12661,N_12270,N_12425);
xnor U12662 (N_12662,N_12437,N_12322);
nand U12663 (N_12663,N_12465,N_12412);
and U12664 (N_12664,N_12326,N_12458);
and U12665 (N_12665,N_12306,N_12309);
xnor U12666 (N_12666,N_12267,N_12301);
and U12667 (N_12667,N_12323,N_12394);
xor U12668 (N_12668,N_12324,N_12451);
and U12669 (N_12669,N_12268,N_12495);
xnor U12670 (N_12670,N_12431,N_12290);
nand U12671 (N_12671,N_12351,N_12328);
xor U12672 (N_12672,N_12391,N_12374);
nand U12673 (N_12673,N_12332,N_12343);
or U12674 (N_12674,N_12415,N_12372);
nand U12675 (N_12675,N_12389,N_12388);
nor U12676 (N_12676,N_12464,N_12298);
xor U12677 (N_12677,N_12261,N_12254);
nand U12678 (N_12678,N_12462,N_12439);
nor U12679 (N_12679,N_12258,N_12464);
xnor U12680 (N_12680,N_12375,N_12422);
xnor U12681 (N_12681,N_12465,N_12436);
xor U12682 (N_12682,N_12400,N_12288);
xor U12683 (N_12683,N_12496,N_12313);
nor U12684 (N_12684,N_12481,N_12388);
nor U12685 (N_12685,N_12258,N_12297);
and U12686 (N_12686,N_12441,N_12497);
nor U12687 (N_12687,N_12394,N_12491);
or U12688 (N_12688,N_12265,N_12306);
xor U12689 (N_12689,N_12439,N_12481);
and U12690 (N_12690,N_12453,N_12480);
nand U12691 (N_12691,N_12409,N_12451);
nand U12692 (N_12692,N_12279,N_12399);
nor U12693 (N_12693,N_12344,N_12454);
xnor U12694 (N_12694,N_12305,N_12250);
or U12695 (N_12695,N_12311,N_12459);
nand U12696 (N_12696,N_12299,N_12286);
or U12697 (N_12697,N_12470,N_12475);
nor U12698 (N_12698,N_12375,N_12347);
nand U12699 (N_12699,N_12486,N_12443);
nor U12700 (N_12700,N_12472,N_12378);
xnor U12701 (N_12701,N_12478,N_12296);
xnor U12702 (N_12702,N_12414,N_12266);
or U12703 (N_12703,N_12407,N_12384);
xnor U12704 (N_12704,N_12409,N_12482);
nor U12705 (N_12705,N_12333,N_12364);
xnor U12706 (N_12706,N_12442,N_12489);
and U12707 (N_12707,N_12288,N_12323);
or U12708 (N_12708,N_12406,N_12412);
and U12709 (N_12709,N_12388,N_12302);
xor U12710 (N_12710,N_12444,N_12298);
nand U12711 (N_12711,N_12397,N_12275);
nor U12712 (N_12712,N_12440,N_12431);
and U12713 (N_12713,N_12468,N_12294);
nor U12714 (N_12714,N_12318,N_12251);
or U12715 (N_12715,N_12292,N_12489);
and U12716 (N_12716,N_12273,N_12301);
xnor U12717 (N_12717,N_12479,N_12423);
and U12718 (N_12718,N_12378,N_12392);
or U12719 (N_12719,N_12427,N_12448);
xor U12720 (N_12720,N_12369,N_12498);
and U12721 (N_12721,N_12326,N_12479);
and U12722 (N_12722,N_12257,N_12486);
nor U12723 (N_12723,N_12473,N_12414);
or U12724 (N_12724,N_12440,N_12412);
nand U12725 (N_12725,N_12274,N_12335);
and U12726 (N_12726,N_12257,N_12304);
and U12727 (N_12727,N_12470,N_12462);
and U12728 (N_12728,N_12438,N_12490);
xor U12729 (N_12729,N_12328,N_12250);
xor U12730 (N_12730,N_12429,N_12315);
or U12731 (N_12731,N_12484,N_12310);
xor U12732 (N_12732,N_12337,N_12452);
and U12733 (N_12733,N_12478,N_12397);
nor U12734 (N_12734,N_12348,N_12302);
nor U12735 (N_12735,N_12391,N_12320);
nand U12736 (N_12736,N_12437,N_12415);
xnor U12737 (N_12737,N_12365,N_12452);
and U12738 (N_12738,N_12408,N_12337);
nand U12739 (N_12739,N_12364,N_12280);
xor U12740 (N_12740,N_12457,N_12376);
xnor U12741 (N_12741,N_12315,N_12257);
xnor U12742 (N_12742,N_12292,N_12290);
and U12743 (N_12743,N_12377,N_12490);
or U12744 (N_12744,N_12334,N_12417);
xnor U12745 (N_12745,N_12363,N_12331);
and U12746 (N_12746,N_12409,N_12441);
nand U12747 (N_12747,N_12337,N_12405);
xor U12748 (N_12748,N_12334,N_12497);
xor U12749 (N_12749,N_12367,N_12321);
or U12750 (N_12750,N_12643,N_12724);
nor U12751 (N_12751,N_12546,N_12631);
nor U12752 (N_12752,N_12659,N_12652);
nor U12753 (N_12753,N_12737,N_12644);
and U12754 (N_12754,N_12611,N_12610);
xnor U12755 (N_12755,N_12675,N_12674);
or U12756 (N_12756,N_12577,N_12678);
nand U12757 (N_12757,N_12542,N_12656);
and U12758 (N_12758,N_12607,N_12640);
nor U12759 (N_12759,N_12653,N_12556);
or U12760 (N_12760,N_12731,N_12595);
nand U12761 (N_12761,N_12541,N_12707);
and U12762 (N_12762,N_12633,N_12718);
nand U12763 (N_12763,N_12740,N_12580);
nand U12764 (N_12764,N_12635,N_12626);
nand U12765 (N_12765,N_12649,N_12594);
nand U12766 (N_12766,N_12584,N_12661);
xor U12767 (N_12767,N_12651,N_12690);
xnor U12768 (N_12768,N_12551,N_12598);
nor U12769 (N_12769,N_12572,N_12666);
nand U12770 (N_12770,N_12655,N_12641);
nand U12771 (N_12771,N_12713,N_12544);
or U12772 (N_12772,N_12732,N_12579);
nand U12773 (N_12773,N_12695,N_12744);
and U12774 (N_12774,N_12609,N_12711);
or U12775 (N_12775,N_12539,N_12712);
xnor U12776 (N_12776,N_12657,N_12543);
or U12777 (N_12777,N_12682,N_12574);
or U12778 (N_12778,N_12552,N_12683);
xor U12779 (N_12779,N_12538,N_12548);
and U12780 (N_12780,N_12701,N_12527);
or U12781 (N_12781,N_12523,N_12663);
nor U12782 (N_12782,N_12613,N_12619);
or U12783 (N_12783,N_12583,N_12746);
or U12784 (N_12784,N_12730,N_12600);
or U12785 (N_12785,N_12664,N_12559);
nand U12786 (N_12786,N_12634,N_12647);
and U12787 (N_12787,N_12535,N_12654);
nor U12788 (N_12788,N_12504,N_12508);
and U12789 (N_12789,N_12519,N_12608);
and U12790 (N_12790,N_12532,N_12662);
nor U12791 (N_12791,N_12747,N_12550);
nor U12792 (N_12792,N_12710,N_12540);
nand U12793 (N_12793,N_12554,N_12728);
xnor U12794 (N_12794,N_12720,N_12729);
and U12795 (N_12795,N_12517,N_12717);
and U12796 (N_12796,N_12603,N_12699);
xnor U12797 (N_12797,N_12526,N_12698);
xnor U12798 (N_12798,N_12599,N_12529);
and U12799 (N_12799,N_12697,N_12593);
and U12800 (N_12800,N_12560,N_12506);
xnor U12801 (N_12801,N_12692,N_12575);
nor U12802 (N_12802,N_12719,N_12505);
nor U12803 (N_12803,N_12734,N_12687);
nand U12804 (N_12804,N_12676,N_12503);
nand U12805 (N_12805,N_12709,N_12528);
xnor U12806 (N_12806,N_12624,N_12589);
xor U12807 (N_12807,N_12622,N_12512);
xnor U12808 (N_12808,N_12704,N_12563);
nor U12809 (N_12809,N_12537,N_12514);
nand U12810 (N_12810,N_12557,N_12629);
nor U12811 (N_12811,N_12642,N_12616);
or U12812 (N_12812,N_12545,N_12576);
or U12813 (N_12813,N_12587,N_12735);
and U12814 (N_12814,N_12650,N_12721);
xor U12815 (N_12815,N_12715,N_12614);
nand U12816 (N_12816,N_12502,N_12586);
nand U12817 (N_12817,N_12700,N_12590);
nand U12818 (N_12818,N_12568,N_12726);
xor U12819 (N_12819,N_12604,N_12671);
nand U12820 (N_12820,N_12620,N_12686);
xor U12821 (N_12821,N_12605,N_12684);
and U12822 (N_12822,N_12722,N_12628);
nand U12823 (N_12823,N_12667,N_12694);
or U12824 (N_12824,N_12708,N_12693);
and U12825 (N_12825,N_12520,N_12553);
and U12826 (N_12826,N_12591,N_12606);
and U12827 (N_12827,N_12705,N_12518);
nand U12828 (N_12828,N_12602,N_12696);
nor U12829 (N_12829,N_12547,N_12582);
nor U12830 (N_12830,N_12627,N_12688);
nor U12831 (N_12831,N_12534,N_12625);
nand U12832 (N_12832,N_12570,N_12585);
xnor U12833 (N_12833,N_12736,N_12509);
and U12834 (N_12834,N_12672,N_12536);
nand U12835 (N_12835,N_12516,N_12727);
or U12836 (N_12836,N_12562,N_12739);
xor U12837 (N_12837,N_12623,N_12743);
xnor U12838 (N_12838,N_12665,N_12742);
nand U12839 (N_12839,N_12525,N_12630);
and U12840 (N_12840,N_12564,N_12567);
nand U12841 (N_12841,N_12573,N_12617);
and U12842 (N_12842,N_12691,N_12549);
or U12843 (N_12843,N_12510,N_12648);
nand U12844 (N_12844,N_12615,N_12507);
xnor U12845 (N_12845,N_12632,N_12703);
or U12846 (N_12846,N_12501,N_12685);
and U12847 (N_12847,N_12565,N_12588);
xnor U12848 (N_12848,N_12515,N_12500);
xnor U12849 (N_12849,N_12702,N_12511);
nor U12850 (N_12850,N_12596,N_12578);
or U12851 (N_12851,N_12533,N_12660);
nand U12852 (N_12852,N_12592,N_12618);
nor U12853 (N_12853,N_12531,N_12677);
or U12854 (N_12854,N_12524,N_12749);
nand U12855 (N_12855,N_12680,N_12612);
or U12856 (N_12856,N_12714,N_12597);
xnor U12857 (N_12857,N_12716,N_12555);
or U12858 (N_12858,N_12558,N_12638);
and U12859 (N_12859,N_12513,N_12581);
nor U12860 (N_12860,N_12646,N_12741);
and U12861 (N_12861,N_12522,N_12637);
xor U12862 (N_12862,N_12669,N_12725);
or U12863 (N_12863,N_12601,N_12745);
nand U12864 (N_12864,N_12569,N_12561);
nand U12865 (N_12865,N_12658,N_12733);
nand U12866 (N_12866,N_12668,N_12681);
nand U12867 (N_12867,N_12521,N_12706);
nand U12868 (N_12868,N_12670,N_12689);
or U12869 (N_12869,N_12748,N_12679);
and U12870 (N_12870,N_12673,N_12636);
nand U12871 (N_12871,N_12639,N_12621);
or U12872 (N_12872,N_12566,N_12645);
xnor U12873 (N_12873,N_12738,N_12530);
nor U12874 (N_12874,N_12571,N_12723);
nor U12875 (N_12875,N_12740,N_12578);
or U12876 (N_12876,N_12598,N_12671);
and U12877 (N_12877,N_12745,N_12628);
xor U12878 (N_12878,N_12721,N_12686);
xnor U12879 (N_12879,N_12741,N_12652);
nor U12880 (N_12880,N_12597,N_12698);
nand U12881 (N_12881,N_12656,N_12675);
nand U12882 (N_12882,N_12511,N_12577);
nand U12883 (N_12883,N_12681,N_12618);
nor U12884 (N_12884,N_12617,N_12603);
nand U12885 (N_12885,N_12674,N_12551);
nor U12886 (N_12886,N_12598,N_12618);
xor U12887 (N_12887,N_12624,N_12668);
xor U12888 (N_12888,N_12707,N_12678);
and U12889 (N_12889,N_12515,N_12717);
xor U12890 (N_12890,N_12714,N_12525);
nor U12891 (N_12891,N_12659,N_12552);
nor U12892 (N_12892,N_12539,N_12737);
nand U12893 (N_12893,N_12660,N_12562);
or U12894 (N_12894,N_12591,N_12710);
nor U12895 (N_12895,N_12685,N_12539);
nor U12896 (N_12896,N_12517,N_12606);
nand U12897 (N_12897,N_12538,N_12727);
xor U12898 (N_12898,N_12662,N_12732);
or U12899 (N_12899,N_12673,N_12529);
nand U12900 (N_12900,N_12632,N_12504);
xor U12901 (N_12901,N_12666,N_12642);
nor U12902 (N_12902,N_12622,N_12587);
and U12903 (N_12903,N_12732,N_12700);
and U12904 (N_12904,N_12606,N_12544);
or U12905 (N_12905,N_12609,N_12634);
nand U12906 (N_12906,N_12566,N_12517);
or U12907 (N_12907,N_12509,N_12716);
xor U12908 (N_12908,N_12525,N_12571);
and U12909 (N_12909,N_12623,N_12656);
nor U12910 (N_12910,N_12655,N_12599);
nand U12911 (N_12911,N_12659,N_12630);
xor U12912 (N_12912,N_12597,N_12565);
or U12913 (N_12913,N_12679,N_12623);
nor U12914 (N_12914,N_12638,N_12521);
nand U12915 (N_12915,N_12544,N_12685);
or U12916 (N_12916,N_12621,N_12627);
xor U12917 (N_12917,N_12618,N_12670);
xnor U12918 (N_12918,N_12522,N_12724);
nor U12919 (N_12919,N_12561,N_12668);
and U12920 (N_12920,N_12525,N_12606);
xnor U12921 (N_12921,N_12654,N_12712);
and U12922 (N_12922,N_12685,N_12549);
xnor U12923 (N_12923,N_12516,N_12626);
and U12924 (N_12924,N_12543,N_12698);
xnor U12925 (N_12925,N_12555,N_12557);
nand U12926 (N_12926,N_12557,N_12568);
nor U12927 (N_12927,N_12566,N_12710);
xor U12928 (N_12928,N_12506,N_12612);
and U12929 (N_12929,N_12674,N_12593);
xnor U12930 (N_12930,N_12643,N_12522);
nand U12931 (N_12931,N_12686,N_12740);
and U12932 (N_12932,N_12701,N_12523);
and U12933 (N_12933,N_12669,N_12608);
or U12934 (N_12934,N_12527,N_12739);
nor U12935 (N_12935,N_12512,N_12708);
nor U12936 (N_12936,N_12592,N_12655);
and U12937 (N_12937,N_12611,N_12679);
and U12938 (N_12938,N_12539,N_12511);
nor U12939 (N_12939,N_12707,N_12523);
xnor U12940 (N_12940,N_12698,N_12707);
nor U12941 (N_12941,N_12687,N_12594);
and U12942 (N_12942,N_12551,N_12650);
or U12943 (N_12943,N_12723,N_12747);
nand U12944 (N_12944,N_12518,N_12695);
nand U12945 (N_12945,N_12645,N_12507);
or U12946 (N_12946,N_12566,N_12552);
nor U12947 (N_12947,N_12713,N_12574);
nand U12948 (N_12948,N_12682,N_12522);
xnor U12949 (N_12949,N_12631,N_12533);
nand U12950 (N_12950,N_12584,N_12720);
nor U12951 (N_12951,N_12655,N_12626);
or U12952 (N_12952,N_12563,N_12728);
or U12953 (N_12953,N_12671,N_12570);
nand U12954 (N_12954,N_12624,N_12656);
and U12955 (N_12955,N_12523,N_12537);
nand U12956 (N_12956,N_12619,N_12596);
xnor U12957 (N_12957,N_12590,N_12743);
nor U12958 (N_12958,N_12503,N_12601);
nor U12959 (N_12959,N_12561,N_12596);
and U12960 (N_12960,N_12619,N_12679);
or U12961 (N_12961,N_12737,N_12583);
and U12962 (N_12962,N_12690,N_12508);
xor U12963 (N_12963,N_12644,N_12529);
or U12964 (N_12964,N_12533,N_12724);
and U12965 (N_12965,N_12625,N_12666);
or U12966 (N_12966,N_12533,N_12521);
or U12967 (N_12967,N_12743,N_12658);
nand U12968 (N_12968,N_12565,N_12675);
or U12969 (N_12969,N_12739,N_12543);
xor U12970 (N_12970,N_12652,N_12552);
nor U12971 (N_12971,N_12529,N_12543);
nor U12972 (N_12972,N_12631,N_12529);
nand U12973 (N_12973,N_12630,N_12687);
and U12974 (N_12974,N_12687,N_12712);
nand U12975 (N_12975,N_12705,N_12629);
nand U12976 (N_12976,N_12549,N_12703);
nor U12977 (N_12977,N_12523,N_12591);
nand U12978 (N_12978,N_12543,N_12500);
or U12979 (N_12979,N_12698,N_12528);
or U12980 (N_12980,N_12737,N_12673);
nand U12981 (N_12981,N_12698,N_12535);
xnor U12982 (N_12982,N_12705,N_12662);
nor U12983 (N_12983,N_12520,N_12591);
or U12984 (N_12984,N_12550,N_12536);
or U12985 (N_12985,N_12703,N_12723);
or U12986 (N_12986,N_12673,N_12653);
nor U12987 (N_12987,N_12628,N_12546);
xnor U12988 (N_12988,N_12741,N_12727);
nand U12989 (N_12989,N_12580,N_12645);
nor U12990 (N_12990,N_12634,N_12575);
or U12991 (N_12991,N_12618,N_12622);
xor U12992 (N_12992,N_12560,N_12635);
or U12993 (N_12993,N_12675,N_12620);
xor U12994 (N_12994,N_12606,N_12743);
nand U12995 (N_12995,N_12583,N_12738);
and U12996 (N_12996,N_12655,N_12705);
or U12997 (N_12997,N_12658,N_12643);
xnor U12998 (N_12998,N_12655,N_12689);
xor U12999 (N_12999,N_12690,N_12704);
or U13000 (N_13000,N_12987,N_12954);
xnor U13001 (N_13001,N_12786,N_12760);
nor U13002 (N_13002,N_12836,N_12978);
or U13003 (N_13003,N_12977,N_12814);
xnor U13004 (N_13004,N_12888,N_12768);
nor U13005 (N_13005,N_12790,N_12754);
nor U13006 (N_13006,N_12798,N_12780);
and U13007 (N_13007,N_12809,N_12903);
and U13008 (N_13008,N_12924,N_12822);
nor U13009 (N_13009,N_12889,N_12803);
and U13010 (N_13010,N_12905,N_12956);
nand U13011 (N_13011,N_12761,N_12983);
xor U13012 (N_13012,N_12765,N_12864);
and U13013 (N_13013,N_12887,N_12883);
or U13014 (N_13014,N_12753,N_12784);
nor U13015 (N_13015,N_12936,N_12843);
or U13016 (N_13016,N_12929,N_12947);
and U13017 (N_13017,N_12797,N_12859);
nor U13018 (N_13018,N_12962,N_12823);
and U13019 (N_13019,N_12839,N_12853);
and U13020 (N_13020,N_12979,N_12937);
and U13021 (N_13021,N_12911,N_12908);
nand U13022 (N_13022,N_12826,N_12841);
and U13023 (N_13023,N_12831,N_12866);
or U13024 (N_13024,N_12981,N_12915);
xor U13025 (N_13025,N_12909,N_12871);
nand U13026 (N_13026,N_12821,N_12844);
or U13027 (N_13027,N_12945,N_12912);
nand U13028 (N_13028,N_12862,N_12818);
nand U13029 (N_13029,N_12923,N_12976);
nand U13030 (N_13030,N_12820,N_12852);
and U13031 (N_13031,N_12931,N_12840);
nand U13032 (N_13032,N_12833,N_12972);
or U13033 (N_13033,N_12904,N_12794);
nor U13034 (N_13034,N_12933,N_12914);
or U13035 (N_13035,N_12834,N_12763);
or U13036 (N_13036,N_12890,N_12957);
xnor U13037 (N_13037,N_12892,N_12764);
and U13038 (N_13038,N_12808,N_12785);
and U13039 (N_13039,N_12995,N_12845);
nor U13040 (N_13040,N_12932,N_12966);
nor U13041 (N_13041,N_12930,N_12848);
xor U13042 (N_13042,N_12921,N_12842);
and U13043 (N_13043,N_12992,N_12874);
or U13044 (N_13044,N_12771,N_12938);
nand U13045 (N_13045,N_12799,N_12813);
xnor U13046 (N_13046,N_12898,N_12916);
xor U13047 (N_13047,N_12854,N_12830);
nor U13048 (N_13048,N_12884,N_12880);
and U13049 (N_13049,N_12948,N_12944);
nor U13050 (N_13050,N_12800,N_12873);
nand U13051 (N_13051,N_12967,N_12939);
and U13052 (N_13052,N_12832,N_12829);
nor U13053 (N_13053,N_12778,N_12782);
nand U13054 (N_13054,N_12870,N_12913);
nand U13055 (N_13055,N_12949,N_12982);
nand U13056 (N_13056,N_12791,N_12825);
or U13057 (N_13057,N_12993,N_12922);
xnor U13058 (N_13058,N_12940,N_12867);
and U13059 (N_13059,N_12943,N_12868);
nand U13060 (N_13060,N_12918,N_12849);
nand U13061 (N_13061,N_12827,N_12787);
xor U13062 (N_13062,N_12877,N_12881);
and U13063 (N_13063,N_12824,N_12960);
and U13064 (N_13064,N_12838,N_12989);
xnor U13065 (N_13065,N_12958,N_12882);
or U13066 (N_13066,N_12899,N_12974);
or U13067 (N_13067,N_12774,N_12876);
nand U13068 (N_13068,N_12789,N_12946);
nor U13069 (N_13069,N_12807,N_12819);
nor U13070 (N_13070,N_12770,N_12997);
nand U13071 (N_13071,N_12920,N_12991);
or U13072 (N_13072,N_12769,N_12994);
or U13073 (N_13073,N_12773,N_12801);
and U13074 (N_13074,N_12886,N_12795);
xnor U13075 (N_13075,N_12863,N_12968);
nor U13076 (N_13076,N_12980,N_12767);
and U13077 (N_13077,N_12851,N_12896);
or U13078 (N_13078,N_12847,N_12788);
and U13079 (N_13079,N_12891,N_12855);
or U13080 (N_13080,N_12999,N_12828);
and U13081 (N_13081,N_12752,N_12919);
nand U13082 (N_13082,N_12781,N_12965);
and U13083 (N_13083,N_12893,N_12928);
xor U13084 (N_13084,N_12846,N_12941);
xnor U13085 (N_13085,N_12857,N_12996);
xnor U13086 (N_13086,N_12860,N_12806);
and U13087 (N_13087,N_12835,N_12772);
and U13088 (N_13088,N_12777,N_12776);
nand U13089 (N_13089,N_12988,N_12985);
or U13090 (N_13090,N_12906,N_12973);
nor U13091 (N_13091,N_12856,N_12804);
and U13092 (N_13092,N_12872,N_12775);
nor U13093 (N_13093,N_12757,N_12926);
nor U13094 (N_13094,N_12885,N_12984);
xor U13095 (N_13095,N_12766,N_12964);
xnor U13096 (N_13096,N_12812,N_12894);
nor U13097 (N_13097,N_12955,N_12837);
nand U13098 (N_13098,N_12751,N_12792);
xnor U13099 (N_13099,N_12961,N_12917);
and U13100 (N_13100,N_12758,N_12796);
nand U13101 (N_13101,N_12756,N_12969);
nand U13102 (N_13102,N_12953,N_12986);
nand U13103 (N_13103,N_12971,N_12895);
nand U13104 (N_13104,N_12998,N_12865);
nor U13105 (N_13105,N_12759,N_12805);
nand U13106 (N_13106,N_12750,N_12910);
nor U13107 (N_13107,N_12935,N_12990);
nor U13108 (N_13108,N_12815,N_12755);
or U13109 (N_13109,N_12942,N_12907);
nand U13110 (N_13110,N_12850,N_12875);
and U13111 (N_13111,N_12793,N_12963);
nor U13112 (N_13112,N_12927,N_12975);
nand U13113 (N_13113,N_12925,N_12950);
or U13114 (N_13114,N_12762,N_12879);
nand U13115 (N_13115,N_12878,N_12970);
nand U13116 (N_13116,N_12869,N_12900);
nand U13117 (N_13117,N_12952,N_12810);
nand U13118 (N_13118,N_12934,N_12902);
and U13119 (N_13119,N_12783,N_12816);
nor U13120 (N_13120,N_12811,N_12817);
or U13121 (N_13121,N_12901,N_12802);
and U13122 (N_13122,N_12858,N_12861);
nand U13123 (N_13123,N_12779,N_12959);
and U13124 (N_13124,N_12951,N_12897);
or U13125 (N_13125,N_12896,N_12964);
nand U13126 (N_13126,N_12854,N_12801);
and U13127 (N_13127,N_12817,N_12901);
or U13128 (N_13128,N_12817,N_12935);
or U13129 (N_13129,N_12787,N_12781);
nand U13130 (N_13130,N_12976,N_12885);
xnor U13131 (N_13131,N_12973,N_12892);
nand U13132 (N_13132,N_12882,N_12953);
or U13133 (N_13133,N_12842,N_12923);
or U13134 (N_13134,N_12890,N_12785);
nand U13135 (N_13135,N_12914,N_12997);
nand U13136 (N_13136,N_12920,N_12929);
xor U13137 (N_13137,N_12765,N_12866);
xnor U13138 (N_13138,N_12812,N_12882);
nand U13139 (N_13139,N_12838,N_12909);
and U13140 (N_13140,N_12970,N_12989);
nor U13141 (N_13141,N_12762,N_12794);
nand U13142 (N_13142,N_12858,N_12968);
or U13143 (N_13143,N_12825,N_12934);
nand U13144 (N_13144,N_12805,N_12864);
and U13145 (N_13145,N_12872,N_12780);
or U13146 (N_13146,N_12940,N_12929);
or U13147 (N_13147,N_12940,N_12799);
nand U13148 (N_13148,N_12811,N_12931);
xnor U13149 (N_13149,N_12889,N_12896);
and U13150 (N_13150,N_12999,N_12801);
nand U13151 (N_13151,N_12862,N_12755);
nor U13152 (N_13152,N_12884,N_12853);
and U13153 (N_13153,N_12956,N_12909);
xnor U13154 (N_13154,N_12885,N_12847);
xor U13155 (N_13155,N_12869,N_12967);
or U13156 (N_13156,N_12999,N_12866);
or U13157 (N_13157,N_12989,N_12798);
nand U13158 (N_13158,N_12775,N_12823);
or U13159 (N_13159,N_12889,N_12962);
nand U13160 (N_13160,N_12903,N_12912);
nor U13161 (N_13161,N_12780,N_12783);
nand U13162 (N_13162,N_12874,N_12810);
or U13163 (N_13163,N_12964,N_12876);
nand U13164 (N_13164,N_12976,N_12795);
or U13165 (N_13165,N_12790,N_12836);
nand U13166 (N_13166,N_12824,N_12838);
xnor U13167 (N_13167,N_12999,N_12815);
xnor U13168 (N_13168,N_12817,N_12822);
nand U13169 (N_13169,N_12915,N_12888);
or U13170 (N_13170,N_12823,N_12781);
or U13171 (N_13171,N_12816,N_12934);
or U13172 (N_13172,N_12955,N_12961);
xnor U13173 (N_13173,N_12967,N_12903);
xor U13174 (N_13174,N_12826,N_12830);
or U13175 (N_13175,N_12983,N_12776);
and U13176 (N_13176,N_12781,N_12907);
nor U13177 (N_13177,N_12998,N_12987);
or U13178 (N_13178,N_12777,N_12854);
nand U13179 (N_13179,N_12921,N_12811);
nand U13180 (N_13180,N_12806,N_12933);
xnor U13181 (N_13181,N_12941,N_12954);
or U13182 (N_13182,N_12979,N_12787);
and U13183 (N_13183,N_12875,N_12924);
nor U13184 (N_13184,N_12888,N_12830);
nor U13185 (N_13185,N_12977,N_12868);
nand U13186 (N_13186,N_12896,N_12919);
and U13187 (N_13187,N_12778,N_12926);
nor U13188 (N_13188,N_12970,N_12767);
nand U13189 (N_13189,N_12812,N_12800);
nand U13190 (N_13190,N_12907,N_12918);
nand U13191 (N_13191,N_12823,N_12798);
and U13192 (N_13192,N_12876,N_12973);
and U13193 (N_13193,N_12930,N_12816);
and U13194 (N_13194,N_12851,N_12919);
xor U13195 (N_13195,N_12871,N_12956);
and U13196 (N_13196,N_12784,N_12950);
xor U13197 (N_13197,N_12800,N_12831);
or U13198 (N_13198,N_12788,N_12887);
and U13199 (N_13199,N_12934,N_12759);
or U13200 (N_13200,N_12878,N_12903);
nor U13201 (N_13201,N_12796,N_12897);
nand U13202 (N_13202,N_12805,N_12764);
nand U13203 (N_13203,N_12809,N_12900);
and U13204 (N_13204,N_12821,N_12950);
or U13205 (N_13205,N_12945,N_12889);
nor U13206 (N_13206,N_12978,N_12802);
nand U13207 (N_13207,N_12856,N_12969);
and U13208 (N_13208,N_12888,N_12862);
nand U13209 (N_13209,N_12944,N_12865);
and U13210 (N_13210,N_12960,N_12790);
nor U13211 (N_13211,N_12910,N_12927);
or U13212 (N_13212,N_12913,N_12884);
nor U13213 (N_13213,N_12898,N_12879);
nor U13214 (N_13214,N_12906,N_12946);
xnor U13215 (N_13215,N_12764,N_12913);
nand U13216 (N_13216,N_12941,N_12928);
or U13217 (N_13217,N_12821,N_12778);
nor U13218 (N_13218,N_12883,N_12853);
xnor U13219 (N_13219,N_12888,N_12884);
or U13220 (N_13220,N_12755,N_12880);
or U13221 (N_13221,N_12969,N_12980);
nor U13222 (N_13222,N_12777,N_12927);
nor U13223 (N_13223,N_12965,N_12917);
or U13224 (N_13224,N_12879,N_12946);
and U13225 (N_13225,N_12757,N_12959);
or U13226 (N_13226,N_12931,N_12852);
or U13227 (N_13227,N_12963,N_12846);
or U13228 (N_13228,N_12807,N_12912);
nand U13229 (N_13229,N_12930,N_12939);
nand U13230 (N_13230,N_12786,N_12962);
or U13231 (N_13231,N_12961,N_12845);
and U13232 (N_13232,N_12945,N_12941);
and U13233 (N_13233,N_12931,N_12865);
or U13234 (N_13234,N_12991,N_12842);
and U13235 (N_13235,N_12923,N_12796);
nor U13236 (N_13236,N_12981,N_12780);
or U13237 (N_13237,N_12773,N_12835);
nand U13238 (N_13238,N_12851,N_12924);
nand U13239 (N_13239,N_12945,N_12943);
or U13240 (N_13240,N_12977,N_12941);
and U13241 (N_13241,N_12844,N_12920);
nand U13242 (N_13242,N_12750,N_12849);
and U13243 (N_13243,N_12786,N_12797);
or U13244 (N_13244,N_12845,N_12969);
or U13245 (N_13245,N_12926,N_12867);
xor U13246 (N_13246,N_12872,N_12754);
nand U13247 (N_13247,N_12756,N_12888);
xor U13248 (N_13248,N_12907,N_12807);
nor U13249 (N_13249,N_12821,N_12776);
nor U13250 (N_13250,N_13067,N_13145);
or U13251 (N_13251,N_13182,N_13209);
or U13252 (N_13252,N_13000,N_13138);
or U13253 (N_13253,N_13035,N_13133);
nand U13254 (N_13254,N_13164,N_13108);
or U13255 (N_13255,N_13063,N_13029);
xor U13256 (N_13256,N_13070,N_13012);
xor U13257 (N_13257,N_13093,N_13077);
nand U13258 (N_13258,N_13002,N_13064);
nand U13259 (N_13259,N_13230,N_13191);
nor U13260 (N_13260,N_13197,N_13105);
xor U13261 (N_13261,N_13073,N_13054);
nand U13262 (N_13262,N_13192,N_13090);
xor U13263 (N_13263,N_13226,N_13113);
and U13264 (N_13264,N_13058,N_13129);
nand U13265 (N_13265,N_13050,N_13086);
nand U13266 (N_13266,N_13109,N_13183);
and U13267 (N_13267,N_13205,N_13084);
xnor U13268 (N_13268,N_13136,N_13008);
nor U13269 (N_13269,N_13114,N_13224);
nor U13270 (N_13270,N_13082,N_13166);
nand U13271 (N_13271,N_13232,N_13227);
xnor U13272 (N_13272,N_13185,N_13229);
xnor U13273 (N_13273,N_13017,N_13184);
nand U13274 (N_13274,N_13053,N_13047);
xor U13275 (N_13275,N_13112,N_13195);
or U13276 (N_13276,N_13021,N_13228);
xor U13277 (N_13277,N_13031,N_13141);
and U13278 (N_13278,N_13171,N_13236);
xor U13279 (N_13279,N_13135,N_13121);
nand U13280 (N_13280,N_13103,N_13152);
xor U13281 (N_13281,N_13083,N_13239);
xor U13282 (N_13282,N_13242,N_13179);
nor U13283 (N_13283,N_13009,N_13019);
nor U13284 (N_13284,N_13099,N_13231);
and U13285 (N_13285,N_13010,N_13092);
nand U13286 (N_13286,N_13217,N_13087);
xnor U13287 (N_13287,N_13127,N_13215);
nand U13288 (N_13288,N_13049,N_13162);
nand U13289 (N_13289,N_13204,N_13167);
or U13290 (N_13290,N_13023,N_13212);
nor U13291 (N_13291,N_13168,N_13153);
xnor U13292 (N_13292,N_13072,N_13174);
and U13293 (N_13293,N_13024,N_13188);
or U13294 (N_13294,N_13071,N_13196);
and U13295 (N_13295,N_13249,N_13040);
xor U13296 (N_13296,N_13225,N_13187);
xnor U13297 (N_13297,N_13006,N_13078);
and U13298 (N_13298,N_13115,N_13247);
or U13299 (N_13299,N_13007,N_13235);
or U13300 (N_13300,N_13246,N_13101);
or U13301 (N_13301,N_13146,N_13213);
or U13302 (N_13302,N_13016,N_13038);
nand U13303 (N_13303,N_13122,N_13085);
xnor U13304 (N_13304,N_13223,N_13243);
and U13305 (N_13305,N_13181,N_13199);
xor U13306 (N_13306,N_13044,N_13148);
nor U13307 (N_13307,N_13045,N_13154);
xnor U13308 (N_13308,N_13068,N_13005);
nor U13309 (N_13309,N_13140,N_13046);
and U13310 (N_13310,N_13074,N_13159);
nand U13311 (N_13311,N_13248,N_13139);
nor U13312 (N_13312,N_13222,N_13052);
and U13313 (N_13313,N_13116,N_13094);
nand U13314 (N_13314,N_13175,N_13028);
nand U13315 (N_13315,N_13033,N_13208);
xor U13316 (N_13316,N_13219,N_13111);
and U13317 (N_13317,N_13034,N_13206);
and U13318 (N_13318,N_13124,N_13169);
nand U13319 (N_13319,N_13080,N_13027);
nand U13320 (N_13320,N_13014,N_13118);
and U13321 (N_13321,N_13170,N_13055);
and U13322 (N_13322,N_13151,N_13075);
nand U13323 (N_13323,N_13155,N_13131);
nand U13324 (N_13324,N_13081,N_13123);
xor U13325 (N_13325,N_13020,N_13180);
or U13326 (N_13326,N_13200,N_13061);
xor U13327 (N_13327,N_13041,N_13233);
or U13328 (N_13328,N_13186,N_13143);
xor U13329 (N_13329,N_13237,N_13158);
xnor U13330 (N_13330,N_13126,N_13190);
or U13331 (N_13331,N_13176,N_13178);
and U13332 (N_13332,N_13095,N_13194);
nor U13333 (N_13333,N_13244,N_13102);
or U13334 (N_13334,N_13234,N_13004);
or U13335 (N_13335,N_13032,N_13240);
and U13336 (N_13336,N_13089,N_13100);
and U13337 (N_13337,N_13091,N_13051);
nor U13338 (N_13338,N_13193,N_13043);
xor U13339 (N_13339,N_13001,N_13156);
nand U13340 (N_13340,N_13098,N_13202);
or U13341 (N_13341,N_13048,N_13241);
and U13342 (N_13342,N_13039,N_13128);
or U13343 (N_13343,N_13037,N_13218);
or U13344 (N_13344,N_13201,N_13238);
xor U13345 (N_13345,N_13104,N_13211);
xor U13346 (N_13346,N_13110,N_13069);
nor U13347 (N_13347,N_13157,N_13198);
xor U13348 (N_13348,N_13216,N_13207);
nand U13349 (N_13349,N_13062,N_13214);
or U13350 (N_13350,N_13022,N_13134);
nor U13351 (N_13351,N_13056,N_13160);
or U13352 (N_13352,N_13130,N_13142);
and U13353 (N_13353,N_13013,N_13163);
or U13354 (N_13354,N_13210,N_13117);
nor U13355 (N_13355,N_13079,N_13189);
or U13356 (N_13356,N_13107,N_13106);
or U13357 (N_13357,N_13076,N_13132);
and U13358 (N_13358,N_13161,N_13220);
nand U13359 (N_13359,N_13026,N_13096);
or U13360 (N_13360,N_13150,N_13120);
and U13361 (N_13361,N_13057,N_13030);
or U13362 (N_13362,N_13003,N_13042);
nor U13363 (N_13363,N_13245,N_13173);
nor U13364 (N_13364,N_13203,N_13172);
nor U13365 (N_13365,N_13137,N_13036);
nand U13366 (N_13366,N_13149,N_13011);
xor U13367 (N_13367,N_13015,N_13125);
nor U13368 (N_13368,N_13060,N_13147);
or U13369 (N_13369,N_13097,N_13066);
nand U13370 (N_13370,N_13065,N_13088);
and U13371 (N_13371,N_13059,N_13119);
or U13372 (N_13372,N_13025,N_13221);
xnor U13373 (N_13373,N_13165,N_13177);
nand U13374 (N_13374,N_13144,N_13018);
nor U13375 (N_13375,N_13127,N_13227);
nand U13376 (N_13376,N_13096,N_13040);
nor U13377 (N_13377,N_13117,N_13014);
nor U13378 (N_13378,N_13031,N_13137);
nor U13379 (N_13379,N_13030,N_13083);
and U13380 (N_13380,N_13159,N_13180);
nor U13381 (N_13381,N_13196,N_13088);
xnor U13382 (N_13382,N_13051,N_13070);
nor U13383 (N_13383,N_13027,N_13161);
nor U13384 (N_13384,N_13073,N_13077);
and U13385 (N_13385,N_13159,N_13022);
or U13386 (N_13386,N_13112,N_13086);
or U13387 (N_13387,N_13002,N_13165);
nand U13388 (N_13388,N_13246,N_13008);
nand U13389 (N_13389,N_13005,N_13133);
nand U13390 (N_13390,N_13107,N_13231);
nor U13391 (N_13391,N_13121,N_13015);
or U13392 (N_13392,N_13244,N_13213);
xnor U13393 (N_13393,N_13022,N_13114);
xnor U13394 (N_13394,N_13244,N_13093);
and U13395 (N_13395,N_13036,N_13078);
or U13396 (N_13396,N_13018,N_13166);
or U13397 (N_13397,N_13249,N_13011);
nand U13398 (N_13398,N_13148,N_13007);
nand U13399 (N_13399,N_13100,N_13043);
nand U13400 (N_13400,N_13203,N_13246);
xnor U13401 (N_13401,N_13001,N_13135);
nor U13402 (N_13402,N_13061,N_13150);
xor U13403 (N_13403,N_13084,N_13131);
nand U13404 (N_13404,N_13217,N_13001);
nand U13405 (N_13405,N_13175,N_13033);
nor U13406 (N_13406,N_13018,N_13020);
xnor U13407 (N_13407,N_13184,N_13127);
nor U13408 (N_13408,N_13158,N_13046);
or U13409 (N_13409,N_13015,N_13067);
xnor U13410 (N_13410,N_13160,N_13088);
and U13411 (N_13411,N_13056,N_13205);
and U13412 (N_13412,N_13004,N_13014);
or U13413 (N_13413,N_13106,N_13058);
nor U13414 (N_13414,N_13087,N_13003);
xor U13415 (N_13415,N_13214,N_13012);
xor U13416 (N_13416,N_13009,N_13226);
or U13417 (N_13417,N_13003,N_13117);
or U13418 (N_13418,N_13141,N_13195);
or U13419 (N_13419,N_13043,N_13091);
nor U13420 (N_13420,N_13045,N_13007);
or U13421 (N_13421,N_13007,N_13202);
nand U13422 (N_13422,N_13029,N_13003);
nand U13423 (N_13423,N_13208,N_13070);
nand U13424 (N_13424,N_13045,N_13000);
xor U13425 (N_13425,N_13044,N_13246);
and U13426 (N_13426,N_13000,N_13085);
or U13427 (N_13427,N_13162,N_13192);
nor U13428 (N_13428,N_13191,N_13221);
xor U13429 (N_13429,N_13236,N_13201);
or U13430 (N_13430,N_13166,N_13059);
or U13431 (N_13431,N_13172,N_13013);
nor U13432 (N_13432,N_13060,N_13067);
or U13433 (N_13433,N_13008,N_13031);
nand U13434 (N_13434,N_13110,N_13232);
xnor U13435 (N_13435,N_13134,N_13057);
nand U13436 (N_13436,N_13097,N_13035);
xor U13437 (N_13437,N_13190,N_13151);
nor U13438 (N_13438,N_13143,N_13247);
and U13439 (N_13439,N_13205,N_13127);
or U13440 (N_13440,N_13204,N_13025);
xnor U13441 (N_13441,N_13086,N_13146);
and U13442 (N_13442,N_13141,N_13051);
nand U13443 (N_13443,N_13142,N_13200);
or U13444 (N_13444,N_13085,N_13134);
nand U13445 (N_13445,N_13054,N_13124);
and U13446 (N_13446,N_13230,N_13008);
nor U13447 (N_13447,N_13159,N_13038);
xor U13448 (N_13448,N_13245,N_13044);
xnor U13449 (N_13449,N_13191,N_13086);
and U13450 (N_13450,N_13196,N_13126);
and U13451 (N_13451,N_13042,N_13171);
xor U13452 (N_13452,N_13193,N_13156);
nor U13453 (N_13453,N_13068,N_13108);
xor U13454 (N_13454,N_13183,N_13058);
xnor U13455 (N_13455,N_13201,N_13039);
and U13456 (N_13456,N_13103,N_13025);
xnor U13457 (N_13457,N_13249,N_13074);
and U13458 (N_13458,N_13114,N_13196);
xnor U13459 (N_13459,N_13117,N_13144);
or U13460 (N_13460,N_13052,N_13056);
nor U13461 (N_13461,N_13038,N_13145);
nand U13462 (N_13462,N_13107,N_13126);
or U13463 (N_13463,N_13059,N_13182);
nor U13464 (N_13464,N_13179,N_13013);
and U13465 (N_13465,N_13039,N_13024);
or U13466 (N_13466,N_13000,N_13197);
xor U13467 (N_13467,N_13229,N_13066);
or U13468 (N_13468,N_13195,N_13144);
and U13469 (N_13469,N_13048,N_13039);
and U13470 (N_13470,N_13145,N_13161);
nand U13471 (N_13471,N_13156,N_13030);
nand U13472 (N_13472,N_13238,N_13023);
nand U13473 (N_13473,N_13132,N_13189);
nor U13474 (N_13474,N_13177,N_13080);
xor U13475 (N_13475,N_13156,N_13013);
and U13476 (N_13476,N_13236,N_13009);
xnor U13477 (N_13477,N_13041,N_13159);
nor U13478 (N_13478,N_13190,N_13062);
nor U13479 (N_13479,N_13153,N_13142);
nand U13480 (N_13480,N_13086,N_13043);
nor U13481 (N_13481,N_13022,N_13121);
and U13482 (N_13482,N_13051,N_13181);
nor U13483 (N_13483,N_13019,N_13160);
nand U13484 (N_13484,N_13128,N_13158);
nor U13485 (N_13485,N_13084,N_13225);
nor U13486 (N_13486,N_13176,N_13222);
or U13487 (N_13487,N_13023,N_13147);
and U13488 (N_13488,N_13238,N_13234);
or U13489 (N_13489,N_13050,N_13212);
or U13490 (N_13490,N_13192,N_13222);
nor U13491 (N_13491,N_13248,N_13094);
and U13492 (N_13492,N_13190,N_13096);
nor U13493 (N_13493,N_13065,N_13025);
or U13494 (N_13494,N_13164,N_13201);
xor U13495 (N_13495,N_13084,N_13080);
or U13496 (N_13496,N_13060,N_13142);
xor U13497 (N_13497,N_13102,N_13191);
nand U13498 (N_13498,N_13133,N_13095);
and U13499 (N_13499,N_13245,N_13226);
and U13500 (N_13500,N_13414,N_13365);
xnor U13501 (N_13501,N_13324,N_13326);
and U13502 (N_13502,N_13296,N_13336);
nand U13503 (N_13503,N_13449,N_13377);
and U13504 (N_13504,N_13343,N_13445);
nand U13505 (N_13505,N_13436,N_13468);
and U13506 (N_13506,N_13390,N_13293);
nand U13507 (N_13507,N_13359,N_13423);
nand U13508 (N_13508,N_13415,N_13300);
or U13509 (N_13509,N_13405,N_13430);
and U13510 (N_13510,N_13346,N_13372);
xnor U13511 (N_13511,N_13478,N_13354);
nand U13512 (N_13512,N_13317,N_13490);
nor U13513 (N_13513,N_13328,N_13371);
nor U13514 (N_13514,N_13435,N_13498);
xnor U13515 (N_13515,N_13404,N_13262);
xor U13516 (N_13516,N_13442,N_13374);
or U13517 (N_13517,N_13261,N_13484);
xnor U13518 (N_13518,N_13408,N_13489);
nor U13519 (N_13519,N_13320,N_13264);
or U13520 (N_13520,N_13287,N_13376);
or U13521 (N_13521,N_13274,N_13389);
xnor U13522 (N_13522,N_13263,N_13378);
or U13523 (N_13523,N_13322,N_13416);
nor U13524 (N_13524,N_13422,N_13411);
and U13525 (N_13525,N_13480,N_13494);
and U13526 (N_13526,N_13323,N_13309);
and U13527 (N_13527,N_13310,N_13260);
or U13528 (N_13528,N_13339,N_13410);
xor U13529 (N_13529,N_13402,N_13453);
nand U13530 (N_13530,N_13294,N_13265);
or U13531 (N_13531,N_13426,N_13458);
xor U13532 (N_13532,N_13456,N_13470);
and U13533 (N_13533,N_13252,N_13318);
nor U13534 (N_13534,N_13403,N_13362);
nor U13535 (N_13535,N_13392,N_13454);
nor U13536 (N_13536,N_13434,N_13305);
nand U13537 (N_13537,N_13394,N_13387);
and U13538 (N_13538,N_13283,N_13462);
nand U13539 (N_13539,N_13427,N_13363);
xnor U13540 (N_13540,N_13250,N_13255);
and U13541 (N_13541,N_13425,N_13257);
nor U13542 (N_13542,N_13353,N_13472);
nor U13543 (N_13543,N_13474,N_13492);
nor U13544 (N_13544,N_13461,N_13373);
xor U13545 (N_13545,N_13301,N_13455);
nor U13546 (N_13546,N_13497,N_13340);
nand U13547 (N_13547,N_13382,N_13496);
nand U13548 (N_13548,N_13285,N_13348);
and U13549 (N_13549,N_13443,N_13441);
and U13550 (N_13550,N_13417,N_13401);
or U13551 (N_13551,N_13447,N_13483);
nor U13552 (N_13552,N_13457,N_13380);
xor U13553 (N_13553,N_13428,N_13407);
nor U13554 (N_13554,N_13276,N_13491);
nor U13555 (N_13555,N_13463,N_13286);
and U13556 (N_13556,N_13406,N_13440);
or U13557 (N_13557,N_13412,N_13475);
nand U13558 (N_13558,N_13292,N_13493);
or U13559 (N_13559,N_13476,N_13269);
or U13560 (N_13560,N_13393,N_13288);
or U13561 (N_13561,N_13295,N_13280);
nor U13562 (N_13562,N_13289,N_13367);
and U13563 (N_13563,N_13381,N_13277);
nand U13564 (N_13564,N_13379,N_13333);
nand U13565 (N_13565,N_13281,N_13312);
or U13566 (N_13566,N_13388,N_13334);
or U13567 (N_13567,N_13444,N_13477);
nor U13568 (N_13568,N_13398,N_13421);
nand U13569 (N_13569,N_13375,N_13298);
nand U13570 (N_13570,N_13448,N_13306);
or U13571 (N_13571,N_13256,N_13383);
nor U13572 (N_13572,N_13345,N_13357);
xnor U13573 (N_13573,N_13327,N_13400);
nand U13574 (N_13574,N_13251,N_13438);
nand U13575 (N_13575,N_13271,N_13282);
xor U13576 (N_13576,N_13465,N_13429);
or U13577 (N_13577,N_13495,N_13499);
and U13578 (N_13578,N_13433,N_13284);
nand U13579 (N_13579,N_13337,N_13291);
xnor U13580 (N_13580,N_13473,N_13330);
nand U13581 (N_13581,N_13409,N_13308);
nand U13582 (N_13582,N_13267,N_13259);
xnor U13583 (N_13583,N_13360,N_13395);
nor U13584 (N_13584,N_13299,N_13446);
xor U13585 (N_13585,N_13464,N_13303);
nand U13586 (N_13586,N_13278,N_13397);
xor U13587 (N_13587,N_13467,N_13342);
nor U13588 (N_13588,N_13486,N_13266);
xnor U13589 (N_13589,N_13431,N_13471);
and U13590 (N_13590,N_13419,N_13418);
nand U13591 (N_13591,N_13451,N_13344);
or U13592 (N_13592,N_13459,N_13460);
and U13593 (N_13593,N_13349,N_13368);
or U13594 (N_13594,N_13297,N_13335);
nor U13595 (N_13595,N_13352,N_13313);
xnor U13596 (N_13596,N_13258,N_13314);
xor U13597 (N_13597,N_13254,N_13439);
or U13598 (N_13598,N_13432,N_13332);
nand U13599 (N_13599,N_13355,N_13479);
or U13600 (N_13600,N_13290,N_13485);
nor U13601 (N_13601,N_13279,N_13307);
nand U13602 (N_13602,N_13391,N_13350);
nor U13603 (N_13603,N_13396,N_13356);
nor U13604 (N_13604,N_13272,N_13329);
xnor U13605 (N_13605,N_13316,N_13452);
xnor U13606 (N_13606,N_13424,N_13386);
nand U13607 (N_13607,N_13325,N_13315);
or U13608 (N_13608,N_13370,N_13481);
and U13609 (N_13609,N_13275,N_13273);
nor U13610 (N_13610,N_13361,N_13321);
nand U13611 (N_13611,N_13253,N_13331);
or U13612 (N_13612,N_13487,N_13347);
nand U13613 (N_13613,N_13369,N_13302);
nor U13614 (N_13614,N_13385,N_13366);
and U13615 (N_13615,N_13469,N_13319);
xor U13616 (N_13616,N_13270,N_13311);
and U13617 (N_13617,N_13364,N_13466);
nor U13618 (N_13618,N_13341,N_13420);
nor U13619 (N_13619,N_13482,N_13338);
and U13620 (N_13620,N_13351,N_13384);
and U13621 (N_13621,N_13304,N_13358);
or U13622 (N_13622,N_13488,N_13399);
xor U13623 (N_13623,N_13413,N_13268);
or U13624 (N_13624,N_13437,N_13450);
xor U13625 (N_13625,N_13262,N_13497);
nor U13626 (N_13626,N_13372,N_13275);
nor U13627 (N_13627,N_13318,N_13259);
nor U13628 (N_13628,N_13282,N_13410);
nor U13629 (N_13629,N_13437,N_13426);
or U13630 (N_13630,N_13465,N_13307);
xnor U13631 (N_13631,N_13347,N_13376);
xnor U13632 (N_13632,N_13403,N_13266);
nor U13633 (N_13633,N_13421,N_13304);
nor U13634 (N_13634,N_13328,N_13298);
and U13635 (N_13635,N_13344,N_13407);
or U13636 (N_13636,N_13454,N_13389);
or U13637 (N_13637,N_13418,N_13264);
and U13638 (N_13638,N_13455,N_13447);
and U13639 (N_13639,N_13405,N_13274);
nand U13640 (N_13640,N_13434,N_13287);
or U13641 (N_13641,N_13263,N_13343);
nor U13642 (N_13642,N_13421,N_13419);
or U13643 (N_13643,N_13415,N_13451);
or U13644 (N_13644,N_13333,N_13290);
nor U13645 (N_13645,N_13355,N_13415);
or U13646 (N_13646,N_13488,N_13323);
and U13647 (N_13647,N_13320,N_13392);
xor U13648 (N_13648,N_13340,N_13448);
nor U13649 (N_13649,N_13277,N_13378);
and U13650 (N_13650,N_13379,N_13366);
nor U13651 (N_13651,N_13258,N_13441);
nand U13652 (N_13652,N_13456,N_13357);
and U13653 (N_13653,N_13271,N_13477);
or U13654 (N_13654,N_13332,N_13314);
xnor U13655 (N_13655,N_13452,N_13455);
and U13656 (N_13656,N_13426,N_13288);
nor U13657 (N_13657,N_13405,N_13273);
nand U13658 (N_13658,N_13454,N_13321);
nor U13659 (N_13659,N_13332,N_13259);
or U13660 (N_13660,N_13408,N_13462);
xnor U13661 (N_13661,N_13396,N_13388);
nor U13662 (N_13662,N_13275,N_13485);
or U13663 (N_13663,N_13351,N_13257);
nand U13664 (N_13664,N_13425,N_13452);
nor U13665 (N_13665,N_13389,N_13426);
xor U13666 (N_13666,N_13402,N_13455);
xor U13667 (N_13667,N_13321,N_13366);
and U13668 (N_13668,N_13444,N_13457);
nand U13669 (N_13669,N_13409,N_13262);
and U13670 (N_13670,N_13324,N_13361);
or U13671 (N_13671,N_13275,N_13439);
or U13672 (N_13672,N_13260,N_13328);
xor U13673 (N_13673,N_13380,N_13433);
and U13674 (N_13674,N_13310,N_13415);
xor U13675 (N_13675,N_13474,N_13418);
xor U13676 (N_13676,N_13282,N_13307);
xor U13677 (N_13677,N_13348,N_13352);
nand U13678 (N_13678,N_13301,N_13287);
or U13679 (N_13679,N_13410,N_13485);
nor U13680 (N_13680,N_13471,N_13277);
nor U13681 (N_13681,N_13414,N_13339);
and U13682 (N_13682,N_13325,N_13412);
nor U13683 (N_13683,N_13340,N_13381);
and U13684 (N_13684,N_13370,N_13304);
xor U13685 (N_13685,N_13373,N_13326);
nor U13686 (N_13686,N_13332,N_13390);
or U13687 (N_13687,N_13308,N_13292);
xnor U13688 (N_13688,N_13453,N_13370);
and U13689 (N_13689,N_13400,N_13317);
or U13690 (N_13690,N_13456,N_13410);
or U13691 (N_13691,N_13461,N_13289);
nand U13692 (N_13692,N_13483,N_13322);
xor U13693 (N_13693,N_13398,N_13476);
xnor U13694 (N_13694,N_13372,N_13348);
xnor U13695 (N_13695,N_13368,N_13419);
and U13696 (N_13696,N_13355,N_13335);
nor U13697 (N_13697,N_13265,N_13499);
xnor U13698 (N_13698,N_13330,N_13257);
nor U13699 (N_13699,N_13310,N_13361);
and U13700 (N_13700,N_13262,N_13259);
nor U13701 (N_13701,N_13421,N_13491);
nand U13702 (N_13702,N_13400,N_13459);
nor U13703 (N_13703,N_13354,N_13355);
nand U13704 (N_13704,N_13308,N_13475);
or U13705 (N_13705,N_13465,N_13342);
nand U13706 (N_13706,N_13384,N_13261);
and U13707 (N_13707,N_13483,N_13381);
and U13708 (N_13708,N_13490,N_13440);
or U13709 (N_13709,N_13401,N_13415);
or U13710 (N_13710,N_13418,N_13292);
nor U13711 (N_13711,N_13309,N_13466);
nand U13712 (N_13712,N_13360,N_13493);
or U13713 (N_13713,N_13410,N_13457);
nor U13714 (N_13714,N_13301,N_13300);
and U13715 (N_13715,N_13352,N_13276);
and U13716 (N_13716,N_13403,N_13305);
or U13717 (N_13717,N_13413,N_13331);
xor U13718 (N_13718,N_13366,N_13315);
nor U13719 (N_13719,N_13375,N_13441);
nand U13720 (N_13720,N_13300,N_13309);
and U13721 (N_13721,N_13482,N_13479);
xnor U13722 (N_13722,N_13285,N_13301);
xor U13723 (N_13723,N_13352,N_13472);
and U13724 (N_13724,N_13326,N_13438);
or U13725 (N_13725,N_13352,N_13279);
nand U13726 (N_13726,N_13478,N_13293);
or U13727 (N_13727,N_13364,N_13422);
and U13728 (N_13728,N_13422,N_13496);
and U13729 (N_13729,N_13361,N_13370);
or U13730 (N_13730,N_13393,N_13495);
and U13731 (N_13731,N_13290,N_13271);
xor U13732 (N_13732,N_13482,N_13488);
xnor U13733 (N_13733,N_13466,N_13422);
or U13734 (N_13734,N_13292,N_13267);
xor U13735 (N_13735,N_13365,N_13434);
or U13736 (N_13736,N_13400,N_13264);
nor U13737 (N_13737,N_13461,N_13434);
or U13738 (N_13738,N_13406,N_13284);
xor U13739 (N_13739,N_13493,N_13288);
xnor U13740 (N_13740,N_13373,N_13302);
or U13741 (N_13741,N_13407,N_13255);
and U13742 (N_13742,N_13307,N_13439);
and U13743 (N_13743,N_13273,N_13385);
or U13744 (N_13744,N_13406,N_13456);
and U13745 (N_13745,N_13455,N_13403);
or U13746 (N_13746,N_13361,N_13294);
xnor U13747 (N_13747,N_13413,N_13385);
nor U13748 (N_13748,N_13302,N_13401);
and U13749 (N_13749,N_13308,N_13284);
xnor U13750 (N_13750,N_13685,N_13717);
and U13751 (N_13751,N_13525,N_13603);
xnor U13752 (N_13752,N_13719,N_13690);
nand U13753 (N_13753,N_13732,N_13671);
nand U13754 (N_13754,N_13625,N_13540);
and U13755 (N_13755,N_13512,N_13569);
and U13756 (N_13756,N_13749,N_13709);
and U13757 (N_13757,N_13500,N_13530);
or U13758 (N_13758,N_13707,N_13579);
nand U13759 (N_13759,N_13616,N_13511);
and U13760 (N_13760,N_13740,N_13651);
xor U13761 (N_13761,N_13666,N_13661);
nor U13762 (N_13762,N_13515,N_13593);
or U13763 (N_13763,N_13665,N_13710);
nor U13764 (N_13764,N_13712,N_13583);
or U13765 (N_13765,N_13574,N_13708);
nor U13766 (N_13766,N_13509,N_13586);
or U13767 (N_13767,N_13736,N_13532);
nor U13768 (N_13768,N_13571,N_13675);
or U13769 (N_13769,N_13611,N_13597);
nor U13770 (N_13770,N_13513,N_13562);
nand U13771 (N_13771,N_13702,N_13678);
xnor U13772 (N_13772,N_13699,N_13522);
nor U13773 (N_13773,N_13725,N_13563);
nand U13774 (N_13774,N_13703,N_13738);
and U13775 (N_13775,N_13589,N_13682);
and U13776 (N_13776,N_13565,N_13731);
nand U13777 (N_13777,N_13559,N_13581);
or U13778 (N_13778,N_13729,N_13693);
or U13779 (N_13779,N_13692,N_13573);
nand U13780 (N_13780,N_13668,N_13646);
nor U13781 (N_13781,N_13541,N_13592);
and U13782 (N_13782,N_13686,N_13608);
or U13783 (N_13783,N_13560,N_13526);
nand U13784 (N_13784,N_13676,N_13544);
xor U13785 (N_13785,N_13527,N_13720);
nor U13786 (N_13786,N_13727,N_13683);
xor U13787 (N_13787,N_13715,N_13529);
nand U13788 (N_13788,N_13714,N_13663);
nand U13789 (N_13789,N_13730,N_13572);
nor U13790 (N_13790,N_13520,N_13590);
xor U13791 (N_13791,N_13582,N_13548);
nor U13792 (N_13792,N_13672,N_13722);
xnor U13793 (N_13793,N_13609,N_13735);
xnor U13794 (N_13794,N_13521,N_13612);
or U13795 (N_13795,N_13704,N_13652);
nand U13796 (N_13796,N_13568,N_13687);
nor U13797 (N_13797,N_13524,N_13543);
nor U13798 (N_13798,N_13649,N_13564);
and U13799 (N_13799,N_13528,N_13645);
nor U13800 (N_13800,N_13567,N_13728);
nor U13801 (N_13801,N_13673,N_13739);
or U13802 (N_13802,N_13632,N_13667);
nand U13803 (N_13803,N_13618,N_13637);
nand U13804 (N_13804,N_13650,N_13633);
nor U13805 (N_13805,N_13677,N_13587);
or U13806 (N_13806,N_13552,N_13734);
xnor U13807 (N_13807,N_13600,N_13596);
xor U13808 (N_13808,N_13654,N_13629);
and U13809 (N_13809,N_13584,N_13580);
nand U13810 (N_13810,N_13670,N_13549);
or U13811 (N_13811,N_13626,N_13721);
and U13812 (N_13812,N_13605,N_13598);
xor U13813 (N_13813,N_13578,N_13501);
xnor U13814 (N_13814,N_13523,N_13507);
nand U13815 (N_13815,N_13554,N_13553);
nor U13816 (N_13816,N_13504,N_13733);
and U13817 (N_13817,N_13658,N_13698);
nand U13818 (N_13818,N_13711,N_13510);
or U13819 (N_13819,N_13705,N_13607);
and U13820 (N_13820,N_13614,N_13506);
and U13821 (N_13821,N_13631,N_13701);
and U13822 (N_13822,N_13546,N_13588);
or U13823 (N_13823,N_13724,N_13595);
nand U13824 (N_13824,N_13662,N_13669);
and U13825 (N_13825,N_13674,N_13716);
or U13826 (N_13826,N_13648,N_13660);
or U13827 (N_13827,N_13636,N_13599);
nand U13828 (N_13828,N_13566,N_13591);
xnor U13829 (N_13829,N_13517,N_13640);
or U13830 (N_13830,N_13534,N_13689);
xor U13831 (N_13831,N_13748,N_13634);
and U13832 (N_13832,N_13570,N_13635);
or U13833 (N_13833,N_13621,N_13615);
or U13834 (N_13834,N_13697,N_13531);
xor U13835 (N_13835,N_13575,N_13518);
xor U13836 (N_13836,N_13718,N_13539);
nor U13837 (N_13837,N_13743,N_13537);
nor U13838 (N_13838,N_13516,N_13688);
nor U13839 (N_13839,N_13606,N_13545);
or U13840 (N_13840,N_13653,N_13726);
nand U13841 (N_13841,N_13627,N_13503);
or U13842 (N_13842,N_13679,N_13542);
and U13843 (N_13843,N_13514,N_13742);
xnor U13844 (N_13844,N_13551,N_13502);
and U13845 (N_13845,N_13713,N_13638);
and U13846 (N_13846,N_13576,N_13602);
or U13847 (N_13847,N_13684,N_13594);
and U13848 (N_13848,N_13577,N_13555);
xnor U13849 (N_13849,N_13610,N_13585);
and U13850 (N_13850,N_13622,N_13741);
or U13851 (N_13851,N_13533,N_13550);
xnor U13852 (N_13852,N_13505,N_13659);
xnor U13853 (N_13853,N_13613,N_13604);
xnor U13854 (N_13854,N_13691,N_13655);
and U13855 (N_13855,N_13680,N_13695);
xor U13856 (N_13856,N_13536,N_13519);
or U13857 (N_13857,N_13558,N_13737);
nor U13858 (N_13858,N_13694,N_13657);
and U13859 (N_13859,N_13745,N_13620);
and U13860 (N_13860,N_13639,N_13641);
nor U13861 (N_13861,N_13664,N_13557);
or U13862 (N_13862,N_13706,N_13556);
nor U13863 (N_13863,N_13561,N_13747);
xnor U13864 (N_13864,N_13617,N_13623);
and U13865 (N_13865,N_13535,N_13630);
and U13866 (N_13866,N_13508,N_13547);
nor U13867 (N_13867,N_13696,N_13681);
xnor U13868 (N_13868,N_13624,N_13538);
and U13869 (N_13869,N_13628,N_13700);
nor U13870 (N_13870,N_13644,N_13643);
or U13871 (N_13871,N_13656,N_13647);
nor U13872 (N_13872,N_13601,N_13619);
xnor U13873 (N_13873,N_13642,N_13746);
nand U13874 (N_13874,N_13744,N_13723);
and U13875 (N_13875,N_13521,N_13746);
or U13876 (N_13876,N_13624,N_13601);
xnor U13877 (N_13877,N_13731,N_13670);
or U13878 (N_13878,N_13562,N_13733);
or U13879 (N_13879,N_13729,N_13606);
xor U13880 (N_13880,N_13585,N_13677);
and U13881 (N_13881,N_13609,N_13724);
nor U13882 (N_13882,N_13550,N_13553);
and U13883 (N_13883,N_13573,N_13714);
xnor U13884 (N_13884,N_13649,N_13597);
nor U13885 (N_13885,N_13732,N_13741);
xnor U13886 (N_13886,N_13736,N_13630);
or U13887 (N_13887,N_13511,N_13651);
nor U13888 (N_13888,N_13551,N_13664);
and U13889 (N_13889,N_13615,N_13557);
nand U13890 (N_13890,N_13618,N_13548);
and U13891 (N_13891,N_13724,N_13678);
xor U13892 (N_13892,N_13566,N_13745);
xnor U13893 (N_13893,N_13573,N_13657);
xnor U13894 (N_13894,N_13688,N_13600);
xnor U13895 (N_13895,N_13686,N_13705);
nor U13896 (N_13896,N_13509,N_13630);
nand U13897 (N_13897,N_13695,N_13674);
nand U13898 (N_13898,N_13712,N_13622);
nand U13899 (N_13899,N_13638,N_13704);
or U13900 (N_13900,N_13679,N_13686);
and U13901 (N_13901,N_13721,N_13656);
nor U13902 (N_13902,N_13569,N_13721);
nand U13903 (N_13903,N_13748,N_13681);
or U13904 (N_13904,N_13656,N_13603);
nor U13905 (N_13905,N_13670,N_13711);
and U13906 (N_13906,N_13554,N_13673);
nor U13907 (N_13907,N_13660,N_13720);
or U13908 (N_13908,N_13539,N_13515);
nor U13909 (N_13909,N_13505,N_13708);
and U13910 (N_13910,N_13561,N_13630);
or U13911 (N_13911,N_13559,N_13575);
or U13912 (N_13912,N_13649,N_13637);
or U13913 (N_13913,N_13697,N_13661);
and U13914 (N_13914,N_13575,N_13558);
xor U13915 (N_13915,N_13624,N_13530);
xor U13916 (N_13916,N_13586,N_13643);
nand U13917 (N_13917,N_13585,N_13605);
xnor U13918 (N_13918,N_13721,N_13579);
nand U13919 (N_13919,N_13652,N_13723);
nand U13920 (N_13920,N_13644,N_13552);
xor U13921 (N_13921,N_13673,N_13626);
or U13922 (N_13922,N_13545,N_13674);
and U13923 (N_13923,N_13573,N_13623);
xnor U13924 (N_13924,N_13559,N_13527);
and U13925 (N_13925,N_13647,N_13609);
nor U13926 (N_13926,N_13549,N_13567);
xnor U13927 (N_13927,N_13746,N_13713);
and U13928 (N_13928,N_13668,N_13703);
nor U13929 (N_13929,N_13532,N_13743);
xnor U13930 (N_13930,N_13547,N_13698);
or U13931 (N_13931,N_13538,N_13736);
and U13932 (N_13932,N_13613,N_13550);
xnor U13933 (N_13933,N_13695,N_13702);
and U13934 (N_13934,N_13655,N_13628);
nand U13935 (N_13935,N_13571,N_13741);
and U13936 (N_13936,N_13621,N_13561);
or U13937 (N_13937,N_13666,N_13627);
and U13938 (N_13938,N_13521,N_13588);
and U13939 (N_13939,N_13561,N_13717);
and U13940 (N_13940,N_13542,N_13539);
and U13941 (N_13941,N_13647,N_13700);
and U13942 (N_13942,N_13565,N_13660);
or U13943 (N_13943,N_13523,N_13686);
nor U13944 (N_13944,N_13668,N_13558);
or U13945 (N_13945,N_13666,N_13745);
and U13946 (N_13946,N_13596,N_13558);
nor U13947 (N_13947,N_13563,N_13533);
and U13948 (N_13948,N_13522,N_13595);
or U13949 (N_13949,N_13641,N_13678);
xnor U13950 (N_13950,N_13740,N_13593);
and U13951 (N_13951,N_13603,N_13581);
xnor U13952 (N_13952,N_13740,N_13555);
nand U13953 (N_13953,N_13746,N_13531);
or U13954 (N_13954,N_13530,N_13699);
xor U13955 (N_13955,N_13711,N_13557);
or U13956 (N_13956,N_13610,N_13594);
xnor U13957 (N_13957,N_13629,N_13592);
and U13958 (N_13958,N_13685,N_13633);
xor U13959 (N_13959,N_13580,N_13686);
and U13960 (N_13960,N_13601,N_13541);
and U13961 (N_13961,N_13551,N_13705);
nand U13962 (N_13962,N_13570,N_13543);
nor U13963 (N_13963,N_13592,N_13528);
nand U13964 (N_13964,N_13525,N_13662);
or U13965 (N_13965,N_13675,N_13501);
nand U13966 (N_13966,N_13658,N_13541);
nand U13967 (N_13967,N_13556,N_13547);
nand U13968 (N_13968,N_13566,N_13652);
xor U13969 (N_13969,N_13535,N_13672);
xor U13970 (N_13970,N_13667,N_13623);
nor U13971 (N_13971,N_13559,N_13610);
nor U13972 (N_13972,N_13647,N_13622);
xnor U13973 (N_13973,N_13670,N_13541);
nand U13974 (N_13974,N_13627,N_13590);
xnor U13975 (N_13975,N_13632,N_13525);
nor U13976 (N_13976,N_13684,N_13734);
xnor U13977 (N_13977,N_13630,N_13546);
nor U13978 (N_13978,N_13610,N_13526);
or U13979 (N_13979,N_13706,N_13514);
or U13980 (N_13980,N_13713,N_13628);
nand U13981 (N_13981,N_13655,N_13738);
or U13982 (N_13982,N_13651,N_13524);
nor U13983 (N_13983,N_13702,N_13661);
or U13984 (N_13984,N_13651,N_13687);
and U13985 (N_13985,N_13501,N_13632);
nor U13986 (N_13986,N_13703,N_13560);
or U13987 (N_13987,N_13573,N_13642);
nor U13988 (N_13988,N_13580,N_13510);
and U13989 (N_13989,N_13682,N_13732);
nor U13990 (N_13990,N_13668,N_13553);
nor U13991 (N_13991,N_13634,N_13525);
nand U13992 (N_13992,N_13531,N_13727);
nand U13993 (N_13993,N_13532,N_13597);
or U13994 (N_13994,N_13741,N_13686);
and U13995 (N_13995,N_13641,N_13545);
nand U13996 (N_13996,N_13572,N_13614);
or U13997 (N_13997,N_13740,N_13634);
nand U13998 (N_13998,N_13746,N_13648);
and U13999 (N_13999,N_13658,N_13537);
xnor U14000 (N_14000,N_13998,N_13822);
and U14001 (N_14001,N_13781,N_13755);
nand U14002 (N_14002,N_13901,N_13884);
xnor U14003 (N_14003,N_13805,N_13871);
nor U14004 (N_14004,N_13962,N_13970);
or U14005 (N_14005,N_13761,N_13810);
xnor U14006 (N_14006,N_13931,N_13846);
and U14007 (N_14007,N_13937,N_13869);
nand U14008 (N_14008,N_13857,N_13953);
nand U14009 (N_14009,N_13992,N_13995);
and U14010 (N_14010,N_13835,N_13927);
and U14011 (N_14011,N_13957,N_13950);
and U14012 (N_14012,N_13837,N_13788);
and U14013 (N_14013,N_13851,N_13896);
and U14014 (N_14014,N_13772,N_13844);
and U14015 (N_14015,N_13819,N_13787);
and U14016 (N_14016,N_13887,N_13866);
nand U14017 (N_14017,N_13838,N_13754);
and U14018 (N_14018,N_13867,N_13806);
or U14019 (N_14019,N_13941,N_13989);
nand U14020 (N_14020,N_13952,N_13840);
xor U14021 (N_14021,N_13983,N_13796);
or U14022 (N_14022,N_13834,N_13906);
nor U14023 (N_14023,N_13809,N_13881);
xor U14024 (N_14024,N_13969,N_13874);
or U14025 (N_14025,N_13888,N_13766);
nand U14026 (N_14026,N_13774,N_13780);
nand U14027 (N_14027,N_13948,N_13795);
or U14028 (N_14028,N_13939,N_13807);
nand U14029 (N_14029,N_13966,N_13875);
or U14030 (N_14030,N_13764,N_13895);
and U14031 (N_14031,N_13849,N_13843);
nor U14032 (N_14032,N_13975,N_13827);
and U14033 (N_14033,N_13990,N_13828);
nor U14034 (N_14034,N_13885,N_13980);
xnor U14035 (N_14035,N_13758,N_13911);
xor U14036 (N_14036,N_13776,N_13815);
and U14037 (N_14037,N_13945,N_13845);
and U14038 (N_14038,N_13899,N_13856);
and U14039 (N_14039,N_13812,N_13824);
nor U14040 (N_14040,N_13913,N_13797);
xnor U14041 (N_14041,N_13942,N_13930);
nor U14042 (N_14042,N_13790,N_13935);
nand U14043 (N_14043,N_13979,N_13928);
or U14044 (N_14044,N_13907,N_13829);
and U14045 (N_14045,N_13929,N_13919);
nor U14046 (N_14046,N_13977,N_13798);
and U14047 (N_14047,N_13753,N_13870);
nor U14048 (N_14048,N_13802,N_13876);
xnor U14049 (N_14049,N_13916,N_13804);
or U14050 (N_14050,N_13816,N_13771);
or U14051 (N_14051,N_13750,N_13852);
nand U14052 (N_14052,N_13792,N_13830);
and U14053 (N_14053,N_13985,N_13842);
xnor U14054 (N_14054,N_13892,N_13920);
and U14055 (N_14055,N_13861,N_13826);
or U14056 (N_14056,N_13974,N_13756);
nand U14057 (N_14057,N_13760,N_13784);
or U14058 (N_14058,N_13823,N_13894);
or U14059 (N_14059,N_13877,N_13794);
nand U14060 (N_14060,N_13978,N_13793);
nand U14061 (N_14061,N_13914,N_13959);
nor U14062 (N_14062,N_13799,N_13994);
xnor U14063 (N_14063,N_13751,N_13864);
and U14064 (N_14064,N_13841,N_13768);
xor U14065 (N_14065,N_13904,N_13882);
or U14066 (N_14066,N_13891,N_13854);
and U14067 (N_14067,N_13860,N_13820);
xnor U14068 (N_14068,N_13893,N_13847);
and U14069 (N_14069,N_13997,N_13988);
and U14070 (N_14070,N_13900,N_13924);
nor U14071 (N_14071,N_13909,N_13991);
and U14072 (N_14072,N_13859,N_13968);
and U14073 (N_14073,N_13855,N_13897);
nand U14074 (N_14074,N_13903,N_13850);
xnor U14075 (N_14075,N_13918,N_13915);
and U14076 (N_14076,N_13831,N_13848);
and U14077 (N_14077,N_13825,N_13936);
nand U14078 (N_14078,N_13814,N_13883);
xor U14079 (N_14079,N_13955,N_13946);
and U14080 (N_14080,N_13811,N_13785);
nand U14081 (N_14081,N_13808,N_13905);
and U14082 (N_14082,N_13961,N_13986);
xor U14083 (N_14083,N_13757,N_13763);
xor U14084 (N_14084,N_13973,N_13908);
nand U14085 (N_14085,N_13886,N_13777);
nand U14086 (N_14086,N_13917,N_13984);
xnor U14087 (N_14087,N_13933,N_13912);
nor U14088 (N_14088,N_13836,N_13821);
nand U14089 (N_14089,N_13921,N_13954);
and U14090 (N_14090,N_13898,N_13947);
and U14091 (N_14091,N_13976,N_13902);
nor U14092 (N_14092,N_13938,N_13981);
nor U14093 (N_14093,N_13934,N_13865);
nand U14094 (N_14094,N_13863,N_13789);
and U14095 (N_14095,N_13803,N_13775);
xor U14096 (N_14096,N_13996,N_13993);
nor U14097 (N_14097,N_13832,N_13925);
or U14098 (N_14098,N_13926,N_13786);
nand U14099 (N_14099,N_13778,N_13767);
nor U14100 (N_14100,N_13765,N_13999);
nor U14101 (N_14101,N_13872,N_13862);
nand U14102 (N_14102,N_13972,N_13773);
xnor U14103 (N_14103,N_13967,N_13982);
nand U14104 (N_14104,N_13880,N_13960);
nor U14105 (N_14105,N_13868,N_13759);
or U14106 (N_14106,N_13833,N_13964);
or U14107 (N_14107,N_13940,N_13951);
or U14108 (N_14108,N_13963,N_13958);
xnor U14109 (N_14109,N_13987,N_13879);
xnor U14110 (N_14110,N_13890,N_13752);
or U14111 (N_14111,N_13858,N_13922);
nor U14112 (N_14112,N_13853,N_13932);
or U14113 (N_14113,N_13944,N_13965);
or U14114 (N_14114,N_13801,N_13791);
and U14115 (N_14115,N_13762,N_13873);
xnor U14116 (N_14116,N_13783,N_13769);
nor U14117 (N_14117,N_13782,N_13923);
nand U14118 (N_14118,N_13949,N_13817);
xor U14119 (N_14119,N_13943,N_13770);
xor U14120 (N_14120,N_13818,N_13971);
nor U14121 (N_14121,N_13800,N_13910);
nor U14122 (N_14122,N_13839,N_13956);
and U14123 (N_14123,N_13779,N_13813);
nor U14124 (N_14124,N_13878,N_13889);
and U14125 (N_14125,N_13889,N_13994);
xnor U14126 (N_14126,N_13869,N_13764);
or U14127 (N_14127,N_13889,N_13873);
and U14128 (N_14128,N_13823,N_13918);
xnor U14129 (N_14129,N_13856,N_13763);
xnor U14130 (N_14130,N_13924,N_13865);
and U14131 (N_14131,N_13960,N_13918);
or U14132 (N_14132,N_13792,N_13850);
or U14133 (N_14133,N_13861,N_13846);
nand U14134 (N_14134,N_13973,N_13775);
and U14135 (N_14135,N_13995,N_13808);
nor U14136 (N_14136,N_13902,N_13838);
xnor U14137 (N_14137,N_13998,N_13897);
xor U14138 (N_14138,N_13868,N_13879);
xnor U14139 (N_14139,N_13828,N_13897);
nand U14140 (N_14140,N_13785,N_13987);
xor U14141 (N_14141,N_13910,N_13849);
nand U14142 (N_14142,N_13924,N_13810);
nor U14143 (N_14143,N_13770,N_13773);
xor U14144 (N_14144,N_13928,N_13974);
xor U14145 (N_14145,N_13798,N_13926);
xor U14146 (N_14146,N_13951,N_13986);
nor U14147 (N_14147,N_13985,N_13955);
nor U14148 (N_14148,N_13879,N_13859);
nor U14149 (N_14149,N_13803,N_13924);
nor U14150 (N_14150,N_13897,N_13764);
or U14151 (N_14151,N_13783,N_13976);
xor U14152 (N_14152,N_13765,N_13963);
nor U14153 (N_14153,N_13811,N_13777);
or U14154 (N_14154,N_13954,N_13926);
or U14155 (N_14155,N_13932,N_13860);
and U14156 (N_14156,N_13765,N_13870);
and U14157 (N_14157,N_13763,N_13878);
nor U14158 (N_14158,N_13980,N_13789);
xnor U14159 (N_14159,N_13847,N_13855);
and U14160 (N_14160,N_13866,N_13935);
or U14161 (N_14161,N_13769,N_13971);
or U14162 (N_14162,N_13863,N_13784);
nor U14163 (N_14163,N_13831,N_13853);
xnor U14164 (N_14164,N_13974,N_13800);
nand U14165 (N_14165,N_13968,N_13954);
or U14166 (N_14166,N_13829,N_13752);
or U14167 (N_14167,N_13859,N_13878);
nand U14168 (N_14168,N_13841,N_13968);
or U14169 (N_14169,N_13999,N_13854);
and U14170 (N_14170,N_13894,N_13965);
nand U14171 (N_14171,N_13963,N_13858);
xor U14172 (N_14172,N_13879,N_13889);
nand U14173 (N_14173,N_13760,N_13851);
xnor U14174 (N_14174,N_13939,N_13814);
nor U14175 (N_14175,N_13923,N_13999);
nor U14176 (N_14176,N_13825,N_13918);
nand U14177 (N_14177,N_13787,N_13891);
nand U14178 (N_14178,N_13755,N_13964);
and U14179 (N_14179,N_13956,N_13827);
or U14180 (N_14180,N_13843,N_13895);
nor U14181 (N_14181,N_13785,N_13831);
and U14182 (N_14182,N_13960,N_13869);
xor U14183 (N_14183,N_13991,N_13821);
xor U14184 (N_14184,N_13859,N_13987);
and U14185 (N_14185,N_13899,N_13852);
and U14186 (N_14186,N_13794,N_13951);
xor U14187 (N_14187,N_13997,N_13984);
or U14188 (N_14188,N_13990,N_13989);
nor U14189 (N_14189,N_13934,N_13926);
xor U14190 (N_14190,N_13774,N_13827);
xor U14191 (N_14191,N_13948,N_13857);
xor U14192 (N_14192,N_13834,N_13893);
or U14193 (N_14193,N_13828,N_13838);
nand U14194 (N_14194,N_13924,N_13967);
nor U14195 (N_14195,N_13906,N_13982);
nor U14196 (N_14196,N_13847,N_13829);
xor U14197 (N_14197,N_13913,N_13941);
or U14198 (N_14198,N_13752,N_13827);
or U14199 (N_14199,N_13901,N_13949);
nor U14200 (N_14200,N_13859,N_13991);
nand U14201 (N_14201,N_13846,N_13893);
or U14202 (N_14202,N_13942,N_13967);
or U14203 (N_14203,N_13837,N_13758);
xnor U14204 (N_14204,N_13964,N_13888);
nand U14205 (N_14205,N_13950,N_13780);
and U14206 (N_14206,N_13846,N_13969);
nor U14207 (N_14207,N_13798,N_13888);
xnor U14208 (N_14208,N_13888,N_13852);
nand U14209 (N_14209,N_13841,N_13933);
nand U14210 (N_14210,N_13975,N_13823);
nor U14211 (N_14211,N_13946,N_13774);
and U14212 (N_14212,N_13885,N_13843);
nor U14213 (N_14213,N_13931,N_13873);
or U14214 (N_14214,N_13983,N_13995);
and U14215 (N_14215,N_13802,N_13996);
xnor U14216 (N_14216,N_13945,N_13967);
or U14217 (N_14217,N_13808,N_13853);
nand U14218 (N_14218,N_13873,N_13756);
xnor U14219 (N_14219,N_13960,N_13851);
nor U14220 (N_14220,N_13853,N_13787);
nor U14221 (N_14221,N_13886,N_13882);
nand U14222 (N_14222,N_13929,N_13772);
nand U14223 (N_14223,N_13979,N_13777);
or U14224 (N_14224,N_13930,N_13778);
nor U14225 (N_14225,N_13962,N_13802);
nor U14226 (N_14226,N_13937,N_13838);
nor U14227 (N_14227,N_13825,N_13874);
nand U14228 (N_14228,N_13890,N_13783);
nand U14229 (N_14229,N_13919,N_13853);
nor U14230 (N_14230,N_13919,N_13822);
nor U14231 (N_14231,N_13797,N_13832);
or U14232 (N_14232,N_13993,N_13941);
nor U14233 (N_14233,N_13883,N_13767);
nand U14234 (N_14234,N_13962,N_13912);
and U14235 (N_14235,N_13772,N_13763);
nand U14236 (N_14236,N_13873,N_13890);
or U14237 (N_14237,N_13774,N_13872);
and U14238 (N_14238,N_13930,N_13914);
nand U14239 (N_14239,N_13765,N_13780);
or U14240 (N_14240,N_13917,N_13931);
or U14241 (N_14241,N_13849,N_13832);
nand U14242 (N_14242,N_13845,N_13834);
nand U14243 (N_14243,N_13756,N_13768);
xnor U14244 (N_14244,N_13923,N_13815);
xor U14245 (N_14245,N_13931,N_13912);
or U14246 (N_14246,N_13789,N_13920);
nand U14247 (N_14247,N_13813,N_13997);
nor U14248 (N_14248,N_13952,N_13786);
xnor U14249 (N_14249,N_13761,N_13857);
or U14250 (N_14250,N_14237,N_14127);
and U14251 (N_14251,N_14036,N_14118);
or U14252 (N_14252,N_14082,N_14229);
and U14253 (N_14253,N_14193,N_14031);
nand U14254 (N_14254,N_14246,N_14125);
xnor U14255 (N_14255,N_14037,N_14012);
nor U14256 (N_14256,N_14241,N_14227);
and U14257 (N_14257,N_14184,N_14014);
nand U14258 (N_14258,N_14016,N_14130);
nor U14259 (N_14259,N_14232,N_14168);
xor U14260 (N_14260,N_14033,N_14039);
xnor U14261 (N_14261,N_14211,N_14077);
or U14262 (N_14262,N_14226,N_14142);
nor U14263 (N_14263,N_14165,N_14126);
xnor U14264 (N_14264,N_14078,N_14170);
nor U14265 (N_14265,N_14138,N_14162);
nand U14266 (N_14266,N_14054,N_14045);
nand U14267 (N_14267,N_14236,N_14104);
nor U14268 (N_14268,N_14102,N_14148);
and U14269 (N_14269,N_14063,N_14018);
nand U14270 (N_14270,N_14121,N_14160);
xor U14271 (N_14271,N_14084,N_14005);
nor U14272 (N_14272,N_14188,N_14136);
or U14273 (N_14273,N_14020,N_14052);
and U14274 (N_14274,N_14115,N_14047);
nor U14275 (N_14275,N_14083,N_14153);
xor U14276 (N_14276,N_14097,N_14240);
and U14277 (N_14277,N_14145,N_14096);
or U14278 (N_14278,N_14141,N_14124);
nor U14279 (N_14279,N_14057,N_14200);
or U14280 (N_14280,N_14003,N_14175);
nand U14281 (N_14281,N_14166,N_14189);
or U14282 (N_14282,N_14080,N_14172);
xor U14283 (N_14283,N_14212,N_14247);
nand U14284 (N_14284,N_14181,N_14085);
xor U14285 (N_14285,N_14008,N_14041);
xnor U14286 (N_14286,N_14025,N_14056);
nor U14287 (N_14287,N_14233,N_14049);
nor U14288 (N_14288,N_14196,N_14028);
or U14289 (N_14289,N_14143,N_14167);
nand U14290 (N_14290,N_14004,N_14040);
and U14291 (N_14291,N_14109,N_14244);
and U14292 (N_14292,N_14207,N_14019);
and U14293 (N_14293,N_14069,N_14242);
and U14294 (N_14294,N_14191,N_14195);
nor U14295 (N_14295,N_14027,N_14216);
xor U14296 (N_14296,N_14000,N_14190);
and U14297 (N_14297,N_14058,N_14133);
and U14298 (N_14298,N_14098,N_14199);
or U14299 (N_14299,N_14068,N_14208);
nor U14300 (N_14300,N_14197,N_14100);
or U14301 (N_14301,N_14156,N_14220);
nor U14302 (N_14302,N_14013,N_14228);
nor U14303 (N_14303,N_14214,N_14095);
xnor U14304 (N_14304,N_14128,N_14223);
nand U14305 (N_14305,N_14131,N_14092);
nand U14306 (N_14306,N_14137,N_14174);
or U14307 (N_14307,N_14001,N_14169);
nor U14308 (N_14308,N_14091,N_14202);
nand U14309 (N_14309,N_14177,N_14009);
or U14310 (N_14310,N_14029,N_14094);
and U14311 (N_14311,N_14178,N_14221);
xnor U14312 (N_14312,N_14132,N_14024);
nand U14313 (N_14313,N_14122,N_14144);
or U14314 (N_14314,N_14210,N_14180);
nor U14315 (N_14315,N_14134,N_14140);
and U14316 (N_14316,N_14204,N_14061);
and U14317 (N_14317,N_14203,N_14176);
xor U14318 (N_14318,N_14044,N_14042);
nand U14319 (N_14319,N_14217,N_14030);
nand U14320 (N_14320,N_14116,N_14113);
and U14321 (N_14321,N_14230,N_14087);
nand U14322 (N_14322,N_14002,N_14157);
xnor U14323 (N_14323,N_14205,N_14225);
nor U14324 (N_14324,N_14108,N_14067);
and U14325 (N_14325,N_14158,N_14201);
nor U14326 (N_14326,N_14119,N_14219);
nor U14327 (N_14327,N_14163,N_14192);
and U14328 (N_14328,N_14171,N_14007);
nor U14329 (N_14329,N_14173,N_14011);
xor U14330 (N_14330,N_14086,N_14146);
and U14331 (N_14331,N_14046,N_14218);
nor U14332 (N_14332,N_14187,N_14070);
nor U14333 (N_14333,N_14238,N_14035);
nor U14334 (N_14334,N_14053,N_14198);
and U14335 (N_14335,N_14185,N_14164);
xor U14336 (N_14336,N_14129,N_14151);
and U14337 (N_14337,N_14159,N_14038);
xnor U14338 (N_14338,N_14183,N_14234);
xnor U14339 (N_14339,N_14074,N_14114);
xor U14340 (N_14340,N_14017,N_14065);
and U14341 (N_14341,N_14186,N_14235);
nor U14342 (N_14342,N_14182,N_14006);
and U14343 (N_14343,N_14051,N_14071);
and U14344 (N_14344,N_14064,N_14110);
nor U14345 (N_14345,N_14248,N_14072);
xor U14346 (N_14346,N_14215,N_14015);
and U14347 (N_14347,N_14161,N_14079);
and U14348 (N_14348,N_14123,N_14093);
and U14349 (N_14349,N_14105,N_14066);
xnor U14350 (N_14350,N_14152,N_14103);
nor U14351 (N_14351,N_14073,N_14107);
and U14352 (N_14352,N_14101,N_14075);
or U14353 (N_14353,N_14023,N_14088);
xnor U14354 (N_14354,N_14010,N_14090);
and U14355 (N_14355,N_14194,N_14055);
nand U14356 (N_14356,N_14048,N_14213);
nor U14357 (N_14357,N_14249,N_14076);
and U14358 (N_14358,N_14022,N_14050);
xor U14359 (N_14359,N_14139,N_14099);
and U14360 (N_14360,N_14209,N_14021);
xor U14361 (N_14361,N_14149,N_14060);
or U14362 (N_14362,N_14026,N_14117);
nand U14363 (N_14363,N_14147,N_14179);
and U14364 (N_14364,N_14120,N_14206);
or U14365 (N_14365,N_14032,N_14222);
nor U14366 (N_14366,N_14111,N_14150);
xor U14367 (N_14367,N_14043,N_14239);
xor U14368 (N_14368,N_14059,N_14155);
xor U14369 (N_14369,N_14062,N_14224);
or U14370 (N_14370,N_14135,N_14112);
or U14371 (N_14371,N_14081,N_14231);
and U14372 (N_14372,N_14089,N_14245);
nor U14373 (N_14373,N_14034,N_14243);
nand U14374 (N_14374,N_14106,N_14154);
nand U14375 (N_14375,N_14067,N_14135);
or U14376 (N_14376,N_14046,N_14123);
nand U14377 (N_14377,N_14071,N_14133);
nand U14378 (N_14378,N_14050,N_14072);
and U14379 (N_14379,N_14080,N_14233);
or U14380 (N_14380,N_14181,N_14067);
and U14381 (N_14381,N_14149,N_14225);
nand U14382 (N_14382,N_14091,N_14089);
or U14383 (N_14383,N_14087,N_14202);
nand U14384 (N_14384,N_14115,N_14124);
or U14385 (N_14385,N_14075,N_14144);
xnor U14386 (N_14386,N_14110,N_14186);
and U14387 (N_14387,N_14184,N_14095);
or U14388 (N_14388,N_14049,N_14086);
nor U14389 (N_14389,N_14245,N_14247);
or U14390 (N_14390,N_14192,N_14131);
nand U14391 (N_14391,N_14239,N_14154);
xnor U14392 (N_14392,N_14204,N_14080);
or U14393 (N_14393,N_14137,N_14163);
xnor U14394 (N_14394,N_14208,N_14193);
xor U14395 (N_14395,N_14007,N_14239);
or U14396 (N_14396,N_14211,N_14008);
or U14397 (N_14397,N_14101,N_14225);
nor U14398 (N_14398,N_14162,N_14043);
or U14399 (N_14399,N_14161,N_14040);
xor U14400 (N_14400,N_14180,N_14033);
nor U14401 (N_14401,N_14148,N_14022);
xor U14402 (N_14402,N_14209,N_14102);
xor U14403 (N_14403,N_14172,N_14089);
or U14404 (N_14404,N_14111,N_14195);
and U14405 (N_14405,N_14155,N_14192);
xnor U14406 (N_14406,N_14185,N_14129);
nor U14407 (N_14407,N_14140,N_14052);
nor U14408 (N_14408,N_14024,N_14214);
xor U14409 (N_14409,N_14147,N_14056);
nor U14410 (N_14410,N_14120,N_14236);
and U14411 (N_14411,N_14224,N_14246);
xor U14412 (N_14412,N_14000,N_14010);
or U14413 (N_14413,N_14062,N_14163);
and U14414 (N_14414,N_14023,N_14066);
nor U14415 (N_14415,N_14053,N_14246);
nor U14416 (N_14416,N_14081,N_14002);
xor U14417 (N_14417,N_14038,N_14085);
nand U14418 (N_14418,N_14108,N_14178);
and U14419 (N_14419,N_14164,N_14220);
or U14420 (N_14420,N_14047,N_14135);
xor U14421 (N_14421,N_14191,N_14219);
xor U14422 (N_14422,N_14052,N_14132);
or U14423 (N_14423,N_14107,N_14212);
or U14424 (N_14424,N_14188,N_14114);
xor U14425 (N_14425,N_14115,N_14133);
or U14426 (N_14426,N_14164,N_14086);
and U14427 (N_14427,N_14125,N_14175);
nor U14428 (N_14428,N_14189,N_14177);
nor U14429 (N_14429,N_14126,N_14149);
or U14430 (N_14430,N_14149,N_14143);
xnor U14431 (N_14431,N_14202,N_14088);
xor U14432 (N_14432,N_14146,N_14142);
and U14433 (N_14433,N_14171,N_14193);
and U14434 (N_14434,N_14218,N_14050);
xnor U14435 (N_14435,N_14099,N_14044);
nand U14436 (N_14436,N_14207,N_14150);
and U14437 (N_14437,N_14014,N_14144);
or U14438 (N_14438,N_14021,N_14235);
or U14439 (N_14439,N_14175,N_14037);
and U14440 (N_14440,N_14057,N_14125);
nand U14441 (N_14441,N_14181,N_14071);
and U14442 (N_14442,N_14076,N_14243);
and U14443 (N_14443,N_14063,N_14107);
nor U14444 (N_14444,N_14134,N_14080);
xor U14445 (N_14445,N_14141,N_14233);
and U14446 (N_14446,N_14167,N_14189);
xnor U14447 (N_14447,N_14038,N_14032);
xnor U14448 (N_14448,N_14152,N_14062);
nand U14449 (N_14449,N_14224,N_14152);
and U14450 (N_14450,N_14088,N_14135);
nor U14451 (N_14451,N_14036,N_14038);
nor U14452 (N_14452,N_14234,N_14223);
and U14453 (N_14453,N_14137,N_14108);
nand U14454 (N_14454,N_14073,N_14230);
nand U14455 (N_14455,N_14213,N_14210);
nor U14456 (N_14456,N_14035,N_14246);
xor U14457 (N_14457,N_14000,N_14197);
and U14458 (N_14458,N_14112,N_14115);
or U14459 (N_14459,N_14172,N_14012);
nand U14460 (N_14460,N_14077,N_14080);
nand U14461 (N_14461,N_14213,N_14052);
and U14462 (N_14462,N_14217,N_14067);
xor U14463 (N_14463,N_14072,N_14101);
nand U14464 (N_14464,N_14219,N_14062);
and U14465 (N_14465,N_14247,N_14092);
nor U14466 (N_14466,N_14129,N_14220);
nand U14467 (N_14467,N_14240,N_14037);
nand U14468 (N_14468,N_14142,N_14194);
xnor U14469 (N_14469,N_14242,N_14001);
or U14470 (N_14470,N_14019,N_14008);
and U14471 (N_14471,N_14151,N_14207);
nand U14472 (N_14472,N_14225,N_14056);
nand U14473 (N_14473,N_14194,N_14211);
nand U14474 (N_14474,N_14164,N_14189);
nor U14475 (N_14475,N_14066,N_14100);
nor U14476 (N_14476,N_14097,N_14058);
xor U14477 (N_14477,N_14096,N_14238);
or U14478 (N_14478,N_14081,N_14166);
or U14479 (N_14479,N_14117,N_14231);
nor U14480 (N_14480,N_14040,N_14169);
and U14481 (N_14481,N_14214,N_14035);
xnor U14482 (N_14482,N_14189,N_14147);
or U14483 (N_14483,N_14085,N_14156);
and U14484 (N_14484,N_14000,N_14218);
or U14485 (N_14485,N_14179,N_14025);
xnor U14486 (N_14486,N_14186,N_14032);
xor U14487 (N_14487,N_14036,N_14140);
xor U14488 (N_14488,N_14225,N_14067);
or U14489 (N_14489,N_14177,N_14151);
nand U14490 (N_14490,N_14121,N_14126);
nand U14491 (N_14491,N_14219,N_14004);
xnor U14492 (N_14492,N_14175,N_14050);
nand U14493 (N_14493,N_14226,N_14000);
nor U14494 (N_14494,N_14147,N_14021);
or U14495 (N_14495,N_14040,N_14248);
and U14496 (N_14496,N_14067,N_14229);
nor U14497 (N_14497,N_14087,N_14219);
nand U14498 (N_14498,N_14118,N_14024);
nand U14499 (N_14499,N_14113,N_14096);
nor U14500 (N_14500,N_14314,N_14396);
xnor U14501 (N_14501,N_14413,N_14408);
nor U14502 (N_14502,N_14387,N_14497);
nand U14503 (N_14503,N_14337,N_14435);
or U14504 (N_14504,N_14361,N_14395);
nand U14505 (N_14505,N_14482,N_14400);
or U14506 (N_14506,N_14464,N_14283);
and U14507 (N_14507,N_14309,N_14367);
xnor U14508 (N_14508,N_14407,N_14363);
or U14509 (N_14509,N_14439,N_14455);
and U14510 (N_14510,N_14307,N_14305);
xor U14511 (N_14511,N_14419,N_14404);
or U14512 (N_14512,N_14493,N_14294);
xnor U14513 (N_14513,N_14284,N_14452);
nor U14514 (N_14514,N_14274,N_14290);
nand U14515 (N_14515,N_14374,N_14441);
or U14516 (N_14516,N_14425,N_14470);
nand U14517 (N_14517,N_14299,N_14368);
xor U14518 (N_14518,N_14357,N_14479);
or U14519 (N_14519,N_14401,N_14383);
or U14520 (N_14520,N_14466,N_14465);
nor U14521 (N_14521,N_14446,N_14444);
and U14522 (N_14522,N_14477,N_14471);
nor U14523 (N_14523,N_14454,N_14457);
nand U14524 (N_14524,N_14376,N_14463);
or U14525 (N_14525,N_14293,N_14494);
and U14526 (N_14526,N_14336,N_14285);
nand U14527 (N_14527,N_14366,N_14453);
nand U14528 (N_14528,N_14297,N_14442);
xnor U14529 (N_14529,N_14420,N_14349);
nand U14530 (N_14530,N_14438,N_14409);
and U14531 (N_14531,N_14476,N_14369);
nor U14532 (N_14532,N_14449,N_14310);
nor U14533 (N_14533,N_14430,N_14346);
and U14534 (N_14534,N_14286,N_14263);
and U14535 (N_14535,N_14300,N_14418);
and U14536 (N_14536,N_14484,N_14333);
nand U14537 (N_14537,N_14252,N_14478);
or U14538 (N_14538,N_14377,N_14498);
nand U14539 (N_14539,N_14354,N_14436);
nor U14540 (N_14540,N_14386,N_14417);
nor U14541 (N_14541,N_14358,N_14338);
and U14542 (N_14542,N_14474,N_14277);
and U14543 (N_14543,N_14316,N_14332);
or U14544 (N_14544,N_14375,N_14469);
or U14545 (N_14545,N_14372,N_14384);
and U14546 (N_14546,N_14485,N_14467);
and U14547 (N_14547,N_14313,N_14301);
nor U14548 (N_14548,N_14398,N_14259);
xnor U14549 (N_14549,N_14412,N_14276);
xnor U14550 (N_14550,N_14262,N_14495);
nor U14551 (N_14551,N_14379,N_14257);
nand U14552 (N_14552,N_14350,N_14339);
and U14553 (N_14553,N_14326,N_14391);
nor U14554 (N_14554,N_14403,N_14272);
nand U14555 (N_14555,N_14320,N_14415);
or U14556 (N_14556,N_14496,N_14296);
nor U14557 (N_14557,N_14311,N_14424);
and U14558 (N_14558,N_14260,N_14289);
nor U14559 (N_14559,N_14322,N_14399);
and U14560 (N_14560,N_14472,N_14380);
and U14561 (N_14561,N_14440,N_14458);
xor U14562 (N_14562,N_14448,N_14251);
or U14563 (N_14563,N_14393,N_14394);
or U14564 (N_14564,N_14483,N_14266);
nand U14565 (N_14565,N_14288,N_14388);
and U14566 (N_14566,N_14342,N_14315);
or U14567 (N_14567,N_14433,N_14373);
nor U14568 (N_14568,N_14302,N_14268);
xnor U14569 (N_14569,N_14382,N_14278);
xnor U14570 (N_14570,N_14319,N_14267);
or U14571 (N_14571,N_14328,N_14253);
nor U14572 (N_14572,N_14422,N_14261);
nand U14573 (N_14573,N_14329,N_14456);
and U14574 (N_14574,N_14352,N_14287);
xor U14575 (N_14575,N_14281,N_14371);
and U14576 (N_14576,N_14345,N_14324);
xor U14577 (N_14577,N_14450,N_14460);
nand U14578 (N_14578,N_14423,N_14256);
nor U14579 (N_14579,N_14325,N_14321);
or U14580 (N_14580,N_14347,N_14416);
xor U14581 (N_14581,N_14364,N_14429);
nor U14582 (N_14582,N_14434,N_14356);
or U14583 (N_14583,N_14254,N_14280);
nor U14584 (N_14584,N_14317,N_14392);
or U14585 (N_14585,N_14335,N_14491);
and U14586 (N_14586,N_14462,N_14327);
nand U14587 (N_14587,N_14437,N_14303);
and U14588 (N_14588,N_14406,N_14431);
xor U14589 (N_14589,N_14432,N_14397);
or U14590 (N_14590,N_14273,N_14421);
and U14591 (N_14591,N_14298,N_14308);
or U14592 (N_14592,N_14343,N_14330);
nor U14593 (N_14593,N_14473,N_14334);
nand U14594 (N_14594,N_14265,N_14370);
nor U14595 (N_14595,N_14411,N_14295);
xnor U14596 (N_14596,N_14323,N_14447);
nand U14597 (N_14597,N_14258,N_14427);
nand U14598 (N_14598,N_14255,N_14306);
and U14599 (N_14599,N_14492,N_14481);
xor U14600 (N_14600,N_14410,N_14348);
nand U14601 (N_14601,N_14385,N_14443);
nand U14602 (N_14602,N_14459,N_14291);
xnor U14603 (N_14603,N_14351,N_14362);
or U14604 (N_14604,N_14468,N_14405);
nand U14605 (N_14605,N_14487,N_14360);
or U14606 (N_14606,N_14340,N_14359);
or U14607 (N_14607,N_14426,N_14490);
or U14608 (N_14608,N_14275,N_14445);
nand U14609 (N_14609,N_14381,N_14292);
xor U14610 (N_14610,N_14499,N_14355);
or U14611 (N_14611,N_14312,N_14389);
and U14612 (N_14612,N_14378,N_14270);
or U14613 (N_14613,N_14250,N_14264);
and U14614 (N_14614,N_14344,N_14331);
nor U14615 (N_14615,N_14269,N_14451);
or U14616 (N_14616,N_14304,N_14365);
nor U14617 (N_14617,N_14480,N_14271);
and U14618 (N_14618,N_14318,N_14279);
nor U14619 (N_14619,N_14461,N_14489);
xor U14620 (N_14620,N_14428,N_14353);
or U14621 (N_14621,N_14475,N_14414);
xnor U14622 (N_14622,N_14341,N_14488);
xnor U14623 (N_14623,N_14402,N_14486);
nor U14624 (N_14624,N_14282,N_14390);
xor U14625 (N_14625,N_14329,N_14410);
nand U14626 (N_14626,N_14403,N_14301);
nor U14627 (N_14627,N_14343,N_14425);
nand U14628 (N_14628,N_14268,N_14447);
and U14629 (N_14629,N_14325,N_14300);
nand U14630 (N_14630,N_14322,N_14423);
xnor U14631 (N_14631,N_14496,N_14309);
and U14632 (N_14632,N_14479,N_14457);
nor U14633 (N_14633,N_14460,N_14393);
nor U14634 (N_14634,N_14396,N_14495);
nor U14635 (N_14635,N_14439,N_14459);
nor U14636 (N_14636,N_14452,N_14454);
nor U14637 (N_14637,N_14383,N_14400);
xnor U14638 (N_14638,N_14423,N_14461);
nor U14639 (N_14639,N_14274,N_14349);
xnor U14640 (N_14640,N_14356,N_14404);
and U14641 (N_14641,N_14299,N_14290);
nand U14642 (N_14642,N_14314,N_14261);
nand U14643 (N_14643,N_14293,N_14362);
xnor U14644 (N_14644,N_14359,N_14405);
and U14645 (N_14645,N_14494,N_14298);
nand U14646 (N_14646,N_14392,N_14484);
nand U14647 (N_14647,N_14273,N_14449);
nand U14648 (N_14648,N_14487,N_14345);
xor U14649 (N_14649,N_14303,N_14465);
and U14650 (N_14650,N_14344,N_14417);
xnor U14651 (N_14651,N_14486,N_14376);
and U14652 (N_14652,N_14429,N_14305);
or U14653 (N_14653,N_14296,N_14277);
nor U14654 (N_14654,N_14479,N_14303);
xor U14655 (N_14655,N_14451,N_14434);
and U14656 (N_14656,N_14268,N_14453);
and U14657 (N_14657,N_14359,N_14346);
nand U14658 (N_14658,N_14471,N_14343);
or U14659 (N_14659,N_14390,N_14499);
nand U14660 (N_14660,N_14478,N_14364);
xnor U14661 (N_14661,N_14316,N_14309);
xnor U14662 (N_14662,N_14376,N_14340);
xor U14663 (N_14663,N_14328,N_14371);
nor U14664 (N_14664,N_14271,N_14494);
nand U14665 (N_14665,N_14403,N_14392);
and U14666 (N_14666,N_14435,N_14277);
xor U14667 (N_14667,N_14256,N_14381);
xnor U14668 (N_14668,N_14484,N_14355);
nor U14669 (N_14669,N_14285,N_14447);
and U14670 (N_14670,N_14284,N_14456);
or U14671 (N_14671,N_14411,N_14409);
nand U14672 (N_14672,N_14288,N_14368);
xnor U14673 (N_14673,N_14402,N_14269);
xnor U14674 (N_14674,N_14440,N_14312);
nand U14675 (N_14675,N_14474,N_14258);
or U14676 (N_14676,N_14271,N_14428);
xnor U14677 (N_14677,N_14446,N_14391);
nand U14678 (N_14678,N_14493,N_14271);
or U14679 (N_14679,N_14290,N_14305);
or U14680 (N_14680,N_14320,N_14479);
or U14681 (N_14681,N_14487,N_14394);
xnor U14682 (N_14682,N_14459,N_14301);
or U14683 (N_14683,N_14369,N_14286);
nor U14684 (N_14684,N_14485,N_14306);
xor U14685 (N_14685,N_14392,N_14291);
nor U14686 (N_14686,N_14274,N_14379);
and U14687 (N_14687,N_14296,N_14369);
or U14688 (N_14688,N_14400,N_14285);
xor U14689 (N_14689,N_14311,N_14455);
and U14690 (N_14690,N_14394,N_14332);
nor U14691 (N_14691,N_14332,N_14354);
nor U14692 (N_14692,N_14267,N_14491);
and U14693 (N_14693,N_14312,N_14263);
nor U14694 (N_14694,N_14428,N_14425);
xnor U14695 (N_14695,N_14422,N_14352);
or U14696 (N_14696,N_14293,N_14468);
nand U14697 (N_14697,N_14482,N_14288);
xor U14698 (N_14698,N_14416,N_14393);
xor U14699 (N_14699,N_14269,N_14398);
xor U14700 (N_14700,N_14305,N_14356);
xnor U14701 (N_14701,N_14428,N_14340);
and U14702 (N_14702,N_14264,N_14391);
xor U14703 (N_14703,N_14380,N_14307);
nor U14704 (N_14704,N_14260,N_14415);
and U14705 (N_14705,N_14442,N_14440);
nor U14706 (N_14706,N_14260,N_14421);
nand U14707 (N_14707,N_14376,N_14455);
or U14708 (N_14708,N_14302,N_14413);
xnor U14709 (N_14709,N_14484,N_14365);
xor U14710 (N_14710,N_14397,N_14462);
xor U14711 (N_14711,N_14394,N_14409);
nor U14712 (N_14712,N_14363,N_14395);
or U14713 (N_14713,N_14442,N_14269);
nor U14714 (N_14714,N_14461,N_14409);
and U14715 (N_14715,N_14278,N_14264);
xnor U14716 (N_14716,N_14258,N_14359);
or U14717 (N_14717,N_14334,N_14268);
nor U14718 (N_14718,N_14390,N_14300);
nand U14719 (N_14719,N_14346,N_14437);
nor U14720 (N_14720,N_14435,N_14456);
and U14721 (N_14721,N_14453,N_14450);
xor U14722 (N_14722,N_14457,N_14306);
or U14723 (N_14723,N_14454,N_14496);
nor U14724 (N_14724,N_14296,N_14469);
xnor U14725 (N_14725,N_14338,N_14400);
nand U14726 (N_14726,N_14443,N_14494);
xor U14727 (N_14727,N_14276,N_14457);
nand U14728 (N_14728,N_14308,N_14313);
xor U14729 (N_14729,N_14370,N_14375);
or U14730 (N_14730,N_14415,N_14453);
or U14731 (N_14731,N_14302,N_14375);
xnor U14732 (N_14732,N_14398,N_14263);
xor U14733 (N_14733,N_14448,N_14252);
xor U14734 (N_14734,N_14463,N_14471);
nand U14735 (N_14735,N_14284,N_14280);
or U14736 (N_14736,N_14398,N_14325);
xnor U14737 (N_14737,N_14401,N_14348);
xnor U14738 (N_14738,N_14276,N_14324);
or U14739 (N_14739,N_14366,N_14384);
xnor U14740 (N_14740,N_14474,N_14412);
nor U14741 (N_14741,N_14256,N_14398);
or U14742 (N_14742,N_14442,N_14284);
or U14743 (N_14743,N_14326,N_14390);
xor U14744 (N_14744,N_14431,N_14334);
xnor U14745 (N_14745,N_14376,N_14353);
nor U14746 (N_14746,N_14348,N_14266);
nor U14747 (N_14747,N_14461,N_14456);
nand U14748 (N_14748,N_14377,N_14477);
nor U14749 (N_14749,N_14287,N_14351);
and U14750 (N_14750,N_14723,N_14716);
or U14751 (N_14751,N_14678,N_14706);
xnor U14752 (N_14752,N_14739,N_14525);
or U14753 (N_14753,N_14652,N_14609);
nand U14754 (N_14754,N_14559,N_14568);
nor U14755 (N_14755,N_14746,N_14726);
or U14756 (N_14756,N_14547,N_14731);
xor U14757 (N_14757,N_14643,N_14654);
nor U14758 (N_14758,N_14552,N_14719);
nor U14759 (N_14759,N_14651,N_14641);
xnor U14760 (N_14760,N_14701,N_14680);
nor U14761 (N_14761,N_14734,N_14614);
and U14762 (N_14762,N_14712,N_14695);
xnor U14763 (N_14763,N_14686,N_14645);
and U14764 (N_14764,N_14621,N_14561);
or U14765 (N_14765,N_14676,N_14692);
and U14766 (N_14766,N_14586,N_14718);
nand U14767 (N_14767,N_14679,N_14633);
or U14768 (N_14768,N_14704,N_14653);
nand U14769 (N_14769,N_14579,N_14589);
nor U14770 (N_14770,N_14717,N_14632);
xor U14771 (N_14771,N_14616,N_14677);
xor U14772 (N_14772,N_14593,N_14603);
xor U14773 (N_14773,N_14598,N_14542);
or U14774 (N_14774,N_14737,N_14736);
or U14775 (N_14775,N_14530,N_14630);
xor U14776 (N_14776,N_14534,N_14658);
xor U14777 (N_14777,N_14562,N_14650);
nor U14778 (N_14778,N_14671,N_14572);
xor U14779 (N_14779,N_14606,N_14560);
and U14780 (N_14780,N_14690,N_14748);
or U14781 (N_14781,N_14691,N_14688);
xnor U14782 (N_14782,N_14631,N_14683);
nor U14783 (N_14783,N_14520,N_14581);
and U14784 (N_14784,N_14573,N_14604);
nor U14785 (N_14785,N_14710,N_14529);
xnor U14786 (N_14786,N_14556,N_14564);
nand U14787 (N_14787,N_14672,N_14503);
and U14788 (N_14788,N_14514,N_14656);
and U14789 (N_14789,N_14709,N_14519);
and U14790 (N_14790,N_14728,N_14588);
nand U14791 (N_14791,N_14636,N_14613);
or U14792 (N_14792,N_14545,N_14620);
nand U14793 (N_14793,N_14662,N_14724);
xor U14794 (N_14794,N_14700,N_14553);
and U14795 (N_14795,N_14504,N_14533);
nand U14796 (N_14796,N_14655,N_14659);
and U14797 (N_14797,N_14502,N_14660);
nand U14798 (N_14798,N_14707,N_14565);
xor U14799 (N_14799,N_14708,N_14526);
nor U14800 (N_14800,N_14634,N_14647);
nor U14801 (N_14801,N_14539,N_14596);
nand U14802 (N_14802,N_14580,N_14681);
nor U14803 (N_14803,N_14570,N_14721);
xor U14804 (N_14804,N_14749,N_14578);
or U14805 (N_14805,N_14535,N_14732);
xnor U14806 (N_14806,N_14575,N_14527);
and U14807 (N_14807,N_14674,N_14583);
and U14808 (N_14808,N_14735,N_14720);
or U14809 (N_14809,N_14624,N_14550);
nor U14810 (N_14810,N_14531,N_14639);
nor U14811 (N_14811,N_14536,N_14644);
xor U14812 (N_14812,N_14571,N_14538);
nand U14813 (N_14813,N_14508,N_14629);
or U14814 (N_14814,N_14699,N_14515);
nand U14815 (N_14815,N_14648,N_14611);
nand U14816 (N_14816,N_14738,N_14626);
or U14817 (N_14817,N_14505,N_14500);
nor U14818 (N_14818,N_14698,N_14741);
and U14819 (N_14819,N_14602,N_14615);
nor U14820 (N_14820,N_14541,N_14554);
nand U14821 (N_14821,N_14663,N_14740);
nor U14822 (N_14822,N_14666,N_14612);
or U14823 (N_14823,N_14747,N_14521);
or U14824 (N_14824,N_14516,N_14714);
nand U14825 (N_14825,N_14569,N_14622);
nand U14826 (N_14826,N_14507,N_14585);
xor U14827 (N_14827,N_14594,N_14696);
or U14828 (N_14828,N_14745,N_14694);
nor U14829 (N_14829,N_14517,N_14673);
xor U14830 (N_14830,N_14638,N_14668);
and U14831 (N_14831,N_14591,N_14506);
nor U14832 (N_14832,N_14510,N_14601);
and U14833 (N_14833,N_14693,N_14627);
or U14834 (N_14834,N_14640,N_14744);
nor U14835 (N_14835,N_14513,N_14649);
or U14836 (N_14836,N_14667,N_14608);
or U14837 (N_14837,N_14607,N_14684);
or U14838 (N_14838,N_14628,N_14548);
and U14839 (N_14839,N_14619,N_14544);
nand U14840 (N_14840,N_14713,N_14555);
and U14841 (N_14841,N_14646,N_14549);
nor U14842 (N_14842,N_14528,N_14511);
xor U14843 (N_14843,N_14567,N_14697);
or U14844 (N_14844,N_14635,N_14670);
nand U14845 (N_14845,N_14730,N_14675);
or U14846 (N_14846,N_14543,N_14600);
nor U14847 (N_14847,N_14532,N_14563);
nor U14848 (N_14848,N_14587,N_14623);
and U14849 (N_14849,N_14577,N_14722);
xor U14850 (N_14850,N_14729,N_14566);
or U14851 (N_14851,N_14743,N_14657);
nand U14852 (N_14852,N_14537,N_14509);
and U14853 (N_14853,N_14540,N_14590);
or U14854 (N_14854,N_14557,N_14703);
xnor U14855 (N_14855,N_14551,N_14597);
nand U14856 (N_14856,N_14625,N_14637);
or U14857 (N_14857,N_14733,N_14584);
nor U14858 (N_14858,N_14582,N_14702);
nor U14859 (N_14859,N_14576,N_14642);
nor U14860 (N_14860,N_14661,N_14523);
or U14861 (N_14861,N_14664,N_14727);
nand U14862 (N_14862,N_14558,N_14522);
xnor U14863 (N_14863,N_14574,N_14669);
and U14864 (N_14864,N_14599,N_14711);
and U14865 (N_14865,N_14682,N_14705);
xnor U14866 (N_14866,N_14592,N_14665);
and U14867 (N_14867,N_14689,N_14524);
and U14868 (N_14868,N_14617,N_14725);
xnor U14869 (N_14869,N_14610,N_14501);
xnor U14870 (N_14870,N_14595,N_14605);
nand U14871 (N_14871,N_14518,N_14618);
nand U14872 (N_14872,N_14512,N_14546);
xor U14873 (N_14873,N_14685,N_14742);
or U14874 (N_14874,N_14687,N_14715);
xor U14875 (N_14875,N_14742,N_14650);
or U14876 (N_14876,N_14704,N_14502);
or U14877 (N_14877,N_14553,N_14576);
and U14878 (N_14878,N_14510,N_14722);
or U14879 (N_14879,N_14654,N_14673);
nor U14880 (N_14880,N_14611,N_14515);
and U14881 (N_14881,N_14615,N_14589);
or U14882 (N_14882,N_14611,N_14696);
nor U14883 (N_14883,N_14673,N_14664);
xor U14884 (N_14884,N_14546,N_14659);
and U14885 (N_14885,N_14695,N_14590);
or U14886 (N_14886,N_14685,N_14737);
xnor U14887 (N_14887,N_14684,N_14565);
nor U14888 (N_14888,N_14506,N_14724);
xnor U14889 (N_14889,N_14727,N_14705);
xnor U14890 (N_14890,N_14743,N_14545);
nor U14891 (N_14891,N_14500,N_14512);
and U14892 (N_14892,N_14748,N_14522);
and U14893 (N_14893,N_14509,N_14712);
or U14894 (N_14894,N_14713,N_14526);
xor U14895 (N_14895,N_14520,N_14683);
xor U14896 (N_14896,N_14686,N_14531);
xnor U14897 (N_14897,N_14537,N_14612);
nand U14898 (N_14898,N_14500,N_14593);
nand U14899 (N_14899,N_14551,N_14617);
xnor U14900 (N_14900,N_14685,N_14649);
or U14901 (N_14901,N_14586,N_14739);
nand U14902 (N_14902,N_14717,N_14705);
xor U14903 (N_14903,N_14597,N_14502);
nand U14904 (N_14904,N_14675,N_14683);
or U14905 (N_14905,N_14625,N_14537);
and U14906 (N_14906,N_14579,N_14729);
nor U14907 (N_14907,N_14707,N_14651);
xor U14908 (N_14908,N_14649,N_14726);
nor U14909 (N_14909,N_14740,N_14687);
xor U14910 (N_14910,N_14710,N_14676);
and U14911 (N_14911,N_14737,N_14542);
nand U14912 (N_14912,N_14651,N_14676);
or U14913 (N_14913,N_14558,N_14655);
and U14914 (N_14914,N_14645,N_14579);
and U14915 (N_14915,N_14544,N_14561);
xor U14916 (N_14916,N_14630,N_14737);
nor U14917 (N_14917,N_14610,N_14655);
nor U14918 (N_14918,N_14623,N_14574);
xor U14919 (N_14919,N_14517,N_14741);
nand U14920 (N_14920,N_14666,N_14551);
nor U14921 (N_14921,N_14516,N_14672);
nor U14922 (N_14922,N_14609,N_14690);
nand U14923 (N_14923,N_14714,N_14651);
xor U14924 (N_14924,N_14561,N_14726);
nand U14925 (N_14925,N_14603,N_14621);
and U14926 (N_14926,N_14680,N_14622);
or U14927 (N_14927,N_14647,N_14706);
nand U14928 (N_14928,N_14607,N_14701);
xnor U14929 (N_14929,N_14650,N_14698);
or U14930 (N_14930,N_14732,N_14544);
nor U14931 (N_14931,N_14692,N_14691);
nor U14932 (N_14932,N_14566,N_14743);
nand U14933 (N_14933,N_14512,N_14603);
xnor U14934 (N_14934,N_14532,N_14521);
nor U14935 (N_14935,N_14582,N_14668);
xnor U14936 (N_14936,N_14535,N_14575);
and U14937 (N_14937,N_14712,N_14572);
or U14938 (N_14938,N_14709,N_14664);
and U14939 (N_14939,N_14667,N_14536);
and U14940 (N_14940,N_14623,N_14593);
xnor U14941 (N_14941,N_14631,N_14624);
or U14942 (N_14942,N_14641,N_14739);
or U14943 (N_14943,N_14635,N_14694);
or U14944 (N_14944,N_14665,N_14608);
or U14945 (N_14945,N_14674,N_14642);
nand U14946 (N_14946,N_14577,N_14711);
or U14947 (N_14947,N_14604,N_14650);
and U14948 (N_14948,N_14594,N_14597);
xor U14949 (N_14949,N_14689,N_14611);
or U14950 (N_14950,N_14736,N_14586);
nor U14951 (N_14951,N_14658,N_14645);
nor U14952 (N_14952,N_14581,N_14664);
nand U14953 (N_14953,N_14542,N_14662);
xnor U14954 (N_14954,N_14610,N_14719);
xor U14955 (N_14955,N_14596,N_14589);
or U14956 (N_14956,N_14742,N_14724);
and U14957 (N_14957,N_14581,N_14528);
or U14958 (N_14958,N_14597,N_14729);
xnor U14959 (N_14959,N_14510,N_14727);
or U14960 (N_14960,N_14541,N_14583);
xor U14961 (N_14961,N_14676,N_14622);
xor U14962 (N_14962,N_14611,N_14587);
xnor U14963 (N_14963,N_14562,N_14553);
nor U14964 (N_14964,N_14612,N_14722);
or U14965 (N_14965,N_14729,N_14719);
nor U14966 (N_14966,N_14659,N_14684);
nor U14967 (N_14967,N_14738,N_14541);
and U14968 (N_14968,N_14673,N_14737);
and U14969 (N_14969,N_14718,N_14507);
xnor U14970 (N_14970,N_14717,N_14589);
xnor U14971 (N_14971,N_14728,N_14687);
nor U14972 (N_14972,N_14674,N_14719);
nor U14973 (N_14973,N_14608,N_14576);
and U14974 (N_14974,N_14747,N_14558);
or U14975 (N_14975,N_14746,N_14617);
and U14976 (N_14976,N_14665,N_14548);
nor U14977 (N_14977,N_14730,N_14670);
and U14978 (N_14978,N_14533,N_14527);
or U14979 (N_14979,N_14690,N_14696);
or U14980 (N_14980,N_14641,N_14552);
nand U14981 (N_14981,N_14610,N_14731);
nor U14982 (N_14982,N_14572,N_14706);
or U14983 (N_14983,N_14519,N_14653);
xor U14984 (N_14984,N_14598,N_14736);
nor U14985 (N_14985,N_14660,N_14639);
nand U14986 (N_14986,N_14637,N_14653);
nand U14987 (N_14987,N_14548,N_14706);
or U14988 (N_14988,N_14627,N_14670);
nand U14989 (N_14989,N_14520,N_14647);
and U14990 (N_14990,N_14697,N_14531);
nand U14991 (N_14991,N_14518,N_14700);
nand U14992 (N_14992,N_14567,N_14725);
or U14993 (N_14993,N_14509,N_14526);
xor U14994 (N_14994,N_14625,N_14660);
and U14995 (N_14995,N_14712,N_14709);
and U14996 (N_14996,N_14532,N_14723);
xor U14997 (N_14997,N_14537,N_14579);
nand U14998 (N_14998,N_14654,N_14619);
nand U14999 (N_14999,N_14630,N_14543);
or U15000 (N_15000,N_14922,N_14789);
and U15001 (N_15001,N_14897,N_14819);
or U15002 (N_15002,N_14987,N_14860);
nand U15003 (N_15003,N_14785,N_14930);
xor U15004 (N_15004,N_14841,N_14985);
nand U15005 (N_15005,N_14852,N_14793);
and U15006 (N_15006,N_14847,N_14936);
xnor U15007 (N_15007,N_14774,N_14782);
nor U15008 (N_15008,N_14772,N_14815);
or U15009 (N_15009,N_14857,N_14984);
and U15010 (N_15010,N_14812,N_14754);
and U15011 (N_15011,N_14794,N_14907);
nor U15012 (N_15012,N_14769,N_14947);
nand U15013 (N_15013,N_14955,N_14993);
or U15014 (N_15014,N_14824,N_14872);
or U15015 (N_15015,N_14874,N_14864);
or U15016 (N_15016,N_14898,N_14931);
or U15017 (N_15017,N_14953,N_14879);
nor U15018 (N_15018,N_14952,N_14972);
and U15019 (N_15019,N_14834,N_14763);
nor U15020 (N_15020,N_14918,N_14884);
xnor U15021 (N_15021,N_14883,N_14989);
xor U15022 (N_15022,N_14753,N_14777);
or U15023 (N_15023,N_14968,N_14944);
nand U15024 (N_15024,N_14980,N_14795);
nor U15025 (N_15025,N_14771,N_14758);
nor U15026 (N_15026,N_14784,N_14896);
nand U15027 (N_15027,N_14928,N_14837);
and U15028 (N_15028,N_14926,N_14895);
and U15029 (N_15029,N_14958,N_14919);
or U15030 (N_15030,N_14942,N_14781);
nand U15031 (N_15031,N_14813,N_14760);
or U15032 (N_15032,N_14877,N_14996);
or U15033 (N_15033,N_14957,N_14975);
and U15034 (N_15034,N_14910,N_14773);
or U15035 (N_15035,N_14988,N_14850);
nor U15036 (N_15036,N_14970,N_14808);
or U15037 (N_15037,N_14783,N_14962);
nand U15038 (N_15038,N_14807,N_14855);
and U15039 (N_15039,N_14776,N_14854);
nor U15040 (N_15040,N_14779,N_14905);
xnor U15041 (N_15041,N_14961,N_14849);
xor U15042 (N_15042,N_14890,N_14868);
xnor U15043 (N_15043,N_14971,N_14799);
nand U15044 (N_15044,N_14950,N_14899);
nor U15045 (N_15045,N_14888,N_14938);
or U15046 (N_15046,N_14792,N_14940);
and U15047 (N_15047,N_14796,N_14933);
nor U15048 (N_15048,N_14932,N_14904);
nor U15049 (N_15049,N_14999,N_14983);
nand U15050 (N_15050,N_14851,N_14903);
xor U15051 (N_15051,N_14966,N_14889);
nand U15052 (N_15052,N_14780,N_14979);
and U15053 (N_15053,N_14960,N_14752);
and U15054 (N_15054,N_14762,N_14863);
nand U15055 (N_15055,N_14786,N_14892);
nor U15056 (N_15056,N_14801,N_14924);
nor U15057 (N_15057,N_14990,N_14790);
or U15058 (N_15058,N_14916,N_14912);
and U15059 (N_15059,N_14839,N_14973);
and U15060 (N_15060,N_14943,N_14830);
nor U15061 (N_15061,N_14964,N_14963);
or U15062 (N_15062,N_14817,N_14775);
nor U15063 (N_15063,N_14804,N_14859);
nor U15064 (N_15064,N_14937,N_14818);
or U15065 (N_15065,N_14978,N_14767);
nand U15066 (N_15066,N_14981,N_14836);
or U15067 (N_15067,N_14921,N_14814);
nor U15068 (N_15068,N_14977,N_14894);
and U15069 (N_15069,N_14831,N_14967);
nand U15070 (N_15070,N_14828,N_14913);
or U15071 (N_15071,N_14842,N_14810);
nand U15072 (N_15072,N_14951,N_14846);
nand U15073 (N_15073,N_14909,N_14923);
xnor U15074 (N_15074,N_14927,N_14991);
and U15075 (N_15075,N_14756,N_14976);
or U15076 (N_15076,N_14862,N_14750);
nor U15077 (N_15077,N_14866,N_14901);
xor U15078 (N_15078,N_14833,N_14844);
or U15079 (N_15079,N_14875,N_14994);
nand U15080 (N_15080,N_14803,N_14838);
and U15081 (N_15081,N_14856,N_14827);
or U15082 (N_15082,N_14759,N_14823);
nand U15083 (N_15083,N_14885,N_14881);
nor U15084 (N_15084,N_14802,N_14992);
nand U15085 (N_15085,N_14997,N_14826);
nand U15086 (N_15086,N_14969,N_14959);
nand U15087 (N_15087,N_14805,N_14878);
nor U15088 (N_15088,N_14925,N_14867);
nor U15089 (N_15089,N_14800,N_14766);
and U15090 (N_15090,N_14935,N_14788);
nor U15091 (N_15091,N_14954,N_14755);
or U15092 (N_15092,N_14797,N_14900);
or U15093 (N_15093,N_14920,N_14809);
or U15094 (N_15094,N_14914,N_14902);
and U15095 (N_15095,N_14848,N_14886);
nor U15096 (N_15096,N_14853,N_14820);
or U15097 (N_15097,N_14858,N_14845);
nor U15098 (N_15098,N_14840,N_14939);
nor U15099 (N_15099,N_14761,N_14934);
xor U15100 (N_15100,N_14843,N_14765);
or U15101 (N_15101,N_14751,N_14880);
and U15102 (N_15102,N_14948,N_14757);
xor U15103 (N_15103,N_14806,N_14816);
and U15104 (N_15104,N_14891,N_14835);
nor U15105 (N_15105,N_14882,N_14825);
xnor U15106 (N_15106,N_14869,N_14941);
xor U15107 (N_15107,N_14873,N_14821);
nor U15108 (N_15108,N_14798,N_14945);
nand U15109 (N_15109,N_14871,N_14764);
or U15110 (N_15110,N_14887,N_14956);
or U15111 (N_15111,N_14768,N_14865);
nand U15112 (N_15112,N_14949,N_14995);
or U15113 (N_15113,N_14893,N_14998);
or U15114 (N_15114,N_14787,N_14811);
xor U15115 (N_15115,N_14908,N_14876);
xnor U15116 (N_15116,N_14915,N_14986);
nor U15117 (N_15117,N_14861,N_14778);
and U15118 (N_15118,N_14982,N_14965);
xnor U15119 (N_15119,N_14822,N_14906);
nor U15120 (N_15120,N_14832,N_14829);
or U15121 (N_15121,N_14974,N_14917);
nand U15122 (N_15122,N_14929,N_14870);
nor U15123 (N_15123,N_14791,N_14911);
xor U15124 (N_15124,N_14946,N_14770);
nand U15125 (N_15125,N_14785,N_14791);
nor U15126 (N_15126,N_14774,N_14894);
or U15127 (N_15127,N_14966,N_14998);
xor U15128 (N_15128,N_14803,N_14856);
nor U15129 (N_15129,N_14911,N_14998);
nand U15130 (N_15130,N_14801,N_14850);
and U15131 (N_15131,N_14894,N_14982);
xor U15132 (N_15132,N_14802,N_14977);
or U15133 (N_15133,N_14952,N_14980);
nor U15134 (N_15134,N_14903,N_14935);
nor U15135 (N_15135,N_14882,N_14842);
nand U15136 (N_15136,N_14812,N_14960);
nor U15137 (N_15137,N_14927,N_14887);
xnor U15138 (N_15138,N_14825,N_14960);
nand U15139 (N_15139,N_14861,N_14876);
nor U15140 (N_15140,N_14977,N_14784);
xor U15141 (N_15141,N_14944,N_14793);
xnor U15142 (N_15142,N_14911,N_14854);
nand U15143 (N_15143,N_14856,N_14844);
and U15144 (N_15144,N_14801,N_14786);
nor U15145 (N_15145,N_14998,N_14974);
xnor U15146 (N_15146,N_14830,N_14762);
xnor U15147 (N_15147,N_14900,N_14927);
nor U15148 (N_15148,N_14825,N_14856);
nand U15149 (N_15149,N_14762,N_14876);
and U15150 (N_15150,N_14793,N_14809);
nand U15151 (N_15151,N_14800,N_14750);
nand U15152 (N_15152,N_14766,N_14857);
and U15153 (N_15153,N_14783,N_14844);
xnor U15154 (N_15154,N_14830,N_14978);
xor U15155 (N_15155,N_14941,N_14820);
nand U15156 (N_15156,N_14873,N_14946);
xnor U15157 (N_15157,N_14908,N_14937);
nand U15158 (N_15158,N_14760,N_14931);
or U15159 (N_15159,N_14971,N_14871);
xor U15160 (N_15160,N_14861,N_14912);
and U15161 (N_15161,N_14826,N_14996);
xnor U15162 (N_15162,N_14850,N_14813);
and U15163 (N_15163,N_14963,N_14871);
nor U15164 (N_15164,N_14758,N_14897);
nor U15165 (N_15165,N_14753,N_14885);
and U15166 (N_15166,N_14789,N_14803);
nand U15167 (N_15167,N_14998,N_14764);
and U15168 (N_15168,N_14955,N_14981);
or U15169 (N_15169,N_14786,N_14777);
nand U15170 (N_15170,N_14980,N_14854);
xor U15171 (N_15171,N_14823,N_14939);
xnor U15172 (N_15172,N_14754,N_14974);
xor U15173 (N_15173,N_14992,N_14979);
nor U15174 (N_15174,N_14778,N_14780);
or U15175 (N_15175,N_14750,N_14787);
nand U15176 (N_15176,N_14849,N_14881);
nor U15177 (N_15177,N_14918,N_14852);
or U15178 (N_15178,N_14783,N_14840);
or U15179 (N_15179,N_14871,N_14781);
xor U15180 (N_15180,N_14956,N_14874);
or U15181 (N_15181,N_14949,N_14866);
nand U15182 (N_15182,N_14780,N_14976);
nor U15183 (N_15183,N_14932,N_14992);
nor U15184 (N_15184,N_14755,N_14913);
nand U15185 (N_15185,N_14905,N_14971);
nand U15186 (N_15186,N_14758,N_14930);
nor U15187 (N_15187,N_14967,N_14771);
or U15188 (N_15188,N_14857,N_14922);
xor U15189 (N_15189,N_14765,N_14866);
or U15190 (N_15190,N_14916,N_14809);
nand U15191 (N_15191,N_14966,N_14957);
nand U15192 (N_15192,N_14927,N_14820);
nand U15193 (N_15193,N_14961,N_14921);
nor U15194 (N_15194,N_14821,N_14924);
xor U15195 (N_15195,N_14785,N_14877);
and U15196 (N_15196,N_14916,N_14982);
nand U15197 (N_15197,N_14791,N_14957);
xnor U15198 (N_15198,N_14861,N_14879);
nor U15199 (N_15199,N_14917,N_14837);
nor U15200 (N_15200,N_14952,N_14985);
and U15201 (N_15201,N_14842,N_14868);
nand U15202 (N_15202,N_14771,N_14965);
or U15203 (N_15203,N_14836,N_14917);
xnor U15204 (N_15204,N_14792,N_14875);
and U15205 (N_15205,N_14948,N_14778);
xor U15206 (N_15206,N_14948,N_14998);
and U15207 (N_15207,N_14903,N_14889);
nor U15208 (N_15208,N_14832,N_14870);
xnor U15209 (N_15209,N_14998,N_14793);
or U15210 (N_15210,N_14850,N_14847);
or U15211 (N_15211,N_14843,N_14874);
nand U15212 (N_15212,N_14899,N_14775);
or U15213 (N_15213,N_14807,N_14769);
nor U15214 (N_15214,N_14905,N_14984);
or U15215 (N_15215,N_14997,N_14812);
or U15216 (N_15216,N_14945,N_14869);
xor U15217 (N_15217,N_14966,N_14902);
or U15218 (N_15218,N_14977,N_14758);
xor U15219 (N_15219,N_14796,N_14767);
nor U15220 (N_15220,N_14912,N_14997);
nand U15221 (N_15221,N_14930,N_14789);
or U15222 (N_15222,N_14842,N_14763);
and U15223 (N_15223,N_14756,N_14901);
nand U15224 (N_15224,N_14907,N_14965);
xnor U15225 (N_15225,N_14822,N_14839);
xor U15226 (N_15226,N_14811,N_14904);
and U15227 (N_15227,N_14927,N_14788);
and U15228 (N_15228,N_14825,N_14788);
nor U15229 (N_15229,N_14870,N_14861);
nor U15230 (N_15230,N_14899,N_14838);
nand U15231 (N_15231,N_14947,N_14856);
xnor U15232 (N_15232,N_14915,N_14875);
or U15233 (N_15233,N_14901,N_14879);
nor U15234 (N_15234,N_14836,N_14761);
nand U15235 (N_15235,N_14794,N_14770);
nor U15236 (N_15236,N_14925,N_14817);
nor U15237 (N_15237,N_14900,N_14798);
nor U15238 (N_15238,N_14761,N_14984);
or U15239 (N_15239,N_14944,N_14876);
and U15240 (N_15240,N_14886,N_14891);
nand U15241 (N_15241,N_14886,N_14857);
and U15242 (N_15242,N_14874,N_14989);
nand U15243 (N_15243,N_14933,N_14961);
xnor U15244 (N_15244,N_14844,N_14966);
nor U15245 (N_15245,N_14846,N_14845);
xor U15246 (N_15246,N_14831,N_14764);
or U15247 (N_15247,N_14752,N_14776);
and U15248 (N_15248,N_14931,N_14817);
and U15249 (N_15249,N_14951,N_14959);
nor U15250 (N_15250,N_15144,N_15200);
xor U15251 (N_15251,N_15019,N_15039);
nor U15252 (N_15252,N_15156,N_15176);
xnor U15253 (N_15253,N_15004,N_15230);
xor U15254 (N_15254,N_15160,N_15115);
xnor U15255 (N_15255,N_15161,N_15110);
nor U15256 (N_15256,N_15113,N_15243);
and U15257 (N_15257,N_15009,N_15193);
nand U15258 (N_15258,N_15090,N_15025);
xnor U15259 (N_15259,N_15136,N_15005);
or U15260 (N_15260,N_15049,N_15219);
xnor U15261 (N_15261,N_15105,N_15178);
and U15262 (N_15262,N_15024,N_15124);
and U15263 (N_15263,N_15053,N_15184);
nand U15264 (N_15264,N_15187,N_15033);
xor U15265 (N_15265,N_15083,N_15194);
xor U15266 (N_15266,N_15235,N_15065);
xor U15267 (N_15267,N_15223,N_15006);
or U15268 (N_15268,N_15060,N_15249);
xor U15269 (N_15269,N_15035,N_15102);
nand U15270 (N_15270,N_15153,N_15190);
nand U15271 (N_15271,N_15087,N_15179);
and U15272 (N_15272,N_15042,N_15239);
nor U15273 (N_15273,N_15040,N_15133);
and U15274 (N_15274,N_15180,N_15037);
xnor U15275 (N_15275,N_15198,N_15245);
nand U15276 (N_15276,N_15028,N_15181);
nor U15277 (N_15277,N_15012,N_15208);
or U15278 (N_15278,N_15112,N_15203);
nand U15279 (N_15279,N_15212,N_15150);
xnor U15280 (N_15280,N_15206,N_15071);
and U15281 (N_15281,N_15074,N_15159);
and U15282 (N_15282,N_15134,N_15072);
and U15283 (N_15283,N_15224,N_15000);
nand U15284 (N_15284,N_15215,N_15027);
nand U15285 (N_15285,N_15056,N_15097);
xnor U15286 (N_15286,N_15066,N_15158);
nand U15287 (N_15287,N_15069,N_15070);
xnor U15288 (N_15288,N_15022,N_15142);
xor U15289 (N_15289,N_15196,N_15141);
or U15290 (N_15290,N_15020,N_15058);
and U15291 (N_15291,N_15104,N_15084);
xor U15292 (N_15292,N_15211,N_15163);
nand U15293 (N_15293,N_15234,N_15085);
xnor U15294 (N_15294,N_15011,N_15120);
nand U15295 (N_15295,N_15086,N_15157);
or U15296 (N_15296,N_15242,N_15041);
nor U15297 (N_15297,N_15057,N_15067);
and U15298 (N_15298,N_15147,N_15199);
nor U15299 (N_15299,N_15207,N_15076);
xor U15300 (N_15300,N_15015,N_15244);
nor U15301 (N_15301,N_15195,N_15095);
nor U15302 (N_15302,N_15192,N_15117);
or U15303 (N_15303,N_15061,N_15197);
xor U15304 (N_15304,N_15132,N_15055);
nor U15305 (N_15305,N_15233,N_15118);
nand U15306 (N_15306,N_15143,N_15127);
and U15307 (N_15307,N_15201,N_15099);
and U15308 (N_15308,N_15229,N_15031);
or U15309 (N_15309,N_15044,N_15050);
nand U15310 (N_15310,N_15106,N_15247);
nor U15311 (N_15311,N_15016,N_15107);
and U15312 (N_15312,N_15029,N_15231);
and U15313 (N_15313,N_15240,N_15214);
nand U15314 (N_15314,N_15051,N_15092);
xor U15315 (N_15315,N_15116,N_15126);
nor U15316 (N_15316,N_15226,N_15149);
and U15317 (N_15317,N_15202,N_15173);
or U15318 (N_15318,N_15155,N_15222);
nor U15319 (N_15319,N_15248,N_15008);
xor U15320 (N_15320,N_15034,N_15032);
nand U15321 (N_15321,N_15013,N_15186);
nor U15322 (N_15322,N_15236,N_15122);
or U15323 (N_15323,N_15175,N_15183);
and U15324 (N_15324,N_15209,N_15169);
nand U15325 (N_15325,N_15054,N_15036);
and U15326 (N_15326,N_15172,N_15177);
nand U15327 (N_15327,N_15148,N_15062);
xor U15328 (N_15328,N_15026,N_15114);
and U15329 (N_15329,N_15128,N_15129);
nor U15330 (N_15330,N_15137,N_15080);
nor U15331 (N_15331,N_15052,N_15100);
and U15332 (N_15332,N_15151,N_15213);
and U15333 (N_15333,N_15185,N_15079);
nor U15334 (N_15334,N_15154,N_15189);
xnor U15335 (N_15335,N_15135,N_15131);
and U15336 (N_15336,N_15123,N_15089);
xnor U15337 (N_15337,N_15002,N_15077);
and U15338 (N_15338,N_15017,N_15125);
and U15339 (N_15339,N_15038,N_15010);
xor U15340 (N_15340,N_15238,N_15188);
xor U15341 (N_15341,N_15146,N_15237);
nor U15342 (N_15342,N_15216,N_15210);
or U15343 (N_15343,N_15059,N_15218);
xnor U15344 (N_15344,N_15164,N_15167);
or U15345 (N_15345,N_15093,N_15109);
xor U15346 (N_15346,N_15241,N_15166);
or U15347 (N_15347,N_15182,N_15003);
nand U15348 (N_15348,N_15217,N_15007);
xor U15349 (N_15349,N_15101,N_15048);
or U15350 (N_15350,N_15171,N_15023);
or U15351 (N_15351,N_15030,N_15091);
or U15352 (N_15352,N_15227,N_15073);
xor U15353 (N_15353,N_15021,N_15111);
xor U15354 (N_15354,N_15145,N_15168);
nor U15355 (N_15355,N_15043,N_15221);
nor U15356 (N_15356,N_15191,N_15121);
xor U15357 (N_15357,N_15170,N_15139);
nand U15358 (N_15358,N_15047,N_15075);
or U15359 (N_15359,N_15068,N_15063);
xnor U15360 (N_15360,N_15119,N_15246);
or U15361 (N_15361,N_15018,N_15205);
nor U15362 (N_15362,N_15096,N_15064);
nor U15363 (N_15363,N_15045,N_15001);
nor U15364 (N_15364,N_15232,N_15152);
nor U15365 (N_15365,N_15228,N_15140);
nor U15366 (N_15366,N_15165,N_15204);
or U15367 (N_15367,N_15138,N_15098);
nand U15368 (N_15368,N_15088,N_15082);
nor U15369 (N_15369,N_15046,N_15103);
or U15370 (N_15370,N_15108,N_15094);
xnor U15371 (N_15371,N_15225,N_15220);
nor U15372 (N_15372,N_15081,N_15174);
nand U15373 (N_15373,N_15130,N_15078);
and U15374 (N_15374,N_15014,N_15162);
or U15375 (N_15375,N_15019,N_15065);
nand U15376 (N_15376,N_15085,N_15025);
xnor U15377 (N_15377,N_15187,N_15107);
and U15378 (N_15378,N_15135,N_15108);
xor U15379 (N_15379,N_15006,N_15153);
and U15380 (N_15380,N_15234,N_15203);
and U15381 (N_15381,N_15156,N_15070);
or U15382 (N_15382,N_15096,N_15093);
and U15383 (N_15383,N_15125,N_15165);
nor U15384 (N_15384,N_15081,N_15138);
nor U15385 (N_15385,N_15056,N_15163);
nor U15386 (N_15386,N_15058,N_15195);
nand U15387 (N_15387,N_15055,N_15007);
nand U15388 (N_15388,N_15106,N_15238);
xnor U15389 (N_15389,N_15187,N_15002);
and U15390 (N_15390,N_15055,N_15161);
and U15391 (N_15391,N_15122,N_15042);
or U15392 (N_15392,N_15121,N_15144);
xnor U15393 (N_15393,N_15055,N_15054);
or U15394 (N_15394,N_15096,N_15160);
nor U15395 (N_15395,N_15083,N_15161);
and U15396 (N_15396,N_15143,N_15163);
nor U15397 (N_15397,N_15015,N_15223);
nand U15398 (N_15398,N_15110,N_15102);
nand U15399 (N_15399,N_15096,N_15050);
or U15400 (N_15400,N_15174,N_15121);
or U15401 (N_15401,N_15067,N_15244);
nand U15402 (N_15402,N_15208,N_15182);
nor U15403 (N_15403,N_15149,N_15049);
or U15404 (N_15404,N_15230,N_15211);
nor U15405 (N_15405,N_15223,N_15134);
or U15406 (N_15406,N_15158,N_15065);
xnor U15407 (N_15407,N_15039,N_15237);
and U15408 (N_15408,N_15199,N_15009);
or U15409 (N_15409,N_15116,N_15104);
or U15410 (N_15410,N_15013,N_15065);
xor U15411 (N_15411,N_15182,N_15199);
xor U15412 (N_15412,N_15089,N_15088);
nor U15413 (N_15413,N_15140,N_15017);
or U15414 (N_15414,N_15070,N_15030);
nand U15415 (N_15415,N_15126,N_15110);
xor U15416 (N_15416,N_15123,N_15199);
nor U15417 (N_15417,N_15007,N_15077);
xor U15418 (N_15418,N_15247,N_15149);
or U15419 (N_15419,N_15168,N_15215);
xor U15420 (N_15420,N_15093,N_15076);
nor U15421 (N_15421,N_15180,N_15031);
or U15422 (N_15422,N_15122,N_15068);
nor U15423 (N_15423,N_15081,N_15013);
or U15424 (N_15424,N_15171,N_15098);
xor U15425 (N_15425,N_15105,N_15146);
nor U15426 (N_15426,N_15024,N_15039);
or U15427 (N_15427,N_15188,N_15244);
nor U15428 (N_15428,N_15194,N_15147);
and U15429 (N_15429,N_15188,N_15139);
or U15430 (N_15430,N_15127,N_15102);
nor U15431 (N_15431,N_15114,N_15021);
and U15432 (N_15432,N_15140,N_15034);
xnor U15433 (N_15433,N_15248,N_15074);
nand U15434 (N_15434,N_15051,N_15137);
and U15435 (N_15435,N_15137,N_15188);
or U15436 (N_15436,N_15157,N_15111);
nor U15437 (N_15437,N_15055,N_15120);
xnor U15438 (N_15438,N_15058,N_15189);
nor U15439 (N_15439,N_15237,N_15012);
nor U15440 (N_15440,N_15234,N_15191);
xnor U15441 (N_15441,N_15067,N_15010);
nand U15442 (N_15442,N_15091,N_15044);
or U15443 (N_15443,N_15170,N_15231);
nand U15444 (N_15444,N_15001,N_15007);
and U15445 (N_15445,N_15120,N_15242);
or U15446 (N_15446,N_15156,N_15238);
xor U15447 (N_15447,N_15016,N_15113);
nand U15448 (N_15448,N_15111,N_15175);
nor U15449 (N_15449,N_15187,N_15106);
nor U15450 (N_15450,N_15106,N_15230);
nor U15451 (N_15451,N_15000,N_15164);
nor U15452 (N_15452,N_15182,N_15228);
nand U15453 (N_15453,N_15107,N_15125);
and U15454 (N_15454,N_15133,N_15215);
nand U15455 (N_15455,N_15038,N_15245);
nand U15456 (N_15456,N_15198,N_15012);
nor U15457 (N_15457,N_15014,N_15066);
or U15458 (N_15458,N_15236,N_15006);
nor U15459 (N_15459,N_15234,N_15099);
or U15460 (N_15460,N_15009,N_15068);
nor U15461 (N_15461,N_15142,N_15101);
xor U15462 (N_15462,N_15066,N_15169);
nand U15463 (N_15463,N_15150,N_15067);
nor U15464 (N_15464,N_15105,N_15022);
and U15465 (N_15465,N_15028,N_15154);
xor U15466 (N_15466,N_15013,N_15187);
or U15467 (N_15467,N_15144,N_15033);
nand U15468 (N_15468,N_15091,N_15204);
or U15469 (N_15469,N_15182,N_15122);
xnor U15470 (N_15470,N_15234,N_15216);
xor U15471 (N_15471,N_15011,N_15170);
nor U15472 (N_15472,N_15064,N_15033);
and U15473 (N_15473,N_15024,N_15063);
xor U15474 (N_15474,N_15178,N_15131);
nor U15475 (N_15475,N_15183,N_15249);
xnor U15476 (N_15476,N_15232,N_15235);
and U15477 (N_15477,N_15083,N_15204);
nor U15478 (N_15478,N_15150,N_15130);
nand U15479 (N_15479,N_15062,N_15200);
nor U15480 (N_15480,N_15015,N_15051);
nand U15481 (N_15481,N_15060,N_15049);
nand U15482 (N_15482,N_15010,N_15044);
nor U15483 (N_15483,N_15176,N_15208);
and U15484 (N_15484,N_15148,N_15015);
and U15485 (N_15485,N_15129,N_15153);
nand U15486 (N_15486,N_15074,N_15111);
xor U15487 (N_15487,N_15236,N_15050);
and U15488 (N_15488,N_15017,N_15036);
or U15489 (N_15489,N_15014,N_15153);
or U15490 (N_15490,N_15164,N_15233);
and U15491 (N_15491,N_15208,N_15004);
and U15492 (N_15492,N_15150,N_15041);
or U15493 (N_15493,N_15040,N_15230);
nand U15494 (N_15494,N_15204,N_15052);
and U15495 (N_15495,N_15202,N_15121);
nor U15496 (N_15496,N_15073,N_15110);
or U15497 (N_15497,N_15205,N_15083);
and U15498 (N_15498,N_15078,N_15154);
nor U15499 (N_15499,N_15127,N_15005);
and U15500 (N_15500,N_15455,N_15357);
or U15501 (N_15501,N_15396,N_15361);
or U15502 (N_15502,N_15443,N_15330);
xnor U15503 (N_15503,N_15311,N_15351);
nor U15504 (N_15504,N_15288,N_15360);
or U15505 (N_15505,N_15260,N_15449);
xnor U15506 (N_15506,N_15477,N_15444);
nand U15507 (N_15507,N_15334,N_15306);
xnor U15508 (N_15508,N_15358,N_15349);
nand U15509 (N_15509,N_15251,N_15340);
nand U15510 (N_15510,N_15400,N_15370);
xnor U15511 (N_15511,N_15322,N_15498);
or U15512 (N_15512,N_15406,N_15258);
nor U15513 (N_15513,N_15347,N_15293);
nand U15514 (N_15514,N_15423,N_15331);
nor U15515 (N_15515,N_15422,N_15289);
xor U15516 (N_15516,N_15494,N_15415);
and U15517 (N_15517,N_15426,N_15384);
nor U15518 (N_15518,N_15395,N_15467);
nand U15519 (N_15519,N_15453,N_15442);
and U15520 (N_15520,N_15424,N_15259);
nand U15521 (N_15521,N_15333,N_15393);
nor U15522 (N_15522,N_15417,N_15488);
xnor U15523 (N_15523,N_15475,N_15389);
nor U15524 (N_15524,N_15405,N_15362);
nor U15525 (N_15525,N_15277,N_15356);
and U15526 (N_15526,N_15425,N_15404);
or U15527 (N_15527,N_15294,N_15390);
and U15528 (N_15528,N_15471,N_15374);
or U15529 (N_15529,N_15397,N_15271);
xnor U15530 (N_15530,N_15250,N_15491);
xor U15531 (N_15531,N_15428,N_15391);
nor U15532 (N_15532,N_15291,N_15399);
and U15533 (N_15533,N_15269,N_15355);
nand U15534 (N_15534,N_15452,N_15383);
nand U15535 (N_15535,N_15478,N_15278);
or U15536 (N_15536,N_15286,N_15439);
nand U15537 (N_15537,N_15285,N_15401);
or U15538 (N_15538,N_15495,N_15298);
nor U15539 (N_15539,N_15261,N_15433);
nand U15540 (N_15540,N_15377,N_15480);
xor U15541 (N_15541,N_15402,N_15466);
xnor U15542 (N_15542,N_15359,N_15486);
xnor U15543 (N_15543,N_15382,N_15420);
and U15544 (N_15544,N_15499,N_15380);
or U15545 (N_15545,N_15476,N_15308);
xor U15546 (N_15546,N_15493,N_15348);
xor U15547 (N_15547,N_15469,N_15437);
and U15548 (N_15548,N_15295,N_15473);
nand U15549 (N_15549,N_15350,N_15353);
and U15550 (N_15550,N_15314,N_15465);
xor U15551 (N_15551,N_15373,N_15416);
or U15552 (N_15552,N_15345,N_15497);
nand U15553 (N_15553,N_15335,N_15323);
nor U15554 (N_15554,N_15301,N_15409);
and U15555 (N_15555,N_15315,N_15454);
or U15556 (N_15556,N_15440,N_15435);
nor U15557 (N_15557,N_15307,N_15273);
and U15558 (N_15558,N_15328,N_15282);
and U15559 (N_15559,N_15253,N_15341);
nor U15560 (N_15560,N_15317,N_15367);
xnor U15561 (N_15561,N_15281,N_15385);
or U15562 (N_15562,N_15290,N_15318);
and U15563 (N_15563,N_15324,N_15411);
nor U15564 (N_15564,N_15352,N_15427);
nor U15565 (N_15565,N_15303,N_15487);
nand U15566 (N_15566,N_15448,N_15305);
xor U15567 (N_15567,N_15490,N_15263);
xnor U15568 (N_15568,N_15387,N_15421);
xnor U15569 (N_15569,N_15326,N_15280);
nand U15570 (N_15570,N_15458,N_15388);
or U15571 (N_15571,N_15252,N_15403);
xor U15572 (N_15572,N_15254,N_15354);
xor U15573 (N_15573,N_15451,N_15375);
nor U15574 (N_15574,N_15284,N_15394);
nor U15575 (N_15575,N_15321,N_15434);
xor U15576 (N_15576,N_15343,N_15468);
or U15577 (N_15577,N_15445,N_15381);
nor U15578 (N_15578,N_15472,N_15392);
and U15579 (N_15579,N_15429,N_15386);
and U15580 (N_15580,N_15270,N_15274);
or U15581 (N_15581,N_15398,N_15272);
and U15582 (N_15582,N_15310,N_15446);
or U15583 (N_15583,N_15257,N_15438);
xor U15584 (N_15584,N_15264,N_15456);
nor U15585 (N_15585,N_15275,N_15297);
nor U15586 (N_15586,N_15329,N_15292);
and U15587 (N_15587,N_15459,N_15408);
nand U15588 (N_15588,N_15450,N_15484);
and U15589 (N_15589,N_15441,N_15460);
or U15590 (N_15590,N_15346,N_15461);
and U15591 (N_15591,N_15489,N_15332);
xnor U15592 (N_15592,N_15363,N_15463);
nor U15593 (N_15593,N_15312,N_15481);
and U15594 (N_15594,N_15483,N_15365);
and U15595 (N_15595,N_15485,N_15430);
and U15596 (N_15596,N_15319,N_15320);
or U15597 (N_15597,N_15267,N_15470);
nor U15598 (N_15598,N_15302,N_15464);
or U15599 (N_15599,N_15378,N_15407);
xor U15600 (N_15600,N_15496,N_15457);
nand U15601 (N_15601,N_15304,N_15342);
xnor U15602 (N_15602,N_15283,N_15418);
and U15603 (N_15603,N_15431,N_15279);
xor U15604 (N_15604,N_15276,N_15265);
xor U15605 (N_15605,N_15339,N_15338);
and U15606 (N_15606,N_15432,N_15366);
and U15607 (N_15607,N_15337,N_15410);
nor U15608 (N_15608,N_15364,N_15413);
xnor U15609 (N_15609,N_15325,N_15419);
nand U15610 (N_15610,N_15462,N_15256);
xor U15611 (N_15611,N_15379,N_15376);
xor U15612 (N_15612,N_15492,N_15296);
or U15613 (N_15613,N_15371,N_15336);
or U15614 (N_15614,N_15299,N_15447);
and U15615 (N_15615,N_15316,N_15479);
xor U15616 (N_15616,N_15268,N_15309);
or U15617 (N_15617,N_15300,N_15262);
and U15618 (N_15618,N_15344,N_15474);
nand U15619 (N_15619,N_15436,N_15327);
and U15620 (N_15620,N_15412,N_15368);
nor U15621 (N_15621,N_15482,N_15266);
xor U15622 (N_15622,N_15372,N_15414);
nand U15623 (N_15623,N_15369,N_15287);
or U15624 (N_15624,N_15255,N_15313);
nand U15625 (N_15625,N_15409,N_15321);
xnor U15626 (N_15626,N_15346,N_15368);
or U15627 (N_15627,N_15421,N_15408);
or U15628 (N_15628,N_15285,N_15261);
and U15629 (N_15629,N_15370,N_15420);
nand U15630 (N_15630,N_15479,N_15270);
and U15631 (N_15631,N_15444,N_15283);
and U15632 (N_15632,N_15489,N_15434);
and U15633 (N_15633,N_15463,N_15382);
xor U15634 (N_15634,N_15289,N_15423);
and U15635 (N_15635,N_15254,N_15429);
xor U15636 (N_15636,N_15265,N_15342);
nor U15637 (N_15637,N_15489,N_15450);
xnor U15638 (N_15638,N_15398,N_15408);
or U15639 (N_15639,N_15328,N_15450);
nand U15640 (N_15640,N_15428,N_15360);
nand U15641 (N_15641,N_15370,N_15347);
and U15642 (N_15642,N_15471,N_15349);
nor U15643 (N_15643,N_15449,N_15482);
xor U15644 (N_15644,N_15411,N_15417);
or U15645 (N_15645,N_15332,N_15486);
nand U15646 (N_15646,N_15485,N_15396);
nand U15647 (N_15647,N_15491,N_15349);
and U15648 (N_15648,N_15278,N_15312);
xnor U15649 (N_15649,N_15311,N_15338);
or U15650 (N_15650,N_15358,N_15480);
nand U15651 (N_15651,N_15359,N_15262);
and U15652 (N_15652,N_15364,N_15298);
nor U15653 (N_15653,N_15341,N_15390);
and U15654 (N_15654,N_15262,N_15263);
or U15655 (N_15655,N_15295,N_15353);
nor U15656 (N_15656,N_15407,N_15471);
nor U15657 (N_15657,N_15410,N_15349);
nand U15658 (N_15658,N_15309,N_15288);
and U15659 (N_15659,N_15308,N_15468);
xnor U15660 (N_15660,N_15447,N_15404);
nand U15661 (N_15661,N_15386,N_15331);
nand U15662 (N_15662,N_15363,N_15432);
or U15663 (N_15663,N_15404,N_15470);
xor U15664 (N_15664,N_15412,N_15349);
or U15665 (N_15665,N_15404,N_15323);
nand U15666 (N_15666,N_15419,N_15427);
nand U15667 (N_15667,N_15317,N_15432);
nand U15668 (N_15668,N_15388,N_15391);
or U15669 (N_15669,N_15291,N_15287);
nor U15670 (N_15670,N_15404,N_15460);
and U15671 (N_15671,N_15398,N_15273);
or U15672 (N_15672,N_15263,N_15497);
or U15673 (N_15673,N_15410,N_15266);
nor U15674 (N_15674,N_15391,N_15496);
or U15675 (N_15675,N_15477,N_15483);
or U15676 (N_15676,N_15477,N_15487);
xnor U15677 (N_15677,N_15299,N_15456);
nor U15678 (N_15678,N_15449,N_15257);
and U15679 (N_15679,N_15319,N_15454);
and U15680 (N_15680,N_15407,N_15493);
or U15681 (N_15681,N_15452,N_15356);
nor U15682 (N_15682,N_15254,N_15253);
or U15683 (N_15683,N_15432,N_15324);
nor U15684 (N_15684,N_15299,N_15430);
xnor U15685 (N_15685,N_15264,N_15409);
xnor U15686 (N_15686,N_15450,N_15279);
nand U15687 (N_15687,N_15393,N_15388);
nand U15688 (N_15688,N_15276,N_15497);
or U15689 (N_15689,N_15395,N_15458);
nor U15690 (N_15690,N_15424,N_15438);
nand U15691 (N_15691,N_15382,N_15364);
nor U15692 (N_15692,N_15478,N_15435);
and U15693 (N_15693,N_15293,N_15392);
nor U15694 (N_15694,N_15285,N_15477);
and U15695 (N_15695,N_15473,N_15264);
and U15696 (N_15696,N_15438,N_15459);
or U15697 (N_15697,N_15400,N_15272);
xnor U15698 (N_15698,N_15486,N_15451);
and U15699 (N_15699,N_15324,N_15298);
or U15700 (N_15700,N_15451,N_15460);
nand U15701 (N_15701,N_15294,N_15368);
nand U15702 (N_15702,N_15488,N_15264);
nor U15703 (N_15703,N_15346,N_15433);
xnor U15704 (N_15704,N_15498,N_15274);
or U15705 (N_15705,N_15349,N_15273);
or U15706 (N_15706,N_15495,N_15399);
and U15707 (N_15707,N_15355,N_15402);
nand U15708 (N_15708,N_15354,N_15369);
nor U15709 (N_15709,N_15397,N_15314);
or U15710 (N_15710,N_15443,N_15465);
nor U15711 (N_15711,N_15335,N_15358);
nor U15712 (N_15712,N_15485,N_15427);
nor U15713 (N_15713,N_15264,N_15302);
and U15714 (N_15714,N_15341,N_15263);
or U15715 (N_15715,N_15336,N_15495);
nor U15716 (N_15716,N_15446,N_15271);
nand U15717 (N_15717,N_15498,N_15447);
or U15718 (N_15718,N_15381,N_15312);
nand U15719 (N_15719,N_15339,N_15318);
nand U15720 (N_15720,N_15481,N_15377);
nor U15721 (N_15721,N_15496,N_15371);
xor U15722 (N_15722,N_15383,N_15416);
nor U15723 (N_15723,N_15289,N_15438);
nand U15724 (N_15724,N_15388,N_15386);
and U15725 (N_15725,N_15266,N_15250);
or U15726 (N_15726,N_15287,N_15427);
or U15727 (N_15727,N_15346,N_15410);
nand U15728 (N_15728,N_15322,N_15267);
or U15729 (N_15729,N_15383,N_15415);
or U15730 (N_15730,N_15441,N_15318);
and U15731 (N_15731,N_15475,N_15266);
and U15732 (N_15732,N_15421,N_15339);
xor U15733 (N_15733,N_15257,N_15389);
xor U15734 (N_15734,N_15276,N_15397);
nand U15735 (N_15735,N_15364,N_15449);
and U15736 (N_15736,N_15325,N_15459);
xor U15737 (N_15737,N_15467,N_15431);
xnor U15738 (N_15738,N_15336,N_15407);
nand U15739 (N_15739,N_15326,N_15313);
nor U15740 (N_15740,N_15427,N_15385);
nor U15741 (N_15741,N_15374,N_15470);
xnor U15742 (N_15742,N_15451,N_15346);
nor U15743 (N_15743,N_15486,N_15340);
and U15744 (N_15744,N_15498,N_15344);
nand U15745 (N_15745,N_15355,N_15373);
or U15746 (N_15746,N_15332,N_15415);
nand U15747 (N_15747,N_15445,N_15266);
xor U15748 (N_15748,N_15317,N_15273);
nand U15749 (N_15749,N_15489,N_15488);
nand U15750 (N_15750,N_15694,N_15566);
and U15751 (N_15751,N_15710,N_15583);
and U15752 (N_15752,N_15728,N_15607);
or U15753 (N_15753,N_15556,N_15727);
and U15754 (N_15754,N_15595,N_15513);
nor U15755 (N_15755,N_15729,N_15636);
nand U15756 (N_15756,N_15613,N_15514);
nor U15757 (N_15757,N_15647,N_15702);
xor U15758 (N_15758,N_15604,N_15601);
or U15759 (N_15759,N_15718,N_15635);
and U15760 (N_15760,N_15697,N_15691);
nor U15761 (N_15761,N_15650,N_15708);
nand U15762 (N_15762,N_15540,N_15505);
and U15763 (N_15763,N_15734,N_15696);
and U15764 (N_15764,N_15700,N_15609);
and U15765 (N_15765,N_15543,N_15677);
xnor U15766 (N_15766,N_15510,N_15568);
xnor U15767 (N_15767,N_15532,N_15633);
xor U15768 (N_15768,N_15588,N_15507);
xor U15769 (N_15769,N_15640,N_15748);
nor U15770 (N_15770,N_15567,N_15648);
nand U15771 (N_15771,N_15564,N_15531);
or U15772 (N_15772,N_15693,N_15602);
xnor U15773 (N_15773,N_15544,N_15587);
nand U15774 (N_15774,N_15589,N_15664);
xor U15775 (N_15775,N_15547,N_15713);
nand U15776 (N_15776,N_15711,N_15598);
nor U15777 (N_15777,N_15606,N_15652);
nand U15778 (N_15778,N_15577,N_15662);
nand U15779 (N_15779,N_15715,N_15709);
xnor U15780 (N_15780,N_15525,N_15580);
xor U15781 (N_15781,N_15743,N_15590);
xnor U15782 (N_15782,N_15665,N_15659);
nand U15783 (N_15783,N_15611,N_15625);
xnor U15784 (N_15784,N_15720,N_15667);
nand U15785 (N_15785,N_15546,N_15703);
or U15786 (N_15786,N_15627,N_15533);
xnor U15787 (N_15787,N_15511,N_15725);
xnor U15788 (N_15788,N_15653,N_15615);
and U15789 (N_15789,N_15554,N_15585);
or U15790 (N_15790,N_15529,N_15535);
nor U15791 (N_15791,N_15731,N_15733);
xnor U15792 (N_15792,N_15634,N_15736);
and U15793 (N_15793,N_15534,N_15501);
xor U15794 (N_15794,N_15737,N_15658);
and U15795 (N_15795,N_15669,N_15698);
nor U15796 (N_15796,N_15572,N_15545);
and U15797 (N_15797,N_15742,N_15624);
xnor U15798 (N_15798,N_15536,N_15539);
xnor U15799 (N_15799,N_15555,N_15631);
nor U15800 (N_15800,N_15746,N_15724);
nor U15801 (N_15801,N_15643,N_15628);
xor U15802 (N_15802,N_15672,N_15557);
nor U15803 (N_15803,N_15522,N_15674);
or U15804 (N_15804,N_15684,N_15586);
nand U15805 (N_15805,N_15508,N_15654);
or U15806 (N_15806,N_15623,N_15550);
or U15807 (N_15807,N_15560,N_15706);
nor U15808 (N_15808,N_15503,N_15578);
nor U15809 (N_15809,N_15518,N_15569);
and U15810 (N_15810,N_15579,N_15553);
nand U15811 (N_15811,N_15515,N_15558);
nor U15812 (N_15812,N_15681,N_15668);
or U15813 (N_15813,N_15597,N_15745);
nor U15814 (N_15814,N_15638,N_15626);
nand U15815 (N_15815,N_15678,N_15670);
xor U15816 (N_15816,N_15632,N_15732);
and U15817 (N_15817,N_15639,N_15721);
or U15818 (N_15818,N_15740,N_15646);
and U15819 (N_15819,N_15500,N_15517);
xor U15820 (N_15820,N_15530,N_15679);
or U15821 (N_15821,N_15663,N_15594);
or U15822 (N_15822,N_15584,N_15712);
xor U15823 (N_15823,N_15645,N_15656);
nor U15824 (N_15824,N_15561,N_15600);
and U15825 (N_15825,N_15707,N_15739);
nand U15826 (N_15826,N_15621,N_15749);
and U15827 (N_15827,N_15570,N_15747);
nor U15828 (N_15828,N_15608,N_15717);
nor U15829 (N_15829,N_15661,N_15673);
nor U15830 (N_15830,N_15719,N_15573);
or U15831 (N_15831,N_15520,N_15537);
nor U15832 (N_15832,N_15575,N_15692);
or U15833 (N_15833,N_15565,N_15683);
or U15834 (N_15834,N_15716,N_15622);
or U15835 (N_15835,N_15552,N_15576);
or U15836 (N_15836,N_15704,N_15741);
xor U15837 (N_15837,N_15689,N_15548);
or U15838 (N_15838,N_15680,N_15549);
or U15839 (N_15839,N_15571,N_15651);
nand U15840 (N_15840,N_15574,N_15562);
and U15841 (N_15841,N_15605,N_15541);
xnor U15842 (N_15842,N_15642,N_15676);
xor U15843 (N_15843,N_15730,N_15701);
and U15844 (N_15844,N_15649,N_15516);
nor U15845 (N_15845,N_15699,N_15523);
xor U15846 (N_15846,N_15528,N_15592);
xnor U15847 (N_15847,N_15591,N_15685);
nand U15848 (N_15848,N_15524,N_15690);
xnor U15849 (N_15849,N_15512,N_15705);
and U15850 (N_15850,N_15596,N_15506);
nand U15851 (N_15851,N_15687,N_15660);
and U15852 (N_15852,N_15619,N_15675);
or U15853 (N_15853,N_15644,N_15502);
and U15854 (N_15854,N_15582,N_15526);
nand U15855 (N_15855,N_15738,N_15612);
xor U15856 (N_15856,N_15695,N_15735);
nand U15857 (N_15857,N_15630,N_15614);
nor U15858 (N_15858,N_15599,N_15542);
xnor U15859 (N_15859,N_15519,N_15714);
nor U15860 (N_15860,N_15657,N_15618);
nand U15861 (N_15861,N_15610,N_15688);
nor U15862 (N_15862,N_15538,N_15726);
or U15863 (N_15863,N_15686,N_15616);
nor U15864 (N_15864,N_15744,N_15603);
and U15865 (N_15865,N_15722,N_15581);
nand U15866 (N_15866,N_15655,N_15551);
xor U15867 (N_15867,N_15682,N_15559);
nor U15868 (N_15868,N_15617,N_15723);
nor U15869 (N_15869,N_15504,N_15671);
nand U15870 (N_15870,N_15629,N_15593);
nand U15871 (N_15871,N_15509,N_15637);
nor U15872 (N_15872,N_15620,N_15641);
and U15873 (N_15873,N_15527,N_15666);
nand U15874 (N_15874,N_15563,N_15521);
or U15875 (N_15875,N_15572,N_15742);
nand U15876 (N_15876,N_15600,N_15691);
nand U15877 (N_15877,N_15749,N_15518);
and U15878 (N_15878,N_15662,N_15665);
xor U15879 (N_15879,N_15522,N_15708);
and U15880 (N_15880,N_15548,N_15649);
and U15881 (N_15881,N_15521,N_15585);
and U15882 (N_15882,N_15696,N_15534);
and U15883 (N_15883,N_15538,N_15718);
nor U15884 (N_15884,N_15595,N_15748);
nand U15885 (N_15885,N_15618,N_15632);
or U15886 (N_15886,N_15716,N_15593);
or U15887 (N_15887,N_15615,N_15630);
nor U15888 (N_15888,N_15576,N_15503);
or U15889 (N_15889,N_15612,N_15529);
nand U15890 (N_15890,N_15685,N_15571);
or U15891 (N_15891,N_15571,N_15509);
nor U15892 (N_15892,N_15641,N_15706);
nor U15893 (N_15893,N_15675,N_15615);
or U15894 (N_15894,N_15500,N_15666);
xnor U15895 (N_15895,N_15505,N_15703);
nand U15896 (N_15896,N_15556,N_15532);
and U15897 (N_15897,N_15574,N_15616);
nor U15898 (N_15898,N_15671,N_15605);
and U15899 (N_15899,N_15687,N_15696);
nor U15900 (N_15900,N_15568,N_15654);
xnor U15901 (N_15901,N_15585,N_15689);
xnor U15902 (N_15902,N_15561,N_15552);
and U15903 (N_15903,N_15712,N_15664);
or U15904 (N_15904,N_15677,N_15634);
nor U15905 (N_15905,N_15635,N_15645);
or U15906 (N_15906,N_15583,N_15674);
nor U15907 (N_15907,N_15564,N_15502);
nor U15908 (N_15908,N_15608,N_15632);
or U15909 (N_15909,N_15713,N_15666);
and U15910 (N_15910,N_15711,N_15629);
nand U15911 (N_15911,N_15550,N_15585);
and U15912 (N_15912,N_15687,N_15718);
nand U15913 (N_15913,N_15639,N_15731);
xnor U15914 (N_15914,N_15506,N_15553);
xor U15915 (N_15915,N_15648,N_15507);
xor U15916 (N_15916,N_15540,N_15593);
xnor U15917 (N_15917,N_15720,N_15575);
nor U15918 (N_15918,N_15742,N_15520);
or U15919 (N_15919,N_15619,N_15652);
nor U15920 (N_15920,N_15520,N_15626);
or U15921 (N_15921,N_15600,N_15718);
nor U15922 (N_15922,N_15523,N_15737);
xnor U15923 (N_15923,N_15679,N_15548);
and U15924 (N_15924,N_15525,N_15621);
and U15925 (N_15925,N_15572,N_15675);
nor U15926 (N_15926,N_15579,N_15511);
xor U15927 (N_15927,N_15663,N_15514);
or U15928 (N_15928,N_15666,N_15528);
xnor U15929 (N_15929,N_15693,N_15580);
nor U15930 (N_15930,N_15742,N_15677);
nor U15931 (N_15931,N_15669,N_15521);
or U15932 (N_15932,N_15613,N_15560);
nor U15933 (N_15933,N_15531,N_15510);
or U15934 (N_15934,N_15589,N_15689);
or U15935 (N_15935,N_15683,N_15555);
and U15936 (N_15936,N_15534,N_15551);
and U15937 (N_15937,N_15596,N_15526);
and U15938 (N_15938,N_15604,N_15585);
or U15939 (N_15939,N_15651,N_15589);
or U15940 (N_15940,N_15631,N_15667);
nor U15941 (N_15941,N_15699,N_15620);
xnor U15942 (N_15942,N_15558,N_15503);
nor U15943 (N_15943,N_15704,N_15681);
and U15944 (N_15944,N_15556,N_15627);
nor U15945 (N_15945,N_15724,N_15625);
xor U15946 (N_15946,N_15537,N_15689);
xnor U15947 (N_15947,N_15603,N_15504);
or U15948 (N_15948,N_15542,N_15627);
xor U15949 (N_15949,N_15517,N_15650);
nand U15950 (N_15950,N_15567,N_15741);
and U15951 (N_15951,N_15615,N_15621);
and U15952 (N_15952,N_15718,N_15720);
xor U15953 (N_15953,N_15592,N_15651);
nor U15954 (N_15954,N_15612,N_15585);
xnor U15955 (N_15955,N_15586,N_15582);
and U15956 (N_15956,N_15547,N_15513);
nand U15957 (N_15957,N_15519,N_15566);
xnor U15958 (N_15958,N_15651,N_15727);
and U15959 (N_15959,N_15641,N_15696);
nor U15960 (N_15960,N_15578,N_15652);
nand U15961 (N_15961,N_15530,N_15708);
xnor U15962 (N_15962,N_15692,N_15718);
and U15963 (N_15963,N_15692,N_15568);
nor U15964 (N_15964,N_15644,N_15598);
nand U15965 (N_15965,N_15723,N_15536);
nor U15966 (N_15966,N_15576,N_15531);
xnor U15967 (N_15967,N_15569,N_15586);
or U15968 (N_15968,N_15609,N_15644);
nand U15969 (N_15969,N_15739,N_15616);
and U15970 (N_15970,N_15644,N_15650);
and U15971 (N_15971,N_15617,N_15741);
or U15972 (N_15972,N_15595,N_15697);
and U15973 (N_15973,N_15514,N_15577);
nor U15974 (N_15974,N_15640,N_15702);
xnor U15975 (N_15975,N_15574,N_15687);
nor U15976 (N_15976,N_15696,N_15714);
and U15977 (N_15977,N_15599,N_15576);
or U15978 (N_15978,N_15651,N_15516);
nor U15979 (N_15979,N_15673,N_15749);
nand U15980 (N_15980,N_15522,N_15679);
nand U15981 (N_15981,N_15643,N_15734);
nand U15982 (N_15982,N_15612,N_15550);
and U15983 (N_15983,N_15619,N_15718);
nand U15984 (N_15984,N_15617,N_15501);
nor U15985 (N_15985,N_15689,N_15609);
or U15986 (N_15986,N_15686,N_15712);
and U15987 (N_15987,N_15632,N_15726);
xor U15988 (N_15988,N_15644,N_15568);
or U15989 (N_15989,N_15601,N_15721);
nor U15990 (N_15990,N_15551,N_15746);
and U15991 (N_15991,N_15728,N_15561);
or U15992 (N_15992,N_15715,N_15722);
xor U15993 (N_15993,N_15725,N_15503);
nand U15994 (N_15994,N_15741,N_15649);
nand U15995 (N_15995,N_15720,N_15530);
or U15996 (N_15996,N_15658,N_15514);
nand U15997 (N_15997,N_15571,N_15708);
xnor U15998 (N_15998,N_15561,N_15719);
xor U15999 (N_15999,N_15617,N_15704);
nand U16000 (N_16000,N_15945,N_15843);
nor U16001 (N_16001,N_15977,N_15781);
nor U16002 (N_16002,N_15866,N_15988);
xnor U16003 (N_16003,N_15833,N_15954);
and U16004 (N_16004,N_15853,N_15935);
nor U16005 (N_16005,N_15993,N_15881);
nor U16006 (N_16006,N_15985,N_15760);
nor U16007 (N_16007,N_15793,N_15766);
or U16008 (N_16008,N_15816,N_15914);
and U16009 (N_16009,N_15778,N_15824);
and U16010 (N_16010,N_15911,N_15888);
nand U16011 (N_16011,N_15909,N_15956);
or U16012 (N_16012,N_15927,N_15856);
nand U16013 (N_16013,N_15846,N_15889);
nand U16014 (N_16014,N_15883,N_15862);
nor U16015 (N_16015,N_15942,N_15970);
and U16016 (N_16016,N_15929,N_15763);
nor U16017 (N_16017,N_15978,N_15857);
nor U16018 (N_16018,N_15772,N_15795);
xnor U16019 (N_16019,N_15870,N_15844);
and U16020 (N_16020,N_15940,N_15799);
nand U16021 (N_16021,N_15976,N_15769);
nand U16022 (N_16022,N_15765,N_15959);
and U16023 (N_16023,N_15801,N_15958);
nand U16024 (N_16024,N_15851,N_15926);
and U16025 (N_16025,N_15949,N_15854);
or U16026 (N_16026,N_15823,N_15786);
xnor U16027 (N_16027,N_15810,N_15832);
and U16028 (N_16028,N_15775,N_15903);
nand U16029 (N_16029,N_15828,N_15934);
or U16030 (N_16030,N_15966,N_15754);
nor U16031 (N_16031,N_15753,N_15867);
and U16032 (N_16032,N_15868,N_15879);
and U16033 (N_16033,N_15841,N_15916);
or U16034 (N_16034,N_15905,N_15825);
nand U16035 (N_16035,N_15807,N_15834);
or U16036 (N_16036,N_15939,N_15917);
or U16037 (N_16037,N_15776,N_15974);
xnor U16038 (N_16038,N_15971,N_15839);
nand U16039 (N_16039,N_15811,N_15864);
xor U16040 (N_16040,N_15931,N_15751);
nor U16041 (N_16041,N_15941,N_15882);
xor U16042 (N_16042,N_15968,N_15890);
or U16043 (N_16043,N_15863,N_15980);
xnor U16044 (N_16044,N_15947,N_15830);
and U16045 (N_16045,N_15814,N_15913);
nor U16046 (N_16046,N_15805,N_15933);
xor U16047 (N_16047,N_15788,N_15948);
nor U16048 (N_16048,N_15878,N_15928);
nor U16049 (N_16049,N_15922,N_15984);
nor U16050 (N_16050,N_15898,N_15899);
nand U16051 (N_16051,N_15983,N_15806);
and U16052 (N_16052,N_15923,N_15831);
nor U16053 (N_16053,N_15845,N_15908);
nand U16054 (N_16054,N_15904,N_15794);
and U16055 (N_16055,N_15758,N_15755);
or U16056 (N_16056,N_15887,N_15975);
or U16057 (N_16057,N_15798,N_15787);
xnor U16058 (N_16058,N_15907,N_15943);
nor U16059 (N_16059,N_15797,N_15919);
nand U16060 (N_16060,N_15790,N_15885);
nor U16061 (N_16061,N_15906,N_15809);
or U16062 (N_16062,N_15821,N_15803);
and U16063 (N_16063,N_15930,N_15802);
and U16064 (N_16064,N_15981,N_15871);
nor U16065 (N_16065,N_15872,N_15915);
nor U16066 (N_16066,N_15835,N_15989);
nor U16067 (N_16067,N_15876,N_15759);
or U16068 (N_16068,N_15900,N_15994);
or U16069 (N_16069,N_15952,N_15842);
nor U16070 (N_16070,N_15895,N_15991);
nor U16071 (N_16071,N_15986,N_15955);
and U16072 (N_16072,N_15762,N_15998);
nand U16073 (N_16073,N_15858,N_15861);
and U16074 (N_16074,N_15827,N_15865);
or U16075 (N_16075,N_15946,N_15838);
and U16076 (N_16076,N_15757,N_15804);
nor U16077 (N_16077,N_15783,N_15964);
or U16078 (N_16078,N_15820,N_15785);
or U16079 (N_16079,N_15829,N_15789);
and U16080 (N_16080,N_15819,N_15996);
xor U16081 (N_16081,N_15936,N_15910);
or U16082 (N_16082,N_15997,N_15893);
and U16083 (N_16083,N_15850,N_15847);
nor U16084 (N_16084,N_15951,N_15880);
and U16085 (N_16085,N_15920,N_15950);
xnor U16086 (N_16086,N_15771,N_15875);
xor U16087 (N_16087,N_15937,N_15869);
nor U16088 (N_16088,N_15884,N_15896);
xnor U16089 (N_16089,N_15967,N_15808);
nor U16090 (N_16090,N_15918,N_15902);
and U16091 (N_16091,N_15770,N_15992);
xor U16092 (N_16092,N_15960,N_15874);
xnor U16093 (N_16093,N_15768,N_15873);
nor U16094 (N_16094,N_15855,N_15773);
xor U16095 (N_16095,N_15953,N_15921);
nor U16096 (N_16096,N_15990,N_15812);
and U16097 (N_16097,N_15979,N_15774);
nor U16098 (N_16098,N_15796,N_15784);
xor U16099 (N_16099,N_15901,N_15892);
xnor U16100 (N_16100,N_15836,N_15779);
and U16101 (N_16101,N_15782,N_15818);
nand U16102 (N_16102,N_15891,N_15963);
and U16103 (N_16103,N_15969,N_15860);
xnor U16104 (N_16104,N_15924,N_15886);
and U16105 (N_16105,N_15944,N_15792);
nand U16106 (N_16106,N_15826,N_15800);
or U16107 (N_16107,N_15813,N_15925);
or U16108 (N_16108,N_15780,N_15972);
nand U16109 (N_16109,N_15877,N_15965);
or U16110 (N_16110,N_15962,N_15761);
or U16111 (N_16111,N_15764,N_15837);
xor U16112 (N_16112,N_15938,N_15750);
or U16113 (N_16113,N_15973,N_15995);
or U16114 (N_16114,N_15822,N_15894);
nand U16115 (N_16115,N_15767,N_15897);
xnor U16116 (N_16116,N_15999,N_15957);
nor U16117 (N_16117,N_15756,N_15912);
or U16118 (N_16118,N_15815,N_15859);
or U16119 (N_16119,N_15791,N_15848);
or U16120 (N_16120,N_15777,N_15987);
xnor U16121 (N_16121,N_15817,N_15982);
and U16122 (N_16122,N_15852,N_15849);
nor U16123 (N_16123,N_15752,N_15840);
or U16124 (N_16124,N_15961,N_15932);
or U16125 (N_16125,N_15779,N_15803);
nor U16126 (N_16126,N_15993,N_15944);
nand U16127 (N_16127,N_15847,N_15764);
nand U16128 (N_16128,N_15993,N_15802);
and U16129 (N_16129,N_15972,N_15868);
nor U16130 (N_16130,N_15982,N_15877);
and U16131 (N_16131,N_15868,N_15978);
xor U16132 (N_16132,N_15821,N_15980);
or U16133 (N_16133,N_15902,N_15885);
nor U16134 (N_16134,N_15838,N_15845);
nand U16135 (N_16135,N_15980,N_15948);
nor U16136 (N_16136,N_15997,N_15847);
and U16137 (N_16137,N_15950,N_15907);
nand U16138 (N_16138,N_15993,N_15780);
nor U16139 (N_16139,N_15919,N_15849);
nand U16140 (N_16140,N_15775,N_15822);
or U16141 (N_16141,N_15995,N_15781);
nor U16142 (N_16142,N_15789,N_15951);
xor U16143 (N_16143,N_15876,N_15817);
nor U16144 (N_16144,N_15863,N_15911);
xor U16145 (N_16145,N_15992,N_15875);
or U16146 (N_16146,N_15773,N_15876);
xnor U16147 (N_16147,N_15803,N_15828);
nor U16148 (N_16148,N_15836,N_15766);
nor U16149 (N_16149,N_15965,N_15947);
nor U16150 (N_16150,N_15881,N_15947);
nand U16151 (N_16151,N_15756,N_15963);
nand U16152 (N_16152,N_15943,N_15900);
or U16153 (N_16153,N_15847,N_15751);
and U16154 (N_16154,N_15889,N_15892);
or U16155 (N_16155,N_15833,N_15953);
xnor U16156 (N_16156,N_15916,N_15919);
xor U16157 (N_16157,N_15785,N_15827);
nor U16158 (N_16158,N_15983,N_15977);
xnor U16159 (N_16159,N_15947,N_15902);
nand U16160 (N_16160,N_15875,N_15905);
and U16161 (N_16161,N_15874,N_15843);
nor U16162 (N_16162,N_15968,N_15762);
or U16163 (N_16163,N_15883,N_15821);
nand U16164 (N_16164,N_15831,N_15848);
xor U16165 (N_16165,N_15937,N_15944);
and U16166 (N_16166,N_15862,N_15795);
xor U16167 (N_16167,N_15889,N_15756);
or U16168 (N_16168,N_15836,N_15769);
nand U16169 (N_16169,N_15781,N_15757);
and U16170 (N_16170,N_15956,N_15922);
nor U16171 (N_16171,N_15890,N_15912);
xor U16172 (N_16172,N_15982,N_15816);
xnor U16173 (N_16173,N_15825,N_15923);
nand U16174 (N_16174,N_15997,N_15947);
and U16175 (N_16175,N_15810,N_15949);
and U16176 (N_16176,N_15973,N_15787);
nand U16177 (N_16177,N_15765,N_15892);
and U16178 (N_16178,N_15883,N_15786);
nor U16179 (N_16179,N_15811,N_15907);
or U16180 (N_16180,N_15793,N_15915);
and U16181 (N_16181,N_15940,N_15833);
nand U16182 (N_16182,N_15874,N_15791);
nand U16183 (N_16183,N_15874,N_15810);
xor U16184 (N_16184,N_15805,N_15958);
nand U16185 (N_16185,N_15910,N_15828);
or U16186 (N_16186,N_15800,N_15908);
nand U16187 (N_16187,N_15800,N_15953);
xnor U16188 (N_16188,N_15755,N_15887);
or U16189 (N_16189,N_15806,N_15877);
and U16190 (N_16190,N_15838,N_15868);
xor U16191 (N_16191,N_15898,N_15865);
nand U16192 (N_16192,N_15982,N_15967);
nand U16193 (N_16193,N_15883,N_15866);
or U16194 (N_16194,N_15896,N_15777);
or U16195 (N_16195,N_15780,N_15798);
and U16196 (N_16196,N_15751,N_15775);
xor U16197 (N_16197,N_15751,N_15838);
and U16198 (N_16198,N_15868,N_15903);
or U16199 (N_16199,N_15982,N_15912);
nor U16200 (N_16200,N_15829,N_15940);
or U16201 (N_16201,N_15869,N_15782);
or U16202 (N_16202,N_15967,N_15919);
xnor U16203 (N_16203,N_15935,N_15798);
xor U16204 (N_16204,N_15974,N_15801);
and U16205 (N_16205,N_15917,N_15991);
xnor U16206 (N_16206,N_15909,N_15779);
xor U16207 (N_16207,N_15772,N_15901);
nor U16208 (N_16208,N_15811,N_15852);
or U16209 (N_16209,N_15827,N_15825);
and U16210 (N_16210,N_15917,N_15892);
or U16211 (N_16211,N_15938,N_15857);
nor U16212 (N_16212,N_15803,N_15888);
nand U16213 (N_16213,N_15802,N_15865);
nand U16214 (N_16214,N_15958,N_15955);
and U16215 (N_16215,N_15913,N_15771);
nand U16216 (N_16216,N_15997,N_15925);
xor U16217 (N_16217,N_15859,N_15890);
xor U16218 (N_16218,N_15897,N_15913);
and U16219 (N_16219,N_15820,N_15812);
nand U16220 (N_16220,N_15987,N_15770);
nor U16221 (N_16221,N_15835,N_15787);
nand U16222 (N_16222,N_15925,N_15975);
nand U16223 (N_16223,N_15843,N_15834);
xnor U16224 (N_16224,N_15923,N_15790);
or U16225 (N_16225,N_15869,N_15935);
nor U16226 (N_16226,N_15778,N_15750);
or U16227 (N_16227,N_15953,N_15827);
nand U16228 (N_16228,N_15786,N_15920);
xor U16229 (N_16229,N_15891,N_15777);
or U16230 (N_16230,N_15981,N_15874);
nand U16231 (N_16231,N_15753,N_15964);
nor U16232 (N_16232,N_15836,N_15750);
xor U16233 (N_16233,N_15866,N_15909);
nor U16234 (N_16234,N_15872,N_15951);
or U16235 (N_16235,N_15991,N_15816);
xnor U16236 (N_16236,N_15811,N_15767);
nor U16237 (N_16237,N_15994,N_15997);
nand U16238 (N_16238,N_15948,N_15919);
xor U16239 (N_16239,N_15835,N_15890);
xor U16240 (N_16240,N_15771,N_15898);
nor U16241 (N_16241,N_15786,N_15827);
xor U16242 (N_16242,N_15814,N_15846);
nor U16243 (N_16243,N_15963,N_15765);
and U16244 (N_16244,N_15808,N_15906);
xor U16245 (N_16245,N_15765,N_15954);
nor U16246 (N_16246,N_15761,N_15791);
or U16247 (N_16247,N_15913,N_15783);
or U16248 (N_16248,N_15889,N_15869);
xnor U16249 (N_16249,N_15987,N_15882);
nand U16250 (N_16250,N_16166,N_16097);
and U16251 (N_16251,N_16093,N_16018);
nor U16252 (N_16252,N_16228,N_16116);
nand U16253 (N_16253,N_16025,N_16057);
nand U16254 (N_16254,N_16085,N_16130);
or U16255 (N_16255,N_16182,N_16139);
xor U16256 (N_16256,N_16033,N_16245);
nor U16257 (N_16257,N_16092,N_16168);
xnor U16258 (N_16258,N_16239,N_16240);
nand U16259 (N_16259,N_16035,N_16193);
and U16260 (N_16260,N_16249,N_16223);
and U16261 (N_16261,N_16089,N_16060);
or U16262 (N_16262,N_16099,N_16062);
nor U16263 (N_16263,N_16069,N_16129);
nor U16264 (N_16264,N_16019,N_16244);
xor U16265 (N_16265,N_16241,N_16145);
nor U16266 (N_16266,N_16225,N_16013);
or U16267 (N_16267,N_16140,N_16045);
nand U16268 (N_16268,N_16243,N_16242);
xnor U16269 (N_16269,N_16084,N_16103);
and U16270 (N_16270,N_16164,N_16210);
nor U16271 (N_16271,N_16006,N_16142);
and U16272 (N_16272,N_16088,N_16022);
nor U16273 (N_16273,N_16004,N_16180);
nand U16274 (N_16274,N_16217,N_16010);
nand U16275 (N_16275,N_16221,N_16199);
or U16276 (N_16276,N_16232,N_16151);
or U16277 (N_16277,N_16065,N_16152);
and U16278 (N_16278,N_16190,N_16165);
nand U16279 (N_16279,N_16247,N_16061);
or U16280 (N_16280,N_16195,N_16076);
or U16281 (N_16281,N_16183,N_16012);
nor U16282 (N_16282,N_16162,N_16067);
xnor U16283 (N_16283,N_16222,N_16203);
and U16284 (N_16284,N_16023,N_16185);
or U16285 (N_16285,N_16172,N_16169);
nor U16286 (N_16286,N_16079,N_16021);
nand U16287 (N_16287,N_16095,N_16024);
and U16288 (N_16288,N_16214,N_16136);
nand U16289 (N_16289,N_16248,N_16051);
or U16290 (N_16290,N_16147,N_16118);
nor U16291 (N_16291,N_16167,N_16213);
xnor U16292 (N_16292,N_16011,N_16090);
or U16293 (N_16293,N_16111,N_16120);
nand U16294 (N_16294,N_16078,N_16072);
nor U16295 (N_16295,N_16037,N_16144);
or U16296 (N_16296,N_16132,N_16154);
or U16297 (N_16297,N_16157,N_16071);
xor U16298 (N_16298,N_16191,N_16075);
or U16299 (N_16299,N_16224,N_16115);
xor U16300 (N_16300,N_16209,N_16208);
xnor U16301 (N_16301,N_16114,N_16187);
or U16302 (N_16302,N_16015,N_16211);
nand U16303 (N_16303,N_16204,N_16094);
nand U16304 (N_16304,N_16124,N_16073);
and U16305 (N_16305,N_16083,N_16031);
and U16306 (N_16306,N_16104,N_16181);
nor U16307 (N_16307,N_16007,N_16036);
or U16308 (N_16308,N_16212,N_16246);
nand U16309 (N_16309,N_16163,N_16016);
xor U16310 (N_16310,N_16029,N_16039);
and U16311 (N_16311,N_16091,N_16158);
or U16312 (N_16312,N_16200,N_16231);
nand U16313 (N_16313,N_16175,N_16000);
nor U16314 (N_16314,N_16137,N_16192);
xor U16315 (N_16315,N_16082,N_16066);
nand U16316 (N_16316,N_16096,N_16063);
xor U16317 (N_16317,N_16236,N_16017);
or U16318 (N_16318,N_16048,N_16008);
nor U16319 (N_16319,N_16178,N_16184);
nand U16320 (N_16320,N_16227,N_16146);
and U16321 (N_16321,N_16064,N_16068);
nor U16322 (N_16322,N_16171,N_16127);
and U16323 (N_16323,N_16027,N_16206);
or U16324 (N_16324,N_16102,N_16216);
and U16325 (N_16325,N_16028,N_16100);
and U16326 (N_16326,N_16050,N_16009);
nor U16327 (N_16327,N_16081,N_16109);
or U16328 (N_16328,N_16198,N_16189);
and U16329 (N_16329,N_16044,N_16135);
nand U16330 (N_16330,N_16014,N_16156);
or U16331 (N_16331,N_16149,N_16001);
or U16332 (N_16332,N_16002,N_16020);
xor U16333 (N_16333,N_16119,N_16196);
nor U16334 (N_16334,N_16141,N_16155);
or U16335 (N_16335,N_16070,N_16122);
xor U16336 (N_16336,N_16026,N_16042);
nor U16337 (N_16337,N_16047,N_16230);
and U16338 (N_16338,N_16143,N_16107);
or U16339 (N_16339,N_16220,N_16188);
nor U16340 (N_16340,N_16153,N_16056);
or U16341 (N_16341,N_16179,N_16113);
nand U16342 (N_16342,N_16054,N_16098);
or U16343 (N_16343,N_16205,N_16229);
nor U16344 (N_16344,N_16032,N_16074);
nor U16345 (N_16345,N_16034,N_16218);
nor U16346 (N_16346,N_16197,N_16219);
nand U16347 (N_16347,N_16125,N_16117);
or U16348 (N_16348,N_16128,N_16207);
and U16349 (N_16349,N_16101,N_16170);
xor U16350 (N_16350,N_16133,N_16202);
or U16351 (N_16351,N_16043,N_16159);
nand U16352 (N_16352,N_16138,N_16052);
or U16353 (N_16353,N_16053,N_16005);
or U16354 (N_16354,N_16040,N_16134);
nor U16355 (N_16355,N_16112,N_16237);
and U16356 (N_16356,N_16150,N_16087);
xor U16357 (N_16357,N_16123,N_16058);
nand U16358 (N_16358,N_16086,N_16126);
or U16359 (N_16359,N_16046,N_16201);
or U16360 (N_16360,N_16055,N_16106);
and U16361 (N_16361,N_16186,N_16234);
nand U16362 (N_16362,N_16238,N_16059);
nor U16363 (N_16363,N_16131,N_16003);
and U16364 (N_16364,N_16160,N_16049);
nor U16365 (N_16365,N_16173,N_16215);
and U16366 (N_16366,N_16194,N_16110);
or U16367 (N_16367,N_16177,N_16108);
or U16368 (N_16368,N_16161,N_16148);
nand U16369 (N_16369,N_16121,N_16080);
and U16370 (N_16370,N_16233,N_16038);
nor U16371 (N_16371,N_16235,N_16105);
nand U16372 (N_16372,N_16226,N_16174);
and U16373 (N_16373,N_16077,N_16030);
xnor U16374 (N_16374,N_16176,N_16041);
or U16375 (N_16375,N_16026,N_16034);
or U16376 (N_16376,N_16223,N_16113);
or U16377 (N_16377,N_16027,N_16214);
nand U16378 (N_16378,N_16238,N_16239);
nor U16379 (N_16379,N_16243,N_16092);
nand U16380 (N_16380,N_16239,N_16231);
and U16381 (N_16381,N_16127,N_16186);
nor U16382 (N_16382,N_16178,N_16230);
or U16383 (N_16383,N_16163,N_16060);
or U16384 (N_16384,N_16013,N_16031);
or U16385 (N_16385,N_16233,N_16006);
or U16386 (N_16386,N_16216,N_16215);
and U16387 (N_16387,N_16131,N_16241);
nand U16388 (N_16388,N_16179,N_16097);
xnor U16389 (N_16389,N_16143,N_16041);
xnor U16390 (N_16390,N_16083,N_16212);
nand U16391 (N_16391,N_16087,N_16064);
and U16392 (N_16392,N_16062,N_16142);
or U16393 (N_16393,N_16015,N_16173);
nand U16394 (N_16394,N_16083,N_16241);
and U16395 (N_16395,N_16164,N_16064);
nor U16396 (N_16396,N_16245,N_16133);
nor U16397 (N_16397,N_16192,N_16158);
and U16398 (N_16398,N_16228,N_16122);
or U16399 (N_16399,N_16150,N_16097);
or U16400 (N_16400,N_16227,N_16210);
xor U16401 (N_16401,N_16097,N_16019);
or U16402 (N_16402,N_16066,N_16065);
nand U16403 (N_16403,N_16143,N_16204);
xor U16404 (N_16404,N_16124,N_16149);
and U16405 (N_16405,N_16174,N_16165);
xnor U16406 (N_16406,N_16053,N_16057);
and U16407 (N_16407,N_16133,N_16239);
nand U16408 (N_16408,N_16219,N_16193);
nand U16409 (N_16409,N_16176,N_16096);
or U16410 (N_16410,N_16249,N_16056);
xor U16411 (N_16411,N_16157,N_16011);
nand U16412 (N_16412,N_16132,N_16135);
xor U16413 (N_16413,N_16132,N_16169);
nand U16414 (N_16414,N_16015,N_16135);
and U16415 (N_16415,N_16046,N_16123);
nand U16416 (N_16416,N_16212,N_16150);
xnor U16417 (N_16417,N_16197,N_16120);
or U16418 (N_16418,N_16140,N_16241);
nor U16419 (N_16419,N_16132,N_16044);
nand U16420 (N_16420,N_16168,N_16239);
nor U16421 (N_16421,N_16092,N_16050);
and U16422 (N_16422,N_16199,N_16198);
nand U16423 (N_16423,N_16020,N_16047);
or U16424 (N_16424,N_16249,N_16188);
nor U16425 (N_16425,N_16153,N_16162);
and U16426 (N_16426,N_16246,N_16035);
xnor U16427 (N_16427,N_16106,N_16240);
and U16428 (N_16428,N_16065,N_16238);
xnor U16429 (N_16429,N_16229,N_16240);
xor U16430 (N_16430,N_16190,N_16221);
nor U16431 (N_16431,N_16098,N_16168);
or U16432 (N_16432,N_16128,N_16028);
xor U16433 (N_16433,N_16033,N_16048);
nor U16434 (N_16434,N_16176,N_16224);
nor U16435 (N_16435,N_16117,N_16233);
and U16436 (N_16436,N_16068,N_16214);
nor U16437 (N_16437,N_16108,N_16101);
nand U16438 (N_16438,N_16031,N_16103);
and U16439 (N_16439,N_16000,N_16006);
nand U16440 (N_16440,N_16151,N_16235);
nor U16441 (N_16441,N_16085,N_16080);
nand U16442 (N_16442,N_16221,N_16029);
xnor U16443 (N_16443,N_16033,N_16220);
or U16444 (N_16444,N_16222,N_16126);
or U16445 (N_16445,N_16060,N_16144);
nor U16446 (N_16446,N_16122,N_16144);
nand U16447 (N_16447,N_16150,N_16064);
and U16448 (N_16448,N_16226,N_16210);
or U16449 (N_16449,N_16009,N_16246);
nor U16450 (N_16450,N_16020,N_16066);
nand U16451 (N_16451,N_16228,N_16129);
nand U16452 (N_16452,N_16103,N_16101);
xor U16453 (N_16453,N_16110,N_16002);
xnor U16454 (N_16454,N_16092,N_16136);
nor U16455 (N_16455,N_16125,N_16131);
and U16456 (N_16456,N_16085,N_16082);
nor U16457 (N_16457,N_16012,N_16031);
or U16458 (N_16458,N_16195,N_16208);
xnor U16459 (N_16459,N_16160,N_16064);
or U16460 (N_16460,N_16169,N_16240);
and U16461 (N_16461,N_16010,N_16001);
or U16462 (N_16462,N_16008,N_16026);
nor U16463 (N_16463,N_16040,N_16181);
nor U16464 (N_16464,N_16061,N_16066);
nor U16465 (N_16465,N_16118,N_16030);
or U16466 (N_16466,N_16238,N_16087);
xnor U16467 (N_16467,N_16173,N_16111);
and U16468 (N_16468,N_16069,N_16076);
and U16469 (N_16469,N_16062,N_16121);
nor U16470 (N_16470,N_16024,N_16219);
nand U16471 (N_16471,N_16085,N_16211);
nor U16472 (N_16472,N_16139,N_16241);
and U16473 (N_16473,N_16036,N_16035);
xor U16474 (N_16474,N_16081,N_16051);
nor U16475 (N_16475,N_16213,N_16058);
nand U16476 (N_16476,N_16212,N_16013);
nand U16477 (N_16477,N_16175,N_16249);
xnor U16478 (N_16478,N_16036,N_16019);
xnor U16479 (N_16479,N_16013,N_16205);
nand U16480 (N_16480,N_16009,N_16225);
and U16481 (N_16481,N_16176,N_16012);
nor U16482 (N_16482,N_16230,N_16037);
nand U16483 (N_16483,N_16130,N_16144);
and U16484 (N_16484,N_16082,N_16077);
nand U16485 (N_16485,N_16078,N_16115);
and U16486 (N_16486,N_16158,N_16225);
or U16487 (N_16487,N_16009,N_16089);
nor U16488 (N_16488,N_16026,N_16165);
nor U16489 (N_16489,N_16200,N_16163);
xor U16490 (N_16490,N_16050,N_16112);
nand U16491 (N_16491,N_16155,N_16112);
nor U16492 (N_16492,N_16191,N_16233);
or U16493 (N_16493,N_16076,N_16144);
and U16494 (N_16494,N_16240,N_16153);
or U16495 (N_16495,N_16058,N_16094);
xnor U16496 (N_16496,N_16087,N_16116);
and U16497 (N_16497,N_16024,N_16218);
and U16498 (N_16498,N_16048,N_16161);
or U16499 (N_16499,N_16117,N_16245);
or U16500 (N_16500,N_16339,N_16368);
xnor U16501 (N_16501,N_16322,N_16491);
and U16502 (N_16502,N_16289,N_16316);
nand U16503 (N_16503,N_16420,N_16330);
xor U16504 (N_16504,N_16348,N_16478);
nand U16505 (N_16505,N_16477,N_16430);
xnor U16506 (N_16506,N_16421,N_16352);
or U16507 (N_16507,N_16253,N_16455);
and U16508 (N_16508,N_16338,N_16302);
and U16509 (N_16509,N_16408,N_16334);
nor U16510 (N_16510,N_16274,N_16268);
xor U16511 (N_16511,N_16323,N_16254);
xnor U16512 (N_16512,N_16300,N_16272);
xor U16513 (N_16513,N_16305,N_16394);
nand U16514 (N_16514,N_16402,N_16311);
nor U16515 (N_16515,N_16447,N_16418);
and U16516 (N_16516,N_16284,N_16483);
nor U16517 (N_16517,N_16457,N_16412);
nor U16518 (N_16518,N_16359,N_16269);
nand U16519 (N_16519,N_16397,N_16364);
xor U16520 (N_16520,N_16297,N_16286);
and U16521 (N_16521,N_16309,N_16470);
nand U16522 (N_16522,N_16446,N_16260);
nor U16523 (N_16523,N_16403,N_16489);
nand U16524 (N_16524,N_16479,N_16376);
or U16525 (N_16525,N_16357,N_16451);
nor U16526 (N_16526,N_16367,N_16429);
nor U16527 (N_16527,N_16458,N_16282);
nor U16528 (N_16528,N_16392,N_16431);
or U16529 (N_16529,N_16319,N_16422);
nand U16530 (N_16530,N_16321,N_16370);
nand U16531 (N_16531,N_16425,N_16276);
nand U16532 (N_16532,N_16303,N_16313);
or U16533 (N_16533,N_16285,N_16461);
or U16534 (N_16534,N_16486,N_16460);
or U16535 (N_16535,N_16354,N_16469);
xnor U16536 (N_16536,N_16317,N_16329);
or U16537 (N_16537,N_16391,N_16474);
xnor U16538 (N_16538,N_16490,N_16310);
xor U16539 (N_16539,N_16328,N_16335);
xnor U16540 (N_16540,N_16440,N_16320);
or U16541 (N_16541,N_16383,N_16463);
nor U16542 (N_16542,N_16405,N_16307);
nor U16543 (N_16543,N_16462,N_16445);
and U16544 (N_16544,N_16304,N_16351);
nand U16545 (N_16545,N_16433,N_16281);
nand U16546 (N_16546,N_16389,N_16251);
and U16547 (N_16547,N_16365,N_16390);
xnor U16548 (N_16548,N_16366,N_16312);
xnor U16549 (N_16549,N_16273,N_16318);
xnor U16550 (N_16550,N_16387,N_16496);
nand U16551 (N_16551,N_16417,N_16471);
xnor U16552 (N_16552,N_16277,N_16407);
and U16553 (N_16553,N_16344,N_16404);
nor U16554 (N_16554,N_16473,N_16441);
or U16555 (N_16555,N_16413,N_16279);
or U16556 (N_16556,N_16349,N_16291);
or U16557 (N_16557,N_16492,N_16416);
nand U16558 (N_16558,N_16258,N_16250);
and U16559 (N_16559,N_16290,N_16399);
and U16560 (N_16560,N_16466,N_16325);
nor U16561 (N_16561,N_16361,N_16427);
nor U16562 (N_16562,N_16371,N_16395);
xnor U16563 (N_16563,N_16375,N_16476);
or U16564 (N_16564,N_16278,N_16481);
and U16565 (N_16565,N_16259,N_16341);
or U16566 (N_16566,N_16373,N_16393);
and U16567 (N_16567,N_16257,N_16424);
nand U16568 (N_16568,N_16271,N_16275);
nor U16569 (N_16569,N_16327,N_16406);
nand U16570 (N_16570,N_16315,N_16343);
nand U16571 (N_16571,N_16332,N_16262);
or U16572 (N_16572,N_16467,N_16434);
nand U16573 (N_16573,N_16423,N_16299);
or U16574 (N_16574,N_16411,N_16443);
or U16575 (N_16575,N_16296,N_16306);
or U16576 (N_16576,N_16453,N_16295);
nand U16577 (N_16577,N_16252,N_16381);
nor U16578 (N_16578,N_16498,N_16409);
nand U16579 (N_16579,N_16380,N_16475);
and U16580 (N_16580,N_16428,N_16353);
and U16581 (N_16581,N_16464,N_16438);
nor U16582 (N_16582,N_16314,N_16465);
nand U16583 (N_16583,N_16324,N_16485);
or U16584 (N_16584,N_16439,N_16355);
and U16585 (N_16585,N_16472,N_16369);
nand U16586 (N_16586,N_16358,N_16267);
nor U16587 (N_16587,N_16326,N_16280);
nor U16588 (N_16588,N_16256,N_16386);
or U16589 (N_16589,N_16298,N_16488);
nand U16590 (N_16590,N_16456,N_16459);
or U16591 (N_16591,N_16377,N_16345);
nor U16592 (N_16592,N_16436,N_16493);
xor U16593 (N_16593,N_16410,N_16264);
xor U16594 (N_16594,N_16494,N_16255);
and U16595 (N_16595,N_16437,N_16263);
and U16596 (N_16596,N_16398,N_16374);
or U16597 (N_16597,N_16432,N_16435);
nor U16598 (N_16598,N_16333,N_16342);
nor U16599 (N_16599,N_16396,N_16487);
nand U16600 (N_16600,N_16452,N_16495);
xnor U16601 (N_16601,N_16360,N_16497);
nand U16602 (N_16602,N_16414,N_16442);
or U16603 (N_16603,N_16468,N_16347);
nor U16604 (N_16604,N_16265,N_16266);
or U16605 (N_16605,N_16499,N_16340);
or U16606 (N_16606,N_16385,N_16293);
and U16607 (N_16607,N_16292,N_16363);
and U16608 (N_16608,N_16480,N_16350);
nor U16609 (N_16609,N_16482,N_16426);
or U16610 (N_16610,N_16454,N_16379);
xnor U16611 (N_16611,N_16337,N_16331);
and U16612 (N_16612,N_16336,N_16288);
xnor U16613 (N_16613,N_16449,N_16450);
or U16614 (N_16614,N_16362,N_16401);
or U16615 (N_16615,N_16261,N_16400);
or U16616 (N_16616,N_16346,N_16484);
xor U16617 (N_16617,N_16378,N_16419);
or U16618 (N_16618,N_16287,N_16444);
xnor U16619 (N_16619,N_16382,N_16388);
and U16620 (N_16620,N_16384,N_16270);
and U16621 (N_16621,N_16301,N_16283);
xor U16622 (N_16622,N_16308,N_16372);
and U16623 (N_16623,N_16415,N_16356);
or U16624 (N_16624,N_16294,N_16448);
nor U16625 (N_16625,N_16344,N_16293);
xor U16626 (N_16626,N_16356,N_16491);
or U16627 (N_16627,N_16476,N_16445);
nand U16628 (N_16628,N_16328,N_16287);
nand U16629 (N_16629,N_16464,N_16253);
or U16630 (N_16630,N_16381,N_16293);
or U16631 (N_16631,N_16438,N_16461);
nor U16632 (N_16632,N_16378,N_16352);
and U16633 (N_16633,N_16287,N_16325);
and U16634 (N_16634,N_16270,N_16450);
nand U16635 (N_16635,N_16473,N_16375);
nand U16636 (N_16636,N_16353,N_16317);
or U16637 (N_16637,N_16278,N_16300);
or U16638 (N_16638,N_16491,N_16422);
nor U16639 (N_16639,N_16405,N_16369);
nand U16640 (N_16640,N_16463,N_16402);
and U16641 (N_16641,N_16407,N_16450);
or U16642 (N_16642,N_16334,N_16348);
and U16643 (N_16643,N_16467,N_16296);
nand U16644 (N_16644,N_16404,N_16439);
or U16645 (N_16645,N_16409,N_16306);
xnor U16646 (N_16646,N_16473,N_16436);
and U16647 (N_16647,N_16490,N_16434);
and U16648 (N_16648,N_16349,N_16478);
nor U16649 (N_16649,N_16388,N_16413);
xor U16650 (N_16650,N_16489,N_16447);
or U16651 (N_16651,N_16301,N_16332);
xor U16652 (N_16652,N_16313,N_16276);
or U16653 (N_16653,N_16417,N_16331);
nor U16654 (N_16654,N_16313,N_16424);
nand U16655 (N_16655,N_16325,N_16352);
nor U16656 (N_16656,N_16471,N_16484);
and U16657 (N_16657,N_16367,N_16412);
nor U16658 (N_16658,N_16476,N_16321);
nor U16659 (N_16659,N_16452,N_16426);
or U16660 (N_16660,N_16376,N_16444);
and U16661 (N_16661,N_16340,N_16345);
xor U16662 (N_16662,N_16305,N_16453);
nor U16663 (N_16663,N_16357,N_16375);
and U16664 (N_16664,N_16366,N_16498);
nor U16665 (N_16665,N_16336,N_16488);
xnor U16666 (N_16666,N_16257,N_16284);
nand U16667 (N_16667,N_16445,N_16458);
or U16668 (N_16668,N_16492,N_16495);
or U16669 (N_16669,N_16326,N_16314);
nor U16670 (N_16670,N_16484,N_16489);
nand U16671 (N_16671,N_16303,N_16261);
nand U16672 (N_16672,N_16439,N_16419);
and U16673 (N_16673,N_16305,N_16289);
xnor U16674 (N_16674,N_16421,N_16392);
or U16675 (N_16675,N_16351,N_16272);
nand U16676 (N_16676,N_16373,N_16346);
and U16677 (N_16677,N_16389,N_16405);
or U16678 (N_16678,N_16458,N_16350);
and U16679 (N_16679,N_16431,N_16490);
and U16680 (N_16680,N_16321,N_16467);
xor U16681 (N_16681,N_16403,N_16406);
xor U16682 (N_16682,N_16469,N_16357);
xnor U16683 (N_16683,N_16299,N_16366);
xor U16684 (N_16684,N_16299,N_16363);
xnor U16685 (N_16685,N_16356,N_16471);
nor U16686 (N_16686,N_16362,N_16290);
nor U16687 (N_16687,N_16283,N_16352);
nor U16688 (N_16688,N_16311,N_16498);
xor U16689 (N_16689,N_16490,N_16492);
and U16690 (N_16690,N_16258,N_16409);
nor U16691 (N_16691,N_16271,N_16291);
nor U16692 (N_16692,N_16397,N_16253);
or U16693 (N_16693,N_16292,N_16374);
nor U16694 (N_16694,N_16365,N_16335);
nand U16695 (N_16695,N_16313,N_16405);
or U16696 (N_16696,N_16344,N_16381);
nor U16697 (N_16697,N_16487,N_16418);
or U16698 (N_16698,N_16335,N_16289);
and U16699 (N_16699,N_16445,N_16305);
and U16700 (N_16700,N_16418,N_16302);
and U16701 (N_16701,N_16380,N_16270);
nand U16702 (N_16702,N_16464,N_16411);
nor U16703 (N_16703,N_16374,N_16378);
nor U16704 (N_16704,N_16264,N_16406);
nand U16705 (N_16705,N_16312,N_16354);
xnor U16706 (N_16706,N_16313,N_16302);
nor U16707 (N_16707,N_16389,N_16452);
nor U16708 (N_16708,N_16457,N_16413);
and U16709 (N_16709,N_16318,N_16314);
xor U16710 (N_16710,N_16269,N_16323);
xor U16711 (N_16711,N_16324,N_16490);
nand U16712 (N_16712,N_16483,N_16440);
and U16713 (N_16713,N_16490,N_16319);
or U16714 (N_16714,N_16384,N_16411);
nor U16715 (N_16715,N_16425,N_16349);
nand U16716 (N_16716,N_16475,N_16463);
nor U16717 (N_16717,N_16314,N_16398);
and U16718 (N_16718,N_16409,N_16488);
xor U16719 (N_16719,N_16410,N_16408);
xnor U16720 (N_16720,N_16465,N_16418);
or U16721 (N_16721,N_16362,N_16266);
nor U16722 (N_16722,N_16444,N_16273);
nor U16723 (N_16723,N_16459,N_16392);
xnor U16724 (N_16724,N_16338,N_16416);
nor U16725 (N_16725,N_16406,N_16262);
and U16726 (N_16726,N_16349,N_16453);
nand U16727 (N_16727,N_16431,N_16337);
nand U16728 (N_16728,N_16285,N_16498);
or U16729 (N_16729,N_16447,N_16337);
xor U16730 (N_16730,N_16276,N_16301);
or U16731 (N_16731,N_16348,N_16376);
nand U16732 (N_16732,N_16371,N_16286);
or U16733 (N_16733,N_16449,N_16414);
nand U16734 (N_16734,N_16497,N_16273);
nor U16735 (N_16735,N_16459,N_16332);
nand U16736 (N_16736,N_16403,N_16421);
nor U16737 (N_16737,N_16424,N_16340);
or U16738 (N_16738,N_16466,N_16486);
nor U16739 (N_16739,N_16391,N_16259);
nand U16740 (N_16740,N_16371,N_16431);
xor U16741 (N_16741,N_16319,N_16408);
and U16742 (N_16742,N_16403,N_16348);
and U16743 (N_16743,N_16292,N_16279);
or U16744 (N_16744,N_16421,N_16490);
nor U16745 (N_16745,N_16487,N_16476);
and U16746 (N_16746,N_16283,N_16317);
xnor U16747 (N_16747,N_16286,N_16262);
nand U16748 (N_16748,N_16278,N_16435);
or U16749 (N_16749,N_16357,N_16265);
nor U16750 (N_16750,N_16674,N_16646);
xnor U16751 (N_16751,N_16560,N_16583);
nor U16752 (N_16752,N_16599,N_16504);
nor U16753 (N_16753,N_16574,N_16555);
nand U16754 (N_16754,N_16729,N_16673);
nand U16755 (N_16755,N_16659,N_16691);
or U16756 (N_16756,N_16618,N_16605);
and U16757 (N_16757,N_16596,N_16679);
nor U16758 (N_16758,N_16669,N_16514);
nor U16759 (N_16759,N_16687,N_16629);
nand U16760 (N_16760,N_16545,N_16732);
and U16761 (N_16761,N_16593,N_16722);
nor U16762 (N_16762,N_16678,N_16620);
nor U16763 (N_16763,N_16578,N_16524);
nand U16764 (N_16764,N_16712,N_16727);
nor U16765 (N_16765,N_16698,N_16619);
and U16766 (N_16766,N_16600,N_16592);
or U16767 (N_16767,N_16503,N_16680);
nor U16768 (N_16768,N_16570,N_16643);
nor U16769 (N_16769,N_16696,N_16531);
nor U16770 (N_16770,N_16628,N_16562);
nor U16771 (N_16771,N_16515,N_16744);
xnor U16772 (N_16772,N_16742,N_16598);
xor U16773 (N_16773,N_16553,N_16601);
nand U16774 (N_16774,N_16533,N_16733);
nand U16775 (N_16775,N_16632,N_16580);
or U16776 (N_16776,N_16509,N_16731);
and U16777 (N_16777,N_16568,N_16645);
nor U16778 (N_16778,N_16611,N_16668);
and U16779 (N_16779,N_16563,N_16682);
nor U16780 (N_16780,N_16718,N_16711);
nand U16781 (N_16781,N_16723,N_16689);
nor U16782 (N_16782,N_16603,N_16644);
or U16783 (N_16783,N_16724,N_16567);
nand U16784 (N_16784,N_16653,N_16706);
nor U16785 (N_16785,N_16538,N_16561);
nor U16786 (N_16786,N_16725,N_16517);
nor U16787 (N_16787,N_16587,N_16667);
nor U16788 (N_16788,N_16702,N_16540);
or U16789 (N_16789,N_16715,N_16565);
nor U16790 (N_16790,N_16695,N_16686);
or U16791 (N_16791,N_16546,N_16735);
nor U16792 (N_16792,N_16683,N_16640);
and U16793 (N_16793,N_16613,N_16681);
or U16794 (N_16794,N_16717,N_16719);
nand U16795 (N_16795,N_16502,N_16526);
xnor U16796 (N_16796,N_16737,N_16595);
and U16797 (N_16797,N_16684,N_16530);
xor U16798 (N_16798,N_16510,N_16641);
or U16799 (N_16799,N_16739,N_16716);
nand U16800 (N_16800,N_16589,N_16720);
or U16801 (N_16801,N_16745,N_16617);
xnor U16802 (N_16802,N_16699,N_16528);
nand U16803 (N_16803,N_16547,N_16747);
and U16804 (N_16804,N_16506,N_16513);
xor U16805 (N_16805,N_16543,N_16606);
xor U16806 (N_16806,N_16590,N_16544);
and U16807 (N_16807,N_16591,N_16571);
nand U16808 (N_16808,N_16736,N_16639);
nand U16809 (N_16809,N_16707,N_16622);
xnor U16810 (N_16810,N_16597,N_16630);
nor U16811 (N_16811,N_16721,N_16521);
or U16812 (N_16812,N_16642,N_16559);
xnor U16813 (N_16813,N_16710,N_16648);
xnor U16814 (N_16814,N_16675,N_16728);
or U16815 (N_16815,N_16584,N_16658);
nand U16816 (N_16816,N_16516,N_16552);
and U16817 (N_16817,N_16505,N_16649);
and U16818 (N_16818,N_16647,N_16607);
nand U16819 (N_16819,N_16652,N_16638);
or U16820 (N_16820,N_16700,N_16581);
and U16821 (N_16821,N_16677,N_16532);
or U16822 (N_16822,N_16633,N_16701);
nand U16823 (N_16823,N_16549,N_16703);
xnor U16824 (N_16824,N_16661,N_16525);
and U16825 (N_16825,N_16650,N_16535);
nor U16826 (N_16826,N_16746,N_16726);
nor U16827 (N_16827,N_16582,N_16522);
nor U16828 (N_16828,N_16748,N_16697);
nand U16829 (N_16829,N_16730,N_16635);
and U16830 (N_16830,N_16738,N_16541);
nand U16831 (N_16831,N_16743,N_16550);
nor U16832 (N_16832,N_16501,N_16670);
nor U16833 (N_16833,N_16602,N_16542);
nand U16834 (N_16834,N_16623,N_16588);
nor U16835 (N_16835,N_16610,N_16539);
xor U16836 (N_16836,N_16564,N_16672);
or U16837 (N_16837,N_16520,N_16709);
nor U16838 (N_16838,N_16604,N_16536);
nor U16839 (N_16839,N_16688,N_16615);
and U16840 (N_16840,N_16627,N_16519);
or U16841 (N_16841,N_16507,N_16631);
and U16842 (N_16842,N_16654,N_16500);
and U16843 (N_16843,N_16566,N_16714);
and U16844 (N_16844,N_16676,N_16556);
and U16845 (N_16845,N_16554,N_16740);
nor U16846 (N_16846,N_16512,N_16609);
and U16847 (N_16847,N_16577,N_16713);
nor U16848 (N_16848,N_16579,N_16612);
and U16849 (N_16849,N_16527,N_16690);
nand U16850 (N_16850,N_16572,N_16508);
or U16851 (N_16851,N_16621,N_16523);
nor U16852 (N_16852,N_16557,N_16663);
or U16853 (N_16853,N_16655,N_16616);
nor U16854 (N_16854,N_16569,N_16624);
and U16855 (N_16855,N_16573,N_16558);
xor U16856 (N_16856,N_16694,N_16518);
xnor U16857 (N_16857,N_16666,N_16551);
nor U16858 (N_16858,N_16664,N_16708);
and U16859 (N_16859,N_16671,N_16705);
and U16860 (N_16860,N_16534,N_16657);
nor U16861 (N_16861,N_16656,N_16637);
xnor U16862 (N_16862,N_16626,N_16693);
nor U16863 (N_16863,N_16651,N_16537);
xor U16864 (N_16864,N_16692,N_16685);
xnor U16865 (N_16865,N_16575,N_16704);
nand U16866 (N_16866,N_16548,N_16529);
and U16867 (N_16867,N_16594,N_16665);
and U16868 (N_16868,N_16585,N_16660);
nand U16869 (N_16869,N_16511,N_16749);
nand U16870 (N_16870,N_16662,N_16625);
xor U16871 (N_16871,N_16614,N_16634);
xnor U16872 (N_16872,N_16636,N_16741);
nor U16873 (N_16873,N_16586,N_16734);
and U16874 (N_16874,N_16576,N_16608);
and U16875 (N_16875,N_16561,N_16533);
and U16876 (N_16876,N_16609,N_16578);
xnor U16877 (N_16877,N_16630,N_16614);
nor U16878 (N_16878,N_16531,N_16541);
and U16879 (N_16879,N_16607,N_16630);
nor U16880 (N_16880,N_16509,N_16634);
and U16881 (N_16881,N_16648,N_16567);
or U16882 (N_16882,N_16593,N_16500);
nand U16883 (N_16883,N_16743,N_16548);
or U16884 (N_16884,N_16704,N_16707);
nor U16885 (N_16885,N_16642,N_16522);
xnor U16886 (N_16886,N_16562,N_16660);
nand U16887 (N_16887,N_16547,N_16544);
and U16888 (N_16888,N_16704,N_16616);
xnor U16889 (N_16889,N_16556,N_16698);
and U16890 (N_16890,N_16728,N_16655);
nand U16891 (N_16891,N_16530,N_16573);
xnor U16892 (N_16892,N_16580,N_16536);
or U16893 (N_16893,N_16683,N_16675);
and U16894 (N_16894,N_16655,N_16511);
and U16895 (N_16895,N_16506,N_16683);
nand U16896 (N_16896,N_16668,N_16533);
nand U16897 (N_16897,N_16626,N_16713);
nor U16898 (N_16898,N_16659,N_16572);
xor U16899 (N_16899,N_16563,N_16705);
nor U16900 (N_16900,N_16577,N_16741);
or U16901 (N_16901,N_16642,N_16632);
nor U16902 (N_16902,N_16723,N_16534);
nor U16903 (N_16903,N_16726,N_16718);
or U16904 (N_16904,N_16670,N_16560);
or U16905 (N_16905,N_16600,N_16737);
nand U16906 (N_16906,N_16710,N_16578);
nand U16907 (N_16907,N_16688,N_16554);
or U16908 (N_16908,N_16639,N_16675);
and U16909 (N_16909,N_16733,N_16647);
xnor U16910 (N_16910,N_16653,N_16603);
and U16911 (N_16911,N_16537,N_16506);
nor U16912 (N_16912,N_16673,N_16628);
xor U16913 (N_16913,N_16642,N_16616);
and U16914 (N_16914,N_16738,N_16718);
nor U16915 (N_16915,N_16564,N_16631);
nor U16916 (N_16916,N_16724,N_16685);
nand U16917 (N_16917,N_16588,N_16574);
xor U16918 (N_16918,N_16735,N_16650);
or U16919 (N_16919,N_16656,N_16560);
and U16920 (N_16920,N_16697,N_16568);
nand U16921 (N_16921,N_16559,N_16538);
or U16922 (N_16922,N_16745,N_16554);
nor U16923 (N_16923,N_16680,N_16717);
nand U16924 (N_16924,N_16699,N_16671);
nand U16925 (N_16925,N_16653,N_16735);
and U16926 (N_16926,N_16738,N_16594);
nand U16927 (N_16927,N_16628,N_16715);
nand U16928 (N_16928,N_16679,N_16550);
xor U16929 (N_16929,N_16515,N_16527);
and U16930 (N_16930,N_16653,N_16675);
or U16931 (N_16931,N_16536,N_16598);
nand U16932 (N_16932,N_16629,N_16583);
nor U16933 (N_16933,N_16629,N_16637);
nor U16934 (N_16934,N_16736,N_16585);
xor U16935 (N_16935,N_16550,N_16672);
or U16936 (N_16936,N_16702,N_16746);
or U16937 (N_16937,N_16633,N_16567);
or U16938 (N_16938,N_16663,N_16742);
nor U16939 (N_16939,N_16707,N_16665);
and U16940 (N_16940,N_16616,N_16571);
xor U16941 (N_16941,N_16733,N_16508);
nand U16942 (N_16942,N_16587,N_16687);
or U16943 (N_16943,N_16661,N_16703);
and U16944 (N_16944,N_16545,N_16660);
xor U16945 (N_16945,N_16508,N_16622);
nor U16946 (N_16946,N_16564,N_16532);
nor U16947 (N_16947,N_16514,N_16564);
xnor U16948 (N_16948,N_16699,N_16584);
nor U16949 (N_16949,N_16738,N_16674);
or U16950 (N_16950,N_16589,N_16733);
and U16951 (N_16951,N_16569,N_16710);
and U16952 (N_16952,N_16654,N_16612);
xor U16953 (N_16953,N_16675,N_16531);
or U16954 (N_16954,N_16536,N_16714);
and U16955 (N_16955,N_16675,N_16591);
xnor U16956 (N_16956,N_16686,N_16548);
nor U16957 (N_16957,N_16657,N_16608);
xor U16958 (N_16958,N_16705,N_16651);
nand U16959 (N_16959,N_16637,N_16517);
or U16960 (N_16960,N_16724,N_16535);
xnor U16961 (N_16961,N_16541,N_16540);
xnor U16962 (N_16962,N_16675,N_16636);
and U16963 (N_16963,N_16549,N_16593);
nand U16964 (N_16964,N_16665,N_16529);
and U16965 (N_16965,N_16657,N_16555);
nor U16966 (N_16966,N_16706,N_16678);
or U16967 (N_16967,N_16688,N_16604);
xor U16968 (N_16968,N_16734,N_16648);
and U16969 (N_16969,N_16604,N_16583);
xnor U16970 (N_16970,N_16544,N_16645);
and U16971 (N_16971,N_16749,N_16720);
nor U16972 (N_16972,N_16624,N_16737);
nor U16973 (N_16973,N_16598,N_16522);
or U16974 (N_16974,N_16523,N_16709);
and U16975 (N_16975,N_16737,N_16711);
and U16976 (N_16976,N_16705,N_16531);
and U16977 (N_16977,N_16556,N_16675);
xnor U16978 (N_16978,N_16534,N_16716);
and U16979 (N_16979,N_16640,N_16694);
nor U16980 (N_16980,N_16696,N_16583);
nor U16981 (N_16981,N_16526,N_16604);
nor U16982 (N_16982,N_16570,N_16511);
or U16983 (N_16983,N_16607,N_16717);
and U16984 (N_16984,N_16619,N_16647);
nor U16985 (N_16985,N_16690,N_16593);
nor U16986 (N_16986,N_16695,N_16621);
or U16987 (N_16987,N_16539,N_16698);
nand U16988 (N_16988,N_16652,N_16522);
and U16989 (N_16989,N_16574,N_16680);
and U16990 (N_16990,N_16694,N_16716);
or U16991 (N_16991,N_16614,N_16655);
or U16992 (N_16992,N_16589,N_16701);
or U16993 (N_16993,N_16511,N_16521);
or U16994 (N_16994,N_16538,N_16539);
nand U16995 (N_16995,N_16738,N_16621);
nor U16996 (N_16996,N_16611,N_16729);
nand U16997 (N_16997,N_16536,N_16539);
nor U16998 (N_16998,N_16522,N_16654);
or U16999 (N_16999,N_16523,N_16681);
xor U17000 (N_17000,N_16914,N_16782);
and U17001 (N_17001,N_16826,N_16961);
or U17002 (N_17002,N_16817,N_16976);
or U17003 (N_17003,N_16863,N_16770);
or U17004 (N_17004,N_16904,N_16780);
xor U17005 (N_17005,N_16963,N_16991);
or U17006 (N_17006,N_16879,N_16762);
or U17007 (N_17007,N_16870,N_16835);
nand U17008 (N_17008,N_16752,N_16843);
and U17009 (N_17009,N_16801,N_16853);
and U17010 (N_17010,N_16769,N_16758);
nand U17011 (N_17011,N_16791,N_16775);
nor U17012 (N_17012,N_16829,N_16921);
nor U17013 (N_17013,N_16908,N_16873);
or U17014 (N_17014,N_16905,N_16966);
nand U17015 (N_17015,N_16947,N_16882);
and U17016 (N_17016,N_16916,N_16925);
nand U17017 (N_17017,N_16819,N_16959);
nand U17018 (N_17018,N_16943,N_16811);
xor U17019 (N_17019,N_16836,N_16955);
nor U17020 (N_17020,N_16933,N_16844);
nor U17021 (N_17021,N_16761,N_16849);
nor U17022 (N_17022,N_16831,N_16965);
and U17023 (N_17023,N_16755,N_16964);
xor U17024 (N_17024,N_16796,N_16804);
nand U17025 (N_17025,N_16894,N_16909);
and U17026 (N_17026,N_16907,N_16893);
and U17027 (N_17027,N_16917,N_16821);
or U17028 (N_17028,N_16828,N_16987);
and U17029 (N_17029,N_16753,N_16846);
xor U17030 (N_17030,N_16865,N_16932);
or U17031 (N_17031,N_16906,N_16954);
and U17032 (N_17032,N_16881,N_16875);
xor U17033 (N_17033,N_16872,N_16839);
xor U17034 (N_17034,N_16986,N_16931);
xnor U17035 (N_17035,N_16998,N_16866);
xnor U17036 (N_17036,N_16812,N_16915);
xor U17037 (N_17037,N_16969,N_16878);
xnor U17038 (N_17038,N_16850,N_16999);
and U17039 (N_17039,N_16759,N_16785);
and U17040 (N_17040,N_16869,N_16848);
or U17041 (N_17041,N_16860,N_16800);
or U17042 (N_17042,N_16806,N_16945);
and U17043 (N_17043,N_16897,N_16951);
nor U17044 (N_17044,N_16940,N_16838);
or U17045 (N_17045,N_16950,N_16797);
nor U17046 (N_17046,N_16868,N_16901);
xor U17047 (N_17047,N_16939,N_16934);
and U17048 (N_17048,N_16985,N_16818);
xnor U17049 (N_17049,N_16960,N_16974);
or U17050 (N_17050,N_16781,N_16900);
or U17051 (N_17051,N_16874,N_16816);
nor U17052 (N_17052,N_16920,N_16927);
xor U17053 (N_17053,N_16751,N_16994);
and U17054 (N_17054,N_16795,N_16984);
and U17055 (N_17055,N_16980,N_16786);
nor U17056 (N_17056,N_16792,N_16822);
nand U17057 (N_17057,N_16857,N_16810);
and U17058 (N_17058,N_16824,N_16832);
and U17059 (N_17059,N_16855,N_16938);
nand U17060 (N_17060,N_16990,N_16793);
and U17061 (N_17061,N_16929,N_16978);
nor U17062 (N_17062,N_16772,N_16983);
nand U17063 (N_17063,N_16776,N_16956);
xor U17064 (N_17064,N_16837,N_16884);
or U17065 (N_17065,N_16820,N_16883);
and U17066 (N_17066,N_16750,N_16948);
and U17067 (N_17067,N_16852,N_16970);
nor U17068 (N_17068,N_16937,N_16977);
nand U17069 (N_17069,N_16973,N_16913);
nor U17070 (N_17070,N_16975,N_16841);
nor U17071 (N_17071,N_16787,N_16981);
xor U17072 (N_17072,N_16946,N_16996);
and U17073 (N_17073,N_16774,N_16859);
nand U17074 (N_17074,N_16888,N_16936);
xnor U17075 (N_17075,N_16886,N_16988);
nand U17076 (N_17076,N_16896,N_16842);
and U17077 (N_17077,N_16845,N_16766);
nand U17078 (N_17078,N_16840,N_16771);
nand U17079 (N_17079,N_16928,N_16808);
and U17080 (N_17080,N_16911,N_16784);
nor U17081 (N_17081,N_16899,N_16757);
nor U17082 (N_17082,N_16861,N_16887);
nand U17083 (N_17083,N_16891,N_16760);
or U17084 (N_17084,N_16944,N_16789);
or U17085 (N_17085,N_16778,N_16813);
xor U17086 (N_17086,N_16754,N_16779);
nand U17087 (N_17087,N_16919,N_16799);
xnor U17088 (N_17088,N_16967,N_16885);
nand U17089 (N_17089,N_16924,N_16807);
and U17090 (N_17090,N_16773,N_16968);
nand U17091 (N_17091,N_16798,N_16935);
or U17092 (N_17092,N_16823,N_16867);
xnor U17093 (N_17093,N_16902,N_16982);
nand U17094 (N_17094,N_16877,N_16972);
xor U17095 (N_17095,N_16993,N_16992);
xnor U17096 (N_17096,N_16858,N_16949);
or U17097 (N_17097,N_16788,N_16802);
nor U17098 (N_17098,N_16790,N_16912);
and U17099 (N_17099,N_16803,N_16922);
or U17100 (N_17100,N_16847,N_16989);
and U17101 (N_17101,N_16809,N_16903);
or U17102 (N_17102,N_16815,N_16756);
and U17103 (N_17103,N_16825,N_16856);
and U17104 (N_17104,N_16995,N_16962);
nor U17105 (N_17105,N_16864,N_16997);
or U17106 (N_17106,N_16830,N_16923);
and U17107 (N_17107,N_16918,N_16805);
xor U17108 (N_17108,N_16910,N_16880);
and U17109 (N_17109,N_16767,N_16765);
xor U17110 (N_17110,N_16763,N_16930);
nor U17111 (N_17111,N_16890,N_16898);
nor U17112 (N_17112,N_16876,N_16889);
nor U17113 (N_17113,N_16926,N_16854);
and U17114 (N_17114,N_16892,N_16777);
or U17115 (N_17115,N_16952,N_16768);
nor U17116 (N_17116,N_16827,N_16794);
and U17117 (N_17117,N_16833,N_16871);
xnor U17118 (N_17118,N_16834,N_16941);
nor U17119 (N_17119,N_16979,N_16957);
nor U17120 (N_17120,N_16958,N_16942);
nand U17121 (N_17121,N_16971,N_16851);
or U17122 (N_17122,N_16862,N_16764);
or U17123 (N_17123,N_16783,N_16953);
or U17124 (N_17124,N_16814,N_16895);
nand U17125 (N_17125,N_16830,N_16909);
xor U17126 (N_17126,N_16929,N_16861);
and U17127 (N_17127,N_16940,N_16754);
or U17128 (N_17128,N_16779,N_16913);
or U17129 (N_17129,N_16904,N_16806);
nand U17130 (N_17130,N_16882,N_16943);
nand U17131 (N_17131,N_16818,N_16955);
nand U17132 (N_17132,N_16857,N_16883);
or U17133 (N_17133,N_16914,N_16750);
and U17134 (N_17134,N_16895,N_16759);
and U17135 (N_17135,N_16863,N_16857);
nand U17136 (N_17136,N_16936,N_16754);
and U17137 (N_17137,N_16949,N_16961);
nor U17138 (N_17138,N_16918,N_16968);
and U17139 (N_17139,N_16851,N_16759);
or U17140 (N_17140,N_16772,N_16868);
nand U17141 (N_17141,N_16824,N_16893);
or U17142 (N_17142,N_16987,N_16892);
and U17143 (N_17143,N_16908,N_16905);
or U17144 (N_17144,N_16770,N_16873);
xor U17145 (N_17145,N_16893,N_16865);
xor U17146 (N_17146,N_16963,N_16757);
and U17147 (N_17147,N_16965,N_16851);
and U17148 (N_17148,N_16779,N_16912);
and U17149 (N_17149,N_16805,N_16986);
nand U17150 (N_17150,N_16808,N_16888);
nand U17151 (N_17151,N_16838,N_16830);
nand U17152 (N_17152,N_16774,N_16816);
nand U17153 (N_17153,N_16923,N_16915);
nand U17154 (N_17154,N_16962,N_16752);
nand U17155 (N_17155,N_16841,N_16942);
xnor U17156 (N_17156,N_16911,N_16922);
nor U17157 (N_17157,N_16972,N_16973);
nand U17158 (N_17158,N_16808,N_16964);
or U17159 (N_17159,N_16774,N_16939);
xor U17160 (N_17160,N_16908,N_16927);
nor U17161 (N_17161,N_16855,N_16876);
nor U17162 (N_17162,N_16754,N_16858);
xnor U17163 (N_17163,N_16878,N_16819);
xor U17164 (N_17164,N_16984,N_16814);
or U17165 (N_17165,N_16976,N_16806);
or U17166 (N_17166,N_16832,N_16924);
nand U17167 (N_17167,N_16966,N_16907);
or U17168 (N_17168,N_16915,N_16760);
and U17169 (N_17169,N_16994,N_16817);
nand U17170 (N_17170,N_16833,N_16928);
and U17171 (N_17171,N_16763,N_16940);
and U17172 (N_17172,N_16992,N_16985);
nor U17173 (N_17173,N_16870,N_16776);
xnor U17174 (N_17174,N_16937,N_16820);
nor U17175 (N_17175,N_16967,N_16853);
or U17176 (N_17176,N_16902,N_16761);
nand U17177 (N_17177,N_16900,N_16863);
xor U17178 (N_17178,N_16916,N_16879);
and U17179 (N_17179,N_16817,N_16991);
nand U17180 (N_17180,N_16757,N_16869);
nor U17181 (N_17181,N_16801,N_16948);
xor U17182 (N_17182,N_16983,N_16908);
and U17183 (N_17183,N_16980,N_16845);
nor U17184 (N_17184,N_16930,N_16954);
nand U17185 (N_17185,N_16983,N_16762);
nand U17186 (N_17186,N_16970,N_16936);
nand U17187 (N_17187,N_16787,N_16881);
nand U17188 (N_17188,N_16937,N_16818);
and U17189 (N_17189,N_16803,N_16985);
nor U17190 (N_17190,N_16819,N_16809);
xnor U17191 (N_17191,N_16817,N_16770);
nand U17192 (N_17192,N_16971,N_16989);
and U17193 (N_17193,N_16958,N_16937);
or U17194 (N_17194,N_16919,N_16842);
nor U17195 (N_17195,N_16829,N_16781);
nor U17196 (N_17196,N_16874,N_16795);
or U17197 (N_17197,N_16907,N_16752);
nor U17198 (N_17198,N_16758,N_16916);
or U17199 (N_17199,N_16821,N_16791);
xor U17200 (N_17200,N_16782,N_16964);
and U17201 (N_17201,N_16778,N_16948);
or U17202 (N_17202,N_16830,N_16861);
and U17203 (N_17203,N_16969,N_16760);
xor U17204 (N_17204,N_16787,N_16816);
nor U17205 (N_17205,N_16800,N_16895);
and U17206 (N_17206,N_16886,N_16890);
and U17207 (N_17207,N_16986,N_16824);
or U17208 (N_17208,N_16805,N_16976);
xnor U17209 (N_17209,N_16778,N_16801);
xnor U17210 (N_17210,N_16804,N_16883);
nor U17211 (N_17211,N_16939,N_16838);
and U17212 (N_17212,N_16789,N_16773);
nand U17213 (N_17213,N_16805,N_16756);
or U17214 (N_17214,N_16976,N_16760);
nor U17215 (N_17215,N_16839,N_16798);
nand U17216 (N_17216,N_16920,N_16765);
and U17217 (N_17217,N_16857,N_16939);
nor U17218 (N_17218,N_16964,N_16954);
nand U17219 (N_17219,N_16858,N_16873);
or U17220 (N_17220,N_16837,N_16980);
nand U17221 (N_17221,N_16908,N_16887);
or U17222 (N_17222,N_16894,N_16752);
xnor U17223 (N_17223,N_16879,N_16805);
nor U17224 (N_17224,N_16802,N_16860);
or U17225 (N_17225,N_16763,N_16856);
nor U17226 (N_17226,N_16913,N_16934);
nor U17227 (N_17227,N_16887,N_16949);
or U17228 (N_17228,N_16901,N_16963);
nor U17229 (N_17229,N_16905,N_16929);
or U17230 (N_17230,N_16925,N_16824);
nand U17231 (N_17231,N_16951,N_16880);
nor U17232 (N_17232,N_16904,N_16900);
and U17233 (N_17233,N_16782,N_16801);
xnor U17234 (N_17234,N_16924,N_16908);
xnor U17235 (N_17235,N_16925,N_16760);
xnor U17236 (N_17236,N_16920,N_16893);
xnor U17237 (N_17237,N_16938,N_16785);
xor U17238 (N_17238,N_16788,N_16980);
or U17239 (N_17239,N_16820,N_16948);
nand U17240 (N_17240,N_16819,N_16811);
nand U17241 (N_17241,N_16919,N_16920);
nand U17242 (N_17242,N_16807,N_16901);
and U17243 (N_17243,N_16986,N_16774);
nor U17244 (N_17244,N_16954,N_16806);
or U17245 (N_17245,N_16765,N_16903);
nand U17246 (N_17246,N_16946,N_16942);
or U17247 (N_17247,N_16825,N_16834);
and U17248 (N_17248,N_16995,N_16953);
nand U17249 (N_17249,N_16930,N_16894);
or U17250 (N_17250,N_17022,N_17012);
nand U17251 (N_17251,N_17002,N_17231);
xor U17252 (N_17252,N_17114,N_17135);
nor U17253 (N_17253,N_17161,N_17194);
or U17254 (N_17254,N_17168,N_17040);
nand U17255 (N_17255,N_17075,N_17056);
or U17256 (N_17256,N_17226,N_17133);
nor U17257 (N_17257,N_17191,N_17013);
or U17258 (N_17258,N_17240,N_17156);
and U17259 (N_17259,N_17228,N_17110);
nand U17260 (N_17260,N_17151,N_17188);
xor U17261 (N_17261,N_17158,N_17139);
nor U17262 (N_17262,N_17061,N_17180);
xnor U17263 (N_17263,N_17234,N_17044);
or U17264 (N_17264,N_17189,N_17082);
and U17265 (N_17265,N_17247,N_17121);
nor U17266 (N_17266,N_17091,N_17236);
and U17267 (N_17267,N_17214,N_17016);
and U17268 (N_17268,N_17045,N_17073);
nand U17269 (N_17269,N_17124,N_17178);
nor U17270 (N_17270,N_17097,N_17205);
or U17271 (N_17271,N_17068,N_17127);
nand U17272 (N_17272,N_17193,N_17120);
and U17273 (N_17273,N_17185,N_17209);
nor U17274 (N_17274,N_17020,N_17103);
and U17275 (N_17275,N_17108,N_17212);
nand U17276 (N_17276,N_17017,N_17142);
nand U17277 (N_17277,N_17187,N_17059);
xnor U17278 (N_17278,N_17245,N_17119);
nor U17279 (N_17279,N_17003,N_17229);
nand U17280 (N_17280,N_17057,N_17049);
xnor U17281 (N_17281,N_17177,N_17223);
and U17282 (N_17282,N_17125,N_17140);
xnor U17283 (N_17283,N_17102,N_17159);
and U17284 (N_17284,N_17173,N_17208);
and U17285 (N_17285,N_17046,N_17227);
xor U17286 (N_17286,N_17146,N_17081);
nor U17287 (N_17287,N_17170,N_17089);
nor U17288 (N_17288,N_17101,N_17238);
nor U17289 (N_17289,N_17080,N_17216);
or U17290 (N_17290,N_17006,N_17217);
or U17291 (N_17291,N_17092,N_17064);
nor U17292 (N_17292,N_17077,N_17203);
and U17293 (N_17293,N_17136,N_17035);
or U17294 (N_17294,N_17220,N_17066);
nand U17295 (N_17295,N_17011,N_17079);
nand U17296 (N_17296,N_17036,N_17113);
or U17297 (N_17297,N_17009,N_17184);
xor U17298 (N_17298,N_17069,N_17058);
and U17299 (N_17299,N_17005,N_17087);
and U17300 (N_17300,N_17129,N_17083);
and U17301 (N_17301,N_17132,N_17128);
and U17302 (N_17302,N_17162,N_17175);
xnor U17303 (N_17303,N_17242,N_17026);
xor U17304 (N_17304,N_17050,N_17048);
or U17305 (N_17305,N_17222,N_17152);
and U17306 (N_17306,N_17138,N_17106);
nand U17307 (N_17307,N_17165,N_17027);
nor U17308 (N_17308,N_17169,N_17105);
xor U17309 (N_17309,N_17099,N_17034);
or U17310 (N_17310,N_17218,N_17207);
or U17311 (N_17311,N_17112,N_17248);
and U17312 (N_17312,N_17211,N_17055);
xor U17313 (N_17313,N_17153,N_17015);
or U17314 (N_17314,N_17190,N_17210);
nor U17315 (N_17315,N_17021,N_17104);
nand U17316 (N_17316,N_17241,N_17024);
and U17317 (N_17317,N_17008,N_17031);
xor U17318 (N_17318,N_17116,N_17143);
or U17319 (N_17319,N_17230,N_17070);
xor U17320 (N_17320,N_17076,N_17160);
and U17321 (N_17321,N_17171,N_17122);
xor U17322 (N_17322,N_17225,N_17232);
or U17323 (N_17323,N_17086,N_17233);
and U17324 (N_17324,N_17038,N_17117);
or U17325 (N_17325,N_17172,N_17023);
nand U17326 (N_17326,N_17157,N_17237);
nor U17327 (N_17327,N_17004,N_17001);
nand U17328 (N_17328,N_17098,N_17192);
or U17329 (N_17329,N_17224,N_17088);
xor U17330 (N_17330,N_17052,N_17130);
nand U17331 (N_17331,N_17196,N_17033);
nor U17332 (N_17332,N_17067,N_17145);
nand U17333 (N_17333,N_17246,N_17032);
nor U17334 (N_17334,N_17197,N_17094);
xor U17335 (N_17335,N_17018,N_17063);
nor U17336 (N_17336,N_17164,N_17167);
and U17337 (N_17337,N_17141,N_17147);
nor U17338 (N_17338,N_17007,N_17215);
and U17339 (N_17339,N_17085,N_17176);
xor U17340 (N_17340,N_17239,N_17029);
nand U17341 (N_17341,N_17243,N_17093);
nand U17342 (N_17342,N_17062,N_17039);
or U17343 (N_17343,N_17201,N_17144);
or U17344 (N_17344,N_17150,N_17047);
nor U17345 (N_17345,N_17221,N_17131);
nand U17346 (N_17346,N_17219,N_17134);
and U17347 (N_17347,N_17042,N_17244);
or U17348 (N_17348,N_17014,N_17051);
nor U17349 (N_17349,N_17054,N_17249);
and U17350 (N_17350,N_17149,N_17072);
nand U17351 (N_17351,N_17183,N_17179);
xor U17352 (N_17352,N_17123,N_17090);
xor U17353 (N_17353,N_17053,N_17010);
xor U17354 (N_17354,N_17198,N_17199);
xnor U17355 (N_17355,N_17181,N_17213);
xor U17356 (N_17356,N_17202,N_17019);
and U17357 (N_17357,N_17155,N_17074);
and U17358 (N_17358,N_17100,N_17096);
and U17359 (N_17359,N_17182,N_17030);
or U17360 (N_17360,N_17148,N_17025);
nand U17361 (N_17361,N_17186,N_17206);
xnor U17362 (N_17362,N_17041,N_17071);
nor U17363 (N_17363,N_17078,N_17118);
and U17364 (N_17364,N_17043,N_17137);
xor U17365 (N_17365,N_17028,N_17111);
nor U17366 (N_17366,N_17107,N_17060);
xor U17367 (N_17367,N_17163,N_17095);
nor U17368 (N_17368,N_17000,N_17166);
nand U17369 (N_17369,N_17065,N_17084);
and U17370 (N_17370,N_17109,N_17154);
xnor U17371 (N_17371,N_17126,N_17204);
nand U17372 (N_17372,N_17200,N_17195);
nor U17373 (N_17373,N_17235,N_17115);
nand U17374 (N_17374,N_17174,N_17037);
or U17375 (N_17375,N_17180,N_17168);
nor U17376 (N_17376,N_17094,N_17246);
nand U17377 (N_17377,N_17228,N_17162);
and U17378 (N_17378,N_17222,N_17099);
and U17379 (N_17379,N_17165,N_17047);
and U17380 (N_17380,N_17175,N_17194);
xor U17381 (N_17381,N_17019,N_17217);
and U17382 (N_17382,N_17025,N_17142);
and U17383 (N_17383,N_17238,N_17022);
nand U17384 (N_17384,N_17179,N_17160);
and U17385 (N_17385,N_17214,N_17137);
or U17386 (N_17386,N_17201,N_17000);
nand U17387 (N_17387,N_17001,N_17147);
xnor U17388 (N_17388,N_17234,N_17178);
or U17389 (N_17389,N_17014,N_17130);
nor U17390 (N_17390,N_17232,N_17067);
xor U17391 (N_17391,N_17208,N_17176);
nand U17392 (N_17392,N_17120,N_17215);
or U17393 (N_17393,N_17111,N_17047);
xnor U17394 (N_17394,N_17204,N_17177);
nor U17395 (N_17395,N_17044,N_17133);
and U17396 (N_17396,N_17230,N_17139);
xor U17397 (N_17397,N_17209,N_17241);
nand U17398 (N_17398,N_17012,N_17218);
and U17399 (N_17399,N_17216,N_17008);
or U17400 (N_17400,N_17236,N_17099);
and U17401 (N_17401,N_17026,N_17053);
nor U17402 (N_17402,N_17011,N_17134);
or U17403 (N_17403,N_17089,N_17060);
xnor U17404 (N_17404,N_17092,N_17163);
xnor U17405 (N_17405,N_17088,N_17035);
xor U17406 (N_17406,N_17031,N_17188);
nand U17407 (N_17407,N_17224,N_17013);
nand U17408 (N_17408,N_17141,N_17156);
or U17409 (N_17409,N_17190,N_17074);
nand U17410 (N_17410,N_17072,N_17243);
and U17411 (N_17411,N_17211,N_17213);
and U17412 (N_17412,N_17137,N_17215);
and U17413 (N_17413,N_17120,N_17118);
xnor U17414 (N_17414,N_17107,N_17170);
or U17415 (N_17415,N_17114,N_17028);
xor U17416 (N_17416,N_17027,N_17086);
nor U17417 (N_17417,N_17054,N_17048);
xnor U17418 (N_17418,N_17013,N_17027);
nor U17419 (N_17419,N_17109,N_17053);
xor U17420 (N_17420,N_17155,N_17181);
nand U17421 (N_17421,N_17085,N_17155);
and U17422 (N_17422,N_17041,N_17209);
nor U17423 (N_17423,N_17221,N_17124);
nor U17424 (N_17424,N_17109,N_17144);
xor U17425 (N_17425,N_17169,N_17179);
nand U17426 (N_17426,N_17139,N_17165);
and U17427 (N_17427,N_17221,N_17187);
nor U17428 (N_17428,N_17106,N_17110);
or U17429 (N_17429,N_17145,N_17014);
xnor U17430 (N_17430,N_17156,N_17030);
and U17431 (N_17431,N_17122,N_17133);
xor U17432 (N_17432,N_17230,N_17232);
nor U17433 (N_17433,N_17134,N_17170);
nand U17434 (N_17434,N_17060,N_17233);
nand U17435 (N_17435,N_17135,N_17002);
nand U17436 (N_17436,N_17014,N_17112);
xnor U17437 (N_17437,N_17248,N_17045);
xnor U17438 (N_17438,N_17199,N_17239);
or U17439 (N_17439,N_17191,N_17037);
nand U17440 (N_17440,N_17015,N_17194);
and U17441 (N_17441,N_17212,N_17246);
nand U17442 (N_17442,N_17213,N_17138);
nand U17443 (N_17443,N_17097,N_17046);
and U17444 (N_17444,N_17182,N_17137);
nor U17445 (N_17445,N_17055,N_17034);
xor U17446 (N_17446,N_17002,N_17037);
xor U17447 (N_17447,N_17111,N_17219);
or U17448 (N_17448,N_17231,N_17134);
nand U17449 (N_17449,N_17155,N_17094);
or U17450 (N_17450,N_17185,N_17053);
nor U17451 (N_17451,N_17207,N_17085);
and U17452 (N_17452,N_17189,N_17192);
xor U17453 (N_17453,N_17215,N_17121);
xor U17454 (N_17454,N_17063,N_17180);
nand U17455 (N_17455,N_17227,N_17057);
nand U17456 (N_17456,N_17067,N_17002);
xnor U17457 (N_17457,N_17022,N_17247);
nor U17458 (N_17458,N_17196,N_17039);
and U17459 (N_17459,N_17118,N_17178);
and U17460 (N_17460,N_17048,N_17122);
or U17461 (N_17461,N_17225,N_17024);
nor U17462 (N_17462,N_17249,N_17087);
and U17463 (N_17463,N_17096,N_17058);
or U17464 (N_17464,N_17192,N_17175);
or U17465 (N_17465,N_17228,N_17222);
and U17466 (N_17466,N_17066,N_17035);
nor U17467 (N_17467,N_17117,N_17232);
nand U17468 (N_17468,N_17028,N_17136);
nor U17469 (N_17469,N_17225,N_17168);
and U17470 (N_17470,N_17206,N_17096);
nand U17471 (N_17471,N_17081,N_17046);
or U17472 (N_17472,N_17139,N_17030);
and U17473 (N_17473,N_17037,N_17089);
nor U17474 (N_17474,N_17231,N_17091);
nor U17475 (N_17475,N_17022,N_17099);
nor U17476 (N_17476,N_17184,N_17150);
xor U17477 (N_17477,N_17241,N_17158);
xnor U17478 (N_17478,N_17053,N_17056);
or U17479 (N_17479,N_17245,N_17097);
and U17480 (N_17480,N_17107,N_17233);
or U17481 (N_17481,N_17241,N_17110);
xnor U17482 (N_17482,N_17194,N_17097);
and U17483 (N_17483,N_17025,N_17223);
nand U17484 (N_17484,N_17006,N_17007);
xnor U17485 (N_17485,N_17034,N_17166);
nor U17486 (N_17486,N_17012,N_17167);
xnor U17487 (N_17487,N_17187,N_17054);
nand U17488 (N_17488,N_17217,N_17095);
xor U17489 (N_17489,N_17082,N_17044);
nand U17490 (N_17490,N_17036,N_17201);
or U17491 (N_17491,N_17173,N_17085);
and U17492 (N_17492,N_17166,N_17142);
nand U17493 (N_17493,N_17225,N_17156);
nor U17494 (N_17494,N_17003,N_17214);
or U17495 (N_17495,N_17176,N_17015);
nand U17496 (N_17496,N_17111,N_17053);
xor U17497 (N_17497,N_17138,N_17170);
nand U17498 (N_17498,N_17044,N_17092);
and U17499 (N_17499,N_17059,N_17066);
xnor U17500 (N_17500,N_17476,N_17304);
xor U17501 (N_17501,N_17486,N_17398);
and U17502 (N_17502,N_17282,N_17350);
nor U17503 (N_17503,N_17359,N_17330);
nor U17504 (N_17504,N_17425,N_17440);
xor U17505 (N_17505,N_17384,N_17268);
nor U17506 (N_17506,N_17441,N_17395);
or U17507 (N_17507,N_17401,N_17275);
nor U17508 (N_17508,N_17494,N_17352);
xor U17509 (N_17509,N_17274,N_17310);
nor U17510 (N_17510,N_17251,N_17323);
nand U17511 (N_17511,N_17293,N_17286);
and U17512 (N_17512,N_17443,N_17387);
nand U17513 (N_17513,N_17250,N_17344);
xnor U17514 (N_17514,N_17396,N_17462);
xnor U17515 (N_17515,N_17355,N_17257);
xor U17516 (N_17516,N_17339,N_17289);
and U17517 (N_17517,N_17382,N_17321);
or U17518 (N_17518,N_17326,N_17393);
xnor U17519 (N_17519,N_17328,N_17356);
and U17520 (N_17520,N_17422,N_17403);
xor U17521 (N_17521,N_17327,N_17402);
and U17522 (N_17522,N_17347,N_17263);
xor U17523 (N_17523,N_17320,N_17270);
or U17524 (N_17524,N_17291,N_17394);
or U17525 (N_17525,N_17271,N_17492);
nor U17526 (N_17526,N_17331,N_17409);
or U17527 (N_17527,N_17253,N_17258);
nand U17528 (N_17528,N_17285,N_17433);
and U17529 (N_17529,N_17435,N_17255);
nand U17530 (N_17530,N_17334,N_17360);
xnor U17531 (N_17531,N_17497,N_17496);
nand U17532 (N_17532,N_17390,N_17485);
nand U17533 (N_17533,N_17333,N_17472);
nand U17534 (N_17534,N_17414,N_17454);
nand U17535 (N_17535,N_17426,N_17442);
xor U17536 (N_17536,N_17340,N_17269);
and U17537 (N_17537,N_17314,N_17256);
nor U17538 (N_17538,N_17421,N_17385);
nand U17539 (N_17539,N_17380,N_17423);
nand U17540 (N_17540,N_17351,N_17439);
xor U17541 (N_17541,N_17300,N_17303);
nor U17542 (N_17542,N_17308,N_17495);
and U17543 (N_17543,N_17365,N_17260);
or U17544 (N_17544,N_17406,N_17436);
xor U17545 (N_17545,N_17397,N_17337);
xor U17546 (N_17546,N_17307,N_17488);
nand U17547 (N_17547,N_17420,N_17467);
nor U17548 (N_17548,N_17287,N_17459);
or U17549 (N_17549,N_17391,N_17348);
nand U17550 (N_17550,N_17312,N_17411);
xnor U17551 (N_17551,N_17335,N_17410);
nand U17552 (N_17552,N_17446,N_17464);
nand U17553 (N_17553,N_17283,N_17273);
nand U17554 (N_17554,N_17315,N_17461);
nand U17555 (N_17555,N_17437,N_17412);
nor U17556 (N_17556,N_17290,N_17279);
nor U17557 (N_17557,N_17288,N_17336);
xnor U17558 (N_17558,N_17392,N_17477);
xor U17559 (N_17559,N_17254,N_17491);
and U17560 (N_17560,N_17295,N_17302);
and U17561 (N_17561,N_17473,N_17487);
nor U17562 (N_17562,N_17267,N_17413);
or U17563 (N_17563,N_17457,N_17319);
xnor U17564 (N_17564,N_17345,N_17316);
nand U17565 (N_17565,N_17311,N_17296);
nand U17566 (N_17566,N_17277,N_17416);
nand U17567 (N_17567,N_17370,N_17354);
or U17568 (N_17568,N_17419,N_17445);
xor U17569 (N_17569,N_17367,N_17322);
nor U17570 (N_17570,N_17294,N_17364);
or U17571 (N_17571,N_17389,N_17456);
xnor U17572 (N_17572,N_17460,N_17415);
or U17573 (N_17573,N_17493,N_17346);
nor U17574 (N_17574,N_17329,N_17427);
xnor U17575 (N_17575,N_17264,N_17463);
or U17576 (N_17576,N_17361,N_17353);
xnor U17577 (N_17577,N_17408,N_17292);
or U17578 (N_17578,N_17266,N_17483);
or U17579 (N_17579,N_17358,N_17388);
nor U17580 (N_17580,N_17465,N_17469);
nor U17581 (N_17581,N_17259,N_17363);
nor U17582 (N_17582,N_17452,N_17470);
or U17583 (N_17583,N_17449,N_17299);
xnor U17584 (N_17584,N_17471,N_17374);
nor U17585 (N_17585,N_17280,N_17265);
xnor U17586 (N_17586,N_17429,N_17430);
nor U17587 (N_17587,N_17418,N_17490);
nand U17588 (N_17588,N_17313,N_17281);
xnor U17589 (N_17589,N_17368,N_17301);
nand U17590 (N_17590,N_17481,N_17261);
or U17591 (N_17591,N_17432,N_17381);
nand U17592 (N_17592,N_17378,N_17343);
nand U17593 (N_17593,N_17297,N_17399);
nand U17594 (N_17594,N_17309,N_17455);
and U17595 (N_17595,N_17444,N_17373);
nor U17596 (N_17596,N_17466,N_17379);
xnor U17597 (N_17597,N_17357,N_17498);
and U17598 (N_17598,N_17468,N_17450);
nand U17599 (N_17599,N_17262,N_17371);
xnor U17600 (N_17600,N_17428,N_17489);
nand U17601 (N_17601,N_17404,N_17484);
or U17602 (N_17602,N_17305,N_17447);
nand U17603 (N_17603,N_17474,N_17400);
xnor U17604 (N_17604,N_17318,N_17369);
nor U17605 (N_17605,N_17417,N_17306);
or U17606 (N_17606,N_17453,N_17278);
nand U17607 (N_17607,N_17276,N_17499);
nor U17608 (N_17608,N_17448,N_17375);
xnor U17609 (N_17609,N_17362,N_17284);
nor U17610 (N_17610,N_17342,N_17480);
nor U17611 (N_17611,N_17324,N_17407);
nand U17612 (N_17612,N_17478,N_17272);
and U17613 (N_17613,N_17424,N_17376);
and U17614 (N_17614,N_17451,N_17434);
nand U17615 (N_17615,N_17377,N_17479);
nand U17616 (N_17616,N_17252,N_17298);
and U17617 (N_17617,N_17325,N_17405);
or U17618 (N_17618,N_17317,N_17475);
nand U17619 (N_17619,N_17372,N_17431);
nand U17620 (N_17620,N_17438,N_17482);
xor U17621 (N_17621,N_17341,N_17366);
or U17622 (N_17622,N_17458,N_17383);
or U17623 (N_17623,N_17349,N_17386);
nor U17624 (N_17624,N_17338,N_17332);
xnor U17625 (N_17625,N_17410,N_17293);
nor U17626 (N_17626,N_17397,N_17274);
nand U17627 (N_17627,N_17478,N_17281);
nor U17628 (N_17628,N_17437,N_17398);
xnor U17629 (N_17629,N_17280,N_17357);
nand U17630 (N_17630,N_17377,N_17458);
xor U17631 (N_17631,N_17362,N_17444);
xnor U17632 (N_17632,N_17348,N_17338);
or U17633 (N_17633,N_17337,N_17484);
and U17634 (N_17634,N_17393,N_17311);
or U17635 (N_17635,N_17352,N_17455);
or U17636 (N_17636,N_17307,N_17379);
nand U17637 (N_17637,N_17410,N_17261);
and U17638 (N_17638,N_17321,N_17421);
or U17639 (N_17639,N_17479,N_17313);
or U17640 (N_17640,N_17412,N_17383);
or U17641 (N_17641,N_17316,N_17324);
nor U17642 (N_17642,N_17479,N_17339);
nand U17643 (N_17643,N_17285,N_17389);
and U17644 (N_17644,N_17477,N_17313);
and U17645 (N_17645,N_17279,N_17456);
nor U17646 (N_17646,N_17444,N_17474);
xnor U17647 (N_17647,N_17310,N_17479);
nand U17648 (N_17648,N_17350,N_17462);
nor U17649 (N_17649,N_17325,N_17285);
nor U17650 (N_17650,N_17407,N_17250);
nor U17651 (N_17651,N_17444,N_17357);
and U17652 (N_17652,N_17333,N_17364);
or U17653 (N_17653,N_17468,N_17498);
nand U17654 (N_17654,N_17253,N_17314);
nand U17655 (N_17655,N_17251,N_17279);
nand U17656 (N_17656,N_17286,N_17284);
and U17657 (N_17657,N_17276,N_17326);
xor U17658 (N_17658,N_17336,N_17256);
or U17659 (N_17659,N_17478,N_17279);
and U17660 (N_17660,N_17458,N_17483);
or U17661 (N_17661,N_17341,N_17337);
nand U17662 (N_17662,N_17368,N_17341);
nand U17663 (N_17663,N_17340,N_17407);
xnor U17664 (N_17664,N_17303,N_17455);
nand U17665 (N_17665,N_17335,N_17403);
xnor U17666 (N_17666,N_17497,N_17332);
xnor U17667 (N_17667,N_17337,N_17299);
xnor U17668 (N_17668,N_17325,N_17340);
nor U17669 (N_17669,N_17413,N_17343);
or U17670 (N_17670,N_17315,N_17445);
and U17671 (N_17671,N_17383,N_17266);
xnor U17672 (N_17672,N_17298,N_17460);
or U17673 (N_17673,N_17394,N_17422);
nor U17674 (N_17674,N_17351,N_17320);
xor U17675 (N_17675,N_17375,N_17338);
xnor U17676 (N_17676,N_17296,N_17423);
nor U17677 (N_17677,N_17280,N_17429);
and U17678 (N_17678,N_17404,N_17492);
nand U17679 (N_17679,N_17318,N_17475);
xor U17680 (N_17680,N_17486,N_17273);
nor U17681 (N_17681,N_17459,N_17303);
and U17682 (N_17682,N_17400,N_17476);
or U17683 (N_17683,N_17480,N_17322);
nand U17684 (N_17684,N_17400,N_17464);
nand U17685 (N_17685,N_17329,N_17320);
and U17686 (N_17686,N_17354,N_17303);
or U17687 (N_17687,N_17485,N_17458);
and U17688 (N_17688,N_17385,N_17290);
nor U17689 (N_17689,N_17303,N_17427);
nand U17690 (N_17690,N_17469,N_17499);
or U17691 (N_17691,N_17430,N_17262);
and U17692 (N_17692,N_17429,N_17255);
or U17693 (N_17693,N_17355,N_17250);
xnor U17694 (N_17694,N_17426,N_17267);
or U17695 (N_17695,N_17348,N_17363);
or U17696 (N_17696,N_17348,N_17310);
nor U17697 (N_17697,N_17400,N_17449);
or U17698 (N_17698,N_17386,N_17332);
xnor U17699 (N_17699,N_17491,N_17490);
nand U17700 (N_17700,N_17270,N_17282);
and U17701 (N_17701,N_17441,N_17359);
and U17702 (N_17702,N_17473,N_17378);
or U17703 (N_17703,N_17308,N_17346);
xnor U17704 (N_17704,N_17450,N_17488);
and U17705 (N_17705,N_17338,N_17269);
nand U17706 (N_17706,N_17261,N_17452);
or U17707 (N_17707,N_17252,N_17339);
nand U17708 (N_17708,N_17290,N_17319);
nand U17709 (N_17709,N_17320,N_17420);
nor U17710 (N_17710,N_17434,N_17342);
and U17711 (N_17711,N_17371,N_17376);
xor U17712 (N_17712,N_17300,N_17268);
nand U17713 (N_17713,N_17252,N_17484);
nand U17714 (N_17714,N_17467,N_17318);
nor U17715 (N_17715,N_17334,N_17271);
nor U17716 (N_17716,N_17349,N_17275);
xor U17717 (N_17717,N_17294,N_17403);
nand U17718 (N_17718,N_17357,N_17261);
nor U17719 (N_17719,N_17312,N_17439);
xnor U17720 (N_17720,N_17274,N_17428);
nand U17721 (N_17721,N_17354,N_17281);
or U17722 (N_17722,N_17431,N_17364);
and U17723 (N_17723,N_17497,N_17285);
nor U17724 (N_17724,N_17311,N_17442);
xnor U17725 (N_17725,N_17312,N_17405);
nor U17726 (N_17726,N_17489,N_17387);
xnor U17727 (N_17727,N_17348,N_17257);
xnor U17728 (N_17728,N_17265,N_17308);
or U17729 (N_17729,N_17480,N_17344);
nor U17730 (N_17730,N_17465,N_17262);
nor U17731 (N_17731,N_17274,N_17383);
nor U17732 (N_17732,N_17334,N_17369);
nand U17733 (N_17733,N_17465,N_17463);
or U17734 (N_17734,N_17475,N_17363);
or U17735 (N_17735,N_17329,N_17371);
nand U17736 (N_17736,N_17479,N_17457);
or U17737 (N_17737,N_17284,N_17281);
or U17738 (N_17738,N_17428,N_17288);
xnor U17739 (N_17739,N_17413,N_17348);
and U17740 (N_17740,N_17480,N_17335);
nand U17741 (N_17741,N_17455,N_17463);
xor U17742 (N_17742,N_17391,N_17250);
xnor U17743 (N_17743,N_17405,N_17419);
xnor U17744 (N_17744,N_17336,N_17404);
nor U17745 (N_17745,N_17455,N_17364);
nor U17746 (N_17746,N_17462,N_17363);
xnor U17747 (N_17747,N_17420,N_17329);
nand U17748 (N_17748,N_17254,N_17317);
and U17749 (N_17749,N_17387,N_17497);
nand U17750 (N_17750,N_17594,N_17730);
and U17751 (N_17751,N_17660,N_17627);
nand U17752 (N_17752,N_17620,N_17638);
or U17753 (N_17753,N_17515,N_17682);
nand U17754 (N_17754,N_17602,N_17546);
nand U17755 (N_17755,N_17530,N_17705);
or U17756 (N_17756,N_17510,N_17504);
nor U17757 (N_17757,N_17670,N_17662);
or U17758 (N_17758,N_17625,N_17727);
nor U17759 (N_17759,N_17694,N_17521);
and U17760 (N_17760,N_17563,N_17595);
or U17761 (N_17761,N_17663,N_17724);
and U17762 (N_17762,N_17518,N_17516);
nand U17763 (N_17763,N_17729,N_17544);
nand U17764 (N_17764,N_17676,N_17734);
xor U17765 (N_17765,N_17689,N_17590);
or U17766 (N_17766,N_17613,N_17744);
xnor U17767 (N_17767,N_17511,N_17557);
and U17768 (N_17768,N_17674,N_17731);
nand U17769 (N_17769,N_17747,N_17733);
and U17770 (N_17770,N_17614,N_17720);
nor U17771 (N_17771,N_17577,N_17743);
and U17772 (N_17772,N_17591,N_17574);
nand U17773 (N_17773,N_17713,N_17600);
nand U17774 (N_17774,N_17526,N_17599);
and U17775 (N_17775,N_17560,N_17533);
xnor U17776 (N_17776,N_17582,N_17529);
or U17777 (N_17777,N_17558,N_17605);
nor U17778 (N_17778,N_17646,N_17608);
nor U17779 (N_17779,N_17505,N_17635);
nor U17780 (N_17780,N_17581,N_17508);
and U17781 (N_17781,N_17623,N_17542);
and U17782 (N_17782,N_17622,N_17619);
nand U17783 (N_17783,N_17652,N_17688);
or U17784 (N_17784,N_17711,N_17579);
xnor U17785 (N_17785,N_17710,N_17572);
nor U17786 (N_17786,N_17683,N_17672);
nand U17787 (N_17787,N_17507,N_17725);
nor U17788 (N_17788,N_17653,N_17617);
nor U17789 (N_17789,N_17669,N_17701);
or U17790 (N_17790,N_17547,N_17650);
and U17791 (N_17791,N_17708,N_17715);
or U17792 (N_17792,N_17681,N_17706);
or U17793 (N_17793,N_17666,N_17592);
nor U17794 (N_17794,N_17540,N_17667);
or U17795 (N_17795,N_17555,N_17728);
or U17796 (N_17796,N_17636,N_17722);
or U17797 (N_17797,N_17687,N_17637);
nor U17798 (N_17798,N_17556,N_17584);
and U17799 (N_17799,N_17621,N_17522);
or U17800 (N_17800,N_17746,N_17665);
nand U17801 (N_17801,N_17677,N_17610);
or U17802 (N_17802,N_17580,N_17640);
nand U17803 (N_17803,N_17644,N_17566);
and U17804 (N_17804,N_17598,N_17553);
nand U17805 (N_17805,N_17576,N_17517);
nor U17806 (N_17806,N_17618,N_17639);
nand U17807 (N_17807,N_17723,N_17626);
nand U17808 (N_17808,N_17655,N_17531);
nor U17809 (N_17809,N_17696,N_17587);
nand U17810 (N_17810,N_17632,N_17679);
nor U17811 (N_17811,N_17514,N_17740);
and U17812 (N_17812,N_17718,N_17721);
or U17813 (N_17813,N_17749,N_17695);
nor U17814 (N_17814,N_17741,N_17520);
xor U17815 (N_17815,N_17545,N_17659);
nor U17816 (N_17816,N_17671,N_17543);
nand U17817 (N_17817,N_17630,N_17714);
nand U17818 (N_17818,N_17700,N_17690);
nand U17819 (N_17819,N_17597,N_17702);
nand U17820 (N_17820,N_17704,N_17596);
or U17821 (N_17821,N_17534,N_17513);
or U17822 (N_17822,N_17634,N_17717);
or U17823 (N_17823,N_17719,N_17649);
or U17824 (N_17824,N_17698,N_17707);
nand U17825 (N_17825,N_17548,N_17680);
xor U17826 (N_17826,N_17551,N_17645);
nand U17827 (N_17827,N_17549,N_17528);
nor U17828 (N_17828,N_17541,N_17568);
or U17829 (N_17829,N_17716,N_17732);
or U17830 (N_17830,N_17506,N_17703);
and U17831 (N_17831,N_17564,N_17607);
nor U17832 (N_17832,N_17527,N_17501);
or U17833 (N_17833,N_17668,N_17503);
nor U17834 (N_17834,N_17697,N_17656);
nand U17835 (N_17835,N_17578,N_17647);
nand U17836 (N_17836,N_17524,N_17601);
nor U17837 (N_17837,N_17603,N_17575);
nor U17838 (N_17838,N_17648,N_17738);
xor U17839 (N_17839,N_17745,N_17684);
or U17840 (N_17840,N_17675,N_17693);
xor U17841 (N_17841,N_17737,N_17735);
or U17842 (N_17842,N_17664,N_17519);
or U17843 (N_17843,N_17616,N_17536);
or U17844 (N_17844,N_17552,N_17748);
and U17845 (N_17845,N_17611,N_17609);
xnor U17846 (N_17846,N_17641,N_17538);
xor U17847 (N_17847,N_17525,N_17532);
nand U17848 (N_17848,N_17565,N_17692);
nand U17849 (N_17849,N_17509,N_17523);
xor U17850 (N_17850,N_17726,N_17554);
and U17851 (N_17851,N_17654,N_17570);
xor U17852 (N_17852,N_17661,N_17512);
and U17853 (N_17853,N_17712,N_17651);
nand U17854 (N_17854,N_17657,N_17500);
nand U17855 (N_17855,N_17561,N_17537);
nor U17856 (N_17856,N_17624,N_17691);
and U17857 (N_17857,N_17739,N_17678);
nor U17858 (N_17858,N_17643,N_17742);
nand U17859 (N_17859,N_17583,N_17562);
nor U17860 (N_17860,N_17586,N_17631);
and U17861 (N_17861,N_17585,N_17686);
and U17862 (N_17862,N_17673,N_17628);
xor U17863 (N_17863,N_17567,N_17604);
or U17864 (N_17864,N_17736,N_17539);
and U17865 (N_17865,N_17573,N_17588);
nand U17866 (N_17866,N_17685,N_17593);
xor U17867 (N_17867,N_17559,N_17615);
nand U17868 (N_17868,N_17633,N_17589);
or U17869 (N_17869,N_17535,N_17629);
and U17870 (N_17870,N_17658,N_17550);
nor U17871 (N_17871,N_17571,N_17606);
and U17872 (N_17872,N_17699,N_17709);
xor U17873 (N_17873,N_17612,N_17502);
or U17874 (N_17874,N_17642,N_17569);
nor U17875 (N_17875,N_17735,N_17588);
and U17876 (N_17876,N_17597,N_17677);
nand U17877 (N_17877,N_17595,N_17743);
xor U17878 (N_17878,N_17500,N_17679);
nor U17879 (N_17879,N_17719,N_17735);
and U17880 (N_17880,N_17598,N_17729);
nor U17881 (N_17881,N_17515,N_17710);
xnor U17882 (N_17882,N_17505,N_17607);
nor U17883 (N_17883,N_17556,N_17616);
and U17884 (N_17884,N_17661,N_17677);
nand U17885 (N_17885,N_17729,N_17663);
nor U17886 (N_17886,N_17630,N_17615);
and U17887 (N_17887,N_17551,N_17709);
and U17888 (N_17888,N_17666,N_17670);
nor U17889 (N_17889,N_17627,N_17727);
and U17890 (N_17890,N_17654,N_17503);
and U17891 (N_17891,N_17682,N_17640);
xnor U17892 (N_17892,N_17524,N_17650);
or U17893 (N_17893,N_17645,N_17577);
xnor U17894 (N_17894,N_17501,N_17623);
nand U17895 (N_17895,N_17702,N_17584);
nand U17896 (N_17896,N_17709,N_17621);
nand U17897 (N_17897,N_17524,N_17682);
or U17898 (N_17898,N_17705,N_17562);
xor U17899 (N_17899,N_17732,N_17737);
and U17900 (N_17900,N_17549,N_17712);
or U17901 (N_17901,N_17611,N_17620);
and U17902 (N_17902,N_17652,N_17742);
nor U17903 (N_17903,N_17685,N_17518);
xnor U17904 (N_17904,N_17740,N_17526);
nor U17905 (N_17905,N_17740,N_17550);
or U17906 (N_17906,N_17516,N_17501);
nand U17907 (N_17907,N_17504,N_17707);
or U17908 (N_17908,N_17548,N_17685);
or U17909 (N_17909,N_17612,N_17645);
nand U17910 (N_17910,N_17715,N_17594);
xnor U17911 (N_17911,N_17580,N_17718);
nor U17912 (N_17912,N_17530,N_17745);
or U17913 (N_17913,N_17658,N_17557);
or U17914 (N_17914,N_17706,N_17544);
and U17915 (N_17915,N_17697,N_17740);
xor U17916 (N_17916,N_17531,N_17588);
or U17917 (N_17917,N_17520,N_17542);
xnor U17918 (N_17918,N_17669,N_17538);
nor U17919 (N_17919,N_17670,N_17642);
or U17920 (N_17920,N_17519,N_17568);
xnor U17921 (N_17921,N_17727,N_17671);
or U17922 (N_17922,N_17584,N_17565);
xnor U17923 (N_17923,N_17537,N_17725);
nor U17924 (N_17924,N_17579,N_17558);
nand U17925 (N_17925,N_17522,N_17559);
xnor U17926 (N_17926,N_17567,N_17518);
nor U17927 (N_17927,N_17645,N_17636);
xor U17928 (N_17928,N_17632,N_17672);
or U17929 (N_17929,N_17680,N_17605);
and U17930 (N_17930,N_17534,N_17640);
nor U17931 (N_17931,N_17735,N_17651);
or U17932 (N_17932,N_17733,N_17701);
or U17933 (N_17933,N_17716,N_17639);
xor U17934 (N_17934,N_17712,N_17609);
and U17935 (N_17935,N_17592,N_17571);
and U17936 (N_17936,N_17724,N_17507);
or U17937 (N_17937,N_17617,N_17747);
and U17938 (N_17938,N_17745,N_17636);
xnor U17939 (N_17939,N_17563,N_17746);
and U17940 (N_17940,N_17694,N_17713);
nand U17941 (N_17941,N_17507,N_17661);
nand U17942 (N_17942,N_17526,N_17500);
or U17943 (N_17943,N_17554,N_17545);
nor U17944 (N_17944,N_17718,N_17701);
or U17945 (N_17945,N_17520,N_17666);
xor U17946 (N_17946,N_17685,N_17735);
nand U17947 (N_17947,N_17649,N_17584);
nor U17948 (N_17948,N_17640,N_17681);
nand U17949 (N_17949,N_17630,N_17688);
nor U17950 (N_17950,N_17745,N_17507);
and U17951 (N_17951,N_17561,N_17611);
or U17952 (N_17952,N_17575,N_17693);
nand U17953 (N_17953,N_17669,N_17648);
and U17954 (N_17954,N_17540,N_17561);
xnor U17955 (N_17955,N_17501,N_17665);
or U17956 (N_17956,N_17600,N_17699);
xor U17957 (N_17957,N_17567,N_17577);
xnor U17958 (N_17958,N_17665,N_17543);
nor U17959 (N_17959,N_17613,N_17582);
nor U17960 (N_17960,N_17703,N_17631);
nand U17961 (N_17961,N_17541,N_17594);
or U17962 (N_17962,N_17579,N_17695);
nor U17963 (N_17963,N_17721,N_17619);
xnor U17964 (N_17964,N_17579,N_17746);
or U17965 (N_17965,N_17726,N_17703);
and U17966 (N_17966,N_17619,N_17558);
or U17967 (N_17967,N_17606,N_17569);
and U17968 (N_17968,N_17554,N_17669);
and U17969 (N_17969,N_17698,N_17671);
xor U17970 (N_17970,N_17707,N_17638);
or U17971 (N_17971,N_17707,N_17628);
or U17972 (N_17972,N_17633,N_17557);
xor U17973 (N_17973,N_17567,N_17721);
and U17974 (N_17974,N_17654,N_17727);
nor U17975 (N_17975,N_17636,N_17589);
xor U17976 (N_17976,N_17524,N_17629);
nand U17977 (N_17977,N_17578,N_17590);
nand U17978 (N_17978,N_17518,N_17574);
or U17979 (N_17979,N_17631,N_17665);
xnor U17980 (N_17980,N_17626,N_17589);
nand U17981 (N_17981,N_17630,N_17687);
nor U17982 (N_17982,N_17707,N_17667);
nand U17983 (N_17983,N_17692,N_17717);
nor U17984 (N_17984,N_17700,N_17674);
or U17985 (N_17985,N_17699,N_17695);
nor U17986 (N_17986,N_17525,N_17509);
and U17987 (N_17987,N_17666,N_17587);
or U17988 (N_17988,N_17511,N_17521);
xnor U17989 (N_17989,N_17536,N_17735);
nor U17990 (N_17990,N_17526,N_17717);
nor U17991 (N_17991,N_17542,N_17687);
and U17992 (N_17992,N_17612,N_17687);
or U17993 (N_17993,N_17744,N_17578);
and U17994 (N_17994,N_17624,N_17545);
and U17995 (N_17995,N_17541,N_17551);
nand U17996 (N_17996,N_17640,N_17655);
nor U17997 (N_17997,N_17736,N_17685);
nand U17998 (N_17998,N_17700,N_17701);
and U17999 (N_17999,N_17528,N_17721);
or U18000 (N_18000,N_17968,N_17873);
nand U18001 (N_18001,N_17964,N_17905);
xor U18002 (N_18002,N_17833,N_17845);
xor U18003 (N_18003,N_17755,N_17894);
nor U18004 (N_18004,N_17859,N_17960);
and U18005 (N_18005,N_17784,N_17796);
nor U18006 (N_18006,N_17813,N_17983);
nor U18007 (N_18007,N_17935,N_17972);
or U18008 (N_18008,N_17950,N_17778);
or U18009 (N_18009,N_17947,N_17812);
and U18010 (N_18010,N_17849,N_17787);
nor U18011 (N_18011,N_17830,N_17760);
nor U18012 (N_18012,N_17906,N_17998);
nand U18013 (N_18013,N_17761,N_17896);
nor U18014 (N_18014,N_17893,N_17752);
nand U18015 (N_18015,N_17821,N_17908);
or U18016 (N_18016,N_17993,N_17865);
and U18017 (N_18017,N_17802,N_17772);
xor U18018 (N_18018,N_17892,N_17939);
nand U18019 (N_18019,N_17858,N_17995);
nand U18020 (N_18020,N_17801,N_17878);
nand U18021 (N_18021,N_17882,N_17827);
nand U18022 (N_18022,N_17957,N_17879);
and U18023 (N_18023,N_17980,N_17840);
or U18024 (N_18024,N_17822,N_17829);
nand U18025 (N_18025,N_17867,N_17852);
and U18026 (N_18026,N_17977,N_17843);
and U18027 (N_18027,N_17994,N_17814);
and U18028 (N_18028,N_17792,N_17958);
or U18029 (N_18029,N_17953,N_17954);
xnor U18030 (N_18030,N_17756,N_17970);
nand U18031 (N_18031,N_17911,N_17959);
nand U18032 (N_18032,N_17770,N_17955);
xnor U18033 (N_18033,N_17769,N_17810);
xor U18034 (N_18034,N_17971,N_17860);
or U18035 (N_18035,N_17899,N_17823);
and U18036 (N_18036,N_17976,N_17777);
or U18037 (N_18037,N_17890,N_17969);
and U18038 (N_18038,N_17779,N_17961);
nor U18039 (N_18039,N_17923,N_17788);
or U18040 (N_18040,N_17759,N_17811);
xnor U18041 (N_18041,N_17921,N_17790);
xor U18042 (N_18042,N_17985,N_17825);
and U18043 (N_18043,N_17835,N_17758);
nand U18044 (N_18044,N_17984,N_17864);
nand U18045 (N_18045,N_17832,N_17986);
xnor U18046 (N_18046,N_17773,N_17938);
and U18047 (N_18047,N_17774,N_17952);
and U18048 (N_18048,N_17862,N_17848);
or U18049 (N_18049,N_17987,N_17880);
xnor U18050 (N_18050,N_17978,N_17928);
nand U18051 (N_18051,N_17951,N_17926);
or U18052 (N_18052,N_17871,N_17751);
and U18053 (N_18053,N_17791,N_17850);
nor U18054 (N_18054,N_17956,N_17824);
or U18055 (N_18055,N_17780,N_17803);
nor U18056 (N_18056,N_17988,N_17750);
or U18057 (N_18057,N_17883,N_17974);
and U18058 (N_18058,N_17909,N_17889);
xor U18059 (N_18059,N_17925,N_17929);
or U18060 (N_18060,N_17819,N_17967);
xor U18061 (N_18061,N_17794,N_17945);
xor U18062 (N_18062,N_17886,N_17920);
nor U18063 (N_18063,N_17913,N_17838);
and U18064 (N_18064,N_17931,N_17965);
and U18065 (N_18065,N_17839,N_17818);
nor U18066 (N_18066,N_17762,N_17775);
or U18067 (N_18067,N_17948,N_17876);
nor U18068 (N_18068,N_17903,N_17863);
nand U18069 (N_18069,N_17932,N_17834);
and U18070 (N_18070,N_17897,N_17870);
nor U18071 (N_18071,N_17875,N_17884);
or U18072 (N_18072,N_17765,N_17927);
or U18073 (N_18073,N_17895,N_17866);
and U18074 (N_18074,N_17981,N_17910);
xnor U18075 (N_18075,N_17898,N_17855);
nand U18076 (N_18076,N_17754,N_17874);
nand U18077 (N_18077,N_17949,N_17782);
nand U18078 (N_18078,N_17776,N_17789);
or U18079 (N_18079,N_17842,N_17937);
nand U18080 (N_18080,N_17912,N_17943);
nor U18081 (N_18081,N_17936,N_17861);
xnor U18082 (N_18082,N_17992,N_17800);
or U18083 (N_18083,N_17805,N_17795);
and U18084 (N_18084,N_17919,N_17856);
and U18085 (N_18085,N_17817,N_17900);
and U18086 (N_18086,N_17804,N_17902);
or U18087 (N_18087,N_17885,N_17806);
nor U18088 (N_18088,N_17922,N_17914);
xor U18089 (N_18089,N_17815,N_17826);
nand U18090 (N_18090,N_17973,N_17844);
xor U18091 (N_18091,N_17793,N_17888);
nor U18092 (N_18092,N_17996,N_17753);
and U18093 (N_18093,N_17851,N_17757);
nand U18094 (N_18094,N_17877,N_17836);
or U18095 (N_18095,N_17767,N_17915);
nor U18096 (N_18096,N_17997,N_17887);
xnor U18097 (N_18097,N_17828,N_17963);
and U18098 (N_18098,N_17869,N_17771);
or U18099 (N_18099,N_17891,N_17868);
nand U18100 (N_18100,N_17941,N_17807);
nor U18101 (N_18101,N_17831,N_17846);
nor U18102 (N_18102,N_17966,N_17904);
nor U18103 (N_18103,N_17847,N_17930);
nor U18104 (N_18104,N_17797,N_17854);
nand U18105 (N_18105,N_17901,N_17857);
xor U18106 (N_18106,N_17940,N_17763);
and U18107 (N_18107,N_17820,N_17917);
xor U18108 (N_18108,N_17809,N_17946);
nor U18109 (N_18109,N_17918,N_17881);
or U18110 (N_18110,N_17916,N_17907);
nand U18111 (N_18111,N_17783,N_17837);
nor U18112 (N_18112,N_17989,N_17962);
nor U18113 (N_18113,N_17764,N_17768);
nand U18114 (N_18114,N_17979,N_17934);
nor U18115 (N_18115,N_17841,N_17991);
or U18116 (N_18116,N_17942,N_17816);
xnor U18117 (N_18117,N_17808,N_17990);
and U18118 (N_18118,N_17853,N_17999);
or U18119 (N_18119,N_17799,N_17766);
nand U18120 (N_18120,N_17781,N_17944);
nand U18121 (N_18121,N_17924,N_17982);
nand U18122 (N_18122,N_17785,N_17872);
nand U18123 (N_18123,N_17975,N_17933);
or U18124 (N_18124,N_17786,N_17798);
or U18125 (N_18125,N_17894,N_17952);
or U18126 (N_18126,N_17787,N_17812);
nand U18127 (N_18127,N_17796,N_17865);
or U18128 (N_18128,N_17898,N_17991);
nand U18129 (N_18129,N_17900,N_17820);
nor U18130 (N_18130,N_17885,N_17932);
xnor U18131 (N_18131,N_17904,N_17968);
and U18132 (N_18132,N_17967,N_17830);
xnor U18133 (N_18133,N_17883,N_17908);
or U18134 (N_18134,N_17863,N_17832);
nor U18135 (N_18135,N_17751,N_17760);
nor U18136 (N_18136,N_17802,N_17921);
xor U18137 (N_18137,N_17992,N_17946);
or U18138 (N_18138,N_17951,N_17802);
and U18139 (N_18139,N_17959,N_17966);
nand U18140 (N_18140,N_17797,N_17940);
and U18141 (N_18141,N_17885,N_17831);
and U18142 (N_18142,N_17930,N_17796);
nand U18143 (N_18143,N_17795,N_17983);
xor U18144 (N_18144,N_17760,N_17856);
xor U18145 (N_18145,N_17824,N_17862);
nand U18146 (N_18146,N_17755,N_17953);
or U18147 (N_18147,N_17793,N_17829);
xnor U18148 (N_18148,N_17934,N_17831);
nand U18149 (N_18149,N_17919,N_17845);
or U18150 (N_18150,N_17758,N_17868);
nand U18151 (N_18151,N_17797,N_17895);
nor U18152 (N_18152,N_17956,N_17998);
nand U18153 (N_18153,N_17853,N_17844);
nand U18154 (N_18154,N_17941,N_17903);
xor U18155 (N_18155,N_17873,N_17870);
and U18156 (N_18156,N_17938,N_17827);
nand U18157 (N_18157,N_17781,N_17832);
or U18158 (N_18158,N_17925,N_17901);
and U18159 (N_18159,N_17942,N_17966);
and U18160 (N_18160,N_17963,N_17780);
nand U18161 (N_18161,N_17955,N_17813);
nand U18162 (N_18162,N_17778,N_17760);
nor U18163 (N_18163,N_17965,N_17791);
or U18164 (N_18164,N_17906,N_17780);
nand U18165 (N_18165,N_17936,N_17843);
nor U18166 (N_18166,N_17916,N_17829);
xor U18167 (N_18167,N_17931,N_17907);
and U18168 (N_18168,N_17798,N_17934);
and U18169 (N_18169,N_17862,N_17867);
nor U18170 (N_18170,N_17967,N_17838);
and U18171 (N_18171,N_17933,N_17881);
xnor U18172 (N_18172,N_17932,N_17978);
nor U18173 (N_18173,N_17854,N_17782);
xor U18174 (N_18174,N_17976,N_17802);
or U18175 (N_18175,N_17930,N_17912);
nand U18176 (N_18176,N_17977,N_17969);
xnor U18177 (N_18177,N_17925,N_17922);
or U18178 (N_18178,N_17787,N_17766);
and U18179 (N_18179,N_17849,N_17848);
or U18180 (N_18180,N_17758,N_17752);
nand U18181 (N_18181,N_17927,N_17922);
nand U18182 (N_18182,N_17827,N_17788);
xnor U18183 (N_18183,N_17902,N_17896);
xor U18184 (N_18184,N_17996,N_17968);
or U18185 (N_18185,N_17971,N_17981);
xor U18186 (N_18186,N_17959,N_17768);
nor U18187 (N_18187,N_17794,N_17971);
nor U18188 (N_18188,N_17850,N_17952);
nor U18189 (N_18189,N_17755,N_17836);
nand U18190 (N_18190,N_17849,N_17780);
and U18191 (N_18191,N_17839,N_17763);
nand U18192 (N_18192,N_17826,N_17851);
and U18193 (N_18193,N_17992,N_17750);
xnor U18194 (N_18194,N_17867,N_17907);
or U18195 (N_18195,N_17774,N_17973);
or U18196 (N_18196,N_17902,N_17824);
nor U18197 (N_18197,N_17787,N_17922);
xor U18198 (N_18198,N_17805,N_17910);
and U18199 (N_18199,N_17811,N_17998);
and U18200 (N_18200,N_17853,N_17885);
nor U18201 (N_18201,N_17992,N_17801);
and U18202 (N_18202,N_17751,N_17997);
and U18203 (N_18203,N_17777,N_17859);
nor U18204 (N_18204,N_17910,N_17952);
xor U18205 (N_18205,N_17798,N_17981);
or U18206 (N_18206,N_17854,N_17789);
or U18207 (N_18207,N_17956,N_17974);
and U18208 (N_18208,N_17911,N_17815);
nand U18209 (N_18209,N_17872,N_17765);
or U18210 (N_18210,N_17883,N_17973);
nand U18211 (N_18211,N_17986,N_17915);
nand U18212 (N_18212,N_17925,N_17763);
xor U18213 (N_18213,N_17838,N_17953);
nor U18214 (N_18214,N_17836,N_17940);
or U18215 (N_18215,N_17911,N_17787);
or U18216 (N_18216,N_17897,N_17979);
nor U18217 (N_18217,N_17877,N_17837);
or U18218 (N_18218,N_17929,N_17753);
nor U18219 (N_18219,N_17979,N_17957);
xor U18220 (N_18220,N_17925,N_17762);
nor U18221 (N_18221,N_17764,N_17803);
or U18222 (N_18222,N_17988,N_17880);
or U18223 (N_18223,N_17917,N_17928);
nor U18224 (N_18224,N_17760,N_17867);
xor U18225 (N_18225,N_17895,N_17795);
xnor U18226 (N_18226,N_17789,N_17754);
nand U18227 (N_18227,N_17846,N_17783);
or U18228 (N_18228,N_17876,N_17815);
and U18229 (N_18229,N_17946,N_17915);
xor U18230 (N_18230,N_17986,N_17980);
or U18231 (N_18231,N_17806,N_17867);
nand U18232 (N_18232,N_17787,N_17800);
and U18233 (N_18233,N_17761,N_17973);
xor U18234 (N_18234,N_17896,N_17900);
or U18235 (N_18235,N_17847,N_17807);
nand U18236 (N_18236,N_17762,N_17986);
or U18237 (N_18237,N_17946,N_17943);
nand U18238 (N_18238,N_17797,N_17881);
or U18239 (N_18239,N_17868,N_17980);
nand U18240 (N_18240,N_17903,N_17953);
or U18241 (N_18241,N_17910,N_17785);
nor U18242 (N_18242,N_17944,N_17809);
nand U18243 (N_18243,N_17786,N_17825);
nor U18244 (N_18244,N_17766,N_17865);
xor U18245 (N_18245,N_17810,N_17850);
and U18246 (N_18246,N_17928,N_17927);
or U18247 (N_18247,N_17940,N_17851);
and U18248 (N_18248,N_17994,N_17866);
nand U18249 (N_18249,N_17809,N_17952);
or U18250 (N_18250,N_18044,N_18072);
nor U18251 (N_18251,N_18127,N_18216);
or U18252 (N_18252,N_18215,N_18244);
nand U18253 (N_18253,N_18219,N_18008);
xor U18254 (N_18254,N_18033,N_18227);
or U18255 (N_18255,N_18161,N_18026);
or U18256 (N_18256,N_18193,N_18014);
nor U18257 (N_18257,N_18240,N_18200);
and U18258 (N_18258,N_18147,N_18126);
or U18259 (N_18259,N_18144,N_18197);
nor U18260 (N_18260,N_18025,N_18209);
xnor U18261 (N_18261,N_18097,N_18217);
nand U18262 (N_18262,N_18043,N_18162);
nor U18263 (N_18263,N_18140,N_18007);
and U18264 (N_18264,N_18153,N_18202);
xnor U18265 (N_18265,N_18168,N_18213);
xor U18266 (N_18266,N_18089,N_18045);
nor U18267 (N_18267,N_18034,N_18011);
nand U18268 (N_18268,N_18064,N_18024);
nand U18269 (N_18269,N_18165,N_18015);
and U18270 (N_18270,N_18092,N_18074);
or U18271 (N_18271,N_18048,N_18096);
and U18272 (N_18272,N_18194,N_18159);
or U18273 (N_18273,N_18171,N_18116);
xor U18274 (N_18274,N_18190,N_18241);
and U18275 (N_18275,N_18204,N_18038);
or U18276 (N_18276,N_18141,N_18223);
or U18277 (N_18277,N_18136,N_18146);
nor U18278 (N_18278,N_18139,N_18125);
xor U18279 (N_18279,N_18201,N_18207);
or U18280 (N_18280,N_18110,N_18176);
or U18281 (N_18281,N_18067,N_18137);
or U18282 (N_18282,N_18128,N_18001);
xnor U18283 (N_18283,N_18095,N_18138);
nand U18284 (N_18284,N_18065,N_18199);
nor U18285 (N_18285,N_18177,N_18221);
or U18286 (N_18286,N_18247,N_18013);
nand U18287 (N_18287,N_18224,N_18233);
nor U18288 (N_18288,N_18101,N_18087);
and U18289 (N_18289,N_18052,N_18068);
xor U18290 (N_18290,N_18090,N_18218);
nor U18291 (N_18291,N_18053,N_18031);
xnor U18292 (N_18292,N_18169,N_18054);
and U18293 (N_18293,N_18086,N_18027);
nand U18294 (N_18294,N_18061,N_18149);
or U18295 (N_18295,N_18220,N_18238);
nand U18296 (N_18296,N_18131,N_18022);
and U18297 (N_18297,N_18040,N_18205);
and U18298 (N_18298,N_18198,N_18206);
and U18299 (N_18299,N_18214,N_18192);
or U18300 (N_18300,N_18155,N_18000);
nand U18301 (N_18301,N_18021,N_18010);
and U18302 (N_18302,N_18157,N_18212);
nand U18303 (N_18303,N_18041,N_18173);
nand U18304 (N_18304,N_18150,N_18099);
nand U18305 (N_18305,N_18123,N_18106);
nand U18306 (N_18306,N_18183,N_18049);
xor U18307 (N_18307,N_18180,N_18191);
nor U18308 (N_18308,N_18167,N_18081);
nand U18309 (N_18309,N_18170,N_18036);
nor U18310 (N_18310,N_18058,N_18166);
xor U18311 (N_18311,N_18047,N_18175);
nand U18312 (N_18312,N_18181,N_18222);
nand U18313 (N_18313,N_18164,N_18226);
nand U18314 (N_18314,N_18046,N_18069);
nand U18315 (N_18315,N_18182,N_18083);
and U18316 (N_18316,N_18103,N_18077);
and U18317 (N_18317,N_18249,N_18225);
nor U18318 (N_18318,N_18179,N_18245);
or U18319 (N_18319,N_18108,N_18084);
or U18320 (N_18320,N_18028,N_18109);
nor U18321 (N_18321,N_18154,N_18093);
or U18322 (N_18322,N_18080,N_18237);
and U18323 (N_18323,N_18210,N_18035);
nand U18324 (N_18324,N_18232,N_18019);
nor U18325 (N_18325,N_18060,N_18009);
and U18326 (N_18326,N_18134,N_18023);
and U18327 (N_18327,N_18102,N_18057);
nor U18328 (N_18328,N_18230,N_18196);
xor U18329 (N_18329,N_18235,N_18188);
nor U18330 (N_18330,N_18094,N_18071);
xnor U18331 (N_18331,N_18078,N_18012);
or U18332 (N_18332,N_18018,N_18195);
xnor U18333 (N_18333,N_18063,N_18130);
nor U18334 (N_18334,N_18148,N_18005);
and U18335 (N_18335,N_18158,N_18051);
and U18336 (N_18336,N_18187,N_18120);
nand U18337 (N_18337,N_18133,N_18020);
or U18338 (N_18338,N_18231,N_18234);
or U18339 (N_18339,N_18152,N_18107);
and U18340 (N_18340,N_18059,N_18211);
nand U18341 (N_18341,N_18104,N_18124);
and U18342 (N_18342,N_18085,N_18032);
xnor U18343 (N_18343,N_18088,N_18143);
xor U18344 (N_18344,N_18062,N_18055);
nor U18345 (N_18345,N_18016,N_18135);
nor U18346 (N_18346,N_18174,N_18242);
nand U18347 (N_18347,N_18243,N_18163);
and U18348 (N_18348,N_18186,N_18098);
xor U18349 (N_18349,N_18037,N_18075);
nand U18350 (N_18350,N_18017,N_18050);
or U18351 (N_18351,N_18172,N_18105);
nor U18352 (N_18352,N_18076,N_18042);
nand U18353 (N_18353,N_18208,N_18119);
or U18354 (N_18354,N_18079,N_18006);
or U18355 (N_18355,N_18073,N_18132);
or U18356 (N_18356,N_18070,N_18030);
xor U18357 (N_18357,N_18114,N_18003);
xnor U18358 (N_18358,N_18115,N_18112);
xnor U18359 (N_18359,N_18156,N_18142);
xor U18360 (N_18360,N_18121,N_18246);
nor U18361 (N_18361,N_18002,N_18239);
or U18362 (N_18362,N_18189,N_18228);
nor U18363 (N_18363,N_18039,N_18145);
nor U18364 (N_18364,N_18118,N_18111);
nand U18365 (N_18365,N_18004,N_18236);
and U18366 (N_18366,N_18117,N_18178);
or U18367 (N_18367,N_18091,N_18185);
and U18368 (N_18368,N_18029,N_18056);
nor U18369 (N_18369,N_18151,N_18066);
or U18370 (N_18370,N_18184,N_18248);
or U18371 (N_18371,N_18129,N_18203);
and U18372 (N_18372,N_18229,N_18082);
nand U18373 (N_18373,N_18160,N_18100);
xor U18374 (N_18374,N_18113,N_18122);
xnor U18375 (N_18375,N_18212,N_18198);
and U18376 (N_18376,N_18107,N_18233);
nand U18377 (N_18377,N_18171,N_18218);
xnor U18378 (N_18378,N_18049,N_18003);
nand U18379 (N_18379,N_18197,N_18099);
and U18380 (N_18380,N_18134,N_18248);
xor U18381 (N_18381,N_18201,N_18225);
and U18382 (N_18382,N_18176,N_18198);
or U18383 (N_18383,N_18096,N_18074);
or U18384 (N_18384,N_18016,N_18180);
nor U18385 (N_18385,N_18231,N_18224);
or U18386 (N_18386,N_18110,N_18124);
nor U18387 (N_18387,N_18033,N_18110);
xnor U18388 (N_18388,N_18065,N_18084);
xnor U18389 (N_18389,N_18060,N_18160);
and U18390 (N_18390,N_18198,N_18148);
nor U18391 (N_18391,N_18092,N_18165);
xnor U18392 (N_18392,N_18102,N_18178);
xnor U18393 (N_18393,N_18004,N_18205);
nor U18394 (N_18394,N_18219,N_18014);
and U18395 (N_18395,N_18152,N_18044);
nand U18396 (N_18396,N_18075,N_18031);
or U18397 (N_18397,N_18042,N_18217);
or U18398 (N_18398,N_18234,N_18083);
nand U18399 (N_18399,N_18159,N_18033);
and U18400 (N_18400,N_18020,N_18191);
and U18401 (N_18401,N_18041,N_18156);
xnor U18402 (N_18402,N_18183,N_18162);
and U18403 (N_18403,N_18164,N_18209);
nand U18404 (N_18404,N_18027,N_18170);
nand U18405 (N_18405,N_18000,N_18173);
or U18406 (N_18406,N_18226,N_18163);
and U18407 (N_18407,N_18229,N_18002);
or U18408 (N_18408,N_18220,N_18003);
or U18409 (N_18409,N_18130,N_18090);
nor U18410 (N_18410,N_18178,N_18051);
nand U18411 (N_18411,N_18214,N_18112);
nand U18412 (N_18412,N_18143,N_18165);
or U18413 (N_18413,N_18203,N_18123);
nor U18414 (N_18414,N_18035,N_18239);
or U18415 (N_18415,N_18149,N_18193);
or U18416 (N_18416,N_18047,N_18127);
or U18417 (N_18417,N_18068,N_18096);
and U18418 (N_18418,N_18245,N_18088);
and U18419 (N_18419,N_18139,N_18127);
nor U18420 (N_18420,N_18096,N_18142);
nand U18421 (N_18421,N_18131,N_18018);
xnor U18422 (N_18422,N_18050,N_18135);
or U18423 (N_18423,N_18248,N_18130);
and U18424 (N_18424,N_18015,N_18156);
and U18425 (N_18425,N_18049,N_18225);
nor U18426 (N_18426,N_18075,N_18063);
nand U18427 (N_18427,N_18171,N_18173);
or U18428 (N_18428,N_18221,N_18106);
nand U18429 (N_18429,N_18026,N_18031);
nand U18430 (N_18430,N_18042,N_18000);
or U18431 (N_18431,N_18123,N_18003);
nor U18432 (N_18432,N_18245,N_18055);
nand U18433 (N_18433,N_18206,N_18171);
xor U18434 (N_18434,N_18070,N_18116);
nand U18435 (N_18435,N_18029,N_18227);
nor U18436 (N_18436,N_18235,N_18125);
nand U18437 (N_18437,N_18069,N_18154);
nand U18438 (N_18438,N_18040,N_18091);
xor U18439 (N_18439,N_18221,N_18212);
nor U18440 (N_18440,N_18110,N_18197);
xnor U18441 (N_18441,N_18106,N_18131);
or U18442 (N_18442,N_18233,N_18080);
or U18443 (N_18443,N_18160,N_18198);
nor U18444 (N_18444,N_18070,N_18169);
or U18445 (N_18445,N_18143,N_18098);
nand U18446 (N_18446,N_18160,N_18106);
nand U18447 (N_18447,N_18176,N_18001);
nor U18448 (N_18448,N_18141,N_18145);
and U18449 (N_18449,N_18043,N_18166);
nand U18450 (N_18450,N_18018,N_18063);
and U18451 (N_18451,N_18195,N_18227);
nand U18452 (N_18452,N_18024,N_18246);
or U18453 (N_18453,N_18147,N_18166);
xnor U18454 (N_18454,N_18108,N_18087);
xnor U18455 (N_18455,N_18153,N_18055);
xor U18456 (N_18456,N_18021,N_18161);
nand U18457 (N_18457,N_18059,N_18044);
xor U18458 (N_18458,N_18136,N_18236);
and U18459 (N_18459,N_18032,N_18013);
and U18460 (N_18460,N_18248,N_18099);
nand U18461 (N_18461,N_18089,N_18141);
nor U18462 (N_18462,N_18082,N_18167);
xor U18463 (N_18463,N_18036,N_18231);
nor U18464 (N_18464,N_18224,N_18161);
xor U18465 (N_18465,N_18029,N_18243);
xnor U18466 (N_18466,N_18248,N_18006);
or U18467 (N_18467,N_18233,N_18060);
or U18468 (N_18468,N_18106,N_18219);
or U18469 (N_18469,N_18197,N_18037);
nand U18470 (N_18470,N_18021,N_18154);
nand U18471 (N_18471,N_18205,N_18241);
and U18472 (N_18472,N_18019,N_18149);
xor U18473 (N_18473,N_18192,N_18026);
nor U18474 (N_18474,N_18004,N_18164);
nor U18475 (N_18475,N_18171,N_18026);
or U18476 (N_18476,N_18015,N_18046);
xnor U18477 (N_18477,N_18048,N_18192);
and U18478 (N_18478,N_18199,N_18034);
or U18479 (N_18479,N_18164,N_18199);
or U18480 (N_18480,N_18122,N_18094);
xnor U18481 (N_18481,N_18141,N_18110);
nor U18482 (N_18482,N_18122,N_18085);
or U18483 (N_18483,N_18247,N_18194);
and U18484 (N_18484,N_18138,N_18131);
nor U18485 (N_18485,N_18136,N_18150);
nor U18486 (N_18486,N_18013,N_18132);
xnor U18487 (N_18487,N_18242,N_18246);
nor U18488 (N_18488,N_18098,N_18122);
and U18489 (N_18489,N_18130,N_18037);
xnor U18490 (N_18490,N_18015,N_18076);
or U18491 (N_18491,N_18126,N_18170);
or U18492 (N_18492,N_18121,N_18062);
xnor U18493 (N_18493,N_18167,N_18017);
or U18494 (N_18494,N_18082,N_18192);
nor U18495 (N_18495,N_18035,N_18141);
nand U18496 (N_18496,N_18055,N_18108);
nand U18497 (N_18497,N_18145,N_18233);
nand U18498 (N_18498,N_18167,N_18042);
xnor U18499 (N_18499,N_18079,N_18200);
nor U18500 (N_18500,N_18427,N_18385);
and U18501 (N_18501,N_18386,N_18281);
and U18502 (N_18502,N_18345,N_18415);
nor U18503 (N_18503,N_18474,N_18397);
and U18504 (N_18504,N_18380,N_18424);
nor U18505 (N_18505,N_18387,N_18264);
and U18506 (N_18506,N_18352,N_18443);
nand U18507 (N_18507,N_18362,N_18355);
nor U18508 (N_18508,N_18425,N_18325);
nor U18509 (N_18509,N_18261,N_18278);
or U18510 (N_18510,N_18310,N_18480);
xor U18511 (N_18511,N_18250,N_18426);
and U18512 (N_18512,N_18360,N_18406);
xor U18513 (N_18513,N_18407,N_18453);
or U18514 (N_18514,N_18495,N_18297);
or U18515 (N_18515,N_18314,N_18470);
and U18516 (N_18516,N_18321,N_18370);
xnor U18517 (N_18517,N_18464,N_18266);
or U18518 (N_18518,N_18330,N_18296);
nor U18519 (N_18519,N_18322,N_18458);
nand U18520 (N_18520,N_18326,N_18409);
nor U18521 (N_18521,N_18431,N_18399);
nor U18522 (N_18522,N_18350,N_18364);
xnor U18523 (N_18523,N_18492,N_18294);
and U18524 (N_18524,N_18391,N_18320);
or U18525 (N_18525,N_18469,N_18371);
nand U18526 (N_18526,N_18252,N_18462);
nor U18527 (N_18527,N_18339,N_18289);
xor U18528 (N_18528,N_18319,N_18260);
nand U18529 (N_18529,N_18412,N_18288);
xor U18530 (N_18530,N_18335,N_18304);
or U18531 (N_18531,N_18276,N_18490);
and U18532 (N_18532,N_18340,N_18446);
xor U18533 (N_18533,N_18465,N_18479);
nand U18534 (N_18534,N_18299,N_18444);
and U18535 (N_18535,N_18405,N_18253);
nor U18536 (N_18536,N_18318,N_18308);
and U18537 (N_18537,N_18302,N_18344);
nor U18538 (N_18538,N_18393,N_18270);
or U18539 (N_18539,N_18347,N_18494);
nand U18540 (N_18540,N_18417,N_18259);
nand U18541 (N_18541,N_18284,N_18400);
or U18542 (N_18542,N_18373,N_18434);
and U18543 (N_18543,N_18354,N_18287);
nor U18544 (N_18544,N_18309,N_18333);
xor U18545 (N_18545,N_18324,N_18413);
xnor U18546 (N_18546,N_18461,N_18483);
nand U18547 (N_18547,N_18430,N_18428);
nor U18548 (N_18548,N_18481,N_18251);
xor U18549 (N_18549,N_18376,N_18312);
or U18550 (N_18550,N_18291,N_18423);
or U18551 (N_18551,N_18496,N_18436);
xnor U18552 (N_18552,N_18338,N_18429);
or U18553 (N_18553,N_18459,N_18300);
and U18554 (N_18554,N_18404,N_18381);
or U18555 (N_18555,N_18452,N_18295);
nor U18556 (N_18556,N_18293,N_18432);
nor U18557 (N_18557,N_18372,N_18383);
nand U18558 (N_18558,N_18499,N_18279);
and U18559 (N_18559,N_18467,N_18472);
nand U18560 (N_18560,N_18369,N_18445);
and U18561 (N_18561,N_18317,N_18390);
xnor U18562 (N_18562,N_18331,N_18377);
nand U18563 (N_18563,N_18382,N_18267);
xnor U18564 (N_18564,N_18454,N_18475);
nor U18565 (N_18565,N_18498,N_18379);
xor U18566 (N_18566,N_18334,N_18460);
or U18567 (N_18567,N_18487,N_18477);
and U18568 (N_18568,N_18363,N_18274);
nor U18569 (N_18569,N_18484,N_18466);
nand U18570 (N_18570,N_18327,N_18343);
and U18571 (N_18571,N_18262,N_18421);
xnor U18572 (N_18572,N_18447,N_18440);
nand U18573 (N_18573,N_18396,N_18263);
nand U18574 (N_18574,N_18455,N_18328);
and U18575 (N_18575,N_18367,N_18265);
nand U18576 (N_18576,N_18254,N_18442);
xnor U18577 (N_18577,N_18482,N_18449);
nand U18578 (N_18578,N_18378,N_18282);
nand U18579 (N_18579,N_18468,N_18488);
and U18580 (N_18580,N_18456,N_18457);
xnor U18581 (N_18581,N_18313,N_18336);
nand U18582 (N_18582,N_18348,N_18418);
nand U18583 (N_18583,N_18332,N_18358);
nand U18584 (N_18584,N_18485,N_18257);
or U18585 (N_18585,N_18361,N_18411);
nand U18586 (N_18586,N_18486,N_18476);
and U18587 (N_18587,N_18375,N_18290);
and U18588 (N_18588,N_18497,N_18306);
nor U18589 (N_18589,N_18384,N_18353);
and U18590 (N_18590,N_18368,N_18256);
xor U18591 (N_18591,N_18271,N_18422);
xnor U18592 (N_18592,N_18311,N_18398);
nor U18593 (N_18593,N_18341,N_18269);
nor U18594 (N_18594,N_18356,N_18301);
xor U18595 (N_18595,N_18403,N_18286);
or U18596 (N_18596,N_18365,N_18478);
nor U18597 (N_18597,N_18463,N_18394);
and U18598 (N_18598,N_18471,N_18441);
and U18599 (N_18599,N_18323,N_18389);
nor U18600 (N_18600,N_18416,N_18285);
nand U18601 (N_18601,N_18402,N_18473);
nor U18602 (N_18602,N_18292,N_18258);
nand U18603 (N_18603,N_18357,N_18283);
xor U18604 (N_18604,N_18392,N_18491);
and U18605 (N_18605,N_18303,N_18410);
nand U18606 (N_18606,N_18433,N_18275);
nand U18607 (N_18607,N_18493,N_18315);
nor U18608 (N_18608,N_18268,N_18307);
and U18609 (N_18609,N_18437,N_18305);
nand U18610 (N_18610,N_18395,N_18451);
and U18611 (N_18611,N_18298,N_18277);
or U18612 (N_18612,N_18414,N_18388);
or U18613 (N_18613,N_18489,N_18435);
nand U18614 (N_18614,N_18255,N_18439);
nor U18615 (N_18615,N_18419,N_18346);
xnor U18616 (N_18616,N_18420,N_18273);
nand U18617 (N_18617,N_18280,N_18448);
nor U18618 (N_18618,N_18349,N_18329);
nor U18619 (N_18619,N_18450,N_18272);
or U18620 (N_18620,N_18438,N_18408);
or U18621 (N_18621,N_18374,N_18316);
nand U18622 (N_18622,N_18351,N_18337);
nand U18623 (N_18623,N_18366,N_18342);
and U18624 (N_18624,N_18401,N_18359);
xor U18625 (N_18625,N_18466,N_18462);
and U18626 (N_18626,N_18450,N_18455);
nor U18627 (N_18627,N_18497,N_18297);
and U18628 (N_18628,N_18262,N_18291);
xor U18629 (N_18629,N_18396,N_18424);
or U18630 (N_18630,N_18381,N_18326);
xnor U18631 (N_18631,N_18282,N_18356);
xor U18632 (N_18632,N_18292,N_18423);
nand U18633 (N_18633,N_18404,N_18475);
nand U18634 (N_18634,N_18355,N_18383);
xnor U18635 (N_18635,N_18418,N_18497);
nand U18636 (N_18636,N_18315,N_18437);
and U18637 (N_18637,N_18363,N_18282);
nand U18638 (N_18638,N_18421,N_18454);
or U18639 (N_18639,N_18341,N_18438);
or U18640 (N_18640,N_18411,N_18496);
or U18641 (N_18641,N_18453,N_18355);
xnor U18642 (N_18642,N_18424,N_18371);
and U18643 (N_18643,N_18328,N_18437);
or U18644 (N_18644,N_18269,N_18344);
xor U18645 (N_18645,N_18275,N_18456);
nand U18646 (N_18646,N_18273,N_18433);
or U18647 (N_18647,N_18424,N_18314);
nand U18648 (N_18648,N_18460,N_18412);
xnor U18649 (N_18649,N_18297,N_18366);
and U18650 (N_18650,N_18393,N_18307);
and U18651 (N_18651,N_18303,N_18480);
and U18652 (N_18652,N_18389,N_18386);
or U18653 (N_18653,N_18493,N_18339);
nand U18654 (N_18654,N_18498,N_18355);
nor U18655 (N_18655,N_18340,N_18395);
xnor U18656 (N_18656,N_18372,N_18254);
nor U18657 (N_18657,N_18483,N_18296);
nor U18658 (N_18658,N_18284,N_18295);
nor U18659 (N_18659,N_18351,N_18491);
nor U18660 (N_18660,N_18430,N_18355);
and U18661 (N_18661,N_18474,N_18450);
nand U18662 (N_18662,N_18483,N_18342);
nand U18663 (N_18663,N_18263,N_18375);
xnor U18664 (N_18664,N_18331,N_18262);
nor U18665 (N_18665,N_18448,N_18453);
and U18666 (N_18666,N_18389,N_18480);
xnor U18667 (N_18667,N_18338,N_18362);
or U18668 (N_18668,N_18474,N_18377);
nor U18669 (N_18669,N_18420,N_18386);
nor U18670 (N_18670,N_18417,N_18411);
nand U18671 (N_18671,N_18312,N_18263);
xnor U18672 (N_18672,N_18466,N_18281);
and U18673 (N_18673,N_18352,N_18343);
nor U18674 (N_18674,N_18453,N_18471);
nor U18675 (N_18675,N_18340,N_18291);
nor U18676 (N_18676,N_18448,N_18333);
nor U18677 (N_18677,N_18270,N_18478);
or U18678 (N_18678,N_18273,N_18459);
nand U18679 (N_18679,N_18316,N_18367);
nand U18680 (N_18680,N_18438,N_18425);
and U18681 (N_18681,N_18444,N_18285);
xor U18682 (N_18682,N_18315,N_18282);
or U18683 (N_18683,N_18289,N_18439);
nor U18684 (N_18684,N_18372,N_18387);
nor U18685 (N_18685,N_18410,N_18292);
xnor U18686 (N_18686,N_18300,N_18369);
xnor U18687 (N_18687,N_18301,N_18268);
nor U18688 (N_18688,N_18300,N_18489);
or U18689 (N_18689,N_18261,N_18473);
or U18690 (N_18690,N_18325,N_18289);
nor U18691 (N_18691,N_18446,N_18399);
nor U18692 (N_18692,N_18266,N_18302);
xnor U18693 (N_18693,N_18453,N_18449);
xor U18694 (N_18694,N_18260,N_18410);
nand U18695 (N_18695,N_18330,N_18405);
or U18696 (N_18696,N_18306,N_18333);
xnor U18697 (N_18697,N_18269,N_18297);
xnor U18698 (N_18698,N_18429,N_18463);
and U18699 (N_18699,N_18269,N_18412);
or U18700 (N_18700,N_18445,N_18443);
and U18701 (N_18701,N_18406,N_18464);
or U18702 (N_18702,N_18432,N_18291);
or U18703 (N_18703,N_18360,N_18401);
or U18704 (N_18704,N_18498,N_18490);
xnor U18705 (N_18705,N_18401,N_18423);
nor U18706 (N_18706,N_18271,N_18349);
xor U18707 (N_18707,N_18499,N_18375);
nor U18708 (N_18708,N_18272,N_18388);
nor U18709 (N_18709,N_18345,N_18271);
or U18710 (N_18710,N_18338,N_18300);
nand U18711 (N_18711,N_18380,N_18346);
nand U18712 (N_18712,N_18448,N_18490);
nor U18713 (N_18713,N_18451,N_18369);
xnor U18714 (N_18714,N_18488,N_18295);
and U18715 (N_18715,N_18319,N_18263);
or U18716 (N_18716,N_18488,N_18277);
nand U18717 (N_18717,N_18464,N_18355);
and U18718 (N_18718,N_18367,N_18418);
or U18719 (N_18719,N_18307,N_18329);
or U18720 (N_18720,N_18464,N_18280);
nand U18721 (N_18721,N_18334,N_18385);
xor U18722 (N_18722,N_18269,N_18480);
nor U18723 (N_18723,N_18381,N_18353);
nand U18724 (N_18724,N_18472,N_18355);
nand U18725 (N_18725,N_18336,N_18398);
nand U18726 (N_18726,N_18277,N_18395);
nor U18727 (N_18727,N_18494,N_18436);
xor U18728 (N_18728,N_18292,N_18427);
and U18729 (N_18729,N_18474,N_18449);
xnor U18730 (N_18730,N_18306,N_18374);
nor U18731 (N_18731,N_18253,N_18436);
nor U18732 (N_18732,N_18362,N_18345);
or U18733 (N_18733,N_18326,N_18372);
nand U18734 (N_18734,N_18307,N_18306);
or U18735 (N_18735,N_18443,N_18337);
xnor U18736 (N_18736,N_18331,N_18318);
nor U18737 (N_18737,N_18300,N_18381);
and U18738 (N_18738,N_18392,N_18454);
xor U18739 (N_18739,N_18469,N_18365);
xor U18740 (N_18740,N_18401,N_18277);
and U18741 (N_18741,N_18426,N_18445);
nor U18742 (N_18742,N_18446,N_18331);
xnor U18743 (N_18743,N_18369,N_18388);
or U18744 (N_18744,N_18412,N_18325);
nand U18745 (N_18745,N_18259,N_18360);
or U18746 (N_18746,N_18407,N_18258);
and U18747 (N_18747,N_18485,N_18251);
xnor U18748 (N_18748,N_18435,N_18407);
nor U18749 (N_18749,N_18364,N_18311);
nand U18750 (N_18750,N_18544,N_18714);
or U18751 (N_18751,N_18562,N_18652);
or U18752 (N_18752,N_18502,N_18598);
and U18753 (N_18753,N_18619,N_18533);
nor U18754 (N_18754,N_18550,N_18737);
and U18755 (N_18755,N_18724,N_18697);
xnor U18756 (N_18756,N_18545,N_18593);
nor U18757 (N_18757,N_18564,N_18575);
nor U18758 (N_18758,N_18704,N_18520);
nor U18759 (N_18759,N_18688,N_18509);
and U18760 (N_18760,N_18569,N_18504);
nand U18761 (N_18761,N_18603,N_18648);
and U18762 (N_18762,N_18551,N_18730);
nand U18763 (N_18763,N_18525,N_18604);
and U18764 (N_18764,N_18613,N_18515);
nor U18765 (N_18765,N_18541,N_18620);
nand U18766 (N_18766,N_18543,N_18679);
and U18767 (N_18767,N_18549,N_18727);
nor U18768 (N_18768,N_18723,N_18703);
xnor U18769 (N_18769,N_18728,N_18553);
xnor U18770 (N_18770,N_18673,N_18686);
and U18771 (N_18771,N_18529,N_18660);
and U18772 (N_18772,N_18634,N_18701);
and U18773 (N_18773,N_18552,N_18505);
or U18774 (N_18774,N_18537,N_18744);
or U18775 (N_18775,N_18700,N_18725);
or U18776 (N_18776,N_18616,N_18694);
nand U18777 (N_18777,N_18611,N_18710);
or U18778 (N_18778,N_18623,N_18641);
nor U18779 (N_18779,N_18582,N_18542);
xor U18780 (N_18780,N_18540,N_18632);
or U18781 (N_18781,N_18693,N_18628);
nor U18782 (N_18782,N_18610,N_18731);
xnor U18783 (N_18783,N_18548,N_18666);
and U18784 (N_18784,N_18718,N_18567);
xor U18785 (N_18785,N_18584,N_18655);
or U18786 (N_18786,N_18659,N_18500);
xnor U18787 (N_18787,N_18699,N_18661);
nor U18788 (N_18788,N_18594,N_18713);
xnor U18789 (N_18789,N_18558,N_18635);
nand U18790 (N_18790,N_18748,N_18735);
or U18791 (N_18791,N_18706,N_18637);
xor U18792 (N_18792,N_18747,N_18521);
nand U18793 (N_18793,N_18615,N_18506);
xor U18794 (N_18794,N_18579,N_18514);
or U18795 (N_18795,N_18707,N_18586);
and U18796 (N_18796,N_18588,N_18678);
and U18797 (N_18797,N_18547,N_18539);
nor U18798 (N_18798,N_18617,N_18527);
nor U18799 (N_18799,N_18646,N_18683);
and U18800 (N_18800,N_18740,N_18702);
and U18801 (N_18801,N_18669,N_18689);
nand U18802 (N_18802,N_18599,N_18519);
nor U18803 (N_18803,N_18696,N_18522);
xnor U18804 (N_18804,N_18501,N_18528);
and U18805 (N_18805,N_18530,N_18614);
and U18806 (N_18806,N_18535,N_18680);
and U18807 (N_18807,N_18577,N_18578);
nor U18808 (N_18808,N_18722,N_18517);
and U18809 (N_18809,N_18605,N_18555);
nor U18810 (N_18810,N_18560,N_18631);
xor U18811 (N_18811,N_18587,N_18656);
or U18812 (N_18812,N_18576,N_18622);
and U18813 (N_18813,N_18624,N_18667);
and U18814 (N_18814,N_18717,N_18636);
xor U18815 (N_18815,N_18523,N_18513);
nor U18816 (N_18816,N_18671,N_18556);
or U18817 (N_18817,N_18531,N_18732);
nand U18818 (N_18818,N_18565,N_18695);
xnor U18819 (N_18819,N_18658,N_18526);
xnor U18820 (N_18820,N_18573,N_18626);
or U18821 (N_18821,N_18709,N_18566);
xor U18822 (N_18822,N_18650,N_18609);
xor U18823 (N_18823,N_18601,N_18612);
and U18824 (N_18824,N_18649,N_18534);
nor U18825 (N_18825,N_18677,N_18682);
xnor U18826 (N_18826,N_18745,N_18524);
xor U18827 (N_18827,N_18716,N_18705);
or U18828 (N_18828,N_18643,N_18625);
and U18829 (N_18829,N_18657,N_18674);
nand U18830 (N_18830,N_18585,N_18712);
xor U18831 (N_18831,N_18607,N_18568);
and U18832 (N_18832,N_18670,N_18561);
nor U18833 (N_18833,N_18639,N_18721);
and U18834 (N_18834,N_18608,N_18738);
nand U18835 (N_18835,N_18672,N_18690);
and U18836 (N_18836,N_18736,N_18726);
nor U18837 (N_18837,N_18651,N_18600);
and U18838 (N_18838,N_18741,N_18572);
nor U18839 (N_18839,N_18581,N_18580);
xor U18840 (N_18840,N_18681,N_18729);
nand U18841 (N_18841,N_18536,N_18597);
or U18842 (N_18842,N_18692,N_18583);
nand U18843 (N_18843,N_18592,N_18645);
nor U18844 (N_18844,N_18675,N_18621);
xor U18845 (N_18845,N_18512,N_18596);
nor U18846 (N_18846,N_18629,N_18691);
nor U18847 (N_18847,N_18685,N_18734);
and U18848 (N_18848,N_18590,N_18739);
xor U18849 (N_18849,N_18640,N_18654);
nand U18850 (N_18850,N_18507,N_18638);
nor U18851 (N_18851,N_18510,N_18570);
and U18852 (N_18852,N_18733,N_18664);
nor U18853 (N_18853,N_18743,N_18627);
xor U18854 (N_18854,N_18546,N_18589);
and U18855 (N_18855,N_18653,N_18538);
nand U18856 (N_18856,N_18559,N_18662);
nor U18857 (N_18857,N_18602,N_18715);
nand U18858 (N_18858,N_18571,N_18595);
nor U18859 (N_18859,N_18633,N_18708);
nand U18860 (N_18860,N_18618,N_18711);
or U18861 (N_18861,N_18511,N_18720);
or U18862 (N_18862,N_18532,N_18630);
or U18863 (N_18863,N_18518,N_18749);
nand U18864 (N_18864,N_18719,N_18687);
or U18865 (N_18865,N_18554,N_18644);
nand U18866 (N_18866,N_18684,N_18668);
nor U18867 (N_18867,N_18698,N_18606);
or U18868 (N_18868,N_18591,N_18742);
nor U18869 (N_18869,N_18516,N_18676);
nor U18870 (N_18870,N_18503,N_18746);
or U18871 (N_18871,N_18508,N_18665);
nor U18872 (N_18872,N_18557,N_18647);
xor U18873 (N_18873,N_18574,N_18563);
and U18874 (N_18874,N_18642,N_18663);
xor U18875 (N_18875,N_18682,N_18712);
nor U18876 (N_18876,N_18670,N_18611);
xnor U18877 (N_18877,N_18614,N_18599);
xnor U18878 (N_18878,N_18614,N_18534);
nand U18879 (N_18879,N_18639,N_18678);
xnor U18880 (N_18880,N_18509,N_18500);
and U18881 (N_18881,N_18581,N_18716);
and U18882 (N_18882,N_18519,N_18640);
nand U18883 (N_18883,N_18560,N_18659);
xnor U18884 (N_18884,N_18560,N_18535);
nand U18885 (N_18885,N_18566,N_18588);
or U18886 (N_18886,N_18600,N_18625);
xnor U18887 (N_18887,N_18641,N_18537);
or U18888 (N_18888,N_18632,N_18522);
or U18889 (N_18889,N_18745,N_18556);
xor U18890 (N_18890,N_18505,N_18515);
or U18891 (N_18891,N_18735,N_18642);
or U18892 (N_18892,N_18648,N_18601);
nor U18893 (N_18893,N_18684,N_18526);
xnor U18894 (N_18894,N_18565,N_18642);
nand U18895 (N_18895,N_18570,N_18607);
xor U18896 (N_18896,N_18667,N_18715);
and U18897 (N_18897,N_18643,N_18537);
xnor U18898 (N_18898,N_18521,N_18624);
nor U18899 (N_18899,N_18597,N_18558);
xor U18900 (N_18900,N_18672,N_18524);
nand U18901 (N_18901,N_18540,N_18610);
or U18902 (N_18902,N_18671,N_18598);
and U18903 (N_18903,N_18605,N_18748);
nor U18904 (N_18904,N_18608,N_18609);
and U18905 (N_18905,N_18715,N_18671);
xnor U18906 (N_18906,N_18505,N_18614);
nor U18907 (N_18907,N_18699,N_18566);
nor U18908 (N_18908,N_18708,N_18725);
and U18909 (N_18909,N_18539,N_18638);
nor U18910 (N_18910,N_18695,N_18624);
nor U18911 (N_18911,N_18589,N_18533);
and U18912 (N_18912,N_18639,N_18690);
and U18913 (N_18913,N_18508,N_18731);
nand U18914 (N_18914,N_18648,N_18593);
or U18915 (N_18915,N_18633,N_18660);
nor U18916 (N_18916,N_18531,N_18724);
xnor U18917 (N_18917,N_18643,N_18554);
nand U18918 (N_18918,N_18556,N_18560);
nor U18919 (N_18919,N_18559,N_18712);
nor U18920 (N_18920,N_18511,N_18654);
nor U18921 (N_18921,N_18592,N_18517);
nand U18922 (N_18922,N_18616,N_18535);
or U18923 (N_18923,N_18585,N_18633);
nand U18924 (N_18924,N_18629,N_18634);
and U18925 (N_18925,N_18544,N_18549);
xnor U18926 (N_18926,N_18629,N_18523);
nor U18927 (N_18927,N_18524,N_18713);
and U18928 (N_18928,N_18602,N_18576);
nor U18929 (N_18929,N_18665,N_18705);
and U18930 (N_18930,N_18510,N_18560);
nor U18931 (N_18931,N_18592,N_18694);
nor U18932 (N_18932,N_18714,N_18553);
or U18933 (N_18933,N_18566,N_18662);
nand U18934 (N_18934,N_18521,N_18678);
nor U18935 (N_18935,N_18651,N_18700);
or U18936 (N_18936,N_18682,N_18633);
nand U18937 (N_18937,N_18612,N_18662);
nor U18938 (N_18938,N_18670,N_18591);
nor U18939 (N_18939,N_18739,N_18605);
nor U18940 (N_18940,N_18566,N_18739);
or U18941 (N_18941,N_18718,N_18527);
and U18942 (N_18942,N_18719,N_18572);
xor U18943 (N_18943,N_18566,N_18519);
nor U18944 (N_18944,N_18664,N_18647);
and U18945 (N_18945,N_18548,N_18562);
and U18946 (N_18946,N_18551,N_18518);
or U18947 (N_18947,N_18637,N_18636);
nand U18948 (N_18948,N_18511,N_18740);
xor U18949 (N_18949,N_18697,N_18666);
and U18950 (N_18950,N_18520,N_18589);
or U18951 (N_18951,N_18535,N_18595);
and U18952 (N_18952,N_18599,N_18506);
nor U18953 (N_18953,N_18564,N_18685);
and U18954 (N_18954,N_18697,N_18650);
nand U18955 (N_18955,N_18590,N_18618);
nand U18956 (N_18956,N_18582,N_18681);
and U18957 (N_18957,N_18710,N_18549);
or U18958 (N_18958,N_18558,N_18515);
nor U18959 (N_18959,N_18600,N_18634);
and U18960 (N_18960,N_18575,N_18511);
nand U18961 (N_18961,N_18740,N_18629);
or U18962 (N_18962,N_18747,N_18665);
and U18963 (N_18963,N_18518,N_18507);
nand U18964 (N_18964,N_18719,N_18723);
nor U18965 (N_18965,N_18602,N_18742);
xnor U18966 (N_18966,N_18679,N_18674);
nand U18967 (N_18967,N_18533,N_18503);
nor U18968 (N_18968,N_18511,N_18716);
nor U18969 (N_18969,N_18671,N_18702);
xor U18970 (N_18970,N_18661,N_18659);
nor U18971 (N_18971,N_18537,N_18742);
xnor U18972 (N_18972,N_18516,N_18690);
nor U18973 (N_18973,N_18531,N_18680);
and U18974 (N_18974,N_18550,N_18747);
nor U18975 (N_18975,N_18555,N_18603);
and U18976 (N_18976,N_18521,N_18641);
nor U18977 (N_18977,N_18609,N_18519);
or U18978 (N_18978,N_18731,N_18739);
and U18979 (N_18979,N_18648,N_18519);
or U18980 (N_18980,N_18619,N_18583);
and U18981 (N_18981,N_18659,N_18539);
xnor U18982 (N_18982,N_18666,N_18546);
nor U18983 (N_18983,N_18636,N_18576);
and U18984 (N_18984,N_18729,N_18661);
or U18985 (N_18985,N_18545,N_18675);
xor U18986 (N_18986,N_18542,N_18550);
nand U18987 (N_18987,N_18562,N_18535);
nor U18988 (N_18988,N_18721,N_18599);
nand U18989 (N_18989,N_18511,N_18725);
xnor U18990 (N_18990,N_18592,N_18640);
nor U18991 (N_18991,N_18564,N_18586);
and U18992 (N_18992,N_18616,N_18536);
or U18993 (N_18993,N_18693,N_18558);
and U18994 (N_18994,N_18665,N_18741);
or U18995 (N_18995,N_18514,N_18610);
nor U18996 (N_18996,N_18676,N_18683);
nand U18997 (N_18997,N_18693,N_18747);
nand U18998 (N_18998,N_18720,N_18742);
and U18999 (N_18999,N_18692,N_18669);
and U19000 (N_19000,N_18977,N_18907);
nand U19001 (N_19001,N_18825,N_18864);
nand U19002 (N_19002,N_18779,N_18955);
or U19003 (N_19003,N_18998,N_18934);
nor U19004 (N_19004,N_18992,N_18892);
xnor U19005 (N_19005,N_18914,N_18827);
xnor U19006 (N_19006,N_18958,N_18860);
nand U19007 (N_19007,N_18789,N_18803);
nand U19008 (N_19008,N_18840,N_18869);
xor U19009 (N_19009,N_18900,N_18973);
or U19010 (N_19010,N_18935,N_18929);
or U19011 (N_19011,N_18817,N_18888);
or U19012 (N_19012,N_18926,N_18780);
xor U19013 (N_19013,N_18906,N_18889);
and U19014 (N_19014,N_18752,N_18867);
nor U19015 (N_19015,N_18815,N_18863);
xor U19016 (N_19016,N_18836,N_18925);
nand U19017 (N_19017,N_18823,N_18950);
or U19018 (N_19018,N_18875,N_18849);
and U19019 (N_19019,N_18795,N_18757);
xnor U19020 (N_19020,N_18865,N_18902);
or U19021 (N_19021,N_18982,N_18932);
nor U19022 (N_19022,N_18931,N_18763);
nor U19023 (N_19023,N_18927,N_18801);
and U19024 (N_19024,N_18845,N_18847);
and U19025 (N_19025,N_18981,N_18966);
nand U19026 (N_19026,N_18756,N_18873);
nor U19027 (N_19027,N_18921,N_18793);
nor U19028 (N_19028,N_18799,N_18974);
nor U19029 (N_19029,N_18897,N_18874);
nand U19030 (N_19030,N_18798,N_18913);
or U19031 (N_19031,N_18947,N_18945);
and U19032 (N_19032,N_18922,N_18937);
xnor U19033 (N_19033,N_18933,N_18987);
nor U19034 (N_19034,N_18970,N_18991);
nor U19035 (N_19035,N_18884,N_18818);
nand U19036 (N_19036,N_18995,N_18936);
and U19037 (N_19037,N_18866,N_18954);
and U19038 (N_19038,N_18814,N_18963);
or U19039 (N_19039,N_18809,N_18972);
or U19040 (N_19040,N_18766,N_18854);
or U19041 (N_19041,N_18846,N_18880);
nor U19042 (N_19042,N_18841,N_18968);
xor U19043 (N_19043,N_18885,N_18843);
or U19044 (N_19044,N_18871,N_18834);
xor U19045 (N_19045,N_18750,N_18917);
nor U19046 (N_19046,N_18794,N_18760);
or U19047 (N_19047,N_18772,N_18877);
nand U19048 (N_19048,N_18790,N_18753);
or U19049 (N_19049,N_18961,N_18764);
and U19050 (N_19050,N_18946,N_18942);
nor U19051 (N_19051,N_18797,N_18923);
nor U19052 (N_19052,N_18759,N_18876);
nand U19053 (N_19053,N_18890,N_18870);
and U19054 (N_19054,N_18915,N_18879);
nor U19055 (N_19055,N_18829,N_18769);
or U19056 (N_19056,N_18957,N_18909);
or U19057 (N_19057,N_18788,N_18819);
or U19058 (N_19058,N_18959,N_18978);
nand U19059 (N_19059,N_18859,N_18979);
or U19060 (N_19060,N_18895,N_18887);
nand U19061 (N_19061,N_18761,N_18988);
or U19062 (N_19062,N_18878,N_18810);
and U19063 (N_19063,N_18778,N_18953);
nand U19064 (N_19064,N_18853,N_18912);
nand U19065 (N_19065,N_18898,N_18872);
and U19066 (N_19066,N_18904,N_18808);
and U19067 (N_19067,N_18883,N_18768);
nand U19068 (N_19068,N_18903,N_18850);
and U19069 (N_19069,N_18944,N_18813);
and U19070 (N_19070,N_18777,N_18997);
and U19071 (N_19071,N_18905,N_18886);
xor U19072 (N_19072,N_18824,N_18857);
nand U19073 (N_19073,N_18800,N_18767);
xnor U19074 (N_19074,N_18938,N_18868);
and U19075 (N_19075,N_18983,N_18891);
or U19076 (N_19076,N_18821,N_18838);
nand U19077 (N_19077,N_18758,N_18893);
nor U19078 (N_19078,N_18916,N_18774);
or U19079 (N_19079,N_18831,N_18771);
and U19080 (N_19080,N_18993,N_18920);
nor U19081 (N_19081,N_18773,N_18861);
and U19082 (N_19082,N_18828,N_18969);
xor U19083 (N_19083,N_18984,N_18822);
nand U19084 (N_19084,N_18855,N_18930);
and U19085 (N_19085,N_18996,N_18911);
or U19086 (N_19086,N_18899,N_18783);
nand U19087 (N_19087,N_18852,N_18805);
nand U19088 (N_19088,N_18960,N_18802);
nand U19089 (N_19089,N_18806,N_18786);
nand U19090 (N_19090,N_18762,N_18994);
xor U19091 (N_19091,N_18775,N_18796);
or U19092 (N_19092,N_18751,N_18989);
and U19093 (N_19093,N_18755,N_18948);
or U19094 (N_19094,N_18943,N_18882);
or U19095 (N_19095,N_18791,N_18826);
nor U19096 (N_19096,N_18842,N_18962);
and U19097 (N_19097,N_18862,N_18881);
xor U19098 (N_19098,N_18928,N_18952);
and U19099 (N_19099,N_18782,N_18941);
or U19100 (N_19100,N_18910,N_18951);
nor U19101 (N_19101,N_18811,N_18901);
xnor U19102 (N_19102,N_18833,N_18765);
or U19103 (N_19103,N_18844,N_18939);
nand U19104 (N_19104,N_18999,N_18830);
xor U19105 (N_19105,N_18754,N_18851);
and U19106 (N_19106,N_18856,N_18785);
nand U19107 (N_19107,N_18792,N_18896);
or U19108 (N_19108,N_18807,N_18986);
or U19109 (N_19109,N_18980,N_18816);
xor U19110 (N_19110,N_18985,N_18781);
nor U19111 (N_19111,N_18848,N_18967);
nand U19112 (N_19112,N_18835,N_18812);
nor U19113 (N_19113,N_18858,N_18776);
or U19114 (N_19114,N_18949,N_18908);
or U19115 (N_19115,N_18976,N_18975);
xnor U19116 (N_19116,N_18940,N_18990);
xor U19117 (N_19117,N_18924,N_18918);
nor U19118 (N_19118,N_18837,N_18839);
or U19119 (N_19119,N_18787,N_18971);
or U19120 (N_19120,N_18820,N_18919);
nor U19121 (N_19121,N_18770,N_18956);
or U19122 (N_19122,N_18784,N_18894);
xnor U19123 (N_19123,N_18832,N_18964);
nor U19124 (N_19124,N_18965,N_18804);
nand U19125 (N_19125,N_18948,N_18788);
xnor U19126 (N_19126,N_18978,N_18786);
nor U19127 (N_19127,N_18893,N_18928);
and U19128 (N_19128,N_18819,N_18842);
or U19129 (N_19129,N_18766,N_18799);
xnor U19130 (N_19130,N_18901,N_18852);
nand U19131 (N_19131,N_18870,N_18926);
nand U19132 (N_19132,N_18973,N_18856);
nor U19133 (N_19133,N_18886,N_18988);
and U19134 (N_19134,N_18966,N_18990);
nor U19135 (N_19135,N_18795,N_18882);
xor U19136 (N_19136,N_18844,N_18853);
and U19137 (N_19137,N_18916,N_18877);
xor U19138 (N_19138,N_18855,N_18889);
nor U19139 (N_19139,N_18938,N_18843);
nand U19140 (N_19140,N_18757,N_18838);
nand U19141 (N_19141,N_18921,N_18846);
and U19142 (N_19142,N_18773,N_18877);
or U19143 (N_19143,N_18991,N_18921);
nor U19144 (N_19144,N_18901,N_18785);
nor U19145 (N_19145,N_18993,N_18996);
nand U19146 (N_19146,N_18942,N_18781);
xnor U19147 (N_19147,N_18883,N_18859);
and U19148 (N_19148,N_18967,N_18860);
and U19149 (N_19149,N_18824,N_18760);
nand U19150 (N_19150,N_18851,N_18816);
nand U19151 (N_19151,N_18987,N_18982);
or U19152 (N_19152,N_18893,N_18855);
nor U19153 (N_19153,N_18899,N_18933);
xnor U19154 (N_19154,N_18979,N_18792);
or U19155 (N_19155,N_18931,N_18877);
nand U19156 (N_19156,N_18818,N_18988);
nand U19157 (N_19157,N_18775,N_18883);
and U19158 (N_19158,N_18914,N_18829);
and U19159 (N_19159,N_18831,N_18839);
nand U19160 (N_19160,N_18968,N_18872);
and U19161 (N_19161,N_18756,N_18858);
xnor U19162 (N_19162,N_18801,N_18790);
and U19163 (N_19163,N_18860,N_18936);
and U19164 (N_19164,N_18825,N_18977);
xor U19165 (N_19165,N_18844,N_18896);
xor U19166 (N_19166,N_18794,N_18844);
xor U19167 (N_19167,N_18835,N_18998);
and U19168 (N_19168,N_18824,N_18872);
or U19169 (N_19169,N_18775,N_18843);
nand U19170 (N_19170,N_18846,N_18820);
and U19171 (N_19171,N_18853,N_18934);
nand U19172 (N_19172,N_18848,N_18762);
or U19173 (N_19173,N_18793,N_18861);
and U19174 (N_19174,N_18887,N_18785);
nand U19175 (N_19175,N_18989,N_18902);
or U19176 (N_19176,N_18826,N_18792);
and U19177 (N_19177,N_18985,N_18894);
nand U19178 (N_19178,N_18831,N_18846);
nand U19179 (N_19179,N_18802,N_18766);
nor U19180 (N_19180,N_18820,N_18824);
nor U19181 (N_19181,N_18760,N_18763);
nand U19182 (N_19182,N_18861,N_18909);
or U19183 (N_19183,N_18785,N_18905);
nand U19184 (N_19184,N_18939,N_18954);
nor U19185 (N_19185,N_18827,N_18979);
nor U19186 (N_19186,N_18941,N_18806);
or U19187 (N_19187,N_18968,N_18812);
and U19188 (N_19188,N_18850,N_18832);
nand U19189 (N_19189,N_18881,N_18905);
and U19190 (N_19190,N_18964,N_18954);
xor U19191 (N_19191,N_18794,N_18818);
xnor U19192 (N_19192,N_18945,N_18872);
xnor U19193 (N_19193,N_18869,N_18884);
nand U19194 (N_19194,N_18822,N_18963);
and U19195 (N_19195,N_18837,N_18895);
nor U19196 (N_19196,N_18842,N_18990);
nand U19197 (N_19197,N_18876,N_18784);
nand U19198 (N_19198,N_18989,N_18856);
xor U19199 (N_19199,N_18945,N_18975);
nand U19200 (N_19200,N_18873,N_18971);
and U19201 (N_19201,N_18755,N_18995);
nor U19202 (N_19202,N_18835,N_18997);
and U19203 (N_19203,N_18851,N_18934);
nand U19204 (N_19204,N_18971,N_18786);
nor U19205 (N_19205,N_18898,N_18976);
nand U19206 (N_19206,N_18804,N_18936);
nand U19207 (N_19207,N_18750,N_18915);
xor U19208 (N_19208,N_18830,N_18821);
nor U19209 (N_19209,N_18787,N_18814);
nor U19210 (N_19210,N_18802,N_18780);
nand U19211 (N_19211,N_18946,N_18815);
nor U19212 (N_19212,N_18766,N_18805);
xor U19213 (N_19213,N_18981,N_18833);
nor U19214 (N_19214,N_18989,N_18984);
nand U19215 (N_19215,N_18820,N_18775);
xor U19216 (N_19216,N_18826,N_18880);
xnor U19217 (N_19217,N_18912,N_18955);
nor U19218 (N_19218,N_18876,N_18810);
or U19219 (N_19219,N_18905,N_18774);
nor U19220 (N_19220,N_18980,N_18896);
nor U19221 (N_19221,N_18772,N_18820);
nand U19222 (N_19222,N_18836,N_18762);
nand U19223 (N_19223,N_18801,N_18985);
and U19224 (N_19224,N_18779,N_18867);
or U19225 (N_19225,N_18886,N_18794);
xnor U19226 (N_19226,N_18773,N_18879);
nor U19227 (N_19227,N_18803,N_18839);
and U19228 (N_19228,N_18911,N_18858);
nand U19229 (N_19229,N_18756,N_18855);
xor U19230 (N_19230,N_18871,N_18756);
nand U19231 (N_19231,N_18911,N_18762);
nand U19232 (N_19232,N_18995,N_18820);
nand U19233 (N_19233,N_18848,N_18962);
or U19234 (N_19234,N_18778,N_18995);
nand U19235 (N_19235,N_18804,N_18909);
xor U19236 (N_19236,N_18883,N_18987);
and U19237 (N_19237,N_18815,N_18958);
nor U19238 (N_19238,N_18903,N_18907);
xnor U19239 (N_19239,N_18822,N_18912);
xnor U19240 (N_19240,N_18914,N_18758);
nand U19241 (N_19241,N_18871,N_18803);
and U19242 (N_19242,N_18970,N_18786);
and U19243 (N_19243,N_18955,N_18907);
or U19244 (N_19244,N_18781,N_18916);
nor U19245 (N_19245,N_18830,N_18879);
xnor U19246 (N_19246,N_18996,N_18976);
nor U19247 (N_19247,N_18876,N_18990);
and U19248 (N_19248,N_18993,N_18895);
nand U19249 (N_19249,N_18806,N_18855);
nor U19250 (N_19250,N_19171,N_19155);
xor U19251 (N_19251,N_19103,N_19043);
or U19252 (N_19252,N_19143,N_19176);
and U19253 (N_19253,N_19080,N_19170);
nor U19254 (N_19254,N_19180,N_19196);
nor U19255 (N_19255,N_19087,N_19088);
nand U19256 (N_19256,N_19082,N_19092);
xor U19257 (N_19257,N_19131,N_19248);
or U19258 (N_19258,N_19157,N_19240);
nor U19259 (N_19259,N_19095,N_19216);
nand U19260 (N_19260,N_19219,N_19089);
nor U19261 (N_19261,N_19137,N_19182);
xor U19262 (N_19262,N_19034,N_19029);
nor U19263 (N_19263,N_19208,N_19084);
nor U19264 (N_19264,N_19153,N_19159);
and U19265 (N_19265,N_19236,N_19207);
xor U19266 (N_19266,N_19183,N_19017);
nor U19267 (N_19267,N_19169,N_19122);
xor U19268 (N_19268,N_19147,N_19053);
nand U19269 (N_19269,N_19086,N_19192);
xor U19270 (N_19270,N_19133,N_19058);
xnor U19271 (N_19271,N_19060,N_19209);
nor U19272 (N_19272,N_19128,N_19054);
and U19273 (N_19273,N_19041,N_19066);
or U19274 (N_19274,N_19116,N_19142);
nand U19275 (N_19275,N_19063,N_19015);
nand U19276 (N_19276,N_19098,N_19028);
nor U19277 (N_19277,N_19065,N_19056);
nor U19278 (N_19278,N_19109,N_19174);
xnor U19279 (N_19279,N_19213,N_19106);
or U19280 (N_19280,N_19019,N_19190);
xor U19281 (N_19281,N_19023,N_19117);
or U19282 (N_19282,N_19102,N_19038);
xor U19283 (N_19283,N_19186,N_19107);
or U19284 (N_19284,N_19242,N_19024);
nand U19285 (N_19285,N_19198,N_19051);
and U19286 (N_19286,N_19026,N_19111);
xnor U19287 (N_19287,N_19225,N_19090);
nand U19288 (N_19288,N_19123,N_19185);
or U19289 (N_19289,N_19203,N_19067);
xor U19290 (N_19290,N_19246,N_19140);
xor U19291 (N_19291,N_19114,N_19126);
nand U19292 (N_19292,N_19184,N_19244);
nand U19293 (N_19293,N_19221,N_19188);
or U19294 (N_19294,N_19223,N_19230);
nand U19295 (N_19295,N_19162,N_19181);
xor U19296 (N_19296,N_19218,N_19108);
and U19297 (N_19297,N_19073,N_19050);
xor U19298 (N_19298,N_19004,N_19007);
xor U19299 (N_19299,N_19070,N_19206);
and U19300 (N_19300,N_19138,N_19195);
nor U19301 (N_19301,N_19167,N_19201);
xor U19302 (N_19302,N_19168,N_19212);
nor U19303 (N_19303,N_19074,N_19215);
or U19304 (N_19304,N_19172,N_19036);
xor U19305 (N_19305,N_19227,N_19130);
xnor U19306 (N_19306,N_19046,N_19217);
nor U19307 (N_19307,N_19151,N_19222);
nor U19308 (N_19308,N_19234,N_19048);
nand U19309 (N_19309,N_19042,N_19228);
nor U19310 (N_19310,N_19068,N_19178);
nand U19311 (N_19311,N_19165,N_19112);
nor U19312 (N_19312,N_19239,N_19166);
or U19313 (N_19313,N_19160,N_19132);
or U19314 (N_19314,N_19064,N_19161);
and U19315 (N_19315,N_19049,N_19158);
nand U19316 (N_19316,N_19135,N_19055);
or U19317 (N_19317,N_19245,N_19009);
and U19318 (N_19318,N_19241,N_19083);
or U19319 (N_19319,N_19104,N_19220);
or U19320 (N_19320,N_19016,N_19033);
nor U19321 (N_19321,N_19232,N_19096);
or U19322 (N_19322,N_19145,N_19205);
nand U19323 (N_19323,N_19008,N_19075);
or U19324 (N_19324,N_19211,N_19076);
and U19325 (N_19325,N_19022,N_19121);
xnor U19326 (N_19326,N_19148,N_19020);
nand U19327 (N_19327,N_19071,N_19224);
or U19328 (N_19328,N_19079,N_19124);
and U19329 (N_19329,N_19175,N_19040);
nor U19330 (N_19330,N_19005,N_19139);
nand U19331 (N_19331,N_19057,N_19177);
or U19332 (N_19332,N_19163,N_19091);
nor U19333 (N_19333,N_19129,N_19035);
and U19334 (N_19334,N_19031,N_19204);
nand U19335 (N_19335,N_19100,N_19173);
nor U19336 (N_19336,N_19105,N_19110);
and U19337 (N_19337,N_19141,N_19039);
xor U19338 (N_19338,N_19136,N_19237);
or U19339 (N_19339,N_19062,N_19010);
xor U19340 (N_19340,N_19189,N_19018);
or U19341 (N_19341,N_19006,N_19179);
nand U19342 (N_19342,N_19013,N_19037);
or U19343 (N_19343,N_19059,N_19187);
or U19344 (N_19344,N_19078,N_19032);
nor U19345 (N_19345,N_19202,N_19115);
xor U19346 (N_19346,N_19238,N_19120);
and U19347 (N_19347,N_19027,N_19003);
xnor U19348 (N_19348,N_19030,N_19149);
xor U19349 (N_19349,N_19156,N_19072);
nand U19350 (N_19350,N_19200,N_19146);
nor U19351 (N_19351,N_19247,N_19194);
and U19352 (N_19352,N_19052,N_19197);
and U19353 (N_19353,N_19214,N_19085);
or U19354 (N_19354,N_19012,N_19069);
nor U19355 (N_19355,N_19011,N_19014);
xor U19356 (N_19356,N_19233,N_19081);
or U19357 (N_19357,N_19118,N_19249);
and U19358 (N_19358,N_19193,N_19001);
or U19359 (N_19359,N_19101,N_19047);
or U19360 (N_19360,N_19119,N_19113);
or U19361 (N_19361,N_19164,N_19127);
xor U19362 (N_19362,N_19093,N_19154);
or U19363 (N_19363,N_19000,N_19097);
nand U19364 (N_19364,N_19191,N_19125);
xor U19365 (N_19365,N_19044,N_19021);
nor U19366 (N_19366,N_19025,N_19134);
xor U19367 (N_19367,N_19045,N_19229);
and U19368 (N_19368,N_19150,N_19152);
or U19369 (N_19369,N_19099,N_19235);
nor U19370 (N_19370,N_19226,N_19002);
nand U19371 (N_19371,N_19210,N_19094);
nand U19372 (N_19372,N_19231,N_19199);
and U19373 (N_19373,N_19144,N_19061);
and U19374 (N_19374,N_19077,N_19243);
or U19375 (N_19375,N_19218,N_19085);
xnor U19376 (N_19376,N_19106,N_19132);
or U19377 (N_19377,N_19148,N_19190);
xnor U19378 (N_19378,N_19124,N_19249);
or U19379 (N_19379,N_19233,N_19214);
nor U19380 (N_19380,N_19213,N_19224);
xnor U19381 (N_19381,N_19221,N_19129);
nor U19382 (N_19382,N_19018,N_19194);
or U19383 (N_19383,N_19211,N_19207);
nor U19384 (N_19384,N_19197,N_19204);
xor U19385 (N_19385,N_19155,N_19209);
xor U19386 (N_19386,N_19123,N_19189);
or U19387 (N_19387,N_19115,N_19193);
or U19388 (N_19388,N_19245,N_19128);
nand U19389 (N_19389,N_19119,N_19108);
nor U19390 (N_19390,N_19107,N_19120);
nor U19391 (N_19391,N_19057,N_19101);
and U19392 (N_19392,N_19095,N_19091);
xnor U19393 (N_19393,N_19165,N_19240);
and U19394 (N_19394,N_19185,N_19121);
nor U19395 (N_19395,N_19165,N_19191);
nor U19396 (N_19396,N_19047,N_19225);
xnor U19397 (N_19397,N_19125,N_19207);
nand U19398 (N_19398,N_19247,N_19007);
nand U19399 (N_19399,N_19186,N_19247);
and U19400 (N_19400,N_19159,N_19135);
and U19401 (N_19401,N_19000,N_19199);
nor U19402 (N_19402,N_19038,N_19046);
nand U19403 (N_19403,N_19126,N_19052);
nand U19404 (N_19404,N_19175,N_19185);
xnor U19405 (N_19405,N_19197,N_19225);
nand U19406 (N_19406,N_19135,N_19079);
xnor U19407 (N_19407,N_19157,N_19222);
or U19408 (N_19408,N_19004,N_19240);
or U19409 (N_19409,N_19089,N_19182);
and U19410 (N_19410,N_19044,N_19179);
nor U19411 (N_19411,N_19008,N_19146);
nor U19412 (N_19412,N_19083,N_19060);
xnor U19413 (N_19413,N_19182,N_19154);
nor U19414 (N_19414,N_19172,N_19038);
or U19415 (N_19415,N_19156,N_19057);
xor U19416 (N_19416,N_19230,N_19146);
nor U19417 (N_19417,N_19244,N_19139);
or U19418 (N_19418,N_19053,N_19061);
xnor U19419 (N_19419,N_19216,N_19197);
and U19420 (N_19420,N_19221,N_19247);
and U19421 (N_19421,N_19042,N_19018);
and U19422 (N_19422,N_19067,N_19046);
xnor U19423 (N_19423,N_19201,N_19075);
xnor U19424 (N_19424,N_19063,N_19123);
nor U19425 (N_19425,N_19121,N_19134);
or U19426 (N_19426,N_19105,N_19014);
xor U19427 (N_19427,N_19155,N_19005);
nand U19428 (N_19428,N_19185,N_19146);
nand U19429 (N_19429,N_19143,N_19074);
nor U19430 (N_19430,N_19002,N_19233);
nor U19431 (N_19431,N_19002,N_19160);
xor U19432 (N_19432,N_19162,N_19057);
nand U19433 (N_19433,N_19039,N_19109);
nand U19434 (N_19434,N_19214,N_19053);
and U19435 (N_19435,N_19164,N_19153);
xor U19436 (N_19436,N_19087,N_19012);
nor U19437 (N_19437,N_19122,N_19032);
or U19438 (N_19438,N_19223,N_19193);
nand U19439 (N_19439,N_19118,N_19148);
and U19440 (N_19440,N_19106,N_19237);
nor U19441 (N_19441,N_19165,N_19176);
nor U19442 (N_19442,N_19055,N_19108);
nor U19443 (N_19443,N_19024,N_19228);
xor U19444 (N_19444,N_19060,N_19157);
and U19445 (N_19445,N_19102,N_19123);
and U19446 (N_19446,N_19027,N_19139);
xor U19447 (N_19447,N_19002,N_19239);
or U19448 (N_19448,N_19165,N_19037);
or U19449 (N_19449,N_19099,N_19197);
or U19450 (N_19450,N_19205,N_19000);
or U19451 (N_19451,N_19057,N_19158);
or U19452 (N_19452,N_19045,N_19007);
xor U19453 (N_19453,N_19151,N_19215);
or U19454 (N_19454,N_19078,N_19119);
nand U19455 (N_19455,N_19227,N_19182);
nor U19456 (N_19456,N_19013,N_19238);
nor U19457 (N_19457,N_19008,N_19084);
xnor U19458 (N_19458,N_19237,N_19059);
nor U19459 (N_19459,N_19193,N_19089);
nor U19460 (N_19460,N_19132,N_19135);
and U19461 (N_19461,N_19127,N_19150);
and U19462 (N_19462,N_19054,N_19146);
and U19463 (N_19463,N_19077,N_19201);
nand U19464 (N_19464,N_19209,N_19180);
or U19465 (N_19465,N_19114,N_19160);
or U19466 (N_19466,N_19183,N_19008);
xnor U19467 (N_19467,N_19160,N_19061);
nand U19468 (N_19468,N_19171,N_19131);
or U19469 (N_19469,N_19193,N_19013);
nand U19470 (N_19470,N_19015,N_19086);
nand U19471 (N_19471,N_19249,N_19174);
xnor U19472 (N_19472,N_19162,N_19035);
or U19473 (N_19473,N_19195,N_19129);
nor U19474 (N_19474,N_19158,N_19093);
and U19475 (N_19475,N_19108,N_19048);
nand U19476 (N_19476,N_19220,N_19140);
or U19477 (N_19477,N_19018,N_19248);
xnor U19478 (N_19478,N_19067,N_19223);
xor U19479 (N_19479,N_19098,N_19038);
nor U19480 (N_19480,N_19233,N_19246);
xor U19481 (N_19481,N_19011,N_19099);
nor U19482 (N_19482,N_19013,N_19160);
xnor U19483 (N_19483,N_19156,N_19061);
and U19484 (N_19484,N_19188,N_19147);
and U19485 (N_19485,N_19194,N_19009);
or U19486 (N_19486,N_19027,N_19187);
nand U19487 (N_19487,N_19186,N_19138);
and U19488 (N_19488,N_19225,N_19056);
nand U19489 (N_19489,N_19171,N_19168);
nand U19490 (N_19490,N_19212,N_19041);
nand U19491 (N_19491,N_19100,N_19112);
nand U19492 (N_19492,N_19162,N_19242);
nor U19493 (N_19493,N_19186,N_19097);
or U19494 (N_19494,N_19204,N_19186);
nand U19495 (N_19495,N_19168,N_19049);
and U19496 (N_19496,N_19182,N_19166);
nand U19497 (N_19497,N_19029,N_19150);
nand U19498 (N_19498,N_19097,N_19172);
or U19499 (N_19499,N_19057,N_19203);
or U19500 (N_19500,N_19399,N_19312);
nand U19501 (N_19501,N_19317,N_19320);
or U19502 (N_19502,N_19323,N_19290);
nand U19503 (N_19503,N_19345,N_19339);
and U19504 (N_19504,N_19456,N_19461);
xor U19505 (N_19505,N_19486,N_19369);
and U19506 (N_19506,N_19485,N_19268);
nand U19507 (N_19507,N_19492,N_19370);
or U19508 (N_19508,N_19460,N_19340);
xnor U19509 (N_19509,N_19360,N_19447);
nand U19510 (N_19510,N_19310,N_19455);
xnor U19511 (N_19511,N_19436,N_19265);
nor U19512 (N_19512,N_19349,N_19273);
nor U19513 (N_19513,N_19391,N_19427);
nand U19514 (N_19514,N_19338,N_19477);
and U19515 (N_19515,N_19352,N_19286);
xor U19516 (N_19516,N_19300,N_19260);
nor U19517 (N_19517,N_19489,N_19495);
or U19518 (N_19518,N_19258,N_19481);
or U19519 (N_19519,N_19269,N_19379);
xnor U19520 (N_19520,N_19403,N_19380);
or U19521 (N_19521,N_19498,N_19424);
nor U19522 (N_19522,N_19421,N_19362);
nand U19523 (N_19523,N_19284,N_19439);
and U19524 (N_19524,N_19448,N_19425);
and U19525 (N_19525,N_19444,N_19253);
or U19526 (N_19526,N_19388,N_19264);
nor U19527 (N_19527,N_19346,N_19442);
nor U19528 (N_19528,N_19306,N_19381);
nand U19529 (N_19529,N_19304,N_19356);
and U19530 (N_19530,N_19416,N_19285);
and U19531 (N_19531,N_19333,N_19266);
nor U19532 (N_19532,N_19279,N_19445);
nor U19533 (N_19533,N_19329,N_19396);
nand U19534 (N_19534,N_19301,N_19468);
and U19535 (N_19535,N_19252,N_19274);
or U19536 (N_19536,N_19365,N_19366);
or U19537 (N_19537,N_19457,N_19420);
nand U19538 (N_19538,N_19450,N_19400);
nand U19539 (N_19539,N_19355,N_19322);
nand U19540 (N_19540,N_19401,N_19411);
and U19541 (N_19541,N_19465,N_19282);
and U19542 (N_19542,N_19354,N_19415);
xor U19543 (N_19543,N_19383,N_19350);
and U19544 (N_19544,N_19307,N_19288);
xnor U19545 (N_19545,N_19315,N_19385);
nor U19546 (N_19546,N_19446,N_19433);
nand U19547 (N_19547,N_19407,N_19335);
and U19548 (N_19548,N_19499,N_19294);
nand U19549 (N_19549,N_19287,N_19261);
or U19550 (N_19550,N_19372,N_19490);
nor U19551 (N_19551,N_19437,N_19363);
xnor U19552 (N_19552,N_19262,N_19434);
and U19553 (N_19553,N_19475,N_19443);
or U19554 (N_19554,N_19466,N_19484);
or U19555 (N_19555,N_19334,N_19324);
nand U19556 (N_19556,N_19493,N_19358);
nand U19557 (N_19557,N_19394,N_19361);
nor U19558 (N_19558,N_19257,N_19298);
xnor U19559 (N_19559,N_19326,N_19478);
and U19560 (N_19560,N_19470,N_19325);
nand U19561 (N_19561,N_19263,N_19308);
xnor U19562 (N_19562,N_19480,N_19463);
or U19563 (N_19563,N_19458,N_19395);
xor U19564 (N_19564,N_19452,N_19410);
xor U19565 (N_19565,N_19289,N_19336);
or U19566 (N_19566,N_19429,N_19293);
nor U19567 (N_19567,N_19494,N_19419);
nand U19568 (N_19568,N_19296,N_19454);
or U19569 (N_19569,N_19283,N_19471);
or U19570 (N_19570,N_19297,N_19414);
or U19571 (N_19571,N_19319,N_19314);
and U19572 (N_19572,N_19343,N_19344);
or U19573 (N_19573,N_19377,N_19311);
nor U19574 (N_19574,N_19422,N_19408);
nand U19575 (N_19575,N_19390,N_19412);
nor U19576 (N_19576,N_19278,N_19459);
and U19577 (N_19577,N_19382,N_19341);
and U19578 (N_19578,N_19357,N_19426);
xor U19579 (N_19579,N_19280,N_19402);
or U19580 (N_19580,N_19389,N_19386);
and U19581 (N_19581,N_19413,N_19272);
and U19582 (N_19582,N_19467,N_19309);
and U19583 (N_19583,N_19368,N_19250);
xor U19584 (N_19584,N_19430,N_19275);
and U19585 (N_19585,N_19404,N_19378);
nor U19586 (N_19586,N_19438,N_19418);
nor U19587 (N_19587,N_19276,N_19337);
nand U19588 (N_19588,N_19267,N_19487);
nor U19589 (N_19589,N_19330,N_19318);
nor U19590 (N_19590,N_19496,N_19299);
and U19591 (N_19591,N_19351,N_19367);
xor U19592 (N_19592,N_19464,N_19392);
nand U19593 (N_19593,N_19479,N_19374);
nand U19594 (N_19594,N_19393,N_19302);
nor U19595 (N_19595,N_19321,N_19347);
xnor U19596 (N_19596,N_19431,N_19488);
nor U19597 (N_19597,N_19295,N_19359);
and U19598 (N_19598,N_19441,N_19474);
nor U19599 (N_19599,N_19476,N_19406);
and U19600 (N_19600,N_19255,N_19482);
nor U19601 (N_19601,N_19423,N_19472);
xor U19602 (N_19602,N_19259,N_19364);
and U19603 (N_19603,N_19270,N_19398);
or U19604 (N_19604,N_19353,N_19428);
nor U19605 (N_19605,N_19348,N_19291);
nand U19606 (N_19606,N_19331,N_19483);
xor U19607 (N_19607,N_19373,N_19342);
and U19608 (N_19608,N_19277,N_19449);
nand U19609 (N_19609,N_19256,N_19405);
xor U19610 (N_19610,N_19305,N_19303);
or U19611 (N_19611,N_19409,N_19313);
or U19612 (N_19612,N_19328,N_19473);
nor U19613 (N_19613,N_19453,N_19491);
or U19614 (N_19614,N_19251,N_19327);
or U19615 (N_19615,N_19451,N_19316);
or U19616 (N_19616,N_19254,N_19397);
nor U19617 (N_19617,N_19435,N_19387);
and U19618 (N_19618,N_19292,N_19469);
nand U19619 (N_19619,N_19432,N_19440);
or U19620 (N_19620,N_19497,N_19375);
and U19621 (N_19621,N_19384,N_19271);
or U19622 (N_19622,N_19376,N_19417);
nand U19623 (N_19623,N_19281,N_19371);
or U19624 (N_19624,N_19332,N_19462);
or U19625 (N_19625,N_19449,N_19424);
xnor U19626 (N_19626,N_19463,N_19375);
xnor U19627 (N_19627,N_19460,N_19343);
nor U19628 (N_19628,N_19251,N_19478);
and U19629 (N_19629,N_19439,N_19431);
nor U19630 (N_19630,N_19494,N_19267);
and U19631 (N_19631,N_19361,N_19344);
nor U19632 (N_19632,N_19492,N_19429);
xor U19633 (N_19633,N_19288,N_19252);
or U19634 (N_19634,N_19424,N_19492);
or U19635 (N_19635,N_19275,N_19441);
nor U19636 (N_19636,N_19326,N_19312);
and U19637 (N_19637,N_19453,N_19433);
nor U19638 (N_19638,N_19492,N_19365);
xor U19639 (N_19639,N_19467,N_19470);
nor U19640 (N_19640,N_19491,N_19494);
nor U19641 (N_19641,N_19254,N_19386);
nor U19642 (N_19642,N_19450,N_19347);
or U19643 (N_19643,N_19473,N_19492);
and U19644 (N_19644,N_19323,N_19307);
xor U19645 (N_19645,N_19326,N_19464);
nor U19646 (N_19646,N_19315,N_19320);
nor U19647 (N_19647,N_19467,N_19405);
nor U19648 (N_19648,N_19440,N_19441);
xnor U19649 (N_19649,N_19281,N_19263);
nand U19650 (N_19650,N_19275,N_19487);
and U19651 (N_19651,N_19412,N_19259);
and U19652 (N_19652,N_19272,N_19267);
nand U19653 (N_19653,N_19432,N_19457);
and U19654 (N_19654,N_19487,N_19423);
nand U19655 (N_19655,N_19266,N_19419);
xor U19656 (N_19656,N_19374,N_19278);
or U19657 (N_19657,N_19418,N_19331);
nand U19658 (N_19658,N_19332,N_19340);
or U19659 (N_19659,N_19475,N_19455);
xor U19660 (N_19660,N_19286,N_19290);
or U19661 (N_19661,N_19474,N_19272);
xor U19662 (N_19662,N_19302,N_19499);
nor U19663 (N_19663,N_19412,N_19404);
nor U19664 (N_19664,N_19343,N_19353);
nor U19665 (N_19665,N_19496,N_19464);
xor U19666 (N_19666,N_19378,N_19440);
and U19667 (N_19667,N_19296,N_19286);
and U19668 (N_19668,N_19250,N_19488);
nand U19669 (N_19669,N_19361,N_19437);
and U19670 (N_19670,N_19268,N_19341);
nor U19671 (N_19671,N_19327,N_19485);
xor U19672 (N_19672,N_19270,N_19312);
xor U19673 (N_19673,N_19408,N_19380);
nor U19674 (N_19674,N_19460,N_19367);
xnor U19675 (N_19675,N_19489,N_19441);
or U19676 (N_19676,N_19381,N_19480);
nor U19677 (N_19677,N_19453,N_19324);
or U19678 (N_19678,N_19268,N_19396);
nor U19679 (N_19679,N_19368,N_19461);
xor U19680 (N_19680,N_19252,N_19492);
xnor U19681 (N_19681,N_19498,N_19490);
and U19682 (N_19682,N_19342,N_19261);
nor U19683 (N_19683,N_19313,N_19439);
nor U19684 (N_19684,N_19343,N_19411);
or U19685 (N_19685,N_19496,N_19427);
xnor U19686 (N_19686,N_19456,N_19489);
or U19687 (N_19687,N_19499,N_19380);
and U19688 (N_19688,N_19382,N_19347);
nand U19689 (N_19689,N_19363,N_19300);
xor U19690 (N_19690,N_19334,N_19361);
or U19691 (N_19691,N_19280,N_19429);
or U19692 (N_19692,N_19477,N_19291);
and U19693 (N_19693,N_19487,N_19309);
or U19694 (N_19694,N_19312,N_19413);
nor U19695 (N_19695,N_19372,N_19423);
and U19696 (N_19696,N_19327,N_19407);
nor U19697 (N_19697,N_19420,N_19424);
xor U19698 (N_19698,N_19274,N_19434);
xor U19699 (N_19699,N_19329,N_19491);
xor U19700 (N_19700,N_19315,N_19413);
and U19701 (N_19701,N_19330,N_19465);
xnor U19702 (N_19702,N_19329,N_19418);
xnor U19703 (N_19703,N_19406,N_19255);
or U19704 (N_19704,N_19466,N_19313);
or U19705 (N_19705,N_19373,N_19265);
nor U19706 (N_19706,N_19453,N_19319);
nand U19707 (N_19707,N_19378,N_19476);
nand U19708 (N_19708,N_19429,N_19398);
nand U19709 (N_19709,N_19498,N_19373);
nand U19710 (N_19710,N_19353,N_19324);
nand U19711 (N_19711,N_19316,N_19262);
or U19712 (N_19712,N_19358,N_19287);
xnor U19713 (N_19713,N_19367,N_19343);
and U19714 (N_19714,N_19308,N_19290);
and U19715 (N_19715,N_19268,N_19331);
nand U19716 (N_19716,N_19494,N_19492);
xnor U19717 (N_19717,N_19346,N_19476);
nand U19718 (N_19718,N_19451,N_19428);
nand U19719 (N_19719,N_19421,N_19461);
nand U19720 (N_19720,N_19397,N_19301);
xnor U19721 (N_19721,N_19352,N_19267);
and U19722 (N_19722,N_19252,N_19399);
nand U19723 (N_19723,N_19349,N_19252);
nand U19724 (N_19724,N_19384,N_19479);
nand U19725 (N_19725,N_19311,N_19483);
xor U19726 (N_19726,N_19446,N_19448);
or U19727 (N_19727,N_19363,N_19484);
or U19728 (N_19728,N_19373,N_19318);
nand U19729 (N_19729,N_19304,N_19435);
xnor U19730 (N_19730,N_19427,N_19400);
and U19731 (N_19731,N_19336,N_19434);
nand U19732 (N_19732,N_19358,N_19254);
nand U19733 (N_19733,N_19314,N_19349);
nor U19734 (N_19734,N_19429,N_19404);
or U19735 (N_19735,N_19302,N_19253);
nor U19736 (N_19736,N_19391,N_19337);
xnor U19737 (N_19737,N_19310,N_19257);
nor U19738 (N_19738,N_19476,N_19421);
nand U19739 (N_19739,N_19401,N_19423);
and U19740 (N_19740,N_19467,N_19319);
nand U19741 (N_19741,N_19277,N_19473);
or U19742 (N_19742,N_19284,N_19425);
and U19743 (N_19743,N_19480,N_19275);
xnor U19744 (N_19744,N_19427,N_19473);
nand U19745 (N_19745,N_19476,N_19479);
nand U19746 (N_19746,N_19322,N_19458);
and U19747 (N_19747,N_19461,N_19328);
or U19748 (N_19748,N_19482,N_19323);
and U19749 (N_19749,N_19344,N_19272);
or U19750 (N_19750,N_19621,N_19566);
nand U19751 (N_19751,N_19653,N_19584);
nor U19752 (N_19752,N_19542,N_19635);
xnor U19753 (N_19753,N_19689,N_19527);
nand U19754 (N_19754,N_19615,N_19719);
nand U19755 (N_19755,N_19531,N_19565);
or U19756 (N_19756,N_19613,N_19505);
xor U19757 (N_19757,N_19659,N_19504);
and U19758 (N_19758,N_19521,N_19548);
and U19759 (N_19759,N_19559,N_19603);
xnor U19760 (N_19760,N_19668,N_19681);
xor U19761 (N_19761,N_19647,N_19502);
xnor U19762 (N_19762,N_19720,N_19725);
nor U19763 (N_19763,N_19693,N_19588);
nand U19764 (N_19764,N_19656,N_19544);
xnor U19765 (N_19765,N_19590,N_19508);
or U19766 (N_19766,N_19589,N_19545);
xnor U19767 (N_19767,N_19537,N_19543);
nand U19768 (N_19768,N_19575,N_19553);
nand U19769 (N_19769,N_19726,N_19688);
xnor U19770 (N_19770,N_19662,N_19592);
xnor U19771 (N_19771,N_19516,N_19650);
or U19772 (N_19772,N_19706,N_19591);
nor U19773 (N_19773,N_19711,N_19517);
nor U19774 (N_19774,N_19707,N_19538);
xnor U19775 (N_19775,N_19649,N_19604);
nor U19776 (N_19776,N_19637,N_19568);
nor U19777 (N_19777,N_19666,N_19593);
xnor U19778 (N_19778,N_19709,N_19510);
nand U19779 (N_19779,N_19539,N_19571);
or U19780 (N_19780,N_19535,N_19675);
and U19781 (N_19781,N_19680,N_19525);
and U19782 (N_19782,N_19500,N_19570);
nand U19783 (N_19783,N_19617,N_19567);
nand U19784 (N_19784,N_19587,N_19651);
nor U19785 (N_19785,N_19550,N_19741);
xnor U19786 (N_19786,N_19736,N_19702);
xnor U19787 (N_19787,N_19507,N_19514);
nor U19788 (N_19788,N_19515,N_19657);
and U19789 (N_19789,N_19534,N_19669);
and U19790 (N_19790,N_19735,N_19679);
or U19791 (N_19791,N_19581,N_19512);
or U19792 (N_19792,N_19556,N_19547);
or U19793 (N_19793,N_19583,N_19697);
xor U19794 (N_19794,N_19729,N_19541);
nand U19795 (N_19795,N_19602,N_19718);
nor U19796 (N_19796,N_19749,N_19745);
nand U19797 (N_19797,N_19742,N_19564);
and U19798 (N_19798,N_19686,N_19738);
nor U19799 (N_19799,N_19616,N_19552);
and U19800 (N_19800,N_19608,N_19610);
or U19801 (N_19801,N_19597,N_19578);
and U19802 (N_19802,N_19577,N_19727);
and U19803 (N_19803,N_19596,N_19579);
and U19804 (N_19804,N_19580,N_19696);
xnor U19805 (N_19805,N_19663,N_19710);
nand U19806 (N_19806,N_19661,N_19678);
or U19807 (N_19807,N_19682,N_19572);
nor U19808 (N_19808,N_19609,N_19713);
nor U19809 (N_19809,N_19503,N_19739);
xor U19810 (N_19810,N_19730,N_19555);
and U19811 (N_19811,N_19665,N_19594);
nand U19812 (N_19812,N_19618,N_19501);
and U19813 (N_19813,N_19700,N_19694);
nor U19814 (N_19814,N_19513,N_19532);
and U19815 (N_19815,N_19554,N_19582);
nor U19816 (N_19816,N_19667,N_19626);
and U19817 (N_19817,N_19728,N_19524);
xnor U19818 (N_19818,N_19598,N_19683);
and U19819 (N_19819,N_19530,N_19714);
xnor U19820 (N_19820,N_19712,N_19641);
and U19821 (N_19821,N_19574,N_19721);
nand U19822 (N_19822,N_19743,N_19573);
xnor U19823 (N_19823,N_19642,N_19648);
or U19824 (N_19824,N_19607,N_19640);
xnor U19825 (N_19825,N_19606,N_19520);
nor U19826 (N_19826,N_19732,N_19747);
xnor U19827 (N_19827,N_19644,N_19601);
nor U19828 (N_19828,N_19599,N_19660);
and U19829 (N_19829,N_19698,N_19562);
or U19830 (N_19830,N_19687,N_19529);
xor U19831 (N_19831,N_19646,N_19672);
and U19832 (N_19832,N_19655,N_19708);
and U19833 (N_19833,N_19563,N_19540);
xnor U19834 (N_19834,N_19585,N_19674);
and U19835 (N_19835,N_19723,N_19724);
and U19836 (N_19836,N_19619,N_19734);
and U19837 (N_19837,N_19628,N_19627);
nor U19838 (N_19838,N_19636,N_19701);
or U19839 (N_19839,N_19549,N_19671);
nand U19840 (N_19840,N_19676,N_19528);
or U19841 (N_19841,N_19731,N_19611);
nor U19842 (N_19842,N_19634,N_19595);
nor U19843 (N_19843,N_19620,N_19526);
and U19844 (N_19844,N_19643,N_19658);
nor U19845 (N_19845,N_19685,N_19737);
xnor U19846 (N_19846,N_19673,N_19690);
and U19847 (N_19847,N_19740,N_19677);
nor U19848 (N_19848,N_19561,N_19518);
or U19849 (N_19849,N_19654,N_19546);
nand U19850 (N_19850,N_19605,N_19509);
and U19851 (N_19851,N_19746,N_19632);
and U19852 (N_19852,N_19576,N_19631);
or U19853 (N_19853,N_19633,N_19522);
or U19854 (N_19854,N_19625,N_19684);
nor U19855 (N_19855,N_19704,N_19511);
nor U19856 (N_19856,N_19705,N_19569);
nand U19857 (N_19857,N_19722,N_19614);
xor U19858 (N_19858,N_19519,N_19699);
or U19859 (N_19859,N_19600,N_19630);
xnor U19860 (N_19860,N_19691,N_19695);
and U19861 (N_19861,N_19664,N_19558);
nor U19862 (N_19862,N_19523,N_19670);
nor U19863 (N_19863,N_19692,N_19717);
or U19864 (N_19864,N_19638,N_19533);
nand U19865 (N_19865,N_19716,N_19645);
or U19866 (N_19866,N_19612,N_19748);
xor U19867 (N_19867,N_19560,N_19629);
xnor U19868 (N_19868,N_19536,N_19703);
or U19869 (N_19869,N_19622,N_19623);
and U19870 (N_19870,N_19715,N_19557);
or U19871 (N_19871,N_19744,N_19639);
nand U19872 (N_19872,N_19733,N_19624);
nor U19873 (N_19873,N_19586,N_19506);
nor U19874 (N_19874,N_19551,N_19652);
and U19875 (N_19875,N_19635,N_19615);
and U19876 (N_19876,N_19742,N_19509);
and U19877 (N_19877,N_19547,N_19599);
and U19878 (N_19878,N_19634,N_19605);
nor U19879 (N_19879,N_19605,N_19510);
xor U19880 (N_19880,N_19559,N_19514);
nor U19881 (N_19881,N_19623,N_19627);
and U19882 (N_19882,N_19580,N_19702);
nand U19883 (N_19883,N_19742,N_19706);
and U19884 (N_19884,N_19541,N_19554);
nand U19885 (N_19885,N_19662,N_19720);
or U19886 (N_19886,N_19508,N_19556);
nor U19887 (N_19887,N_19534,N_19559);
nand U19888 (N_19888,N_19717,N_19577);
xor U19889 (N_19889,N_19694,N_19609);
or U19890 (N_19890,N_19568,N_19683);
or U19891 (N_19891,N_19600,N_19667);
nor U19892 (N_19892,N_19722,N_19627);
nor U19893 (N_19893,N_19737,N_19688);
or U19894 (N_19894,N_19719,N_19689);
nor U19895 (N_19895,N_19655,N_19580);
nand U19896 (N_19896,N_19530,N_19694);
xor U19897 (N_19897,N_19521,N_19720);
or U19898 (N_19898,N_19608,N_19692);
or U19899 (N_19899,N_19584,N_19517);
nor U19900 (N_19900,N_19668,N_19736);
xnor U19901 (N_19901,N_19736,N_19529);
nand U19902 (N_19902,N_19571,N_19677);
or U19903 (N_19903,N_19749,N_19578);
nand U19904 (N_19904,N_19695,N_19602);
nor U19905 (N_19905,N_19734,N_19534);
xor U19906 (N_19906,N_19694,N_19632);
nor U19907 (N_19907,N_19724,N_19631);
and U19908 (N_19908,N_19710,N_19569);
xnor U19909 (N_19909,N_19631,N_19708);
xor U19910 (N_19910,N_19640,N_19681);
nor U19911 (N_19911,N_19572,N_19591);
or U19912 (N_19912,N_19527,N_19662);
or U19913 (N_19913,N_19534,N_19737);
or U19914 (N_19914,N_19561,N_19601);
or U19915 (N_19915,N_19740,N_19678);
or U19916 (N_19916,N_19686,N_19571);
and U19917 (N_19917,N_19686,N_19735);
or U19918 (N_19918,N_19544,N_19541);
or U19919 (N_19919,N_19716,N_19558);
nor U19920 (N_19920,N_19707,N_19619);
xnor U19921 (N_19921,N_19649,N_19643);
xor U19922 (N_19922,N_19741,N_19570);
nor U19923 (N_19923,N_19656,N_19527);
nand U19924 (N_19924,N_19551,N_19596);
and U19925 (N_19925,N_19655,N_19522);
and U19926 (N_19926,N_19676,N_19601);
nor U19927 (N_19927,N_19516,N_19718);
nand U19928 (N_19928,N_19652,N_19736);
xor U19929 (N_19929,N_19611,N_19575);
xor U19930 (N_19930,N_19693,N_19540);
xnor U19931 (N_19931,N_19633,N_19651);
or U19932 (N_19932,N_19707,N_19674);
nor U19933 (N_19933,N_19520,N_19649);
or U19934 (N_19934,N_19702,N_19660);
nand U19935 (N_19935,N_19529,N_19701);
and U19936 (N_19936,N_19630,N_19656);
and U19937 (N_19937,N_19598,N_19718);
or U19938 (N_19938,N_19709,N_19582);
or U19939 (N_19939,N_19578,N_19734);
xor U19940 (N_19940,N_19588,N_19696);
and U19941 (N_19941,N_19634,N_19540);
nand U19942 (N_19942,N_19635,N_19562);
nand U19943 (N_19943,N_19575,N_19562);
or U19944 (N_19944,N_19711,N_19507);
and U19945 (N_19945,N_19650,N_19748);
xor U19946 (N_19946,N_19664,N_19640);
nor U19947 (N_19947,N_19688,N_19685);
xor U19948 (N_19948,N_19649,N_19677);
nor U19949 (N_19949,N_19656,N_19501);
and U19950 (N_19950,N_19510,N_19748);
or U19951 (N_19951,N_19626,N_19572);
or U19952 (N_19952,N_19666,N_19545);
and U19953 (N_19953,N_19568,N_19691);
nand U19954 (N_19954,N_19643,N_19502);
nor U19955 (N_19955,N_19550,N_19549);
or U19956 (N_19956,N_19652,N_19655);
and U19957 (N_19957,N_19681,N_19624);
or U19958 (N_19958,N_19542,N_19734);
and U19959 (N_19959,N_19692,N_19703);
and U19960 (N_19960,N_19540,N_19742);
nor U19961 (N_19961,N_19716,N_19735);
xnor U19962 (N_19962,N_19685,N_19607);
nor U19963 (N_19963,N_19659,N_19706);
xnor U19964 (N_19964,N_19576,N_19602);
nand U19965 (N_19965,N_19669,N_19658);
nand U19966 (N_19966,N_19537,N_19749);
and U19967 (N_19967,N_19654,N_19602);
or U19968 (N_19968,N_19744,N_19671);
nand U19969 (N_19969,N_19686,N_19526);
or U19970 (N_19970,N_19555,N_19630);
and U19971 (N_19971,N_19594,N_19714);
xor U19972 (N_19972,N_19516,N_19551);
nor U19973 (N_19973,N_19616,N_19608);
xor U19974 (N_19974,N_19591,N_19623);
and U19975 (N_19975,N_19680,N_19730);
and U19976 (N_19976,N_19570,N_19565);
nor U19977 (N_19977,N_19628,N_19517);
nor U19978 (N_19978,N_19654,N_19549);
nand U19979 (N_19979,N_19746,N_19637);
or U19980 (N_19980,N_19581,N_19645);
and U19981 (N_19981,N_19591,N_19503);
nand U19982 (N_19982,N_19680,N_19618);
and U19983 (N_19983,N_19533,N_19544);
nand U19984 (N_19984,N_19744,N_19723);
or U19985 (N_19985,N_19728,N_19525);
nand U19986 (N_19986,N_19521,N_19735);
nand U19987 (N_19987,N_19581,N_19657);
xnor U19988 (N_19988,N_19522,N_19682);
nor U19989 (N_19989,N_19652,N_19739);
nor U19990 (N_19990,N_19523,N_19502);
xnor U19991 (N_19991,N_19685,N_19623);
or U19992 (N_19992,N_19526,N_19639);
and U19993 (N_19993,N_19584,N_19623);
or U19994 (N_19994,N_19575,N_19528);
nor U19995 (N_19995,N_19532,N_19551);
xor U19996 (N_19996,N_19521,N_19743);
and U19997 (N_19997,N_19536,N_19732);
nor U19998 (N_19998,N_19619,N_19645);
and U19999 (N_19999,N_19505,N_19681);
nand UO_0 (O_0,N_19761,N_19914);
nor UO_1 (O_1,N_19945,N_19812);
nand UO_2 (O_2,N_19895,N_19920);
nor UO_3 (O_3,N_19906,N_19881);
or UO_4 (O_4,N_19849,N_19868);
and UO_5 (O_5,N_19927,N_19925);
nor UO_6 (O_6,N_19976,N_19896);
nor UO_7 (O_7,N_19969,N_19891);
nor UO_8 (O_8,N_19943,N_19955);
and UO_9 (O_9,N_19781,N_19785);
nor UO_10 (O_10,N_19915,N_19751);
or UO_11 (O_11,N_19837,N_19764);
and UO_12 (O_12,N_19942,N_19949);
nand UO_13 (O_13,N_19898,N_19900);
xnor UO_14 (O_14,N_19816,N_19829);
and UO_15 (O_15,N_19833,N_19804);
xnor UO_16 (O_16,N_19771,N_19779);
or UO_17 (O_17,N_19784,N_19758);
xnor UO_18 (O_18,N_19913,N_19807);
and UO_19 (O_19,N_19924,N_19893);
and UO_20 (O_20,N_19912,N_19865);
or UO_21 (O_21,N_19994,N_19933);
nand UO_22 (O_22,N_19767,N_19902);
nand UO_23 (O_23,N_19797,N_19862);
nand UO_24 (O_24,N_19907,N_19793);
or UO_25 (O_25,N_19889,N_19860);
xnor UO_26 (O_26,N_19988,N_19997);
and UO_27 (O_27,N_19821,N_19773);
nand UO_28 (O_28,N_19871,N_19790);
and UO_29 (O_29,N_19929,N_19931);
and UO_30 (O_30,N_19867,N_19956);
nor UO_31 (O_31,N_19753,N_19822);
xnor UO_32 (O_32,N_19855,N_19880);
and UO_33 (O_33,N_19788,N_19783);
xnor UO_34 (O_34,N_19834,N_19778);
xnor UO_35 (O_35,N_19842,N_19810);
nor UO_36 (O_36,N_19869,N_19995);
or UO_37 (O_37,N_19996,N_19904);
xor UO_38 (O_38,N_19762,N_19879);
or UO_39 (O_39,N_19911,N_19886);
nand UO_40 (O_40,N_19755,N_19990);
or UO_41 (O_41,N_19872,N_19941);
nor UO_42 (O_42,N_19776,N_19859);
or UO_43 (O_43,N_19908,N_19918);
or UO_44 (O_44,N_19938,N_19809);
or UO_45 (O_45,N_19939,N_19883);
or UO_46 (O_46,N_19854,N_19806);
xnor UO_47 (O_47,N_19970,N_19839);
and UO_48 (O_48,N_19989,N_19866);
nor UO_49 (O_49,N_19968,N_19992);
or UO_50 (O_50,N_19818,N_19815);
and UO_51 (O_51,N_19825,N_19813);
and UO_52 (O_52,N_19979,N_19999);
xnor UO_53 (O_53,N_19917,N_19959);
nand UO_54 (O_54,N_19946,N_19986);
xor UO_55 (O_55,N_19921,N_19894);
xnor UO_56 (O_56,N_19841,N_19966);
nand UO_57 (O_57,N_19984,N_19763);
and UO_58 (O_58,N_19960,N_19888);
nor UO_59 (O_59,N_19885,N_19858);
xor UO_60 (O_60,N_19808,N_19802);
or UO_61 (O_61,N_19750,N_19847);
nand UO_62 (O_62,N_19948,N_19963);
or UO_63 (O_63,N_19974,N_19861);
and UO_64 (O_64,N_19853,N_19782);
nor UO_65 (O_65,N_19830,N_19798);
xor UO_66 (O_66,N_19982,N_19954);
and UO_67 (O_67,N_19874,N_19801);
nor UO_68 (O_68,N_19814,N_19774);
nand UO_69 (O_69,N_19940,N_19965);
nor UO_70 (O_70,N_19787,N_19851);
or UO_71 (O_71,N_19967,N_19897);
and UO_72 (O_72,N_19870,N_19971);
or UO_73 (O_73,N_19985,N_19786);
nor UO_74 (O_74,N_19775,N_19882);
and UO_75 (O_75,N_19823,N_19903);
xnor UO_76 (O_76,N_19757,N_19768);
and UO_77 (O_77,N_19811,N_19799);
and UO_78 (O_78,N_19972,N_19958);
nor UO_79 (O_79,N_19840,N_19832);
nor UO_80 (O_80,N_19791,N_19857);
xnor UO_81 (O_81,N_19877,N_19827);
and UO_82 (O_82,N_19919,N_19953);
nor UO_83 (O_83,N_19961,N_19901);
nor UO_84 (O_84,N_19887,N_19957);
nand UO_85 (O_85,N_19789,N_19973);
or UO_86 (O_86,N_19934,N_19846);
nor UO_87 (O_87,N_19844,N_19831);
nor UO_88 (O_88,N_19843,N_19993);
nor UO_89 (O_89,N_19852,N_19944);
or UO_90 (O_90,N_19777,N_19826);
nor UO_91 (O_91,N_19803,N_19952);
or UO_92 (O_92,N_19980,N_19765);
nor UO_93 (O_93,N_19937,N_19769);
and UO_94 (O_94,N_19795,N_19892);
or UO_95 (O_95,N_19962,N_19987);
or UO_96 (O_96,N_19800,N_19998);
xor UO_97 (O_97,N_19873,N_19876);
nor UO_98 (O_98,N_19752,N_19863);
or UO_99 (O_99,N_19964,N_19875);
xnor UO_100 (O_100,N_19910,N_19950);
and UO_101 (O_101,N_19981,N_19932);
or UO_102 (O_102,N_19850,N_19916);
xnor UO_103 (O_103,N_19796,N_19905);
or UO_104 (O_104,N_19770,N_19856);
and UO_105 (O_105,N_19923,N_19909);
xnor UO_106 (O_106,N_19805,N_19754);
or UO_107 (O_107,N_19884,N_19991);
nor UO_108 (O_108,N_19890,N_19978);
nor UO_109 (O_109,N_19928,N_19930);
nand UO_110 (O_110,N_19760,N_19824);
nand UO_111 (O_111,N_19947,N_19951);
nor UO_112 (O_112,N_19845,N_19975);
nor UO_113 (O_113,N_19838,N_19835);
and UO_114 (O_114,N_19936,N_19926);
or UO_115 (O_115,N_19766,N_19780);
or UO_116 (O_116,N_19772,N_19759);
or UO_117 (O_117,N_19836,N_19794);
and UO_118 (O_118,N_19848,N_19899);
or UO_119 (O_119,N_19864,N_19878);
nand UO_120 (O_120,N_19817,N_19977);
xnor UO_121 (O_121,N_19756,N_19922);
nand UO_122 (O_122,N_19792,N_19819);
or UO_123 (O_123,N_19983,N_19828);
nor UO_124 (O_124,N_19820,N_19935);
xnor UO_125 (O_125,N_19804,N_19847);
nor UO_126 (O_126,N_19998,N_19947);
nand UO_127 (O_127,N_19988,N_19929);
nand UO_128 (O_128,N_19842,N_19866);
xor UO_129 (O_129,N_19857,N_19849);
nor UO_130 (O_130,N_19956,N_19820);
or UO_131 (O_131,N_19836,N_19974);
and UO_132 (O_132,N_19818,N_19816);
and UO_133 (O_133,N_19780,N_19918);
and UO_134 (O_134,N_19869,N_19790);
nand UO_135 (O_135,N_19864,N_19789);
nor UO_136 (O_136,N_19947,N_19767);
nor UO_137 (O_137,N_19798,N_19989);
or UO_138 (O_138,N_19850,N_19760);
xnor UO_139 (O_139,N_19814,N_19842);
nor UO_140 (O_140,N_19887,N_19889);
nand UO_141 (O_141,N_19841,N_19922);
or UO_142 (O_142,N_19936,N_19912);
nor UO_143 (O_143,N_19789,N_19953);
nand UO_144 (O_144,N_19995,N_19979);
nor UO_145 (O_145,N_19823,N_19877);
or UO_146 (O_146,N_19784,N_19794);
and UO_147 (O_147,N_19887,N_19861);
or UO_148 (O_148,N_19803,N_19795);
nor UO_149 (O_149,N_19843,N_19869);
or UO_150 (O_150,N_19847,N_19989);
and UO_151 (O_151,N_19940,N_19924);
or UO_152 (O_152,N_19972,N_19925);
xnor UO_153 (O_153,N_19862,N_19832);
or UO_154 (O_154,N_19837,N_19868);
xor UO_155 (O_155,N_19940,N_19808);
nand UO_156 (O_156,N_19941,N_19830);
xnor UO_157 (O_157,N_19756,N_19885);
nand UO_158 (O_158,N_19937,N_19821);
nand UO_159 (O_159,N_19782,N_19993);
xor UO_160 (O_160,N_19854,N_19897);
and UO_161 (O_161,N_19814,N_19920);
nand UO_162 (O_162,N_19965,N_19904);
nor UO_163 (O_163,N_19949,N_19912);
xnor UO_164 (O_164,N_19979,N_19802);
nand UO_165 (O_165,N_19884,N_19817);
nand UO_166 (O_166,N_19984,N_19862);
or UO_167 (O_167,N_19918,N_19806);
or UO_168 (O_168,N_19930,N_19914);
xnor UO_169 (O_169,N_19816,N_19837);
xnor UO_170 (O_170,N_19778,N_19946);
nand UO_171 (O_171,N_19982,N_19986);
or UO_172 (O_172,N_19847,N_19940);
nor UO_173 (O_173,N_19804,N_19773);
and UO_174 (O_174,N_19914,N_19959);
nand UO_175 (O_175,N_19778,N_19815);
nand UO_176 (O_176,N_19936,N_19860);
nand UO_177 (O_177,N_19910,N_19828);
and UO_178 (O_178,N_19903,N_19923);
nor UO_179 (O_179,N_19977,N_19763);
or UO_180 (O_180,N_19999,N_19969);
and UO_181 (O_181,N_19994,N_19987);
or UO_182 (O_182,N_19804,N_19873);
and UO_183 (O_183,N_19908,N_19882);
and UO_184 (O_184,N_19809,N_19940);
nand UO_185 (O_185,N_19901,N_19990);
xor UO_186 (O_186,N_19989,N_19928);
and UO_187 (O_187,N_19850,N_19927);
and UO_188 (O_188,N_19779,N_19876);
nand UO_189 (O_189,N_19823,N_19998);
nor UO_190 (O_190,N_19781,N_19908);
or UO_191 (O_191,N_19779,N_19933);
or UO_192 (O_192,N_19877,N_19936);
nor UO_193 (O_193,N_19816,N_19950);
xor UO_194 (O_194,N_19797,N_19751);
or UO_195 (O_195,N_19813,N_19771);
nand UO_196 (O_196,N_19753,N_19845);
nor UO_197 (O_197,N_19854,N_19757);
nand UO_198 (O_198,N_19758,N_19873);
nor UO_199 (O_199,N_19794,N_19950);
and UO_200 (O_200,N_19906,N_19846);
or UO_201 (O_201,N_19923,N_19928);
or UO_202 (O_202,N_19831,N_19963);
nor UO_203 (O_203,N_19824,N_19811);
nor UO_204 (O_204,N_19849,N_19939);
and UO_205 (O_205,N_19795,N_19839);
or UO_206 (O_206,N_19776,N_19898);
xor UO_207 (O_207,N_19914,N_19924);
or UO_208 (O_208,N_19914,N_19963);
xor UO_209 (O_209,N_19993,N_19954);
or UO_210 (O_210,N_19891,N_19771);
or UO_211 (O_211,N_19855,N_19854);
nand UO_212 (O_212,N_19772,N_19825);
or UO_213 (O_213,N_19879,N_19792);
xnor UO_214 (O_214,N_19994,N_19938);
nor UO_215 (O_215,N_19958,N_19880);
or UO_216 (O_216,N_19982,N_19859);
and UO_217 (O_217,N_19985,N_19848);
nand UO_218 (O_218,N_19837,N_19999);
nor UO_219 (O_219,N_19810,N_19977);
xor UO_220 (O_220,N_19979,N_19785);
nand UO_221 (O_221,N_19822,N_19833);
nand UO_222 (O_222,N_19826,N_19958);
nor UO_223 (O_223,N_19916,N_19804);
nand UO_224 (O_224,N_19920,N_19925);
nand UO_225 (O_225,N_19885,N_19958);
xor UO_226 (O_226,N_19952,N_19958);
xnor UO_227 (O_227,N_19973,N_19980);
xor UO_228 (O_228,N_19851,N_19919);
and UO_229 (O_229,N_19963,N_19875);
nand UO_230 (O_230,N_19856,N_19911);
nor UO_231 (O_231,N_19760,N_19801);
or UO_232 (O_232,N_19911,N_19879);
nand UO_233 (O_233,N_19993,N_19933);
and UO_234 (O_234,N_19845,N_19860);
and UO_235 (O_235,N_19936,N_19762);
and UO_236 (O_236,N_19876,N_19808);
and UO_237 (O_237,N_19991,N_19957);
nor UO_238 (O_238,N_19937,N_19764);
and UO_239 (O_239,N_19935,N_19779);
xnor UO_240 (O_240,N_19924,N_19773);
or UO_241 (O_241,N_19816,N_19891);
or UO_242 (O_242,N_19835,N_19923);
xor UO_243 (O_243,N_19965,N_19916);
nand UO_244 (O_244,N_19995,N_19944);
and UO_245 (O_245,N_19818,N_19918);
and UO_246 (O_246,N_19961,N_19789);
nor UO_247 (O_247,N_19882,N_19838);
and UO_248 (O_248,N_19864,N_19782);
xnor UO_249 (O_249,N_19869,N_19912);
or UO_250 (O_250,N_19899,N_19889);
xnor UO_251 (O_251,N_19946,N_19850);
or UO_252 (O_252,N_19886,N_19794);
nor UO_253 (O_253,N_19816,N_19866);
nor UO_254 (O_254,N_19907,N_19816);
nor UO_255 (O_255,N_19999,N_19827);
or UO_256 (O_256,N_19800,N_19981);
and UO_257 (O_257,N_19965,N_19931);
nand UO_258 (O_258,N_19984,N_19894);
xor UO_259 (O_259,N_19874,N_19954);
nand UO_260 (O_260,N_19980,N_19871);
nand UO_261 (O_261,N_19934,N_19808);
and UO_262 (O_262,N_19973,N_19925);
nand UO_263 (O_263,N_19962,N_19834);
nand UO_264 (O_264,N_19764,N_19768);
xnor UO_265 (O_265,N_19883,N_19780);
nand UO_266 (O_266,N_19776,N_19814);
nand UO_267 (O_267,N_19873,N_19765);
or UO_268 (O_268,N_19839,N_19946);
nand UO_269 (O_269,N_19821,N_19851);
or UO_270 (O_270,N_19915,N_19805);
or UO_271 (O_271,N_19933,N_19834);
and UO_272 (O_272,N_19983,N_19964);
xnor UO_273 (O_273,N_19954,N_19926);
and UO_274 (O_274,N_19760,N_19952);
xnor UO_275 (O_275,N_19769,N_19924);
nand UO_276 (O_276,N_19964,N_19956);
nand UO_277 (O_277,N_19803,N_19766);
nand UO_278 (O_278,N_19983,N_19959);
xnor UO_279 (O_279,N_19750,N_19955);
nor UO_280 (O_280,N_19785,N_19844);
nand UO_281 (O_281,N_19920,N_19961);
nor UO_282 (O_282,N_19803,N_19869);
nand UO_283 (O_283,N_19891,N_19897);
or UO_284 (O_284,N_19910,N_19998);
or UO_285 (O_285,N_19826,N_19796);
and UO_286 (O_286,N_19816,N_19811);
xnor UO_287 (O_287,N_19898,N_19996);
xor UO_288 (O_288,N_19824,N_19988);
nor UO_289 (O_289,N_19987,N_19855);
xnor UO_290 (O_290,N_19814,N_19783);
or UO_291 (O_291,N_19813,N_19762);
or UO_292 (O_292,N_19924,N_19802);
or UO_293 (O_293,N_19870,N_19750);
nand UO_294 (O_294,N_19967,N_19996);
and UO_295 (O_295,N_19835,N_19946);
and UO_296 (O_296,N_19806,N_19995);
xor UO_297 (O_297,N_19804,N_19979);
or UO_298 (O_298,N_19798,N_19795);
nand UO_299 (O_299,N_19862,N_19836);
xor UO_300 (O_300,N_19756,N_19802);
or UO_301 (O_301,N_19784,N_19938);
xnor UO_302 (O_302,N_19783,N_19939);
or UO_303 (O_303,N_19767,N_19946);
and UO_304 (O_304,N_19892,N_19963);
xor UO_305 (O_305,N_19798,N_19842);
xnor UO_306 (O_306,N_19846,N_19826);
or UO_307 (O_307,N_19984,N_19973);
xor UO_308 (O_308,N_19751,N_19977);
and UO_309 (O_309,N_19788,N_19917);
nand UO_310 (O_310,N_19886,N_19785);
and UO_311 (O_311,N_19978,N_19790);
and UO_312 (O_312,N_19899,N_19983);
nand UO_313 (O_313,N_19754,N_19781);
nor UO_314 (O_314,N_19783,N_19925);
xnor UO_315 (O_315,N_19871,N_19775);
nand UO_316 (O_316,N_19990,N_19888);
nor UO_317 (O_317,N_19812,N_19835);
and UO_318 (O_318,N_19938,N_19803);
nor UO_319 (O_319,N_19771,N_19938);
or UO_320 (O_320,N_19754,N_19785);
nand UO_321 (O_321,N_19830,N_19822);
and UO_322 (O_322,N_19848,N_19755);
or UO_323 (O_323,N_19780,N_19929);
nand UO_324 (O_324,N_19827,N_19863);
nor UO_325 (O_325,N_19936,N_19939);
nand UO_326 (O_326,N_19789,N_19761);
nand UO_327 (O_327,N_19902,N_19780);
nor UO_328 (O_328,N_19880,N_19864);
xor UO_329 (O_329,N_19835,N_19850);
xnor UO_330 (O_330,N_19928,N_19819);
nor UO_331 (O_331,N_19764,N_19864);
nand UO_332 (O_332,N_19832,N_19903);
and UO_333 (O_333,N_19773,N_19944);
and UO_334 (O_334,N_19925,N_19851);
nand UO_335 (O_335,N_19955,N_19751);
xnor UO_336 (O_336,N_19796,N_19836);
nand UO_337 (O_337,N_19761,N_19892);
or UO_338 (O_338,N_19918,N_19882);
xor UO_339 (O_339,N_19902,N_19750);
xor UO_340 (O_340,N_19937,N_19832);
nor UO_341 (O_341,N_19788,N_19908);
and UO_342 (O_342,N_19832,N_19877);
and UO_343 (O_343,N_19782,N_19894);
or UO_344 (O_344,N_19772,N_19758);
and UO_345 (O_345,N_19919,N_19833);
nor UO_346 (O_346,N_19843,N_19759);
nand UO_347 (O_347,N_19813,N_19754);
xnor UO_348 (O_348,N_19754,N_19905);
and UO_349 (O_349,N_19916,N_19964);
and UO_350 (O_350,N_19932,N_19963);
or UO_351 (O_351,N_19756,N_19827);
xor UO_352 (O_352,N_19963,N_19961);
nand UO_353 (O_353,N_19813,N_19902);
nor UO_354 (O_354,N_19818,N_19761);
and UO_355 (O_355,N_19844,N_19932);
nor UO_356 (O_356,N_19753,N_19934);
xor UO_357 (O_357,N_19939,N_19865);
xor UO_358 (O_358,N_19792,N_19989);
nand UO_359 (O_359,N_19833,N_19828);
nand UO_360 (O_360,N_19751,N_19787);
and UO_361 (O_361,N_19956,N_19919);
or UO_362 (O_362,N_19788,N_19807);
or UO_363 (O_363,N_19888,N_19899);
xor UO_364 (O_364,N_19900,N_19929);
xnor UO_365 (O_365,N_19990,N_19839);
or UO_366 (O_366,N_19936,N_19770);
and UO_367 (O_367,N_19976,N_19924);
xor UO_368 (O_368,N_19803,N_19915);
nor UO_369 (O_369,N_19919,N_19945);
or UO_370 (O_370,N_19932,N_19794);
or UO_371 (O_371,N_19828,N_19889);
xor UO_372 (O_372,N_19814,N_19854);
nand UO_373 (O_373,N_19973,N_19801);
xnor UO_374 (O_374,N_19846,N_19944);
xnor UO_375 (O_375,N_19802,N_19830);
or UO_376 (O_376,N_19768,N_19914);
and UO_377 (O_377,N_19925,N_19966);
nand UO_378 (O_378,N_19995,N_19974);
xnor UO_379 (O_379,N_19764,N_19972);
or UO_380 (O_380,N_19797,N_19872);
nand UO_381 (O_381,N_19930,N_19802);
xnor UO_382 (O_382,N_19949,N_19783);
or UO_383 (O_383,N_19923,N_19854);
nor UO_384 (O_384,N_19910,N_19942);
and UO_385 (O_385,N_19900,N_19980);
and UO_386 (O_386,N_19866,N_19821);
nand UO_387 (O_387,N_19873,N_19827);
and UO_388 (O_388,N_19793,N_19833);
nor UO_389 (O_389,N_19837,N_19911);
and UO_390 (O_390,N_19998,N_19955);
and UO_391 (O_391,N_19886,N_19973);
or UO_392 (O_392,N_19754,N_19965);
or UO_393 (O_393,N_19862,N_19982);
or UO_394 (O_394,N_19752,N_19979);
nand UO_395 (O_395,N_19762,N_19802);
nor UO_396 (O_396,N_19824,N_19781);
nor UO_397 (O_397,N_19946,N_19756);
xnor UO_398 (O_398,N_19757,N_19959);
nand UO_399 (O_399,N_19833,N_19817);
or UO_400 (O_400,N_19827,N_19803);
or UO_401 (O_401,N_19879,N_19967);
nand UO_402 (O_402,N_19941,N_19803);
nor UO_403 (O_403,N_19820,N_19998);
nor UO_404 (O_404,N_19831,N_19878);
xnor UO_405 (O_405,N_19887,N_19966);
xor UO_406 (O_406,N_19764,N_19842);
and UO_407 (O_407,N_19878,N_19955);
xnor UO_408 (O_408,N_19942,N_19952);
xor UO_409 (O_409,N_19856,N_19807);
and UO_410 (O_410,N_19963,N_19750);
xnor UO_411 (O_411,N_19908,N_19812);
nand UO_412 (O_412,N_19935,N_19885);
and UO_413 (O_413,N_19962,N_19844);
xnor UO_414 (O_414,N_19759,N_19777);
nand UO_415 (O_415,N_19802,N_19799);
xor UO_416 (O_416,N_19882,N_19890);
or UO_417 (O_417,N_19791,N_19758);
xnor UO_418 (O_418,N_19810,N_19866);
nand UO_419 (O_419,N_19865,N_19831);
xor UO_420 (O_420,N_19995,N_19765);
xor UO_421 (O_421,N_19953,N_19812);
nand UO_422 (O_422,N_19778,N_19805);
nor UO_423 (O_423,N_19909,N_19805);
nor UO_424 (O_424,N_19934,N_19953);
and UO_425 (O_425,N_19799,N_19999);
nor UO_426 (O_426,N_19924,N_19986);
or UO_427 (O_427,N_19936,N_19895);
or UO_428 (O_428,N_19950,N_19793);
nand UO_429 (O_429,N_19755,N_19949);
nand UO_430 (O_430,N_19942,N_19903);
xor UO_431 (O_431,N_19857,N_19852);
or UO_432 (O_432,N_19783,N_19780);
xor UO_433 (O_433,N_19820,N_19858);
and UO_434 (O_434,N_19911,N_19799);
and UO_435 (O_435,N_19887,N_19972);
nor UO_436 (O_436,N_19952,N_19753);
nor UO_437 (O_437,N_19788,N_19907);
or UO_438 (O_438,N_19961,N_19758);
xnor UO_439 (O_439,N_19907,N_19851);
nor UO_440 (O_440,N_19775,N_19988);
xnor UO_441 (O_441,N_19958,N_19861);
xnor UO_442 (O_442,N_19855,N_19961);
nand UO_443 (O_443,N_19760,N_19775);
and UO_444 (O_444,N_19905,N_19948);
xnor UO_445 (O_445,N_19945,N_19815);
or UO_446 (O_446,N_19754,N_19858);
nand UO_447 (O_447,N_19971,N_19821);
or UO_448 (O_448,N_19801,N_19900);
nand UO_449 (O_449,N_19757,N_19913);
nand UO_450 (O_450,N_19784,N_19823);
and UO_451 (O_451,N_19888,N_19930);
xor UO_452 (O_452,N_19964,N_19976);
xor UO_453 (O_453,N_19756,N_19920);
nor UO_454 (O_454,N_19779,N_19801);
or UO_455 (O_455,N_19963,N_19995);
nand UO_456 (O_456,N_19880,N_19793);
nor UO_457 (O_457,N_19925,N_19835);
xnor UO_458 (O_458,N_19884,N_19986);
nor UO_459 (O_459,N_19844,N_19750);
xor UO_460 (O_460,N_19784,N_19902);
nand UO_461 (O_461,N_19853,N_19908);
or UO_462 (O_462,N_19773,N_19846);
xnor UO_463 (O_463,N_19992,N_19960);
xnor UO_464 (O_464,N_19815,N_19785);
or UO_465 (O_465,N_19793,N_19919);
nand UO_466 (O_466,N_19842,N_19933);
nor UO_467 (O_467,N_19950,N_19791);
or UO_468 (O_468,N_19909,N_19957);
nand UO_469 (O_469,N_19867,N_19889);
and UO_470 (O_470,N_19977,N_19933);
or UO_471 (O_471,N_19891,N_19756);
xnor UO_472 (O_472,N_19779,N_19915);
or UO_473 (O_473,N_19784,N_19883);
and UO_474 (O_474,N_19912,N_19838);
nand UO_475 (O_475,N_19879,N_19870);
nand UO_476 (O_476,N_19861,N_19866);
nor UO_477 (O_477,N_19851,N_19965);
or UO_478 (O_478,N_19752,N_19818);
nand UO_479 (O_479,N_19880,N_19832);
nor UO_480 (O_480,N_19935,N_19867);
and UO_481 (O_481,N_19963,N_19870);
or UO_482 (O_482,N_19948,N_19832);
nor UO_483 (O_483,N_19917,N_19923);
and UO_484 (O_484,N_19992,N_19882);
and UO_485 (O_485,N_19763,N_19896);
nand UO_486 (O_486,N_19870,N_19904);
or UO_487 (O_487,N_19880,N_19951);
or UO_488 (O_488,N_19803,N_19933);
and UO_489 (O_489,N_19848,N_19860);
xor UO_490 (O_490,N_19954,N_19758);
nor UO_491 (O_491,N_19815,N_19871);
nand UO_492 (O_492,N_19992,N_19911);
xor UO_493 (O_493,N_19833,N_19872);
nand UO_494 (O_494,N_19773,N_19777);
or UO_495 (O_495,N_19921,N_19757);
or UO_496 (O_496,N_19842,N_19867);
nor UO_497 (O_497,N_19837,N_19895);
nand UO_498 (O_498,N_19901,N_19924);
nor UO_499 (O_499,N_19833,N_19957);
xor UO_500 (O_500,N_19794,N_19899);
or UO_501 (O_501,N_19802,N_19974);
or UO_502 (O_502,N_19800,N_19915);
and UO_503 (O_503,N_19822,N_19982);
xor UO_504 (O_504,N_19884,N_19750);
xnor UO_505 (O_505,N_19754,N_19988);
or UO_506 (O_506,N_19948,N_19954);
xor UO_507 (O_507,N_19922,N_19822);
nand UO_508 (O_508,N_19800,N_19763);
xor UO_509 (O_509,N_19881,N_19856);
and UO_510 (O_510,N_19838,N_19890);
xor UO_511 (O_511,N_19861,N_19908);
xnor UO_512 (O_512,N_19898,N_19815);
nor UO_513 (O_513,N_19810,N_19915);
nor UO_514 (O_514,N_19899,N_19797);
nor UO_515 (O_515,N_19908,N_19975);
nor UO_516 (O_516,N_19958,N_19870);
nor UO_517 (O_517,N_19867,N_19903);
xor UO_518 (O_518,N_19906,N_19874);
xnor UO_519 (O_519,N_19950,N_19973);
and UO_520 (O_520,N_19796,N_19811);
xor UO_521 (O_521,N_19947,N_19843);
xor UO_522 (O_522,N_19889,N_19799);
nand UO_523 (O_523,N_19967,N_19849);
and UO_524 (O_524,N_19862,N_19828);
xnor UO_525 (O_525,N_19908,N_19876);
xnor UO_526 (O_526,N_19964,N_19877);
nor UO_527 (O_527,N_19757,N_19903);
or UO_528 (O_528,N_19765,N_19808);
nand UO_529 (O_529,N_19755,N_19903);
or UO_530 (O_530,N_19843,N_19954);
nor UO_531 (O_531,N_19789,N_19897);
nor UO_532 (O_532,N_19920,N_19854);
nor UO_533 (O_533,N_19853,N_19902);
xor UO_534 (O_534,N_19988,N_19905);
nand UO_535 (O_535,N_19964,N_19842);
and UO_536 (O_536,N_19911,N_19750);
nor UO_537 (O_537,N_19911,N_19956);
or UO_538 (O_538,N_19856,N_19961);
xor UO_539 (O_539,N_19838,N_19937);
xor UO_540 (O_540,N_19782,N_19869);
xor UO_541 (O_541,N_19977,N_19945);
xnor UO_542 (O_542,N_19911,N_19900);
nand UO_543 (O_543,N_19797,N_19978);
and UO_544 (O_544,N_19786,N_19753);
nand UO_545 (O_545,N_19965,N_19992);
nor UO_546 (O_546,N_19861,N_19845);
or UO_547 (O_547,N_19828,N_19957);
and UO_548 (O_548,N_19753,N_19811);
nor UO_549 (O_549,N_19869,N_19990);
nor UO_550 (O_550,N_19803,N_19960);
or UO_551 (O_551,N_19818,N_19777);
and UO_552 (O_552,N_19868,N_19901);
nand UO_553 (O_553,N_19834,N_19775);
nor UO_554 (O_554,N_19988,N_19980);
nand UO_555 (O_555,N_19783,N_19849);
nor UO_556 (O_556,N_19753,N_19931);
or UO_557 (O_557,N_19758,N_19965);
and UO_558 (O_558,N_19858,N_19971);
and UO_559 (O_559,N_19937,N_19763);
and UO_560 (O_560,N_19872,N_19894);
nand UO_561 (O_561,N_19834,N_19909);
and UO_562 (O_562,N_19751,N_19918);
xor UO_563 (O_563,N_19803,N_19901);
nor UO_564 (O_564,N_19750,N_19818);
xor UO_565 (O_565,N_19873,N_19760);
nand UO_566 (O_566,N_19891,N_19912);
and UO_567 (O_567,N_19994,N_19803);
xor UO_568 (O_568,N_19751,N_19910);
xor UO_569 (O_569,N_19897,N_19778);
and UO_570 (O_570,N_19923,N_19853);
nor UO_571 (O_571,N_19789,N_19791);
and UO_572 (O_572,N_19871,N_19799);
or UO_573 (O_573,N_19906,N_19828);
nor UO_574 (O_574,N_19963,N_19760);
nor UO_575 (O_575,N_19781,N_19834);
nand UO_576 (O_576,N_19961,N_19844);
nor UO_577 (O_577,N_19753,N_19885);
or UO_578 (O_578,N_19819,N_19848);
or UO_579 (O_579,N_19967,N_19968);
xor UO_580 (O_580,N_19824,N_19905);
and UO_581 (O_581,N_19863,N_19996);
or UO_582 (O_582,N_19847,N_19759);
nand UO_583 (O_583,N_19932,N_19837);
or UO_584 (O_584,N_19963,N_19811);
xnor UO_585 (O_585,N_19791,N_19891);
and UO_586 (O_586,N_19974,N_19784);
and UO_587 (O_587,N_19837,N_19854);
nand UO_588 (O_588,N_19996,N_19879);
and UO_589 (O_589,N_19897,N_19907);
nor UO_590 (O_590,N_19840,N_19861);
xor UO_591 (O_591,N_19949,N_19955);
nor UO_592 (O_592,N_19760,N_19763);
nor UO_593 (O_593,N_19880,N_19860);
and UO_594 (O_594,N_19839,N_19763);
xnor UO_595 (O_595,N_19779,N_19990);
or UO_596 (O_596,N_19837,N_19910);
or UO_597 (O_597,N_19762,N_19994);
xnor UO_598 (O_598,N_19840,N_19770);
and UO_599 (O_599,N_19805,N_19901);
or UO_600 (O_600,N_19875,N_19796);
or UO_601 (O_601,N_19938,N_19840);
or UO_602 (O_602,N_19945,N_19820);
and UO_603 (O_603,N_19904,N_19763);
xnor UO_604 (O_604,N_19822,N_19818);
or UO_605 (O_605,N_19890,N_19794);
and UO_606 (O_606,N_19843,N_19879);
nand UO_607 (O_607,N_19856,N_19995);
or UO_608 (O_608,N_19785,N_19845);
nor UO_609 (O_609,N_19874,N_19904);
nand UO_610 (O_610,N_19858,N_19976);
nand UO_611 (O_611,N_19766,N_19948);
or UO_612 (O_612,N_19987,N_19891);
xnor UO_613 (O_613,N_19963,N_19998);
nor UO_614 (O_614,N_19812,N_19931);
xnor UO_615 (O_615,N_19803,N_19843);
or UO_616 (O_616,N_19793,N_19792);
nor UO_617 (O_617,N_19866,N_19788);
nor UO_618 (O_618,N_19903,N_19946);
nor UO_619 (O_619,N_19880,N_19873);
and UO_620 (O_620,N_19834,N_19794);
nand UO_621 (O_621,N_19973,N_19890);
nand UO_622 (O_622,N_19951,N_19892);
and UO_623 (O_623,N_19918,N_19975);
or UO_624 (O_624,N_19897,N_19835);
or UO_625 (O_625,N_19868,N_19857);
nor UO_626 (O_626,N_19824,N_19907);
nor UO_627 (O_627,N_19796,N_19842);
and UO_628 (O_628,N_19824,N_19903);
or UO_629 (O_629,N_19874,N_19829);
nor UO_630 (O_630,N_19802,N_19758);
or UO_631 (O_631,N_19985,N_19832);
nand UO_632 (O_632,N_19978,N_19816);
and UO_633 (O_633,N_19860,N_19758);
or UO_634 (O_634,N_19762,N_19806);
xnor UO_635 (O_635,N_19815,N_19839);
xnor UO_636 (O_636,N_19997,N_19778);
xor UO_637 (O_637,N_19922,N_19878);
or UO_638 (O_638,N_19776,N_19920);
nor UO_639 (O_639,N_19992,N_19849);
or UO_640 (O_640,N_19793,N_19871);
xor UO_641 (O_641,N_19789,N_19861);
and UO_642 (O_642,N_19931,N_19752);
nand UO_643 (O_643,N_19941,N_19783);
or UO_644 (O_644,N_19822,N_19803);
nor UO_645 (O_645,N_19853,N_19788);
nor UO_646 (O_646,N_19972,N_19796);
and UO_647 (O_647,N_19862,N_19771);
nor UO_648 (O_648,N_19878,N_19852);
and UO_649 (O_649,N_19926,N_19848);
xnor UO_650 (O_650,N_19858,N_19948);
or UO_651 (O_651,N_19935,N_19907);
or UO_652 (O_652,N_19975,N_19790);
nor UO_653 (O_653,N_19992,N_19936);
xor UO_654 (O_654,N_19800,N_19773);
and UO_655 (O_655,N_19907,N_19769);
nor UO_656 (O_656,N_19788,N_19909);
nor UO_657 (O_657,N_19950,N_19801);
and UO_658 (O_658,N_19759,N_19774);
nor UO_659 (O_659,N_19808,N_19801);
or UO_660 (O_660,N_19973,N_19979);
nor UO_661 (O_661,N_19777,N_19793);
nor UO_662 (O_662,N_19976,N_19981);
nand UO_663 (O_663,N_19796,N_19979);
nor UO_664 (O_664,N_19911,N_19896);
or UO_665 (O_665,N_19848,N_19965);
xnor UO_666 (O_666,N_19807,N_19918);
or UO_667 (O_667,N_19811,N_19916);
or UO_668 (O_668,N_19759,N_19816);
nand UO_669 (O_669,N_19874,N_19868);
xor UO_670 (O_670,N_19782,N_19816);
and UO_671 (O_671,N_19834,N_19823);
nand UO_672 (O_672,N_19753,N_19967);
and UO_673 (O_673,N_19823,N_19765);
nand UO_674 (O_674,N_19767,N_19897);
and UO_675 (O_675,N_19813,N_19792);
and UO_676 (O_676,N_19830,N_19803);
nor UO_677 (O_677,N_19940,N_19760);
nand UO_678 (O_678,N_19772,N_19794);
or UO_679 (O_679,N_19991,N_19845);
nand UO_680 (O_680,N_19955,N_19846);
or UO_681 (O_681,N_19773,N_19999);
xor UO_682 (O_682,N_19888,N_19957);
nand UO_683 (O_683,N_19770,N_19777);
xnor UO_684 (O_684,N_19790,N_19942);
nor UO_685 (O_685,N_19999,N_19932);
xor UO_686 (O_686,N_19931,N_19910);
or UO_687 (O_687,N_19986,N_19885);
nor UO_688 (O_688,N_19999,N_19910);
and UO_689 (O_689,N_19784,N_19773);
nand UO_690 (O_690,N_19807,N_19848);
nand UO_691 (O_691,N_19946,N_19920);
nand UO_692 (O_692,N_19911,N_19810);
nand UO_693 (O_693,N_19959,N_19804);
or UO_694 (O_694,N_19929,N_19791);
and UO_695 (O_695,N_19778,N_19926);
xnor UO_696 (O_696,N_19814,N_19936);
xnor UO_697 (O_697,N_19907,N_19944);
nor UO_698 (O_698,N_19755,N_19918);
nor UO_699 (O_699,N_19933,N_19864);
and UO_700 (O_700,N_19935,N_19948);
nor UO_701 (O_701,N_19895,N_19994);
or UO_702 (O_702,N_19762,N_19846);
nand UO_703 (O_703,N_19928,N_19785);
or UO_704 (O_704,N_19761,N_19921);
and UO_705 (O_705,N_19786,N_19781);
nand UO_706 (O_706,N_19808,N_19752);
xor UO_707 (O_707,N_19788,N_19944);
nand UO_708 (O_708,N_19801,N_19836);
or UO_709 (O_709,N_19808,N_19958);
nor UO_710 (O_710,N_19761,N_19829);
or UO_711 (O_711,N_19868,N_19927);
and UO_712 (O_712,N_19786,N_19761);
nand UO_713 (O_713,N_19820,N_19905);
xor UO_714 (O_714,N_19804,N_19929);
or UO_715 (O_715,N_19870,N_19869);
nand UO_716 (O_716,N_19769,N_19877);
and UO_717 (O_717,N_19913,N_19836);
and UO_718 (O_718,N_19996,N_19777);
xor UO_719 (O_719,N_19791,N_19827);
xnor UO_720 (O_720,N_19918,N_19815);
nand UO_721 (O_721,N_19788,N_19847);
nand UO_722 (O_722,N_19906,N_19802);
xor UO_723 (O_723,N_19844,N_19786);
xnor UO_724 (O_724,N_19750,N_19905);
and UO_725 (O_725,N_19958,N_19844);
nor UO_726 (O_726,N_19762,N_19777);
or UO_727 (O_727,N_19795,N_19829);
or UO_728 (O_728,N_19885,N_19852);
or UO_729 (O_729,N_19984,N_19998);
nor UO_730 (O_730,N_19972,N_19831);
nand UO_731 (O_731,N_19750,N_19842);
nor UO_732 (O_732,N_19924,N_19759);
or UO_733 (O_733,N_19787,N_19877);
xor UO_734 (O_734,N_19992,N_19788);
nand UO_735 (O_735,N_19759,N_19807);
and UO_736 (O_736,N_19968,N_19797);
nand UO_737 (O_737,N_19839,N_19860);
and UO_738 (O_738,N_19930,N_19989);
xor UO_739 (O_739,N_19965,N_19864);
nand UO_740 (O_740,N_19836,N_19909);
or UO_741 (O_741,N_19834,N_19761);
xnor UO_742 (O_742,N_19770,N_19847);
and UO_743 (O_743,N_19866,N_19939);
nor UO_744 (O_744,N_19806,N_19751);
nand UO_745 (O_745,N_19988,N_19976);
and UO_746 (O_746,N_19841,N_19809);
xnor UO_747 (O_747,N_19999,N_19985);
nor UO_748 (O_748,N_19910,N_19834);
and UO_749 (O_749,N_19843,N_19995);
xor UO_750 (O_750,N_19958,N_19887);
nand UO_751 (O_751,N_19814,N_19798);
nand UO_752 (O_752,N_19790,N_19761);
and UO_753 (O_753,N_19890,N_19809);
or UO_754 (O_754,N_19930,N_19935);
and UO_755 (O_755,N_19808,N_19753);
xor UO_756 (O_756,N_19761,N_19832);
nor UO_757 (O_757,N_19914,N_19913);
xor UO_758 (O_758,N_19806,N_19876);
xor UO_759 (O_759,N_19761,N_19964);
and UO_760 (O_760,N_19908,N_19756);
nor UO_761 (O_761,N_19888,N_19764);
xnor UO_762 (O_762,N_19823,N_19788);
nand UO_763 (O_763,N_19905,N_19815);
xnor UO_764 (O_764,N_19946,N_19930);
and UO_765 (O_765,N_19875,N_19838);
xor UO_766 (O_766,N_19915,N_19928);
or UO_767 (O_767,N_19909,N_19895);
and UO_768 (O_768,N_19905,N_19957);
nor UO_769 (O_769,N_19940,N_19870);
and UO_770 (O_770,N_19893,N_19988);
nand UO_771 (O_771,N_19909,N_19760);
and UO_772 (O_772,N_19997,N_19948);
nor UO_773 (O_773,N_19785,N_19876);
xor UO_774 (O_774,N_19775,N_19800);
or UO_775 (O_775,N_19897,N_19888);
and UO_776 (O_776,N_19967,N_19756);
nor UO_777 (O_777,N_19779,N_19982);
and UO_778 (O_778,N_19920,N_19926);
nor UO_779 (O_779,N_19755,N_19772);
nor UO_780 (O_780,N_19999,N_19768);
or UO_781 (O_781,N_19924,N_19859);
and UO_782 (O_782,N_19828,N_19970);
nor UO_783 (O_783,N_19946,N_19884);
nand UO_784 (O_784,N_19813,N_19777);
nor UO_785 (O_785,N_19911,N_19855);
xor UO_786 (O_786,N_19905,N_19829);
nand UO_787 (O_787,N_19997,N_19842);
nand UO_788 (O_788,N_19948,N_19907);
and UO_789 (O_789,N_19856,N_19903);
or UO_790 (O_790,N_19987,N_19864);
or UO_791 (O_791,N_19799,N_19758);
xnor UO_792 (O_792,N_19994,N_19919);
nor UO_793 (O_793,N_19850,N_19785);
and UO_794 (O_794,N_19853,N_19832);
and UO_795 (O_795,N_19887,N_19875);
and UO_796 (O_796,N_19766,N_19782);
nor UO_797 (O_797,N_19857,N_19903);
nor UO_798 (O_798,N_19870,N_19821);
nand UO_799 (O_799,N_19789,N_19878);
and UO_800 (O_800,N_19806,N_19988);
nor UO_801 (O_801,N_19793,N_19807);
nor UO_802 (O_802,N_19828,N_19798);
or UO_803 (O_803,N_19961,N_19990);
or UO_804 (O_804,N_19787,N_19938);
xor UO_805 (O_805,N_19768,N_19890);
xor UO_806 (O_806,N_19932,N_19765);
and UO_807 (O_807,N_19972,N_19930);
or UO_808 (O_808,N_19780,N_19815);
or UO_809 (O_809,N_19797,N_19783);
nand UO_810 (O_810,N_19983,N_19768);
xnor UO_811 (O_811,N_19911,N_19932);
nand UO_812 (O_812,N_19985,N_19772);
or UO_813 (O_813,N_19821,N_19799);
nand UO_814 (O_814,N_19877,N_19846);
nor UO_815 (O_815,N_19983,N_19782);
nand UO_816 (O_816,N_19956,N_19903);
or UO_817 (O_817,N_19759,N_19884);
nand UO_818 (O_818,N_19912,N_19956);
nor UO_819 (O_819,N_19866,N_19800);
nor UO_820 (O_820,N_19772,N_19859);
and UO_821 (O_821,N_19874,N_19900);
or UO_822 (O_822,N_19833,N_19945);
or UO_823 (O_823,N_19981,N_19808);
and UO_824 (O_824,N_19899,N_19755);
nor UO_825 (O_825,N_19972,N_19836);
and UO_826 (O_826,N_19944,N_19904);
and UO_827 (O_827,N_19928,N_19842);
and UO_828 (O_828,N_19899,N_19866);
and UO_829 (O_829,N_19903,N_19969);
xor UO_830 (O_830,N_19921,N_19811);
or UO_831 (O_831,N_19759,N_19839);
nor UO_832 (O_832,N_19914,N_19937);
nor UO_833 (O_833,N_19927,N_19993);
xor UO_834 (O_834,N_19906,N_19799);
and UO_835 (O_835,N_19892,N_19913);
or UO_836 (O_836,N_19958,N_19975);
nand UO_837 (O_837,N_19805,N_19904);
or UO_838 (O_838,N_19867,N_19884);
and UO_839 (O_839,N_19923,N_19931);
nand UO_840 (O_840,N_19898,N_19847);
nor UO_841 (O_841,N_19943,N_19882);
xor UO_842 (O_842,N_19967,N_19982);
nor UO_843 (O_843,N_19861,N_19941);
and UO_844 (O_844,N_19816,N_19965);
xor UO_845 (O_845,N_19918,N_19796);
or UO_846 (O_846,N_19963,N_19810);
nand UO_847 (O_847,N_19925,N_19778);
or UO_848 (O_848,N_19849,N_19872);
nor UO_849 (O_849,N_19803,N_19982);
or UO_850 (O_850,N_19819,N_19856);
nor UO_851 (O_851,N_19841,N_19963);
xor UO_852 (O_852,N_19943,N_19774);
nand UO_853 (O_853,N_19840,N_19871);
nand UO_854 (O_854,N_19766,N_19905);
xnor UO_855 (O_855,N_19932,N_19899);
nand UO_856 (O_856,N_19801,N_19854);
nor UO_857 (O_857,N_19820,N_19809);
or UO_858 (O_858,N_19828,N_19938);
or UO_859 (O_859,N_19807,N_19832);
and UO_860 (O_860,N_19942,N_19954);
and UO_861 (O_861,N_19966,N_19931);
and UO_862 (O_862,N_19824,N_19778);
xnor UO_863 (O_863,N_19826,N_19781);
and UO_864 (O_864,N_19948,N_19827);
nor UO_865 (O_865,N_19880,N_19899);
or UO_866 (O_866,N_19885,N_19859);
or UO_867 (O_867,N_19917,N_19856);
xnor UO_868 (O_868,N_19801,N_19769);
or UO_869 (O_869,N_19932,N_19789);
and UO_870 (O_870,N_19957,N_19895);
xor UO_871 (O_871,N_19830,N_19799);
nand UO_872 (O_872,N_19988,N_19823);
nor UO_873 (O_873,N_19844,N_19983);
xnor UO_874 (O_874,N_19987,N_19801);
and UO_875 (O_875,N_19976,N_19972);
nand UO_876 (O_876,N_19860,N_19941);
or UO_877 (O_877,N_19839,N_19938);
and UO_878 (O_878,N_19911,N_19864);
xor UO_879 (O_879,N_19779,N_19957);
nor UO_880 (O_880,N_19977,N_19880);
and UO_881 (O_881,N_19902,N_19844);
nand UO_882 (O_882,N_19919,N_19843);
xor UO_883 (O_883,N_19812,N_19798);
xor UO_884 (O_884,N_19852,N_19880);
xor UO_885 (O_885,N_19875,N_19917);
xor UO_886 (O_886,N_19951,N_19955);
nand UO_887 (O_887,N_19951,N_19817);
or UO_888 (O_888,N_19960,N_19818);
or UO_889 (O_889,N_19963,N_19868);
nand UO_890 (O_890,N_19827,N_19883);
or UO_891 (O_891,N_19994,N_19836);
and UO_892 (O_892,N_19798,N_19973);
nand UO_893 (O_893,N_19838,N_19819);
nand UO_894 (O_894,N_19767,N_19848);
or UO_895 (O_895,N_19756,N_19867);
or UO_896 (O_896,N_19874,N_19757);
or UO_897 (O_897,N_19928,N_19913);
nand UO_898 (O_898,N_19845,N_19990);
xor UO_899 (O_899,N_19765,N_19901);
xor UO_900 (O_900,N_19866,N_19864);
and UO_901 (O_901,N_19998,N_19980);
xor UO_902 (O_902,N_19758,N_19968);
or UO_903 (O_903,N_19898,N_19887);
nor UO_904 (O_904,N_19797,N_19888);
nor UO_905 (O_905,N_19899,N_19893);
xnor UO_906 (O_906,N_19767,N_19915);
nor UO_907 (O_907,N_19801,N_19766);
xor UO_908 (O_908,N_19902,N_19815);
and UO_909 (O_909,N_19858,N_19999);
or UO_910 (O_910,N_19857,N_19756);
xnor UO_911 (O_911,N_19953,N_19836);
nor UO_912 (O_912,N_19865,N_19814);
and UO_913 (O_913,N_19877,N_19882);
nor UO_914 (O_914,N_19969,N_19905);
xor UO_915 (O_915,N_19814,N_19902);
or UO_916 (O_916,N_19760,N_19998);
xnor UO_917 (O_917,N_19936,N_19952);
and UO_918 (O_918,N_19836,N_19820);
nand UO_919 (O_919,N_19882,N_19970);
or UO_920 (O_920,N_19776,N_19780);
nand UO_921 (O_921,N_19968,N_19906);
nor UO_922 (O_922,N_19941,N_19864);
nand UO_923 (O_923,N_19895,N_19810);
and UO_924 (O_924,N_19850,N_19826);
nor UO_925 (O_925,N_19852,N_19993);
or UO_926 (O_926,N_19770,N_19812);
or UO_927 (O_927,N_19864,N_19908);
nand UO_928 (O_928,N_19774,N_19758);
xnor UO_929 (O_929,N_19960,N_19842);
and UO_930 (O_930,N_19765,N_19918);
and UO_931 (O_931,N_19992,N_19974);
xnor UO_932 (O_932,N_19995,N_19897);
or UO_933 (O_933,N_19829,N_19907);
nand UO_934 (O_934,N_19773,N_19805);
nor UO_935 (O_935,N_19774,N_19999);
nor UO_936 (O_936,N_19999,N_19941);
nor UO_937 (O_937,N_19918,N_19759);
nand UO_938 (O_938,N_19890,N_19845);
xnor UO_939 (O_939,N_19869,N_19957);
and UO_940 (O_940,N_19905,N_19813);
nand UO_941 (O_941,N_19770,N_19854);
nor UO_942 (O_942,N_19947,N_19959);
nor UO_943 (O_943,N_19856,N_19933);
xnor UO_944 (O_944,N_19804,N_19943);
nor UO_945 (O_945,N_19852,N_19814);
nor UO_946 (O_946,N_19830,N_19787);
nand UO_947 (O_947,N_19823,N_19826);
or UO_948 (O_948,N_19755,N_19808);
and UO_949 (O_949,N_19972,N_19859);
or UO_950 (O_950,N_19802,N_19755);
or UO_951 (O_951,N_19938,N_19958);
and UO_952 (O_952,N_19842,N_19853);
or UO_953 (O_953,N_19828,N_19787);
xor UO_954 (O_954,N_19878,N_19851);
xnor UO_955 (O_955,N_19769,N_19980);
or UO_956 (O_956,N_19935,N_19931);
or UO_957 (O_957,N_19841,N_19965);
xnor UO_958 (O_958,N_19981,N_19822);
and UO_959 (O_959,N_19776,N_19834);
xor UO_960 (O_960,N_19782,N_19878);
nand UO_961 (O_961,N_19775,N_19767);
or UO_962 (O_962,N_19904,N_19811);
or UO_963 (O_963,N_19823,N_19807);
nor UO_964 (O_964,N_19876,N_19938);
and UO_965 (O_965,N_19763,N_19993);
xnor UO_966 (O_966,N_19979,N_19961);
nor UO_967 (O_967,N_19785,N_19906);
xor UO_968 (O_968,N_19929,N_19803);
nand UO_969 (O_969,N_19829,N_19759);
nor UO_970 (O_970,N_19941,N_19862);
nand UO_971 (O_971,N_19797,N_19918);
nor UO_972 (O_972,N_19781,N_19750);
nand UO_973 (O_973,N_19978,N_19859);
nor UO_974 (O_974,N_19950,N_19889);
xnor UO_975 (O_975,N_19775,N_19900);
xor UO_976 (O_976,N_19769,N_19818);
or UO_977 (O_977,N_19933,N_19774);
xor UO_978 (O_978,N_19793,N_19971);
nand UO_979 (O_979,N_19889,N_19966);
nand UO_980 (O_980,N_19818,N_19778);
nand UO_981 (O_981,N_19951,N_19833);
and UO_982 (O_982,N_19762,N_19784);
nor UO_983 (O_983,N_19767,N_19942);
nor UO_984 (O_984,N_19826,N_19928);
or UO_985 (O_985,N_19845,N_19897);
nand UO_986 (O_986,N_19780,N_19831);
and UO_987 (O_987,N_19994,N_19798);
or UO_988 (O_988,N_19843,N_19834);
nor UO_989 (O_989,N_19800,N_19794);
and UO_990 (O_990,N_19758,N_19854);
nand UO_991 (O_991,N_19952,N_19888);
or UO_992 (O_992,N_19792,N_19853);
nor UO_993 (O_993,N_19882,N_19962);
xnor UO_994 (O_994,N_19850,N_19972);
nor UO_995 (O_995,N_19859,N_19755);
and UO_996 (O_996,N_19953,N_19804);
or UO_997 (O_997,N_19906,N_19992);
nand UO_998 (O_998,N_19877,N_19835);
nand UO_999 (O_999,N_19811,N_19846);
or UO_1000 (O_1000,N_19814,N_19855);
or UO_1001 (O_1001,N_19788,N_19981);
and UO_1002 (O_1002,N_19897,N_19961);
and UO_1003 (O_1003,N_19922,N_19912);
nor UO_1004 (O_1004,N_19914,N_19843);
nand UO_1005 (O_1005,N_19815,N_19928);
or UO_1006 (O_1006,N_19803,N_19842);
xnor UO_1007 (O_1007,N_19973,N_19894);
nor UO_1008 (O_1008,N_19750,N_19766);
or UO_1009 (O_1009,N_19824,N_19750);
nor UO_1010 (O_1010,N_19874,N_19957);
xnor UO_1011 (O_1011,N_19804,N_19842);
nor UO_1012 (O_1012,N_19792,N_19872);
or UO_1013 (O_1013,N_19788,N_19868);
and UO_1014 (O_1014,N_19997,N_19785);
or UO_1015 (O_1015,N_19867,N_19910);
nand UO_1016 (O_1016,N_19814,N_19773);
nor UO_1017 (O_1017,N_19764,N_19968);
xor UO_1018 (O_1018,N_19758,N_19857);
nand UO_1019 (O_1019,N_19878,N_19905);
and UO_1020 (O_1020,N_19762,N_19801);
nand UO_1021 (O_1021,N_19858,N_19771);
and UO_1022 (O_1022,N_19826,N_19900);
or UO_1023 (O_1023,N_19817,N_19792);
xor UO_1024 (O_1024,N_19995,N_19880);
and UO_1025 (O_1025,N_19846,N_19979);
or UO_1026 (O_1026,N_19971,N_19799);
xor UO_1027 (O_1027,N_19783,N_19860);
nand UO_1028 (O_1028,N_19876,N_19863);
and UO_1029 (O_1029,N_19805,N_19975);
xnor UO_1030 (O_1030,N_19989,N_19755);
nand UO_1031 (O_1031,N_19848,N_19811);
or UO_1032 (O_1032,N_19987,N_19890);
nor UO_1033 (O_1033,N_19801,N_19806);
and UO_1034 (O_1034,N_19853,N_19833);
or UO_1035 (O_1035,N_19761,N_19876);
xor UO_1036 (O_1036,N_19915,N_19870);
and UO_1037 (O_1037,N_19752,N_19924);
xnor UO_1038 (O_1038,N_19805,N_19823);
xor UO_1039 (O_1039,N_19804,N_19807);
and UO_1040 (O_1040,N_19842,N_19789);
nor UO_1041 (O_1041,N_19880,N_19945);
nor UO_1042 (O_1042,N_19940,N_19980);
xor UO_1043 (O_1043,N_19991,N_19799);
nand UO_1044 (O_1044,N_19966,N_19809);
xnor UO_1045 (O_1045,N_19761,N_19849);
nand UO_1046 (O_1046,N_19824,N_19819);
xor UO_1047 (O_1047,N_19912,N_19831);
nor UO_1048 (O_1048,N_19906,N_19798);
or UO_1049 (O_1049,N_19904,N_19817);
and UO_1050 (O_1050,N_19768,N_19781);
nor UO_1051 (O_1051,N_19845,N_19790);
nand UO_1052 (O_1052,N_19974,N_19983);
nand UO_1053 (O_1053,N_19948,N_19786);
nor UO_1054 (O_1054,N_19988,N_19834);
or UO_1055 (O_1055,N_19758,N_19951);
or UO_1056 (O_1056,N_19882,N_19888);
nor UO_1057 (O_1057,N_19820,N_19996);
or UO_1058 (O_1058,N_19953,N_19995);
nor UO_1059 (O_1059,N_19944,N_19982);
or UO_1060 (O_1060,N_19897,N_19973);
nor UO_1061 (O_1061,N_19768,N_19889);
nand UO_1062 (O_1062,N_19874,N_19837);
or UO_1063 (O_1063,N_19801,N_19800);
or UO_1064 (O_1064,N_19822,N_19942);
nand UO_1065 (O_1065,N_19956,N_19910);
and UO_1066 (O_1066,N_19837,N_19790);
nand UO_1067 (O_1067,N_19995,N_19980);
nor UO_1068 (O_1068,N_19756,N_19878);
nor UO_1069 (O_1069,N_19802,N_19995);
xnor UO_1070 (O_1070,N_19890,N_19821);
xnor UO_1071 (O_1071,N_19847,N_19872);
and UO_1072 (O_1072,N_19774,N_19983);
nand UO_1073 (O_1073,N_19808,N_19966);
xor UO_1074 (O_1074,N_19794,N_19948);
or UO_1075 (O_1075,N_19824,N_19942);
nand UO_1076 (O_1076,N_19840,N_19964);
or UO_1077 (O_1077,N_19794,N_19985);
nand UO_1078 (O_1078,N_19997,N_19975);
nand UO_1079 (O_1079,N_19984,N_19925);
and UO_1080 (O_1080,N_19967,N_19865);
xor UO_1081 (O_1081,N_19753,N_19762);
nand UO_1082 (O_1082,N_19763,N_19921);
nor UO_1083 (O_1083,N_19804,N_19859);
nor UO_1084 (O_1084,N_19974,N_19986);
xnor UO_1085 (O_1085,N_19905,N_19828);
and UO_1086 (O_1086,N_19779,N_19987);
or UO_1087 (O_1087,N_19937,N_19768);
nand UO_1088 (O_1088,N_19982,N_19853);
xnor UO_1089 (O_1089,N_19837,N_19870);
nor UO_1090 (O_1090,N_19896,N_19862);
or UO_1091 (O_1091,N_19871,N_19830);
nor UO_1092 (O_1092,N_19944,N_19918);
nand UO_1093 (O_1093,N_19992,N_19880);
or UO_1094 (O_1094,N_19945,N_19917);
nor UO_1095 (O_1095,N_19832,N_19932);
or UO_1096 (O_1096,N_19921,N_19807);
nor UO_1097 (O_1097,N_19890,N_19861);
nand UO_1098 (O_1098,N_19991,N_19864);
and UO_1099 (O_1099,N_19758,N_19956);
nor UO_1100 (O_1100,N_19950,N_19774);
nor UO_1101 (O_1101,N_19810,N_19868);
xor UO_1102 (O_1102,N_19863,N_19957);
nor UO_1103 (O_1103,N_19756,N_19970);
or UO_1104 (O_1104,N_19977,N_19868);
nor UO_1105 (O_1105,N_19832,N_19916);
or UO_1106 (O_1106,N_19977,N_19985);
or UO_1107 (O_1107,N_19989,N_19962);
xor UO_1108 (O_1108,N_19765,N_19756);
or UO_1109 (O_1109,N_19850,N_19792);
xor UO_1110 (O_1110,N_19834,N_19904);
xor UO_1111 (O_1111,N_19778,N_19767);
nand UO_1112 (O_1112,N_19893,N_19968);
nor UO_1113 (O_1113,N_19957,N_19971);
xor UO_1114 (O_1114,N_19945,N_19854);
xor UO_1115 (O_1115,N_19813,N_19850);
and UO_1116 (O_1116,N_19756,N_19783);
nor UO_1117 (O_1117,N_19895,N_19814);
and UO_1118 (O_1118,N_19894,N_19839);
and UO_1119 (O_1119,N_19888,N_19836);
and UO_1120 (O_1120,N_19902,N_19850);
xor UO_1121 (O_1121,N_19927,N_19846);
or UO_1122 (O_1122,N_19909,N_19999);
nor UO_1123 (O_1123,N_19848,N_19934);
and UO_1124 (O_1124,N_19955,N_19896);
xor UO_1125 (O_1125,N_19978,N_19980);
nor UO_1126 (O_1126,N_19915,N_19764);
nand UO_1127 (O_1127,N_19906,N_19854);
xor UO_1128 (O_1128,N_19846,N_19894);
xor UO_1129 (O_1129,N_19766,N_19936);
or UO_1130 (O_1130,N_19991,N_19831);
nand UO_1131 (O_1131,N_19847,N_19948);
nand UO_1132 (O_1132,N_19913,N_19941);
and UO_1133 (O_1133,N_19910,N_19784);
or UO_1134 (O_1134,N_19780,N_19887);
xnor UO_1135 (O_1135,N_19852,N_19764);
xnor UO_1136 (O_1136,N_19757,N_19915);
nor UO_1137 (O_1137,N_19878,N_19817);
and UO_1138 (O_1138,N_19806,N_19802);
nand UO_1139 (O_1139,N_19768,N_19987);
xnor UO_1140 (O_1140,N_19785,N_19977);
nor UO_1141 (O_1141,N_19770,N_19853);
nand UO_1142 (O_1142,N_19769,N_19967);
and UO_1143 (O_1143,N_19928,N_19786);
nand UO_1144 (O_1144,N_19768,N_19831);
xnor UO_1145 (O_1145,N_19964,N_19817);
nor UO_1146 (O_1146,N_19810,N_19799);
and UO_1147 (O_1147,N_19889,N_19872);
nand UO_1148 (O_1148,N_19762,N_19837);
xnor UO_1149 (O_1149,N_19983,N_19921);
nand UO_1150 (O_1150,N_19888,N_19999);
nor UO_1151 (O_1151,N_19795,N_19868);
or UO_1152 (O_1152,N_19828,N_19949);
and UO_1153 (O_1153,N_19858,N_19919);
or UO_1154 (O_1154,N_19997,N_19924);
or UO_1155 (O_1155,N_19861,N_19947);
and UO_1156 (O_1156,N_19999,N_19889);
or UO_1157 (O_1157,N_19751,N_19972);
or UO_1158 (O_1158,N_19916,N_19780);
xor UO_1159 (O_1159,N_19771,N_19860);
xor UO_1160 (O_1160,N_19830,N_19991);
nand UO_1161 (O_1161,N_19804,N_19894);
xor UO_1162 (O_1162,N_19962,N_19772);
xor UO_1163 (O_1163,N_19883,N_19841);
nor UO_1164 (O_1164,N_19870,N_19913);
and UO_1165 (O_1165,N_19950,N_19902);
nand UO_1166 (O_1166,N_19765,N_19977);
nand UO_1167 (O_1167,N_19956,N_19905);
nor UO_1168 (O_1168,N_19841,N_19953);
nand UO_1169 (O_1169,N_19873,N_19776);
or UO_1170 (O_1170,N_19909,N_19936);
nor UO_1171 (O_1171,N_19902,N_19886);
nand UO_1172 (O_1172,N_19821,N_19928);
nand UO_1173 (O_1173,N_19956,N_19863);
and UO_1174 (O_1174,N_19985,N_19814);
nor UO_1175 (O_1175,N_19899,N_19847);
nand UO_1176 (O_1176,N_19979,N_19760);
or UO_1177 (O_1177,N_19866,N_19882);
and UO_1178 (O_1178,N_19765,N_19875);
xor UO_1179 (O_1179,N_19850,N_19896);
nand UO_1180 (O_1180,N_19771,N_19944);
nor UO_1181 (O_1181,N_19978,N_19780);
or UO_1182 (O_1182,N_19892,N_19814);
and UO_1183 (O_1183,N_19964,N_19865);
nor UO_1184 (O_1184,N_19787,N_19879);
and UO_1185 (O_1185,N_19809,N_19865);
or UO_1186 (O_1186,N_19939,N_19892);
and UO_1187 (O_1187,N_19937,N_19930);
xnor UO_1188 (O_1188,N_19985,N_19820);
nor UO_1189 (O_1189,N_19804,N_19770);
nor UO_1190 (O_1190,N_19759,N_19830);
nand UO_1191 (O_1191,N_19876,N_19917);
nor UO_1192 (O_1192,N_19786,N_19861);
xor UO_1193 (O_1193,N_19979,N_19887);
nor UO_1194 (O_1194,N_19818,N_19992);
xnor UO_1195 (O_1195,N_19773,N_19929);
nand UO_1196 (O_1196,N_19874,N_19788);
nand UO_1197 (O_1197,N_19942,N_19909);
nor UO_1198 (O_1198,N_19972,N_19906);
or UO_1199 (O_1199,N_19900,N_19945);
or UO_1200 (O_1200,N_19782,N_19880);
nand UO_1201 (O_1201,N_19910,N_19853);
or UO_1202 (O_1202,N_19951,N_19752);
nor UO_1203 (O_1203,N_19905,N_19909);
nand UO_1204 (O_1204,N_19903,N_19973);
and UO_1205 (O_1205,N_19940,N_19987);
and UO_1206 (O_1206,N_19751,N_19857);
or UO_1207 (O_1207,N_19935,N_19839);
xor UO_1208 (O_1208,N_19842,N_19994);
or UO_1209 (O_1209,N_19913,N_19866);
or UO_1210 (O_1210,N_19763,N_19810);
xnor UO_1211 (O_1211,N_19945,N_19912);
nand UO_1212 (O_1212,N_19961,N_19918);
xor UO_1213 (O_1213,N_19826,N_19873);
xor UO_1214 (O_1214,N_19899,N_19971);
xnor UO_1215 (O_1215,N_19752,N_19764);
and UO_1216 (O_1216,N_19860,N_19967);
nor UO_1217 (O_1217,N_19931,N_19954);
nor UO_1218 (O_1218,N_19802,N_19937);
xor UO_1219 (O_1219,N_19995,N_19926);
nand UO_1220 (O_1220,N_19805,N_19781);
or UO_1221 (O_1221,N_19980,N_19839);
nand UO_1222 (O_1222,N_19803,N_19835);
nor UO_1223 (O_1223,N_19961,N_19783);
xnor UO_1224 (O_1224,N_19750,N_19762);
or UO_1225 (O_1225,N_19946,N_19784);
and UO_1226 (O_1226,N_19834,N_19873);
nand UO_1227 (O_1227,N_19936,N_19801);
or UO_1228 (O_1228,N_19768,N_19860);
and UO_1229 (O_1229,N_19863,N_19763);
xnor UO_1230 (O_1230,N_19929,N_19762);
nand UO_1231 (O_1231,N_19874,N_19847);
or UO_1232 (O_1232,N_19807,N_19999);
xnor UO_1233 (O_1233,N_19848,N_19945);
nor UO_1234 (O_1234,N_19943,N_19766);
xor UO_1235 (O_1235,N_19893,N_19793);
nor UO_1236 (O_1236,N_19877,N_19775);
or UO_1237 (O_1237,N_19945,N_19762);
or UO_1238 (O_1238,N_19770,N_19998);
or UO_1239 (O_1239,N_19751,N_19912);
nand UO_1240 (O_1240,N_19970,N_19944);
nand UO_1241 (O_1241,N_19931,N_19995);
xnor UO_1242 (O_1242,N_19829,N_19967);
nand UO_1243 (O_1243,N_19750,N_19786);
or UO_1244 (O_1244,N_19998,N_19911);
nand UO_1245 (O_1245,N_19883,N_19856);
xnor UO_1246 (O_1246,N_19862,N_19790);
and UO_1247 (O_1247,N_19921,N_19971);
nor UO_1248 (O_1248,N_19889,N_19942);
or UO_1249 (O_1249,N_19819,N_19882);
and UO_1250 (O_1250,N_19861,N_19939);
nor UO_1251 (O_1251,N_19789,N_19778);
nand UO_1252 (O_1252,N_19990,N_19757);
nand UO_1253 (O_1253,N_19814,N_19917);
or UO_1254 (O_1254,N_19952,N_19786);
nor UO_1255 (O_1255,N_19940,N_19932);
nand UO_1256 (O_1256,N_19931,N_19852);
and UO_1257 (O_1257,N_19915,N_19960);
nand UO_1258 (O_1258,N_19926,N_19787);
nand UO_1259 (O_1259,N_19777,N_19949);
or UO_1260 (O_1260,N_19811,N_19948);
or UO_1261 (O_1261,N_19903,N_19802);
or UO_1262 (O_1262,N_19869,N_19905);
or UO_1263 (O_1263,N_19820,N_19894);
or UO_1264 (O_1264,N_19846,N_19839);
and UO_1265 (O_1265,N_19830,N_19939);
nand UO_1266 (O_1266,N_19966,N_19857);
xor UO_1267 (O_1267,N_19833,N_19933);
nor UO_1268 (O_1268,N_19916,N_19830);
xnor UO_1269 (O_1269,N_19858,N_19932);
nand UO_1270 (O_1270,N_19997,N_19963);
nand UO_1271 (O_1271,N_19796,N_19873);
and UO_1272 (O_1272,N_19843,N_19813);
nor UO_1273 (O_1273,N_19831,N_19766);
and UO_1274 (O_1274,N_19970,N_19897);
nand UO_1275 (O_1275,N_19918,N_19853);
xnor UO_1276 (O_1276,N_19791,N_19928);
nor UO_1277 (O_1277,N_19919,N_19995);
nand UO_1278 (O_1278,N_19826,N_19890);
nand UO_1279 (O_1279,N_19875,N_19972);
nor UO_1280 (O_1280,N_19910,N_19819);
nand UO_1281 (O_1281,N_19845,N_19884);
nand UO_1282 (O_1282,N_19812,N_19811);
xor UO_1283 (O_1283,N_19814,N_19812);
or UO_1284 (O_1284,N_19787,N_19752);
or UO_1285 (O_1285,N_19858,N_19879);
and UO_1286 (O_1286,N_19955,N_19841);
nor UO_1287 (O_1287,N_19797,N_19985);
xor UO_1288 (O_1288,N_19932,N_19980);
or UO_1289 (O_1289,N_19772,N_19930);
nand UO_1290 (O_1290,N_19868,N_19939);
and UO_1291 (O_1291,N_19795,N_19824);
nand UO_1292 (O_1292,N_19827,N_19837);
or UO_1293 (O_1293,N_19827,N_19799);
nand UO_1294 (O_1294,N_19800,N_19833);
and UO_1295 (O_1295,N_19862,N_19826);
and UO_1296 (O_1296,N_19966,N_19763);
or UO_1297 (O_1297,N_19959,N_19998);
xor UO_1298 (O_1298,N_19871,N_19937);
nor UO_1299 (O_1299,N_19762,N_19779);
or UO_1300 (O_1300,N_19928,N_19778);
nand UO_1301 (O_1301,N_19809,N_19932);
and UO_1302 (O_1302,N_19933,N_19867);
nor UO_1303 (O_1303,N_19756,N_19876);
and UO_1304 (O_1304,N_19975,N_19770);
and UO_1305 (O_1305,N_19755,N_19778);
nor UO_1306 (O_1306,N_19841,N_19755);
and UO_1307 (O_1307,N_19925,N_19978);
nor UO_1308 (O_1308,N_19898,N_19807);
or UO_1309 (O_1309,N_19866,N_19895);
or UO_1310 (O_1310,N_19814,N_19888);
and UO_1311 (O_1311,N_19837,N_19857);
nor UO_1312 (O_1312,N_19886,N_19873);
and UO_1313 (O_1313,N_19890,N_19977);
and UO_1314 (O_1314,N_19935,N_19982);
nand UO_1315 (O_1315,N_19809,N_19777);
nand UO_1316 (O_1316,N_19861,N_19988);
nand UO_1317 (O_1317,N_19808,N_19892);
or UO_1318 (O_1318,N_19847,N_19825);
nor UO_1319 (O_1319,N_19987,N_19826);
xor UO_1320 (O_1320,N_19913,N_19991);
xor UO_1321 (O_1321,N_19780,N_19953);
or UO_1322 (O_1322,N_19759,N_19853);
nor UO_1323 (O_1323,N_19908,N_19796);
and UO_1324 (O_1324,N_19901,N_19967);
and UO_1325 (O_1325,N_19870,N_19908);
and UO_1326 (O_1326,N_19826,N_19830);
nor UO_1327 (O_1327,N_19965,N_19913);
nand UO_1328 (O_1328,N_19871,N_19894);
nor UO_1329 (O_1329,N_19869,N_19893);
nand UO_1330 (O_1330,N_19772,N_19875);
and UO_1331 (O_1331,N_19770,N_19787);
nand UO_1332 (O_1332,N_19911,N_19950);
nor UO_1333 (O_1333,N_19833,N_19999);
xnor UO_1334 (O_1334,N_19851,N_19902);
xor UO_1335 (O_1335,N_19783,N_19804);
nand UO_1336 (O_1336,N_19904,N_19760);
or UO_1337 (O_1337,N_19772,N_19840);
nor UO_1338 (O_1338,N_19937,N_19941);
and UO_1339 (O_1339,N_19948,N_19919);
and UO_1340 (O_1340,N_19898,N_19785);
or UO_1341 (O_1341,N_19924,N_19994);
nor UO_1342 (O_1342,N_19994,N_19756);
or UO_1343 (O_1343,N_19885,N_19997);
and UO_1344 (O_1344,N_19914,N_19845);
or UO_1345 (O_1345,N_19871,N_19898);
xor UO_1346 (O_1346,N_19972,N_19899);
xor UO_1347 (O_1347,N_19872,N_19928);
nor UO_1348 (O_1348,N_19953,N_19902);
nor UO_1349 (O_1349,N_19938,N_19881);
xnor UO_1350 (O_1350,N_19825,N_19959);
nand UO_1351 (O_1351,N_19989,N_19793);
and UO_1352 (O_1352,N_19801,N_19944);
nor UO_1353 (O_1353,N_19781,N_19917);
xor UO_1354 (O_1354,N_19936,N_19925);
nand UO_1355 (O_1355,N_19901,N_19754);
or UO_1356 (O_1356,N_19790,N_19879);
or UO_1357 (O_1357,N_19821,N_19791);
nor UO_1358 (O_1358,N_19855,N_19849);
nor UO_1359 (O_1359,N_19990,N_19978);
or UO_1360 (O_1360,N_19925,N_19828);
nand UO_1361 (O_1361,N_19811,N_19973);
or UO_1362 (O_1362,N_19951,N_19915);
xnor UO_1363 (O_1363,N_19937,N_19803);
xor UO_1364 (O_1364,N_19806,N_19753);
nand UO_1365 (O_1365,N_19870,N_19917);
nor UO_1366 (O_1366,N_19759,N_19855);
nand UO_1367 (O_1367,N_19800,N_19858);
or UO_1368 (O_1368,N_19895,N_19973);
nand UO_1369 (O_1369,N_19842,N_19824);
nor UO_1370 (O_1370,N_19967,N_19861);
xnor UO_1371 (O_1371,N_19986,N_19815);
xor UO_1372 (O_1372,N_19817,N_19750);
or UO_1373 (O_1373,N_19807,N_19937);
or UO_1374 (O_1374,N_19764,N_19806);
nor UO_1375 (O_1375,N_19913,N_19956);
or UO_1376 (O_1376,N_19965,N_19909);
nand UO_1377 (O_1377,N_19807,N_19770);
nand UO_1378 (O_1378,N_19767,N_19751);
xor UO_1379 (O_1379,N_19820,N_19764);
or UO_1380 (O_1380,N_19896,N_19819);
nand UO_1381 (O_1381,N_19816,N_19770);
xnor UO_1382 (O_1382,N_19806,N_19792);
xor UO_1383 (O_1383,N_19976,N_19818);
and UO_1384 (O_1384,N_19752,N_19837);
and UO_1385 (O_1385,N_19983,N_19816);
nand UO_1386 (O_1386,N_19993,N_19920);
nor UO_1387 (O_1387,N_19783,N_19852);
nand UO_1388 (O_1388,N_19770,N_19872);
nand UO_1389 (O_1389,N_19995,N_19976);
nand UO_1390 (O_1390,N_19851,N_19898);
xnor UO_1391 (O_1391,N_19937,N_19750);
nor UO_1392 (O_1392,N_19811,N_19843);
or UO_1393 (O_1393,N_19961,N_19817);
or UO_1394 (O_1394,N_19763,N_19876);
xnor UO_1395 (O_1395,N_19835,N_19799);
or UO_1396 (O_1396,N_19927,N_19951);
nand UO_1397 (O_1397,N_19790,N_19870);
xor UO_1398 (O_1398,N_19875,N_19974);
nand UO_1399 (O_1399,N_19928,N_19887);
and UO_1400 (O_1400,N_19758,N_19848);
nor UO_1401 (O_1401,N_19788,N_19789);
nor UO_1402 (O_1402,N_19933,N_19975);
nand UO_1403 (O_1403,N_19840,N_19932);
nor UO_1404 (O_1404,N_19925,N_19816);
and UO_1405 (O_1405,N_19897,N_19770);
nor UO_1406 (O_1406,N_19979,N_19877);
nor UO_1407 (O_1407,N_19887,N_19951);
and UO_1408 (O_1408,N_19797,N_19996);
and UO_1409 (O_1409,N_19808,N_19948);
or UO_1410 (O_1410,N_19870,N_19814);
nand UO_1411 (O_1411,N_19865,N_19944);
nor UO_1412 (O_1412,N_19865,N_19824);
or UO_1413 (O_1413,N_19810,N_19771);
xor UO_1414 (O_1414,N_19966,N_19914);
nor UO_1415 (O_1415,N_19856,N_19935);
nor UO_1416 (O_1416,N_19813,N_19892);
and UO_1417 (O_1417,N_19814,N_19935);
or UO_1418 (O_1418,N_19753,N_19835);
xnor UO_1419 (O_1419,N_19866,N_19915);
or UO_1420 (O_1420,N_19926,N_19958);
nor UO_1421 (O_1421,N_19939,N_19755);
or UO_1422 (O_1422,N_19973,N_19963);
or UO_1423 (O_1423,N_19871,N_19938);
and UO_1424 (O_1424,N_19763,N_19916);
xnor UO_1425 (O_1425,N_19801,N_19867);
or UO_1426 (O_1426,N_19933,N_19821);
and UO_1427 (O_1427,N_19863,N_19902);
xor UO_1428 (O_1428,N_19781,N_19816);
and UO_1429 (O_1429,N_19890,N_19857);
and UO_1430 (O_1430,N_19822,N_19795);
nand UO_1431 (O_1431,N_19916,N_19995);
or UO_1432 (O_1432,N_19758,N_19909);
nor UO_1433 (O_1433,N_19944,N_19886);
nand UO_1434 (O_1434,N_19947,N_19773);
nand UO_1435 (O_1435,N_19761,N_19810);
xnor UO_1436 (O_1436,N_19784,N_19844);
nor UO_1437 (O_1437,N_19921,N_19849);
or UO_1438 (O_1438,N_19763,N_19910);
nand UO_1439 (O_1439,N_19981,N_19844);
xnor UO_1440 (O_1440,N_19900,N_19831);
or UO_1441 (O_1441,N_19764,N_19808);
xor UO_1442 (O_1442,N_19999,N_19872);
and UO_1443 (O_1443,N_19936,N_19967);
nand UO_1444 (O_1444,N_19903,N_19984);
nor UO_1445 (O_1445,N_19930,N_19838);
xor UO_1446 (O_1446,N_19920,N_19930);
nand UO_1447 (O_1447,N_19859,N_19792);
and UO_1448 (O_1448,N_19959,N_19840);
nor UO_1449 (O_1449,N_19946,N_19758);
nor UO_1450 (O_1450,N_19886,N_19757);
nor UO_1451 (O_1451,N_19843,N_19771);
nand UO_1452 (O_1452,N_19837,N_19830);
xnor UO_1453 (O_1453,N_19853,N_19816);
and UO_1454 (O_1454,N_19972,N_19931);
and UO_1455 (O_1455,N_19752,N_19809);
or UO_1456 (O_1456,N_19830,N_19868);
nand UO_1457 (O_1457,N_19855,N_19981);
xor UO_1458 (O_1458,N_19809,N_19914);
or UO_1459 (O_1459,N_19772,N_19785);
xnor UO_1460 (O_1460,N_19883,N_19895);
nor UO_1461 (O_1461,N_19911,N_19980);
or UO_1462 (O_1462,N_19996,N_19906);
or UO_1463 (O_1463,N_19992,N_19925);
nor UO_1464 (O_1464,N_19758,N_19825);
nor UO_1465 (O_1465,N_19886,N_19812);
nand UO_1466 (O_1466,N_19793,N_19794);
nand UO_1467 (O_1467,N_19924,N_19896);
xor UO_1468 (O_1468,N_19777,N_19852);
or UO_1469 (O_1469,N_19850,N_19790);
or UO_1470 (O_1470,N_19766,N_19912);
xor UO_1471 (O_1471,N_19813,N_19768);
nor UO_1472 (O_1472,N_19771,N_19963);
or UO_1473 (O_1473,N_19832,N_19865);
xor UO_1474 (O_1474,N_19948,N_19964);
nor UO_1475 (O_1475,N_19830,N_19909);
and UO_1476 (O_1476,N_19766,N_19834);
nor UO_1477 (O_1477,N_19890,N_19912);
nor UO_1478 (O_1478,N_19922,N_19761);
nor UO_1479 (O_1479,N_19821,N_19750);
nor UO_1480 (O_1480,N_19927,N_19860);
and UO_1481 (O_1481,N_19841,N_19823);
or UO_1482 (O_1482,N_19915,N_19963);
nor UO_1483 (O_1483,N_19768,N_19877);
nand UO_1484 (O_1484,N_19940,N_19793);
or UO_1485 (O_1485,N_19954,N_19909);
and UO_1486 (O_1486,N_19822,N_19935);
or UO_1487 (O_1487,N_19771,N_19949);
nand UO_1488 (O_1488,N_19847,N_19793);
nor UO_1489 (O_1489,N_19970,N_19826);
xnor UO_1490 (O_1490,N_19768,N_19758);
and UO_1491 (O_1491,N_19900,N_19897);
nand UO_1492 (O_1492,N_19939,N_19902);
or UO_1493 (O_1493,N_19814,N_19825);
nor UO_1494 (O_1494,N_19768,N_19924);
and UO_1495 (O_1495,N_19925,N_19949);
or UO_1496 (O_1496,N_19955,N_19937);
xnor UO_1497 (O_1497,N_19876,N_19892);
and UO_1498 (O_1498,N_19976,N_19750);
and UO_1499 (O_1499,N_19808,N_19794);
and UO_1500 (O_1500,N_19872,N_19843);
and UO_1501 (O_1501,N_19900,N_19778);
or UO_1502 (O_1502,N_19966,N_19783);
and UO_1503 (O_1503,N_19828,N_19986);
and UO_1504 (O_1504,N_19797,N_19782);
nor UO_1505 (O_1505,N_19776,N_19865);
xor UO_1506 (O_1506,N_19750,N_19864);
nor UO_1507 (O_1507,N_19756,N_19752);
or UO_1508 (O_1508,N_19765,N_19772);
nand UO_1509 (O_1509,N_19929,N_19920);
xnor UO_1510 (O_1510,N_19912,N_19930);
nand UO_1511 (O_1511,N_19820,N_19796);
or UO_1512 (O_1512,N_19824,N_19847);
or UO_1513 (O_1513,N_19769,N_19770);
and UO_1514 (O_1514,N_19815,N_19840);
nor UO_1515 (O_1515,N_19834,N_19915);
nand UO_1516 (O_1516,N_19902,N_19854);
or UO_1517 (O_1517,N_19754,N_19870);
nand UO_1518 (O_1518,N_19875,N_19767);
nor UO_1519 (O_1519,N_19835,N_19787);
or UO_1520 (O_1520,N_19885,N_19883);
and UO_1521 (O_1521,N_19976,N_19970);
nand UO_1522 (O_1522,N_19883,N_19840);
nand UO_1523 (O_1523,N_19886,N_19816);
nor UO_1524 (O_1524,N_19952,N_19834);
and UO_1525 (O_1525,N_19875,N_19754);
nand UO_1526 (O_1526,N_19925,N_19877);
xor UO_1527 (O_1527,N_19984,N_19906);
and UO_1528 (O_1528,N_19763,N_19798);
xnor UO_1529 (O_1529,N_19959,N_19933);
nand UO_1530 (O_1530,N_19937,N_19861);
and UO_1531 (O_1531,N_19862,N_19952);
nor UO_1532 (O_1532,N_19892,N_19826);
or UO_1533 (O_1533,N_19767,N_19771);
and UO_1534 (O_1534,N_19762,N_19849);
and UO_1535 (O_1535,N_19998,N_19771);
nand UO_1536 (O_1536,N_19757,N_19870);
or UO_1537 (O_1537,N_19812,N_19833);
xor UO_1538 (O_1538,N_19756,N_19761);
or UO_1539 (O_1539,N_19959,N_19854);
nand UO_1540 (O_1540,N_19794,N_19996);
and UO_1541 (O_1541,N_19762,N_19809);
and UO_1542 (O_1542,N_19780,N_19889);
nand UO_1543 (O_1543,N_19861,N_19753);
and UO_1544 (O_1544,N_19798,N_19931);
nor UO_1545 (O_1545,N_19871,N_19944);
or UO_1546 (O_1546,N_19799,N_19770);
and UO_1547 (O_1547,N_19752,N_19807);
and UO_1548 (O_1548,N_19923,N_19825);
nand UO_1549 (O_1549,N_19796,N_19754);
xor UO_1550 (O_1550,N_19890,N_19814);
xor UO_1551 (O_1551,N_19753,N_19855);
or UO_1552 (O_1552,N_19801,N_19970);
xnor UO_1553 (O_1553,N_19750,N_19945);
xor UO_1554 (O_1554,N_19825,N_19982);
xor UO_1555 (O_1555,N_19972,N_19879);
and UO_1556 (O_1556,N_19879,N_19928);
nand UO_1557 (O_1557,N_19878,N_19907);
xnor UO_1558 (O_1558,N_19832,N_19872);
nand UO_1559 (O_1559,N_19920,N_19810);
nand UO_1560 (O_1560,N_19840,N_19943);
or UO_1561 (O_1561,N_19957,N_19966);
or UO_1562 (O_1562,N_19834,N_19980);
xnor UO_1563 (O_1563,N_19853,N_19914);
nand UO_1564 (O_1564,N_19841,N_19868);
nor UO_1565 (O_1565,N_19827,N_19847);
nand UO_1566 (O_1566,N_19863,N_19916);
nand UO_1567 (O_1567,N_19909,N_19865);
xnor UO_1568 (O_1568,N_19752,N_19907);
nand UO_1569 (O_1569,N_19781,N_19954);
or UO_1570 (O_1570,N_19914,N_19939);
nand UO_1571 (O_1571,N_19932,N_19759);
xnor UO_1572 (O_1572,N_19940,N_19963);
nand UO_1573 (O_1573,N_19781,N_19877);
or UO_1574 (O_1574,N_19909,N_19883);
and UO_1575 (O_1575,N_19755,N_19876);
nor UO_1576 (O_1576,N_19807,N_19881);
nand UO_1577 (O_1577,N_19896,N_19990);
and UO_1578 (O_1578,N_19847,N_19769);
nor UO_1579 (O_1579,N_19837,N_19982);
and UO_1580 (O_1580,N_19846,N_19995);
and UO_1581 (O_1581,N_19911,N_19753);
nand UO_1582 (O_1582,N_19792,N_19750);
or UO_1583 (O_1583,N_19898,N_19841);
nand UO_1584 (O_1584,N_19908,N_19885);
nor UO_1585 (O_1585,N_19882,N_19979);
and UO_1586 (O_1586,N_19915,N_19759);
and UO_1587 (O_1587,N_19796,N_19821);
xnor UO_1588 (O_1588,N_19796,N_19784);
nand UO_1589 (O_1589,N_19916,N_19767);
and UO_1590 (O_1590,N_19896,N_19962);
xnor UO_1591 (O_1591,N_19912,N_19915);
xnor UO_1592 (O_1592,N_19912,N_19916);
or UO_1593 (O_1593,N_19796,N_19890);
xor UO_1594 (O_1594,N_19952,N_19820);
nor UO_1595 (O_1595,N_19980,N_19912);
nand UO_1596 (O_1596,N_19852,N_19859);
nor UO_1597 (O_1597,N_19837,N_19968);
nand UO_1598 (O_1598,N_19831,N_19883);
nor UO_1599 (O_1599,N_19827,N_19858);
and UO_1600 (O_1600,N_19851,N_19985);
nor UO_1601 (O_1601,N_19908,N_19760);
nor UO_1602 (O_1602,N_19881,N_19855);
xnor UO_1603 (O_1603,N_19859,N_19795);
nand UO_1604 (O_1604,N_19750,N_19759);
or UO_1605 (O_1605,N_19932,N_19901);
nand UO_1606 (O_1606,N_19881,N_19972);
nor UO_1607 (O_1607,N_19869,N_19916);
xor UO_1608 (O_1608,N_19850,N_19829);
xnor UO_1609 (O_1609,N_19805,N_19982);
and UO_1610 (O_1610,N_19800,N_19812);
and UO_1611 (O_1611,N_19918,N_19943);
nor UO_1612 (O_1612,N_19891,N_19818);
or UO_1613 (O_1613,N_19768,N_19762);
and UO_1614 (O_1614,N_19820,N_19910);
xor UO_1615 (O_1615,N_19762,N_19975);
nand UO_1616 (O_1616,N_19798,N_19939);
nor UO_1617 (O_1617,N_19927,N_19813);
nand UO_1618 (O_1618,N_19952,N_19909);
or UO_1619 (O_1619,N_19987,N_19930);
nor UO_1620 (O_1620,N_19960,N_19907);
nand UO_1621 (O_1621,N_19907,N_19936);
or UO_1622 (O_1622,N_19856,N_19861);
nor UO_1623 (O_1623,N_19885,N_19924);
nand UO_1624 (O_1624,N_19964,N_19985);
nor UO_1625 (O_1625,N_19791,N_19848);
nand UO_1626 (O_1626,N_19935,N_19875);
nor UO_1627 (O_1627,N_19783,N_19974);
xor UO_1628 (O_1628,N_19816,N_19911);
nand UO_1629 (O_1629,N_19953,N_19803);
xnor UO_1630 (O_1630,N_19819,N_19954);
or UO_1631 (O_1631,N_19773,N_19965);
xnor UO_1632 (O_1632,N_19934,N_19756);
nor UO_1633 (O_1633,N_19971,N_19761);
nor UO_1634 (O_1634,N_19799,N_19862);
nand UO_1635 (O_1635,N_19799,N_19899);
nor UO_1636 (O_1636,N_19902,N_19961);
and UO_1637 (O_1637,N_19905,N_19760);
nor UO_1638 (O_1638,N_19756,N_19975);
and UO_1639 (O_1639,N_19791,N_19943);
and UO_1640 (O_1640,N_19992,N_19883);
xor UO_1641 (O_1641,N_19979,N_19969);
nor UO_1642 (O_1642,N_19917,N_19773);
nor UO_1643 (O_1643,N_19913,N_19886);
and UO_1644 (O_1644,N_19760,N_19910);
and UO_1645 (O_1645,N_19876,N_19858);
nand UO_1646 (O_1646,N_19942,N_19915);
or UO_1647 (O_1647,N_19823,N_19754);
nand UO_1648 (O_1648,N_19767,N_19796);
nand UO_1649 (O_1649,N_19849,N_19882);
nor UO_1650 (O_1650,N_19940,N_19810);
or UO_1651 (O_1651,N_19776,N_19772);
xnor UO_1652 (O_1652,N_19865,N_19983);
nand UO_1653 (O_1653,N_19759,N_19770);
nand UO_1654 (O_1654,N_19932,N_19933);
and UO_1655 (O_1655,N_19755,N_19974);
nand UO_1656 (O_1656,N_19771,N_19895);
nor UO_1657 (O_1657,N_19886,N_19994);
nand UO_1658 (O_1658,N_19850,N_19791);
xor UO_1659 (O_1659,N_19852,N_19989);
xor UO_1660 (O_1660,N_19755,N_19773);
nand UO_1661 (O_1661,N_19811,N_19766);
nand UO_1662 (O_1662,N_19870,N_19956);
xor UO_1663 (O_1663,N_19970,N_19943);
and UO_1664 (O_1664,N_19895,N_19870);
and UO_1665 (O_1665,N_19866,N_19813);
or UO_1666 (O_1666,N_19924,N_19922);
nor UO_1667 (O_1667,N_19799,N_19970);
nand UO_1668 (O_1668,N_19980,N_19925);
or UO_1669 (O_1669,N_19869,N_19908);
or UO_1670 (O_1670,N_19756,N_19997);
nand UO_1671 (O_1671,N_19755,N_19971);
nand UO_1672 (O_1672,N_19956,N_19932);
or UO_1673 (O_1673,N_19775,N_19855);
and UO_1674 (O_1674,N_19844,N_19925);
nor UO_1675 (O_1675,N_19880,N_19993);
nand UO_1676 (O_1676,N_19808,N_19905);
and UO_1677 (O_1677,N_19968,N_19845);
nor UO_1678 (O_1678,N_19888,N_19832);
nand UO_1679 (O_1679,N_19968,N_19947);
nand UO_1680 (O_1680,N_19852,N_19754);
or UO_1681 (O_1681,N_19861,N_19959);
or UO_1682 (O_1682,N_19908,N_19913);
xor UO_1683 (O_1683,N_19924,N_19910);
xor UO_1684 (O_1684,N_19963,N_19804);
or UO_1685 (O_1685,N_19907,N_19973);
and UO_1686 (O_1686,N_19942,N_19817);
or UO_1687 (O_1687,N_19846,N_19825);
or UO_1688 (O_1688,N_19898,N_19984);
and UO_1689 (O_1689,N_19979,N_19914);
or UO_1690 (O_1690,N_19890,N_19787);
nor UO_1691 (O_1691,N_19972,N_19934);
and UO_1692 (O_1692,N_19833,N_19913);
xor UO_1693 (O_1693,N_19986,N_19859);
xor UO_1694 (O_1694,N_19955,N_19894);
or UO_1695 (O_1695,N_19774,N_19968);
xnor UO_1696 (O_1696,N_19933,N_19920);
or UO_1697 (O_1697,N_19842,N_19808);
and UO_1698 (O_1698,N_19757,N_19910);
nor UO_1699 (O_1699,N_19986,N_19985);
nand UO_1700 (O_1700,N_19842,N_19952);
nand UO_1701 (O_1701,N_19799,N_19957);
nand UO_1702 (O_1702,N_19853,N_19941);
and UO_1703 (O_1703,N_19834,N_19925);
nand UO_1704 (O_1704,N_19896,N_19983);
and UO_1705 (O_1705,N_19770,N_19864);
nand UO_1706 (O_1706,N_19860,N_19811);
or UO_1707 (O_1707,N_19899,N_19802);
nor UO_1708 (O_1708,N_19920,N_19849);
and UO_1709 (O_1709,N_19994,N_19932);
and UO_1710 (O_1710,N_19781,N_19880);
xor UO_1711 (O_1711,N_19766,N_19871);
nand UO_1712 (O_1712,N_19874,N_19753);
or UO_1713 (O_1713,N_19976,N_19908);
xor UO_1714 (O_1714,N_19802,N_19765);
nand UO_1715 (O_1715,N_19764,N_19824);
xor UO_1716 (O_1716,N_19926,N_19983);
nor UO_1717 (O_1717,N_19850,N_19828);
or UO_1718 (O_1718,N_19980,N_19788);
nand UO_1719 (O_1719,N_19819,N_19760);
nor UO_1720 (O_1720,N_19902,N_19768);
or UO_1721 (O_1721,N_19948,N_19767);
nor UO_1722 (O_1722,N_19860,N_19878);
xnor UO_1723 (O_1723,N_19853,N_19752);
xor UO_1724 (O_1724,N_19764,N_19753);
nand UO_1725 (O_1725,N_19977,N_19804);
and UO_1726 (O_1726,N_19907,N_19771);
and UO_1727 (O_1727,N_19750,N_19961);
nor UO_1728 (O_1728,N_19786,N_19792);
nor UO_1729 (O_1729,N_19979,N_19974);
nand UO_1730 (O_1730,N_19860,N_19881);
nand UO_1731 (O_1731,N_19813,N_19785);
nor UO_1732 (O_1732,N_19793,N_19874);
nor UO_1733 (O_1733,N_19839,N_19819);
nand UO_1734 (O_1734,N_19909,N_19831);
and UO_1735 (O_1735,N_19845,N_19969);
and UO_1736 (O_1736,N_19994,N_19948);
xor UO_1737 (O_1737,N_19915,N_19796);
nand UO_1738 (O_1738,N_19820,N_19860);
nand UO_1739 (O_1739,N_19879,N_19893);
nor UO_1740 (O_1740,N_19917,N_19980);
nor UO_1741 (O_1741,N_19835,N_19995);
nand UO_1742 (O_1742,N_19945,N_19953);
and UO_1743 (O_1743,N_19956,N_19826);
nor UO_1744 (O_1744,N_19913,N_19905);
nand UO_1745 (O_1745,N_19757,N_19914);
nand UO_1746 (O_1746,N_19767,N_19856);
or UO_1747 (O_1747,N_19845,N_19983);
and UO_1748 (O_1748,N_19958,N_19895);
nor UO_1749 (O_1749,N_19874,N_19853);
and UO_1750 (O_1750,N_19792,N_19883);
nor UO_1751 (O_1751,N_19957,N_19815);
nor UO_1752 (O_1752,N_19786,N_19778);
and UO_1753 (O_1753,N_19945,N_19927);
xor UO_1754 (O_1754,N_19971,N_19880);
or UO_1755 (O_1755,N_19792,N_19968);
xnor UO_1756 (O_1756,N_19991,N_19900);
or UO_1757 (O_1757,N_19801,N_19998);
or UO_1758 (O_1758,N_19981,N_19802);
and UO_1759 (O_1759,N_19824,N_19769);
nor UO_1760 (O_1760,N_19943,N_19816);
or UO_1761 (O_1761,N_19849,N_19962);
and UO_1762 (O_1762,N_19980,N_19958);
and UO_1763 (O_1763,N_19960,N_19824);
nand UO_1764 (O_1764,N_19928,N_19770);
xor UO_1765 (O_1765,N_19957,N_19914);
and UO_1766 (O_1766,N_19970,N_19875);
and UO_1767 (O_1767,N_19893,N_19983);
and UO_1768 (O_1768,N_19879,N_19817);
and UO_1769 (O_1769,N_19826,N_19997);
or UO_1770 (O_1770,N_19843,N_19796);
xor UO_1771 (O_1771,N_19827,N_19751);
nor UO_1772 (O_1772,N_19983,N_19937);
nand UO_1773 (O_1773,N_19922,N_19792);
nor UO_1774 (O_1774,N_19858,N_19834);
or UO_1775 (O_1775,N_19921,N_19898);
nand UO_1776 (O_1776,N_19985,N_19995);
and UO_1777 (O_1777,N_19909,N_19961);
xor UO_1778 (O_1778,N_19778,N_19884);
or UO_1779 (O_1779,N_19947,N_19980);
xnor UO_1780 (O_1780,N_19801,N_19897);
xor UO_1781 (O_1781,N_19755,N_19946);
and UO_1782 (O_1782,N_19990,N_19791);
xnor UO_1783 (O_1783,N_19771,N_19830);
and UO_1784 (O_1784,N_19853,N_19954);
nand UO_1785 (O_1785,N_19893,N_19978);
xor UO_1786 (O_1786,N_19786,N_19951);
nor UO_1787 (O_1787,N_19898,N_19840);
nand UO_1788 (O_1788,N_19862,N_19893);
xnor UO_1789 (O_1789,N_19970,N_19998);
nand UO_1790 (O_1790,N_19968,N_19788);
xnor UO_1791 (O_1791,N_19898,N_19850);
or UO_1792 (O_1792,N_19891,N_19956);
nand UO_1793 (O_1793,N_19956,N_19965);
nor UO_1794 (O_1794,N_19949,N_19803);
nand UO_1795 (O_1795,N_19855,N_19973);
xor UO_1796 (O_1796,N_19803,N_19867);
nor UO_1797 (O_1797,N_19959,N_19994);
nor UO_1798 (O_1798,N_19850,N_19841);
xor UO_1799 (O_1799,N_19903,N_19809);
xor UO_1800 (O_1800,N_19848,N_19761);
and UO_1801 (O_1801,N_19892,N_19907);
xnor UO_1802 (O_1802,N_19923,N_19859);
and UO_1803 (O_1803,N_19823,N_19772);
xnor UO_1804 (O_1804,N_19926,N_19955);
nand UO_1805 (O_1805,N_19896,N_19878);
nor UO_1806 (O_1806,N_19841,N_19960);
or UO_1807 (O_1807,N_19773,N_19883);
and UO_1808 (O_1808,N_19805,N_19896);
and UO_1809 (O_1809,N_19826,N_19897);
xor UO_1810 (O_1810,N_19846,N_19932);
nor UO_1811 (O_1811,N_19911,N_19872);
or UO_1812 (O_1812,N_19891,N_19976);
nor UO_1813 (O_1813,N_19919,N_19878);
or UO_1814 (O_1814,N_19825,N_19934);
nor UO_1815 (O_1815,N_19950,N_19888);
nor UO_1816 (O_1816,N_19845,N_19806);
or UO_1817 (O_1817,N_19829,N_19955);
and UO_1818 (O_1818,N_19919,N_19928);
nor UO_1819 (O_1819,N_19963,N_19782);
xor UO_1820 (O_1820,N_19882,N_19868);
nand UO_1821 (O_1821,N_19936,N_19881);
and UO_1822 (O_1822,N_19772,N_19792);
nand UO_1823 (O_1823,N_19971,N_19915);
nor UO_1824 (O_1824,N_19767,N_19937);
xnor UO_1825 (O_1825,N_19833,N_19816);
or UO_1826 (O_1826,N_19888,N_19917);
nand UO_1827 (O_1827,N_19932,N_19849);
nand UO_1828 (O_1828,N_19838,N_19858);
nand UO_1829 (O_1829,N_19993,N_19882);
nor UO_1830 (O_1830,N_19835,N_19780);
nor UO_1831 (O_1831,N_19811,N_19850);
or UO_1832 (O_1832,N_19988,N_19760);
and UO_1833 (O_1833,N_19989,N_19908);
xor UO_1834 (O_1834,N_19796,N_19766);
and UO_1835 (O_1835,N_19829,N_19781);
nand UO_1836 (O_1836,N_19818,N_19826);
or UO_1837 (O_1837,N_19771,N_19993);
nor UO_1838 (O_1838,N_19957,N_19983);
xor UO_1839 (O_1839,N_19953,N_19956);
xor UO_1840 (O_1840,N_19916,N_19908);
nand UO_1841 (O_1841,N_19962,N_19964);
xnor UO_1842 (O_1842,N_19848,N_19822);
or UO_1843 (O_1843,N_19936,N_19951);
or UO_1844 (O_1844,N_19821,N_19988);
nand UO_1845 (O_1845,N_19891,N_19834);
or UO_1846 (O_1846,N_19973,N_19930);
nor UO_1847 (O_1847,N_19848,N_19997);
nor UO_1848 (O_1848,N_19808,N_19780);
nand UO_1849 (O_1849,N_19963,N_19809);
nand UO_1850 (O_1850,N_19760,N_19822);
and UO_1851 (O_1851,N_19929,N_19810);
and UO_1852 (O_1852,N_19751,N_19825);
xor UO_1853 (O_1853,N_19927,N_19937);
nor UO_1854 (O_1854,N_19800,N_19849);
xor UO_1855 (O_1855,N_19965,N_19823);
and UO_1856 (O_1856,N_19799,N_19847);
xnor UO_1857 (O_1857,N_19774,N_19883);
xor UO_1858 (O_1858,N_19889,N_19953);
nor UO_1859 (O_1859,N_19854,N_19999);
xor UO_1860 (O_1860,N_19886,N_19962);
or UO_1861 (O_1861,N_19894,N_19840);
and UO_1862 (O_1862,N_19942,N_19857);
nand UO_1863 (O_1863,N_19954,N_19877);
or UO_1864 (O_1864,N_19970,N_19899);
and UO_1865 (O_1865,N_19863,N_19987);
nand UO_1866 (O_1866,N_19888,N_19982);
nand UO_1867 (O_1867,N_19791,N_19941);
or UO_1868 (O_1868,N_19777,N_19823);
or UO_1869 (O_1869,N_19872,N_19841);
and UO_1870 (O_1870,N_19867,N_19851);
and UO_1871 (O_1871,N_19856,N_19979);
nand UO_1872 (O_1872,N_19794,N_19799);
and UO_1873 (O_1873,N_19944,N_19774);
nor UO_1874 (O_1874,N_19848,N_19788);
nand UO_1875 (O_1875,N_19904,N_19937);
xnor UO_1876 (O_1876,N_19781,N_19914);
nor UO_1877 (O_1877,N_19958,N_19757);
and UO_1878 (O_1878,N_19949,N_19909);
nand UO_1879 (O_1879,N_19860,N_19952);
nand UO_1880 (O_1880,N_19851,N_19899);
and UO_1881 (O_1881,N_19979,N_19893);
nand UO_1882 (O_1882,N_19809,N_19978);
xnor UO_1883 (O_1883,N_19889,N_19893);
nor UO_1884 (O_1884,N_19794,N_19895);
nand UO_1885 (O_1885,N_19756,N_19998);
or UO_1886 (O_1886,N_19819,N_19809);
nand UO_1887 (O_1887,N_19788,N_19775);
nand UO_1888 (O_1888,N_19964,N_19791);
and UO_1889 (O_1889,N_19867,N_19983);
xnor UO_1890 (O_1890,N_19877,N_19844);
xor UO_1891 (O_1891,N_19852,N_19970);
nor UO_1892 (O_1892,N_19754,N_19919);
nand UO_1893 (O_1893,N_19940,N_19881);
nor UO_1894 (O_1894,N_19792,N_19967);
nand UO_1895 (O_1895,N_19820,N_19946);
and UO_1896 (O_1896,N_19823,N_19982);
and UO_1897 (O_1897,N_19811,N_19797);
or UO_1898 (O_1898,N_19959,N_19760);
nand UO_1899 (O_1899,N_19911,N_19802);
xnor UO_1900 (O_1900,N_19800,N_19784);
nor UO_1901 (O_1901,N_19803,N_19757);
and UO_1902 (O_1902,N_19823,N_19934);
nor UO_1903 (O_1903,N_19924,N_19957);
nand UO_1904 (O_1904,N_19825,N_19882);
xnor UO_1905 (O_1905,N_19858,N_19942);
nor UO_1906 (O_1906,N_19850,N_19985);
xnor UO_1907 (O_1907,N_19772,N_19904);
nor UO_1908 (O_1908,N_19946,N_19848);
xnor UO_1909 (O_1909,N_19986,N_19968);
and UO_1910 (O_1910,N_19992,N_19869);
and UO_1911 (O_1911,N_19971,N_19888);
nand UO_1912 (O_1912,N_19787,N_19971);
nand UO_1913 (O_1913,N_19759,N_19937);
nor UO_1914 (O_1914,N_19962,N_19900);
nor UO_1915 (O_1915,N_19973,N_19869);
xnor UO_1916 (O_1916,N_19912,N_19990);
xnor UO_1917 (O_1917,N_19794,N_19960);
nand UO_1918 (O_1918,N_19777,N_19838);
and UO_1919 (O_1919,N_19943,N_19851);
or UO_1920 (O_1920,N_19917,N_19769);
nand UO_1921 (O_1921,N_19779,N_19841);
and UO_1922 (O_1922,N_19825,N_19902);
nand UO_1923 (O_1923,N_19795,N_19935);
and UO_1924 (O_1924,N_19890,N_19966);
and UO_1925 (O_1925,N_19774,N_19965);
and UO_1926 (O_1926,N_19933,N_19965);
nand UO_1927 (O_1927,N_19880,N_19962);
and UO_1928 (O_1928,N_19765,N_19838);
or UO_1929 (O_1929,N_19962,N_19775);
nand UO_1930 (O_1930,N_19867,N_19778);
nor UO_1931 (O_1931,N_19830,N_19925);
nand UO_1932 (O_1932,N_19961,N_19999);
xnor UO_1933 (O_1933,N_19875,N_19898);
xor UO_1934 (O_1934,N_19847,N_19963);
xnor UO_1935 (O_1935,N_19867,N_19752);
xor UO_1936 (O_1936,N_19874,N_19918);
or UO_1937 (O_1937,N_19996,N_19751);
or UO_1938 (O_1938,N_19773,N_19778);
or UO_1939 (O_1939,N_19827,N_19903);
and UO_1940 (O_1940,N_19948,N_19924);
and UO_1941 (O_1941,N_19795,N_19953);
nor UO_1942 (O_1942,N_19792,N_19986);
nand UO_1943 (O_1943,N_19973,N_19916);
xor UO_1944 (O_1944,N_19904,N_19974);
nor UO_1945 (O_1945,N_19905,N_19977);
or UO_1946 (O_1946,N_19893,N_19976);
nand UO_1947 (O_1947,N_19753,N_19914);
nor UO_1948 (O_1948,N_19783,N_19768);
nor UO_1949 (O_1949,N_19803,N_19852);
xnor UO_1950 (O_1950,N_19808,N_19996);
nand UO_1951 (O_1951,N_19956,N_19833);
and UO_1952 (O_1952,N_19823,N_19883);
nor UO_1953 (O_1953,N_19958,N_19768);
and UO_1954 (O_1954,N_19831,N_19814);
nor UO_1955 (O_1955,N_19939,N_19770);
nor UO_1956 (O_1956,N_19837,N_19943);
and UO_1957 (O_1957,N_19879,N_19780);
or UO_1958 (O_1958,N_19960,N_19957);
xor UO_1959 (O_1959,N_19780,N_19983);
nand UO_1960 (O_1960,N_19991,N_19933);
nor UO_1961 (O_1961,N_19886,N_19917);
nor UO_1962 (O_1962,N_19945,N_19782);
nor UO_1963 (O_1963,N_19914,N_19878);
nand UO_1964 (O_1964,N_19804,N_19857);
xor UO_1965 (O_1965,N_19852,N_19917);
or UO_1966 (O_1966,N_19853,N_19991);
nor UO_1967 (O_1967,N_19825,N_19759);
and UO_1968 (O_1968,N_19829,N_19993);
xnor UO_1969 (O_1969,N_19965,N_19799);
nor UO_1970 (O_1970,N_19793,N_19873);
or UO_1971 (O_1971,N_19896,N_19870);
nand UO_1972 (O_1972,N_19808,N_19763);
nand UO_1973 (O_1973,N_19800,N_19818);
and UO_1974 (O_1974,N_19875,N_19996);
nor UO_1975 (O_1975,N_19870,N_19798);
or UO_1976 (O_1976,N_19891,N_19760);
xnor UO_1977 (O_1977,N_19873,N_19878);
nor UO_1978 (O_1978,N_19945,N_19803);
xor UO_1979 (O_1979,N_19974,N_19769);
or UO_1980 (O_1980,N_19881,N_19947);
nand UO_1981 (O_1981,N_19765,N_19771);
and UO_1982 (O_1982,N_19773,N_19849);
nor UO_1983 (O_1983,N_19935,N_19756);
or UO_1984 (O_1984,N_19974,N_19834);
nand UO_1985 (O_1985,N_19902,N_19861);
nand UO_1986 (O_1986,N_19803,N_19936);
or UO_1987 (O_1987,N_19958,N_19815);
and UO_1988 (O_1988,N_19847,N_19794);
or UO_1989 (O_1989,N_19846,N_19767);
xor UO_1990 (O_1990,N_19908,N_19751);
or UO_1991 (O_1991,N_19944,N_19799);
nand UO_1992 (O_1992,N_19942,N_19975);
xnor UO_1993 (O_1993,N_19752,N_19774);
and UO_1994 (O_1994,N_19779,N_19776);
and UO_1995 (O_1995,N_19951,N_19878);
nand UO_1996 (O_1996,N_19918,N_19799);
or UO_1997 (O_1997,N_19995,N_19787);
nand UO_1998 (O_1998,N_19902,N_19862);
nand UO_1999 (O_1999,N_19813,N_19805);
nand UO_2000 (O_2000,N_19964,N_19826);
nand UO_2001 (O_2001,N_19944,N_19762);
xnor UO_2002 (O_2002,N_19901,N_19891);
nand UO_2003 (O_2003,N_19837,N_19831);
xnor UO_2004 (O_2004,N_19958,N_19923);
xor UO_2005 (O_2005,N_19843,N_19815);
and UO_2006 (O_2006,N_19918,N_19953);
xnor UO_2007 (O_2007,N_19892,N_19771);
nor UO_2008 (O_2008,N_19936,N_19756);
nand UO_2009 (O_2009,N_19804,N_19865);
nand UO_2010 (O_2010,N_19783,N_19930);
xor UO_2011 (O_2011,N_19883,N_19976);
xnor UO_2012 (O_2012,N_19803,N_19817);
or UO_2013 (O_2013,N_19978,N_19820);
nor UO_2014 (O_2014,N_19904,N_19753);
nand UO_2015 (O_2015,N_19779,N_19832);
or UO_2016 (O_2016,N_19790,N_19809);
or UO_2017 (O_2017,N_19987,N_19790);
nand UO_2018 (O_2018,N_19864,N_19969);
nand UO_2019 (O_2019,N_19893,N_19771);
and UO_2020 (O_2020,N_19833,N_19867);
nand UO_2021 (O_2021,N_19957,N_19950);
and UO_2022 (O_2022,N_19957,N_19926);
and UO_2023 (O_2023,N_19858,N_19882);
nand UO_2024 (O_2024,N_19761,N_19937);
or UO_2025 (O_2025,N_19956,N_19764);
xor UO_2026 (O_2026,N_19832,N_19998);
or UO_2027 (O_2027,N_19792,N_19852);
nor UO_2028 (O_2028,N_19860,N_19998);
nand UO_2029 (O_2029,N_19917,N_19895);
or UO_2030 (O_2030,N_19825,N_19989);
or UO_2031 (O_2031,N_19875,N_19858);
or UO_2032 (O_2032,N_19990,N_19874);
or UO_2033 (O_2033,N_19769,N_19782);
and UO_2034 (O_2034,N_19922,N_19907);
or UO_2035 (O_2035,N_19801,N_19827);
xnor UO_2036 (O_2036,N_19880,N_19897);
xor UO_2037 (O_2037,N_19792,N_19776);
nor UO_2038 (O_2038,N_19962,N_19798);
or UO_2039 (O_2039,N_19919,N_19771);
and UO_2040 (O_2040,N_19839,N_19975);
nand UO_2041 (O_2041,N_19969,N_19971);
and UO_2042 (O_2042,N_19897,N_19879);
xor UO_2043 (O_2043,N_19812,N_19824);
or UO_2044 (O_2044,N_19996,N_19978);
or UO_2045 (O_2045,N_19750,N_19843);
and UO_2046 (O_2046,N_19816,N_19924);
nand UO_2047 (O_2047,N_19902,N_19909);
nand UO_2048 (O_2048,N_19877,N_19806);
xor UO_2049 (O_2049,N_19869,N_19755);
or UO_2050 (O_2050,N_19984,N_19804);
xnor UO_2051 (O_2051,N_19829,N_19897);
xnor UO_2052 (O_2052,N_19814,N_19964);
nand UO_2053 (O_2053,N_19963,N_19853);
xnor UO_2054 (O_2054,N_19971,N_19978);
nand UO_2055 (O_2055,N_19959,N_19792);
nand UO_2056 (O_2056,N_19850,N_19866);
and UO_2057 (O_2057,N_19786,N_19869);
nand UO_2058 (O_2058,N_19859,N_19880);
nand UO_2059 (O_2059,N_19855,N_19986);
nand UO_2060 (O_2060,N_19941,N_19916);
and UO_2061 (O_2061,N_19893,N_19815);
and UO_2062 (O_2062,N_19793,N_19832);
and UO_2063 (O_2063,N_19923,N_19881);
nor UO_2064 (O_2064,N_19857,N_19851);
or UO_2065 (O_2065,N_19765,N_19957);
xnor UO_2066 (O_2066,N_19805,N_19980);
xor UO_2067 (O_2067,N_19881,N_19994);
or UO_2068 (O_2068,N_19996,N_19768);
or UO_2069 (O_2069,N_19801,N_19843);
nor UO_2070 (O_2070,N_19860,N_19913);
or UO_2071 (O_2071,N_19867,N_19926);
nor UO_2072 (O_2072,N_19934,N_19968);
xor UO_2073 (O_2073,N_19953,N_19942);
xnor UO_2074 (O_2074,N_19794,N_19900);
nand UO_2075 (O_2075,N_19829,N_19985);
nand UO_2076 (O_2076,N_19926,N_19928);
or UO_2077 (O_2077,N_19872,N_19822);
and UO_2078 (O_2078,N_19783,N_19970);
or UO_2079 (O_2079,N_19885,N_19968);
xnor UO_2080 (O_2080,N_19936,N_19916);
nor UO_2081 (O_2081,N_19835,N_19914);
nor UO_2082 (O_2082,N_19892,N_19780);
nor UO_2083 (O_2083,N_19812,N_19821);
xnor UO_2084 (O_2084,N_19751,N_19904);
nand UO_2085 (O_2085,N_19917,N_19790);
or UO_2086 (O_2086,N_19881,N_19978);
xnor UO_2087 (O_2087,N_19930,N_19910);
nor UO_2088 (O_2088,N_19786,N_19808);
nand UO_2089 (O_2089,N_19946,N_19960);
nand UO_2090 (O_2090,N_19782,N_19750);
or UO_2091 (O_2091,N_19841,N_19778);
and UO_2092 (O_2092,N_19875,N_19969);
xnor UO_2093 (O_2093,N_19856,N_19882);
xnor UO_2094 (O_2094,N_19858,N_19933);
and UO_2095 (O_2095,N_19777,N_19873);
xnor UO_2096 (O_2096,N_19850,N_19853);
nand UO_2097 (O_2097,N_19929,N_19952);
nor UO_2098 (O_2098,N_19797,N_19963);
and UO_2099 (O_2099,N_19885,N_19810);
and UO_2100 (O_2100,N_19940,N_19792);
xnor UO_2101 (O_2101,N_19789,N_19794);
nand UO_2102 (O_2102,N_19854,N_19917);
and UO_2103 (O_2103,N_19882,N_19976);
nand UO_2104 (O_2104,N_19940,N_19879);
nor UO_2105 (O_2105,N_19791,N_19766);
nor UO_2106 (O_2106,N_19836,N_19889);
nor UO_2107 (O_2107,N_19960,N_19847);
nand UO_2108 (O_2108,N_19840,N_19866);
nand UO_2109 (O_2109,N_19921,N_19966);
nor UO_2110 (O_2110,N_19885,N_19779);
nand UO_2111 (O_2111,N_19816,N_19963);
nand UO_2112 (O_2112,N_19786,N_19919);
and UO_2113 (O_2113,N_19760,N_19881);
xnor UO_2114 (O_2114,N_19922,N_19788);
or UO_2115 (O_2115,N_19938,N_19893);
and UO_2116 (O_2116,N_19848,N_19871);
and UO_2117 (O_2117,N_19842,N_19989);
nand UO_2118 (O_2118,N_19995,N_19798);
or UO_2119 (O_2119,N_19924,N_19811);
xor UO_2120 (O_2120,N_19827,N_19798);
and UO_2121 (O_2121,N_19774,N_19833);
xor UO_2122 (O_2122,N_19947,N_19796);
and UO_2123 (O_2123,N_19773,N_19976);
nor UO_2124 (O_2124,N_19969,N_19771);
nand UO_2125 (O_2125,N_19861,N_19769);
nand UO_2126 (O_2126,N_19927,N_19893);
xnor UO_2127 (O_2127,N_19862,N_19980);
nor UO_2128 (O_2128,N_19875,N_19864);
or UO_2129 (O_2129,N_19935,N_19942);
nand UO_2130 (O_2130,N_19991,N_19761);
or UO_2131 (O_2131,N_19912,N_19953);
or UO_2132 (O_2132,N_19936,N_19796);
nand UO_2133 (O_2133,N_19888,N_19935);
or UO_2134 (O_2134,N_19771,N_19909);
nor UO_2135 (O_2135,N_19872,N_19787);
xor UO_2136 (O_2136,N_19760,N_19985);
or UO_2137 (O_2137,N_19796,N_19895);
or UO_2138 (O_2138,N_19910,N_19987);
and UO_2139 (O_2139,N_19758,N_19801);
nor UO_2140 (O_2140,N_19797,N_19976);
nor UO_2141 (O_2141,N_19831,N_19987);
nand UO_2142 (O_2142,N_19898,N_19884);
nand UO_2143 (O_2143,N_19950,N_19997);
or UO_2144 (O_2144,N_19919,N_19909);
or UO_2145 (O_2145,N_19841,N_19752);
nand UO_2146 (O_2146,N_19763,N_19818);
nand UO_2147 (O_2147,N_19842,N_19769);
nand UO_2148 (O_2148,N_19857,N_19858);
nor UO_2149 (O_2149,N_19759,N_19780);
xnor UO_2150 (O_2150,N_19773,N_19930);
nand UO_2151 (O_2151,N_19871,N_19945);
or UO_2152 (O_2152,N_19865,N_19807);
nor UO_2153 (O_2153,N_19871,N_19880);
and UO_2154 (O_2154,N_19944,N_19816);
nand UO_2155 (O_2155,N_19994,N_19757);
or UO_2156 (O_2156,N_19919,N_19985);
nor UO_2157 (O_2157,N_19750,N_19966);
nand UO_2158 (O_2158,N_19887,N_19960);
xor UO_2159 (O_2159,N_19877,N_19790);
nor UO_2160 (O_2160,N_19904,N_19782);
xor UO_2161 (O_2161,N_19982,N_19895);
nand UO_2162 (O_2162,N_19858,N_19892);
nand UO_2163 (O_2163,N_19938,N_19832);
nand UO_2164 (O_2164,N_19962,N_19839);
and UO_2165 (O_2165,N_19832,N_19822);
nand UO_2166 (O_2166,N_19983,N_19917);
xnor UO_2167 (O_2167,N_19775,N_19879);
xor UO_2168 (O_2168,N_19945,N_19882);
nand UO_2169 (O_2169,N_19949,N_19929);
nand UO_2170 (O_2170,N_19834,N_19782);
nor UO_2171 (O_2171,N_19770,N_19867);
and UO_2172 (O_2172,N_19952,N_19898);
xor UO_2173 (O_2173,N_19827,N_19805);
nor UO_2174 (O_2174,N_19799,N_19921);
nor UO_2175 (O_2175,N_19873,N_19753);
or UO_2176 (O_2176,N_19944,N_19829);
xor UO_2177 (O_2177,N_19892,N_19863);
xnor UO_2178 (O_2178,N_19770,N_19988);
nor UO_2179 (O_2179,N_19967,N_19868);
or UO_2180 (O_2180,N_19857,N_19757);
nor UO_2181 (O_2181,N_19849,N_19915);
nor UO_2182 (O_2182,N_19987,N_19813);
nor UO_2183 (O_2183,N_19759,N_19859);
or UO_2184 (O_2184,N_19843,N_19925);
xor UO_2185 (O_2185,N_19766,N_19995);
xnor UO_2186 (O_2186,N_19876,N_19813);
nor UO_2187 (O_2187,N_19911,N_19848);
xor UO_2188 (O_2188,N_19884,N_19997);
or UO_2189 (O_2189,N_19773,N_19854);
xor UO_2190 (O_2190,N_19886,N_19768);
xnor UO_2191 (O_2191,N_19823,N_19787);
xnor UO_2192 (O_2192,N_19910,N_19774);
and UO_2193 (O_2193,N_19878,N_19968);
and UO_2194 (O_2194,N_19831,N_19889);
or UO_2195 (O_2195,N_19923,N_19819);
xor UO_2196 (O_2196,N_19823,N_19808);
xnor UO_2197 (O_2197,N_19809,N_19832);
or UO_2198 (O_2198,N_19769,N_19889);
nor UO_2199 (O_2199,N_19979,N_19945);
nor UO_2200 (O_2200,N_19915,N_19861);
xor UO_2201 (O_2201,N_19824,N_19862);
or UO_2202 (O_2202,N_19780,N_19857);
and UO_2203 (O_2203,N_19852,N_19939);
nand UO_2204 (O_2204,N_19972,N_19984);
nand UO_2205 (O_2205,N_19852,N_19901);
nor UO_2206 (O_2206,N_19877,N_19984);
and UO_2207 (O_2207,N_19809,N_19792);
and UO_2208 (O_2208,N_19784,N_19792);
nor UO_2209 (O_2209,N_19771,N_19900);
and UO_2210 (O_2210,N_19977,N_19941);
and UO_2211 (O_2211,N_19965,N_19874);
and UO_2212 (O_2212,N_19817,N_19901);
nor UO_2213 (O_2213,N_19935,N_19854);
and UO_2214 (O_2214,N_19860,N_19944);
and UO_2215 (O_2215,N_19898,N_19792);
nand UO_2216 (O_2216,N_19775,N_19829);
nand UO_2217 (O_2217,N_19781,N_19982);
nor UO_2218 (O_2218,N_19839,N_19976);
nand UO_2219 (O_2219,N_19927,N_19900);
xnor UO_2220 (O_2220,N_19858,N_19959);
and UO_2221 (O_2221,N_19869,N_19898);
or UO_2222 (O_2222,N_19982,N_19751);
xnor UO_2223 (O_2223,N_19934,N_19793);
and UO_2224 (O_2224,N_19867,N_19773);
or UO_2225 (O_2225,N_19845,N_19954);
and UO_2226 (O_2226,N_19771,N_19890);
nand UO_2227 (O_2227,N_19924,N_19800);
xnor UO_2228 (O_2228,N_19760,N_19960);
or UO_2229 (O_2229,N_19838,N_19778);
nand UO_2230 (O_2230,N_19915,N_19815);
and UO_2231 (O_2231,N_19912,N_19914);
nor UO_2232 (O_2232,N_19995,N_19819);
or UO_2233 (O_2233,N_19933,N_19852);
nand UO_2234 (O_2234,N_19808,N_19844);
nor UO_2235 (O_2235,N_19836,N_19825);
xnor UO_2236 (O_2236,N_19758,N_19852);
xor UO_2237 (O_2237,N_19953,N_19970);
and UO_2238 (O_2238,N_19830,N_19948);
xnor UO_2239 (O_2239,N_19917,N_19925);
xnor UO_2240 (O_2240,N_19823,N_19909);
and UO_2241 (O_2241,N_19996,N_19843);
and UO_2242 (O_2242,N_19981,N_19817);
nand UO_2243 (O_2243,N_19812,N_19975);
xnor UO_2244 (O_2244,N_19953,N_19779);
nand UO_2245 (O_2245,N_19918,N_19863);
or UO_2246 (O_2246,N_19909,N_19762);
xnor UO_2247 (O_2247,N_19897,N_19974);
nand UO_2248 (O_2248,N_19891,N_19827);
or UO_2249 (O_2249,N_19918,N_19979);
xnor UO_2250 (O_2250,N_19885,N_19970);
or UO_2251 (O_2251,N_19790,N_19900);
or UO_2252 (O_2252,N_19825,N_19806);
xor UO_2253 (O_2253,N_19872,N_19981);
and UO_2254 (O_2254,N_19996,N_19787);
xnor UO_2255 (O_2255,N_19895,N_19933);
nand UO_2256 (O_2256,N_19842,N_19771);
nor UO_2257 (O_2257,N_19877,N_19926);
nand UO_2258 (O_2258,N_19960,N_19977);
nor UO_2259 (O_2259,N_19982,N_19800);
xor UO_2260 (O_2260,N_19946,N_19826);
nor UO_2261 (O_2261,N_19830,N_19997);
nor UO_2262 (O_2262,N_19871,N_19920);
nor UO_2263 (O_2263,N_19751,N_19870);
nand UO_2264 (O_2264,N_19886,N_19898);
nor UO_2265 (O_2265,N_19858,N_19908);
xnor UO_2266 (O_2266,N_19867,N_19830);
xnor UO_2267 (O_2267,N_19801,N_19990);
nor UO_2268 (O_2268,N_19865,N_19919);
nor UO_2269 (O_2269,N_19830,N_19896);
and UO_2270 (O_2270,N_19826,N_19863);
nand UO_2271 (O_2271,N_19953,N_19767);
nand UO_2272 (O_2272,N_19868,N_19750);
and UO_2273 (O_2273,N_19975,N_19910);
nor UO_2274 (O_2274,N_19968,N_19856);
nor UO_2275 (O_2275,N_19799,N_19854);
xor UO_2276 (O_2276,N_19932,N_19943);
and UO_2277 (O_2277,N_19797,N_19979);
or UO_2278 (O_2278,N_19812,N_19757);
and UO_2279 (O_2279,N_19904,N_19900);
nand UO_2280 (O_2280,N_19864,N_19889);
and UO_2281 (O_2281,N_19798,N_19843);
xor UO_2282 (O_2282,N_19860,N_19851);
nand UO_2283 (O_2283,N_19883,N_19912);
xnor UO_2284 (O_2284,N_19854,N_19921);
and UO_2285 (O_2285,N_19766,N_19972);
or UO_2286 (O_2286,N_19762,N_19912);
or UO_2287 (O_2287,N_19841,N_19843);
and UO_2288 (O_2288,N_19922,N_19797);
nand UO_2289 (O_2289,N_19844,N_19948);
or UO_2290 (O_2290,N_19932,N_19808);
nand UO_2291 (O_2291,N_19800,N_19901);
and UO_2292 (O_2292,N_19984,N_19941);
or UO_2293 (O_2293,N_19808,N_19805);
nor UO_2294 (O_2294,N_19840,N_19838);
or UO_2295 (O_2295,N_19793,N_19920);
xor UO_2296 (O_2296,N_19991,N_19932);
or UO_2297 (O_2297,N_19957,N_19901);
nand UO_2298 (O_2298,N_19869,N_19846);
nand UO_2299 (O_2299,N_19765,N_19929);
xor UO_2300 (O_2300,N_19755,N_19901);
nand UO_2301 (O_2301,N_19888,N_19986);
and UO_2302 (O_2302,N_19923,N_19831);
nand UO_2303 (O_2303,N_19981,N_19889);
or UO_2304 (O_2304,N_19773,N_19902);
and UO_2305 (O_2305,N_19995,N_19833);
nor UO_2306 (O_2306,N_19931,N_19881);
and UO_2307 (O_2307,N_19913,N_19874);
and UO_2308 (O_2308,N_19797,N_19849);
nor UO_2309 (O_2309,N_19907,N_19932);
xnor UO_2310 (O_2310,N_19987,N_19933);
or UO_2311 (O_2311,N_19750,N_19960);
nand UO_2312 (O_2312,N_19815,N_19777);
or UO_2313 (O_2313,N_19996,N_19802);
or UO_2314 (O_2314,N_19816,N_19865);
xor UO_2315 (O_2315,N_19901,N_19793);
and UO_2316 (O_2316,N_19926,N_19779);
and UO_2317 (O_2317,N_19931,N_19769);
nor UO_2318 (O_2318,N_19845,N_19959);
and UO_2319 (O_2319,N_19753,N_19781);
nand UO_2320 (O_2320,N_19850,N_19998);
xor UO_2321 (O_2321,N_19832,N_19860);
or UO_2322 (O_2322,N_19942,N_19927);
or UO_2323 (O_2323,N_19887,N_19924);
xnor UO_2324 (O_2324,N_19868,N_19838);
xor UO_2325 (O_2325,N_19934,N_19884);
xor UO_2326 (O_2326,N_19896,N_19871);
and UO_2327 (O_2327,N_19959,N_19961);
xnor UO_2328 (O_2328,N_19996,N_19792);
or UO_2329 (O_2329,N_19948,N_19852);
and UO_2330 (O_2330,N_19873,N_19911);
or UO_2331 (O_2331,N_19955,N_19942);
or UO_2332 (O_2332,N_19949,N_19892);
and UO_2333 (O_2333,N_19928,N_19980);
xor UO_2334 (O_2334,N_19985,N_19890);
nor UO_2335 (O_2335,N_19878,N_19753);
or UO_2336 (O_2336,N_19806,N_19810);
or UO_2337 (O_2337,N_19816,N_19846);
or UO_2338 (O_2338,N_19888,N_19805);
xor UO_2339 (O_2339,N_19984,N_19886);
nand UO_2340 (O_2340,N_19893,N_19822);
and UO_2341 (O_2341,N_19809,N_19840);
xor UO_2342 (O_2342,N_19803,N_19908);
or UO_2343 (O_2343,N_19814,N_19905);
nand UO_2344 (O_2344,N_19985,N_19937);
or UO_2345 (O_2345,N_19901,N_19779);
and UO_2346 (O_2346,N_19861,N_19763);
or UO_2347 (O_2347,N_19901,N_19821);
and UO_2348 (O_2348,N_19952,N_19961);
nand UO_2349 (O_2349,N_19951,N_19775);
xnor UO_2350 (O_2350,N_19959,N_19859);
or UO_2351 (O_2351,N_19985,N_19864);
nor UO_2352 (O_2352,N_19901,N_19759);
and UO_2353 (O_2353,N_19958,N_19835);
or UO_2354 (O_2354,N_19884,N_19844);
or UO_2355 (O_2355,N_19825,N_19992);
xnor UO_2356 (O_2356,N_19899,N_19996);
xor UO_2357 (O_2357,N_19862,N_19932);
nor UO_2358 (O_2358,N_19783,N_19916);
and UO_2359 (O_2359,N_19916,N_19880);
xnor UO_2360 (O_2360,N_19858,N_19997);
nor UO_2361 (O_2361,N_19986,N_19905);
and UO_2362 (O_2362,N_19867,N_19878);
xor UO_2363 (O_2363,N_19952,N_19990);
xnor UO_2364 (O_2364,N_19764,N_19883);
xor UO_2365 (O_2365,N_19972,N_19914);
and UO_2366 (O_2366,N_19897,N_19960);
and UO_2367 (O_2367,N_19843,N_19866);
or UO_2368 (O_2368,N_19955,N_19758);
and UO_2369 (O_2369,N_19820,N_19928);
nor UO_2370 (O_2370,N_19842,N_19857);
nand UO_2371 (O_2371,N_19848,N_19993);
nand UO_2372 (O_2372,N_19901,N_19876);
nor UO_2373 (O_2373,N_19834,N_19879);
nor UO_2374 (O_2374,N_19844,N_19788);
xnor UO_2375 (O_2375,N_19924,N_19956);
and UO_2376 (O_2376,N_19880,N_19848);
nand UO_2377 (O_2377,N_19839,N_19864);
nor UO_2378 (O_2378,N_19826,N_19905);
or UO_2379 (O_2379,N_19894,N_19774);
nor UO_2380 (O_2380,N_19808,N_19756);
xnor UO_2381 (O_2381,N_19835,N_19968);
nor UO_2382 (O_2382,N_19924,N_19965);
nor UO_2383 (O_2383,N_19794,N_19759);
nand UO_2384 (O_2384,N_19777,N_19850);
or UO_2385 (O_2385,N_19977,N_19963);
nor UO_2386 (O_2386,N_19766,N_19804);
or UO_2387 (O_2387,N_19780,N_19753);
nor UO_2388 (O_2388,N_19917,N_19907);
or UO_2389 (O_2389,N_19857,N_19927);
or UO_2390 (O_2390,N_19869,N_19788);
or UO_2391 (O_2391,N_19952,N_19921);
and UO_2392 (O_2392,N_19764,N_19898);
or UO_2393 (O_2393,N_19904,N_19859);
nand UO_2394 (O_2394,N_19949,N_19937);
or UO_2395 (O_2395,N_19961,N_19782);
and UO_2396 (O_2396,N_19834,N_19828);
xor UO_2397 (O_2397,N_19956,N_19874);
nor UO_2398 (O_2398,N_19836,N_19861);
and UO_2399 (O_2399,N_19842,N_19924);
and UO_2400 (O_2400,N_19788,N_19778);
xnor UO_2401 (O_2401,N_19998,N_19969);
and UO_2402 (O_2402,N_19977,N_19975);
nor UO_2403 (O_2403,N_19792,N_19861);
nor UO_2404 (O_2404,N_19912,N_19819);
and UO_2405 (O_2405,N_19844,N_19830);
xnor UO_2406 (O_2406,N_19955,N_19753);
nand UO_2407 (O_2407,N_19821,N_19986);
nor UO_2408 (O_2408,N_19983,N_19817);
or UO_2409 (O_2409,N_19890,N_19813);
xnor UO_2410 (O_2410,N_19870,N_19768);
and UO_2411 (O_2411,N_19854,N_19785);
nor UO_2412 (O_2412,N_19857,N_19841);
nand UO_2413 (O_2413,N_19895,N_19913);
or UO_2414 (O_2414,N_19904,N_19842);
xor UO_2415 (O_2415,N_19931,N_19944);
and UO_2416 (O_2416,N_19895,N_19840);
xnor UO_2417 (O_2417,N_19922,N_19866);
or UO_2418 (O_2418,N_19859,N_19969);
nor UO_2419 (O_2419,N_19964,N_19853);
xor UO_2420 (O_2420,N_19817,N_19822);
or UO_2421 (O_2421,N_19889,N_19957);
or UO_2422 (O_2422,N_19878,N_19773);
nand UO_2423 (O_2423,N_19878,N_19834);
or UO_2424 (O_2424,N_19952,N_19819);
nand UO_2425 (O_2425,N_19992,N_19979);
or UO_2426 (O_2426,N_19809,N_19761);
or UO_2427 (O_2427,N_19880,N_19903);
nand UO_2428 (O_2428,N_19916,N_19926);
or UO_2429 (O_2429,N_19751,N_19762);
and UO_2430 (O_2430,N_19987,N_19923);
and UO_2431 (O_2431,N_19904,N_19789);
nor UO_2432 (O_2432,N_19816,N_19918);
xor UO_2433 (O_2433,N_19945,N_19896);
or UO_2434 (O_2434,N_19975,N_19888);
and UO_2435 (O_2435,N_19994,N_19802);
and UO_2436 (O_2436,N_19975,N_19873);
nand UO_2437 (O_2437,N_19840,N_19946);
and UO_2438 (O_2438,N_19756,N_19757);
xnor UO_2439 (O_2439,N_19868,N_19799);
or UO_2440 (O_2440,N_19763,N_19885);
or UO_2441 (O_2441,N_19967,N_19819);
xor UO_2442 (O_2442,N_19800,N_19942);
nand UO_2443 (O_2443,N_19808,N_19898);
nor UO_2444 (O_2444,N_19788,N_19852);
and UO_2445 (O_2445,N_19862,N_19849);
or UO_2446 (O_2446,N_19921,N_19998);
and UO_2447 (O_2447,N_19762,N_19986);
xor UO_2448 (O_2448,N_19830,N_19933);
nor UO_2449 (O_2449,N_19921,N_19946);
nand UO_2450 (O_2450,N_19893,N_19926);
xor UO_2451 (O_2451,N_19887,N_19864);
nand UO_2452 (O_2452,N_19772,N_19879);
or UO_2453 (O_2453,N_19910,N_19979);
xnor UO_2454 (O_2454,N_19776,N_19891);
xnor UO_2455 (O_2455,N_19881,N_19960);
xnor UO_2456 (O_2456,N_19983,N_19831);
and UO_2457 (O_2457,N_19839,N_19902);
nand UO_2458 (O_2458,N_19980,N_19859);
or UO_2459 (O_2459,N_19965,N_19756);
or UO_2460 (O_2460,N_19794,N_19841);
and UO_2461 (O_2461,N_19836,N_19826);
or UO_2462 (O_2462,N_19879,N_19862);
nor UO_2463 (O_2463,N_19820,N_19817);
or UO_2464 (O_2464,N_19875,N_19968);
and UO_2465 (O_2465,N_19980,N_19962);
nand UO_2466 (O_2466,N_19811,N_19912);
and UO_2467 (O_2467,N_19883,N_19916);
or UO_2468 (O_2468,N_19843,N_19810);
and UO_2469 (O_2469,N_19771,N_19861);
and UO_2470 (O_2470,N_19957,N_19952);
and UO_2471 (O_2471,N_19825,N_19819);
and UO_2472 (O_2472,N_19952,N_19960);
and UO_2473 (O_2473,N_19929,N_19993);
nor UO_2474 (O_2474,N_19871,N_19868);
xnor UO_2475 (O_2475,N_19851,N_19987);
and UO_2476 (O_2476,N_19849,N_19993);
and UO_2477 (O_2477,N_19908,N_19825);
xnor UO_2478 (O_2478,N_19756,N_19893);
nand UO_2479 (O_2479,N_19806,N_19996);
nor UO_2480 (O_2480,N_19865,N_19889);
and UO_2481 (O_2481,N_19935,N_19993);
nand UO_2482 (O_2482,N_19926,N_19874);
or UO_2483 (O_2483,N_19844,N_19943);
nor UO_2484 (O_2484,N_19770,N_19755);
nand UO_2485 (O_2485,N_19794,N_19936);
or UO_2486 (O_2486,N_19802,N_19805);
and UO_2487 (O_2487,N_19942,N_19855);
nand UO_2488 (O_2488,N_19842,N_19844);
nor UO_2489 (O_2489,N_19966,N_19899);
and UO_2490 (O_2490,N_19976,N_19956);
nand UO_2491 (O_2491,N_19903,N_19852);
xnor UO_2492 (O_2492,N_19977,N_19789);
nand UO_2493 (O_2493,N_19846,N_19918);
or UO_2494 (O_2494,N_19942,N_19973);
xnor UO_2495 (O_2495,N_19859,N_19966);
and UO_2496 (O_2496,N_19850,N_19861);
xor UO_2497 (O_2497,N_19789,N_19970);
or UO_2498 (O_2498,N_19796,N_19869);
xnor UO_2499 (O_2499,N_19967,N_19895);
endmodule