module basic_500_3000_500_6_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_411,In_317);
and U1 (N_1,In_446,In_104);
or U2 (N_2,In_266,In_129);
or U3 (N_3,In_54,In_123);
nand U4 (N_4,In_73,In_227);
nand U5 (N_5,In_118,In_16);
or U6 (N_6,In_346,In_109);
nor U7 (N_7,In_248,In_238);
and U8 (N_8,In_311,In_42);
and U9 (N_9,In_468,In_30);
nor U10 (N_10,In_98,In_170);
nand U11 (N_11,In_82,In_377);
or U12 (N_12,In_190,In_243);
nor U13 (N_13,In_172,In_130);
nor U14 (N_14,In_110,In_239);
and U15 (N_15,In_309,In_384);
xor U16 (N_16,In_473,In_20);
or U17 (N_17,In_373,In_162);
and U18 (N_18,In_114,In_58);
or U19 (N_19,In_481,In_32);
nand U20 (N_20,In_440,In_462);
or U21 (N_21,In_211,In_43);
and U22 (N_22,In_390,In_307);
nor U23 (N_23,In_124,In_93);
or U24 (N_24,In_328,In_482);
nor U25 (N_25,In_35,In_256);
or U26 (N_26,In_220,In_92);
xor U27 (N_27,In_278,In_204);
or U28 (N_28,In_269,In_194);
nor U29 (N_29,In_492,In_436);
xor U30 (N_30,In_324,In_378);
nor U31 (N_31,In_415,In_60);
or U32 (N_32,In_210,In_424);
and U33 (N_33,In_437,In_363);
or U34 (N_34,In_380,In_300);
nand U35 (N_35,In_120,In_361);
or U36 (N_36,In_155,In_267);
or U37 (N_37,In_460,In_27);
or U38 (N_38,In_394,In_439);
nand U39 (N_39,In_165,In_486);
xor U40 (N_40,In_87,In_485);
and U41 (N_41,In_405,In_251);
nand U42 (N_42,In_96,In_416);
xnor U43 (N_43,In_398,In_188);
nor U44 (N_44,In_189,In_258);
nor U45 (N_45,In_133,In_400);
or U46 (N_46,In_385,In_325);
or U47 (N_47,In_465,In_6);
or U48 (N_48,In_297,In_444);
nand U49 (N_49,In_438,In_177);
or U50 (N_50,In_55,In_15);
nand U51 (N_51,In_432,In_11);
nor U52 (N_52,In_289,In_364);
xnor U53 (N_53,In_44,In_496);
nor U54 (N_54,In_180,In_184);
nand U55 (N_55,In_4,In_223);
nor U56 (N_56,In_487,In_393);
or U57 (N_57,In_351,In_467);
nand U58 (N_58,In_339,In_260);
and U59 (N_59,In_218,In_141);
nand U60 (N_60,In_131,In_428);
xnor U61 (N_61,In_352,In_274);
or U62 (N_62,In_222,In_434);
nor U63 (N_63,In_163,In_368);
xnor U64 (N_64,In_312,In_259);
nand U65 (N_65,In_85,In_206);
nor U66 (N_66,In_75,In_216);
and U67 (N_67,In_374,In_139);
nand U68 (N_68,In_391,In_288);
nor U69 (N_69,In_335,In_302);
or U70 (N_70,In_349,In_91);
nor U71 (N_71,In_198,In_175);
and U72 (N_72,In_254,In_119);
or U73 (N_73,In_397,In_94);
and U74 (N_74,In_367,In_402);
xnor U75 (N_75,In_301,In_66);
nand U76 (N_76,In_376,In_408);
and U77 (N_77,In_217,In_145);
nand U78 (N_78,In_414,In_365);
or U79 (N_79,In_413,In_225);
or U80 (N_80,In_321,In_38);
nor U81 (N_81,In_455,In_379);
nand U82 (N_82,In_280,In_318);
nand U83 (N_83,In_423,In_137);
nor U84 (N_84,In_125,In_226);
and U85 (N_85,In_168,In_80);
or U86 (N_86,In_354,In_95);
xor U87 (N_87,In_334,In_371);
and U88 (N_88,In_375,In_24);
nor U89 (N_89,In_26,In_116);
nand U90 (N_90,In_427,In_151);
nand U91 (N_91,In_331,In_268);
nand U92 (N_92,In_138,In_315);
nand U93 (N_93,In_340,In_53);
nand U94 (N_94,In_51,In_112);
nand U95 (N_95,In_264,In_5);
nand U96 (N_96,In_186,In_196);
nand U97 (N_97,In_156,In_199);
nor U98 (N_98,In_357,In_244);
nor U99 (N_99,In_57,In_422);
nand U100 (N_100,In_111,In_341);
or U101 (N_101,In_290,In_359);
nand U102 (N_102,In_136,In_454);
nand U103 (N_103,In_452,In_466);
or U104 (N_104,In_193,In_203);
nand U105 (N_105,In_158,In_285);
nand U106 (N_106,In_355,In_291);
nor U107 (N_107,In_224,In_50);
xor U108 (N_108,In_313,In_445);
nand U109 (N_109,In_430,In_143);
nand U110 (N_110,In_208,In_67);
nor U111 (N_111,In_65,In_74);
nand U112 (N_112,In_488,In_314);
nand U113 (N_113,In_295,In_221);
and U114 (N_114,In_435,In_347);
or U115 (N_115,In_242,In_276);
nand U116 (N_116,In_306,In_237);
nor U117 (N_117,In_146,In_490);
nand U118 (N_118,In_447,In_261);
and U119 (N_119,In_212,In_426);
nand U120 (N_120,In_76,In_161);
or U121 (N_121,In_240,In_275);
nand U122 (N_122,In_78,In_395);
xor U123 (N_123,In_420,In_272);
or U124 (N_124,In_499,In_353);
nand U125 (N_125,In_21,In_281);
nand U126 (N_126,In_322,In_279);
nor U127 (N_127,In_250,In_2);
xnor U128 (N_128,In_149,In_388);
nand U129 (N_129,In_182,In_456);
and U130 (N_130,In_25,In_326);
or U131 (N_131,In_484,In_294);
nand U132 (N_132,In_8,In_336);
nand U133 (N_133,In_106,In_386);
nor U134 (N_134,In_406,In_89);
and U135 (N_135,In_201,In_305);
nand U136 (N_136,In_476,In_333);
nand U137 (N_137,In_234,In_407);
nand U138 (N_138,In_19,In_152);
nor U139 (N_139,In_22,In_40);
and U140 (N_140,In_134,In_122);
nor U141 (N_141,In_419,In_231);
or U142 (N_142,In_296,In_113);
nand U143 (N_143,In_257,In_270);
nor U144 (N_144,In_245,In_431);
or U145 (N_145,In_115,In_381);
xor U146 (N_146,In_404,In_86);
nor U147 (N_147,In_392,In_195);
and U148 (N_148,In_358,In_255);
and U149 (N_149,In_207,In_62);
and U150 (N_150,In_327,In_167);
nand U151 (N_151,In_483,In_160);
or U152 (N_152,In_107,In_63);
or U153 (N_153,In_39,In_173);
nand U154 (N_154,In_34,In_29);
nand U155 (N_155,In_79,In_215);
or U156 (N_156,In_299,In_448);
nand U157 (N_157,In_214,In_491);
nor U158 (N_158,In_37,In_253);
and U159 (N_159,In_200,In_101);
and U160 (N_160,In_304,In_479);
or U161 (N_161,In_83,In_497);
or U162 (N_162,In_219,In_425);
and U163 (N_163,In_362,In_442);
nand U164 (N_164,In_443,In_310);
nor U165 (N_165,In_337,In_81);
or U166 (N_166,In_97,In_399);
or U167 (N_167,In_382,In_401);
or U168 (N_168,In_247,In_178);
or U169 (N_169,In_117,In_265);
xor U170 (N_170,In_495,In_417);
and U171 (N_171,In_235,In_232);
or U172 (N_172,In_478,In_451);
nand U173 (N_173,In_153,In_45);
nor U174 (N_174,In_99,In_480);
nor U175 (N_175,In_142,In_360);
or U176 (N_176,In_271,In_458);
nor U177 (N_177,In_418,In_56);
and U178 (N_178,In_179,In_3);
nand U179 (N_179,In_286,In_68);
nand U180 (N_180,In_100,In_103);
and U181 (N_181,In_409,In_154);
xor U182 (N_182,In_69,In_148);
and U183 (N_183,In_52,In_472);
nand U184 (N_184,In_370,In_213);
nor U185 (N_185,In_150,In_433);
xor U186 (N_186,In_36,In_412);
nand U187 (N_187,In_429,In_41);
nor U188 (N_188,In_246,In_183);
and U189 (N_189,In_157,In_338);
nor U190 (N_190,In_469,In_230);
and U191 (N_191,In_229,In_498);
and U192 (N_192,In_46,In_228);
or U193 (N_193,In_369,In_33);
xor U194 (N_194,In_461,In_263);
nand U195 (N_195,In_166,In_12);
nand U196 (N_196,In_77,In_298);
nor U197 (N_197,In_316,In_459);
nor U198 (N_198,In_197,In_7);
or U199 (N_199,In_132,In_241);
xor U200 (N_200,In_185,In_273);
and U201 (N_201,In_320,In_372);
or U202 (N_202,In_323,In_171);
nor U203 (N_203,In_31,In_453);
and U204 (N_204,In_292,In_48);
xor U205 (N_205,In_9,In_348);
and U206 (N_206,In_191,In_205);
nor U207 (N_207,In_277,In_90);
nor U208 (N_208,In_47,In_421);
nor U209 (N_209,In_61,In_174);
nor U210 (N_210,In_463,In_236);
and U211 (N_211,In_303,In_252);
nor U212 (N_212,In_383,In_181);
nand U213 (N_213,In_159,In_449);
and U214 (N_214,In_342,In_147);
or U215 (N_215,In_282,In_88);
and U216 (N_216,In_329,In_344);
or U217 (N_217,In_441,In_64);
and U218 (N_218,In_350,In_283);
or U219 (N_219,In_319,In_450);
nor U220 (N_220,In_493,In_471);
nor U221 (N_221,In_49,In_284);
or U222 (N_222,In_10,In_262);
and U223 (N_223,In_0,In_387);
nand U224 (N_224,In_477,In_192);
or U225 (N_225,In_356,In_489);
xnor U226 (N_226,In_71,In_202);
nor U227 (N_227,In_14,In_403);
and U228 (N_228,In_293,In_135);
nand U229 (N_229,In_164,In_70);
and U230 (N_230,In_470,In_249);
or U231 (N_231,In_72,In_18);
nor U232 (N_232,In_287,In_345);
nor U233 (N_233,In_474,In_187);
or U234 (N_234,In_366,In_102);
xnor U235 (N_235,In_457,In_308);
nand U236 (N_236,In_121,In_105);
and U237 (N_237,In_84,In_59);
and U238 (N_238,In_330,In_126);
nand U239 (N_239,In_464,In_140);
or U240 (N_240,In_396,In_17);
nand U241 (N_241,In_108,In_209);
nand U242 (N_242,In_332,In_1);
and U243 (N_243,In_343,In_28);
nand U244 (N_244,In_233,In_144);
nand U245 (N_245,In_23,In_176);
and U246 (N_246,In_127,In_494);
nor U247 (N_247,In_128,In_13);
and U248 (N_248,In_410,In_475);
or U249 (N_249,In_389,In_169);
xor U250 (N_250,In_388,In_30);
or U251 (N_251,In_124,In_320);
nand U252 (N_252,In_452,In_110);
xnor U253 (N_253,In_87,In_247);
or U254 (N_254,In_310,In_29);
or U255 (N_255,In_455,In_302);
nor U256 (N_256,In_3,In_89);
nand U257 (N_257,In_312,In_61);
nand U258 (N_258,In_131,In_263);
nor U259 (N_259,In_377,In_424);
nor U260 (N_260,In_225,In_269);
nor U261 (N_261,In_39,In_52);
or U262 (N_262,In_392,In_342);
and U263 (N_263,In_269,In_493);
or U264 (N_264,In_454,In_55);
nand U265 (N_265,In_293,In_48);
or U266 (N_266,In_281,In_473);
nand U267 (N_267,In_405,In_58);
nand U268 (N_268,In_35,In_32);
or U269 (N_269,In_52,In_251);
and U270 (N_270,In_21,In_172);
nor U271 (N_271,In_242,In_370);
and U272 (N_272,In_71,In_62);
nand U273 (N_273,In_51,In_65);
nand U274 (N_274,In_227,In_75);
nor U275 (N_275,In_277,In_175);
and U276 (N_276,In_258,In_205);
nand U277 (N_277,In_341,In_312);
or U278 (N_278,In_139,In_292);
nor U279 (N_279,In_398,In_88);
and U280 (N_280,In_433,In_158);
nand U281 (N_281,In_381,In_475);
and U282 (N_282,In_461,In_67);
and U283 (N_283,In_114,In_328);
nor U284 (N_284,In_439,In_440);
xor U285 (N_285,In_305,In_158);
nand U286 (N_286,In_288,In_82);
or U287 (N_287,In_269,In_169);
nor U288 (N_288,In_15,In_166);
and U289 (N_289,In_246,In_231);
or U290 (N_290,In_432,In_167);
nand U291 (N_291,In_96,In_474);
or U292 (N_292,In_416,In_173);
or U293 (N_293,In_171,In_216);
or U294 (N_294,In_169,In_64);
or U295 (N_295,In_425,In_74);
nor U296 (N_296,In_137,In_494);
xnor U297 (N_297,In_6,In_241);
or U298 (N_298,In_395,In_155);
nand U299 (N_299,In_205,In_161);
xnor U300 (N_300,In_231,In_289);
nand U301 (N_301,In_308,In_490);
nor U302 (N_302,In_102,In_304);
nor U303 (N_303,In_163,In_408);
nand U304 (N_304,In_265,In_191);
nand U305 (N_305,In_24,In_153);
or U306 (N_306,In_331,In_36);
nand U307 (N_307,In_86,In_443);
nor U308 (N_308,In_350,In_395);
nor U309 (N_309,In_419,In_172);
and U310 (N_310,In_62,In_113);
and U311 (N_311,In_431,In_6);
or U312 (N_312,In_345,In_10);
nand U313 (N_313,In_301,In_78);
xor U314 (N_314,In_72,In_54);
and U315 (N_315,In_60,In_328);
and U316 (N_316,In_418,In_41);
or U317 (N_317,In_284,In_321);
or U318 (N_318,In_106,In_176);
nor U319 (N_319,In_13,In_131);
nor U320 (N_320,In_244,In_455);
nand U321 (N_321,In_420,In_390);
nor U322 (N_322,In_48,In_91);
nor U323 (N_323,In_431,In_37);
and U324 (N_324,In_411,In_193);
xnor U325 (N_325,In_272,In_494);
or U326 (N_326,In_149,In_145);
and U327 (N_327,In_1,In_437);
or U328 (N_328,In_157,In_347);
or U329 (N_329,In_154,In_12);
nand U330 (N_330,In_48,In_402);
xnor U331 (N_331,In_282,In_30);
nor U332 (N_332,In_98,In_253);
nand U333 (N_333,In_373,In_17);
and U334 (N_334,In_342,In_129);
and U335 (N_335,In_394,In_213);
or U336 (N_336,In_446,In_441);
and U337 (N_337,In_498,In_485);
nor U338 (N_338,In_331,In_398);
nor U339 (N_339,In_79,In_385);
or U340 (N_340,In_112,In_353);
or U341 (N_341,In_396,In_322);
or U342 (N_342,In_120,In_204);
nand U343 (N_343,In_416,In_334);
and U344 (N_344,In_329,In_100);
xnor U345 (N_345,In_163,In_146);
or U346 (N_346,In_24,In_274);
or U347 (N_347,In_9,In_67);
nor U348 (N_348,In_418,In_323);
nand U349 (N_349,In_482,In_286);
nand U350 (N_350,In_478,In_334);
nor U351 (N_351,In_313,In_419);
or U352 (N_352,In_50,In_325);
or U353 (N_353,In_258,In_415);
nand U354 (N_354,In_343,In_66);
nor U355 (N_355,In_354,In_383);
and U356 (N_356,In_344,In_448);
and U357 (N_357,In_41,In_260);
and U358 (N_358,In_314,In_2);
or U359 (N_359,In_380,In_179);
nor U360 (N_360,In_186,In_197);
nand U361 (N_361,In_138,In_349);
nand U362 (N_362,In_93,In_439);
or U363 (N_363,In_410,In_402);
nand U364 (N_364,In_150,In_344);
or U365 (N_365,In_183,In_214);
and U366 (N_366,In_257,In_404);
and U367 (N_367,In_113,In_327);
nor U368 (N_368,In_455,In_422);
nor U369 (N_369,In_320,In_244);
nor U370 (N_370,In_154,In_482);
nand U371 (N_371,In_251,In_397);
or U372 (N_372,In_149,In_458);
nand U373 (N_373,In_463,In_176);
or U374 (N_374,In_240,In_466);
nand U375 (N_375,In_328,In_181);
nand U376 (N_376,In_284,In_357);
nor U377 (N_377,In_81,In_96);
or U378 (N_378,In_379,In_227);
nand U379 (N_379,In_46,In_474);
and U380 (N_380,In_210,In_470);
nand U381 (N_381,In_284,In_177);
nor U382 (N_382,In_428,In_262);
nand U383 (N_383,In_182,In_118);
xor U384 (N_384,In_103,In_237);
and U385 (N_385,In_273,In_413);
nand U386 (N_386,In_105,In_252);
or U387 (N_387,In_203,In_266);
and U388 (N_388,In_108,In_366);
or U389 (N_389,In_299,In_43);
xnor U390 (N_390,In_112,In_26);
nor U391 (N_391,In_122,In_21);
nor U392 (N_392,In_15,In_121);
xor U393 (N_393,In_360,In_258);
nor U394 (N_394,In_400,In_88);
or U395 (N_395,In_400,In_99);
nand U396 (N_396,In_471,In_475);
nor U397 (N_397,In_220,In_335);
and U398 (N_398,In_57,In_488);
nand U399 (N_399,In_11,In_81);
and U400 (N_400,In_177,In_25);
and U401 (N_401,In_280,In_51);
or U402 (N_402,In_94,In_491);
nand U403 (N_403,In_0,In_86);
and U404 (N_404,In_48,In_357);
or U405 (N_405,In_434,In_48);
nor U406 (N_406,In_181,In_331);
nand U407 (N_407,In_370,In_210);
xor U408 (N_408,In_110,In_180);
and U409 (N_409,In_475,In_170);
nor U410 (N_410,In_325,In_96);
xor U411 (N_411,In_286,In_345);
and U412 (N_412,In_297,In_163);
nor U413 (N_413,In_337,In_6);
nor U414 (N_414,In_402,In_403);
xor U415 (N_415,In_314,In_136);
nand U416 (N_416,In_272,In_10);
nor U417 (N_417,In_233,In_45);
and U418 (N_418,In_473,In_471);
nand U419 (N_419,In_426,In_78);
nor U420 (N_420,In_77,In_197);
and U421 (N_421,In_418,In_184);
nand U422 (N_422,In_167,In_348);
nand U423 (N_423,In_283,In_299);
nand U424 (N_424,In_271,In_198);
or U425 (N_425,In_433,In_253);
and U426 (N_426,In_417,In_127);
or U427 (N_427,In_51,In_308);
or U428 (N_428,In_389,In_317);
nand U429 (N_429,In_345,In_299);
xnor U430 (N_430,In_301,In_312);
and U431 (N_431,In_405,In_73);
nand U432 (N_432,In_291,In_43);
or U433 (N_433,In_236,In_337);
and U434 (N_434,In_462,In_475);
nand U435 (N_435,In_313,In_91);
and U436 (N_436,In_352,In_290);
nand U437 (N_437,In_165,In_429);
and U438 (N_438,In_156,In_186);
xor U439 (N_439,In_73,In_176);
or U440 (N_440,In_123,In_232);
and U441 (N_441,In_32,In_402);
nor U442 (N_442,In_5,In_2);
nor U443 (N_443,In_247,In_383);
or U444 (N_444,In_95,In_161);
or U445 (N_445,In_327,In_283);
or U446 (N_446,In_3,In_17);
and U447 (N_447,In_213,In_153);
or U448 (N_448,In_347,In_167);
and U449 (N_449,In_6,In_139);
nand U450 (N_450,In_282,In_443);
nor U451 (N_451,In_390,In_289);
nand U452 (N_452,In_451,In_323);
xor U453 (N_453,In_297,In_183);
nand U454 (N_454,In_167,In_285);
or U455 (N_455,In_423,In_419);
nand U456 (N_456,In_379,In_392);
nand U457 (N_457,In_40,In_208);
nand U458 (N_458,In_287,In_25);
and U459 (N_459,In_141,In_339);
nor U460 (N_460,In_51,In_358);
or U461 (N_461,In_422,In_71);
nor U462 (N_462,In_388,In_220);
and U463 (N_463,In_460,In_353);
and U464 (N_464,In_127,In_77);
and U465 (N_465,In_494,In_95);
nor U466 (N_466,In_289,In_186);
nand U467 (N_467,In_165,In_164);
or U468 (N_468,In_45,In_210);
nand U469 (N_469,In_203,In_6);
or U470 (N_470,In_460,In_325);
and U471 (N_471,In_381,In_367);
or U472 (N_472,In_115,In_377);
or U473 (N_473,In_25,In_407);
or U474 (N_474,In_167,In_94);
xor U475 (N_475,In_92,In_446);
nand U476 (N_476,In_363,In_477);
or U477 (N_477,In_380,In_91);
or U478 (N_478,In_45,In_171);
and U479 (N_479,In_466,In_31);
nor U480 (N_480,In_380,In_367);
nor U481 (N_481,In_384,In_444);
and U482 (N_482,In_179,In_493);
nand U483 (N_483,In_489,In_333);
or U484 (N_484,In_410,In_318);
nor U485 (N_485,In_133,In_438);
nand U486 (N_486,In_138,In_68);
and U487 (N_487,In_310,In_95);
nor U488 (N_488,In_292,In_256);
xor U489 (N_489,In_152,In_224);
nor U490 (N_490,In_158,In_301);
nand U491 (N_491,In_350,In_330);
nand U492 (N_492,In_205,In_369);
xor U493 (N_493,In_239,In_194);
and U494 (N_494,In_490,In_59);
nand U495 (N_495,In_48,In_16);
nand U496 (N_496,In_248,In_64);
or U497 (N_497,In_207,In_286);
nand U498 (N_498,In_70,In_493);
or U499 (N_499,In_482,In_475);
nor U500 (N_500,N_305,N_261);
and U501 (N_501,N_446,N_14);
or U502 (N_502,N_189,N_490);
xnor U503 (N_503,N_70,N_416);
and U504 (N_504,N_160,N_345);
nand U505 (N_505,N_124,N_405);
or U506 (N_506,N_205,N_452);
nand U507 (N_507,N_413,N_142);
xor U508 (N_508,N_482,N_280);
and U509 (N_509,N_204,N_120);
or U510 (N_510,N_302,N_107);
nor U511 (N_511,N_87,N_323);
and U512 (N_512,N_481,N_144);
and U513 (N_513,N_118,N_194);
and U514 (N_514,N_435,N_226);
or U515 (N_515,N_95,N_136);
and U516 (N_516,N_439,N_97);
nand U517 (N_517,N_182,N_440);
and U518 (N_518,N_11,N_38);
nand U519 (N_519,N_290,N_461);
nor U520 (N_520,N_248,N_135);
nor U521 (N_521,N_187,N_495);
or U522 (N_522,N_262,N_195);
xnor U523 (N_523,N_252,N_161);
nand U524 (N_524,N_498,N_67);
xor U525 (N_525,N_377,N_78);
nor U526 (N_526,N_374,N_229);
xnor U527 (N_527,N_279,N_354);
nor U528 (N_528,N_271,N_178);
nand U529 (N_529,N_379,N_167);
or U530 (N_530,N_197,N_111);
nor U531 (N_531,N_286,N_314);
xnor U532 (N_532,N_369,N_464);
nand U533 (N_533,N_311,N_201);
nor U534 (N_534,N_433,N_214);
and U535 (N_535,N_260,N_491);
nand U536 (N_536,N_175,N_384);
nand U537 (N_537,N_173,N_174);
nor U538 (N_538,N_22,N_221);
nor U539 (N_539,N_172,N_73);
or U540 (N_540,N_497,N_283);
nor U541 (N_541,N_364,N_185);
nor U542 (N_542,N_276,N_179);
and U543 (N_543,N_6,N_465);
and U544 (N_544,N_313,N_158);
nor U545 (N_545,N_51,N_163);
and U546 (N_546,N_301,N_449);
or U547 (N_547,N_159,N_150);
nor U548 (N_548,N_391,N_59);
or U549 (N_549,N_53,N_28);
nor U550 (N_550,N_177,N_285);
nand U551 (N_551,N_406,N_386);
or U552 (N_552,N_154,N_35);
xnor U553 (N_553,N_408,N_333);
and U554 (N_554,N_141,N_196);
or U555 (N_555,N_63,N_335);
and U556 (N_556,N_259,N_147);
nor U557 (N_557,N_110,N_164);
nor U558 (N_558,N_417,N_426);
nand U559 (N_559,N_134,N_162);
nand U560 (N_560,N_18,N_102);
and U561 (N_561,N_343,N_37);
nor U562 (N_562,N_385,N_493);
nor U563 (N_563,N_460,N_48);
nand U564 (N_564,N_296,N_222);
nand U565 (N_565,N_451,N_371);
and U566 (N_566,N_100,N_176);
or U567 (N_567,N_308,N_206);
and U568 (N_568,N_93,N_103);
nor U569 (N_569,N_191,N_253);
nand U570 (N_570,N_80,N_246);
nor U571 (N_571,N_424,N_104);
nand U572 (N_572,N_232,N_436);
nor U573 (N_573,N_143,N_486);
xnor U574 (N_574,N_105,N_472);
nor U575 (N_575,N_344,N_348);
and U576 (N_576,N_122,N_133);
nand U577 (N_577,N_12,N_74);
nand U578 (N_578,N_42,N_112);
xor U579 (N_579,N_169,N_34);
or U580 (N_580,N_363,N_299);
nand U581 (N_581,N_129,N_475);
xnor U582 (N_582,N_75,N_289);
nand U583 (N_583,N_145,N_431);
or U584 (N_584,N_456,N_69);
nand U585 (N_585,N_139,N_339);
and U586 (N_586,N_485,N_390);
nand U587 (N_587,N_32,N_429);
xnor U588 (N_588,N_337,N_16);
xnor U589 (N_589,N_89,N_477);
and U590 (N_590,N_101,N_44);
nand U591 (N_591,N_395,N_284);
nand U592 (N_592,N_434,N_338);
and U593 (N_593,N_0,N_373);
xnor U594 (N_594,N_347,N_269);
or U595 (N_595,N_420,N_132);
or U596 (N_596,N_297,N_317);
nand U597 (N_597,N_396,N_309);
xor U598 (N_598,N_245,N_215);
or U599 (N_599,N_84,N_108);
or U600 (N_600,N_499,N_352);
nor U601 (N_601,N_153,N_432);
and U602 (N_602,N_423,N_488);
nor U603 (N_603,N_330,N_468);
and U604 (N_604,N_62,N_404);
or U605 (N_605,N_224,N_326);
or U606 (N_606,N_29,N_184);
nand U607 (N_607,N_457,N_106);
xor U608 (N_608,N_123,N_265);
nor U609 (N_609,N_392,N_65);
nand U610 (N_610,N_151,N_400);
nand U611 (N_611,N_471,N_180);
or U612 (N_612,N_427,N_401);
nand U613 (N_613,N_243,N_361);
or U614 (N_614,N_466,N_264);
or U615 (N_615,N_121,N_444);
and U616 (N_616,N_474,N_447);
or U617 (N_617,N_320,N_1);
nor U618 (N_618,N_362,N_298);
and U619 (N_619,N_17,N_170);
nor U620 (N_620,N_146,N_4);
or U621 (N_621,N_263,N_43);
nand U622 (N_622,N_193,N_86);
and U623 (N_623,N_186,N_99);
nor U624 (N_624,N_138,N_13);
nor U625 (N_625,N_198,N_430);
nand U626 (N_626,N_127,N_351);
nand U627 (N_627,N_119,N_480);
nor U628 (N_628,N_239,N_274);
xnor U629 (N_629,N_47,N_483);
nor U630 (N_630,N_156,N_24);
and U631 (N_631,N_249,N_98);
nor U632 (N_632,N_292,N_220);
nand U633 (N_633,N_453,N_288);
or U634 (N_634,N_428,N_56);
nor U635 (N_635,N_240,N_378);
nand U636 (N_636,N_455,N_212);
or U637 (N_637,N_210,N_46);
or U638 (N_638,N_360,N_237);
nand U639 (N_639,N_470,N_353);
nor U640 (N_640,N_188,N_322);
or U641 (N_641,N_39,N_293);
nor U642 (N_642,N_367,N_382);
nor U643 (N_643,N_61,N_402);
nor U644 (N_644,N_91,N_342);
or U645 (N_645,N_183,N_273);
xnor U646 (N_646,N_45,N_282);
or U647 (N_647,N_281,N_398);
or U648 (N_648,N_7,N_68);
nor U649 (N_649,N_376,N_437);
nand U650 (N_650,N_117,N_64);
and U651 (N_651,N_211,N_3);
and U652 (N_652,N_321,N_278);
or U653 (N_653,N_448,N_368);
or U654 (N_654,N_231,N_41);
or U655 (N_655,N_168,N_213);
nor U656 (N_656,N_409,N_40);
nor U657 (N_657,N_334,N_209);
xnor U658 (N_658,N_350,N_267);
nand U659 (N_659,N_36,N_9);
nor U660 (N_660,N_81,N_469);
nand U661 (N_661,N_90,N_393);
or U662 (N_662,N_58,N_441);
nor U663 (N_663,N_113,N_256);
nand U664 (N_664,N_438,N_203);
nand U665 (N_665,N_319,N_372);
and U666 (N_666,N_190,N_357);
nand U667 (N_667,N_359,N_30);
nor U668 (N_668,N_346,N_60);
nand U669 (N_669,N_230,N_165);
and U670 (N_670,N_83,N_463);
and U671 (N_671,N_19,N_383);
nand U672 (N_672,N_155,N_399);
and U673 (N_673,N_241,N_148);
nand U674 (N_674,N_242,N_238);
xor U675 (N_675,N_49,N_312);
and U676 (N_676,N_15,N_217);
or U677 (N_677,N_31,N_137);
or U678 (N_678,N_26,N_327);
xnor U679 (N_679,N_479,N_387);
xor U680 (N_680,N_496,N_199);
or U681 (N_681,N_459,N_307);
xor U682 (N_682,N_202,N_476);
nand U683 (N_683,N_207,N_216);
nand U684 (N_684,N_96,N_425);
nand U685 (N_685,N_336,N_76);
nand U686 (N_686,N_77,N_192);
or U687 (N_687,N_54,N_130);
nand U688 (N_688,N_380,N_421);
and U689 (N_689,N_445,N_33);
nand U690 (N_690,N_20,N_250);
and U691 (N_691,N_277,N_291);
and U692 (N_692,N_5,N_181);
nand U693 (N_693,N_244,N_478);
nand U694 (N_694,N_272,N_200);
and U695 (N_695,N_487,N_494);
nand U696 (N_696,N_275,N_266);
and U697 (N_697,N_407,N_233);
nand U698 (N_698,N_397,N_255);
and U699 (N_699,N_228,N_473);
and U700 (N_700,N_166,N_462);
or U701 (N_701,N_27,N_318);
nor U702 (N_702,N_55,N_152);
xnor U703 (N_703,N_254,N_450);
or U704 (N_704,N_2,N_410);
nor U705 (N_705,N_8,N_303);
nand U706 (N_706,N_52,N_306);
or U707 (N_707,N_419,N_219);
and U708 (N_708,N_324,N_315);
nand U709 (N_709,N_82,N_109);
and U710 (N_710,N_227,N_114);
or U711 (N_711,N_23,N_389);
nand U712 (N_712,N_10,N_88);
and U713 (N_713,N_458,N_454);
nor U714 (N_714,N_171,N_412);
and U715 (N_715,N_467,N_79);
and U716 (N_716,N_126,N_268);
nand U717 (N_717,N_116,N_251);
or U718 (N_718,N_411,N_85);
nor U719 (N_719,N_415,N_270);
nor U720 (N_720,N_394,N_235);
nor U721 (N_721,N_489,N_365);
or U722 (N_722,N_94,N_115);
and U723 (N_723,N_294,N_25);
or U724 (N_724,N_355,N_418);
or U725 (N_725,N_328,N_92);
nand U726 (N_726,N_388,N_66);
or U727 (N_727,N_304,N_349);
nor U728 (N_728,N_329,N_21);
nand U729 (N_729,N_236,N_341);
nor U730 (N_730,N_414,N_442);
or U731 (N_731,N_234,N_366);
nor U732 (N_732,N_57,N_208);
and U733 (N_733,N_125,N_140);
or U734 (N_734,N_325,N_247);
nand U735 (N_735,N_223,N_484);
and U736 (N_736,N_332,N_443);
xnor U737 (N_737,N_131,N_287);
nor U738 (N_738,N_72,N_295);
or U739 (N_739,N_258,N_370);
xnor U740 (N_740,N_218,N_356);
nand U741 (N_741,N_331,N_340);
xor U742 (N_742,N_316,N_225);
nand U743 (N_743,N_50,N_492);
or U744 (N_744,N_157,N_375);
nand U745 (N_745,N_381,N_300);
nand U746 (N_746,N_358,N_71);
nor U747 (N_747,N_403,N_149);
nor U748 (N_748,N_422,N_310);
xnor U749 (N_749,N_257,N_128);
and U750 (N_750,N_447,N_45);
nand U751 (N_751,N_441,N_193);
and U752 (N_752,N_95,N_495);
and U753 (N_753,N_455,N_90);
and U754 (N_754,N_225,N_32);
or U755 (N_755,N_33,N_133);
nor U756 (N_756,N_434,N_223);
xnor U757 (N_757,N_313,N_76);
nand U758 (N_758,N_51,N_1);
nor U759 (N_759,N_114,N_260);
xnor U760 (N_760,N_153,N_436);
nand U761 (N_761,N_442,N_136);
nor U762 (N_762,N_306,N_454);
nor U763 (N_763,N_143,N_100);
and U764 (N_764,N_245,N_208);
nor U765 (N_765,N_85,N_160);
nor U766 (N_766,N_62,N_480);
xor U767 (N_767,N_5,N_50);
xnor U768 (N_768,N_22,N_168);
and U769 (N_769,N_55,N_54);
nor U770 (N_770,N_86,N_412);
nor U771 (N_771,N_79,N_36);
nor U772 (N_772,N_449,N_270);
or U773 (N_773,N_58,N_111);
xnor U774 (N_774,N_338,N_30);
xor U775 (N_775,N_470,N_463);
nor U776 (N_776,N_288,N_133);
xnor U777 (N_777,N_494,N_34);
nor U778 (N_778,N_390,N_471);
or U779 (N_779,N_413,N_119);
nor U780 (N_780,N_399,N_63);
xnor U781 (N_781,N_455,N_99);
nor U782 (N_782,N_221,N_184);
or U783 (N_783,N_325,N_195);
and U784 (N_784,N_87,N_394);
nand U785 (N_785,N_26,N_352);
nor U786 (N_786,N_209,N_230);
nand U787 (N_787,N_460,N_204);
nor U788 (N_788,N_416,N_421);
nor U789 (N_789,N_78,N_48);
and U790 (N_790,N_296,N_87);
nor U791 (N_791,N_57,N_51);
or U792 (N_792,N_229,N_10);
xor U793 (N_793,N_478,N_496);
xor U794 (N_794,N_63,N_201);
nand U795 (N_795,N_2,N_328);
nor U796 (N_796,N_195,N_360);
and U797 (N_797,N_106,N_393);
xor U798 (N_798,N_414,N_78);
or U799 (N_799,N_19,N_55);
nand U800 (N_800,N_209,N_103);
nand U801 (N_801,N_135,N_438);
or U802 (N_802,N_133,N_459);
nor U803 (N_803,N_477,N_487);
or U804 (N_804,N_76,N_157);
xnor U805 (N_805,N_439,N_374);
or U806 (N_806,N_278,N_341);
nand U807 (N_807,N_249,N_328);
xnor U808 (N_808,N_237,N_97);
and U809 (N_809,N_442,N_214);
or U810 (N_810,N_24,N_332);
or U811 (N_811,N_289,N_20);
nor U812 (N_812,N_325,N_222);
and U813 (N_813,N_472,N_69);
and U814 (N_814,N_285,N_463);
nor U815 (N_815,N_341,N_186);
nand U816 (N_816,N_121,N_257);
nor U817 (N_817,N_391,N_246);
xor U818 (N_818,N_467,N_498);
and U819 (N_819,N_260,N_66);
nor U820 (N_820,N_96,N_491);
xnor U821 (N_821,N_446,N_439);
nand U822 (N_822,N_380,N_334);
nor U823 (N_823,N_91,N_240);
or U824 (N_824,N_294,N_376);
and U825 (N_825,N_61,N_461);
nand U826 (N_826,N_445,N_491);
and U827 (N_827,N_49,N_70);
nand U828 (N_828,N_285,N_389);
and U829 (N_829,N_4,N_47);
and U830 (N_830,N_19,N_104);
and U831 (N_831,N_395,N_381);
or U832 (N_832,N_382,N_470);
nand U833 (N_833,N_400,N_405);
and U834 (N_834,N_252,N_122);
nand U835 (N_835,N_312,N_311);
and U836 (N_836,N_4,N_17);
nor U837 (N_837,N_169,N_350);
nand U838 (N_838,N_160,N_447);
or U839 (N_839,N_323,N_34);
and U840 (N_840,N_353,N_334);
nor U841 (N_841,N_179,N_336);
or U842 (N_842,N_186,N_268);
nand U843 (N_843,N_131,N_249);
xor U844 (N_844,N_499,N_100);
and U845 (N_845,N_350,N_304);
nand U846 (N_846,N_138,N_201);
and U847 (N_847,N_458,N_397);
nor U848 (N_848,N_425,N_493);
nand U849 (N_849,N_22,N_15);
and U850 (N_850,N_281,N_83);
and U851 (N_851,N_193,N_119);
or U852 (N_852,N_50,N_362);
nand U853 (N_853,N_123,N_260);
nor U854 (N_854,N_306,N_286);
nand U855 (N_855,N_480,N_471);
nor U856 (N_856,N_331,N_53);
nor U857 (N_857,N_340,N_153);
and U858 (N_858,N_87,N_345);
nand U859 (N_859,N_89,N_65);
nand U860 (N_860,N_89,N_46);
or U861 (N_861,N_85,N_191);
nand U862 (N_862,N_142,N_146);
nand U863 (N_863,N_136,N_131);
nor U864 (N_864,N_249,N_374);
nor U865 (N_865,N_97,N_95);
nor U866 (N_866,N_132,N_350);
nand U867 (N_867,N_78,N_108);
nor U868 (N_868,N_8,N_98);
nor U869 (N_869,N_14,N_490);
nand U870 (N_870,N_149,N_171);
and U871 (N_871,N_78,N_17);
nor U872 (N_872,N_204,N_234);
nand U873 (N_873,N_121,N_422);
nor U874 (N_874,N_363,N_440);
nand U875 (N_875,N_13,N_294);
nor U876 (N_876,N_113,N_308);
and U877 (N_877,N_249,N_474);
xor U878 (N_878,N_419,N_332);
and U879 (N_879,N_149,N_294);
xor U880 (N_880,N_121,N_280);
nor U881 (N_881,N_347,N_196);
nor U882 (N_882,N_86,N_14);
nand U883 (N_883,N_413,N_2);
nand U884 (N_884,N_381,N_467);
nand U885 (N_885,N_144,N_35);
and U886 (N_886,N_276,N_135);
nand U887 (N_887,N_250,N_24);
or U888 (N_888,N_84,N_347);
xor U889 (N_889,N_379,N_424);
nand U890 (N_890,N_460,N_457);
nor U891 (N_891,N_50,N_319);
or U892 (N_892,N_197,N_248);
nand U893 (N_893,N_183,N_188);
and U894 (N_894,N_304,N_458);
xnor U895 (N_895,N_382,N_298);
nand U896 (N_896,N_449,N_463);
nor U897 (N_897,N_343,N_366);
and U898 (N_898,N_220,N_99);
nand U899 (N_899,N_230,N_6);
or U900 (N_900,N_369,N_442);
or U901 (N_901,N_260,N_435);
nor U902 (N_902,N_237,N_81);
and U903 (N_903,N_0,N_81);
and U904 (N_904,N_2,N_310);
nand U905 (N_905,N_325,N_153);
nor U906 (N_906,N_201,N_14);
or U907 (N_907,N_255,N_224);
and U908 (N_908,N_365,N_235);
nand U909 (N_909,N_129,N_96);
nor U910 (N_910,N_134,N_455);
or U911 (N_911,N_111,N_369);
nor U912 (N_912,N_134,N_153);
nor U913 (N_913,N_188,N_2);
and U914 (N_914,N_108,N_239);
nand U915 (N_915,N_207,N_398);
nand U916 (N_916,N_242,N_135);
nand U917 (N_917,N_218,N_58);
and U918 (N_918,N_270,N_456);
xnor U919 (N_919,N_159,N_395);
xnor U920 (N_920,N_469,N_17);
or U921 (N_921,N_174,N_5);
and U922 (N_922,N_184,N_378);
and U923 (N_923,N_147,N_194);
xor U924 (N_924,N_320,N_408);
or U925 (N_925,N_136,N_353);
and U926 (N_926,N_240,N_64);
and U927 (N_927,N_19,N_127);
nand U928 (N_928,N_298,N_176);
xnor U929 (N_929,N_312,N_288);
nor U930 (N_930,N_190,N_12);
and U931 (N_931,N_25,N_296);
xor U932 (N_932,N_397,N_494);
nand U933 (N_933,N_399,N_374);
and U934 (N_934,N_279,N_485);
nor U935 (N_935,N_86,N_482);
xnor U936 (N_936,N_467,N_165);
xnor U937 (N_937,N_279,N_262);
and U938 (N_938,N_137,N_302);
or U939 (N_939,N_317,N_129);
or U940 (N_940,N_223,N_189);
xnor U941 (N_941,N_430,N_477);
or U942 (N_942,N_484,N_188);
and U943 (N_943,N_401,N_262);
nand U944 (N_944,N_148,N_411);
nor U945 (N_945,N_165,N_100);
nand U946 (N_946,N_454,N_30);
xnor U947 (N_947,N_2,N_469);
nand U948 (N_948,N_414,N_165);
nor U949 (N_949,N_309,N_494);
or U950 (N_950,N_192,N_32);
or U951 (N_951,N_350,N_296);
nand U952 (N_952,N_388,N_67);
nand U953 (N_953,N_200,N_461);
nand U954 (N_954,N_135,N_463);
nor U955 (N_955,N_377,N_152);
or U956 (N_956,N_473,N_9);
or U957 (N_957,N_66,N_454);
nor U958 (N_958,N_284,N_46);
nand U959 (N_959,N_190,N_140);
or U960 (N_960,N_215,N_276);
or U961 (N_961,N_279,N_474);
nor U962 (N_962,N_444,N_10);
or U963 (N_963,N_485,N_283);
nor U964 (N_964,N_368,N_311);
nand U965 (N_965,N_114,N_190);
nor U966 (N_966,N_465,N_428);
and U967 (N_967,N_22,N_17);
or U968 (N_968,N_459,N_476);
nand U969 (N_969,N_194,N_418);
nand U970 (N_970,N_182,N_179);
and U971 (N_971,N_324,N_461);
nor U972 (N_972,N_194,N_279);
nand U973 (N_973,N_185,N_387);
xor U974 (N_974,N_13,N_193);
or U975 (N_975,N_155,N_453);
xnor U976 (N_976,N_280,N_358);
nand U977 (N_977,N_436,N_22);
xnor U978 (N_978,N_145,N_32);
and U979 (N_979,N_228,N_19);
nand U980 (N_980,N_329,N_123);
or U981 (N_981,N_419,N_204);
nand U982 (N_982,N_114,N_187);
xor U983 (N_983,N_321,N_279);
or U984 (N_984,N_199,N_158);
nor U985 (N_985,N_421,N_338);
nand U986 (N_986,N_82,N_125);
and U987 (N_987,N_115,N_95);
nand U988 (N_988,N_350,N_347);
nor U989 (N_989,N_388,N_474);
nor U990 (N_990,N_78,N_193);
nand U991 (N_991,N_262,N_126);
or U992 (N_992,N_435,N_453);
nand U993 (N_993,N_262,N_306);
nor U994 (N_994,N_494,N_10);
nand U995 (N_995,N_295,N_481);
or U996 (N_996,N_326,N_194);
nand U997 (N_997,N_332,N_439);
xnor U998 (N_998,N_325,N_413);
nor U999 (N_999,N_451,N_147);
nand U1000 (N_1000,N_943,N_824);
or U1001 (N_1001,N_823,N_842);
nor U1002 (N_1002,N_846,N_696);
nor U1003 (N_1003,N_795,N_936);
xor U1004 (N_1004,N_892,N_620);
and U1005 (N_1005,N_709,N_714);
and U1006 (N_1006,N_948,N_509);
nand U1007 (N_1007,N_703,N_672);
or U1008 (N_1008,N_661,N_970);
or U1009 (N_1009,N_656,N_651);
or U1010 (N_1010,N_544,N_767);
xnor U1011 (N_1011,N_588,N_616);
nand U1012 (N_1012,N_785,N_799);
and U1013 (N_1013,N_777,N_762);
xor U1014 (N_1014,N_671,N_551);
nor U1015 (N_1015,N_864,N_743);
or U1016 (N_1016,N_815,N_932);
nor U1017 (N_1017,N_708,N_707);
nand U1018 (N_1018,N_764,N_536);
or U1019 (N_1019,N_985,N_880);
and U1020 (N_1020,N_598,N_944);
and U1021 (N_1021,N_581,N_992);
nor U1022 (N_1022,N_918,N_926);
or U1023 (N_1023,N_939,N_821);
xor U1024 (N_1024,N_958,N_641);
nand U1025 (N_1025,N_726,N_582);
nand U1026 (N_1026,N_621,N_908);
or U1027 (N_1027,N_678,N_920);
and U1028 (N_1028,N_951,N_643);
or U1029 (N_1029,N_971,N_910);
nor U1030 (N_1030,N_800,N_954);
nor U1031 (N_1031,N_595,N_505);
nand U1032 (N_1032,N_521,N_534);
nor U1033 (N_1033,N_778,N_520);
or U1034 (N_1034,N_719,N_668);
and U1035 (N_1035,N_510,N_986);
nor U1036 (N_1036,N_749,N_981);
nand U1037 (N_1037,N_638,N_758);
and U1038 (N_1038,N_903,N_727);
xnor U1039 (N_1039,N_818,N_555);
and U1040 (N_1040,N_789,N_816);
nor U1041 (N_1041,N_596,N_828);
and U1042 (N_1042,N_806,N_938);
or U1043 (N_1043,N_655,N_820);
nand U1044 (N_1044,N_791,N_857);
nor U1045 (N_1045,N_997,N_539);
nor U1046 (N_1046,N_574,N_888);
and U1047 (N_1047,N_972,N_569);
and U1048 (N_1048,N_690,N_822);
and U1049 (N_1049,N_859,N_775);
nand U1050 (N_1050,N_950,N_717);
nor U1051 (N_1051,N_852,N_730);
and U1052 (N_1052,N_895,N_511);
and U1053 (N_1053,N_963,N_535);
nor U1054 (N_1054,N_660,N_677);
nor U1055 (N_1055,N_591,N_525);
nor U1056 (N_1056,N_884,N_866);
nand U1057 (N_1057,N_779,N_798);
nand U1058 (N_1058,N_692,N_922);
xor U1059 (N_1059,N_871,N_650);
nand U1060 (N_1060,N_770,N_759);
nor U1061 (N_1061,N_741,N_745);
or U1062 (N_1062,N_504,N_684);
nand U1063 (N_1063,N_604,N_585);
nor U1064 (N_1064,N_648,N_653);
nand U1065 (N_1065,N_645,N_836);
nand U1066 (N_1066,N_814,N_548);
or U1067 (N_1067,N_697,N_603);
nor U1068 (N_1068,N_786,N_945);
and U1069 (N_1069,N_896,N_790);
nand U1070 (N_1070,N_607,N_914);
xor U1071 (N_1071,N_729,N_952);
nor U1072 (N_1072,N_756,N_865);
nor U1073 (N_1073,N_959,N_538);
nand U1074 (N_1074,N_924,N_853);
and U1075 (N_1075,N_652,N_923);
nand U1076 (N_1076,N_832,N_988);
xnor U1077 (N_1077,N_975,N_872);
and U1078 (N_1078,N_769,N_990);
and U1079 (N_1079,N_606,N_722);
nor U1080 (N_1080,N_768,N_813);
nor U1081 (N_1081,N_545,N_506);
nor U1082 (N_1082,N_999,N_894);
nand U1083 (N_1083,N_875,N_565);
and U1084 (N_1084,N_844,N_869);
or U1085 (N_1085,N_782,N_710);
and U1086 (N_1086,N_850,N_568);
and U1087 (N_1087,N_704,N_556);
nand U1088 (N_1088,N_909,N_861);
or U1089 (N_1089,N_962,N_784);
nor U1090 (N_1090,N_517,N_526);
xnor U1091 (N_1091,N_961,N_615);
nor U1092 (N_1092,N_739,N_868);
nand U1093 (N_1093,N_841,N_738);
and U1094 (N_1094,N_883,N_977);
nand U1095 (N_1095,N_724,N_501);
and U1096 (N_1096,N_691,N_642);
nand U1097 (N_1097,N_734,N_874);
nand U1098 (N_1098,N_512,N_531);
nor U1099 (N_1099,N_628,N_564);
and U1100 (N_1100,N_748,N_755);
xnor U1101 (N_1101,N_687,N_601);
or U1102 (N_1102,N_592,N_803);
and U1103 (N_1103,N_984,N_693);
nor U1104 (N_1104,N_576,N_794);
or U1105 (N_1105,N_854,N_580);
nor U1106 (N_1106,N_787,N_974);
and U1107 (N_1107,N_837,N_766);
nor U1108 (N_1108,N_667,N_513);
and U1109 (N_1109,N_797,N_826);
or U1110 (N_1110,N_855,N_774);
nor U1111 (N_1111,N_553,N_674);
or U1112 (N_1112,N_847,N_680);
or U1113 (N_1113,N_560,N_681);
and U1114 (N_1114,N_781,N_978);
nand U1115 (N_1115,N_819,N_830);
and U1116 (N_1116,N_788,N_507);
nor U1117 (N_1117,N_810,N_736);
nand U1118 (N_1118,N_562,N_838);
nor U1119 (N_1119,N_809,N_527);
or U1120 (N_1120,N_503,N_802);
or U1121 (N_1121,N_827,N_715);
xnor U1122 (N_1122,N_662,N_593);
nand U1123 (N_1123,N_614,N_754);
nand U1124 (N_1124,N_751,N_829);
xnor U1125 (N_1125,N_533,N_519);
nor U1126 (N_1126,N_870,N_848);
or U1127 (N_1127,N_554,N_546);
nand U1128 (N_1128,N_969,N_502);
and U1129 (N_1129,N_904,N_612);
nand U1130 (N_1130,N_584,N_947);
nand U1131 (N_1131,N_624,N_608);
xnor U1132 (N_1132,N_522,N_843);
and U1133 (N_1133,N_634,N_640);
and U1134 (N_1134,N_925,N_528);
nand U1135 (N_1135,N_991,N_900);
nand U1136 (N_1136,N_566,N_907);
nor U1137 (N_1137,N_765,N_742);
or U1138 (N_1138,N_550,N_627);
and U1139 (N_1139,N_783,N_516);
and U1140 (N_1140,N_805,N_980);
xnor U1141 (N_1141,N_776,N_905);
nor U1142 (N_1142,N_863,N_801);
nand U1143 (N_1143,N_928,N_515);
xnor U1144 (N_1144,N_937,N_657);
or U1145 (N_1145,N_851,N_732);
nor U1146 (N_1146,N_773,N_597);
nor U1147 (N_1147,N_867,N_817);
nor U1148 (N_1148,N_658,N_839);
or U1149 (N_1149,N_686,N_858);
or U1150 (N_1150,N_699,N_898);
or U1151 (N_1151,N_682,N_740);
or U1152 (N_1152,N_968,N_733);
or U1153 (N_1153,N_639,N_885);
or U1154 (N_1154,N_917,N_600);
nor U1155 (N_1155,N_964,N_599);
and U1156 (N_1156,N_529,N_877);
and U1157 (N_1157,N_577,N_524);
xnor U1158 (N_1158,N_906,N_713);
or U1159 (N_1159,N_626,N_930);
nor U1160 (N_1160,N_889,N_716);
nand U1161 (N_1161,N_629,N_623);
or U1162 (N_1162,N_793,N_812);
or U1163 (N_1163,N_913,N_808);
nor U1164 (N_1164,N_646,N_594);
nand U1165 (N_1165,N_578,N_728);
nand U1166 (N_1166,N_675,N_780);
and U1167 (N_1167,N_664,N_845);
nor U1168 (N_1168,N_967,N_532);
or U1169 (N_1169,N_856,N_935);
nand U1170 (N_1170,N_637,N_747);
nor U1171 (N_1171,N_735,N_543);
nor U1172 (N_1172,N_725,N_698);
and U1173 (N_1173,N_610,N_630);
xor U1174 (N_1174,N_540,N_720);
or U1175 (N_1175,N_700,N_579);
nor U1176 (N_1176,N_583,N_995);
and U1177 (N_1177,N_567,N_835);
nand U1178 (N_1178,N_901,N_514);
nand U1179 (N_1179,N_669,N_609);
nand U1180 (N_1180,N_912,N_804);
xor U1181 (N_1181,N_942,N_763);
and U1182 (N_1182,N_915,N_688);
and U1183 (N_1183,N_929,N_670);
nor U1184 (N_1184,N_983,N_746);
and U1185 (N_1185,N_683,N_590);
and U1186 (N_1186,N_508,N_711);
and U1187 (N_1187,N_530,N_571);
nand U1188 (N_1188,N_941,N_635);
and U1189 (N_1189,N_723,N_994);
nor U1190 (N_1190,N_976,N_633);
or U1191 (N_1191,N_676,N_771);
or U1192 (N_1192,N_833,N_694);
nand U1193 (N_1193,N_622,N_721);
and U1194 (N_1194,N_921,N_993);
nand U1195 (N_1195,N_893,N_573);
nor U1196 (N_1196,N_750,N_831);
nand U1197 (N_1197,N_760,N_899);
and U1198 (N_1198,N_965,N_953);
nor U1199 (N_1199,N_542,N_575);
nor U1200 (N_1200,N_982,N_701);
xor U1201 (N_1201,N_689,N_996);
nor U1202 (N_1202,N_989,N_979);
nand U1203 (N_1203,N_570,N_807);
nand U1204 (N_1204,N_876,N_541);
or U1205 (N_1205,N_949,N_862);
or U1206 (N_1206,N_632,N_718);
nor U1207 (N_1207,N_957,N_523);
and U1208 (N_1208,N_625,N_811);
nand U1209 (N_1209,N_611,N_617);
and U1210 (N_1210,N_631,N_890);
nor U1211 (N_1211,N_879,N_916);
or U1212 (N_1212,N_605,N_860);
nand U1213 (N_1213,N_685,N_840);
and U1214 (N_1214,N_881,N_919);
xnor U1215 (N_1215,N_705,N_702);
or U1216 (N_1216,N_933,N_886);
nand U1217 (N_1217,N_589,N_834);
nor U1218 (N_1218,N_887,N_731);
nor U1219 (N_1219,N_679,N_558);
nand U1220 (N_1220,N_955,N_757);
and U1221 (N_1221,N_659,N_647);
nor U1222 (N_1222,N_761,N_613);
nor U1223 (N_1223,N_563,N_934);
nor U1224 (N_1224,N_602,N_946);
nand U1225 (N_1225,N_960,N_927);
nand U1226 (N_1226,N_618,N_549);
and U1227 (N_1227,N_902,N_940);
or U1228 (N_1228,N_897,N_649);
or U1229 (N_1229,N_644,N_973);
or U1230 (N_1230,N_849,N_636);
or U1231 (N_1231,N_882,N_998);
or U1232 (N_1232,N_737,N_878);
or U1233 (N_1233,N_557,N_911);
nor U1234 (N_1234,N_559,N_673);
nor U1235 (N_1235,N_772,N_931);
nand U1236 (N_1236,N_712,N_537);
and U1237 (N_1237,N_552,N_663);
nor U1238 (N_1238,N_706,N_752);
or U1239 (N_1239,N_666,N_825);
nor U1240 (N_1240,N_547,N_619);
and U1241 (N_1241,N_891,N_873);
and U1242 (N_1242,N_665,N_744);
nand U1243 (N_1243,N_956,N_500);
xor U1244 (N_1244,N_587,N_561);
nor U1245 (N_1245,N_654,N_753);
nand U1246 (N_1246,N_987,N_695);
nor U1247 (N_1247,N_792,N_966);
or U1248 (N_1248,N_572,N_586);
nor U1249 (N_1249,N_796,N_518);
xor U1250 (N_1250,N_914,N_878);
or U1251 (N_1251,N_911,N_807);
nor U1252 (N_1252,N_555,N_723);
xnor U1253 (N_1253,N_689,N_883);
xnor U1254 (N_1254,N_730,N_903);
or U1255 (N_1255,N_535,N_883);
nand U1256 (N_1256,N_698,N_594);
and U1257 (N_1257,N_707,N_529);
xnor U1258 (N_1258,N_890,N_617);
and U1259 (N_1259,N_823,N_989);
or U1260 (N_1260,N_814,N_688);
or U1261 (N_1261,N_663,N_921);
nor U1262 (N_1262,N_566,N_847);
nor U1263 (N_1263,N_869,N_676);
nand U1264 (N_1264,N_517,N_546);
nand U1265 (N_1265,N_772,N_894);
nand U1266 (N_1266,N_595,N_793);
and U1267 (N_1267,N_538,N_601);
nor U1268 (N_1268,N_800,N_647);
and U1269 (N_1269,N_886,N_957);
and U1270 (N_1270,N_565,N_840);
and U1271 (N_1271,N_656,N_838);
nand U1272 (N_1272,N_616,N_624);
and U1273 (N_1273,N_652,N_607);
nor U1274 (N_1274,N_677,N_950);
or U1275 (N_1275,N_660,N_513);
xor U1276 (N_1276,N_630,N_956);
nand U1277 (N_1277,N_741,N_666);
xor U1278 (N_1278,N_959,N_809);
nor U1279 (N_1279,N_586,N_952);
nand U1280 (N_1280,N_869,N_744);
nor U1281 (N_1281,N_618,N_866);
nand U1282 (N_1282,N_668,N_894);
or U1283 (N_1283,N_579,N_803);
nor U1284 (N_1284,N_728,N_554);
nand U1285 (N_1285,N_974,N_507);
nand U1286 (N_1286,N_790,N_702);
nand U1287 (N_1287,N_656,N_520);
or U1288 (N_1288,N_557,N_981);
or U1289 (N_1289,N_971,N_563);
or U1290 (N_1290,N_710,N_625);
and U1291 (N_1291,N_780,N_924);
xnor U1292 (N_1292,N_903,N_656);
or U1293 (N_1293,N_881,N_573);
nand U1294 (N_1294,N_643,N_516);
and U1295 (N_1295,N_887,N_554);
and U1296 (N_1296,N_572,N_776);
xnor U1297 (N_1297,N_975,N_749);
or U1298 (N_1298,N_599,N_825);
nand U1299 (N_1299,N_573,N_770);
nor U1300 (N_1300,N_893,N_998);
or U1301 (N_1301,N_954,N_872);
nand U1302 (N_1302,N_747,N_971);
nand U1303 (N_1303,N_934,N_831);
and U1304 (N_1304,N_875,N_685);
or U1305 (N_1305,N_900,N_769);
or U1306 (N_1306,N_706,N_943);
and U1307 (N_1307,N_848,N_537);
nor U1308 (N_1308,N_633,N_736);
or U1309 (N_1309,N_740,N_555);
and U1310 (N_1310,N_627,N_677);
and U1311 (N_1311,N_995,N_509);
nand U1312 (N_1312,N_734,N_704);
or U1313 (N_1313,N_579,N_598);
xnor U1314 (N_1314,N_954,N_735);
xor U1315 (N_1315,N_553,N_929);
and U1316 (N_1316,N_880,N_921);
and U1317 (N_1317,N_656,N_936);
nand U1318 (N_1318,N_934,N_931);
and U1319 (N_1319,N_578,N_822);
or U1320 (N_1320,N_957,N_782);
or U1321 (N_1321,N_793,N_682);
or U1322 (N_1322,N_851,N_587);
xnor U1323 (N_1323,N_557,N_875);
or U1324 (N_1324,N_625,N_814);
nor U1325 (N_1325,N_998,N_832);
nand U1326 (N_1326,N_665,N_554);
or U1327 (N_1327,N_570,N_642);
and U1328 (N_1328,N_838,N_770);
or U1329 (N_1329,N_573,N_539);
nor U1330 (N_1330,N_736,N_696);
nand U1331 (N_1331,N_524,N_931);
nand U1332 (N_1332,N_968,N_680);
xor U1333 (N_1333,N_654,N_974);
and U1334 (N_1334,N_849,N_572);
or U1335 (N_1335,N_735,N_744);
nand U1336 (N_1336,N_637,N_848);
and U1337 (N_1337,N_729,N_632);
or U1338 (N_1338,N_748,N_782);
nand U1339 (N_1339,N_944,N_784);
nand U1340 (N_1340,N_787,N_794);
and U1341 (N_1341,N_968,N_763);
and U1342 (N_1342,N_659,N_536);
xor U1343 (N_1343,N_662,N_960);
nand U1344 (N_1344,N_903,N_960);
nand U1345 (N_1345,N_936,N_745);
and U1346 (N_1346,N_817,N_970);
nor U1347 (N_1347,N_819,N_874);
and U1348 (N_1348,N_529,N_598);
xnor U1349 (N_1349,N_584,N_596);
or U1350 (N_1350,N_761,N_758);
and U1351 (N_1351,N_545,N_916);
nand U1352 (N_1352,N_652,N_930);
xor U1353 (N_1353,N_791,N_785);
nor U1354 (N_1354,N_535,N_923);
nand U1355 (N_1355,N_843,N_534);
nand U1356 (N_1356,N_526,N_794);
or U1357 (N_1357,N_834,N_690);
nand U1358 (N_1358,N_573,N_948);
and U1359 (N_1359,N_950,N_657);
nor U1360 (N_1360,N_767,N_626);
xor U1361 (N_1361,N_748,N_873);
or U1362 (N_1362,N_972,N_994);
and U1363 (N_1363,N_734,N_706);
and U1364 (N_1364,N_828,N_637);
and U1365 (N_1365,N_956,N_893);
nand U1366 (N_1366,N_584,N_785);
or U1367 (N_1367,N_531,N_735);
or U1368 (N_1368,N_826,N_983);
and U1369 (N_1369,N_525,N_507);
or U1370 (N_1370,N_862,N_693);
nand U1371 (N_1371,N_861,N_514);
nor U1372 (N_1372,N_775,N_776);
nor U1373 (N_1373,N_666,N_613);
nand U1374 (N_1374,N_905,N_688);
xnor U1375 (N_1375,N_734,N_913);
and U1376 (N_1376,N_816,N_802);
and U1377 (N_1377,N_792,N_911);
nor U1378 (N_1378,N_750,N_604);
and U1379 (N_1379,N_948,N_908);
nand U1380 (N_1380,N_633,N_895);
nand U1381 (N_1381,N_914,N_710);
and U1382 (N_1382,N_651,N_950);
and U1383 (N_1383,N_764,N_728);
xnor U1384 (N_1384,N_735,N_763);
nor U1385 (N_1385,N_766,N_665);
and U1386 (N_1386,N_660,N_851);
or U1387 (N_1387,N_831,N_960);
or U1388 (N_1388,N_786,N_518);
and U1389 (N_1389,N_582,N_522);
xor U1390 (N_1390,N_993,N_931);
nand U1391 (N_1391,N_652,N_795);
nor U1392 (N_1392,N_642,N_628);
nor U1393 (N_1393,N_936,N_901);
or U1394 (N_1394,N_632,N_666);
xnor U1395 (N_1395,N_837,N_769);
or U1396 (N_1396,N_536,N_790);
nor U1397 (N_1397,N_981,N_705);
nor U1398 (N_1398,N_952,N_978);
xor U1399 (N_1399,N_569,N_579);
and U1400 (N_1400,N_526,N_936);
nand U1401 (N_1401,N_799,N_830);
nor U1402 (N_1402,N_738,N_781);
nand U1403 (N_1403,N_876,N_824);
or U1404 (N_1404,N_549,N_836);
and U1405 (N_1405,N_982,N_976);
nand U1406 (N_1406,N_783,N_601);
nand U1407 (N_1407,N_569,N_907);
nand U1408 (N_1408,N_856,N_887);
and U1409 (N_1409,N_788,N_831);
or U1410 (N_1410,N_515,N_856);
or U1411 (N_1411,N_747,N_994);
or U1412 (N_1412,N_795,N_721);
nor U1413 (N_1413,N_885,N_973);
or U1414 (N_1414,N_601,N_654);
nor U1415 (N_1415,N_825,N_679);
nor U1416 (N_1416,N_523,N_966);
and U1417 (N_1417,N_977,N_851);
and U1418 (N_1418,N_803,N_993);
or U1419 (N_1419,N_648,N_623);
nand U1420 (N_1420,N_616,N_777);
xor U1421 (N_1421,N_932,N_970);
nand U1422 (N_1422,N_846,N_745);
or U1423 (N_1423,N_508,N_682);
and U1424 (N_1424,N_596,N_570);
or U1425 (N_1425,N_814,N_528);
nand U1426 (N_1426,N_883,N_660);
xnor U1427 (N_1427,N_968,N_737);
nor U1428 (N_1428,N_618,N_608);
or U1429 (N_1429,N_895,N_551);
nand U1430 (N_1430,N_809,N_708);
xnor U1431 (N_1431,N_726,N_671);
or U1432 (N_1432,N_906,N_743);
xor U1433 (N_1433,N_822,N_515);
nand U1434 (N_1434,N_770,N_801);
or U1435 (N_1435,N_804,N_533);
nand U1436 (N_1436,N_989,N_877);
or U1437 (N_1437,N_635,N_877);
and U1438 (N_1438,N_802,N_601);
nor U1439 (N_1439,N_989,N_604);
or U1440 (N_1440,N_653,N_876);
or U1441 (N_1441,N_961,N_899);
or U1442 (N_1442,N_548,N_817);
or U1443 (N_1443,N_771,N_539);
or U1444 (N_1444,N_945,N_669);
and U1445 (N_1445,N_937,N_706);
nand U1446 (N_1446,N_723,N_995);
xor U1447 (N_1447,N_837,N_771);
nand U1448 (N_1448,N_938,N_786);
nand U1449 (N_1449,N_808,N_545);
and U1450 (N_1450,N_846,N_535);
and U1451 (N_1451,N_725,N_918);
xnor U1452 (N_1452,N_766,N_582);
and U1453 (N_1453,N_940,N_971);
nor U1454 (N_1454,N_590,N_745);
nand U1455 (N_1455,N_668,N_522);
nor U1456 (N_1456,N_906,N_712);
and U1457 (N_1457,N_713,N_864);
or U1458 (N_1458,N_966,N_617);
xor U1459 (N_1459,N_725,N_768);
nor U1460 (N_1460,N_946,N_702);
xor U1461 (N_1461,N_993,N_538);
nor U1462 (N_1462,N_775,N_655);
nor U1463 (N_1463,N_839,N_900);
nand U1464 (N_1464,N_943,N_761);
xor U1465 (N_1465,N_791,N_687);
or U1466 (N_1466,N_500,N_511);
nor U1467 (N_1467,N_991,N_948);
nor U1468 (N_1468,N_618,N_578);
nor U1469 (N_1469,N_666,N_758);
xnor U1470 (N_1470,N_586,N_924);
nand U1471 (N_1471,N_786,N_690);
nor U1472 (N_1472,N_689,N_759);
nand U1473 (N_1473,N_534,N_578);
nand U1474 (N_1474,N_565,N_968);
or U1475 (N_1475,N_811,N_805);
nor U1476 (N_1476,N_734,N_737);
and U1477 (N_1477,N_547,N_722);
nor U1478 (N_1478,N_638,N_545);
nand U1479 (N_1479,N_642,N_823);
nand U1480 (N_1480,N_943,N_781);
or U1481 (N_1481,N_593,N_909);
nor U1482 (N_1482,N_804,N_845);
nor U1483 (N_1483,N_905,N_858);
nand U1484 (N_1484,N_896,N_723);
or U1485 (N_1485,N_559,N_860);
nor U1486 (N_1486,N_692,N_958);
nor U1487 (N_1487,N_593,N_526);
and U1488 (N_1488,N_512,N_841);
or U1489 (N_1489,N_876,N_928);
or U1490 (N_1490,N_825,N_579);
nand U1491 (N_1491,N_975,N_931);
and U1492 (N_1492,N_586,N_991);
nor U1493 (N_1493,N_749,N_517);
and U1494 (N_1494,N_949,N_526);
xnor U1495 (N_1495,N_805,N_645);
or U1496 (N_1496,N_991,N_728);
and U1497 (N_1497,N_641,N_775);
nand U1498 (N_1498,N_831,N_865);
or U1499 (N_1499,N_989,N_739);
nand U1500 (N_1500,N_1024,N_1468);
nand U1501 (N_1501,N_1200,N_1148);
or U1502 (N_1502,N_1220,N_1422);
nand U1503 (N_1503,N_1396,N_1231);
xnor U1504 (N_1504,N_1487,N_1262);
and U1505 (N_1505,N_1432,N_1219);
and U1506 (N_1506,N_1031,N_1064);
and U1507 (N_1507,N_1009,N_1176);
nor U1508 (N_1508,N_1165,N_1347);
nand U1509 (N_1509,N_1315,N_1107);
nor U1510 (N_1510,N_1479,N_1384);
nand U1511 (N_1511,N_1074,N_1483);
and U1512 (N_1512,N_1252,N_1195);
and U1513 (N_1513,N_1154,N_1242);
and U1514 (N_1514,N_1232,N_1298);
or U1515 (N_1515,N_1360,N_1039);
xor U1516 (N_1516,N_1060,N_1282);
nor U1517 (N_1517,N_1291,N_1289);
and U1518 (N_1518,N_1378,N_1029);
nand U1519 (N_1519,N_1164,N_1476);
nand U1520 (N_1520,N_1377,N_1265);
or U1521 (N_1521,N_1363,N_1136);
nand U1522 (N_1522,N_1145,N_1144);
nor U1523 (N_1523,N_1425,N_1488);
and U1524 (N_1524,N_1317,N_1052);
and U1525 (N_1525,N_1448,N_1157);
nor U1526 (N_1526,N_1278,N_1383);
or U1527 (N_1527,N_1070,N_1345);
nor U1528 (N_1528,N_1019,N_1301);
nand U1529 (N_1529,N_1130,N_1208);
or U1530 (N_1530,N_1055,N_1050);
nand U1531 (N_1531,N_1350,N_1417);
or U1532 (N_1532,N_1359,N_1201);
nand U1533 (N_1533,N_1471,N_1192);
nand U1534 (N_1534,N_1096,N_1333);
nor U1535 (N_1535,N_1431,N_1123);
nor U1536 (N_1536,N_1057,N_1373);
or U1537 (N_1537,N_1000,N_1270);
and U1538 (N_1538,N_1048,N_1106);
nor U1539 (N_1539,N_1484,N_1076);
or U1540 (N_1540,N_1111,N_1013);
and U1541 (N_1541,N_1305,N_1372);
xnor U1542 (N_1542,N_1427,N_1120);
nor U1543 (N_1543,N_1103,N_1011);
nand U1544 (N_1544,N_1250,N_1126);
nor U1545 (N_1545,N_1433,N_1406);
and U1546 (N_1546,N_1085,N_1086);
and U1547 (N_1547,N_1386,N_1408);
or U1548 (N_1548,N_1400,N_1495);
and U1549 (N_1549,N_1409,N_1131);
xor U1550 (N_1550,N_1253,N_1230);
nand U1551 (N_1551,N_1038,N_1014);
or U1552 (N_1552,N_1261,N_1292);
nor U1553 (N_1553,N_1065,N_1355);
nand U1554 (N_1554,N_1159,N_1216);
nor U1555 (N_1555,N_1303,N_1366);
nand U1556 (N_1556,N_1438,N_1343);
or U1557 (N_1557,N_1444,N_1089);
xnor U1558 (N_1558,N_1385,N_1094);
nand U1559 (N_1559,N_1277,N_1247);
nand U1560 (N_1560,N_1498,N_1135);
xnor U1561 (N_1561,N_1022,N_1117);
nor U1562 (N_1562,N_1239,N_1332);
nand U1563 (N_1563,N_1235,N_1110);
xnor U1564 (N_1564,N_1069,N_1478);
or U1565 (N_1565,N_1229,N_1045);
or U1566 (N_1566,N_1286,N_1274);
and U1567 (N_1567,N_1205,N_1115);
nor U1568 (N_1568,N_1391,N_1420);
or U1569 (N_1569,N_1461,N_1204);
nand U1570 (N_1570,N_1306,N_1424);
and U1571 (N_1571,N_1440,N_1156);
nor U1572 (N_1572,N_1462,N_1358);
or U1573 (N_1573,N_1007,N_1302);
nand U1574 (N_1574,N_1264,N_1403);
nor U1575 (N_1575,N_1179,N_1489);
and U1576 (N_1576,N_1327,N_1132);
and U1577 (N_1577,N_1101,N_1362);
nand U1578 (N_1578,N_1098,N_1062);
nand U1579 (N_1579,N_1356,N_1324);
nand U1580 (N_1580,N_1402,N_1410);
nand U1581 (N_1581,N_1267,N_1017);
xor U1582 (N_1582,N_1442,N_1405);
or U1583 (N_1583,N_1293,N_1049);
and U1584 (N_1584,N_1464,N_1399);
or U1585 (N_1585,N_1199,N_1097);
or U1586 (N_1586,N_1434,N_1341);
or U1587 (N_1587,N_1194,N_1416);
nor U1588 (N_1588,N_1326,N_1349);
or U1589 (N_1589,N_1227,N_1166);
or U1590 (N_1590,N_1281,N_1459);
nand U1591 (N_1591,N_1285,N_1236);
nor U1592 (N_1592,N_1037,N_1351);
nand U1593 (N_1593,N_1380,N_1041);
nor U1594 (N_1594,N_1002,N_1423);
or U1595 (N_1595,N_1241,N_1091);
nor U1596 (N_1596,N_1240,N_1419);
nor U1597 (N_1597,N_1309,N_1173);
nor U1598 (N_1598,N_1088,N_1469);
nor U1599 (N_1599,N_1284,N_1467);
nand U1600 (N_1600,N_1042,N_1397);
nand U1601 (N_1601,N_1214,N_1139);
nor U1602 (N_1602,N_1446,N_1105);
nor U1603 (N_1603,N_1122,N_1246);
and U1604 (N_1604,N_1369,N_1212);
nor U1605 (N_1605,N_1357,N_1388);
nand U1606 (N_1606,N_1348,N_1217);
and U1607 (N_1607,N_1206,N_1001);
nor U1608 (N_1608,N_1087,N_1150);
or U1609 (N_1609,N_1381,N_1251);
nand U1610 (N_1610,N_1485,N_1137);
and U1611 (N_1611,N_1304,N_1268);
xor U1612 (N_1612,N_1053,N_1295);
or U1613 (N_1613,N_1223,N_1497);
or U1614 (N_1614,N_1015,N_1003);
nor U1615 (N_1615,N_1443,N_1193);
nor U1616 (N_1616,N_1140,N_1294);
nand U1617 (N_1617,N_1296,N_1346);
nor U1618 (N_1618,N_1210,N_1340);
xnor U1619 (N_1619,N_1477,N_1414);
xnor U1620 (N_1620,N_1012,N_1496);
nand U1621 (N_1621,N_1028,N_1224);
and U1622 (N_1622,N_1191,N_1319);
nand U1623 (N_1623,N_1170,N_1233);
nand U1624 (N_1624,N_1280,N_1134);
nand U1625 (N_1625,N_1034,N_1389);
or U1626 (N_1626,N_1339,N_1472);
or U1627 (N_1627,N_1260,N_1272);
nand U1628 (N_1628,N_1186,N_1313);
nand U1629 (N_1629,N_1033,N_1175);
nand U1630 (N_1630,N_1300,N_1492);
and U1631 (N_1631,N_1211,N_1474);
xnor U1632 (N_1632,N_1162,N_1411);
or U1633 (N_1633,N_1083,N_1092);
nor U1634 (N_1634,N_1138,N_1177);
nor U1635 (N_1635,N_1256,N_1109);
nor U1636 (N_1636,N_1435,N_1353);
or U1637 (N_1637,N_1008,N_1198);
and U1638 (N_1638,N_1202,N_1452);
nor U1639 (N_1639,N_1401,N_1054);
xor U1640 (N_1640,N_1445,N_1104);
and U1641 (N_1641,N_1382,N_1125);
nand U1642 (N_1642,N_1335,N_1141);
and U1643 (N_1643,N_1451,N_1412);
xor U1644 (N_1644,N_1330,N_1153);
nor U1645 (N_1645,N_1066,N_1259);
xnor U1646 (N_1646,N_1116,N_1093);
nand U1647 (N_1647,N_1393,N_1390);
nand U1648 (N_1648,N_1171,N_1428);
or U1649 (N_1649,N_1430,N_1158);
nor U1650 (N_1650,N_1482,N_1370);
nand U1651 (N_1651,N_1222,N_1079);
and U1652 (N_1652,N_1456,N_1481);
and U1653 (N_1653,N_1082,N_1178);
and U1654 (N_1654,N_1470,N_1119);
nand U1655 (N_1655,N_1203,N_1100);
or U1656 (N_1656,N_1458,N_1245);
nand U1657 (N_1657,N_1290,N_1322);
or U1658 (N_1658,N_1404,N_1344);
and U1659 (N_1659,N_1486,N_1027);
nand U1660 (N_1660,N_1004,N_1398);
and U1661 (N_1661,N_1387,N_1044);
nand U1662 (N_1662,N_1465,N_1318);
and U1663 (N_1663,N_1258,N_1328);
nor U1664 (N_1664,N_1151,N_1321);
and U1665 (N_1665,N_1075,N_1421);
and U1666 (N_1666,N_1226,N_1243);
nor U1667 (N_1667,N_1127,N_1374);
or U1668 (N_1668,N_1121,N_1215);
nand U1669 (N_1669,N_1426,N_1276);
or U1670 (N_1670,N_1187,N_1102);
nand U1671 (N_1671,N_1084,N_1081);
nand U1672 (N_1672,N_1437,N_1006);
or U1673 (N_1673,N_1407,N_1257);
nand U1674 (N_1674,N_1283,N_1189);
nor U1675 (N_1675,N_1297,N_1376);
nand U1676 (N_1676,N_1475,N_1287);
nor U1677 (N_1677,N_1149,N_1018);
nand U1678 (N_1678,N_1196,N_1371);
or U1679 (N_1679,N_1271,N_1334);
nand U1680 (N_1680,N_1180,N_1244);
or U1681 (N_1681,N_1310,N_1112);
nor U1682 (N_1682,N_1168,N_1450);
nand U1683 (N_1683,N_1466,N_1213);
nor U1684 (N_1684,N_1364,N_1061);
and U1685 (N_1685,N_1113,N_1457);
or U1686 (N_1686,N_1128,N_1169);
and U1687 (N_1687,N_1147,N_1368);
and U1688 (N_1688,N_1207,N_1181);
or U1689 (N_1689,N_1172,N_1067);
nand U1690 (N_1690,N_1248,N_1299);
or U1691 (N_1691,N_1020,N_1152);
and U1692 (N_1692,N_1454,N_1323);
nand U1693 (N_1693,N_1026,N_1182);
and U1694 (N_1694,N_1225,N_1439);
or U1695 (N_1695,N_1255,N_1118);
nor U1696 (N_1696,N_1160,N_1447);
or U1697 (N_1697,N_1312,N_1491);
or U1698 (N_1698,N_1030,N_1056);
nor U1699 (N_1699,N_1059,N_1071);
xor U1700 (N_1700,N_1016,N_1392);
nand U1701 (N_1701,N_1249,N_1320);
nand U1702 (N_1702,N_1429,N_1314);
nor U1703 (N_1703,N_1394,N_1367);
nor U1704 (N_1704,N_1036,N_1266);
xor U1705 (N_1705,N_1218,N_1337);
nor U1706 (N_1706,N_1413,N_1190);
and U1707 (N_1707,N_1338,N_1035);
nor U1708 (N_1708,N_1124,N_1418);
or U1709 (N_1709,N_1078,N_1073);
nand U1710 (N_1710,N_1342,N_1209);
nand U1711 (N_1711,N_1493,N_1129);
nand U1712 (N_1712,N_1254,N_1005);
xnor U1713 (N_1713,N_1237,N_1463);
xor U1714 (N_1714,N_1161,N_1032);
or U1715 (N_1715,N_1436,N_1234);
and U1716 (N_1716,N_1269,N_1279);
or U1717 (N_1717,N_1375,N_1114);
nor U1718 (N_1718,N_1494,N_1480);
xor U1719 (N_1719,N_1329,N_1184);
and U1720 (N_1720,N_1490,N_1021);
and U1721 (N_1721,N_1040,N_1415);
or U1722 (N_1722,N_1197,N_1025);
and U1723 (N_1723,N_1188,N_1095);
and U1724 (N_1724,N_1441,N_1099);
nor U1725 (N_1725,N_1307,N_1275);
or U1726 (N_1726,N_1325,N_1072);
nand U1727 (N_1727,N_1288,N_1449);
xor U1728 (N_1728,N_1331,N_1273);
xnor U1729 (N_1729,N_1473,N_1058);
or U1730 (N_1730,N_1395,N_1311);
nor U1731 (N_1731,N_1263,N_1046);
nand U1732 (N_1732,N_1108,N_1185);
or U1733 (N_1733,N_1308,N_1051);
and U1734 (N_1734,N_1047,N_1155);
or U1735 (N_1735,N_1077,N_1221);
nand U1736 (N_1736,N_1174,N_1090);
nor U1737 (N_1737,N_1023,N_1080);
nand U1738 (N_1738,N_1142,N_1365);
or U1739 (N_1739,N_1455,N_1460);
or U1740 (N_1740,N_1453,N_1379);
nor U1741 (N_1741,N_1183,N_1361);
nor U1742 (N_1742,N_1010,N_1228);
or U1743 (N_1743,N_1238,N_1163);
nand U1744 (N_1744,N_1063,N_1068);
or U1745 (N_1745,N_1133,N_1043);
or U1746 (N_1746,N_1143,N_1336);
or U1747 (N_1747,N_1354,N_1146);
nand U1748 (N_1748,N_1316,N_1499);
nand U1749 (N_1749,N_1167,N_1352);
and U1750 (N_1750,N_1491,N_1381);
nand U1751 (N_1751,N_1057,N_1109);
xnor U1752 (N_1752,N_1107,N_1153);
nor U1753 (N_1753,N_1080,N_1094);
nor U1754 (N_1754,N_1394,N_1216);
nand U1755 (N_1755,N_1304,N_1099);
nand U1756 (N_1756,N_1341,N_1139);
or U1757 (N_1757,N_1257,N_1362);
nor U1758 (N_1758,N_1322,N_1029);
xnor U1759 (N_1759,N_1180,N_1427);
and U1760 (N_1760,N_1392,N_1150);
nor U1761 (N_1761,N_1309,N_1080);
nand U1762 (N_1762,N_1357,N_1330);
or U1763 (N_1763,N_1473,N_1216);
nor U1764 (N_1764,N_1085,N_1235);
xor U1765 (N_1765,N_1095,N_1114);
or U1766 (N_1766,N_1003,N_1045);
nor U1767 (N_1767,N_1251,N_1485);
or U1768 (N_1768,N_1169,N_1161);
nor U1769 (N_1769,N_1367,N_1037);
and U1770 (N_1770,N_1112,N_1284);
or U1771 (N_1771,N_1143,N_1092);
and U1772 (N_1772,N_1234,N_1359);
nand U1773 (N_1773,N_1372,N_1192);
or U1774 (N_1774,N_1171,N_1262);
nand U1775 (N_1775,N_1029,N_1321);
nor U1776 (N_1776,N_1139,N_1476);
and U1777 (N_1777,N_1121,N_1345);
or U1778 (N_1778,N_1317,N_1282);
or U1779 (N_1779,N_1217,N_1283);
nor U1780 (N_1780,N_1074,N_1055);
and U1781 (N_1781,N_1390,N_1276);
or U1782 (N_1782,N_1439,N_1482);
nand U1783 (N_1783,N_1286,N_1065);
nor U1784 (N_1784,N_1114,N_1196);
nor U1785 (N_1785,N_1181,N_1031);
nor U1786 (N_1786,N_1178,N_1224);
and U1787 (N_1787,N_1342,N_1244);
and U1788 (N_1788,N_1211,N_1291);
or U1789 (N_1789,N_1338,N_1446);
nor U1790 (N_1790,N_1322,N_1362);
nor U1791 (N_1791,N_1166,N_1440);
xnor U1792 (N_1792,N_1037,N_1011);
or U1793 (N_1793,N_1346,N_1238);
nand U1794 (N_1794,N_1210,N_1416);
or U1795 (N_1795,N_1278,N_1411);
nand U1796 (N_1796,N_1366,N_1460);
and U1797 (N_1797,N_1308,N_1351);
or U1798 (N_1798,N_1283,N_1292);
xnor U1799 (N_1799,N_1247,N_1097);
nor U1800 (N_1800,N_1221,N_1452);
nor U1801 (N_1801,N_1391,N_1168);
and U1802 (N_1802,N_1145,N_1350);
nor U1803 (N_1803,N_1070,N_1131);
and U1804 (N_1804,N_1435,N_1019);
nand U1805 (N_1805,N_1212,N_1240);
or U1806 (N_1806,N_1262,N_1183);
nor U1807 (N_1807,N_1173,N_1187);
nor U1808 (N_1808,N_1140,N_1160);
nand U1809 (N_1809,N_1095,N_1034);
nand U1810 (N_1810,N_1193,N_1325);
xnor U1811 (N_1811,N_1064,N_1072);
nor U1812 (N_1812,N_1465,N_1079);
or U1813 (N_1813,N_1315,N_1386);
and U1814 (N_1814,N_1252,N_1143);
nor U1815 (N_1815,N_1467,N_1120);
nor U1816 (N_1816,N_1217,N_1114);
or U1817 (N_1817,N_1436,N_1136);
or U1818 (N_1818,N_1391,N_1488);
and U1819 (N_1819,N_1260,N_1402);
nand U1820 (N_1820,N_1290,N_1092);
xor U1821 (N_1821,N_1279,N_1367);
xnor U1822 (N_1822,N_1483,N_1078);
or U1823 (N_1823,N_1238,N_1255);
nand U1824 (N_1824,N_1495,N_1134);
nand U1825 (N_1825,N_1105,N_1322);
nand U1826 (N_1826,N_1321,N_1038);
nor U1827 (N_1827,N_1339,N_1060);
or U1828 (N_1828,N_1300,N_1198);
or U1829 (N_1829,N_1229,N_1344);
nand U1830 (N_1830,N_1488,N_1221);
nor U1831 (N_1831,N_1464,N_1417);
nor U1832 (N_1832,N_1349,N_1493);
and U1833 (N_1833,N_1026,N_1020);
or U1834 (N_1834,N_1322,N_1295);
and U1835 (N_1835,N_1495,N_1191);
nor U1836 (N_1836,N_1100,N_1036);
xnor U1837 (N_1837,N_1303,N_1377);
and U1838 (N_1838,N_1477,N_1432);
or U1839 (N_1839,N_1102,N_1315);
nor U1840 (N_1840,N_1048,N_1411);
or U1841 (N_1841,N_1402,N_1132);
nand U1842 (N_1842,N_1241,N_1393);
nor U1843 (N_1843,N_1129,N_1144);
nand U1844 (N_1844,N_1382,N_1035);
nor U1845 (N_1845,N_1492,N_1459);
or U1846 (N_1846,N_1034,N_1237);
and U1847 (N_1847,N_1112,N_1286);
xor U1848 (N_1848,N_1394,N_1264);
or U1849 (N_1849,N_1083,N_1111);
nor U1850 (N_1850,N_1017,N_1083);
nand U1851 (N_1851,N_1161,N_1192);
xnor U1852 (N_1852,N_1294,N_1379);
nand U1853 (N_1853,N_1079,N_1042);
and U1854 (N_1854,N_1011,N_1106);
xor U1855 (N_1855,N_1419,N_1347);
nand U1856 (N_1856,N_1483,N_1300);
nand U1857 (N_1857,N_1118,N_1220);
or U1858 (N_1858,N_1160,N_1133);
and U1859 (N_1859,N_1216,N_1162);
or U1860 (N_1860,N_1487,N_1018);
nor U1861 (N_1861,N_1362,N_1462);
nor U1862 (N_1862,N_1012,N_1291);
nand U1863 (N_1863,N_1485,N_1483);
nor U1864 (N_1864,N_1353,N_1397);
and U1865 (N_1865,N_1436,N_1489);
and U1866 (N_1866,N_1349,N_1298);
or U1867 (N_1867,N_1026,N_1375);
nor U1868 (N_1868,N_1234,N_1313);
nand U1869 (N_1869,N_1050,N_1046);
nor U1870 (N_1870,N_1166,N_1491);
or U1871 (N_1871,N_1332,N_1088);
or U1872 (N_1872,N_1243,N_1475);
and U1873 (N_1873,N_1399,N_1082);
nor U1874 (N_1874,N_1097,N_1228);
nor U1875 (N_1875,N_1317,N_1440);
nand U1876 (N_1876,N_1262,N_1035);
xnor U1877 (N_1877,N_1348,N_1009);
or U1878 (N_1878,N_1084,N_1322);
nor U1879 (N_1879,N_1166,N_1124);
or U1880 (N_1880,N_1419,N_1331);
nor U1881 (N_1881,N_1367,N_1318);
or U1882 (N_1882,N_1011,N_1481);
nand U1883 (N_1883,N_1086,N_1327);
or U1884 (N_1884,N_1133,N_1303);
nand U1885 (N_1885,N_1239,N_1409);
nor U1886 (N_1886,N_1128,N_1284);
xor U1887 (N_1887,N_1008,N_1167);
and U1888 (N_1888,N_1226,N_1382);
nor U1889 (N_1889,N_1366,N_1325);
nor U1890 (N_1890,N_1034,N_1129);
nand U1891 (N_1891,N_1335,N_1492);
and U1892 (N_1892,N_1354,N_1304);
nand U1893 (N_1893,N_1194,N_1418);
nor U1894 (N_1894,N_1055,N_1312);
nand U1895 (N_1895,N_1483,N_1076);
or U1896 (N_1896,N_1199,N_1059);
and U1897 (N_1897,N_1298,N_1240);
nand U1898 (N_1898,N_1178,N_1174);
xnor U1899 (N_1899,N_1161,N_1140);
nand U1900 (N_1900,N_1098,N_1096);
or U1901 (N_1901,N_1227,N_1115);
or U1902 (N_1902,N_1405,N_1318);
nand U1903 (N_1903,N_1138,N_1208);
or U1904 (N_1904,N_1347,N_1156);
or U1905 (N_1905,N_1364,N_1323);
nand U1906 (N_1906,N_1463,N_1234);
and U1907 (N_1907,N_1245,N_1340);
and U1908 (N_1908,N_1078,N_1260);
or U1909 (N_1909,N_1431,N_1459);
nand U1910 (N_1910,N_1351,N_1026);
and U1911 (N_1911,N_1002,N_1080);
nand U1912 (N_1912,N_1110,N_1184);
nand U1913 (N_1913,N_1106,N_1084);
and U1914 (N_1914,N_1469,N_1354);
and U1915 (N_1915,N_1383,N_1164);
nand U1916 (N_1916,N_1052,N_1206);
or U1917 (N_1917,N_1406,N_1079);
nand U1918 (N_1918,N_1038,N_1199);
or U1919 (N_1919,N_1100,N_1027);
nor U1920 (N_1920,N_1205,N_1270);
nor U1921 (N_1921,N_1335,N_1040);
or U1922 (N_1922,N_1310,N_1201);
nor U1923 (N_1923,N_1228,N_1335);
nand U1924 (N_1924,N_1175,N_1170);
nand U1925 (N_1925,N_1079,N_1118);
and U1926 (N_1926,N_1108,N_1388);
nor U1927 (N_1927,N_1054,N_1237);
nor U1928 (N_1928,N_1058,N_1482);
or U1929 (N_1929,N_1136,N_1013);
and U1930 (N_1930,N_1118,N_1404);
nor U1931 (N_1931,N_1371,N_1304);
and U1932 (N_1932,N_1197,N_1301);
and U1933 (N_1933,N_1472,N_1493);
or U1934 (N_1934,N_1073,N_1369);
nand U1935 (N_1935,N_1004,N_1497);
or U1936 (N_1936,N_1376,N_1424);
or U1937 (N_1937,N_1487,N_1306);
or U1938 (N_1938,N_1360,N_1499);
xnor U1939 (N_1939,N_1226,N_1116);
xnor U1940 (N_1940,N_1395,N_1261);
or U1941 (N_1941,N_1122,N_1178);
nand U1942 (N_1942,N_1141,N_1370);
and U1943 (N_1943,N_1133,N_1253);
nor U1944 (N_1944,N_1452,N_1440);
and U1945 (N_1945,N_1111,N_1169);
and U1946 (N_1946,N_1169,N_1438);
and U1947 (N_1947,N_1266,N_1172);
xnor U1948 (N_1948,N_1394,N_1229);
nand U1949 (N_1949,N_1372,N_1385);
and U1950 (N_1950,N_1479,N_1118);
nand U1951 (N_1951,N_1359,N_1266);
xnor U1952 (N_1952,N_1256,N_1369);
and U1953 (N_1953,N_1369,N_1352);
nor U1954 (N_1954,N_1314,N_1233);
xnor U1955 (N_1955,N_1433,N_1098);
nand U1956 (N_1956,N_1080,N_1393);
xor U1957 (N_1957,N_1173,N_1326);
nand U1958 (N_1958,N_1223,N_1426);
nand U1959 (N_1959,N_1073,N_1354);
nand U1960 (N_1960,N_1436,N_1062);
and U1961 (N_1961,N_1035,N_1202);
and U1962 (N_1962,N_1428,N_1215);
xnor U1963 (N_1963,N_1166,N_1318);
nor U1964 (N_1964,N_1017,N_1096);
nor U1965 (N_1965,N_1427,N_1089);
nor U1966 (N_1966,N_1012,N_1136);
nor U1967 (N_1967,N_1417,N_1065);
nand U1968 (N_1968,N_1132,N_1230);
or U1969 (N_1969,N_1044,N_1168);
nor U1970 (N_1970,N_1196,N_1388);
and U1971 (N_1971,N_1118,N_1235);
nand U1972 (N_1972,N_1049,N_1118);
or U1973 (N_1973,N_1462,N_1444);
nor U1974 (N_1974,N_1068,N_1400);
and U1975 (N_1975,N_1224,N_1033);
or U1976 (N_1976,N_1429,N_1223);
nor U1977 (N_1977,N_1057,N_1060);
or U1978 (N_1978,N_1236,N_1136);
or U1979 (N_1979,N_1149,N_1189);
nand U1980 (N_1980,N_1164,N_1236);
nor U1981 (N_1981,N_1451,N_1139);
and U1982 (N_1982,N_1268,N_1065);
nor U1983 (N_1983,N_1237,N_1116);
or U1984 (N_1984,N_1145,N_1200);
or U1985 (N_1985,N_1019,N_1083);
and U1986 (N_1986,N_1202,N_1438);
and U1987 (N_1987,N_1481,N_1029);
nand U1988 (N_1988,N_1230,N_1266);
nor U1989 (N_1989,N_1405,N_1007);
or U1990 (N_1990,N_1320,N_1039);
nand U1991 (N_1991,N_1021,N_1218);
and U1992 (N_1992,N_1128,N_1145);
or U1993 (N_1993,N_1152,N_1241);
or U1994 (N_1994,N_1108,N_1320);
or U1995 (N_1995,N_1372,N_1028);
nand U1996 (N_1996,N_1397,N_1308);
nor U1997 (N_1997,N_1011,N_1282);
nor U1998 (N_1998,N_1329,N_1120);
nand U1999 (N_1999,N_1399,N_1320);
nor U2000 (N_2000,N_1942,N_1876);
and U2001 (N_2001,N_1561,N_1708);
nand U2002 (N_2002,N_1620,N_1526);
and U2003 (N_2003,N_1555,N_1663);
xnor U2004 (N_2004,N_1732,N_1733);
or U2005 (N_2005,N_1913,N_1553);
nand U2006 (N_2006,N_1627,N_1584);
and U2007 (N_2007,N_1803,N_1673);
and U2008 (N_2008,N_1974,N_1583);
and U2009 (N_2009,N_1925,N_1572);
nor U2010 (N_2010,N_1827,N_1843);
nor U2011 (N_2011,N_1749,N_1657);
or U2012 (N_2012,N_1679,N_1850);
xor U2013 (N_2013,N_1748,N_1886);
or U2014 (N_2014,N_1937,N_1637);
nand U2015 (N_2015,N_1807,N_1841);
nor U2016 (N_2016,N_1743,N_1951);
nor U2017 (N_2017,N_1823,N_1845);
and U2018 (N_2018,N_1912,N_1835);
nor U2019 (N_2019,N_1808,N_1800);
nand U2020 (N_2020,N_1781,N_1576);
nor U2021 (N_2021,N_1938,N_1797);
or U2022 (N_2022,N_1933,N_1779);
and U2023 (N_2023,N_1778,N_1722);
or U2024 (N_2024,N_1972,N_1981);
or U2025 (N_2025,N_1777,N_1692);
nand U2026 (N_2026,N_1944,N_1612);
or U2027 (N_2027,N_1889,N_1780);
nor U2028 (N_2028,N_1606,N_1927);
nor U2029 (N_2029,N_1899,N_1961);
nand U2030 (N_2030,N_1514,N_1546);
or U2031 (N_2031,N_1905,N_1932);
nor U2032 (N_2032,N_1742,N_1615);
nand U2033 (N_2033,N_1669,N_1596);
nand U2034 (N_2034,N_1856,N_1658);
or U2035 (N_2035,N_1616,N_1910);
nor U2036 (N_2036,N_1973,N_1618);
nand U2037 (N_2037,N_1790,N_1826);
nand U2038 (N_2038,N_1577,N_1599);
and U2039 (N_2039,N_1765,N_1967);
nor U2040 (N_2040,N_1502,N_1846);
nor U2041 (N_2041,N_1969,N_1870);
and U2042 (N_2042,N_1821,N_1928);
or U2043 (N_2043,N_1683,N_1725);
nand U2044 (N_2044,N_1784,N_1688);
nor U2045 (N_2045,N_1997,N_1659);
nor U2046 (N_2046,N_1684,N_1594);
and U2047 (N_2047,N_1567,N_1704);
or U2048 (N_2048,N_1875,N_1500);
nor U2049 (N_2049,N_1668,N_1560);
nand U2050 (N_2050,N_1509,N_1697);
nor U2051 (N_2051,N_1963,N_1987);
nand U2052 (N_2052,N_1647,N_1792);
and U2053 (N_2053,N_1517,N_1666);
or U2054 (N_2054,N_1943,N_1745);
and U2055 (N_2055,N_1703,N_1760);
nor U2056 (N_2056,N_1775,N_1686);
or U2057 (N_2057,N_1630,N_1994);
nor U2058 (N_2058,N_1855,N_1885);
nor U2059 (N_2059,N_1590,N_1527);
or U2060 (N_2060,N_1550,N_1603);
and U2061 (N_2061,N_1706,N_1948);
nand U2062 (N_2062,N_1665,N_1662);
xnor U2063 (N_2063,N_1557,N_1702);
nand U2064 (N_2064,N_1985,N_1848);
and U2065 (N_2065,N_1971,N_1626);
nor U2066 (N_2066,N_1709,N_1809);
nor U2067 (N_2067,N_1847,N_1523);
nor U2068 (N_2068,N_1986,N_1674);
or U2069 (N_2069,N_1568,N_1602);
nor U2070 (N_2070,N_1955,N_1975);
or U2071 (N_2071,N_1891,N_1931);
and U2072 (N_2072,N_1920,N_1532);
or U2073 (N_2073,N_1818,N_1656);
nor U2074 (N_2074,N_1866,N_1506);
or U2075 (N_2075,N_1719,N_1670);
nand U2076 (N_2076,N_1549,N_1840);
nor U2077 (N_2077,N_1820,N_1598);
xor U2078 (N_2078,N_1595,N_1877);
or U2079 (N_2079,N_1661,N_1543);
nor U2080 (N_2080,N_1727,N_1879);
nand U2081 (N_2081,N_1785,N_1696);
xnor U2082 (N_2082,N_1976,N_1787);
nor U2083 (N_2083,N_1623,N_1610);
and U2084 (N_2084,N_1832,N_1865);
nor U2085 (N_2085,N_1857,N_1978);
nor U2086 (N_2086,N_1565,N_1611);
nor U2087 (N_2087,N_1767,N_1897);
and U2088 (N_2088,N_1958,N_1746);
xor U2089 (N_2089,N_1581,N_1828);
or U2090 (N_2090,N_1660,N_1833);
nand U2091 (N_2091,N_1540,N_1607);
nor U2092 (N_2092,N_1536,N_1864);
and U2093 (N_2093,N_1890,N_1984);
and U2094 (N_2094,N_1874,N_1597);
or U2095 (N_2095,N_1911,N_1924);
xnor U2096 (N_2096,N_1766,N_1991);
or U2097 (N_2097,N_1632,N_1764);
xor U2098 (N_2098,N_1635,N_1521);
nand U2099 (N_2099,N_1545,N_1654);
nor U2100 (N_2100,N_1628,N_1710);
or U2101 (N_2101,N_1600,N_1844);
and U2102 (N_2102,N_1793,N_1547);
or U2103 (N_2103,N_1965,N_1621);
xor U2104 (N_2104,N_1902,N_1960);
xor U2105 (N_2105,N_1592,N_1634);
nor U2106 (N_2106,N_1556,N_1672);
and U2107 (N_2107,N_1993,N_1728);
nand U2108 (N_2108,N_1798,N_1715);
xor U2109 (N_2109,N_1878,N_1587);
xnor U2110 (N_2110,N_1868,N_1939);
nand U2111 (N_2111,N_1935,N_1511);
nand U2112 (N_2112,N_1713,N_1681);
or U2113 (N_2113,N_1753,N_1735);
nand U2114 (N_2114,N_1842,N_1887);
and U2115 (N_2115,N_1544,N_1513);
or U2116 (N_2116,N_1537,N_1625);
or U2117 (N_2117,N_1528,N_1638);
or U2118 (N_2118,N_1811,N_1921);
xor U2119 (N_2119,N_1664,N_1862);
xor U2120 (N_2120,N_1680,N_1586);
nor U2121 (N_2121,N_1731,N_1677);
or U2122 (N_2122,N_1690,N_1691);
or U2123 (N_2123,N_1786,N_1761);
nor U2124 (N_2124,N_1831,N_1949);
or U2125 (N_2125,N_1916,N_1699);
and U2126 (N_2126,N_1573,N_1946);
and U2127 (N_2127,N_1551,N_1756);
and U2128 (N_2128,N_1508,N_1741);
and U2129 (N_2129,N_1919,N_1996);
and U2130 (N_2130,N_1707,N_1529);
nand U2131 (N_2131,N_1768,N_1542);
or U2132 (N_2132,N_1992,N_1882);
nor U2133 (N_2133,N_1554,N_1929);
nor U2134 (N_2134,N_1701,N_1989);
xor U2135 (N_2135,N_1640,N_1518);
or U2136 (N_2136,N_1738,N_1676);
xor U2137 (N_2137,N_1531,N_1569);
or U2138 (N_2138,N_1729,N_1880);
nand U2139 (N_2139,N_1614,N_1830);
nor U2140 (N_2140,N_1711,N_1525);
nor U2141 (N_2141,N_1754,N_1849);
nand U2142 (N_2142,N_1915,N_1801);
or U2143 (N_2143,N_1533,N_1834);
nor U2144 (N_2144,N_1737,N_1964);
nor U2145 (N_2145,N_1655,N_1613);
nand U2146 (N_2146,N_1788,N_1726);
or U2147 (N_2147,N_1716,N_1783);
nor U2148 (N_2148,N_1636,N_1813);
or U2149 (N_2149,N_1582,N_1789);
nand U2150 (N_2150,N_1947,N_1643);
and U2151 (N_2151,N_1712,N_1755);
nor U2152 (N_2152,N_1646,N_1983);
or U2153 (N_2153,N_1950,N_1854);
or U2154 (N_2154,N_1806,N_1837);
nor U2155 (N_2155,N_1999,N_1622);
or U2156 (N_2156,N_1977,N_1585);
nor U2157 (N_2157,N_1945,N_1757);
nand U2158 (N_2158,N_1575,N_1867);
xnor U2159 (N_2159,N_1570,N_1819);
xnor U2160 (N_2160,N_1970,N_1751);
nand U2161 (N_2161,N_1759,N_1605);
and U2162 (N_2162,N_1534,N_1888);
or U2163 (N_2163,N_1648,N_1530);
xnor U2164 (N_2164,N_1571,N_1678);
and U2165 (N_2165,N_1667,N_1990);
nor U2166 (N_2166,N_1520,N_1956);
nor U2167 (N_2167,N_1802,N_1988);
nand U2168 (N_2168,N_1968,N_1898);
nor U2169 (N_2169,N_1979,N_1805);
and U2170 (N_2170,N_1714,N_1515);
and U2171 (N_2171,N_1700,N_1904);
nand U2172 (N_2172,N_1682,N_1624);
xnor U2173 (N_2173,N_1871,N_1941);
nand U2174 (N_2174,N_1541,N_1724);
and U2175 (N_2175,N_1516,N_1752);
nand U2176 (N_2176,N_1601,N_1895);
or U2177 (N_2177,N_1852,N_1907);
nor U2178 (N_2178,N_1894,N_1860);
or U2179 (N_2179,N_1982,N_1644);
or U2180 (N_2180,N_1559,N_1810);
nor U2181 (N_2181,N_1782,N_1861);
xnor U2182 (N_2182,N_1633,N_1817);
or U2183 (N_2183,N_1859,N_1718);
and U2184 (N_2184,N_1671,N_1934);
nor U2185 (N_2185,N_1685,N_1909);
nor U2186 (N_2186,N_1539,N_1796);
xor U2187 (N_2187,N_1900,N_1825);
or U2188 (N_2188,N_1794,N_1650);
nand U2189 (N_2189,N_1591,N_1892);
nand U2190 (N_2190,N_1853,N_1762);
and U2191 (N_2191,N_1698,N_1799);
or U2192 (N_2192,N_1980,N_1769);
nor U2193 (N_2193,N_1881,N_1908);
or U2194 (N_2194,N_1617,N_1535);
xnor U2195 (N_2195,N_1744,N_1816);
nand U2196 (N_2196,N_1901,N_1524);
or U2197 (N_2197,N_1851,N_1770);
xnor U2198 (N_2198,N_1829,N_1578);
and U2199 (N_2199,N_1548,N_1906);
nand U2200 (N_2200,N_1771,N_1922);
or U2201 (N_2201,N_1593,N_1619);
or U2202 (N_2202,N_1930,N_1812);
nand U2203 (N_2203,N_1940,N_1839);
nor U2204 (N_2204,N_1507,N_1566);
and U2205 (N_2205,N_1730,N_1589);
and U2206 (N_2206,N_1720,N_1649);
and U2207 (N_2207,N_1501,N_1772);
nand U2208 (N_2208,N_1952,N_1629);
or U2209 (N_2209,N_1651,N_1824);
and U2210 (N_2210,N_1740,N_1763);
nand U2211 (N_2211,N_1962,N_1774);
nand U2212 (N_2212,N_1923,N_1563);
or U2213 (N_2213,N_1695,N_1562);
xnor U2214 (N_2214,N_1914,N_1608);
nand U2215 (N_2215,N_1936,N_1675);
nor U2216 (N_2216,N_1773,N_1653);
or U2217 (N_2217,N_1588,N_1995);
and U2218 (N_2218,N_1538,N_1815);
nor U2219 (N_2219,N_1869,N_1747);
xor U2220 (N_2220,N_1893,N_1739);
xnor U2221 (N_2221,N_1953,N_1917);
nor U2222 (N_2222,N_1776,N_1734);
xor U2223 (N_2223,N_1903,N_1791);
or U2224 (N_2224,N_1873,N_1884);
or U2225 (N_2225,N_1512,N_1652);
nand U2226 (N_2226,N_1522,N_1694);
or U2227 (N_2227,N_1564,N_1503);
or U2228 (N_2228,N_1926,N_1858);
nand U2229 (N_2229,N_1957,N_1863);
and U2230 (N_2230,N_1872,N_1689);
nor U2231 (N_2231,N_1579,N_1822);
xnor U2232 (N_2232,N_1750,N_1736);
and U2233 (N_2233,N_1609,N_1574);
nor U2234 (N_2234,N_1896,N_1966);
xnor U2235 (N_2235,N_1954,N_1687);
or U2236 (N_2236,N_1693,N_1804);
nand U2237 (N_2237,N_1721,N_1705);
or U2238 (N_2238,N_1814,N_1631);
xnor U2239 (N_2239,N_1645,N_1504);
and U2240 (N_2240,N_1723,N_1883);
nor U2241 (N_2241,N_1505,N_1558);
nor U2242 (N_2242,N_1552,N_1641);
or U2243 (N_2243,N_1519,N_1639);
and U2244 (N_2244,N_1838,N_1580);
or U2245 (N_2245,N_1717,N_1604);
xnor U2246 (N_2246,N_1959,N_1836);
and U2247 (N_2247,N_1918,N_1642);
and U2248 (N_2248,N_1758,N_1998);
xor U2249 (N_2249,N_1795,N_1510);
xnor U2250 (N_2250,N_1961,N_1697);
and U2251 (N_2251,N_1837,N_1712);
or U2252 (N_2252,N_1845,N_1568);
and U2253 (N_2253,N_1596,N_1616);
xor U2254 (N_2254,N_1739,N_1941);
and U2255 (N_2255,N_1659,N_1878);
and U2256 (N_2256,N_1821,N_1783);
nand U2257 (N_2257,N_1764,N_1783);
nor U2258 (N_2258,N_1818,N_1704);
nor U2259 (N_2259,N_1766,N_1677);
or U2260 (N_2260,N_1710,N_1528);
nor U2261 (N_2261,N_1900,N_1586);
or U2262 (N_2262,N_1738,N_1608);
and U2263 (N_2263,N_1897,N_1534);
nor U2264 (N_2264,N_1763,N_1704);
and U2265 (N_2265,N_1685,N_1942);
nand U2266 (N_2266,N_1518,N_1685);
nor U2267 (N_2267,N_1698,N_1529);
and U2268 (N_2268,N_1887,N_1738);
and U2269 (N_2269,N_1688,N_1625);
nand U2270 (N_2270,N_1584,N_1654);
or U2271 (N_2271,N_1663,N_1881);
nand U2272 (N_2272,N_1921,N_1673);
nand U2273 (N_2273,N_1521,N_1607);
and U2274 (N_2274,N_1800,N_1955);
or U2275 (N_2275,N_1906,N_1911);
and U2276 (N_2276,N_1560,N_1543);
nand U2277 (N_2277,N_1874,N_1616);
nor U2278 (N_2278,N_1904,N_1753);
or U2279 (N_2279,N_1764,N_1768);
nand U2280 (N_2280,N_1705,N_1519);
and U2281 (N_2281,N_1503,N_1796);
nor U2282 (N_2282,N_1617,N_1551);
or U2283 (N_2283,N_1786,N_1536);
and U2284 (N_2284,N_1800,N_1799);
or U2285 (N_2285,N_1669,N_1946);
and U2286 (N_2286,N_1902,N_1981);
or U2287 (N_2287,N_1603,N_1725);
nor U2288 (N_2288,N_1828,N_1539);
nor U2289 (N_2289,N_1809,N_1521);
or U2290 (N_2290,N_1587,N_1721);
nand U2291 (N_2291,N_1776,N_1914);
and U2292 (N_2292,N_1809,N_1654);
nor U2293 (N_2293,N_1524,N_1780);
nand U2294 (N_2294,N_1775,N_1765);
and U2295 (N_2295,N_1677,N_1549);
or U2296 (N_2296,N_1531,N_1645);
nand U2297 (N_2297,N_1889,N_1864);
and U2298 (N_2298,N_1708,N_1950);
nand U2299 (N_2299,N_1991,N_1594);
and U2300 (N_2300,N_1829,N_1523);
and U2301 (N_2301,N_1809,N_1515);
or U2302 (N_2302,N_1982,N_1945);
and U2303 (N_2303,N_1688,N_1657);
nor U2304 (N_2304,N_1765,N_1975);
nor U2305 (N_2305,N_1684,N_1583);
nand U2306 (N_2306,N_1831,N_1511);
and U2307 (N_2307,N_1941,N_1942);
nand U2308 (N_2308,N_1878,N_1813);
or U2309 (N_2309,N_1553,N_1575);
and U2310 (N_2310,N_1852,N_1824);
nor U2311 (N_2311,N_1817,N_1956);
nor U2312 (N_2312,N_1674,N_1945);
nor U2313 (N_2313,N_1986,N_1974);
and U2314 (N_2314,N_1539,N_1865);
nand U2315 (N_2315,N_1547,N_1753);
nand U2316 (N_2316,N_1868,N_1851);
and U2317 (N_2317,N_1576,N_1523);
nand U2318 (N_2318,N_1688,N_1610);
and U2319 (N_2319,N_1868,N_1860);
and U2320 (N_2320,N_1967,N_1583);
nor U2321 (N_2321,N_1578,N_1716);
or U2322 (N_2322,N_1512,N_1525);
nor U2323 (N_2323,N_1834,N_1603);
and U2324 (N_2324,N_1685,N_1694);
and U2325 (N_2325,N_1613,N_1787);
xor U2326 (N_2326,N_1661,N_1560);
and U2327 (N_2327,N_1959,N_1841);
xor U2328 (N_2328,N_1654,N_1691);
or U2329 (N_2329,N_1611,N_1875);
nand U2330 (N_2330,N_1976,N_1738);
nand U2331 (N_2331,N_1764,N_1695);
nor U2332 (N_2332,N_1806,N_1588);
nor U2333 (N_2333,N_1787,N_1767);
or U2334 (N_2334,N_1586,N_1556);
or U2335 (N_2335,N_1998,N_1722);
nand U2336 (N_2336,N_1794,N_1886);
nand U2337 (N_2337,N_1720,N_1865);
nand U2338 (N_2338,N_1954,N_1772);
or U2339 (N_2339,N_1633,N_1975);
or U2340 (N_2340,N_1884,N_1810);
xnor U2341 (N_2341,N_1553,N_1866);
xor U2342 (N_2342,N_1918,N_1954);
and U2343 (N_2343,N_1810,N_1790);
or U2344 (N_2344,N_1722,N_1933);
xor U2345 (N_2345,N_1818,N_1666);
or U2346 (N_2346,N_1771,N_1887);
xnor U2347 (N_2347,N_1522,N_1755);
nand U2348 (N_2348,N_1621,N_1501);
and U2349 (N_2349,N_1641,N_1657);
or U2350 (N_2350,N_1844,N_1662);
or U2351 (N_2351,N_1625,N_1779);
nand U2352 (N_2352,N_1727,N_1604);
xor U2353 (N_2353,N_1781,N_1995);
xnor U2354 (N_2354,N_1671,N_1737);
nor U2355 (N_2355,N_1648,N_1841);
and U2356 (N_2356,N_1828,N_1942);
or U2357 (N_2357,N_1605,N_1774);
nand U2358 (N_2358,N_1583,N_1832);
xor U2359 (N_2359,N_1898,N_1711);
nand U2360 (N_2360,N_1781,N_1599);
nor U2361 (N_2361,N_1538,N_1720);
nor U2362 (N_2362,N_1814,N_1880);
and U2363 (N_2363,N_1993,N_1912);
nand U2364 (N_2364,N_1757,N_1712);
and U2365 (N_2365,N_1500,N_1924);
or U2366 (N_2366,N_1678,N_1982);
nor U2367 (N_2367,N_1907,N_1997);
xnor U2368 (N_2368,N_1536,N_1547);
or U2369 (N_2369,N_1947,N_1613);
or U2370 (N_2370,N_1651,N_1793);
or U2371 (N_2371,N_1757,N_1990);
nor U2372 (N_2372,N_1839,N_1505);
xor U2373 (N_2373,N_1932,N_1706);
and U2374 (N_2374,N_1780,N_1693);
or U2375 (N_2375,N_1727,N_1956);
or U2376 (N_2376,N_1766,N_1559);
nor U2377 (N_2377,N_1827,N_1842);
nand U2378 (N_2378,N_1884,N_1865);
nor U2379 (N_2379,N_1912,N_1956);
and U2380 (N_2380,N_1682,N_1876);
nor U2381 (N_2381,N_1870,N_1851);
and U2382 (N_2382,N_1738,N_1993);
and U2383 (N_2383,N_1635,N_1771);
and U2384 (N_2384,N_1729,N_1564);
xor U2385 (N_2385,N_1771,N_1745);
xor U2386 (N_2386,N_1910,N_1981);
xor U2387 (N_2387,N_1972,N_1754);
and U2388 (N_2388,N_1700,N_1559);
or U2389 (N_2389,N_1829,N_1631);
or U2390 (N_2390,N_1808,N_1846);
or U2391 (N_2391,N_1920,N_1866);
or U2392 (N_2392,N_1674,N_1772);
and U2393 (N_2393,N_1844,N_1732);
nand U2394 (N_2394,N_1821,N_1937);
or U2395 (N_2395,N_1972,N_1909);
and U2396 (N_2396,N_1946,N_1804);
or U2397 (N_2397,N_1638,N_1537);
nor U2398 (N_2398,N_1879,N_1782);
and U2399 (N_2399,N_1757,N_1982);
xor U2400 (N_2400,N_1502,N_1949);
or U2401 (N_2401,N_1524,N_1610);
or U2402 (N_2402,N_1601,N_1853);
and U2403 (N_2403,N_1997,N_1979);
or U2404 (N_2404,N_1911,N_1971);
nand U2405 (N_2405,N_1835,N_1692);
nand U2406 (N_2406,N_1916,N_1717);
and U2407 (N_2407,N_1725,N_1942);
xnor U2408 (N_2408,N_1748,N_1753);
and U2409 (N_2409,N_1822,N_1985);
or U2410 (N_2410,N_1672,N_1821);
and U2411 (N_2411,N_1531,N_1885);
nor U2412 (N_2412,N_1867,N_1699);
nor U2413 (N_2413,N_1655,N_1773);
nand U2414 (N_2414,N_1517,N_1816);
nand U2415 (N_2415,N_1782,N_1908);
or U2416 (N_2416,N_1941,N_1709);
nand U2417 (N_2417,N_1969,N_1600);
and U2418 (N_2418,N_1735,N_1718);
and U2419 (N_2419,N_1922,N_1711);
nor U2420 (N_2420,N_1766,N_1688);
nor U2421 (N_2421,N_1624,N_1638);
nor U2422 (N_2422,N_1708,N_1881);
nor U2423 (N_2423,N_1853,N_1692);
or U2424 (N_2424,N_1919,N_1636);
nor U2425 (N_2425,N_1705,N_1762);
and U2426 (N_2426,N_1713,N_1977);
nand U2427 (N_2427,N_1878,N_1728);
nor U2428 (N_2428,N_1848,N_1999);
nor U2429 (N_2429,N_1665,N_1639);
and U2430 (N_2430,N_1572,N_1866);
or U2431 (N_2431,N_1863,N_1660);
xor U2432 (N_2432,N_1887,N_1519);
or U2433 (N_2433,N_1859,N_1526);
nand U2434 (N_2434,N_1743,N_1935);
or U2435 (N_2435,N_1995,N_1997);
nor U2436 (N_2436,N_1577,N_1647);
and U2437 (N_2437,N_1693,N_1710);
nor U2438 (N_2438,N_1775,N_1678);
xnor U2439 (N_2439,N_1873,N_1568);
and U2440 (N_2440,N_1938,N_1769);
xnor U2441 (N_2441,N_1815,N_1534);
or U2442 (N_2442,N_1988,N_1912);
xnor U2443 (N_2443,N_1848,N_1643);
and U2444 (N_2444,N_1659,N_1636);
or U2445 (N_2445,N_1754,N_1755);
or U2446 (N_2446,N_1743,N_1622);
nor U2447 (N_2447,N_1582,N_1948);
xor U2448 (N_2448,N_1570,N_1514);
and U2449 (N_2449,N_1994,N_1821);
xor U2450 (N_2450,N_1847,N_1972);
nand U2451 (N_2451,N_1974,N_1861);
nor U2452 (N_2452,N_1874,N_1785);
nand U2453 (N_2453,N_1807,N_1523);
or U2454 (N_2454,N_1872,N_1548);
xnor U2455 (N_2455,N_1848,N_1712);
or U2456 (N_2456,N_1595,N_1631);
and U2457 (N_2457,N_1736,N_1876);
xor U2458 (N_2458,N_1760,N_1538);
nor U2459 (N_2459,N_1830,N_1674);
nand U2460 (N_2460,N_1570,N_1709);
nor U2461 (N_2461,N_1713,N_1664);
nor U2462 (N_2462,N_1933,N_1696);
xor U2463 (N_2463,N_1921,N_1716);
nor U2464 (N_2464,N_1851,N_1731);
and U2465 (N_2465,N_1946,N_1615);
and U2466 (N_2466,N_1913,N_1729);
xor U2467 (N_2467,N_1881,N_1746);
nand U2468 (N_2468,N_1967,N_1934);
nand U2469 (N_2469,N_1751,N_1907);
and U2470 (N_2470,N_1916,N_1986);
or U2471 (N_2471,N_1958,N_1985);
and U2472 (N_2472,N_1852,N_1709);
nand U2473 (N_2473,N_1830,N_1737);
nand U2474 (N_2474,N_1568,N_1624);
xnor U2475 (N_2475,N_1619,N_1981);
nand U2476 (N_2476,N_1955,N_1530);
or U2477 (N_2477,N_1834,N_1620);
nand U2478 (N_2478,N_1560,N_1657);
nand U2479 (N_2479,N_1645,N_1886);
nand U2480 (N_2480,N_1526,N_1994);
xnor U2481 (N_2481,N_1845,N_1874);
xor U2482 (N_2482,N_1973,N_1622);
and U2483 (N_2483,N_1745,N_1842);
or U2484 (N_2484,N_1693,N_1599);
or U2485 (N_2485,N_1790,N_1833);
and U2486 (N_2486,N_1937,N_1931);
or U2487 (N_2487,N_1554,N_1847);
nor U2488 (N_2488,N_1854,N_1619);
and U2489 (N_2489,N_1527,N_1898);
nand U2490 (N_2490,N_1945,N_1908);
nor U2491 (N_2491,N_1958,N_1528);
nor U2492 (N_2492,N_1872,N_1943);
xor U2493 (N_2493,N_1964,N_1943);
and U2494 (N_2494,N_1735,N_1944);
xor U2495 (N_2495,N_1799,N_1652);
nor U2496 (N_2496,N_1573,N_1751);
nor U2497 (N_2497,N_1749,N_1807);
xnor U2498 (N_2498,N_1575,N_1957);
and U2499 (N_2499,N_1744,N_1594);
nand U2500 (N_2500,N_2458,N_2031);
nor U2501 (N_2501,N_2067,N_2113);
and U2502 (N_2502,N_2279,N_2392);
nand U2503 (N_2503,N_2312,N_2201);
and U2504 (N_2504,N_2361,N_2047);
and U2505 (N_2505,N_2414,N_2336);
and U2506 (N_2506,N_2075,N_2455);
nor U2507 (N_2507,N_2214,N_2474);
nand U2508 (N_2508,N_2266,N_2190);
nor U2509 (N_2509,N_2415,N_2010);
xor U2510 (N_2510,N_2343,N_2131);
and U2511 (N_2511,N_2486,N_2023);
nor U2512 (N_2512,N_2170,N_2286);
and U2513 (N_2513,N_2435,N_2303);
or U2514 (N_2514,N_2161,N_2387);
or U2515 (N_2515,N_2155,N_2102);
nand U2516 (N_2516,N_2186,N_2055);
nor U2517 (N_2517,N_2080,N_2107);
or U2518 (N_2518,N_2138,N_2088);
nor U2519 (N_2519,N_2175,N_2344);
or U2520 (N_2520,N_2464,N_2142);
and U2521 (N_2521,N_2147,N_2222);
nand U2522 (N_2522,N_2444,N_2041);
nor U2523 (N_2523,N_2158,N_2267);
or U2524 (N_2524,N_2276,N_2469);
and U2525 (N_2525,N_2281,N_2254);
xor U2526 (N_2526,N_2262,N_2367);
and U2527 (N_2527,N_2025,N_2079);
and U2528 (N_2528,N_2283,N_2300);
and U2529 (N_2529,N_2439,N_2449);
nor U2530 (N_2530,N_2438,N_2052);
and U2531 (N_2531,N_2132,N_2410);
nand U2532 (N_2532,N_2016,N_2139);
and U2533 (N_2533,N_2364,N_2021);
xnor U2534 (N_2534,N_2110,N_2363);
xor U2535 (N_2535,N_2362,N_2339);
nand U2536 (N_2536,N_2194,N_2454);
nor U2537 (N_2537,N_2168,N_2076);
or U2538 (N_2538,N_2382,N_2407);
or U2539 (N_2539,N_2360,N_2424);
or U2540 (N_2540,N_2372,N_2174);
and U2541 (N_2541,N_2246,N_2430);
nor U2542 (N_2542,N_2348,N_2263);
and U2543 (N_2543,N_2054,N_2207);
nor U2544 (N_2544,N_2095,N_2251);
xor U2545 (N_2545,N_2056,N_2405);
and U2546 (N_2546,N_2004,N_2200);
xnor U2547 (N_2547,N_2329,N_2077);
nand U2548 (N_2548,N_2386,N_2232);
nor U2549 (N_2549,N_2396,N_2125);
nand U2550 (N_2550,N_2053,N_2146);
nand U2551 (N_2551,N_2479,N_2203);
and U2552 (N_2552,N_2422,N_2176);
and U2553 (N_2553,N_2009,N_2093);
or U2554 (N_2554,N_2179,N_2087);
and U2555 (N_2555,N_2085,N_2099);
or U2556 (N_2556,N_2059,N_2256);
or U2557 (N_2557,N_2224,N_2149);
nor U2558 (N_2558,N_2306,N_2390);
nor U2559 (N_2559,N_2319,N_2243);
nand U2560 (N_2560,N_2325,N_2271);
or U2561 (N_2561,N_2191,N_2463);
xor U2562 (N_2562,N_2480,N_2334);
xor U2563 (N_2563,N_2402,N_2115);
and U2564 (N_2564,N_2062,N_2347);
nand U2565 (N_2565,N_2375,N_2134);
and U2566 (N_2566,N_2202,N_2365);
and U2567 (N_2567,N_2022,N_2321);
xnor U2568 (N_2568,N_2377,N_2288);
nand U2569 (N_2569,N_2145,N_2391);
nand U2570 (N_2570,N_2412,N_2282);
and U2571 (N_2571,N_2488,N_2298);
or U2572 (N_2572,N_2295,N_2225);
nand U2573 (N_2573,N_2130,N_2136);
xor U2574 (N_2574,N_2111,N_2216);
nand U2575 (N_2575,N_2233,N_2236);
nand U2576 (N_2576,N_2495,N_2244);
nor U2577 (N_2577,N_2209,N_2215);
xor U2578 (N_2578,N_2210,N_2466);
xor U2579 (N_2579,N_2451,N_2245);
or U2580 (N_2580,N_2090,N_2416);
nand U2581 (N_2581,N_2484,N_2097);
nand U2582 (N_2582,N_2459,N_2489);
nor U2583 (N_2583,N_2137,N_2205);
nand U2584 (N_2584,N_2148,N_2069);
xnor U2585 (N_2585,N_2177,N_2159);
and U2586 (N_2586,N_2292,N_2061);
or U2587 (N_2587,N_2433,N_2259);
nor U2588 (N_2588,N_2434,N_2036);
or U2589 (N_2589,N_2044,N_2452);
or U2590 (N_2590,N_2101,N_2437);
nor U2591 (N_2591,N_2296,N_2260);
xnor U2592 (N_2592,N_2189,N_2291);
or U2593 (N_2593,N_2230,N_2366);
nand U2594 (N_2594,N_2409,N_2490);
and U2595 (N_2595,N_2257,N_2249);
or U2596 (N_2596,N_2445,N_2252);
and U2597 (N_2597,N_2220,N_2420);
xnor U2598 (N_2598,N_2304,N_2398);
or U2599 (N_2599,N_2326,N_2401);
nor U2600 (N_2600,N_2197,N_2431);
nor U2601 (N_2601,N_2269,N_2065);
xnor U2602 (N_2602,N_2465,N_2185);
and U2603 (N_2603,N_2235,N_2285);
or U2604 (N_2604,N_2178,N_2049);
and U2605 (N_2605,N_2265,N_2423);
and U2606 (N_2606,N_2373,N_2311);
and U2607 (N_2607,N_2460,N_2066);
nor U2608 (N_2608,N_2089,N_2289);
and U2609 (N_2609,N_2337,N_2350);
and U2610 (N_2610,N_2166,N_2184);
xor U2611 (N_2611,N_2003,N_2083);
or U2612 (N_2612,N_2371,N_2331);
nand U2613 (N_2613,N_2019,N_2104);
nor U2614 (N_2614,N_2231,N_2494);
xnor U2615 (N_2615,N_2381,N_2014);
xor U2616 (N_2616,N_2324,N_2314);
nand U2617 (N_2617,N_2007,N_2109);
nand U2618 (N_2618,N_2287,N_2105);
and U2619 (N_2619,N_2499,N_2172);
and U2620 (N_2620,N_2317,N_2394);
and U2621 (N_2621,N_2498,N_2408);
and U2622 (N_2622,N_2073,N_2389);
or U2623 (N_2623,N_2204,N_2310);
and U2624 (N_2624,N_2293,N_2413);
or U2625 (N_2625,N_2448,N_2468);
nand U2626 (N_2626,N_2481,N_2057);
nand U2627 (N_2627,N_2120,N_2229);
nand U2628 (N_2628,N_2164,N_2029);
nor U2629 (N_2629,N_2144,N_2126);
or U2630 (N_2630,N_2253,N_2193);
and U2631 (N_2631,N_2006,N_2264);
xor U2632 (N_2632,N_2116,N_2238);
or U2633 (N_2633,N_2497,N_2342);
nand U2634 (N_2634,N_2313,N_2035);
nand U2635 (N_2635,N_2092,N_2211);
and U2636 (N_2636,N_2273,N_2103);
nor U2637 (N_2637,N_2315,N_2033);
xnor U2638 (N_2638,N_2307,N_2258);
nor U2639 (N_2639,N_2124,N_2040);
or U2640 (N_2640,N_2108,N_2028);
nand U2641 (N_2641,N_2359,N_2404);
nor U2642 (N_2642,N_2240,N_2301);
and U2643 (N_2643,N_2411,N_2376);
or U2644 (N_2644,N_2357,N_2268);
and U2645 (N_2645,N_2309,N_2045);
xor U2646 (N_2646,N_2218,N_2345);
nand U2647 (N_2647,N_2017,N_2050);
nor U2648 (N_2648,N_2385,N_2277);
and U2649 (N_2649,N_2026,N_2081);
nor U2650 (N_2650,N_2058,N_2284);
and U2651 (N_2651,N_2199,N_2123);
or U2652 (N_2652,N_2212,N_2034);
xor U2653 (N_2653,N_2461,N_2426);
xor U2654 (N_2654,N_2106,N_2226);
or U2655 (N_2655,N_2478,N_2340);
nand U2656 (N_2656,N_2368,N_2400);
nor U2657 (N_2657,N_2383,N_2446);
or U2658 (N_2658,N_2280,N_2143);
or U2659 (N_2659,N_2487,N_2012);
and U2660 (N_2660,N_2182,N_2117);
nand U2661 (N_2661,N_2261,N_2173);
nor U2662 (N_2662,N_2121,N_2406);
nand U2663 (N_2663,N_2013,N_2213);
and U2664 (N_2664,N_2346,N_2349);
and U2665 (N_2665,N_2421,N_2043);
nand U2666 (N_2666,N_2418,N_2492);
or U2667 (N_2667,N_2378,N_2316);
nor U2668 (N_2668,N_2395,N_2397);
nand U2669 (N_2669,N_2074,N_2086);
or U2670 (N_2670,N_2154,N_2030);
nor U2671 (N_2671,N_2001,N_2471);
or U2672 (N_2672,N_2447,N_2141);
xnor U2673 (N_2673,N_2039,N_2063);
nand U2674 (N_2674,N_2467,N_2358);
nor U2675 (N_2675,N_2477,N_2096);
and U2676 (N_2676,N_2165,N_2196);
or U2677 (N_2677,N_2082,N_2127);
xnor U2678 (N_2678,N_2078,N_2208);
or U2679 (N_2679,N_2046,N_2308);
nor U2680 (N_2680,N_2442,N_2440);
and U2681 (N_2681,N_2020,N_2171);
nand U2682 (N_2682,N_2234,N_2384);
nand U2683 (N_2683,N_2380,N_2135);
nor U2684 (N_2684,N_2157,N_2228);
or U2685 (N_2685,N_2403,N_2335);
nor U2686 (N_2686,N_2242,N_2169);
and U2687 (N_2687,N_2332,N_2354);
and U2688 (N_2688,N_2094,N_2032);
or U2689 (N_2689,N_2485,N_2217);
nand U2690 (N_2690,N_2162,N_2374);
xnor U2691 (N_2691,N_2187,N_2388);
nor U2692 (N_2692,N_2436,N_2338);
or U2693 (N_2693,N_2473,N_2370);
or U2694 (N_2694,N_2167,N_2156);
nand U2695 (N_2695,N_2432,N_2008);
nor U2696 (N_2696,N_2140,N_2163);
nor U2697 (N_2697,N_2419,N_2493);
or U2698 (N_2698,N_2038,N_2129);
nand U2699 (N_2699,N_2475,N_2491);
nand U2700 (N_2700,N_2318,N_2322);
nand U2701 (N_2701,N_2239,N_2305);
nand U2702 (N_2702,N_2302,N_2027);
nor U2703 (N_2703,N_2018,N_2219);
xnor U2704 (N_2704,N_2071,N_2356);
nand U2705 (N_2705,N_2250,N_2278);
nor U2706 (N_2706,N_2482,N_2122);
xnor U2707 (N_2707,N_2353,N_2294);
or U2708 (N_2708,N_2470,N_2330);
and U2709 (N_2709,N_2206,N_2456);
nor U2710 (N_2710,N_2496,N_2299);
and U2711 (N_2711,N_2457,N_2195);
or U2712 (N_2712,N_2188,N_2084);
nand U2713 (N_2713,N_2011,N_2450);
nor U2714 (N_2714,N_2425,N_2133);
xnor U2715 (N_2715,N_2002,N_2462);
nand U2716 (N_2716,N_2000,N_2112);
or U2717 (N_2717,N_2472,N_2327);
nand U2718 (N_2718,N_2181,N_2221);
or U2719 (N_2719,N_2064,N_2379);
nor U2720 (N_2720,N_2060,N_2150);
or U2721 (N_2721,N_2441,N_2015);
and U2722 (N_2722,N_2152,N_2198);
nor U2723 (N_2723,N_2417,N_2248);
nand U2724 (N_2724,N_2241,N_2429);
or U2725 (N_2725,N_2051,N_2048);
and U2726 (N_2726,N_2070,N_2328);
and U2727 (N_2727,N_2192,N_2355);
nor U2728 (N_2728,N_2270,N_2443);
nand U2729 (N_2729,N_2114,N_2341);
and U2730 (N_2730,N_2223,N_2351);
nor U2731 (N_2731,N_2453,N_2333);
or U2732 (N_2732,N_2042,N_2160);
or U2733 (N_2733,N_2024,N_2275);
nand U2734 (N_2734,N_2428,N_2247);
nor U2735 (N_2735,N_2068,N_2128);
and U2736 (N_2736,N_2399,N_2100);
nand U2737 (N_2737,N_2153,N_2272);
and U2738 (N_2738,N_2369,N_2098);
xor U2739 (N_2739,N_2119,N_2393);
xor U2740 (N_2740,N_2180,N_2352);
nor U2741 (N_2741,N_2151,N_2476);
and U2742 (N_2742,N_2118,N_2037);
or U2743 (N_2743,N_2227,N_2005);
and U2744 (N_2744,N_2091,N_2323);
nor U2745 (N_2745,N_2183,N_2237);
xnor U2746 (N_2746,N_2483,N_2072);
and U2747 (N_2747,N_2255,N_2427);
or U2748 (N_2748,N_2297,N_2320);
nand U2749 (N_2749,N_2290,N_2274);
nand U2750 (N_2750,N_2337,N_2309);
and U2751 (N_2751,N_2348,N_2127);
nor U2752 (N_2752,N_2354,N_2492);
nand U2753 (N_2753,N_2312,N_2206);
nor U2754 (N_2754,N_2101,N_2388);
nand U2755 (N_2755,N_2129,N_2223);
xnor U2756 (N_2756,N_2148,N_2117);
nand U2757 (N_2757,N_2358,N_2362);
xnor U2758 (N_2758,N_2059,N_2012);
or U2759 (N_2759,N_2040,N_2166);
nor U2760 (N_2760,N_2413,N_2026);
nand U2761 (N_2761,N_2154,N_2203);
xnor U2762 (N_2762,N_2343,N_2214);
nor U2763 (N_2763,N_2284,N_2010);
and U2764 (N_2764,N_2145,N_2141);
nand U2765 (N_2765,N_2430,N_2405);
and U2766 (N_2766,N_2453,N_2193);
and U2767 (N_2767,N_2108,N_2366);
nand U2768 (N_2768,N_2319,N_2140);
nand U2769 (N_2769,N_2079,N_2364);
nor U2770 (N_2770,N_2099,N_2267);
nand U2771 (N_2771,N_2268,N_2464);
or U2772 (N_2772,N_2211,N_2216);
xnor U2773 (N_2773,N_2098,N_2339);
nor U2774 (N_2774,N_2274,N_2394);
nor U2775 (N_2775,N_2085,N_2332);
nor U2776 (N_2776,N_2174,N_2377);
and U2777 (N_2777,N_2283,N_2090);
xor U2778 (N_2778,N_2459,N_2384);
nor U2779 (N_2779,N_2386,N_2468);
xnor U2780 (N_2780,N_2339,N_2337);
nor U2781 (N_2781,N_2484,N_2274);
or U2782 (N_2782,N_2333,N_2347);
xor U2783 (N_2783,N_2360,N_2164);
nand U2784 (N_2784,N_2131,N_2475);
or U2785 (N_2785,N_2346,N_2229);
nand U2786 (N_2786,N_2062,N_2318);
nor U2787 (N_2787,N_2439,N_2377);
nor U2788 (N_2788,N_2456,N_2256);
nor U2789 (N_2789,N_2260,N_2343);
and U2790 (N_2790,N_2096,N_2253);
nand U2791 (N_2791,N_2424,N_2345);
nand U2792 (N_2792,N_2010,N_2337);
and U2793 (N_2793,N_2322,N_2136);
xor U2794 (N_2794,N_2030,N_2457);
or U2795 (N_2795,N_2224,N_2153);
nor U2796 (N_2796,N_2122,N_2028);
nand U2797 (N_2797,N_2459,N_2303);
and U2798 (N_2798,N_2444,N_2485);
nor U2799 (N_2799,N_2283,N_2350);
nand U2800 (N_2800,N_2213,N_2163);
or U2801 (N_2801,N_2174,N_2055);
nand U2802 (N_2802,N_2154,N_2393);
nand U2803 (N_2803,N_2346,N_2153);
or U2804 (N_2804,N_2271,N_2057);
nand U2805 (N_2805,N_2014,N_2282);
nor U2806 (N_2806,N_2244,N_2476);
or U2807 (N_2807,N_2104,N_2189);
nand U2808 (N_2808,N_2307,N_2297);
and U2809 (N_2809,N_2088,N_2020);
nand U2810 (N_2810,N_2033,N_2165);
nor U2811 (N_2811,N_2033,N_2442);
or U2812 (N_2812,N_2032,N_2119);
or U2813 (N_2813,N_2381,N_2252);
nor U2814 (N_2814,N_2311,N_2482);
nand U2815 (N_2815,N_2400,N_2147);
or U2816 (N_2816,N_2076,N_2151);
nand U2817 (N_2817,N_2395,N_2257);
nor U2818 (N_2818,N_2289,N_2219);
or U2819 (N_2819,N_2051,N_2067);
nor U2820 (N_2820,N_2460,N_2196);
or U2821 (N_2821,N_2220,N_2154);
and U2822 (N_2822,N_2359,N_2204);
nand U2823 (N_2823,N_2368,N_2449);
and U2824 (N_2824,N_2420,N_2117);
nor U2825 (N_2825,N_2332,N_2070);
or U2826 (N_2826,N_2332,N_2382);
nor U2827 (N_2827,N_2425,N_2267);
nand U2828 (N_2828,N_2150,N_2346);
nor U2829 (N_2829,N_2427,N_2327);
nor U2830 (N_2830,N_2281,N_2305);
and U2831 (N_2831,N_2036,N_2320);
nand U2832 (N_2832,N_2424,N_2398);
and U2833 (N_2833,N_2009,N_2247);
xnor U2834 (N_2834,N_2271,N_2053);
or U2835 (N_2835,N_2119,N_2090);
xor U2836 (N_2836,N_2095,N_2216);
or U2837 (N_2837,N_2345,N_2182);
nand U2838 (N_2838,N_2141,N_2306);
or U2839 (N_2839,N_2191,N_2285);
nand U2840 (N_2840,N_2358,N_2407);
and U2841 (N_2841,N_2325,N_2398);
nand U2842 (N_2842,N_2112,N_2455);
or U2843 (N_2843,N_2285,N_2375);
xor U2844 (N_2844,N_2359,N_2465);
nor U2845 (N_2845,N_2155,N_2239);
nand U2846 (N_2846,N_2088,N_2351);
nand U2847 (N_2847,N_2192,N_2025);
nand U2848 (N_2848,N_2204,N_2153);
xnor U2849 (N_2849,N_2151,N_2090);
nor U2850 (N_2850,N_2324,N_2241);
and U2851 (N_2851,N_2413,N_2182);
or U2852 (N_2852,N_2244,N_2188);
nand U2853 (N_2853,N_2356,N_2397);
nand U2854 (N_2854,N_2204,N_2324);
or U2855 (N_2855,N_2388,N_2037);
or U2856 (N_2856,N_2319,N_2185);
nor U2857 (N_2857,N_2235,N_2430);
nor U2858 (N_2858,N_2088,N_2116);
xnor U2859 (N_2859,N_2339,N_2010);
nor U2860 (N_2860,N_2478,N_2217);
nor U2861 (N_2861,N_2039,N_2282);
and U2862 (N_2862,N_2397,N_2179);
and U2863 (N_2863,N_2205,N_2089);
nor U2864 (N_2864,N_2440,N_2431);
and U2865 (N_2865,N_2234,N_2099);
nor U2866 (N_2866,N_2064,N_2477);
nor U2867 (N_2867,N_2222,N_2497);
or U2868 (N_2868,N_2331,N_2238);
and U2869 (N_2869,N_2478,N_2297);
xor U2870 (N_2870,N_2091,N_2482);
xnor U2871 (N_2871,N_2451,N_2002);
and U2872 (N_2872,N_2134,N_2085);
nand U2873 (N_2873,N_2073,N_2187);
or U2874 (N_2874,N_2250,N_2216);
or U2875 (N_2875,N_2121,N_2093);
or U2876 (N_2876,N_2373,N_2423);
or U2877 (N_2877,N_2219,N_2363);
nor U2878 (N_2878,N_2409,N_2305);
nand U2879 (N_2879,N_2204,N_2480);
nand U2880 (N_2880,N_2004,N_2175);
nor U2881 (N_2881,N_2442,N_2128);
and U2882 (N_2882,N_2459,N_2191);
nor U2883 (N_2883,N_2011,N_2048);
or U2884 (N_2884,N_2384,N_2288);
and U2885 (N_2885,N_2101,N_2224);
nand U2886 (N_2886,N_2305,N_2204);
nand U2887 (N_2887,N_2426,N_2221);
nand U2888 (N_2888,N_2155,N_2013);
xnor U2889 (N_2889,N_2021,N_2469);
and U2890 (N_2890,N_2189,N_2108);
or U2891 (N_2891,N_2157,N_2446);
and U2892 (N_2892,N_2437,N_2380);
nor U2893 (N_2893,N_2492,N_2275);
nand U2894 (N_2894,N_2251,N_2031);
nand U2895 (N_2895,N_2429,N_2159);
nand U2896 (N_2896,N_2452,N_2304);
or U2897 (N_2897,N_2440,N_2198);
nor U2898 (N_2898,N_2343,N_2495);
nand U2899 (N_2899,N_2115,N_2015);
nand U2900 (N_2900,N_2126,N_2014);
or U2901 (N_2901,N_2035,N_2300);
and U2902 (N_2902,N_2331,N_2457);
nand U2903 (N_2903,N_2075,N_2226);
nand U2904 (N_2904,N_2450,N_2081);
and U2905 (N_2905,N_2264,N_2064);
xnor U2906 (N_2906,N_2175,N_2341);
nor U2907 (N_2907,N_2206,N_2210);
nand U2908 (N_2908,N_2279,N_2332);
or U2909 (N_2909,N_2464,N_2128);
nand U2910 (N_2910,N_2445,N_2154);
nor U2911 (N_2911,N_2131,N_2018);
nand U2912 (N_2912,N_2429,N_2497);
nor U2913 (N_2913,N_2361,N_2249);
nand U2914 (N_2914,N_2375,N_2450);
or U2915 (N_2915,N_2451,N_2321);
xor U2916 (N_2916,N_2067,N_2275);
nor U2917 (N_2917,N_2322,N_2094);
and U2918 (N_2918,N_2008,N_2363);
nand U2919 (N_2919,N_2170,N_2412);
nor U2920 (N_2920,N_2335,N_2478);
nand U2921 (N_2921,N_2186,N_2083);
or U2922 (N_2922,N_2130,N_2274);
nor U2923 (N_2923,N_2197,N_2030);
nand U2924 (N_2924,N_2417,N_2055);
nand U2925 (N_2925,N_2167,N_2182);
or U2926 (N_2926,N_2369,N_2161);
or U2927 (N_2927,N_2447,N_2273);
or U2928 (N_2928,N_2400,N_2354);
and U2929 (N_2929,N_2392,N_2340);
nand U2930 (N_2930,N_2187,N_2474);
or U2931 (N_2931,N_2271,N_2368);
nand U2932 (N_2932,N_2268,N_2226);
or U2933 (N_2933,N_2481,N_2050);
and U2934 (N_2934,N_2202,N_2263);
nor U2935 (N_2935,N_2310,N_2248);
and U2936 (N_2936,N_2095,N_2464);
or U2937 (N_2937,N_2271,N_2366);
nand U2938 (N_2938,N_2492,N_2318);
nor U2939 (N_2939,N_2440,N_2141);
nand U2940 (N_2940,N_2254,N_2441);
nand U2941 (N_2941,N_2230,N_2319);
or U2942 (N_2942,N_2498,N_2157);
or U2943 (N_2943,N_2018,N_2420);
and U2944 (N_2944,N_2428,N_2392);
nand U2945 (N_2945,N_2331,N_2144);
and U2946 (N_2946,N_2067,N_2358);
nand U2947 (N_2947,N_2242,N_2147);
nand U2948 (N_2948,N_2124,N_2033);
or U2949 (N_2949,N_2242,N_2065);
nor U2950 (N_2950,N_2474,N_2079);
nor U2951 (N_2951,N_2185,N_2373);
xor U2952 (N_2952,N_2252,N_2485);
nor U2953 (N_2953,N_2207,N_2050);
nand U2954 (N_2954,N_2087,N_2249);
or U2955 (N_2955,N_2451,N_2059);
xnor U2956 (N_2956,N_2220,N_2324);
nand U2957 (N_2957,N_2319,N_2481);
nor U2958 (N_2958,N_2490,N_2134);
or U2959 (N_2959,N_2352,N_2247);
and U2960 (N_2960,N_2067,N_2298);
nor U2961 (N_2961,N_2098,N_2138);
nand U2962 (N_2962,N_2062,N_2473);
and U2963 (N_2963,N_2043,N_2305);
or U2964 (N_2964,N_2035,N_2120);
nor U2965 (N_2965,N_2240,N_2335);
or U2966 (N_2966,N_2111,N_2141);
nor U2967 (N_2967,N_2065,N_2010);
xor U2968 (N_2968,N_2074,N_2250);
nand U2969 (N_2969,N_2430,N_2389);
nor U2970 (N_2970,N_2124,N_2270);
nor U2971 (N_2971,N_2108,N_2255);
and U2972 (N_2972,N_2358,N_2232);
and U2973 (N_2973,N_2164,N_2313);
and U2974 (N_2974,N_2446,N_2491);
and U2975 (N_2975,N_2169,N_2303);
and U2976 (N_2976,N_2461,N_2047);
or U2977 (N_2977,N_2173,N_2461);
nor U2978 (N_2978,N_2184,N_2452);
or U2979 (N_2979,N_2446,N_2087);
nor U2980 (N_2980,N_2061,N_2426);
or U2981 (N_2981,N_2114,N_2256);
xnor U2982 (N_2982,N_2184,N_2235);
and U2983 (N_2983,N_2120,N_2065);
and U2984 (N_2984,N_2253,N_2079);
or U2985 (N_2985,N_2360,N_2405);
and U2986 (N_2986,N_2029,N_2256);
and U2987 (N_2987,N_2320,N_2420);
or U2988 (N_2988,N_2082,N_2344);
or U2989 (N_2989,N_2213,N_2374);
or U2990 (N_2990,N_2488,N_2047);
or U2991 (N_2991,N_2087,N_2340);
nor U2992 (N_2992,N_2112,N_2195);
nor U2993 (N_2993,N_2101,N_2331);
xnor U2994 (N_2994,N_2343,N_2113);
and U2995 (N_2995,N_2307,N_2207);
or U2996 (N_2996,N_2195,N_2012);
nand U2997 (N_2997,N_2153,N_2326);
nand U2998 (N_2998,N_2062,N_2477);
xnor U2999 (N_2999,N_2160,N_2398);
nand UO_0 (O_0,N_2577,N_2659);
nor UO_1 (O_1,N_2953,N_2762);
or UO_2 (O_2,N_2984,N_2714);
nand UO_3 (O_3,N_2656,N_2956);
xor UO_4 (O_4,N_2771,N_2825);
nor UO_5 (O_5,N_2649,N_2754);
nand UO_6 (O_6,N_2860,N_2963);
and UO_7 (O_7,N_2863,N_2789);
nor UO_8 (O_8,N_2783,N_2981);
nand UO_9 (O_9,N_2880,N_2598);
and UO_10 (O_10,N_2922,N_2925);
nor UO_11 (O_11,N_2503,N_2615);
nor UO_12 (O_12,N_2988,N_2892);
or UO_13 (O_13,N_2655,N_2673);
xnor UO_14 (O_14,N_2745,N_2926);
and UO_15 (O_15,N_2704,N_2870);
or UO_16 (O_16,N_2816,N_2835);
or UO_17 (O_17,N_2928,N_2998);
or UO_18 (O_18,N_2980,N_2944);
and UO_19 (O_19,N_2541,N_2588);
and UO_20 (O_20,N_2524,N_2942);
and UO_21 (O_21,N_2951,N_2930);
or UO_22 (O_22,N_2778,N_2691);
xnor UO_23 (O_23,N_2583,N_2900);
nor UO_24 (O_24,N_2635,N_2905);
or UO_25 (O_25,N_2525,N_2943);
nor UO_26 (O_26,N_2641,N_2726);
and UO_27 (O_27,N_2558,N_2913);
or UO_28 (O_28,N_2937,N_2510);
nor UO_29 (O_29,N_2580,N_2823);
or UO_30 (O_30,N_2869,N_2872);
xor UO_31 (O_31,N_2533,N_2651);
or UO_32 (O_32,N_2518,N_2740);
and UO_33 (O_33,N_2903,N_2758);
nand UO_34 (O_34,N_2570,N_2698);
nor UO_35 (O_35,N_2877,N_2974);
or UO_36 (O_36,N_2562,N_2677);
nand UO_37 (O_37,N_2664,N_2927);
nor UO_38 (O_38,N_2883,N_2831);
xor UO_39 (O_39,N_2543,N_2808);
or UO_40 (O_40,N_2934,N_2648);
nand UO_41 (O_41,N_2569,N_2993);
nand UO_42 (O_42,N_2721,N_2871);
xnor UO_43 (O_43,N_2520,N_2837);
nand UO_44 (O_44,N_2897,N_2896);
or UO_45 (O_45,N_2895,N_2989);
nor UO_46 (O_46,N_2550,N_2700);
nand UO_47 (O_47,N_2765,N_2555);
or UO_48 (O_48,N_2800,N_2646);
nor UO_49 (O_49,N_2731,N_2626);
and UO_50 (O_50,N_2798,N_2846);
nor UO_51 (O_51,N_2578,N_2878);
nor UO_52 (O_52,N_2889,N_2966);
xnor UO_53 (O_53,N_2729,N_2633);
or UO_54 (O_54,N_2713,N_2637);
nor UO_55 (O_55,N_2694,N_2645);
nor UO_56 (O_56,N_2792,N_2914);
or UO_57 (O_57,N_2596,N_2764);
xor UO_58 (O_58,N_2589,N_2730);
nor UO_59 (O_59,N_2643,N_2805);
nor UO_60 (O_60,N_2938,N_2611);
and UO_61 (O_61,N_2737,N_2865);
nor UO_62 (O_62,N_2920,N_2960);
and UO_63 (O_63,N_2755,N_2716);
and UO_64 (O_64,N_2886,N_2601);
nor UO_65 (O_65,N_2667,N_2513);
or UO_66 (O_66,N_2782,N_2665);
nand UO_67 (O_67,N_2672,N_2802);
nor UO_68 (O_68,N_2618,N_2881);
and UO_69 (O_69,N_2811,N_2662);
xor UO_70 (O_70,N_2723,N_2906);
and UO_71 (O_71,N_2748,N_2508);
nor UO_72 (O_72,N_2709,N_2600);
xnor UO_73 (O_73,N_2627,N_2738);
nand UO_74 (O_74,N_2838,N_2819);
nand UO_75 (O_75,N_2733,N_2606);
nand UO_76 (O_76,N_2822,N_2706);
and UO_77 (O_77,N_2749,N_2836);
and UO_78 (O_78,N_2623,N_2750);
nand UO_79 (O_79,N_2540,N_2609);
nor UO_80 (O_80,N_2931,N_2674);
or UO_81 (O_81,N_2887,N_2506);
or UO_82 (O_82,N_2712,N_2683);
nand UO_83 (O_83,N_2610,N_2532);
or UO_84 (O_84,N_2553,N_2557);
or UO_85 (O_85,N_2638,N_2582);
nand UO_86 (O_86,N_2791,N_2923);
xor UO_87 (O_87,N_2597,N_2720);
and UO_88 (O_88,N_2932,N_2899);
nand UO_89 (O_89,N_2631,N_2797);
and UO_90 (O_90,N_2781,N_2692);
nand UO_91 (O_91,N_2519,N_2718);
or UO_92 (O_92,N_2912,N_2528);
or UO_93 (O_93,N_2563,N_2741);
nand UO_94 (O_94,N_2780,N_2617);
nand UO_95 (O_95,N_2768,N_2565);
or UO_96 (O_96,N_2546,N_2788);
nor UO_97 (O_97,N_2948,N_2708);
and UO_98 (O_98,N_2814,N_2843);
xor UO_99 (O_99,N_2873,N_2803);
and UO_100 (O_100,N_2702,N_2852);
nand UO_101 (O_101,N_2773,N_2859);
and UO_102 (O_102,N_2972,N_2605);
or UO_103 (O_103,N_2977,N_2595);
nand UO_104 (O_104,N_2751,N_2855);
and UO_105 (O_105,N_2534,N_2907);
and UO_106 (O_106,N_2894,N_2940);
nand UO_107 (O_107,N_2945,N_2879);
nand UO_108 (O_108,N_2522,N_2675);
nor UO_109 (O_109,N_2535,N_2959);
nor UO_110 (O_110,N_2970,N_2584);
nor UO_111 (O_111,N_2766,N_2770);
nand UO_112 (O_112,N_2647,N_2629);
nor UO_113 (O_113,N_2893,N_2552);
nand UO_114 (O_114,N_2613,N_2918);
nand UO_115 (O_115,N_2501,N_2668);
xnor UO_116 (O_116,N_2875,N_2538);
and UO_117 (O_117,N_2979,N_2957);
or UO_118 (O_118,N_2884,N_2854);
nand UO_119 (O_119,N_2901,N_2946);
and UO_120 (O_120,N_2747,N_2985);
and UO_121 (O_121,N_2616,N_2642);
or UO_122 (O_122,N_2703,N_2566);
or UO_123 (O_123,N_2699,N_2511);
nor UO_124 (O_124,N_2581,N_2514);
and UO_125 (O_125,N_2560,N_2801);
and UO_126 (O_126,N_2933,N_2834);
nor UO_127 (O_127,N_2844,N_2604);
nor UO_128 (O_128,N_2634,N_2815);
nor UO_129 (O_129,N_2982,N_2971);
nand UO_130 (O_130,N_2504,N_2573);
nand UO_131 (O_131,N_2688,N_2556);
nand UO_132 (O_132,N_2742,N_2575);
nand UO_133 (O_133,N_2572,N_2515);
or UO_134 (O_134,N_2902,N_2696);
or UO_135 (O_135,N_2856,N_2898);
nor UO_136 (O_136,N_2746,N_2772);
or UO_137 (O_137,N_2987,N_2763);
or UO_138 (O_138,N_2628,N_2710);
nor UO_139 (O_139,N_2996,N_2544);
and UO_140 (O_140,N_2851,N_2545);
nor UO_141 (O_141,N_2779,N_2705);
or UO_142 (O_142,N_2752,N_2568);
or UO_143 (O_143,N_2630,N_2796);
xor UO_144 (O_144,N_2861,N_2711);
or UO_145 (O_145,N_2795,N_2950);
or UO_146 (O_146,N_2827,N_2594);
xor UO_147 (O_147,N_2587,N_2728);
nor UO_148 (O_148,N_2916,N_2840);
or UO_149 (O_149,N_2882,N_2567);
and UO_150 (O_150,N_2991,N_2636);
nand UO_151 (O_151,N_2576,N_2620);
and UO_152 (O_152,N_2579,N_2958);
nor UO_153 (O_153,N_2697,N_2727);
nand UO_154 (O_154,N_2978,N_2690);
and UO_155 (O_155,N_2813,N_2622);
or UO_156 (O_156,N_2919,N_2862);
nor UO_157 (O_157,N_2607,N_2810);
xnor UO_158 (O_158,N_2969,N_2857);
nor UO_159 (O_159,N_2640,N_2592);
nand UO_160 (O_160,N_2736,N_2756);
nand UO_161 (O_161,N_2955,N_2542);
or UO_162 (O_162,N_2509,N_2909);
xnor UO_163 (O_163,N_2602,N_2548);
xor UO_164 (O_164,N_2890,N_2876);
or UO_165 (O_165,N_2968,N_2821);
or UO_166 (O_166,N_2841,N_2701);
and UO_167 (O_167,N_2686,N_2830);
and UO_168 (O_168,N_2849,N_2826);
nor UO_169 (O_169,N_2949,N_2654);
nor UO_170 (O_170,N_2910,N_2537);
and UO_171 (O_171,N_2868,N_2523);
xor UO_172 (O_172,N_2531,N_2561);
and UO_173 (O_173,N_2660,N_2512);
and UO_174 (O_174,N_2885,N_2767);
nor UO_175 (O_175,N_2888,N_2739);
nor UO_176 (O_176,N_2769,N_2536);
or UO_177 (O_177,N_2715,N_2551);
or UO_178 (O_178,N_2695,N_2812);
or UO_179 (O_179,N_2936,N_2725);
xor UO_180 (O_180,N_2829,N_2842);
or UO_181 (O_181,N_2624,N_2809);
or UO_182 (O_182,N_2554,N_2921);
xnor UO_183 (O_183,N_2586,N_2612);
or UO_184 (O_184,N_2599,N_2941);
xnor UO_185 (O_185,N_2952,N_2965);
and UO_186 (O_186,N_2845,N_2818);
or UO_187 (O_187,N_2824,N_2983);
xnor UO_188 (O_188,N_2853,N_2679);
nor UO_189 (O_189,N_2687,N_2625);
or UO_190 (O_190,N_2847,N_2593);
or UO_191 (O_191,N_2929,N_2915);
xor UO_192 (O_192,N_2743,N_2689);
nand UO_193 (O_193,N_2759,N_2547);
nor UO_194 (O_194,N_2676,N_2500);
nor UO_195 (O_195,N_2794,N_2817);
or UO_196 (O_196,N_2777,N_2775);
nand UO_197 (O_197,N_2574,N_2517);
xor UO_198 (O_198,N_2776,N_2526);
or UO_199 (O_199,N_2657,N_2680);
or UO_200 (O_200,N_2874,N_2760);
nor UO_201 (O_201,N_2539,N_2924);
nand UO_202 (O_202,N_2935,N_2585);
nor UO_203 (O_203,N_2828,N_2505);
nand UO_204 (O_204,N_2799,N_2911);
xor UO_205 (O_205,N_2790,N_2858);
nor UO_206 (O_206,N_2653,N_2564);
or UO_207 (O_207,N_2848,N_2619);
nor UO_208 (O_208,N_2990,N_2986);
nor UO_209 (O_209,N_2939,N_2785);
and UO_210 (O_210,N_2832,N_2724);
and UO_211 (O_211,N_2682,N_2632);
nor UO_212 (O_212,N_2804,N_2529);
or UO_213 (O_213,N_2549,N_2973);
and UO_214 (O_214,N_2908,N_2820);
xor UO_215 (O_215,N_2644,N_2994);
nor UO_216 (O_216,N_2850,N_2904);
nand UO_217 (O_217,N_2793,N_2867);
or UO_218 (O_218,N_2962,N_2717);
nor UO_219 (O_219,N_2681,N_2693);
nor UO_220 (O_220,N_2707,N_2976);
nand UO_221 (O_221,N_2995,N_2559);
or UO_222 (O_222,N_2590,N_2761);
nand UO_223 (O_223,N_2744,N_2608);
nand UO_224 (O_224,N_2685,N_2722);
or UO_225 (O_225,N_2521,N_2917);
and UO_226 (O_226,N_2735,N_2571);
xor UO_227 (O_227,N_2786,N_2866);
nor UO_228 (O_228,N_2734,N_2753);
and UO_229 (O_229,N_2621,N_2891);
nor UO_230 (O_230,N_2719,N_2954);
nand UO_231 (O_231,N_2975,N_2992);
or UO_232 (O_232,N_2516,N_2757);
xnor UO_233 (O_233,N_2530,N_2678);
and UO_234 (O_234,N_2671,N_2999);
or UO_235 (O_235,N_2507,N_2603);
nand UO_236 (O_236,N_2784,N_2807);
or UO_237 (O_237,N_2591,N_2669);
or UO_238 (O_238,N_2658,N_2774);
xnor UO_239 (O_239,N_2639,N_2652);
or UO_240 (O_240,N_2997,N_2839);
nand UO_241 (O_241,N_2666,N_2961);
nand UO_242 (O_242,N_2806,N_2947);
nor UO_243 (O_243,N_2833,N_2670);
nor UO_244 (O_244,N_2964,N_2864);
nor UO_245 (O_245,N_2684,N_2614);
and UO_246 (O_246,N_2650,N_2787);
and UO_247 (O_247,N_2502,N_2732);
xor UO_248 (O_248,N_2967,N_2527);
and UO_249 (O_249,N_2661,N_2663);
nor UO_250 (O_250,N_2588,N_2626);
or UO_251 (O_251,N_2864,N_2669);
or UO_252 (O_252,N_2870,N_2732);
xnor UO_253 (O_253,N_2817,N_2842);
nand UO_254 (O_254,N_2912,N_2964);
xnor UO_255 (O_255,N_2511,N_2714);
nor UO_256 (O_256,N_2537,N_2784);
and UO_257 (O_257,N_2792,N_2692);
or UO_258 (O_258,N_2870,N_2919);
or UO_259 (O_259,N_2839,N_2656);
xor UO_260 (O_260,N_2542,N_2895);
nand UO_261 (O_261,N_2800,N_2671);
or UO_262 (O_262,N_2617,N_2958);
or UO_263 (O_263,N_2841,N_2959);
xnor UO_264 (O_264,N_2576,N_2715);
nand UO_265 (O_265,N_2683,N_2582);
nor UO_266 (O_266,N_2938,N_2721);
nand UO_267 (O_267,N_2857,N_2882);
and UO_268 (O_268,N_2618,N_2581);
and UO_269 (O_269,N_2590,N_2731);
nand UO_270 (O_270,N_2922,N_2753);
nand UO_271 (O_271,N_2823,N_2953);
nor UO_272 (O_272,N_2879,N_2521);
or UO_273 (O_273,N_2552,N_2619);
and UO_274 (O_274,N_2944,N_2869);
xnor UO_275 (O_275,N_2843,N_2740);
nor UO_276 (O_276,N_2679,N_2906);
or UO_277 (O_277,N_2636,N_2690);
nor UO_278 (O_278,N_2535,N_2788);
xor UO_279 (O_279,N_2767,N_2722);
or UO_280 (O_280,N_2776,N_2722);
and UO_281 (O_281,N_2875,N_2821);
xor UO_282 (O_282,N_2630,N_2905);
and UO_283 (O_283,N_2966,N_2860);
nand UO_284 (O_284,N_2557,N_2587);
nand UO_285 (O_285,N_2530,N_2799);
and UO_286 (O_286,N_2974,N_2907);
nand UO_287 (O_287,N_2920,N_2831);
or UO_288 (O_288,N_2520,N_2693);
nand UO_289 (O_289,N_2791,N_2832);
and UO_290 (O_290,N_2685,N_2889);
or UO_291 (O_291,N_2952,N_2551);
nand UO_292 (O_292,N_2597,N_2978);
and UO_293 (O_293,N_2967,N_2510);
nor UO_294 (O_294,N_2784,N_2977);
nand UO_295 (O_295,N_2597,N_2999);
nand UO_296 (O_296,N_2760,N_2902);
nor UO_297 (O_297,N_2575,N_2619);
or UO_298 (O_298,N_2727,N_2964);
nor UO_299 (O_299,N_2643,N_2683);
or UO_300 (O_300,N_2712,N_2860);
or UO_301 (O_301,N_2967,N_2575);
and UO_302 (O_302,N_2642,N_2826);
and UO_303 (O_303,N_2975,N_2971);
xor UO_304 (O_304,N_2527,N_2678);
nand UO_305 (O_305,N_2932,N_2537);
xnor UO_306 (O_306,N_2557,N_2921);
or UO_307 (O_307,N_2546,N_2557);
xor UO_308 (O_308,N_2827,N_2954);
and UO_309 (O_309,N_2604,N_2921);
and UO_310 (O_310,N_2537,N_2658);
nand UO_311 (O_311,N_2851,N_2899);
nor UO_312 (O_312,N_2686,N_2550);
xnor UO_313 (O_313,N_2784,N_2599);
and UO_314 (O_314,N_2745,N_2585);
and UO_315 (O_315,N_2839,N_2668);
and UO_316 (O_316,N_2852,N_2678);
or UO_317 (O_317,N_2983,N_2573);
and UO_318 (O_318,N_2760,N_2711);
or UO_319 (O_319,N_2565,N_2691);
nor UO_320 (O_320,N_2804,N_2594);
nor UO_321 (O_321,N_2907,N_2727);
or UO_322 (O_322,N_2850,N_2742);
nand UO_323 (O_323,N_2889,N_2542);
nor UO_324 (O_324,N_2852,N_2669);
and UO_325 (O_325,N_2792,N_2547);
xor UO_326 (O_326,N_2802,N_2741);
nand UO_327 (O_327,N_2940,N_2893);
xnor UO_328 (O_328,N_2810,N_2857);
and UO_329 (O_329,N_2716,N_2614);
or UO_330 (O_330,N_2584,N_2775);
and UO_331 (O_331,N_2735,N_2997);
or UO_332 (O_332,N_2590,N_2926);
nor UO_333 (O_333,N_2665,N_2808);
xnor UO_334 (O_334,N_2968,N_2644);
nand UO_335 (O_335,N_2580,N_2547);
or UO_336 (O_336,N_2974,N_2868);
and UO_337 (O_337,N_2852,N_2770);
or UO_338 (O_338,N_2969,N_2793);
or UO_339 (O_339,N_2948,N_2724);
or UO_340 (O_340,N_2822,N_2635);
nor UO_341 (O_341,N_2661,N_2933);
nor UO_342 (O_342,N_2623,N_2811);
and UO_343 (O_343,N_2591,N_2925);
xor UO_344 (O_344,N_2862,N_2551);
nor UO_345 (O_345,N_2988,N_2840);
nor UO_346 (O_346,N_2650,N_2730);
or UO_347 (O_347,N_2600,N_2756);
nor UO_348 (O_348,N_2846,N_2589);
nor UO_349 (O_349,N_2632,N_2614);
or UO_350 (O_350,N_2667,N_2822);
or UO_351 (O_351,N_2946,N_2763);
nand UO_352 (O_352,N_2573,N_2992);
or UO_353 (O_353,N_2902,N_2860);
or UO_354 (O_354,N_2974,N_2769);
and UO_355 (O_355,N_2946,N_2709);
nand UO_356 (O_356,N_2618,N_2587);
nand UO_357 (O_357,N_2631,N_2674);
or UO_358 (O_358,N_2966,N_2826);
nor UO_359 (O_359,N_2694,N_2731);
and UO_360 (O_360,N_2601,N_2713);
nor UO_361 (O_361,N_2735,N_2859);
or UO_362 (O_362,N_2646,N_2628);
xor UO_363 (O_363,N_2508,N_2521);
nor UO_364 (O_364,N_2715,N_2655);
nor UO_365 (O_365,N_2550,N_2733);
or UO_366 (O_366,N_2603,N_2683);
nand UO_367 (O_367,N_2915,N_2717);
nor UO_368 (O_368,N_2803,N_2799);
and UO_369 (O_369,N_2732,N_2939);
and UO_370 (O_370,N_2933,N_2888);
nor UO_371 (O_371,N_2883,N_2613);
and UO_372 (O_372,N_2582,N_2826);
and UO_373 (O_373,N_2835,N_2704);
or UO_374 (O_374,N_2736,N_2572);
or UO_375 (O_375,N_2907,N_2515);
nor UO_376 (O_376,N_2633,N_2572);
nor UO_377 (O_377,N_2980,N_2603);
nor UO_378 (O_378,N_2558,N_2596);
xor UO_379 (O_379,N_2577,N_2904);
nor UO_380 (O_380,N_2941,N_2682);
nand UO_381 (O_381,N_2556,N_2623);
and UO_382 (O_382,N_2722,N_2838);
or UO_383 (O_383,N_2724,N_2586);
or UO_384 (O_384,N_2906,N_2503);
nand UO_385 (O_385,N_2657,N_2826);
or UO_386 (O_386,N_2559,N_2576);
nand UO_387 (O_387,N_2712,N_2749);
or UO_388 (O_388,N_2624,N_2655);
or UO_389 (O_389,N_2986,N_2596);
or UO_390 (O_390,N_2754,N_2741);
nor UO_391 (O_391,N_2929,N_2997);
nand UO_392 (O_392,N_2606,N_2526);
and UO_393 (O_393,N_2645,N_2942);
nor UO_394 (O_394,N_2903,N_2794);
and UO_395 (O_395,N_2736,N_2842);
nand UO_396 (O_396,N_2790,N_2826);
or UO_397 (O_397,N_2827,N_2515);
nand UO_398 (O_398,N_2825,N_2905);
nand UO_399 (O_399,N_2895,N_2849);
xnor UO_400 (O_400,N_2649,N_2954);
xor UO_401 (O_401,N_2883,N_2822);
xor UO_402 (O_402,N_2892,N_2756);
or UO_403 (O_403,N_2713,N_2542);
xnor UO_404 (O_404,N_2762,N_2665);
and UO_405 (O_405,N_2757,N_2748);
nand UO_406 (O_406,N_2710,N_2789);
and UO_407 (O_407,N_2626,N_2837);
nor UO_408 (O_408,N_2743,N_2757);
nand UO_409 (O_409,N_2643,N_2801);
and UO_410 (O_410,N_2586,N_2791);
nand UO_411 (O_411,N_2670,N_2893);
nor UO_412 (O_412,N_2748,N_2893);
xor UO_413 (O_413,N_2624,N_2651);
and UO_414 (O_414,N_2698,N_2579);
nand UO_415 (O_415,N_2610,N_2641);
xor UO_416 (O_416,N_2955,N_2942);
nand UO_417 (O_417,N_2696,N_2971);
xnor UO_418 (O_418,N_2773,N_2863);
nand UO_419 (O_419,N_2666,N_2716);
and UO_420 (O_420,N_2719,N_2654);
nand UO_421 (O_421,N_2622,N_2775);
xor UO_422 (O_422,N_2585,N_2991);
or UO_423 (O_423,N_2692,N_2790);
nor UO_424 (O_424,N_2802,N_2748);
nand UO_425 (O_425,N_2627,N_2527);
or UO_426 (O_426,N_2905,N_2673);
nor UO_427 (O_427,N_2921,N_2774);
or UO_428 (O_428,N_2624,N_2721);
nand UO_429 (O_429,N_2804,N_2961);
nand UO_430 (O_430,N_2564,N_2599);
nand UO_431 (O_431,N_2665,N_2742);
or UO_432 (O_432,N_2569,N_2907);
nor UO_433 (O_433,N_2951,N_2830);
and UO_434 (O_434,N_2709,N_2859);
nand UO_435 (O_435,N_2616,N_2559);
nor UO_436 (O_436,N_2701,N_2599);
or UO_437 (O_437,N_2748,N_2517);
nand UO_438 (O_438,N_2781,N_2653);
and UO_439 (O_439,N_2787,N_2554);
nand UO_440 (O_440,N_2970,N_2919);
nand UO_441 (O_441,N_2558,N_2907);
nand UO_442 (O_442,N_2643,N_2884);
nor UO_443 (O_443,N_2804,N_2724);
nor UO_444 (O_444,N_2787,N_2689);
nand UO_445 (O_445,N_2785,N_2552);
nand UO_446 (O_446,N_2836,N_2676);
nand UO_447 (O_447,N_2747,N_2715);
nand UO_448 (O_448,N_2578,N_2713);
nand UO_449 (O_449,N_2710,N_2821);
nand UO_450 (O_450,N_2722,N_2841);
xnor UO_451 (O_451,N_2972,N_2567);
or UO_452 (O_452,N_2636,N_2655);
or UO_453 (O_453,N_2941,N_2801);
xor UO_454 (O_454,N_2864,N_2501);
nor UO_455 (O_455,N_2844,N_2632);
nor UO_456 (O_456,N_2638,N_2732);
xor UO_457 (O_457,N_2775,N_2507);
or UO_458 (O_458,N_2857,N_2643);
nor UO_459 (O_459,N_2931,N_2598);
and UO_460 (O_460,N_2655,N_2919);
xor UO_461 (O_461,N_2636,N_2935);
nor UO_462 (O_462,N_2744,N_2518);
nor UO_463 (O_463,N_2961,N_2577);
nand UO_464 (O_464,N_2704,N_2681);
nand UO_465 (O_465,N_2963,N_2902);
or UO_466 (O_466,N_2783,N_2617);
or UO_467 (O_467,N_2592,N_2677);
and UO_468 (O_468,N_2926,N_2714);
or UO_469 (O_469,N_2926,N_2552);
and UO_470 (O_470,N_2962,N_2806);
nor UO_471 (O_471,N_2923,N_2685);
and UO_472 (O_472,N_2552,N_2725);
nor UO_473 (O_473,N_2976,N_2856);
nand UO_474 (O_474,N_2545,N_2695);
or UO_475 (O_475,N_2830,N_2671);
nand UO_476 (O_476,N_2807,N_2682);
or UO_477 (O_477,N_2587,N_2989);
and UO_478 (O_478,N_2752,N_2693);
nor UO_479 (O_479,N_2758,N_2597);
nand UO_480 (O_480,N_2916,N_2793);
nand UO_481 (O_481,N_2592,N_2806);
and UO_482 (O_482,N_2704,N_2793);
nand UO_483 (O_483,N_2902,N_2870);
nand UO_484 (O_484,N_2956,N_2634);
nand UO_485 (O_485,N_2513,N_2540);
and UO_486 (O_486,N_2589,N_2618);
and UO_487 (O_487,N_2705,N_2810);
nor UO_488 (O_488,N_2761,N_2535);
and UO_489 (O_489,N_2942,N_2890);
nand UO_490 (O_490,N_2597,N_2909);
nand UO_491 (O_491,N_2966,N_2523);
and UO_492 (O_492,N_2766,N_2594);
nand UO_493 (O_493,N_2574,N_2680);
nand UO_494 (O_494,N_2862,N_2999);
or UO_495 (O_495,N_2584,N_2936);
and UO_496 (O_496,N_2970,N_2917);
nor UO_497 (O_497,N_2988,N_2828);
nand UO_498 (O_498,N_2627,N_2693);
xnor UO_499 (O_499,N_2634,N_2795);
endmodule