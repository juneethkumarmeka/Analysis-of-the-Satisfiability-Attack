module basic_2500_25000_3000_10_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_1347,In_1404);
xnor U1 (N_1,In_2375,In_1594);
or U2 (N_2,In_108,In_625);
or U3 (N_3,In_1604,In_933);
and U4 (N_4,In_83,In_2241);
xor U5 (N_5,In_502,In_1501);
xor U6 (N_6,In_109,In_305);
and U7 (N_7,In_925,In_569);
nor U8 (N_8,In_830,In_41);
nor U9 (N_9,In_1798,In_200);
nor U10 (N_10,In_1768,In_726);
or U11 (N_11,In_78,In_2383);
and U12 (N_12,In_100,In_453);
or U13 (N_13,In_669,In_1640);
nor U14 (N_14,In_827,In_1828);
nor U15 (N_15,In_809,In_2160);
nor U16 (N_16,In_2078,In_2442);
or U17 (N_17,In_752,In_869);
or U18 (N_18,In_1362,In_2485);
or U19 (N_19,In_89,In_604);
or U20 (N_20,In_1164,In_1956);
nor U21 (N_21,In_978,In_1989);
or U22 (N_22,In_1176,In_1556);
xor U23 (N_23,In_340,In_997);
and U24 (N_24,In_1854,In_1023);
xor U25 (N_25,In_374,In_58);
and U26 (N_26,In_2182,In_212);
xor U27 (N_27,In_1535,In_32);
xor U28 (N_28,In_1957,In_1422);
nand U29 (N_29,In_188,In_1134);
nand U30 (N_30,In_1575,In_233);
nand U31 (N_31,In_1651,In_1006);
or U32 (N_32,In_296,In_1786);
xor U33 (N_33,In_2201,In_965);
nor U34 (N_34,In_1787,In_439);
nand U35 (N_35,In_2305,In_337);
nor U36 (N_36,In_1348,In_1197);
or U37 (N_37,In_1985,In_92);
nand U38 (N_38,In_121,In_1799);
and U39 (N_39,In_125,In_1597);
nor U40 (N_40,In_519,In_103);
and U41 (N_41,In_499,In_881);
nor U42 (N_42,In_1552,In_1170);
or U43 (N_43,In_1430,In_90);
or U44 (N_44,In_823,In_2458);
xnor U45 (N_45,In_653,In_1890);
nand U46 (N_46,In_671,In_1187);
or U47 (N_47,In_790,In_274);
nand U48 (N_48,In_369,In_1758);
nand U49 (N_49,In_2450,In_450);
and U50 (N_50,In_306,In_1479);
nand U51 (N_51,In_124,In_1897);
xor U52 (N_52,In_2341,In_2032);
xor U53 (N_53,In_316,In_406);
nor U54 (N_54,In_534,In_1408);
and U55 (N_55,In_2264,In_1109);
or U56 (N_56,In_1064,In_39);
nand U57 (N_57,In_1901,In_596);
nand U58 (N_58,In_244,In_1959);
nand U59 (N_59,In_853,In_434);
or U60 (N_60,In_2126,In_2074);
xnor U61 (N_61,In_2193,In_907);
or U62 (N_62,In_2287,In_1855);
or U63 (N_63,In_936,In_2400);
and U64 (N_64,In_1783,In_2115);
nand U65 (N_65,In_1279,In_1942);
xor U66 (N_66,In_1240,In_1053);
nand U67 (N_67,In_1540,In_1384);
xor U68 (N_68,In_578,In_2213);
nor U69 (N_69,In_350,In_486);
xnor U70 (N_70,In_2202,In_2374);
nor U71 (N_71,In_2357,In_1421);
xnor U72 (N_72,In_1548,In_1813);
and U73 (N_73,In_74,In_440);
xor U74 (N_74,In_1782,In_2415);
nand U75 (N_75,In_242,In_201);
nor U76 (N_76,In_651,In_36);
xor U77 (N_77,In_530,In_2154);
nor U78 (N_78,In_1034,In_1600);
nand U79 (N_79,In_163,In_2354);
xor U80 (N_80,In_1152,In_2421);
nand U81 (N_81,In_1285,In_375);
nand U82 (N_82,In_216,In_182);
xor U83 (N_83,In_798,In_1199);
nand U84 (N_84,In_318,In_1486);
nor U85 (N_85,In_2216,In_57);
or U86 (N_86,In_1297,In_118);
and U87 (N_87,In_821,In_463);
nand U88 (N_88,In_2144,In_65);
nor U89 (N_89,In_2382,In_2416);
or U90 (N_90,In_1533,In_695);
or U91 (N_91,In_1143,In_1774);
nand U92 (N_92,In_2292,In_2176);
nor U93 (N_93,In_1793,In_1983);
xor U94 (N_94,In_693,In_1724);
nand U95 (N_95,In_642,In_2285);
xnor U96 (N_96,In_687,In_102);
nand U97 (N_97,In_592,In_268);
nand U98 (N_98,In_970,In_27);
and U99 (N_99,In_1233,In_1725);
nor U100 (N_100,In_394,In_1731);
xor U101 (N_101,In_1261,In_824);
nand U102 (N_102,In_1491,In_1296);
or U103 (N_103,In_1081,In_929);
and U104 (N_104,In_744,In_1282);
nor U105 (N_105,In_527,In_2000);
nor U106 (N_106,In_1085,In_2271);
or U107 (N_107,In_21,In_1214);
nand U108 (N_108,In_1365,In_2380);
nand U109 (N_109,In_1092,In_1973);
and U110 (N_110,In_889,In_928);
nand U111 (N_111,In_932,In_944);
or U112 (N_112,In_2215,In_553);
or U113 (N_113,In_470,In_52);
and U114 (N_114,In_1172,In_1975);
or U115 (N_115,In_97,In_2304);
nor U116 (N_116,In_1242,In_227);
and U117 (N_117,In_1280,In_1780);
xnor U118 (N_118,In_1505,In_1858);
xor U119 (N_119,In_2166,In_1177);
and U120 (N_120,In_1675,In_1709);
nor U121 (N_121,In_682,In_2082);
nor U122 (N_122,In_1537,In_2147);
and U123 (N_123,In_166,In_1883);
nand U124 (N_124,In_615,In_1070);
nor U125 (N_125,In_1732,In_577);
xor U126 (N_126,In_1551,In_115);
nor U127 (N_127,In_2235,In_1496);
or U128 (N_128,In_2398,In_1200);
nand U129 (N_129,In_430,In_819);
or U130 (N_130,In_205,In_1423);
nand U131 (N_131,In_1390,In_1991);
and U132 (N_132,In_1754,In_1342);
nor U133 (N_133,In_731,In_1254);
xor U134 (N_134,In_354,In_2171);
and U135 (N_135,In_660,In_483);
or U136 (N_136,In_568,In_2262);
and U137 (N_137,In_2351,In_775);
xnor U138 (N_138,In_1628,In_1645);
xnor U139 (N_139,In_105,In_491);
or U140 (N_140,In_2013,In_1232);
xnor U141 (N_141,In_1665,In_1656);
and U142 (N_142,In_1457,In_1616);
nand U143 (N_143,In_1008,In_1874);
or U144 (N_144,In_663,In_1104);
nor U145 (N_145,In_1952,In_1664);
and U146 (N_146,In_648,In_1933);
and U147 (N_147,In_2464,In_938);
or U148 (N_148,In_1898,In_1610);
and U149 (N_149,In_1845,In_1573);
or U150 (N_150,In_88,In_996);
nand U151 (N_151,In_2425,In_1425);
nor U152 (N_152,In_395,In_1075);
and U153 (N_153,In_1831,In_1899);
nor U154 (N_154,In_681,In_1389);
or U155 (N_155,In_110,In_1930);
nor U156 (N_156,In_1945,In_1943);
nand U157 (N_157,In_2343,In_2427);
and U158 (N_158,In_1520,In_2462);
and U159 (N_159,In_1887,In_956);
nand U160 (N_160,In_1843,In_104);
and U161 (N_161,In_1792,In_355);
nand U162 (N_162,In_349,In_570);
xnor U163 (N_163,In_315,In_753);
and U164 (N_164,In_2151,In_1797);
nor U165 (N_165,In_2217,In_1944);
nand U166 (N_166,In_1990,In_66);
or U167 (N_167,In_1161,In_1621);
or U168 (N_168,In_1340,In_23);
or U169 (N_169,In_372,In_1133);
xnor U170 (N_170,In_977,In_714);
xor U171 (N_171,In_1067,In_2163);
nor U172 (N_172,In_150,In_1574);
or U173 (N_173,In_609,In_2052);
nand U174 (N_174,In_1293,In_1881);
xor U175 (N_175,In_649,In_703);
nor U176 (N_176,In_1117,In_407);
xnor U177 (N_177,In_503,In_2258);
nand U178 (N_178,In_1205,In_202);
xnor U179 (N_179,In_1166,In_2021);
nand U180 (N_180,In_2220,In_1720);
or U181 (N_181,In_2306,In_1585);
nand U182 (N_182,In_582,In_1609);
nor U183 (N_183,In_516,In_1019);
xor U184 (N_184,In_1746,In_449);
xor U185 (N_185,In_804,In_178);
xor U186 (N_186,In_2286,In_1914);
nor U187 (N_187,In_898,In_2325);
xnor U188 (N_188,In_284,In_1321);
or U189 (N_189,In_878,In_2066);
and U190 (N_190,In_2247,In_1788);
xor U191 (N_191,In_1542,In_185);
nor U192 (N_192,In_704,In_221);
or U193 (N_193,In_1059,In_618);
or U194 (N_194,In_451,In_1712);
nor U195 (N_195,In_1511,In_1372);
and U196 (N_196,In_2125,In_1777);
and U197 (N_197,In_1114,In_1459);
or U198 (N_198,In_2278,In_1905);
nor U199 (N_199,In_1449,In_967);
xor U200 (N_200,In_1153,In_230);
nand U201 (N_201,In_1028,In_141);
nand U202 (N_202,In_994,In_1156);
nor U203 (N_203,In_2475,In_2498);
and U204 (N_204,In_931,In_1719);
nor U205 (N_205,In_2404,In_2109);
and U206 (N_206,In_1424,In_538);
and U207 (N_207,In_854,In_1212);
nand U208 (N_208,In_1703,In_748);
and U209 (N_209,In_1359,In_299);
nand U210 (N_210,In_2050,In_1235);
or U211 (N_211,In_129,In_1194);
nor U212 (N_212,In_358,In_2091);
xnor U213 (N_213,In_2092,In_1663);
xnor U214 (N_214,In_1693,In_248);
and U215 (N_215,In_1925,In_0);
or U216 (N_216,In_1373,In_431);
or U217 (N_217,In_2494,In_1912);
and U218 (N_218,In_771,In_972);
nor U219 (N_219,In_1658,In_1747);
or U220 (N_220,In_399,In_24);
nand U221 (N_221,In_894,In_688);
xor U222 (N_222,In_1270,In_1497);
or U223 (N_223,In_1592,In_370);
xor U224 (N_224,In_532,In_1318);
nor U225 (N_225,In_1572,In_734);
nand U226 (N_226,In_1795,In_2087);
and U227 (N_227,In_1829,In_958);
nor U228 (N_228,In_1687,In_1637);
or U229 (N_229,In_137,In_1298);
nor U230 (N_230,In_760,In_2489);
nor U231 (N_231,In_2138,In_1826);
or U232 (N_232,In_884,In_2282);
nor U233 (N_233,In_352,In_139);
or U234 (N_234,In_1821,In_1705);
or U235 (N_235,In_1888,In_509);
xor U236 (N_236,In_1623,In_162);
or U237 (N_237,In_1713,In_2332);
nor U238 (N_238,In_1437,In_54);
and U239 (N_239,In_620,In_2101);
and U240 (N_240,In_2227,In_981);
xor U241 (N_241,In_91,In_2452);
or U242 (N_242,In_1872,In_728);
nand U243 (N_243,In_194,In_2408);
xnor U244 (N_244,In_1869,In_1208);
xnor U245 (N_245,In_2157,In_1679);
nand U246 (N_246,In_2010,In_2081);
nor U247 (N_247,In_947,In_1541);
xnor U248 (N_248,In_1891,In_1434);
or U249 (N_249,In_2496,In_2131);
or U250 (N_250,In_1695,In_2379);
and U251 (N_251,In_2367,In_559);
or U252 (N_252,In_258,In_1072);
and U253 (N_253,In_347,In_1095);
xnor U254 (N_254,In_1876,In_14);
xnor U255 (N_255,In_1369,In_2146);
xnor U256 (N_256,In_336,In_1169);
nand U257 (N_257,In_303,In_542);
nor U258 (N_258,In_1866,In_1056);
and U259 (N_259,In_1251,In_1776);
xnor U260 (N_260,In_2495,In_813);
and U261 (N_261,In_617,In_300);
and U262 (N_262,In_801,In_2175);
nand U263 (N_263,In_198,In_1910);
or U264 (N_264,In_1441,In_2386);
nand U265 (N_265,In_1847,In_1032);
or U266 (N_266,In_280,In_1877);
nand U267 (N_267,In_712,In_1288);
and U268 (N_268,In_581,In_1697);
or U269 (N_269,In_839,In_1627);
or U270 (N_270,In_832,In_1311);
and U271 (N_271,In_101,In_2256);
and U272 (N_272,In_2338,In_1010);
or U273 (N_273,In_677,In_1108);
xor U274 (N_274,In_338,In_1393);
nand U275 (N_275,In_1805,In_893);
and U276 (N_276,In_2242,In_2309);
xnor U277 (N_277,In_2037,In_1071);
xor U278 (N_278,In_1779,In_1678);
or U279 (N_279,In_1473,In_2469);
nand U280 (N_280,In_75,In_1988);
or U281 (N_281,In_595,In_1461);
or U282 (N_282,In_951,In_701);
and U283 (N_283,In_1643,In_1642);
xor U284 (N_284,In_1265,In_1455);
and U285 (N_285,In_2244,In_1688);
nand U286 (N_286,In_1699,In_1377);
xnor U287 (N_287,In_1175,In_2);
nand U288 (N_288,In_1916,In_2329);
nand U289 (N_289,In_1512,In_2478);
xor U290 (N_290,In_1385,In_1031);
nand U291 (N_291,In_1918,In_796);
or U292 (N_292,In_2466,In_301);
xnor U293 (N_293,In_259,In_690);
and U294 (N_294,In_179,In_1036);
nand U295 (N_295,In_95,In_1309);
and U296 (N_296,In_1583,In_62);
nand U297 (N_297,In_1727,In_1033);
and U298 (N_298,In_2359,In_1051);
and U299 (N_299,In_2186,In_1859);
nor U300 (N_300,In_339,In_497);
nor U301 (N_301,In_1633,In_1403);
and U302 (N_302,In_650,In_2099);
nand U303 (N_303,In_1084,In_547);
or U304 (N_304,In_706,In_2482);
nor U305 (N_305,In_50,In_2226);
nand U306 (N_306,In_1150,In_1121);
nand U307 (N_307,In_1135,In_586);
nand U308 (N_308,In_2336,In_468);
or U309 (N_309,In_1650,In_1841);
or U310 (N_310,In_366,In_915);
nand U311 (N_311,In_1922,In_2326);
nor U312 (N_312,In_633,In_694);
or U313 (N_313,In_2321,In_1894);
xnor U314 (N_314,In_319,In_1333);
xnor U315 (N_315,In_1846,In_1951);
nand U316 (N_316,In_1063,In_2270);
nor U317 (N_317,In_2016,In_1380);
xnor U318 (N_318,In_1801,In_195);
nand U319 (N_319,In_246,In_1387);
nor U320 (N_320,In_1076,In_1613);
nor U321 (N_321,In_1800,In_2279);
and U322 (N_322,In_999,In_419);
or U323 (N_323,In_1029,In_900);
and U324 (N_324,In_602,In_1742);
or U325 (N_325,In_1954,In_666);
nor U326 (N_326,In_1772,In_2397);
and U327 (N_327,In_721,In_2158);
or U328 (N_328,In_2294,In_2224);
and U329 (N_329,In_335,In_788);
nand U330 (N_330,In_1743,In_456);
or U331 (N_331,In_1304,In_329);
or U332 (N_332,In_870,In_1044);
nand U333 (N_333,In_1183,In_1508);
nand U334 (N_334,In_949,In_1096);
nor U335 (N_335,In_2024,In_659);
nor U336 (N_336,In_657,In_1873);
and U337 (N_337,In_2257,In_1765);
and U338 (N_338,In_2200,In_494);
nor U339 (N_339,In_1677,In_2316);
xor U340 (N_340,In_1494,In_1807);
or U341 (N_341,In_833,In_1701);
or U342 (N_342,In_1868,In_1862);
xnor U343 (N_343,In_224,In_1723);
and U344 (N_344,In_40,In_2246);
and U345 (N_345,In_782,In_2467);
or U346 (N_346,In_1447,In_362);
and U347 (N_347,In_2164,In_2263);
nor U348 (N_348,In_2148,In_909);
nor U349 (N_349,In_1415,In_2364);
and U350 (N_350,In_1935,In_1219);
nor U351 (N_351,In_1790,In_1968);
xor U352 (N_352,In_562,In_756);
nor U353 (N_353,In_1538,In_382);
nor U354 (N_354,In_1560,In_482);
nor U355 (N_355,In_1475,In_2484);
or U356 (N_356,In_1722,In_1634);
or U357 (N_357,In_639,In_2327);
xor U358 (N_358,In_1079,In_147);
xor U359 (N_359,In_2056,In_1181);
or U360 (N_360,In_1301,In_1802);
xnor U361 (N_361,In_2155,In_1875);
and U362 (N_362,In_2077,In_1291);
nor U363 (N_363,In_1198,In_2323);
and U364 (N_364,In_781,In_1635);
xor U365 (N_365,In_10,In_1371);
or U366 (N_366,In_1413,In_1700);
nand U367 (N_367,In_1256,In_1303);
nand U368 (N_368,In_2405,In_767);
or U369 (N_369,In_1769,In_55);
or U370 (N_370,In_556,In_1547);
xor U371 (N_371,In_1416,In_1559);
nand U372 (N_372,In_6,In_848);
and U373 (N_373,In_2080,In_1379);
and U374 (N_374,In_2371,In_656);
nand U375 (N_375,In_184,In_1391);
xnor U376 (N_376,In_1454,In_313);
and U377 (N_377,In_1683,In_203);
nor U378 (N_378,In_2266,In_528);
and U379 (N_379,In_1611,In_1982);
nand U380 (N_380,In_2123,In_1680);
nor U381 (N_381,In_1804,In_1814);
nand U382 (N_382,In_1694,In_2443);
nor U383 (N_383,In_2044,In_1524);
nor U384 (N_384,In_93,In_2018);
or U385 (N_385,In_2236,In_2454);
xnor U386 (N_386,In_1436,In_808);
and U387 (N_387,In_2180,In_1484);
or U388 (N_388,In_598,In_2033);
nand U389 (N_389,In_588,In_739);
nand U390 (N_390,In_806,In_1525);
nand U391 (N_391,In_749,In_1381);
xor U392 (N_392,In_2250,In_902);
xor U393 (N_393,In_85,In_1676);
and U394 (N_394,In_2295,In_696);
or U395 (N_395,In_1103,In_855);
nor U396 (N_396,In_2406,In_1653);
xor U397 (N_397,In_1262,In_1244);
nor U398 (N_398,In_2275,In_1123);
or U399 (N_399,In_2134,In_852);
nor U400 (N_400,In_365,In_1963);
and U401 (N_401,In_1686,In_860);
nor U402 (N_402,In_2497,In_1691);
xor U403 (N_403,In_738,In_444);
nor U404 (N_404,In_2108,In_514);
and U405 (N_405,In_628,In_550);
and U406 (N_406,In_1002,In_2248);
nor U407 (N_407,In_1612,In_1048);
and U408 (N_408,In_292,In_241);
nand U409 (N_409,In_842,In_2387);
nand U410 (N_410,In_183,In_1221);
and U411 (N_411,In_1442,In_1994);
and U412 (N_412,In_1532,In_67);
nand U413 (N_413,In_1138,In_1791);
xnor U414 (N_414,In_1188,In_716);
xor U415 (N_415,In_297,In_177);
or U416 (N_416,In_2280,In_2413);
nand U417 (N_417,In_134,In_408);
xnor U418 (N_418,In_2204,In_799);
or U419 (N_419,In_2401,In_1091);
and U420 (N_420,In_526,In_580);
or U421 (N_421,In_17,In_2090);
and U422 (N_422,In_939,In_43);
xnor U423 (N_423,In_1458,In_2187);
and U424 (N_424,In_1339,In_2065);
and U425 (N_425,In_1139,In_652);
xor U426 (N_426,In_1407,In_2490);
nor U427 (N_427,In_1386,In_2276);
or U428 (N_428,In_142,In_2221);
nor U429 (N_429,In_524,In_86);
nand U430 (N_430,In_1346,In_942);
nand U431 (N_431,In_746,In_426);
xnor U432 (N_432,In_1657,In_1062);
or U433 (N_433,In_1599,In_333);
or U434 (N_434,In_636,In_950);
nand U435 (N_435,In_1764,In_225);
xor U436 (N_436,In_448,In_488);
nand U437 (N_437,In_961,In_792);
xor U438 (N_438,In_1191,In_1632);
nor U439 (N_439,In_1974,In_1025);
nand U440 (N_440,In_2062,In_2222);
nand U441 (N_441,In_1892,In_22);
nor U442 (N_442,In_1966,In_2086);
and U443 (N_443,In_1137,In_831);
and U444 (N_444,In_1741,In_1570);
nor U445 (N_445,In_1196,In_1815);
nor U446 (N_446,In_1825,In_1671);
xnor U447 (N_447,In_1088,In_72);
nand U448 (N_448,In_1539,In_1509);
nor U449 (N_449,In_243,In_637);
or U450 (N_450,In_1328,In_1223);
and U451 (N_451,In_1522,In_857);
nor U452 (N_452,In_149,In_2237);
or U453 (N_453,In_579,In_346);
and U454 (N_454,In_1766,In_247);
or U455 (N_455,In_1770,In_392);
xnor U456 (N_456,In_2345,In_1714);
nand U457 (N_457,In_2433,In_1148);
or U458 (N_458,In_1165,In_152);
and U459 (N_459,In_232,In_635);
and U460 (N_460,In_111,In_1978);
xnor U461 (N_461,In_1065,In_267);
or U462 (N_462,In_1850,In_1852);
or U463 (N_463,In_1314,In_835);
nor U464 (N_464,In_1101,In_447);
and U465 (N_465,In_1106,In_1257);
and U466 (N_466,In_2001,In_851);
and U467 (N_467,In_1299,In_1119);
xor U468 (N_468,In_561,In_2145);
or U469 (N_469,In_1950,In_228);
nand U470 (N_470,In_2407,In_892);
and U471 (N_471,In_1322,In_603);
or U472 (N_472,In_7,In_1294);
nor U473 (N_473,In_989,In_1842);
nor U474 (N_474,In_2277,In_606);
and U475 (N_475,In_460,In_1647);
nor U476 (N_476,In_436,In_828);
or U477 (N_477,In_2274,In_2479);
and U478 (N_478,In_1083,In_1816);
and U479 (N_479,In_192,In_1050);
or U480 (N_480,In_1068,In_822);
nor U481 (N_481,In_2435,In_1498);
xor U482 (N_482,In_12,In_698);
xor U483 (N_483,In_343,In_724);
nand U484 (N_484,In_308,In_2487);
or U485 (N_485,In_1468,In_2419);
nand U486 (N_486,In_116,In_1024);
nor U487 (N_487,In_1606,In_1027);
and U488 (N_488,In_2348,In_2085);
nand U489 (N_489,In_238,In_512);
nand U490 (N_490,In_1907,In_1157);
and U491 (N_491,In_2268,In_275);
nor U492 (N_492,In_2228,In_1042);
and U493 (N_493,In_2358,In_480);
and U494 (N_494,In_2113,In_1364);
and U495 (N_495,In_2194,In_1094);
and U496 (N_496,In_1343,In_2448);
and U497 (N_497,In_2079,In_2255);
xnor U498 (N_498,In_1324,In_2284);
or U499 (N_499,In_1222,In_479);
nor U500 (N_500,In_1480,In_750);
and U501 (N_501,In_218,In_1241);
nand U502 (N_502,In_1544,In_263);
and U503 (N_503,In_1803,In_1558);
nor U504 (N_504,In_2112,In_945);
nand U505 (N_505,In_1217,In_729);
nand U506 (N_506,In_1211,In_1267);
nor U507 (N_507,In_960,In_647);
and U508 (N_508,In_106,In_454);
or U509 (N_509,In_1553,In_1624);
nor U510 (N_510,In_511,In_1168);
nor U511 (N_511,In_986,In_619);
and U512 (N_512,In_993,In_257);
and U513 (N_513,In_2124,In_1105);
xor U514 (N_514,In_172,In_1590);
nor U515 (N_515,In_1243,In_1971);
xnor U516 (N_516,In_1506,In_2005);
and U517 (N_517,In_764,In_190);
nand U518 (N_518,In_373,In_779);
nor U519 (N_519,In_231,In_2003);
and U520 (N_520,In_291,In_260);
nand U521 (N_521,In_461,In_135);
or U522 (N_522,In_638,In_1127);
and U523 (N_523,In_2027,In_334);
nand U524 (N_524,In_458,In_973);
nand U525 (N_525,In_1644,In_35);
nand U526 (N_526,In_2026,In_117);
nand U527 (N_527,In_1470,In_1038);
or U528 (N_528,In_1419,In_1648);
xnor U529 (N_529,In_525,In_722);
and U530 (N_530,In_975,In_1773);
xor U531 (N_531,In_25,In_1682);
and U532 (N_532,In_2206,In_1007);
and U533 (N_533,In_2430,In_1252);
or U534 (N_534,In_1,In_11);
nand U535 (N_535,In_1099,In_1717);
xor U536 (N_536,In_1477,In_843);
and U537 (N_537,In_1625,In_1431);
and U538 (N_538,In_1856,In_1399);
nor U539 (N_539,In_1588,In_181);
or U540 (N_540,In_1760,In_1274);
xnor U541 (N_541,In_1596,In_1041);
nand U542 (N_542,In_1827,In_45);
and U543 (N_543,In_174,In_4);
and U544 (N_544,In_918,In_381);
nand U545 (N_545,In_2423,In_1401);
or U546 (N_546,In_2392,In_1184);
nor U547 (N_547,In_1319,In_279);
and U548 (N_548,In_2483,In_351);
xnor U549 (N_549,In_2355,In_727);
or U550 (N_550,In_811,In_531);
xor U551 (N_551,In_1272,In_1502);
nor U552 (N_552,In_1981,In_107);
or U553 (N_553,In_2061,In_160);
or U554 (N_554,In_2243,In_1681);
xor U555 (N_555,In_2411,In_13);
nand U556 (N_556,In_151,In_368);
xnor U557 (N_557,In_1576,In_1684);
xor U558 (N_558,In_1504,In_2071);
and U559 (N_559,In_2051,In_2028);
and U560 (N_560,In_1237,In_927);
xnor U561 (N_561,In_2162,In_1018);
and U562 (N_562,In_1026,In_1830);
nand U563 (N_563,In_289,In_2456);
nor U564 (N_564,In_146,In_1100);
and U565 (N_565,In_1543,In_590);
xor U566 (N_566,In_1924,In_208);
or U567 (N_567,In_256,In_376);
nand U568 (N_568,In_325,In_1629);
nor U569 (N_569,In_2168,In_1331);
or U570 (N_570,In_2122,In_1667);
and U571 (N_571,In_1039,In_1086);
nor U572 (N_572,In_53,In_2313);
xor U573 (N_573,In_1463,In_1011);
and U574 (N_574,In_560,In_2480);
xnor U575 (N_575,In_2319,In_1716);
nor U576 (N_576,In_196,In_988);
nand U577 (N_577,In_388,In_1639);
nor U578 (N_578,In_1492,In_1771);
xnor U579 (N_579,In_1402,In_611);
or U580 (N_580,In_1054,In_2389);
xor U581 (N_581,In_1921,In_626);
and U582 (N_582,In_130,In_797);
or U583 (N_583,In_393,In_2067);
xnor U584 (N_584,In_661,In_176);
nor U585 (N_585,In_1306,In_2007);
xnor U586 (N_586,In_423,In_1626);
and U587 (N_587,In_475,In_717);
and U588 (N_588,In_543,In_2042);
xor U589 (N_589,In_1735,In_410);
and U590 (N_590,In_2172,In_751);
nor U591 (N_591,In_1213,In_654);
or U592 (N_592,In_2057,In_1248);
nor U593 (N_593,In_1323,In_2429);
or U594 (N_594,In_1140,In_1107);
or U595 (N_595,In_1937,In_1349);
nor U596 (N_596,In_2011,In_1601);
and U597 (N_597,In_1443,In_391);
and U598 (N_598,In_1488,In_1173);
xor U599 (N_599,In_421,In_1972);
nand U600 (N_600,In_1266,In_398);
nor U601 (N_601,In_2130,In_816);
nand U602 (N_602,In_1514,In_1015);
nand U603 (N_603,In_1698,In_2141);
and U604 (N_604,In_546,In_63);
xor U605 (N_605,In_845,In_616);
and U606 (N_606,In_873,In_1513);
and U607 (N_607,In_2149,In_847);
xor U608 (N_608,In_2029,In_2302);
nand U609 (N_609,In_1396,In_457);
or U610 (N_610,In_1097,In_2232);
xor U611 (N_611,In_963,In_883);
or U612 (N_612,In_2403,In_995);
nor U613 (N_613,In_169,In_1395);
or U614 (N_614,In_536,In_171);
nand U615 (N_615,In_442,In_1432);
nand U616 (N_616,In_262,In_1778);
nor U617 (N_617,In_1762,In_1970);
nor U618 (N_618,In_219,In_2234);
nor U619 (N_619,In_2210,In_1130);
and U620 (N_620,In_1569,In_1810);
or U621 (N_621,In_1865,In_281);
nand U622 (N_622,In_1185,In_210);
or U623 (N_623,In_557,In_1263);
nand U624 (N_624,In_572,In_220);
nand U625 (N_625,In_515,In_720);
and U626 (N_626,In_136,In_1929);
and U627 (N_627,In_785,In_1987);
nand U628 (N_628,In_323,In_42);
or U629 (N_629,In_762,In_462);
nand U630 (N_630,In_758,In_2088);
or U631 (N_631,In_1451,In_678);
nor U632 (N_632,In_412,In_2377);
or U633 (N_633,In_1174,In_2009);
or U634 (N_634,In_371,In_2073);
and U635 (N_635,In_411,In_2197);
nor U636 (N_636,In_1450,In_937);
nor U637 (N_637,In_1578,In_1182);
xnor U638 (N_638,In_401,In_1158);
or U639 (N_639,In_156,In_1336);
nor U640 (N_640,In_1965,In_1231);
xnor U641 (N_641,In_1334,In_2097);
nand U642 (N_642,In_679,In_1878);
or U643 (N_643,In_2455,In_138);
or U644 (N_644,In_954,In_2366);
xnor U645 (N_645,In_867,In_1493);
or U646 (N_646,In_396,In_856);
or U647 (N_647,In_912,In_2190);
or U648 (N_648,In_2301,In_1004);
nor U649 (N_649,In_1510,In_1889);
and U650 (N_650,In_1264,In_1500);
xor U651 (N_651,In_2198,In_1745);
nor U652 (N_652,In_282,In_167);
nor U653 (N_653,In_2184,In_2014);
nand U654 (N_654,In_2470,In_715);
or U655 (N_655,In_33,In_207);
xor U656 (N_656,In_1089,In_953);
xnor U657 (N_657,In_272,In_627);
or U658 (N_658,In_276,In_1895);
nor U659 (N_659,In_1195,In_1579);
nor U660 (N_660,In_1489,In_1737);
and U661 (N_661,In_472,In_1886);
nand U662 (N_662,In_699,In_683);
xor U663 (N_663,In_2396,In_26);
xnor U664 (N_664,In_1310,In_484);
and U665 (N_665,In_1726,In_413);
nand U666 (N_666,In_326,In_161);
nand U667 (N_667,In_473,In_77);
nand U668 (N_668,In_2239,In_94);
nand U669 (N_669,In_1113,In_261);
or U670 (N_670,In_1563,In_404);
nand U671 (N_671,In_68,In_921);
or U672 (N_672,In_667,In_18);
or U673 (N_673,In_741,In_1239);
and U674 (N_674,In_1366,In_2240);
or U675 (N_675,In_2472,In_2251);
xnor U676 (N_676,In_1917,In_1409);
and U677 (N_677,In_96,In_1374);
or U678 (N_678,In_676,In_2493);
nor U679 (N_679,In_1131,In_1582);
xnor U680 (N_680,In_1102,In_1186);
xor U681 (N_681,In_48,In_474);
nor U682 (N_682,In_1545,In_1308);
nand U683 (N_683,In_2230,In_197);
or U684 (N_684,In_2173,In_791);
nand U685 (N_685,In_2388,In_612);
nor U686 (N_686,In_903,In_1357);
xnor U687 (N_687,In_1405,In_1268);
nand U688 (N_688,In_1819,In_1673);
and U689 (N_689,In_2344,In_608);
or U690 (N_690,In_307,In_2426);
or U691 (N_691,In_1129,In_2114);
and U692 (N_692,In_971,In_360);
or U693 (N_693,In_1690,In_1439);
xnor U694 (N_694,In_302,In_1203);
and U695 (N_695,In_345,In_1058);
nand U696 (N_696,In_266,In_1111);
nor U697 (N_697,In_1427,In_761);
xor U698 (N_698,In_1962,In_2418);
or U699 (N_699,In_363,In_904);
or U700 (N_700,In_1467,In_644);
nor U701 (N_701,In_1561,In_1849);
nor U702 (N_702,In_1851,In_464);
nand U703 (N_703,In_1110,In_2291);
nor U704 (N_704,In_1740,In_1474);
nor U705 (N_705,In_1281,In_1465);
nand U706 (N_706,In_2225,In_2308);
or U707 (N_707,In_1341,In_1418);
or U708 (N_708,In_2219,In_1589);
nand U709 (N_709,In_778,In_2360);
or U710 (N_710,In_2399,In_1128);
nor U711 (N_711,In_145,In_2471);
nor U712 (N_712,In_1020,In_1204);
xor U713 (N_713,In_29,In_1756);
and U714 (N_714,In_15,In_1955);
xor U715 (N_715,In_613,In_1618);
and U716 (N_716,In_1750,In_1307);
or U717 (N_717,In_784,In_1967);
or U718 (N_718,In_157,In_1523);
nand U719 (N_719,In_836,In_2102);
or U720 (N_720,In_1941,In_1515);
nand U721 (N_721,In_277,In_1225);
nand U722 (N_722,In_424,In_378);
and U723 (N_723,In_159,In_476);
xnor U724 (N_724,In_1730,In_1706);
nor U725 (N_725,In_1550,In_2153);
nor U726 (N_726,In_641,In_1258);
and U727 (N_727,In_686,In_342);
and U728 (N_728,In_87,In_70);
nand U729 (N_729,In_2183,In_1580);
or U730 (N_730,In_1022,In_923);
and U731 (N_731,In_1710,In_2317);
nor U732 (N_732,In_1557,In_2303);
nor U733 (N_733,In_523,In_948);
nand U734 (N_734,In_1755,In_700);
or U735 (N_735,In_552,In_8);
nand U736 (N_736,In_1159,In_2322);
nand U737 (N_737,In_1832,In_213);
xnor U738 (N_738,In_501,In_312);
nor U739 (N_739,In_2296,In_1662);
nand U740 (N_740,In_2440,In_1167);
xor U741 (N_741,In_2349,In_64);
nand U742 (N_742,In_1350,In_776);
and U743 (N_743,In_445,In_1964);
or U744 (N_744,In_1259,In_1605);
and U745 (N_745,In_1247,In_84);
xnor U746 (N_746,In_1316,In_1001);
nor U747 (N_747,In_2055,In_2468);
nand U748 (N_748,In_1253,In_1885);
nor U749 (N_749,In_390,In_1809);
xor U750 (N_750,In_1834,In_1394);
or U751 (N_751,In_1315,In_132);
and U752 (N_752,In_2297,In_2188);
and U753 (N_753,In_322,In_2476);
or U754 (N_754,In_2459,In_1711);
nor U755 (N_755,In_888,In_1005);
and U756 (N_756,In_2330,In_1636);
xor U757 (N_757,In_2075,In_1591);
and U758 (N_758,In_2342,In_874);
nor U759 (N_759,In_1344,In_1228);
or U760 (N_760,In_1670,In_1283);
nor U761 (N_761,In_402,In_1953);
and U762 (N_762,In_1230,In_1685);
or U763 (N_763,In_576,In_2252);
and U764 (N_764,In_493,In_466);
nand U765 (N_765,In_3,In_2096);
xnor U766 (N_766,In_9,In_2409);
nor U767 (N_767,In_838,In_288);
nand U768 (N_768,In_206,In_2127);
xnor U769 (N_769,In_2120,In_452);
nand U770 (N_770,In_887,In_814);
or U771 (N_771,In_1757,In_807);
nor U772 (N_772,In_545,In_2324);
xor U773 (N_773,In_2002,In_222);
nand U774 (N_774,In_1920,In_1271);
and U775 (N_775,In_1749,In_2352);
xnor U776 (N_776,In_1375,In_632);
or U777 (N_777,In_624,In_513);
nor U778 (N_778,In_1516,In_537);
nand U779 (N_779,In_1948,In_1353);
and U780 (N_780,In_2315,In_2362);
or U781 (N_781,In_2298,In_389);
xor U782 (N_782,In_1718,In_769);
xor U783 (N_783,In_359,In_2474);
xnor U784 (N_784,In_2025,In_2107);
and U785 (N_785,In_38,In_199);
and U786 (N_786,In_2207,In_1527);
nor U787 (N_787,In_812,In_2424);
or U788 (N_788,In_446,In_1564);
xnor U789 (N_789,In_314,In_2140);
or U790 (N_790,In_783,In_1429);
and U791 (N_791,In_1702,In_1207);
xnor U792 (N_792,In_1145,In_674);
and U793 (N_793,In_2105,In_1098);
nor U794 (N_794,In_2072,In_492);
xor U795 (N_795,In_574,In_2300);
and U796 (N_796,In_1035,In_630);
nor U797 (N_797,In_332,In_2034);
and U798 (N_798,In_120,In_1060);
nand U799 (N_799,In_891,In_563);
xnor U800 (N_800,In_490,In_1481);
nor U801 (N_801,In_672,In_1057);
nand U802 (N_802,In_481,In_730);
or U803 (N_803,In_1047,In_1595);
nand U804 (N_804,In_911,In_1565);
nand U805 (N_805,In_2178,In_984);
and U806 (N_806,In_723,In_357);
nand U807 (N_807,In_133,In_1880);
nand U808 (N_808,In_685,In_708);
xor U809 (N_809,In_1936,In_429);
or U810 (N_810,In_2192,In_2205);
or U811 (N_811,In_2038,In_414);
and U812 (N_812,In_30,In_2363);
nand U813 (N_813,In_1598,In_1162);
and U814 (N_814,In_665,In_787);
or U815 (N_815,In_1126,In_2293);
xor U816 (N_816,In_800,In_144);
xnor U817 (N_817,In_1784,In_1462);
or U818 (N_818,In_1646,In_879);
and U819 (N_819,In_876,In_713);
nand U820 (N_820,In_2414,In_1517);
xor U821 (N_821,In_1848,In_2039);
xor U822 (N_822,In_2208,In_982);
nand U823 (N_823,In_1668,In_614);
and U824 (N_824,In_1620,In_998);
or U825 (N_825,In_1836,In_2095);
or U826 (N_826,In_1216,In_2150);
and U827 (N_827,In_1812,In_239);
xor U828 (N_828,In_170,In_2040);
or U829 (N_829,In_148,In_691);
or U830 (N_830,In_962,In_465);
nand U831 (N_831,In_793,In_204);
nand U832 (N_832,In_1345,In_126);
or U833 (N_833,In_1833,In_1482);
nand U834 (N_834,In_564,In_1999);
nand U835 (N_835,In_2103,In_2434);
xnor U836 (N_836,In_1017,In_428);
and U837 (N_837,In_2373,In_1947);
nand U838 (N_838,In_2436,In_1124);
and U839 (N_839,In_535,In_571);
or U840 (N_840,In_1857,In_49);
xnor U841 (N_841,In_926,In_2391);
xor U842 (N_842,In_920,In_418);
nand U843 (N_843,In_2310,In_872);
and U844 (N_844,In_215,In_2179);
or U845 (N_845,In_786,In_2070);
or U846 (N_846,In_1567,In_2093);
or U847 (N_847,In_1355,In_420);
nor U848 (N_848,In_969,In_645);
and U849 (N_849,In_1638,In_974);
nand U850 (N_850,In_1986,In_387);
xnor U851 (N_851,In_735,In_901);
nand U852 (N_852,In_240,In_1587);
and U853 (N_853,In_1977,In_2463);
xnor U854 (N_854,In_1151,In_2195);
and U855 (N_855,In_1397,In_1753);
nor U856 (N_856,In_235,In_1021);
or U857 (N_857,In_128,In_1908);
nand U858 (N_858,In_1073,In_500);
or U859 (N_859,In_1245,In_237);
xnor U860 (N_860,In_1013,In_1748);
nand U861 (N_861,In_1360,In_487);
xor U862 (N_862,In_2369,In_2439);
xor U863 (N_863,In_1155,In_20);
and U864 (N_864,In_946,In_871);
nand U865 (N_865,In_1721,In_2488);
nor U866 (N_866,In_2118,In_966);
and U867 (N_867,In_2191,In_1487);
or U868 (N_868,In_69,In_506);
nor U869 (N_869,In_180,In_1751);
nand U870 (N_870,In_992,In_1666);
and U871 (N_871,In_1824,In_692);
and U872 (N_872,In_432,In_757);
nand U873 (N_873,In_1250,In_112);
nand U874 (N_874,In_868,In_384);
nor U875 (N_875,In_1934,In_1376);
xnor U876 (N_876,In_2453,In_1320);
nand U877 (N_877,In_1696,In_1969);
nor U878 (N_878,In_2265,In_1286);
xnor U879 (N_879,In_2152,In_1302);
nand U880 (N_880,In_2169,In_684);
nor U881 (N_881,In_631,In_1400);
and U882 (N_882,In_621,In_702);
nor U883 (N_883,In_585,In_818);
and U884 (N_884,In_916,In_1503);
or U885 (N_885,In_1351,In_1736);
and U886 (N_886,In_2334,In_1926);
nor U887 (N_887,In_2428,In_1446);
xor U888 (N_888,In_19,In_1652);
xor U889 (N_889,In_1093,In_817);
or U890 (N_890,In_1292,In_1932);
xnor U891 (N_891,In_273,In_2390);
nor U892 (N_892,In_2022,In_668);
or U893 (N_893,In_957,In_2119);
nand U894 (N_894,In_846,In_270);
or U895 (N_895,In_607,In_2060);
nor U896 (N_896,In_834,In_485);
or U897 (N_897,In_2238,In_2381);
and U898 (N_898,In_56,In_82);
xnor U899 (N_899,In_1428,In_331);
nand U900 (N_900,In_1466,In_1411);
or U901 (N_901,In_1276,In_1822);
nand U902 (N_902,In_905,In_173);
xor U903 (N_903,In_1236,In_60);
and U904 (N_904,In_2477,In_623);
xnor U905 (N_905,In_1586,In_1210);
or U906 (N_906,In_425,In_510);
and U907 (N_907,In_521,In_1728);
xnor U908 (N_908,In_2394,In_2492);
xnor U909 (N_909,In_2223,In_743);
and U910 (N_910,In_709,In_327);
and U911 (N_911,In_1356,In_1220);
and U912 (N_912,In_840,In_548);
nor U913 (N_913,In_862,In_1003);
xor U914 (N_914,In_2402,In_249);
and U915 (N_915,In_496,In_98);
or U916 (N_916,In_269,In_1074);
or U917 (N_917,In_2384,In_1295);
and U918 (N_918,In_1536,In_689);
or U919 (N_919,In_1144,In_1448);
or U920 (N_920,In_555,In_2350);
or U921 (N_921,In_1870,In_191);
nand U922 (N_922,In_991,In_533);
nor U923 (N_923,In_1414,In_209);
nand U924 (N_924,In_990,In_1260);
nor U925 (N_925,In_815,In_1518);
and U926 (N_926,In_1529,In_353);
nor U927 (N_927,In_985,In_477);
nand U928 (N_928,In_2318,In_155);
xor U929 (N_929,In_1483,In_1410);
nand U930 (N_930,In_1808,In_863);
or U931 (N_931,In_1246,In_1329);
xnor U932 (N_932,In_2212,In_1046);
nor U933 (N_933,In_794,In_1189);
xor U934 (N_934,In_1614,In_1077);
nor U935 (N_935,In_127,In_1202);
nand U936 (N_936,In_81,In_805);
nor U937 (N_937,In_1115,In_600);
nor U938 (N_938,In_441,In_1040);
and U939 (N_939,In_1438,In_861);
nand U940 (N_940,In_2063,In_899);
nand U941 (N_941,In_1289,In_1332);
nand U942 (N_942,In_780,In_1061);
xnor U943 (N_943,In_935,In_2449);
xor U944 (N_944,In_1453,In_309);
nand U945 (N_945,In_1215,In_283);
or U946 (N_946,In_1125,In_2053);
or U947 (N_947,In_1378,In_544);
nor U948 (N_948,In_2137,In_2049);
or U949 (N_949,In_747,In_955);
xor U950 (N_950,In_380,In_1526);
xnor U951 (N_951,In_980,In_114);
or U952 (N_952,In_1122,In_2017);
and U953 (N_953,In_1915,In_1923);
nor U954 (N_954,In_250,In_1938);
xor U955 (N_955,In_1147,In_1913);
or U956 (N_956,In_1476,In_930);
and U957 (N_957,In_478,In_1313);
xor U958 (N_958,In_328,In_1837);
or U959 (N_959,In_2465,In_597);
and U960 (N_960,In_1464,In_1806);
xnor U961 (N_961,In_2170,In_643);
nand U962 (N_962,In_2385,In_1330);
nor U963 (N_963,In_348,In_849);
nor U964 (N_964,In_2272,In_1338);
nand U965 (N_965,In_522,In_710);
or U966 (N_966,In_1000,In_1234);
and U967 (N_967,In_640,In_885);
nand U968 (N_968,In_1546,In_906);
or U969 (N_969,In_2431,In_2008);
xnor U970 (N_970,In_253,In_341);
xnor U971 (N_971,In_2457,In_1055);
xnor U972 (N_972,In_768,In_1838);
nand U973 (N_973,In_864,In_1171);
xnor U974 (N_974,In_1287,In_1577);
and U975 (N_975,In_1811,In_226);
nor U976 (N_976,In_377,In_2036);
nor U977 (N_977,In_1335,In_1568);
and U978 (N_978,In_859,In_841);
xor U979 (N_979,In_1622,In_295);
or U980 (N_980,In_754,In_2491);
nor U981 (N_981,In_2253,In_1440);
nor U982 (N_982,In_397,In_1136);
nor U983 (N_983,In_664,In_2273);
nor U984 (N_984,In_31,In_1863);
and U985 (N_985,In_2417,In_1354);
and U986 (N_986,In_2214,In_304);
and U987 (N_987,In_1227,In_622);
or U988 (N_988,In_1785,In_1818);
nor U989 (N_989,In_680,In_605);
or U990 (N_990,In_2441,In_634);
or U991 (N_991,In_646,In_1692);
and U992 (N_992,In_437,In_193);
and U993 (N_993,In_1661,In_2481);
xor U994 (N_994,In_1659,In_773);
and U995 (N_995,In_2395,In_1337);
nand U996 (N_996,In_1224,In_1566);
or U997 (N_997,In_795,In_1619);
or U998 (N_998,In_79,In_2181);
and U999 (N_999,In_317,In_763);
and U1000 (N_1000,In_386,In_599);
nand U1001 (N_1001,In_330,In_573);
nand U1002 (N_1002,In_2412,In_405);
nor U1003 (N_1003,In_286,In_1444);
xor U1004 (N_1004,In_1902,In_251);
nor U1005 (N_1005,In_1752,In_1193);
nand U1006 (N_1006,In_1269,In_1617);
nor U1007 (N_1007,In_770,In_417);
xnor U1008 (N_1008,In_427,In_2365);
nand U1009 (N_1009,In_1352,In_2376);
or U1010 (N_1010,In_2030,In_1180);
or U1011 (N_1011,In_175,In_73);
xor U1012 (N_1012,In_882,In_164);
or U1013 (N_1013,In_265,In_1796);
xnor U1014 (N_1014,In_1249,In_2035);
and U1015 (N_1015,In_99,In_1879);
or U1016 (N_1016,In_2083,In_2059);
or U1017 (N_1017,In_2047,In_1456);
and U1018 (N_1018,In_2023,In_2233);
nand U1019 (N_1019,In_1445,In_2015);
and U1020 (N_1020,In_2203,In_705);
xnor U1021 (N_1021,In_1078,In_1928);
and U1022 (N_1022,In_264,In_2167);
nor U1023 (N_1023,In_541,In_2098);
nand U1024 (N_1024,In_922,In_2444);
nor U1025 (N_1025,In_1383,In_1154);
or U1026 (N_1026,In_2132,In_1367);
nand U1027 (N_1027,In_1775,In_211);
xnor U1028 (N_1028,In_896,In_2161);
nor U1029 (N_1029,In_1602,In_765);
and U1030 (N_1030,In_1420,In_2045);
nor U1031 (N_1031,In_61,In_1729);
or U1032 (N_1032,In_529,In_217);
nor U1033 (N_1033,In_1052,In_1649);
xor U1034 (N_1034,In_495,In_504);
and U1035 (N_1035,In_46,In_1992);
nor U1036 (N_1036,In_416,In_1738);
nand U1037 (N_1037,In_1118,In_361);
and U1038 (N_1038,In_1069,In_113);
or U1039 (N_1039,In_2378,In_234);
xor U1040 (N_1040,In_539,In_287);
nor U1041 (N_1041,In_875,In_1584);
nor U1042 (N_1042,In_1528,In_1179);
xnor U1043 (N_1043,In_1615,In_1976);
nor U1044 (N_1044,In_583,In_1478);
xnor U1045 (N_1045,In_2094,In_745);
xnor U1046 (N_1046,In_2473,In_1961);
and U1047 (N_1047,In_1763,In_2177);
or U1048 (N_1048,In_1278,In_2048);
nand U1049 (N_1049,In_1382,In_1049);
nand U1050 (N_1050,In_742,In_344);
or U1051 (N_1051,In_2136,In_271);
xnor U1052 (N_1052,In_2361,In_285);
nand U1053 (N_1053,In_1631,In_802);
or U1054 (N_1054,In_566,In_189);
xnor U1055 (N_1055,In_37,In_1884);
or U1056 (N_1056,In_1326,In_385);
and U1057 (N_1057,In_165,In_409);
nor U1058 (N_1058,In_2196,In_1995);
nand U1059 (N_1059,In_1946,In_825);
nor U1060 (N_1060,In_2267,In_214);
xnor U1061 (N_1061,In_2117,In_2004);
and U1062 (N_1062,In_2012,In_1761);
nor U1063 (N_1063,In_438,In_154);
and U1064 (N_1064,In_2111,In_655);
or U1065 (N_1065,In_51,In_589);
nor U1066 (N_1066,In_34,In_415);
and U1067 (N_1067,In_1882,In_1911);
nand U1068 (N_1068,In_2461,In_2328);
or U1069 (N_1069,In_1871,In_1142);
xor U1070 (N_1070,In_2084,In_2259);
nand U1071 (N_1071,In_1860,In_1839);
and U1072 (N_1072,In_2135,In_1120);
and U1073 (N_1073,In_1435,In_2346);
or U1074 (N_1074,In_1132,In_880);
nand U1075 (N_1075,In_987,In_777);
and U1076 (N_1076,In_2420,In_1417);
xor U1077 (N_1077,In_1090,In_2189);
and U1078 (N_1078,In_471,In_1218);
and U1079 (N_1079,In_670,In_1759);
xor U1080 (N_1080,In_1689,In_575);
nand U1081 (N_1081,In_2422,In_565);
and U1082 (N_1082,In_294,In_435);
or U1083 (N_1083,In_1554,In_964);
nor U1084 (N_1084,In_697,In_2290);
and U1085 (N_1085,In_2410,In_143);
nand U1086 (N_1086,In_844,In_1472);
xor U1087 (N_1087,In_2283,In_1853);
and U1088 (N_1088,In_1919,In_732);
xor U1089 (N_1089,In_2174,In_2311);
or U1090 (N_1090,In_1669,In_508);
or U1091 (N_1091,In_140,In_1931);
nand U1092 (N_1092,In_153,In_2337);
nand U1093 (N_1093,In_2128,In_983);
nand U1094 (N_1094,In_1485,In_2312);
nand U1095 (N_1095,In_1835,In_400);
nand U1096 (N_1096,In_1370,In_2133);
xnor U1097 (N_1097,In_1490,In_122);
and U1098 (N_1098,In_507,In_591);
or U1099 (N_1099,In_310,In_2288);
xnor U1100 (N_1100,In_1226,In_1358);
xor U1101 (N_1101,In_943,In_443);
nor U1102 (N_1102,In_422,In_1116);
xnor U1103 (N_1103,In_1209,In_2046);
nor U1104 (N_1104,In_737,In_1460);
xor U1105 (N_1105,In_1996,In_1469);
and U1106 (N_1106,In_952,In_2451);
nor U1107 (N_1107,In_1744,In_1238);
nand U1108 (N_1108,In_910,In_1864);
xor U1109 (N_1109,In_1317,In_1927);
or U1110 (N_1110,In_913,In_2447);
xnor U1111 (N_1111,In_1521,In_934);
and U1112 (N_1112,In_740,In_1471);
nand U1113 (N_1113,In_1368,In_919);
and U1114 (N_1114,In_1958,In_2249);
nor U1115 (N_1115,In_1733,In_187);
nand U1116 (N_1116,In_2064,In_917);
and U1117 (N_1117,In_1707,In_1327);
nand U1118 (N_1118,In_293,In_1190);
or U1119 (N_1119,In_772,In_1275);
xnor U1120 (N_1120,In_736,In_324);
nand U1121 (N_1121,In_403,In_520);
or U1122 (N_1122,In_1433,In_459);
or U1123 (N_1123,In_2347,In_2254);
nand U1124 (N_1124,In_719,In_1160);
xnor U1125 (N_1125,In_498,In_1012);
or U1126 (N_1126,In_1392,In_1844);
xnor U1127 (N_1127,In_1867,In_2100);
nand U1128 (N_1128,In_1654,In_959);
nor U1129 (N_1129,In_2142,In_1593);
nor U1130 (N_1130,In_2432,In_2041);
nand U1131 (N_1131,In_2058,In_829);
xnor U1132 (N_1132,In_505,In_518);
nor U1133 (N_1133,In_1016,In_1840);
xnor U1134 (N_1134,In_2076,In_1789);
or U1135 (N_1135,In_1388,In_321);
or U1136 (N_1136,In_725,In_44);
or U1137 (N_1137,In_2121,In_71);
and U1138 (N_1138,In_774,In_1082);
xor U1139 (N_1139,In_1112,In_1900);
nor U1140 (N_1140,In_1993,In_28);
and U1141 (N_1141,In_2054,In_1206);
or U1142 (N_1142,In_1794,In_2307);
nor U1143 (N_1143,In_1149,In_367);
xnor U1144 (N_1144,In_1426,In_675);
xnor U1145 (N_1145,In_897,In_168);
nor U1146 (N_1146,In_1043,In_80);
or U1147 (N_1147,In_890,In_2339);
and U1148 (N_1148,In_1325,In_1201);
or U1149 (N_1149,In_2486,In_803);
and U1150 (N_1150,In_123,In_364);
nor U1151 (N_1151,In_1607,In_2368);
and U1152 (N_1152,In_610,In_1014);
or U1153 (N_1153,In_2089,In_587);
and U1154 (N_1154,In_2211,In_1141);
or U1155 (N_1155,In_2356,In_1674);
nand U1156 (N_1156,In_2156,In_1412);
xnor U1157 (N_1157,In_2185,In_2331);
or U1158 (N_1158,In_2006,In_1452);
xor U1159 (N_1159,In_601,In_2019);
xnor U1160 (N_1160,In_1555,In_2218);
nand U1161 (N_1161,In_549,In_1767);
xor U1162 (N_1162,In_877,In_1940);
nand U1163 (N_1163,In_1290,In_1660);
nand U1164 (N_1164,In_2340,In_820);
xor U1165 (N_1165,In_540,In_489);
xnor U1166 (N_1166,In_941,In_517);
or U1167 (N_1167,In_2139,In_789);
nor U1168 (N_1168,In_1495,In_1861);
nand U1169 (N_1169,In_1305,In_1896);
and U1170 (N_1170,In_810,In_2370);
or U1171 (N_1171,In_673,In_2281);
and U1172 (N_1172,In_1980,In_1655);
nand U1173 (N_1173,In_1984,In_223);
xnor U1174 (N_1174,In_850,In_826);
nand U1175 (N_1175,In_1704,In_245);
nand U1176 (N_1176,In_1708,In_1300);
or U1177 (N_1177,In_1531,In_551);
nand U1178 (N_1178,In_255,In_290);
xnor U1179 (N_1179,In_1571,In_2245);
or U1180 (N_1180,In_2031,In_467);
and U1181 (N_1181,In_1630,In_2069);
nor U1182 (N_1182,In_1080,In_1361);
or U1183 (N_1183,In_594,In_76);
nand U1184 (N_1184,In_584,In_2229);
and U1185 (N_1185,In_1363,In_895);
nor U1186 (N_1186,In_2231,In_2110);
or U1187 (N_1187,In_755,In_254);
and U1188 (N_1188,In_320,In_1672);
or U1189 (N_1189,In_298,In_5);
or U1190 (N_1190,In_1817,In_1045);
nor U1191 (N_1191,In_1906,In_1641);
xor U1192 (N_1192,In_1998,In_554);
nand U1193 (N_1193,In_1273,In_1904);
nand U1194 (N_1194,In_2445,In_837);
and U1195 (N_1195,In_379,In_1398);
nand U1196 (N_1196,In_2320,In_252);
nand U1197 (N_1197,In_1229,In_968);
nor U1198 (N_1198,In_186,In_311);
nand U1199 (N_1199,In_2393,In_1715);
or U1200 (N_1200,In_1499,In_2068);
xnor U1201 (N_1201,In_1734,In_1549);
nand U1202 (N_1202,In_2269,In_1939);
nor U1203 (N_1203,In_16,In_1562);
xnor U1204 (N_1204,In_2143,In_2289);
nand U1205 (N_1205,In_558,In_2499);
and U1206 (N_1206,In_1037,In_1277);
or U1207 (N_1207,In_658,In_1146);
nor U1208 (N_1208,In_47,In_1530);
xnor U1209 (N_1209,In_2261,In_455);
nand U1210 (N_1210,In_2104,In_865);
nand U1211 (N_1211,In_593,In_976);
nand U1212 (N_1212,In_1066,In_2116);
or U1213 (N_1213,In_119,In_2159);
nand U1214 (N_1214,In_886,In_908);
nand U1215 (N_1215,In_940,In_2353);
or U1216 (N_1216,In_2446,In_629);
nor U1217 (N_1217,In_1519,In_2129);
nand U1218 (N_1218,In_229,In_1255);
and U1219 (N_1219,In_1087,In_2333);
nand U1220 (N_1220,In_2020,In_1178);
xor U1221 (N_1221,In_383,In_2199);
nand U1222 (N_1222,In_1608,In_1903);
or U1223 (N_1223,In_733,In_1960);
nor U1224 (N_1224,In_1009,In_131);
nor U1225 (N_1225,In_1284,In_1997);
or U1226 (N_1226,In_2165,In_2043);
xor U1227 (N_1227,In_433,In_2372);
xnor U1228 (N_1228,In_1823,In_1893);
nand U1229 (N_1229,In_1949,In_2438);
xnor U1230 (N_1230,In_2260,In_2314);
xnor U1231 (N_1231,In_979,In_2209);
nor U1232 (N_1232,In_866,In_707);
xnor U1233 (N_1233,In_1909,In_914);
nand U1234 (N_1234,In_1820,In_356);
nor U1235 (N_1235,In_469,In_59);
or U1236 (N_1236,In_2335,In_2460);
nand U1237 (N_1237,In_158,In_1163);
and U1238 (N_1238,In_1507,In_1603);
or U1239 (N_1239,In_858,In_662);
nor U1240 (N_1240,In_567,In_1979);
xnor U1241 (N_1241,In_236,In_924);
and U1242 (N_1242,In_1781,In_1030);
and U1243 (N_1243,In_2299,In_1192);
xor U1244 (N_1244,In_718,In_278);
nand U1245 (N_1245,In_759,In_766);
xor U1246 (N_1246,In_1534,In_2106);
or U1247 (N_1247,In_1406,In_711);
nand U1248 (N_1248,In_2437,In_1739);
or U1249 (N_1249,In_1312,In_1581);
xor U1250 (N_1250,In_104,In_211);
and U1251 (N_1251,In_1849,In_2240);
xnor U1252 (N_1252,In_391,In_383);
or U1253 (N_1253,In_2352,In_6);
nand U1254 (N_1254,In_1222,In_452);
or U1255 (N_1255,In_705,In_2047);
or U1256 (N_1256,In_1259,In_1859);
xor U1257 (N_1257,In_1073,In_348);
xnor U1258 (N_1258,In_2163,In_375);
and U1259 (N_1259,In_579,In_64);
nand U1260 (N_1260,In_898,In_1169);
xnor U1261 (N_1261,In_1043,In_569);
nand U1262 (N_1262,In_1250,In_6);
or U1263 (N_1263,In_926,In_568);
or U1264 (N_1264,In_1723,In_72);
nor U1265 (N_1265,In_1540,In_603);
xor U1266 (N_1266,In_770,In_1059);
nor U1267 (N_1267,In_2209,In_2489);
nor U1268 (N_1268,In_2027,In_1778);
and U1269 (N_1269,In_1910,In_2093);
and U1270 (N_1270,In_995,In_1218);
nor U1271 (N_1271,In_2445,In_108);
xnor U1272 (N_1272,In_2058,In_1016);
and U1273 (N_1273,In_2053,In_1879);
xor U1274 (N_1274,In_1178,In_1822);
and U1275 (N_1275,In_839,In_1104);
xor U1276 (N_1276,In_792,In_1400);
or U1277 (N_1277,In_1788,In_337);
nor U1278 (N_1278,In_2127,In_283);
nor U1279 (N_1279,In_715,In_159);
or U1280 (N_1280,In_1519,In_200);
nor U1281 (N_1281,In_1509,In_792);
nand U1282 (N_1282,In_567,In_1584);
xnor U1283 (N_1283,In_513,In_478);
xor U1284 (N_1284,In_961,In_1872);
nor U1285 (N_1285,In_1923,In_1540);
and U1286 (N_1286,In_28,In_2463);
or U1287 (N_1287,In_1136,In_1468);
or U1288 (N_1288,In_1547,In_382);
xnor U1289 (N_1289,In_954,In_1087);
nor U1290 (N_1290,In_2197,In_509);
nor U1291 (N_1291,In_1508,In_746);
and U1292 (N_1292,In_2053,In_134);
and U1293 (N_1293,In_1724,In_1990);
or U1294 (N_1294,In_1928,In_1057);
nand U1295 (N_1295,In_727,In_1454);
xnor U1296 (N_1296,In_344,In_2427);
or U1297 (N_1297,In_489,In_1935);
nand U1298 (N_1298,In_1770,In_597);
and U1299 (N_1299,In_218,In_2184);
nand U1300 (N_1300,In_214,In_956);
and U1301 (N_1301,In_248,In_1514);
xnor U1302 (N_1302,In_2055,In_2082);
or U1303 (N_1303,In_287,In_1241);
xnor U1304 (N_1304,In_528,In_1288);
or U1305 (N_1305,In_397,In_73);
xnor U1306 (N_1306,In_562,In_474);
and U1307 (N_1307,In_1851,In_1093);
nor U1308 (N_1308,In_350,In_533);
nand U1309 (N_1309,In_1093,In_1041);
nor U1310 (N_1310,In_2008,In_721);
xor U1311 (N_1311,In_1566,In_898);
nand U1312 (N_1312,In_738,In_961);
nand U1313 (N_1313,In_2215,In_363);
or U1314 (N_1314,In_478,In_26);
nand U1315 (N_1315,In_271,In_762);
nor U1316 (N_1316,In_436,In_116);
nand U1317 (N_1317,In_279,In_407);
and U1318 (N_1318,In_1022,In_2191);
xnor U1319 (N_1319,In_1570,In_1609);
xnor U1320 (N_1320,In_1531,In_2132);
or U1321 (N_1321,In_1986,In_453);
or U1322 (N_1322,In_510,In_986);
nor U1323 (N_1323,In_740,In_268);
nand U1324 (N_1324,In_1746,In_1183);
or U1325 (N_1325,In_69,In_1833);
xor U1326 (N_1326,In_769,In_2416);
nand U1327 (N_1327,In_2180,In_307);
nor U1328 (N_1328,In_536,In_1236);
nor U1329 (N_1329,In_810,In_2125);
nand U1330 (N_1330,In_115,In_838);
nand U1331 (N_1331,In_825,In_296);
and U1332 (N_1332,In_2223,In_1823);
nand U1333 (N_1333,In_1540,In_1180);
and U1334 (N_1334,In_218,In_2042);
nor U1335 (N_1335,In_2092,In_905);
and U1336 (N_1336,In_2320,In_1601);
and U1337 (N_1337,In_517,In_2163);
and U1338 (N_1338,In_815,In_1952);
and U1339 (N_1339,In_1506,In_814);
nand U1340 (N_1340,In_1729,In_1005);
xnor U1341 (N_1341,In_1885,In_938);
or U1342 (N_1342,In_397,In_1663);
nand U1343 (N_1343,In_752,In_239);
xnor U1344 (N_1344,In_1536,In_354);
nor U1345 (N_1345,In_1116,In_535);
and U1346 (N_1346,In_333,In_1803);
and U1347 (N_1347,In_1192,In_1418);
and U1348 (N_1348,In_2131,In_1012);
and U1349 (N_1349,In_863,In_1111);
nor U1350 (N_1350,In_529,In_1137);
nand U1351 (N_1351,In_1014,In_445);
and U1352 (N_1352,In_261,In_614);
xor U1353 (N_1353,In_2363,In_496);
nor U1354 (N_1354,In_1670,In_2374);
and U1355 (N_1355,In_425,In_1669);
or U1356 (N_1356,In_161,In_2152);
xnor U1357 (N_1357,In_1174,In_2317);
nor U1358 (N_1358,In_671,In_948);
nand U1359 (N_1359,In_1393,In_93);
xor U1360 (N_1360,In_460,In_2277);
xnor U1361 (N_1361,In_57,In_2252);
nor U1362 (N_1362,In_190,In_1503);
nor U1363 (N_1363,In_494,In_1514);
and U1364 (N_1364,In_1905,In_1056);
nand U1365 (N_1365,In_2011,In_626);
nand U1366 (N_1366,In_1801,In_17);
nand U1367 (N_1367,In_2437,In_2449);
nor U1368 (N_1368,In_570,In_1298);
nor U1369 (N_1369,In_24,In_2169);
or U1370 (N_1370,In_255,In_1806);
nor U1371 (N_1371,In_160,In_1789);
and U1372 (N_1372,In_377,In_965);
nand U1373 (N_1373,In_1348,In_2289);
or U1374 (N_1374,In_377,In_2455);
nor U1375 (N_1375,In_1576,In_434);
and U1376 (N_1376,In_666,In_1637);
xnor U1377 (N_1377,In_1951,In_2205);
or U1378 (N_1378,In_839,In_2486);
nor U1379 (N_1379,In_1936,In_368);
nand U1380 (N_1380,In_1975,In_465);
nand U1381 (N_1381,In_1283,In_2453);
and U1382 (N_1382,In_1471,In_99);
nor U1383 (N_1383,In_1102,In_1673);
xnor U1384 (N_1384,In_1676,In_596);
or U1385 (N_1385,In_766,In_1856);
and U1386 (N_1386,In_2459,In_1625);
xor U1387 (N_1387,In_2075,In_426);
and U1388 (N_1388,In_2180,In_841);
or U1389 (N_1389,In_1830,In_1081);
nor U1390 (N_1390,In_2150,In_535);
xor U1391 (N_1391,In_1495,In_1217);
and U1392 (N_1392,In_2478,In_1459);
nor U1393 (N_1393,In_1658,In_1721);
and U1394 (N_1394,In_884,In_1346);
and U1395 (N_1395,In_518,In_597);
and U1396 (N_1396,In_65,In_328);
nand U1397 (N_1397,In_1616,In_41);
nand U1398 (N_1398,In_413,In_113);
nand U1399 (N_1399,In_1335,In_1736);
nor U1400 (N_1400,In_2367,In_2259);
nand U1401 (N_1401,In_1769,In_1738);
or U1402 (N_1402,In_737,In_103);
nand U1403 (N_1403,In_586,In_595);
or U1404 (N_1404,In_389,In_1719);
nand U1405 (N_1405,In_1615,In_14);
or U1406 (N_1406,In_713,In_1102);
nand U1407 (N_1407,In_225,In_2423);
and U1408 (N_1408,In_1594,In_912);
nor U1409 (N_1409,In_960,In_351);
and U1410 (N_1410,In_863,In_1163);
nor U1411 (N_1411,In_2143,In_667);
and U1412 (N_1412,In_678,In_2459);
nor U1413 (N_1413,In_194,In_1357);
nand U1414 (N_1414,In_1622,In_56);
nand U1415 (N_1415,In_2415,In_1010);
and U1416 (N_1416,In_1525,In_841);
nor U1417 (N_1417,In_1654,In_1595);
nor U1418 (N_1418,In_498,In_1677);
and U1419 (N_1419,In_1652,In_2057);
nand U1420 (N_1420,In_1045,In_652);
or U1421 (N_1421,In_467,In_1251);
xor U1422 (N_1422,In_971,In_1963);
nor U1423 (N_1423,In_452,In_1424);
and U1424 (N_1424,In_1502,In_1396);
nor U1425 (N_1425,In_997,In_1152);
nand U1426 (N_1426,In_1306,In_2250);
and U1427 (N_1427,In_15,In_1157);
or U1428 (N_1428,In_132,In_1637);
and U1429 (N_1429,In_1513,In_1911);
nand U1430 (N_1430,In_885,In_2148);
nor U1431 (N_1431,In_651,In_2079);
nand U1432 (N_1432,In_2012,In_572);
nor U1433 (N_1433,In_119,In_308);
xnor U1434 (N_1434,In_2281,In_45);
nand U1435 (N_1435,In_939,In_1337);
and U1436 (N_1436,In_879,In_1448);
xor U1437 (N_1437,In_2029,In_427);
nor U1438 (N_1438,In_989,In_508);
nand U1439 (N_1439,In_506,In_670);
or U1440 (N_1440,In_1143,In_291);
xor U1441 (N_1441,In_544,In_1205);
or U1442 (N_1442,In_2078,In_384);
and U1443 (N_1443,In_1996,In_1565);
nand U1444 (N_1444,In_917,In_2274);
nand U1445 (N_1445,In_703,In_1560);
and U1446 (N_1446,In_1863,In_2017);
or U1447 (N_1447,In_347,In_2261);
and U1448 (N_1448,In_1440,In_962);
xor U1449 (N_1449,In_2311,In_1558);
or U1450 (N_1450,In_1016,In_1138);
nand U1451 (N_1451,In_1835,In_432);
and U1452 (N_1452,In_1881,In_179);
nor U1453 (N_1453,In_261,In_903);
or U1454 (N_1454,In_1890,In_1286);
xnor U1455 (N_1455,In_588,In_303);
nor U1456 (N_1456,In_1710,In_2222);
or U1457 (N_1457,In_925,In_1614);
nor U1458 (N_1458,In_2448,In_801);
nand U1459 (N_1459,In_114,In_2282);
nor U1460 (N_1460,In_2321,In_1083);
nor U1461 (N_1461,In_2435,In_2417);
and U1462 (N_1462,In_1445,In_2492);
xor U1463 (N_1463,In_705,In_1445);
or U1464 (N_1464,In_803,In_1462);
or U1465 (N_1465,In_2163,In_1544);
nor U1466 (N_1466,In_947,In_1638);
nand U1467 (N_1467,In_813,In_2218);
nand U1468 (N_1468,In_2168,In_1760);
nor U1469 (N_1469,In_624,In_155);
nor U1470 (N_1470,In_1527,In_484);
xor U1471 (N_1471,In_2369,In_1459);
or U1472 (N_1472,In_2206,In_1589);
xor U1473 (N_1473,In_2170,In_1019);
or U1474 (N_1474,In_312,In_138);
nor U1475 (N_1475,In_1394,In_555);
xnor U1476 (N_1476,In_2106,In_1080);
nor U1477 (N_1477,In_2260,In_1967);
xor U1478 (N_1478,In_1992,In_1781);
xnor U1479 (N_1479,In_1834,In_1666);
or U1480 (N_1480,In_2361,In_1718);
xnor U1481 (N_1481,In_963,In_2368);
or U1482 (N_1482,In_433,In_1433);
or U1483 (N_1483,In_886,In_1255);
nor U1484 (N_1484,In_1495,In_1785);
and U1485 (N_1485,In_1864,In_2252);
nor U1486 (N_1486,In_464,In_1091);
xnor U1487 (N_1487,In_1625,In_2420);
xor U1488 (N_1488,In_938,In_1828);
and U1489 (N_1489,In_1194,In_1993);
nand U1490 (N_1490,In_2441,In_211);
or U1491 (N_1491,In_1412,In_1128);
or U1492 (N_1492,In_342,In_1806);
and U1493 (N_1493,In_1786,In_1638);
nand U1494 (N_1494,In_1879,In_1020);
or U1495 (N_1495,In_575,In_848);
or U1496 (N_1496,In_1712,In_928);
nand U1497 (N_1497,In_317,In_1001);
xor U1498 (N_1498,In_1736,In_65);
nand U1499 (N_1499,In_563,In_1259);
xnor U1500 (N_1500,In_1816,In_2396);
xor U1501 (N_1501,In_818,In_1803);
and U1502 (N_1502,In_1225,In_1707);
nor U1503 (N_1503,In_2052,In_2034);
nand U1504 (N_1504,In_1174,In_680);
nor U1505 (N_1505,In_1224,In_1320);
xor U1506 (N_1506,In_409,In_1502);
nand U1507 (N_1507,In_1249,In_1385);
xnor U1508 (N_1508,In_434,In_1081);
nand U1509 (N_1509,In_311,In_545);
nand U1510 (N_1510,In_1807,In_1564);
and U1511 (N_1511,In_2211,In_2480);
or U1512 (N_1512,In_1966,In_1120);
nand U1513 (N_1513,In_533,In_795);
xor U1514 (N_1514,In_2132,In_774);
and U1515 (N_1515,In_1156,In_1389);
xnor U1516 (N_1516,In_2388,In_1597);
or U1517 (N_1517,In_2208,In_397);
and U1518 (N_1518,In_1339,In_774);
nand U1519 (N_1519,In_331,In_818);
nor U1520 (N_1520,In_1143,In_1019);
xor U1521 (N_1521,In_764,In_2149);
xor U1522 (N_1522,In_1861,In_2398);
nor U1523 (N_1523,In_584,In_685);
and U1524 (N_1524,In_1323,In_1268);
and U1525 (N_1525,In_1408,In_1330);
nand U1526 (N_1526,In_2435,In_2447);
xor U1527 (N_1527,In_1774,In_184);
and U1528 (N_1528,In_2417,In_812);
and U1529 (N_1529,In_554,In_2437);
and U1530 (N_1530,In_679,In_1393);
or U1531 (N_1531,In_1997,In_483);
nand U1532 (N_1532,In_1926,In_651);
nor U1533 (N_1533,In_1582,In_1418);
xor U1534 (N_1534,In_2116,In_1111);
and U1535 (N_1535,In_1273,In_325);
nand U1536 (N_1536,In_1906,In_678);
and U1537 (N_1537,In_540,In_1715);
nand U1538 (N_1538,In_2352,In_843);
nand U1539 (N_1539,In_1863,In_1936);
nand U1540 (N_1540,In_851,In_1906);
or U1541 (N_1541,In_2414,In_1253);
or U1542 (N_1542,In_572,In_1312);
nand U1543 (N_1543,In_1660,In_1276);
nor U1544 (N_1544,In_1095,In_865);
nand U1545 (N_1545,In_2122,In_2426);
nor U1546 (N_1546,In_2198,In_705);
and U1547 (N_1547,In_1906,In_1389);
nand U1548 (N_1548,In_2191,In_2031);
nand U1549 (N_1549,In_2435,In_754);
and U1550 (N_1550,In_27,In_141);
nand U1551 (N_1551,In_2313,In_1586);
nor U1552 (N_1552,In_1517,In_741);
xnor U1553 (N_1553,In_562,In_1149);
or U1554 (N_1554,In_750,In_1149);
nor U1555 (N_1555,In_1188,In_438);
nand U1556 (N_1556,In_392,In_1704);
or U1557 (N_1557,In_2374,In_2383);
and U1558 (N_1558,In_509,In_2286);
nor U1559 (N_1559,In_834,In_608);
nor U1560 (N_1560,In_782,In_1593);
or U1561 (N_1561,In_297,In_1088);
or U1562 (N_1562,In_44,In_201);
xnor U1563 (N_1563,In_2324,In_1082);
or U1564 (N_1564,In_2264,In_1559);
and U1565 (N_1565,In_1603,In_1314);
nand U1566 (N_1566,In_1808,In_812);
or U1567 (N_1567,In_478,In_1807);
nand U1568 (N_1568,In_59,In_1442);
and U1569 (N_1569,In_200,In_1045);
nand U1570 (N_1570,In_2493,In_1997);
or U1571 (N_1571,In_124,In_2269);
and U1572 (N_1572,In_575,In_1473);
nand U1573 (N_1573,In_264,In_1650);
xor U1574 (N_1574,In_2014,In_1254);
xnor U1575 (N_1575,In_2495,In_33);
or U1576 (N_1576,In_1014,In_2207);
nand U1577 (N_1577,In_406,In_1142);
nand U1578 (N_1578,In_370,In_2121);
nor U1579 (N_1579,In_236,In_108);
and U1580 (N_1580,In_62,In_1712);
nand U1581 (N_1581,In_1725,In_354);
nand U1582 (N_1582,In_771,In_2102);
nand U1583 (N_1583,In_151,In_431);
nand U1584 (N_1584,In_268,In_1117);
nand U1585 (N_1585,In_2183,In_2477);
and U1586 (N_1586,In_2449,In_1779);
and U1587 (N_1587,In_407,In_382);
or U1588 (N_1588,In_2265,In_2479);
xor U1589 (N_1589,In_358,In_1183);
xor U1590 (N_1590,In_1961,In_433);
and U1591 (N_1591,In_2250,In_688);
nor U1592 (N_1592,In_1338,In_1082);
nor U1593 (N_1593,In_1391,In_2280);
nor U1594 (N_1594,In_1997,In_1865);
or U1595 (N_1595,In_1673,In_1022);
nand U1596 (N_1596,In_2157,In_276);
nand U1597 (N_1597,In_698,In_980);
nand U1598 (N_1598,In_742,In_579);
or U1599 (N_1599,In_1006,In_2474);
xor U1600 (N_1600,In_1524,In_2241);
and U1601 (N_1601,In_993,In_1237);
or U1602 (N_1602,In_1932,In_621);
nor U1603 (N_1603,In_2132,In_842);
xor U1604 (N_1604,In_1894,In_2242);
nand U1605 (N_1605,In_1046,In_39);
and U1606 (N_1606,In_282,In_1957);
or U1607 (N_1607,In_727,In_1825);
nor U1608 (N_1608,In_173,In_2372);
and U1609 (N_1609,In_1354,In_2258);
or U1610 (N_1610,In_1370,In_367);
nor U1611 (N_1611,In_1443,In_1205);
nand U1612 (N_1612,In_61,In_699);
or U1613 (N_1613,In_329,In_283);
nor U1614 (N_1614,In_323,In_1420);
and U1615 (N_1615,In_1995,In_615);
or U1616 (N_1616,In_1991,In_1261);
nand U1617 (N_1617,In_1554,In_635);
or U1618 (N_1618,In_1801,In_374);
nor U1619 (N_1619,In_1294,In_748);
xnor U1620 (N_1620,In_713,In_1753);
xnor U1621 (N_1621,In_1431,In_700);
and U1622 (N_1622,In_1914,In_156);
nor U1623 (N_1623,In_318,In_949);
nor U1624 (N_1624,In_793,In_1269);
and U1625 (N_1625,In_1427,In_45);
nand U1626 (N_1626,In_976,In_1464);
and U1627 (N_1627,In_264,In_304);
and U1628 (N_1628,In_2409,In_1176);
or U1629 (N_1629,In_2487,In_1145);
nand U1630 (N_1630,In_969,In_1729);
xnor U1631 (N_1631,In_722,In_583);
nor U1632 (N_1632,In_711,In_305);
or U1633 (N_1633,In_293,In_348);
nand U1634 (N_1634,In_1896,In_1411);
nand U1635 (N_1635,In_2406,In_1292);
or U1636 (N_1636,In_650,In_1662);
or U1637 (N_1637,In_1931,In_562);
nor U1638 (N_1638,In_854,In_1478);
or U1639 (N_1639,In_725,In_2437);
nand U1640 (N_1640,In_622,In_1436);
and U1641 (N_1641,In_244,In_2368);
and U1642 (N_1642,In_2378,In_368);
xor U1643 (N_1643,In_2293,In_2325);
and U1644 (N_1644,In_2014,In_1838);
and U1645 (N_1645,In_577,In_1405);
or U1646 (N_1646,In_2462,In_10);
nor U1647 (N_1647,In_163,In_724);
nor U1648 (N_1648,In_980,In_544);
nand U1649 (N_1649,In_775,In_359);
or U1650 (N_1650,In_2185,In_1071);
nand U1651 (N_1651,In_238,In_1796);
nor U1652 (N_1652,In_1940,In_1883);
or U1653 (N_1653,In_1734,In_452);
nand U1654 (N_1654,In_772,In_2435);
or U1655 (N_1655,In_649,In_2400);
xnor U1656 (N_1656,In_965,In_188);
and U1657 (N_1657,In_2104,In_715);
nor U1658 (N_1658,In_714,In_2075);
or U1659 (N_1659,In_1902,In_308);
and U1660 (N_1660,In_198,In_570);
nand U1661 (N_1661,In_105,In_1561);
nand U1662 (N_1662,In_1452,In_1387);
nor U1663 (N_1663,In_1038,In_1788);
or U1664 (N_1664,In_1414,In_2470);
and U1665 (N_1665,In_1845,In_1885);
nand U1666 (N_1666,In_1092,In_2047);
and U1667 (N_1667,In_1498,In_346);
or U1668 (N_1668,In_1990,In_257);
nand U1669 (N_1669,In_14,In_748);
or U1670 (N_1670,In_1679,In_937);
or U1671 (N_1671,In_2128,In_2079);
nand U1672 (N_1672,In_456,In_1059);
xnor U1673 (N_1673,In_118,In_995);
nor U1674 (N_1674,In_1168,In_2002);
nor U1675 (N_1675,In_1627,In_1970);
nand U1676 (N_1676,In_2327,In_1003);
nand U1677 (N_1677,In_2416,In_1593);
nand U1678 (N_1678,In_1254,In_2351);
nor U1679 (N_1679,In_1203,In_852);
xnor U1680 (N_1680,In_59,In_1651);
nand U1681 (N_1681,In_46,In_2286);
or U1682 (N_1682,In_624,In_1515);
or U1683 (N_1683,In_456,In_1323);
or U1684 (N_1684,In_2103,In_1456);
and U1685 (N_1685,In_1470,In_2318);
or U1686 (N_1686,In_609,In_1528);
or U1687 (N_1687,In_887,In_77);
and U1688 (N_1688,In_425,In_553);
xnor U1689 (N_1689,In_275,In_1714);
and U1690 (N_1690,In_1440,In_664);
nand U1691 (N_1691,In_1309,In_2449);
nand U1692 (N_1692,In_705,In_744);
nor U1693 (N_1693,In_1047,In_1487);
xor U1694 (N_1694,In_559,In_2061);
and U1695 (N_1695,In_528,In_1557);
nor U1696 (N_1696,In_1373,In_471);
xnor U1697 (N_1697,In_2427,In_1482);
nand U1698 (N_1698,In_1440,In_849);
nand U1699 (N_1699,In_649,In_1366);
or U1700 (N_1700,In_574,In_508);
nand U1701 (N_1701,In_1107,In_421);
and U1702 (N_1702,In_795,In_318);
nand U1703 (N_1703,In_1723,In_443);
xnor U1704 (N_1704,In_713,In_485);
and U1705 (N_1705,In_655,In_1881);
nor U1706 (N_1706,In_241,In_156);
xnor U1707 (N_1707,In_1541,In_1341);
xor U1708 (N_1708,In_1300,In_1850);
and U1709 (N_1709,In_1505,In_1395);
or U1710 (N_1710,In_735,In_1090);
xor U1711 (N_1711,In_1577,In_1348);
and U1712 (N_1712,In_2252,In_1577);
nand U1713 (N_1713,In_1007,In_324);
nand U1714 (N_1714,In_377,In_1711);
nand U1715 (N_1715,In_1182,In_1597);
nand U1716 (N_1716,In_2436,In_1131);
nand U1717 (N_1717,In_2267,In_1576);
nand U1718 (N_1718,In_1007,In_749);
nand U1719 (N_1719,In_2186,In_1899);
nor U1720 (N_1720,In_1231,In_1489);
or U1721 (N_1721,In_1765,In_1417);
xor U1722 (N_1722,In_163,In_511);
or U1723 (N_1723,In_2306,In_345);
or U1724 (N_1724,In_2120,In_1740);
nand U1725 (N_1725,In_333,In_1777);
or U1726 (N_1726,In_53,In_2322);
or U1727 (N_1727,In_702,In_784);
nand U1728 (N_1728,In_1019,In_2031);
nand U1729 (N_1729,In_1360,In_1926);
nand U1730 (N_1730,In_936,In_2487);
xnor U1731 (N_1731,In_2019,In_726);
or U1732 (N_1732,In_1469,In_50);
nand U1733 (N_1733,In_725,In_167);
xnor U1734 (N_1734,In_1606,In_2386);
and U1735 (N_1735,In_536,In_281);
or U1736 (N_1736,In_1591,In_1763);
xnor U1737 (N_1737,In_44,In_1613);
or U1738 (N_1738,In_797,In_2486);
or U1739 (N_1739,In_1716,In_877);
or U1740 (N_1740,In_636,In_1934);
nor U1741 (N_1741,In_1611,In_850);
xor U1742 (N_1742,In_1802,In_468);
xnor U1743 (N_1743,In_1227,In_2040);
and U1744 (N_1744,In_1156,In_873);
xor U1745 (N_1745,In_508,In_1839);
xor U1746 (N_1746,In_1188,In_1200);
nand U1747 (N_1747,In_2080,In_2173);
or U1748 (N_1748,In_1628,In_2485);
or U1749 (N_1749,In_2381,In_2386);
nor U1750 (N_1750,In_2060,In_1916);
and U1751 (N_1751,In_2437,In_1611);
nand U1752 (N_1752,In_2039,In_1785);
and U1753 (N_1753,In_951,In_360);
nand U1754 (N_1754,In_33,In_2342);
and U1755 (N_1755,In_527,In_2168);
and U1756 (N_1756,In_1218,In_1308);
nand U1757 (N_1757,In_1409,In_2030);
and U1758 (N_1758,In_1968,In_337);
nor U1759 (N_1759,In_2355,In_38);
nor U1760 (N_1760,In_143,In_1827);
nor U1761 (N_1761,In_1243,In_1143);
nor U1762 (N_1762,In_2114,In_1228);
xnor U1763 (N_1763,In_764,In_61);
xnor U1764 (N_1764,In_2325,In_2199);
xnor U1765 (N_1765,In_1119,In_1387);
or U1766 (N_1766,In_296,In_1770);
or U1767 (N_1767,In_942,In_1403);
nor U1768 (N_1768,In_2236,In_362);
nand U1769 (N_1769,In_2197,In_2127);
nor U1770 (N_1770,In_945,In_1672);
and U1771 (N_1771,In_992,In_819);
nor U1772 (N_1772,In_949,In_798);
nor U1773 (N_1773,In_603,In_1286);
or U1774 (N_1774,In_513,In_685);
and U1775 (N_1775,In_1560,In_1658);
nand U1776 (N_1776,In_1366,In_2059);
nand U1777 (N_1777,In_2049,In_2242);
nand U1778 (N_1778,In_592,In_1148);
nand U1779 (N_1779,In_1464,In_943);
nor U1780 (N_1780,In_985,In_973);
xnor U1781 (N_1781,In_2013,In_1885);
or U1782 (N_1782,In_310,In_2180);
nand U1783 (N_1783,In_1690,In_2216);
nor U1784 (N_1784,In_477,In_2255);
and U1785 (N_1785,In_594,In_1525);
xnor U1786 (N_1786,In_2342,In_377);
nor U1787 (N_1787,In_194,In_2091);
nand U1788 (N_1788,In_2155,In_1054);
nand U1789 (N_1789,In_604,In_1469);
or U1790 (N_1790,In_1417,In_206);
and U1791 (N_1791,In_2371,In_302);
xnor U1792 (N_1792,In_1681,In_1787);
xor U1793 (N_1793,In_237,In_657);
and U1794 (N_1794,In_835,In_2401);
nor U1795 (N_1795,In_1993,In_990);
or U1796 (N_1796,In_123,In_389);
nor U1797 (N_1797,In_7,In_1035);
xnor U1798 (N_1798,In_883,In_1084);
and U1799 (N_1799,In_2334,In_16);
nor U1800 (N_1800,In_2391,In_1643);
or U1801 (N_1801,In_65,In_803);
or U1802 (N_1802,In_2262,In_2088);
nor U1803 (N_1803,In_202,In_2080);
xor U1804 (N_1804,In_2201,In_858);
xor U1805 (N_1805,In_1852,In_474);
nor U1806 (N_1806,In_2385,In_105);
or U1807 (N_1807,In_1123,In_1364);
xor U1808 (N_1808,In_1599,In_74);
or U1809 (N_1809,In_234,In_460);
nor U1810 (N_1810,In_1663,In_381);
and U1811 (N_1811,In_1141,In_938);
nor U1812 (N_1812,In_669,In_824);
and U1813 (N_1813,In_2027,In_1416);
xor U1814 (N_1814,In_1599,In_2454);
nand U1815 (N_1815,In_2417,In_1050);
and U1816 (N_1816,In_1996,In_265);
nor U1817 (N_1817,In_1136,In_1554);
nor U1818 (N_1818,In_361,In_753);
nand U1819 (N_1819,In_699,In_154);
nand U1820 (N_1820,In_1354,In_836);
or U1821 (N_1821,In_340,In_809);
or U1822 (N_1822,In_220,In_98);
and U1823 (N_1823,In_1213,In_1308);
and U1824 (N_1824,In_831,In_383);
xnor U1825 (N_1825,In_881,In_632);
nor U1826 (N_1826,In_1259,In_71);
nand U1827 (N_1827,In_123,In_2018);
nor U1828 (N_1828,In_478,In_460);
or U1829 (N_1829,In_2496,In_1100);
xor U1830 (N_1830,In_1564,In_555);
nor U1831 (N_1831,In_793,In_558);
xnor U1832 (N_1832,In_7,In_2092);
and U1833 (N_1833,In_1791,In_1584);
xor U1834 (N_1834,In_1278,In_2138);
or U1835 (N_1835,In_2258,In_512);
nor U1836 (N_1836,In_2449,In_195);
nor U1837 (N_1837,In_1230,In_1361);
and U1838 (N_1838,In_114,In_1273);
xor U1839 (N_1839,In_2179,In_280);
and U1840 (N_1840,In_1975,In_2383);
or U1841 (N_1841,In_1192,In_677);
xnor U1842 (N_1842,In_1484,In_1728);
nor U1843 (N_1843,In_1478,In_2434);
xnor U1844 (N_1844,In_838,In_292);
xor U1845 (N_1845,In_41,In_1384);
xnor U1846 (N_1846,In_1358,In_2162);
or U1847 (N_1847,In_1462,In_1474);
nor U1848 (N_1848,In_330,In_1088);
or U1849 (N_1849,In_222,In_1184);
or U1850 (N_1850,In_2240,In_472);
and U1851 (N_1851,In_2032,In_1592);
nor U1852 (N_1852,In_1585,In_2300);
nor U1853 (N_1853,In_1972,In_258);
nand U1854 (N_1854,In_1458,In_2080);
or U1855 (N_1855,In_2019,In_1846);
nand U1856 (N_1856,In_2480,In_2435);
nor U1857 (N_1857,In_1688,In_356);
nand U1858 (N_1858,In_846,In_1780);
and U1859 (N_1859,In_976,In_1415);
or U1860 (N_1860,In_425,In_511);
xnor U1861 (N_1861,In_2,In_2469);
nand U1862 (N_1862,In_2304,In_814);
nand U1863 (N_1863,In_864,In_1042);
nor U1864 (N_1864,In_1679,In_959);
or U1865 (N_1865,In_827,In_1610);
xor U1866 (N_1866,In_1402,In_1626);
nor U1867 (N_1867,In_1172,In_249);
xor U1868 (N_1868,In_1600,In_531);
nand U1869 (N_1869,In_1960,In_2342);
or U1870 (N_1870,In_1254,In_631);
and U1871 (N_1871,In_1693,In_1401);
nor U1872 (N_1872,In_2108,In_86);
xnor U1873 (N_1873,In_2256,In_144);
or U1874 (N_1874,In_2025,In_563);
nor U1875 (N_1875,In_1254,In_1550);
nor U1876 (N_1876,In_1375,In_2372);
and U1877 (N_1877,In_1035,In_850);
xor U1878 (N_1878,In_909,In_1346);
and U1879 (N_1879,In_2165,In_636);
nand U1880 (N_1880,In_361,In_1596);
nand U1881 (N_1881,In_2432,In_2352);
nand U1882 (N_1882,In_1801,In_800);
xor U1883 (N_1883,In_1350,In_2244);
nand U1884 (N_1884,In_1586,In_2081);
and U1885 (N_1885,In_2390,In_2019);
and U1886 (N_1886,In_1092,In_1569);
and U1887 (N_1887,In_143,In_2393);
nor U1888 (N_1888,In_978,In_1061);
xor U1889 (N_1889,In_633,In_861);
xnor U1890 (N_1890,In_2173,In_173);
or U1891 (N_1891,In_1706,In_2463);
or U1892 (N_1892,In_999,In_1522);
nand U1893 (N_1893,In_660,In_510);
or U1894 (N_1894,In_209,In_218);
nor U1895 (N_1895,In_505,In_1624);
nand U1896 (N_1896,In_1093,In_568);
xor U1897 (N_1897,In_2196,In_757);
or U1898 (N_1898,In_250,In_2433);
or U1899 (N_1899,In_717,In_240);
xnor U1900 (N_1900,In_1795,In_1148);
or U1901 (N_1901,In_2008,In_1426);
nand U1902 (N_1902,In_95,In_1323);
nor U1903 (N_1903,In_1128,In_738);
nand U1904 (N_1904,In_5,In_2464);
or U1905 (N_1905,In_1856,In_1252);
nor U1906 (N_1906,In_1606,In_682);
xnor U1907 (N_1907,In_129,In_2051);
nor U1908 (N_1908,In_2273,In_1961);
xor U1909 (N_1909,In_73,In_2112);
xor U1910 (N_1910,In_1939,In_1218);
xnor U1911 (N_1911,In_1720,In_667);
nand U1912 (N_1912,In_434,In_1797);
and U1913 (N_1913,In_898,In_919);
or U1914 (N_1914,In_2317,In_1175);
nor U1915 (N_1915,In_171,In_839);
nor U1916 (N_1916,In_1400,In_379);
nand U1917 (N_1917,In_1731,In_358);
xor U1918 (N_1918,In_1751,In_2215);
xor U1919 (N_1919,In_95,In_1418);
nand U1920 (N_1920,In_2132,In_21);
nand U1921 (N_1921,In_322,In_1656);
nand U1922 (N_1922,In_28,In_2004);
nor U1923 (N_1923,In_1271,In_463);
nand U1924 (N_1924,In_1975,In_288);
or U1925 (N_1925,In_203,In_1756);
or U1926 (N_1926,In_1980,In_2262);
or U1927 (N_1927,In_2258,In_75);
nor U1928 (N_1928,In_920,In_1198);
and U1929 (N_1929,In_2005,In_666);
and U1930 (N_1930,In_2393,In_1431);
nand U1931 (N_1931,In_1730,In_464);
and U1932 (N_1932,In_1451,In_1651);
and U1933 (N_1933,In_1759,In_1221);
xnor U1934 (N_1934,In_1464,In_111);
nor U1935 (N_1935,In_1061,In_2433);
and U1936 (N_1936,In_915,In_1703);
or U1937 (N_1937,In_1206,In_1749);
and U1938 (N_1938,In_2019,In_236);
xor U1939 (N_1939,In_177,In_1647);
or U1940 (N_1940,In_2419,In_2016);
xnor U1941 (N_1941,In_1794,In_277);
xnor U1942 (N_1942,In_1895,In_1491);
xor U1943 (N_1943,In_1130,In_2234);
nor U1944 (N_1944,In_2417,In_1372);
nor U1945 (N_1945,In_1109,In_179);
nor U1946 (N_1946,In_1265,In_421);
or U1947 (N_1947,In_2115,In_590);
nand U1948 (N_1948,In_2371,In_660);
nand U1949 (N_1949,In_1059,In_619);
nor U1950 (N_1950,In_1368,In_629);
and U1951 (N_1951,In_1817,In_599);
nand U1952 (N_1952,In_2426,In_738);
or U1953 (N_1953,In_1349,In_1067);
nor U1954 (N_1954,In_625,In_1383);
xor U1955 (N_1955,In_131,In_2037);
and U1956 (N_1956,In_2308,In_1289);
or U1957 (N_1957,In_1863,In_1354);
and U1958 (N_1958,In_1521,In_2313);
xor U1959 (N_1959,In_629,In_1663);
or U1960 (N_1960,In_1627,In_840);
xnor U1961 (N_1961,In_1517,In_861);
xor U1962 (N_1962,In_1182,In_1531);
nand U1963 (N_1963,In_191,In_712);
nor U1964 (N_1964,In_1246,In_1797);
or U1965 (N_1965,In_2087,In_618);
nor U1966 (N_1966,In_673,In_1654);
xor U1967 (N_1967,In_2034,In_1831);
or U1968 (N_1968,In_2312,In_2227);
xnor U1969 (N_1969,In_1414,In_645);
nor U1970 (N_1970,In_1980,In_2348);
nand U1971 (N_1971,In_1405,In_566);
xor U1972 (N_1972,In_2340,In_1988);
nor U1973 (N_1973,In_2216,In_1370);
nand U1974 (N_1974,In_993,In_1745);
nand U1975 (N_1975,In_1694,In_2293);
and U1976 (N_1976,In_1973,In_2387);
and U1977 (N_1977,In_609,In_2275);
nand U1978 (N_1978,In_2392,In_2352);
xnor U1979 (N_1979,In_119,In_655);
or U1980 (N_1980,In_2085,In_434);
or U1981 (N_1981,In_1854,In_2252);
xnor U1982 (N_1982,In_2412,In_2121);
and U1983 (N_1983,In_180,In_2078);
and U1984 (N_1984,In_820,In_1596);
nand U1985 (N_1985,In_118,In_1030);
and U1986 (N_1986,In_2462,In_2122);
and U1987 (N_1987,In_568,In_2171);
nor U1988 (N_1988,In_2108,In_2218);
nor U1989 (N_1989,In_2053,In_1313);
and U1990 (N_1990,In_1771,In_2120);
and U1991 (N_1991,In_638,In_2078);
and U1992 (N_1992,In_2448,In_1465);
xnor U1993 (N_1993,In_1938,In_1695);
or U1994 (N_1994,In_1690,In_2301);
or U1995 (N_1995,In_49,In_926);
nand U1996 (N_1996,In_74,In_567);
and U1997 (N_1997,In_2442,In_156);
nor U1998 (N_1998,In_889,In_1232);
and U1999 (N_1999,In_1812,In_805);
nor U2000 (N_2000,In_1283,In_545);
or U2001 (N_2001,In_1995,In_300);
xor U2002 (N_2002,In_1026,In_624);
or U2003 (N_2003,In_2140,In_1070);
xor U2004 (N_2004,In_1221,In_2106);
nand U2005 (N_2005,In_332,In_610);
nor U2006 (N_2006,In_2267,In_1772);
nand U2007 (N_2007,In_2422,In_473);
nor U2008 (N_2008,In_78,In_1818);
xor U2009 (N_2009,In_2292,In_271);
nand U2010 (N_2010,In_2411,In_2478);
nor U2011 (N_2011,In_435,In_1425);
xnor U2012 (N_2012,In_947,In_2081);
and U2013 (N_2013,In_325,In_851);
or U2014 (N_2014,In_979,In_1737);
or U2015 (N_2015,In_2237,In_1238);
nand U2016 (N_2016,In_1770,In_1503);
nor U2017 (N_2017,In_1242,In_1086);
and U2018 (N_2018,In_1968,In_1686);
or U2019 (N_2019,In_179,In_1127);
or U2020 (N_2020,In_2378,In_312);
or U2021 (N_2021,In_2237,In_534);
and U2022 (N_2022,In_1215,In_660);
and U2023 (N_2023,In_57,In_1963);
and U2024 (N_2024,In_53,In_864);
or U2025 (N_2025,In_1167,In_329);
nand U2026 (N_2026,In_2082,In_2039);
nand U2027 (N_2027,In_411,In_1024);
nor U2028 (N_2028,In_416,In_323);
nor U2029 (N_2029,In_1410,In_1172);
nor U2030 (N_2030,In_482,In_1646);
xor U2031 (N_2031,In_953,In_1116);
nor U2032 (N_2032,In_1105,In_2476);
nor U2033 (N_2033,In_1997,In_1461);
or U2034 (N_2034,In_1614,In_1756);
nor U2035 (N_2035,In_908,In_267);
and U2036 (N_2036,In_1168,In_1990);
nor U2037 (N_2037,In_1775,In_922);
nand U2038 (N_2038,In_1376,In_343);
or U2039 (N_2039,In_583,In_491);
nor U2040 (N_2040,In_40,In_1142);
nand U2041 (N_2041,In_394,In_180);
or U2042 (N_2042,In_649,In_1);
xor U2043 (N_2043,In_1119,In_1820);
and U2044 (N_2044,In_2271,In_871);
and U2045 (N_2045,In_305,In_3);
nand U2046 (N_2046,In_2489,In_90);
xor U2047 (N_2047,In_2410,In_812);
and U2048 (N_2048,In_695,In_2001);
nand U2049 (N_2049,In_383,In_1101);
or U2050 (N_2050,In_1490,In_2276);
nand U2051 (N_2051,In_1977,In_70);
or U2052 (N_2052,In_2115,In_668);
nand U2053 (N_2053,In_976,In_458);
or U2054 (N_2054,In_886,In_982);
nor U2055 (N_2055,In_83,In_2494);
nand U2056 (N_2056,In_1781,In_1554);
xnor U2057 (N_2057,In_606,In_286);
or U2058 (N_2058,In_647,In_2203);
nand U2059 (N_2059,In_225,In_1033);
nand U2060 (N_2060,In_2340,In_1961);
nor U2061 (N_2061,In_2108,In_2332);
xnor U2062 (N_2062,In_2299,In_767);
xor U2063 (N_2063,In_125,In_948);
nor U2064 (N_2064,In_1772,In_1038);
and U2065 (N_2065,In_1292,In_882);
nor U2066 (N_2066,In_2464,In_2354);
nor U2067 (N_2067,In_880,In_1991);
nand U2068 (N_2068,In_233,In_267);
nand U2069 (N_2069,In_1504,In_827);
or U2070 (N_2070,In_1564,In_2209);
nor U2071 (N_2071,In_1252,In_1654);
nand U2072 (N_2072,In_2033,In_1207);
xnor U2073 (N_2073,In_1531,In_159);
and U2074 (N_2074,In_1425,In_1553);
and U2075 (N_2075,In_1961,In_1693);
xnor U2076 (N_2076,In_1231,In_1736);
or U2077 (N_2077,In_1979,In_1480);
and U2078 (N_2078,In_741,In_391);
and U2079 (N_2079,In_557,In_2061);
nand U2080 (N_2080,In_692,In_1056);
and U2081 (N_2081,In_116,In_4);
and U2082 (N_2082,In_186,In_1649);
xnor U2083 (N_2083,In_1475,In_231);
xor U2084 (N_2084,In_90,In_2498);
and U2085 (N_2085,In_1031,In_1689);
xor U2086 (N_2086,In_437,In_1691);
and U2087 (N_2087,In_1005,In_1958);
or U2088 (N_2088,In_1114,In_1919);
nor U2089 (N_2089,In_272,In_202);
or U2090 (N_2090,In_971,In_1630);
xnor U2091 (N_2091,In_1173,In_350);
nor U2092 (N_2092,In_2181,In_845);
or U2093 (N_2093,In_2278,In_343);
nand U2094 (N_2094,In_1924,In_1584);
or U2095 (N_2095,In_1244,In_589);
or U2096 (N_2096,In_1035,In_2011);
nor U2097 (N_2097,In_1435,In_746);
and U2098 (N_2098,In_1346,In_1370);
nand U2099 (N_2099,In_2122,In_579);
and U2100 (N_2100,In_1548,In_1810);
nand U2101 (N_2101,In_1961,In_96);
and U2102 (N_2102,In_2344,In_1531);
or U2103 (N_2103,In_533,In_531);
xnor U2104 (N_2104,In_2004,In_2298);
or U2105 (N_2105,In_1359,In_1939);
and U2106 (N_2106,In_2027,In_1823);
nor U2107 (N_2107,In_1296,In_1864);
and U2108 (N_2108,In_1605,In_419);
xor U2109 (N_2109,In_23,In_322);
or U2110 (N_2110,In_2379,In_1561);
xnor U2111 (N_2111,In_1473,In_1389);
or U2112 (N_2112,In_2281,In_720);
nand U2113 (N_2113,In_409,In_1371);
xor U2114 (N_2114,In_1725,In_2353);
and U2115 (N_2115,In_1719,In_1094);
or U2116 (N_2116,In_914,In_2156);
nand U2117 (N_2117,In_417,In_260);
and U2118 (N_2118,In_1424,In_1672);
or U2119 (N_2119,In_1048,In_725);
nand U2120 (N_2120,In_1751,In_1713);
or U2121 (N_2121,In_169,In_1668);
nor U2122 (N_2122,In_1000,In_1019);
and U2123 (N_2123,In_1057,In_1041);
xor U2124 (N_2124,In_1616,In_774);
xnor U2125 (N_2125,In_406,In_247);
xor U2126 (N_2126,In_2356,In_1237);
nor U2127 (N_2127,In_2286,In_567);
and U2128 (N_2128,In_2327,In_39);
or U2129 (N_2129,In_20,In_1943);
nor U2130 (N_2130,In_2472,In_1029);
or U2131 (N_2131,In_546,In_1916);
and U2132 (N_2132,In_490,In_601);
and U2133 (N_2133,In_2436,In_1480);
and U2134 (N_2134,In_1830,In_1532);
or U2135 (N_2135,In_2258,In_1718);
or U2136 (N_2136,In_9,In_1237);
or U2137 (N_2137,In_1720,In_1823);
nand U2138 (N_2138,In_1949,In_186);
nand U2139 (N_2139,In_1887,In_1250);
nand U2140 (N_2140,In_802,In_173);
or U2141 (N_2141,In_1411,In_2451);
or U2142 (N_2142,In_1296,In_1728);
nand U2143 (N_2143,In_106,In_431);
or U2144 (N_2144,In_429,In_2114);
or U2145 (N_2145,In_1696,In_382);
or U2146 (N_2146,In_1507,In_202);
xnor U2147 (N_2147,In_1693,In_1041);
nand U2148 (N_2148,In_1111,In_431);
or U2149 (N_2149,In_2211,In_2315);
or U2150 (N_2150,In_943,In_572);
and U2151 (N_2151,In_2205,In_2089);
xnor U2152 (N_2152,In_1289,In_1506);
xnor U2153 (N_2153,In_1498,In_967);
or U2154 (N_2154,In_1780,In_2076);
and U2155 (N_2155,In_1021,In_2433);
nor U2156 (N_2156,In_2449,In_60);
and U2157 (N_2157,In_1555,In_1687);
nand U2158 (N_2158,In_167,In_2482);
and U2159 (N_2159,In_622,In_1689);
or U2160 (N_2160,In_1682,In_2109);
and U2161 (N_2161,In_397,In_1496);
nand U2162 (N_2162,In_1234,In_1467);
nand U2163 (N_2163,In_1608,In_2308);
nor U2164 (N_2164,In_733,In_2387);
xnor U2165 (N_2165,In_1351,In_170);
or U2166 (N_2166,In_1321,In_2025);
xnor U2167 (N_2167,In_2415,In_325);
or U2168 (N_2168,In_264,In_71);
nand U2169 (N_2169,In_1245,In_120);
nor U2170 (N_2170,In_1771,In_1968);
xnor U2171 (N_2171,In_251,In_1491);
nand U2172 (N_2172,In_1805,In_488);
or U2173 (N_2173,In_299,In_1776);
nand U2174 (N_2174,In_1806,In_1994);
nor U2175 (N_2175,In_2110,In_200);
or U2176 (N_2176,In_2161,In_2179);
nor U2177 (N_2177,In_2443,In_1735);
nor U2178 (N_2178,In_1699,In_1157);
xor U2179 (N_2179,In_972,In_1858);
nor U2180 (N_2180,In_670,In_1645);
xnor U2181 (N_2181,In_1864,In_1843);
nor U2182 (N_2182,In_1124,In_1667);
and U2183 (N_2183,In_814,In_2032);
nor U2184 (N_2184,In_1881,In_497);
and U2185 (N_2185,In_1351,In_922);
or U2186 (N_2186,In_1603,In_101);
nand U2187 (N_2187,In_1945,In_342);
nor U2188 (N_2188,In_1143,In_2040);
nor U2189 (N_2189,In_1413,In_2381);
or U2190 (N_2190,In_1748,In_1302);
or U2191 (N_2191,In_857,In_1720);
or U2192 (N_2192,In_114,In_822);
xor U2193 (N_2193,In_813,In_2348);
nand U2194 (N_2194,In_112,In_2481);
and U2195 (N_2195,In_1586,In_2466);
nand U2196 (N_2196,In_1241,In_1220);
and U2197 (N_2197,In_48,In_2098);
nand U2198 (N_2198,In_2211,In_1192);
xor U2199 (N_2199,In_2199,In_26);
and U2200 (N_2200,In_1723,In_2259);
xor U2201 (N_2201,In_1058,In_818);
nor U2202 (N_2202,In_1140,In_567);
or U2203 (N_2203,In_2432,In_1786);
nand U2204 (N_2204,In_900,In_2198);
nand U2205 (N_2205,In_1884,In_1708);
nor U2206 (N_2206,In_794,In_240);
or U2207 (N_2207,In_1254,In_2069);
xor U2208 (N_2208,In_467,In_643);
xnor U2209 (N_2209,In_320,In_773);
nand U2210 (N_2210,In_42,In_630);
nand U2211 (N_2211,In_1936,In_168);
xnor U2212 (N_2212,In_1630,In_2357);
xor U2213 (N_2213,In_185,In_1369);
nor U2214 (N_2214,In_2424,In_1182);
nor U2215 (N_2215,In_1717,In_2415);
nor U2216 (N_2216,In_2474,In_397);
nor U2217 (N_2217,In_2072,In_368);
nor U2218 (N_2218,In_2261,In_986);
nand U2219 (N_2219,In_408,In_1662);
and U2220 (N_2220,In_284,In_1562);
or U2221 (N_2221,In_1108,In_294);
nand U2222 (N_2222,In_2162,In_851);
and U2223 (N_2223,In_70,In_788);
nor U2224 (N_2224,In_251,In_2076);
nor U2225 (N_2225,In_462,In_1107);
nor U2226 (N_2226,In_1904,In_317);
nand U2227 (N_2227,In_1347,In_2342);
or U2228 (N_2228,In_1730,In_1339);
xor U2229 (N_2229,In_2490,In_1461);
xnor U2230 (N_2230,In_1991,In_1386);
nor U2231 (N_2231,In_166,In_1215);
nand U2232 (N_2232,In_2498,In_2348);
or U2233 (N_2233,In_1789,In_1021);
and U2234 (N_2234,In_261,In_476);
nand U2235 (N_2235,In_818,In_2348);
nor U2236 (N_2236,In_637,In_954);
nor U2237 (N_2237,In_1414,In_2070);
nor U2238 (N_2238,In_759,In_1047);
or U2239 (N_2239,In_1614,In_1031);
nor U2240 (N_2240,In_1081,In_824);
or U2241 (N_2241,In_1297,In_2125);
and U2242 (N_2242,In_721,In_2261);
nand U2243 (N_2243,In_758,In_2019);
and U2244 (N_2244,In_1402,In_226);
nand U2245 (N_2245,In_86,In_2489);
nor U2246 (N_2246,In_1778,In_934);
and U2247 (N_2247,In_2366,In_2149);
xnor U2248 (N_2248,In_2175,In_263);
or U2249 (N_2249,In_110,In_513);
or U2250 (N_2250,In_14,In_1109);
or U2251 (N_2251,In_2133,In_1140);
and U2252 (N_2252,In_1405,In_122);
and U2253 (N_2253,In_2158,In_379);
and U2254 (N_2254,In_1639,In_1510);
and U2255 (N_2255,In_2481,In_1071);
or U2256 (N_2256,In_1498,In_1154);
or U2257 (N_2257,In_114,In_82);
nand U2258 (N_2258,In_841,In_1445);
or U2259 (N_2259,In_1295,In_494);
nor U2260 (N_2260,In_925,In_876);
xor U2261 (N_2261,In_717,In_2382);
nor U2262 (N_2262,In_348,In_251);
nand U2263 (N_2263,In_2233,In_2013);
and U2264 (N_2264,In_1678,In_1034);
nand U2265 (N_2265,In_1450,In_397);
xnor U2266 (N_2266,In_1863,In_1113);
and U2267 (N_2267,In_582,In_204);
and U2268 (N_2268,In_227,In_1134);
xor U2269 (N_2269,In_672,In_1307);
xor U2270 (N_2270,In_2409,In_1729);
or U2271 (N_2271,In_1316,In_2292);
and U2272 (N_2272,In_1653,In_78);
nand U2273 (N_2273,In_995,In_671);
nor U2274 (N_2274,In_309,In_458);
and U2275 (N_2275,In_534,In_2287);
nand U2276 (N_2276,In_1940,In_94);
or U2277 (N_2277,In_1290,In_931);
nand U2278 (N_2278,In_283,In_2187);
nor U2279 (N_2279,In_1125,In_1747);
nor U2280 (N_2280,In_941,In_1563);
xor U2281 (N_2281,In_969,In_578);
nor U2282 (N_2282,In_1471,In_716);
nand U2283 (N_2283,In_2012,In_1045);
nor U2284 (N_2284,In_1412,In_879);
or U2285 (N_2285,In_868,In_306);
and U2286 (N_2286,In_2326,In_1506);
xnor U2287 (N_2287,In_1218,In_1473);
nand U2288 (N_2288,In_2245,In_2313);
and U2289 (N_2289,In_539,In_1168);
nor U2290 (N_2290,In_2054,In_1351);
xnor U2291 (N_2291,In_479,In_2288);
and U2292 (N_2292,In_1869,In_1671);
or U2293 (N_2293,In_2464,In_2470);
nand U2294 (N_2294,In_2037,In_2098);
xor U2295 (N_2295,In_1308,In_586);
xor U2296 (N_2296,In_574,In_2116);
xor U2297 (N_2297,In_2147,In_1625);
nor U2298 (N_2298,In_2405,In_1111);
or U2299 (N_2299,In_1771,In_824);
nand U2300 (N_2300,In_1099,In_192);
and U2301 (N_2301,In_1862,In_1309);
and U2302 (N_2302,In_1114,In_836);
nor U2303 (N_2303,In_1621,In_1031);
nor U2304 (N_2304,In_941,In_352);
nor U2305 (N_2305,In_1353,In_1619);
or U2306 (N_2306,In_2095,In_223);
xnor U2307 (N_2307,In_568,In_1017);
nand U2308 (N_2308,In_521,In_1877);
nand U2309 (N_2309,In_1541,In_46);
and U2310 (N_2310,In_1218,In_365);
nor U2311 (N_2311,In_1711,In_1959);
nor U2312 (N_2312,In_1633,In_990);
nor U2313 (N_2313,In_444,In_1624);
nor U2314 (N_2314,In_1895,In_1067);
nor U2315 (N_2315,In_835,In_1651);
and U2316 (N_2316,In_1386,In_136);
or U2317 (N_2317,In_527,In_234);
nand U2318 (N_2318,In_1864,In_199);
nor U2319 (N_2319,In_169,In_924);
xor U2320 (N_2320,In_85,In_280);
xnor U2321 (N_2321,In_2059,In_1400);
nor U2322 (N_2322,In_2055,In_2043);
xor U2323 (N_2323,In_2178,In_1860);
nor U2324 (N_2324,In_1839,In_1757);
and U2325 (N_2325,In_2379,In_1267);
nand U2326 (N_2326,In_189,In_999);
and U2327 (N_2327,In_1444,In_1832);
nor U2328 (N_2328,In_2460,In_2476);
nand U2329 (N_2329,In_718,In_716);
xor U2330 (N_2330,In_2311,In_2175);
nand U2331 (N_2331,In_2260,In_2456);
xor U2332 (N_2332,In_67,In_578);
or U2333 (N_2333,In_1951,In_1631);
nand U2334 (N_2334,In_434,In_2342);
nor U2335 (N_2335,In_125,In_1156);
xnor U2336 (N_2336,In_885,In_1588);
nand U2337 (N_2337,In_1238,In_2443);
and U2338 (N_2338,In_1496,In_222);
xor U2339 (N_2339,In_1295,In_1453);
nor U2340 (N_2340,In_1945,In_1867);
xor U2341 (N_2341,In_2468,In_646);
and U2342 (N_2342,In_2018,In_231);
and U2343 (N_2343,In_963,In_2397);
or U2344 (N_2344,In_767,In_527);
or U2345 (N_2345,In_1555,In_1288);
or U2346 (N_2346,In_2371,In_1394);
or U2347 (N_2347,In_1650,In_772);
nor U2348 (N_2348,In_726,In_410);
and U2349 (N_2349,In_780,In_794);
or U2350 (N_2350,In_1645,In_2102);
xor U2351 (N_2351,In_2110,In_918);
xnor U2352 (N_2352,In_1013,In_601);
xnor U2353 (N_2353,In_635,In_708);
or U2354 (N_2354,In_2182,In_2342);
xor U2355 (N_2355,In_728,In_927);
xor U2356 (N_2356,In_24,In_2355);
nand U2357 (N_2357,In_1645,In_1621);
and U2358 (N_2358,In_2027,In_2318);
or U2359 (N_2359,In_1978,In_166);
nand U2360 (N_2360,In_443,In_2097);
or U2361 (N_2361,In_900,In_269);
and U2362 (N_2362,In_1731,In_1790);
nand U2363 (N_2363,In_162,In_1281);
nor U2364 (N_2364,In_317,In_539);
or U2365 (N_2365,In_178,In_1996);
and U2366 (N_2366,In_2104,In_225);
xor U2367 (N_2367,In_1199,In_1712);
xnor U2368 (N_2368,In_1370,In_1354);
nor U2369 (N_2369,In_235,In_1690);
or U2370 (N_2370,In_2416,In_2390);
nor U2371 (N_2371,In_262,In_396);
or U2372 (N_2372,In_839,In_985);
xor U2373 (N_2373,In_659,In_727);
and U2374 (N_2374,In_341,In_84);
nand U2375 (N_2375,In_329,In_1345);
or U2376 (N_2376,In_668,In_963);
nor U2377 (N_2377,In_2439,In_1460);
xnor U2378 (N_2378,In_1155,In_1574);
nor U2379 (N_2379,In_2375,In_103);
and U2380 (N_2380,In_1183,In_1637);
xor U2381 (N_2381,In_214,In_326);
and U2382 (N_2382,In_2146,In_1073);
or U2383 (N_2383,In_683,In_2114);
nor U2384 (N_2384,In_1600,In_585);
and U2385 (N_2385,In_1757,In_294);
nand U2386 (N_2386,In_1368,In_1302);
nor U2387 (N_2387,In_1544,In_1946);
nor U2388 (N_2388,In_1025,In_2055);
and U2389 (N_2389,In_448,In_1753);
and U2390 (N_2390,In_1302,In_1184);
and U2391 (N_2391,In_1291,In_100);
or U2392 (N_2392,In_934,In_1976);
or U2393 (N_2393,In_1460,In_745);
nand U2394 (N_2394,In_717,In_1371);
or U2395 (N_2395,In_834,In_1146);
nand U2396 (N_2396,In_35,In_25);
nand U2397 (N_2397,In_1891,In_1299);
nand U2398 (N_2398,In_2287,In_1861);
or U2399 (N_2399,In_43,In_1166);
and U2400 (N_2400,In_2289,In_2183);
and U2401 (N_2401,In_1431,In_716);
nand U2402 (N_2402,In_1592,In_1779);
and U2403 (N_2403,In_1770,In_2023);
and U2404 (N_2404,In_968,In_2272);
or U2405 (N_2405,In_2221,In_541);
or U2406 (N_2406,In_402,In_655);
nand U2407 (N_2407,In_304,In_309);
nand U2408 (N_2408,In_1183,In_1838);
nand U2409 (N_2409,In_10,In_1326);
xor U2410 (N_2410,In_9,In_117);
xnor U2411 (N_2411,In_703,In_599);
and U2412 (N_2412,In_318,In_1336);
or U2413 (N_2413,In_1441,In_1519);
and U2414 (N_2414,In_2425,In_257);
nand U2415 (N_2415,In_1605,In_1648);
and U2416 (N_2416,In_1356,In_1322);
xor U2417 (N_2417,In_801,In_2322);
and U2418 (N_2418,In_1539,In_1802);
xnor U2419 (N_2419,In_849,In_81);
xnor U2420 (N_2420,In_516,In_1125);
nand U2421 (N_2421,In_502,In_1319);
nor U2422 (N_2422,In_2103,In_1782);
nand U2423 (N_2423,In_893,In_386);
xnor U2424 (N_2424,In_1009,In_961);
and U2425 (N_2425,In_2366,In_1092);
or U2426 (N_2426,In_1171,In_1549);
nand U2427 (N_2427,In_2118,In_409);
nand U2428 (N_2428,In_1679,In_968);
or U2429 (N_2429,In_2166,In_297);
or U2430 (N_2430,In_1861,In_203);
nand U2431 (N_2431,In_2382,In_2211);
xnor U2432 (N_2432,In_870,In_829);
and U2433 (N_2433,In_2213,In_153);
and U2434 (N_2434,In_1058,In_2333);
and U2435 (N_2435,In_850,In_1343);
nor U2436 (N_2436,In_1079,In_90);
nand U2437 (N_2437,In_225,In_404);
and U2438 (N_2438,In_782,In_1654);
nor U2439 (N_2439,In_1383,In_771);
nand U2440 (N_2440,In_724,In_1142);
or U2441 (N_2441,In_468,In_810);
nand U2442 (N_2442,In_33,In_1239);
nand U2443 (N_2443,In_937,In_2175);
or U2444 (N_2444,In_1546,In_1990);
and U2445 (N_2445,In_2298,In_134);
xnor U2446 (N_2446,In_1766,In_600);
nand U2447 (N_2447,In_923,In_1467);
nor U2448 (N_2448,In_2490,In_2205);
xnor U2449 (N_2449,In_282,In_444);
and U2450 (N_2450,In_1136,In_1278);
xor U2451 (N_2451,In_2315,In_354);
xor U2452 (N_2452,In_947,In_2403);
or U2453 (N_2453,In_2442,In_1212);
nand U2454 (N_2454,In_341,In_2487);
or U2455 (N_2455,In_680,In_2034);
or U2456 (N_2456,In_2053,In_1265);
xor U2457 (N_2457,In_1888,In_1846);
or U2458 (N_2458,In_1107,In_178);
xnor U2459 (N_2459,In_1423,In_413);
nand U2460 (N_2460,In_1280,In_1052);
or U2461 (N_2461,In_2444,In_1959);
and U2462 (N_2462,In_2338,In_403);
nor U2463 (N_2463,In_1731,In_1019);
or U2464 (N_2464,In_1124,In_292);
nand U2465 (N_2465,In_118,In_1492);
nor U2466 (N_2466,In_1816,In_821);
nand U2467 (N_2467,In_353,In_518);
or U2468 (N_2468,In_990,In_350);
nor U2469 (N_2469,In_1408,In_1835);
and U2470 (N_2470,In_1032,In_828);
nor U2471 (N_2471,In_2412,In_121);
nor U2472 (N_2472,In_393,In_1203);
nand U2473 (N_2473,In_2357,In_1855);
xor U2474 (N_2474,In_1601,In_2237);
xor U2475 (N_2475,In_340,In_2413);
xor U2476 (N_2476,In_1387,In_40);
and U2477 (N_2477,In_114,In_1170);
and U2478 (N_2478,In_1409,In_2204);
or U2479 (N_2479,In_1670,In_969);
or U2480 (N_2480,In_839,In_1633);
xor U2481 (N_2481,In_1363,In_1286);
or U2482 (N_2482,In_586,In_933);
and U2483 (N_2483,In_137,In_392);
nand U2484 (N_2484,In_1592,In_326);
or U2485 (N_2485,In_1822,In_2295);
nand U2486 (N_2486,In_900,In_780);
or U2487 (N_2487,In_1420,In_615);
or U2488 (N_2488,In_218,In_2457);
xnor U2489 (N_2489,In_1406,In_256);
nand U2490 (N_2490,In_1943,In_994);
and U2491 (N_2491,In_994,In_564);
or U2492 (N_2492,In_681,In_2088);
nor U2493 (N_2493,In_1866,In_1066);
nand U2494 (N_2494,In_1230,In_137);
or U2495 (N_2495,In_1633,In_1413);
nand U2496 (N_2496,In_1534,In_1879);
or U2497 (N_2497,In_1610,In_1618);
and U2498 (N_2498,In_1228,In_1338);
and U2499 (N_2499,In_878,In_1195);
xnor U2500 (N_2500,N_1419,N_1226);
and U2501 (N_2501,N_1693,N_1434);
nand U2502 (N_2502,N_1130,N_111);
nand U2503 (N_2503,N_1183,N_290);
nand U2504 (N_2504,N_2386,N_1940);
nand U2505 (N_2505,N_2102,N_342);
or U2506 (N_2506,N_562,N_2228);
nor U2507 (N_2507,N_1902,N_1724);
nor U2508 (N_2508,N_2207,N_204);
or U2509 (N_2509,N_386,N_972);
nand U2510 (N_2510,N_30,N_2375);
xor U2511 (N_2511,N_1321,N_1810);
nand U2512 (N_2512,N_1507,N_818);
nor U2513 (N_2513,N_1243,N_289);
or U2514 (N_2514,N_1158,N_1926);
nand U2515 (N_2515,N_406,N_595);
or U2516 (N_2516,N_361,N_1857);
or U2517 (N_2517,N_2193,N_1137);
and U2518 (N_2518,N_1519,N_566);
nor U2519 (N_2519,N_110,N_2463);
and U2520 (N_2520,N_1392,N_945);
or U2521 (N_2521,N_1475,N_2288);
or U2522 (N_2522,N_515,N_554);
xor U2523 (N_2523,N_490,N_1787);
or U2524 (N_2524,N_1399,N_2256);
xor U2525 (N_2525,N_116,N_193);
nand U2526 (N_2526,N_1109,N_636);
nor U2527 (N_2527,N_114,N_2236);
nand U2528 (N_2528,N_2204,N_849);
or U2529 (N_2529,N_2239,N_367);
xor U2530 (N_2530,N_2246,N_2241);
and U2531 (N_2531,N_1887,N_1054);
and U2532 (N_2532,N_1711,N_485);
xor U2533 (N_2533,N_1676,N_2192);
nand U2534 (N_2534,N_684,N_906);
xor U2535 (N_2535,N_1246,N_2251);
xnor U2536 (N_2536,N_890,N_1598);
nand U2537 (N_2537,N_2449,N_1496);
and U2538 (N_2538,N_205,N_1498);
xnor U2539 (N_2539,N_1445,N_26);
nor U2540 (N_2540,N_789,N_2267);
and U2541 (N_2541,N_378,N_502);
nor U2542 (N_2542,N_824,N_2033);
and U2543 (N_2543,N_1479,N_2437);
and U2544 (N_2544,N_94,N_279);
nand U2545 (N_2545,N_301,N_2380);
nor U2546 (N_2546,N_1455,N_846);
and U2547 (N_2547,N_93,N_2493);
or U2548 (N_2548,N_45,N_2230);
nand U2549 (N_2549,N_2101,N_2354);
nor U2550 (N_2550,N_450,N_1710);
nor U2551 (N_2551,N_804,N_1031);
nor U2552 (N_2552,N_447,N_1915);
xor U2553 (N_2553,N_145,N_2289);
and U2554 (N_2554,N_1992,N_1844);
and U2555 (N_2555,N_1248,N_2427);
and U2556 (N_2556,N_210,N_2304);
xor U2557 (N_2557,N_1714,N_1401);
xnor U2558 (N_2558,N_1013,N_1741);
nor U2559 (N_2559,N_1920,N_1324);
or U2560 (N_2560,N_2495,N_2040);
nor U2561 (N_2561,N_27,N_1783);
nand U2562 (N_2562,N_535,N_692);
xnor U2563 (N_2563,N_982,N_2315);
xnor U2564 (N_2564,N_43,N_531);
and U2565 (N_2565,N_320,N_2051);
xnor U2566 (N_2566,N_1612,N_1922);
or U2567 (N_2567,N_1523,N_816);
or U2568 (N_2568,N_2129,N_396);
or U2569 (N_2569,N_984,N_1981);
or U2570 (N_2570,N_1345,N_1422);
xor U2571 (N_2571,N_2374,N_106);
xnor U2572 (N_2572,N_1500,N_932);
or U2573 (N_2573,N_900,N_1092);
nand U2574 (N_2574,N_1313,N_1805);
nor U2575 (N_2575,N_1831,N_1517);
nor U2576 (N_2576,N_476,N_1095);
or U2577 (N_2577,N_2498,N_1826);
and U2578 (N_2578,N_2244,N_619);
nor U2579 (N_2579,N_1188,N_2370);
or U2580 (N_2580,N_1978,N_1378);
and U2581 (N_2581,N_1256,N_1781);
and U2582 (N_2582,N_2297,N_2287);
nor U2583 (N_2583,N_2229,N_1349);
or U2584 (N_2584,N_1795,N_239);
xnor U2585 (N_2585,N_2015,N_1890);
nand U2586 (N_2586,N_503,N_995);
or U2587 (N_2587,N_1493,N_113);
and U2588 (N_2588,N_2003,N_2063);
and U2589 (N_2589,N_395,N_2301);
or U2590 (N_2590,N_676,N_1760);
nor U2591 (N_2591,N_2171,N_181);
or U2592 (N_2592,N_2472,N_1592);
or U2593 (N_2593,N_1719,N_1625);
nand U2594 (N_2594,N_1735,N_861);
or U2595 (N_2595,N_1149,N_1756);
nand U2596 (N_2596,N_1916,N_1855);
nand U2597 (N_2597,N_305,N_1977);
or U2598 (N_2598,N_338,N_50);
nand U2599 (N_2599,N_126,N_1749);
and U2600 (N_2600,N_214,N_381);
xnor U2601 (N_2601,N_2481,N_518);
or U2602 (N_2602,N_702,N_448);
nor U2603 (N_2603,N_2223,N_2064);
xnor U2604 (N_2604,N_39,N_321);
xor U2605 (N_2605,N_546,N_891);
xor U2606 (N_2606,N_1780,N_840);
nand U2607 (N_2607,N_683,N_1545);
xnor U2608 (N_2608,N_48,N_843);
xnor U2609 (N_2609,N_1373,N_937);
nor U2610 (N_2610,N_577,N_913);
and U2611 (N_2611,N_1597,N_1892);
or U2612 (N_2612,N_1495,N_1393);
nand U2613 (N_2613,N_122,N_2181);
or U2614 (N_2614,N_510,N_1274);
and U2615 (N_2615,N_2242,N_1118);
xnor U2616 (N_2616,N_1073,N_1414);
nand U2617 (N_2617,N_1833,N_1836);
or U2618 (N_2618,N_2099,N_47);
and U2619 (N_2619,N_1593,N_1941);
and U2620 (N_2620,N_1570,N_125);
nor U2621 (N_2621,N_1065,N_1117);
or U2622 (N_2622,N_1763,N_825);
xnor U2623 (N_2623,N_1167,N_1652);
nor U2624 (N_2624,N_613,N_2211);
nand U2625 (N_2625,N_1674,N_1453);
xor U2626 (N_2626,N_1871,N_196);
and U2627 (N_2627,N_1609,N_2235);
nor U2628 (N_2628,N_1712,N_2310);
xnor U2629 (N_2629,N_1681,N_408);
nand U2630 (N_2630,N_1869,N_432);
nor U2631 (N_2631,N_1549,N_2306);
nor U2632 (N_2632,N_2172,N_1627);
or U2633 (N_2633,N_155,N_222);
and U2634 (N_2634,N_426,N_2406);
or U2635 (N_2635,N_71,N_271);
nor U2636 (N_2636,N_349,N_1368);
nor U2637 (N_2637,N_249,N_2443);
or U2638 (N_2638,N_57,N_1056);
xor U2639 (N_2639,N_833,N_917);
and U2640 (N_2640,N_969,N_1666);
xor U2641 (N_2641,N_974,N_1264);
nor U2642 (N_2642,N_2458,N_2081);
and U2643 (N_2643,N_2168,N_1728);
nand U2644 (N_2644,N_1485,N_1649);
or U2645 (N_2645,N_1021,N_99);
nand U2646 (N_2646,N_506,N_2035);
nand U2647 (N_2647,N_1911,N_681);
and U2648 (N_2648,N_2319,N_331);
nand U2649 (N_2649,N_1876,N_1071);
nand U2650 (N_2650,N_284,N_1228);
nor U2651 (N_2651,N_1823,N_1829);
nand U2652 (N_2652,N_1987,N_1659);
xor U2653 (N_2653,N_1234,N_938);
nor U2654 (N_2654,N_1342,N_915);
nor U2655 (N_2655,N_2088,N_128);
nor U2656 (N_2656,N_1096,N_673);
nor U2657 (N_2657,N_1743,N_187);
xnor U2658 (N_2658,N_307,N_2065);
nor U2659 (N_2659,N_778,N_763);
and U2660 (N_2660,N_2083,N_1355);
nor U2661 (N_2661,N_1957,N_2143);
or U2662 (N_2662,N_1614,N_2294);
and U2663 (N_2663,N_653,N_295);
or U2664 (N_2664,N_2044,N_884);
or U2665 (N_2665,N_1762,N_1536);
xor U2666 (N_2666,N_324,N_841);
xnor U2667 (N_2667,N_1830,N_1038);
xor U2668 (N_2668,N_527,N_2453);
and U2669 (N_2669,N_2078,N_2212);
nor U2670 (N_2670,N_724,N_1732);
or U2671 (N_2671,N_2265,N_61);
xnor U2672 (N_2672,N_2270,N_903);
or U2673 (N_2673,N_315,N_2014);
nand U2674 (N_2674,N_56,N_1568);
xor U2675 (N_2675,N_2490,N_2048);
and U2676 (N_2676,N_2266,N_2264);
or U2677 (N_2677,N_1837,N_1600);
nand U2678 (N_2678,N_2434,N_596);
nand U2679 (N_2679,N_1824,N_2188);
and U2680 (N_2680,N_2036,N_2324);
or U2681 (N_2681,N_658,N_870);
or U2682 (N_2682,N_1045,N_2426);
and U2683 (N_2683,N_555,N_1472);
xor U2684 (N_2684,N_904,N_1180);
or U2685 (N_2685,N_1591,N_2070);
xor U2686 (N_2686,N_1459,N_2478);
or U2687 (N_2687,N_780,N_1005);
xor U2688 (N_2688,N_1619,N_1971);
and U2689 (N_2689,N_1573,N_1305);
and U2690 (N_2690,N_388,N_2104);
and U2691 (N_2691,N_2414,N_1935);
and U2692 (N_2692,N_1085,N_102);
xor U2693 (N_2693,N_1034,N_2147);
xnor U2694 (N_2694,N_534,N_1776);
xor U2695 (N_2695,N_799,N_512);
and U2696 (N_2696,N_2157,N_1044);
or U2697 (N_2697,N_137,N_465);
and U2698 (N_2698,N_1299,N_2250);
or U2699 (N_2699,N_1825,N_948);
nand U2700 (N_2700,N_1945,N_2119);
nand U2701 (N_2701,N_557,N_2296);
nand U2702 (N_2702,N_678,N_541);
and U2703 (N_2703,N_9,N_1607);
nor U2704 (N_2704,N_1446,N_700);
xor U2705 (N_2705,N_2150,N_2131);
and U2706 (N_2706,N_507,N_2337);
and U2707 (N_2707,N_1564,N_1577);
xor U2708 (N_2708,N_1984,N_1020);
or U2709 (N_2709,N_1557,N_1939);
nor U2710 (N_2710,N_526,N_2077);
or U2711 (N_2711,N_690,N_16);
nor U2712 (N_2712,N_399,N_1288);
or U2713 (N_2713,N_2384,N_729);
xor U2714 (N_2714,N_2118,N_456);
or U2715 (N_2715,N_1567,N_1884);
or U2716 (N_2716,N_1660,N_277);
and U2717 (N_2717,N_1746,N_1552);
and U2718 (N_2718,N_2444,N_885);
nand U2719 (N_2719,N_2072,N_78);
nor U2720 (N_2720,N_144,N_248);
nor U2721 (N_2721,N_1924,N_1185);
or U2722 (N_2722,N_131,N_1931);
and U2723 (N_2723,N_231,N_109);
nor U2724 (N_2724,N_986,N_1949);
or U2725 (N_2725,N_341,N_655);
or U2726 (N_2726,N_4,N_755);
nand U2727 (N_2727,N_1665,N_2291);
or U2728 (N_2728,N_85,N_2046);
xor U2729 (N_2729,N_2402,N_2385);
and U2730 (N_2730,N_537,N_1819);
nand U2731 (N_2731,N_719,N_1662);
and U2732 (N_2732,N_712,N_1974);
and U2733 (N_2733,N_291,N_979);
or U2734 (N_2734,N_784,N_851);
xnor U2735 (N_2735,N_2120,N_2007);
or U2736 (N_2736,N_1302,N_135);
xor U2737 (N_2737,N_2008,N_208);
xor U2738 (N_2738,N_705,N_251);
and U2739 (N_2739,N_2167,N_177);
nor U2740 (N_2740,N_363,N_1141);
or U2741 (N_2741,N_2316,N_2031);
nor U2742 (N_2742,N_1478,N_568);
and U2743 (N_2743,N_6,N_1590);
or U2744 (N_2744,N_521,N_1629);
xor U2745 (N_2745,N_1412,N_159);
xnor U2746 (N_2746,N_740,N_1983);
or U2747 (N_2747,N_1004,N_588);
nor U2748 (N_2748,N_237,N_2473);
xnor U2749 (N_2749,N_1042,N_264);
xnor U2750 (N_2750,N_1370,N_1166);
nor U2751 (N_2751,N_1168,N_1571);
nor U2752 (N_2752,N_1398,N_1522);
nor U2753 (N_2753,N_766,N_244);
nand U2754 (N_2754,N_796,N_978);
and U2755 (N_2755,N_1326,N_940);
and U2756 (N_2756,N_2082,N_1856);
nand U2757 (N_2757,N_2262,N_617);
and U2758 (N_2758,N_2107,N_2344);
and U2759 (N_2759,N_1845,N_779);
nand U2760 (N_2760,N_1734,N_1895);
or U2761 (N_2761,N_887,N_2238);
nand U2762 (N_2762,N_360,N_1508);
nor U2763 (N_2763,N_312,N_1014);
nor U2764 (N_2764,N_594,N_798);
xnor U2765 (N_2765,N_748,N_1956);
and U2766 (N_2766,N_774,N_1903);
xor U2767 (N_2767,N_180,N_793);
or U2768 (N_2768,N_2182,N_1842);
nor U2769 (N_2769,N_1249,N_487);
nor U2770 (N_2770,N_475,N_2276);
or U2771 (N_2771,N_2448,N_1541);
nand U2772 (N_2772,N_2255,N_2069);
or U2773 (N_2773,N_1145,N_860);
or U2774 (N_2774,N_1319,N_169);
xnor U2775 (N_2775,N_136,N_2020);
or U2776 (N_2776,N_11,N_2342);
or U2777 (N_2777,N_115,N_1875);
or U2778 (N_2778,N_22,N_493);
or U2779 (N_2779,N_2432,N_314);
xnor U2780 (N_2780,N_1539,N_8);
nor U2781 (N_2781,N_1272,N_194);
nand U2782 (N_2782,N_2156,N_1);
xor U2783 (N_2783,N_961,N_1794);
or U2784 (N_2784,N_2038,N_2362);
or U2785 (N_2785,N_672,N_2174);
nor U2786 (N_2786,N_384,N_701);
and U2787 (N_2787,N_765,N_2268);
nor U2788 (N_2788,N_1528,N_470);
nor U2789 (N_2789,N_203,N_1242);
and U2790 (N_2790,N_442,N_2429);
xnor U2791 (N_2791,N_2094,N_715);
and U2792 (N_2792,N_198,N_1040);
xor U2793 (N_2793,N_1839,N_1252);
nor U2794 (N_2794,N_394,N_616);
nand U2795 (N_2795,N_1671,N_2488);
or U2796 (N_2796,N_473,N_1360);
or U2797 (N_2797,N_523,N_153);
nand U2798 (N_2798,N_1329,N_1198);
xnor U2799 (N_2799,N_1047,N_964);
and U2800 (N_2800,N_2371,N_1215);
and U2801 (N_2801,N_539,N_1584);
and U2802 (N_2802,N_1051,N_791);
nor U2803 (N_2803,N_649,N_258);
nand U2804 (N_2804,N_556,N_362);
and U2805 (N_2805,N_190,N_2454);
nor U2806 (N_2806,N_1558,N_618);
and U2807 (N_2807,N_1262,N_192);
nor U2808 (N_2808,N_36,N_1306);
xor U2809 (N_2809,N_745,N_727);
nand U2810 (N_2810,N_570,N_5);
nand U2811 (N_2811,N_971,N_662);
xor U2812 (N_2812,N_1260,N_718);
nand U2813 (N_2813,N_786,N_553);
and U2814 (N_2814,N_2253,N_316);
and U2815 (N_2815,N_1025,N_195);
or U2816 (N_2816,N_1807,N_2042);
nor U2817 (N_2817,N_1396,N_1001);
or U2818 (N_2818,N_1730,N_339);
nor U2819 (N_2819,N_832,N_660);
nor U2820 (N_2820,N_1169,N_572);
or U2821 (N_2821,N_1766,N_720);
nand U2822 (N_2822,N_1151,N_455);
xnor U2823 (N_2823,N_1012,N_278);
nor U2824 (N_2824,N_411,N_1041);
and U2825 (N_2825,N_37,N_654);
nand U2826 (N_2826,N_139,N_771);
and U2827 (N_2827,N_533,N_1438);
or U2828 (N_2828,N_872,N_1340);
xnor U2829 (N_2829,N_346,N_1435);
xor U2830 (N_2830,N_648,N_1269);
xnor U2831 (N_2831,N_1864,N_1699);
or U2832 (N_2832,N_1811,N_1174);
nor U2833 (N_2833,N_578,N_2479);
nand U2834 (N_2834,N_1068,N_2201);
nor U2835 (N_2835,N_1411,N_1284);
nand U2836 (N_2836,N_1703,N_1484);
and U2837 (N_2837,N_1524,N_377);
or U2838 (N_2838,N_2079,N_2247);
nand U2839 (N_2839,N_657,N_1947);
or U2840 (N_2840,N_1525,N_348);
and U2841 (N_2841,N_854,N_1880);
and U2842 (N_2842,N_2122,N_1311);
and U2843 (N_2843,N_2368,N_1191);
nor U2844 (N_2844,N_575,N_1337);
xnor U2845 (N_2845,N_2249,N_703);
nor U2846 (N_2846,N_178,N_625);
and U2847 (N_2847,N_1960,N_2160);
xnor U2848 (N_2848,N_2474,N_1521);
and U2849 (N_2849,N_197,N_2019);
or U2850 (N_2850,N_100,N_345);
and U2851 (N_2851,N_1090,N_430);
xnor U2852 (N_2852,N_2237,N_138);
and U2853 (N_2853,N_524,N_1953);
and U2854 (N_2854,N_95,N_2206);
or U2855 (N_2855,N_1292,N_1206);
xor U2856 (N_2856,N_1696,N_445);
and U2857 (N_2857,N_2224,N_319);
and U2858 (N_2858,N_814,N_2058);
or U2859 (N_2859,N_1036,N_2336);
nor U2860 (N_2860,N_1648,N_542);
or U2861 (N_2861,N_1817,N_154);
xnor U2862 (N_2862,N_2299,N_374);
or U2863 (N_2863,N_2343,N_164);
or U2864 (N_2864,N_434,N_2420);
nand U2865 (N_2865,N_1099,N_698);
nor U2866 (N_2866,N_1861,N_2176);
or U2867 (N_2867,N_1008,N_0);
and U2868 (N_2868,N_354,N_260);
and U2869 (N_2869,N_1542,N_635);
or U2870 (N_2870,N_294,N_2293);
xor U2871 (N_2871,N_1750,N_514);
or U2872 (N_2872,N_1616,N_1362);
or U2873 (N_2873,N_888,N_530);
nand U2874 (N_2874,N_1476,N_1127);
and U2875 (N_2875,N_479,N_1661);
nand U2876 (N_2876,N_1146,N_1737);
or U2877 (N_2877,N_1100,N_525);
and U2878 (N_2878,N_983,N_1480);
and U2879 (N_2879,N_1854,N_1063);
nor U2880 (N_2880,N_1963,N_366);
or U2881 (N_2881,N_28,N_943);
or U2882 (N_2882,N_147,N_2381);
nand U2883 (N_2883,N_1413,N_1473);
nand U2884 (N_2884,N_2028,N_246);
nor U2885 (N_2885,N_2018,N_2334);
or U2886 (N_2886,N_1834,N_1372);
or U2887 (N_2887,N_2,N_902);
nand U2888 (N_2888,N_1996,N_1553);
xnor U2889 (N_2889,N_732,N_223);
and U2890 (N_2890,N_2093,N_1820);
and U2891 (N_2891,N_2074,N_412);
nor U2892 (N_2892,N_1154,N_563);
or U2893 (N_2893,N_268,N_547);
and U2894 (N_2894,N_304,N_696);
or U2895 (N_2895,N_768,N_1395);
and U2896 (N_2896,N_544,N_1588);
and U2897 (N_2897,N_1093,N_1513);
xor U2898 (N_2898,N_83,N_2163);
nor U2899 (N_2899,N_357,N_436);
nand U2900 (N_2900,N_1320,N_1230);
and U2901 (N_2901,N_49,N_519);
and U2902 (N_2902,N_2489,N_2450);
or U2903 (N_2903,N_1785,N_808);
xnor U2904 (N_2904,N_340,N_1959);
nor U2905 (N_2905,N_834,N_1777);
nor U2906 (N_2906,N_1487,N_1675);
or U2907 (N_2907,N_2491,N_2209);
xnor U2908 (N_2908,N_1655,N_1123);
and U2909 (N_2909,N_931,N_1143);
nand U2910 (N_2910,N_1658,N_2480);
nor U2911 (N_2911,N_1219,N_2037);
nor U2912 (N_2912,N_723,N_478);
or U2913 (N_2913,N_601,N_695);
or U2914 (N_2914,N_1367,N_127);
or U2915 (N_2915,N_1387,N_880);
xnor U2916 (N_2916,N_2161,N_1813);
nand U2917 (N_2917,N_1173,N_149);
xnor U2918 (N_2918,N_1454,N_1282);
xor U2919 (N_2919,N_767,N_414);
nand U2920 (N_2920,N_669,N_757);
xor U2921 (N_2921,N_172,N_550);
nor U2922 (N_2922,N_589,N_852);
and U2923 (N_2923,N_1175,N_1980);
nor U2924 (N_2924,N_2445,N_1213);
xnor U2925 (N_2925,N_1418,N_1651);
and U2926 (N_2926,N_1181,N_2034);
or U2927 (N_2927,N_944,N_803);
nand U2928 (N_2928,N_1594,N_444);
or U2929 (N_2929,N_87,N_2284);
xnor U2930 (N_2930,N_1618,N_79);
nor U2931 (N_2931,N_2387,N_928);
nor U2932 (N_2932,N_2396,N_1770);
nand U2933 (N_2933,N_1982,N_240);
xor U2934 (N_2934,N_1682,N_1247);
nor U2935 (N_2935,N_1637,N_714);
nor U2936 (N_2936,N_62,N_581);
xor U2937 (N_2937,N_895,N_1443);
nor U2938 (N_2938,N_1170,N_391);
or U2939 (N_2939,N_1502,N_55);
and U2940 (N_2940,N_1804,N_1867);
and U2941 (N_2941,N_645,N_1858);
and U2942 (N_2942,N_1914,N_865);
or U2943 (N_2943,N_337,N_1474);
nand U2944 (N_2944,N_1801,N_2436);
xnor U2945 (N_2945,N_1491,N_746);
nor U2946 (N_2946,N_1503,N_2067);
xnor U2947 (N_2947,N_211,N_400);
xor U2948 (N_2948,N_431,N_760);
nand U2949 (N_2949,N_2350,N_468);
xnor U2950 (N_2950,N_758,N_382);
xnor U2951 (N_2951,N_2467,N_949);
xnor U2952 (N_2952,N_750,N_2043);
or U2953 (N_2953,N_970,N_202);
nand U2954 (N_2954,N_2009,N_2383);
and U2955 (N_2955,N_1335,N_492);
xor U2956 (N_2956,N_1225,N_132);
nor U2957 (N_2957,N_306,N_2363);
and U2958 (N_2958,N_7,N_1037);
nand U2959 (N_2959,N_930,N_269);
nand U2960 (N_2960,N_741,N_1505);
and U2961 (N_2961,N_879,N_764);
nor U2962 (N_2962,N_491,N_1494);
or U2963 (N_2963,N_1860,N_747);
or U2964 (N_2964,N_276,N_2149);
xnor U2965 (N_2965,N_1217,N_1683);
nand U2966 (N_2966,N_234,N_1448);
or U2967 (N_2967,N_121,N_2485);
nor U2968 (N_2968,N_1547,N_965);
xnor U2969 (N_2969,N_1968,N_797);
nand U2970 (N_2970,N_199,N_280);
nor U2971 (N_2971,N_1548,N_925);
xnor U2972 (N_2972,N_2243,N_1582);
or U2973 (N_2973,N_548,N_1603);
or U2974 (N_2974,N_2105,N_1899);
or U2975 (N_2975,N_75,N_1006);
xnor U2976 (N_2976,N_560,N_2376);
and U2977 (N_2977,N_1798,N_2013);
xor U2978 (N_2978,N_1672,N_730);
nor U2979 (N_2979,N_440,N_1744);
nor U2980 (N_2980,N_2468,N_1194);
xor U2981 (N_2981,N_1461,N_409);
or U2982 (N_2982,N_2257,N_148);
xnor U2983 (N_2983,N_839,N_405);
and U2984 (N_2984,N_97,N_1530);
nor U2985 (N_2985,N_1293,N_460);
and U2986 (N_2986,N_1533,N_1343);
or U2987 (N_2987,N_1896,N_1720);
and U2988 (N_2988,N_90,N_1271);
xor U2989 (N_2989,N_927,N_597);
and U2990 (N_2990,N_532,N_823);
or U2991 (N_2991,N_1874,N_330);
xnor U2992 (N_2992,N_67,N_1554);
or U2993 (N_2993,N_558,N_1492);
nand U2994 (N_2994,N_1602,N_977);
xor U2995 (N_2995,N_751,N_76);
nand U2996 (N_2996,N_82,N_1323);
xnor U2997 (N_2997,N_2017,N_1673);
or U2998 (N_2998,N_371,N_451);
or U2999 (N_2999,N_2245,N_1397);
and U3000 (N_3000,N_924,N_1088);
xor U3001 (N_3001,N_313,N_1080);
or U3002 (N_3002,N_296,N_467);
nor U3003 (N_3003,N_761,N_2189);
nor U3004 (N_3004,N_1344,N_1172);
and U3005 (N_3005,N_2053,N_1713);
and U3006 (N_3006,N_612,N_2179);
xor U3007 (N_3007,N_1210,N_2431);
nor U3008 (N_3008,N_403,N_689);
nand U3009 (N_3009,N_1910,N_387);
nor U3010 (N_3010,N_2111,N_1365);
xnor U3011 (N_3011,N_1440,N_975);
and U3012 (N_3012,N_1462,N_1828);
nand U3013 (N_3013,N_1942,N_1214);
and U3014 (N_3014,N_1300,N_711);
and U3015 (N_3015,N_1792,N_1186);
nor U3016 (N_3016,N_2322,N_867);
nand U3017 (N_3017,N_2418,N_58);
nor U3018 (N_3018,N_1449,N_1268);
nand U3019 (N_3019,N_1259,N_1879);
xor U3020 (N_3020,N_2219,N_73);
or U3021 (N_3021,N_1677,N_708);
nor U3022 (N_3022,N_1509,N_881);
or U3023 (N_3023,N_1295,N_2248);
and U3024 (N_3024,N_2221,N_1410);
or U3025 (N_3025,N_909,N_2208);
xor U3026 (N_3026,N_599,N_1436);
or U3027 (N_3027,N_1067,N_1341);
or U3028 (N_3028,N_217,N_2292);
or U3029 (N_3029,N_1352,N_1752);
xor U3030 (N_3030,N_256,N_787);
nand U3031 (N_3031,N_2130,N_802);
xnor U3032 (N_3032,N_1111,N_2309);
and U3033 (N_3033,N_230,N_150);
xnor U3034 (N_3034,N_2416,N_141);
xnor U3035 (N_3035,N_1531,N_1862);
or U3036 (N_3036,N_2146,N_383);
and U3037 (N_3037,N_586,N_142);
xor U3038 (N_3038,N_108,N_2140);
or U3039 (N_3039,N_934,N_806);
nand U3040 (N_3040,N_1555,N_1684);
nand U3041 (N_3041,N_1359,N_817);
or U3042 (N_3042,N_1447,N_1338);
nand U3043 (N_3043,N_133,N_2422);
or U3044 (N_3044,N_1948,N_300);
nand U3045 (N_3045,N_1722,N_754);
xnor U3046 (N_3046,N_1075,N_1469);
nand U3047 (N_3047,N_1227,N_2290);
xnor U3048 (N_3048,N_1296,N_272);
nor U3049 (N_3049,N_2128,N_1679);
nor U3050 (N_3050,N_2346,N_2190);
and U3051 (N_3051,N_2369,N_1778);
xnor U3052 (N_3052,N_908,N_1791);
and U3053 (N_3053,N_1465,N_1546);
nand U3054 (N_3054,N_2378,N_350);
nor U3055 (N_3055,N_543,N_1551);
xor U3056 (N_3056,N_429,N_2056);
and U3057 (N_3057,N_1189,N_624);
nand U3058 (N_3058,N_1280,N_265);
nand U3059 (N_3059,N_2085,N_2333);
nor U3060 (N_3060,N_2447,N_20);
and U3061 (N_3061,N_2100,N_1089);
or U3062 (N_3062,N_628,N_827);
nor U3063 (N_3063,N_939,N_899);
nand U3064 (N_3064,N_1576,N_600);
nand U3065 (N_3065,N_800,N_1200);
and U3066 (N_3066,N_2185,N_951);
or U3067 (N_3067,N_2282,N_2470);
or U3068 (N_3068,N_2476,N_1371);
and U3069 (N_3069,N_1102,N_721);
nand U3070 (N_3070,N_520,N_1286);
xnor U3071 (N_3071,N_1636,N_282);
nand U3072 (N_3072,N_32,N_1055);
or U3073 (N_3073,N_2016,N_1951);
nor U3074 (N_3074,N_285,N_1779);
or U3075 (N_3075,N_1751,N_2366);
nand U3076 (N_3076,N_92,N_2317);
nand U3077 (N_3077,N_2455,N_2049);
xnor U3078 (N_3078,N_691,N_461);
nor U3079 (N_3079,N_393,N_1694);
nor U3080 (N_3080,N_952,N_1159);
nand U3081 (N_3081,N_1863,N_2068);
xor U3082 (N_3082,N_1512,N_511);
nor U3083 (N_3083,N_513,N_1640);
xor U3084 (N_3084,N_1451,N_716);
xor U3085 (N_3085,N_1644,N_2199);
and U3086 (N_3086,N_480,N_980);
nor U3087 (N_3087,N_1078,N_38);
or U3088 (N_3088,N_2098,N_1772);
nand U3089 (N_3089,N_2177,N_1285);
nand U3090 (N_3090,N_1692,N_253);
nand U3091 (N_3091,N_528,N_845);
nand U3092 (N_3092,N_117,N_2286);
or U3093 (N_3093,N_1182,N_2359);
and U3094 (N_3094,N_343,N_54);
nor U3095 (N_3095,N_2277,N_3);
and U3096 (N_3096,N_218,N_1083);
and U3097 (N_3097,N_1753,N_561);
xor U3098 (N_3098,N_53,N_1430);
or U3099 (N_3099,N_737,N_1587);
nor U3100 (N_3100,N_2278,N_438);
and U3101 (N_3101,N_640,N_2340);
nor U3102 (N_3102,N_40,N_910);
or U3103 (N_3103,N_706,N_151);
or U3104 (N_3104,N_2203,N_962);
xnor U3105 (N_3105,N_1125,N_498);
xnor U3106 (N_3106,N_2144,N_1729);
nor U3107 (N_3107,N_1336,N_1458);
nand U3108 (N_3108,N_425,N_2428);
nor U3109 (N_3109,N_699,N_857);
nor U3110 (N_3110,N_10,N_644);
nor U3111 (N_3111,N_2059,N_1192);
nor U3112 (N_3112,N_80,N_717);
or U3113 (N_3113,N_801,N_2372);
nor U3114 (N_3114,N_229,N_2152);
nand U3115 (N_3115,N_794,N_674);
nand U3116 (N_3116,N_2367,N_1937);
nor U3117 (N_3117,N_170,N_991);
and U3118 (N_3118,N_2154,N_333);
or U3119 (N_3119,N_2173,N_1818);
and U3120 (N_3120,N_2184,N_621);
nor U3121 (N_3121,N_1195,N_1647);
nand U3122 (N_3122,N_992,N_1048);
and U3123 (N_3123,N_2158,N_2132);
nand U3124 (N_3124,N_579,N_59);
xor U3125 (N_3125,N_1878,N_1072);
nor U3126 (N_3126,N_1022,N_1257);
nand U3127 (N_3127,N_65,N_2313);
and U3128 (N_3128,N_1007,N_70);
nor U3129 (N_3129,N_1566,N_667);
nor U3130 (N_3130,N_1082,N_2066);
nand U3131 (N_3131,N_1407,N_186);
or U3132 (N_3132,N_505,N_1156);
nand U3133 (N_3133,N_1966,N_2487);
and U3134 (N_3134,N_2412,N_433);
nand U3135 (N_3135,N_2389,N_1946);
nor U3136 (N_3136,N_2347,N_1165);
and U3137 (N_3137,N_1450,N_2151);
nand U3138 (N_3138,N_936,N_611);
nand U3139 (N_3139,N_1803,N_1906);
nor U3140 (N_3140,N_1617,N_1417);
xnor U3141 (N_3141,N_1140,N_1765);
and U3142 (N_3142,N_1098,N_2148);
or U3143 (N_3143,N_844,N_12);
nor U3144 (N_3144,N_837,N_1301);
nand U3145 (N_3145,N_435,N_1116);
and U3146 (N_3146,N_738,N_474);
and U3147 (N_3147,N_252,N_1281);
nor U3148 (N_3148,N_188,N_344);
nand U3149 (N_3149,N_499,N_1624);
or U3150 (N_3150,N_1477,N_1277);
nor U3151 (N_3151,N_1933,N_2025);
nand U3152 (N_3152,N_1882,N_501);
nor U3153 (N_3153,N_466,N_608);
and U3154 (N_3154,N_847,N_1033);
xnor U3155 (N_3155,N_2113,N_1361);
and U3156 (N_3156,N_569,N_666);
nand U3157 (N_3157,N_2403,N_1515);
nor U3158 (N_3158,N_1913,N_1190);
xnor U3159 (N_3159,N_1275,N_2305);
or U3160 (N_3160,N_1070,N_103);
nor U3161 (N_3161,N_483,N_1482);
xnor U3162 (N_3162,N_775,N_1236);
xor U3163 (N_3163,N_1028,N_1927);
xor U3164 (N_3164,N_1467,N_1543);
nand U3165 (N_3165,N_1870,N_2205);
and U3166 (N_3166,N_44,N_261);
and U3167 (N_3167,N_753,N_1255);
nor U3168 (N_3168,N_359,N_1201);
nand U3169 (N_3169,N_1353,N_916);
nor U3170 (N_3170,N_710,N_826);
nand U3171 (N_3171,N_1529,N_661);
and U3172 (N_3172,N_2280,N_2494);
xor U3173 (N_3173,N_1139,N_1501);
xnor U3174 (N_3174,N_1131,N_250);
nand U3175 (N_3175,N_1702,N_2300);
nand U3176 (N_3176,N_365,N_1216);
and U3177 (N_3177,N_1747,N_1087);
or U3178 (N_3178,N_1322,N_328);
nand U3179 (N_3179,N_1608,N_107);
xor U3180 (N_3180,N_1325,N_2404);
and U3181 (N_3181,N_1218,N_1708);
nor U3182 (N_3182,N_1613,N_1689);
or U3183 (N_3183,N_74,N_1975);
and U3184 (N_3184,N_610,N_1000);
xor U3185 (N_3185,N_1157,N_2045);
and U3186 (N_3186,N_688,N_41);
and U3187 (N_3187,N_1934,N_1898);
nand U3188 (N_3188,N_174,N_266);
xor U3189 (N_3189,N_64,N_369);
nor U3190 (N_3190,N_2377,N_607);
or U3191 (N_3191,N_1688,N_1339);
nand U3192 (N_3192,N_2355,N_2279);
or U3193 (N_3193,N_2071,N_1923);
or U3194 (N_3194,N_953,N_1122);
or U3195 (N_3195,N_1565,N_2232);
nand U3196 (N_3196,N_1912,N_2039);
nor U3197 (N_3197,N_2092,N_1278);
nor U3198 (N_3198,N_1589,N_1560);
and U3199 (N_3199,N_1742,N_323);
and U3200 (N_3200,N_1424,N_1289);
and U3201 (N_3201,N_1764,N_1527);
nor U3202 (N_3202,N_2357,N_1027);
or U3203 (N_3203,N_72,N_1979);
nand U3204 (N_3204,N_1885,N_398);
nor U3205 (N_3205,N_567,N_1897);
and U3206 (N_3206,N_81,N_329);
xor U3207 (N_3207,N_805,N_1488);
nor U3208 (N_3208,N_91,N_413);
nor U3209 (N_3209,N_2475,N_1775);
nor U3210 (N_3210,N_1796,N_855);
nor U3211 (N_3211,N_446,N_1003);
xor U3212 (N_3212,N_224,N_1348);
or U3213 (N_3213,N_1808,N_1628);
xor U3214 (N_3214,N_1009,N_1888);
nand U3215 (N_3215,N_2345,N_2095);
or U3216 (N_3216,N_2331,N_946);
nand U3217 (N_3217,N_351,N_1964);
nand U3218 (N_3218,N_2307,N_2312);
or U3219 (N_3219,N_790,N_232);
or U3220 (N_3220,N_2218,N_84);
xor U3221 (N_3221,N_2259,N_283);
nor U3222 (N_3222,N_209,N_1865);
nor U3223 (N_3223,N_1721,N_647);
and U3224 (N_3224,N_183,N_1754);
and U3225 (N_3225,N_463,N_1929);
nand U3226 (N_3226,N_31,N_2471);
or U3227 (N_3227,N_1908,N_1261);
nand U3228 (N_3228,N_281,N_52);
xnor U3229 (N_3229,N_299,N_1079);
nand U3230 (N_3230,N_2125,N_749);
xor U3231 (N_3231,N_522,N_1866);
and U3232 (N_3232,N_713,N_744);
or U3233 (N_3233,N_876,N_1209);
xnor U3234 (N_3234,N_1738,N_1081);
and U3235 (N_3235,N_2217,N_1768);
or U3236 (N_3236,N_1128,N_293);
nor U3237 (N_3237,N_423,N_1386);
xnor U3238 (N_3238,N_1563,N_2435);
and U3239 (N_3239,N_1086,N_1126);
or U3240 (N_3240,N_2269,N_773);
nand U3241 (N_3241,N_776,N_496);
and U3242 (N_3242,N_1656,N_454);
nand U3243 (N_3243,N_1015,N_777);
or U3244 (N_3244,N_605,N_634);
xnor U3245 (N_3245,N_2227,N_424);
xnor U3246 (N_3246,N_1605,N_2353);
and U3247 (N_3247,N_1019,N_1550);
nor U3248 (N_3248,N_606,N_1486);
nor U3249 (N_3249,N_1112,N_2175);
nor U3250 (N_3250,N_1060,N_372);
nor U3251 (N_3251,N_1208,N_1024);
xnor U3252 (N_3252,N_2320,N_140);
or U3253 (N_3253,N_2202,N_2482);
nor U3254 (N_3254,N_2351,N_665);
nand U3255 (N_3255,N_1394,N_956);
xnor U3256 (N_3256,N_158,N_1663);
or U3257 (N_3257,N_921,N_1026);
nand U3258 (N_3258,N_609,N_1110);
nand U3259 (N_3259,N_2026,N_494);
nor U3260 (N_3260,N_1599,N_1944);
and U3261 (N_3261,N_2254,N_397);
xor U3262 (N_3262,N_1053,N_1700);
nor U3263 (N_3263,N_420,N_273);
nand U3264 (N_3264,N_2097,N_679);
nor U3265 (N_3265,N_1705,N_574);
and U3266 (N_3266,N_1847,N_2440);
and U3267 (N_3267,N_2379,N_1731);
or U3268 (N_3268,N_1506,N_2271);
xor U3269 (N_3269,N_89,N_2273);
and U3270 (N_3270,N_25,N_2464);
nand U3271 (N_3271,N_376,N_1016);
nor U3272 (N_3272,N_1740,N_1229);
or U3273 (N_3273,N_1697,N_592);
xnor U3274 (N_3274,N_830,N_1653);
and U3275 (N_3275,N_146,N_2399);
or U3276 (N_3276,N_51,N_2308);
or U3277 (N_3277,N_402,N_404);
or U3278 (N_3278,N_1685,N_670);
nor U3279 (N_3279,N_254,N_1057);
xnor U3280 (N_3280,N_1532,N_735);
nand U3281 (N_3281,N_1108,N_1930);
or U3282 (N_3282,N_858,N_821);
nand U3283 (N_3283,N_1106,N_1233);
and U3284 (N_3284,N_643,N_263);
nand U3285 (N_3285,N_1585,N_68);
or U3286 (N_3286,N_1457,N_302);
nand U3287 (N_3287,N_1310,N_859);
nor U3288 (N_3288,N_482,N_2425);
nor U3289 (N_3289,N_1972,N_1511);
xor U3290 (N_3290,N_124,N_1832);
nor U3291 (N_3291,N_368,N_901);
or U3292 (N_3292,N_1426,N_1030);
xnor U3293 (N_3293,N_1986,N_1327);
nor U3294 (N_3294,N_274,N_1490);
or U3295 (N_3295,N_1318,N_1312);
nor U3296 (N_3296,N_807,N_1062);
or U3297 (N_3297,N_1103,N_1812);
and U3298 (N_3298,N_1635,N_1620);
or U3299 (N_3299,N_1881,N_1639);
and U3300 (N_3300,N_2075,N_2084);
xnor U3301 (N_3301,N_1997,N_416);
nor U3302 (N_3302,N_1153,N_1084);
xnor U3303 (N_3303,N_1138,N_822);
or U3304 (N_3304,N_1315,N_1851);
nor U3305 (N_3305,N_1580,N_2153);
nand U3306 (N_3306,N_1520,N_877);
nand U3307 (N_3307,N_1267,N_685);
nor U3308 (N_3308,N_457,N_2002);
nand U3309 (N_3309,N_1723,N_2106);
and U3310 (N_3310,N_1429,N_2138);
nor U3311 (N_3311,N_1416,N_742);
nor U3312 (N_3312,N_1375,N_2041);
xnor U3313 (N_3313,N_471,N_309);
or U3314 (N_3314,N_497,N_785);
or U3315 (N_3315,N_923,N_1251);
xor U3316 (N_3316,N_637,N_112);
and U3317 (N_3317,N_1843,N_2222);
xor U3318 (N_3318,N_871,N_2198);
and U3319 (N_3319,N_123,N_2086);
xnor U3320 (N_3320,N_2298,N_2373);
nor U3321 (N_3321,N_1135,N_161);
or U3322 (N_3322,N_1076,N_2186);
nor U3323 (N_3323,N_2210,N_182);
nor U3324 (N_3324,N_2135,N_410);
nor U3325 (N_3325,N_1404,N_896);
xnor U3326 (N_3326,N_1205,N_623);
nand U3327 (N_3327,N_481,N_1354);
nor U3328 (N_3328,N_990,N_35);
or U3329 (N_3329,N_1291,N_1035);
or U3330 (N_3330,N_212,N_171);
xor U3331 (N_3331,N_2492,N_1017);
nor U3332 (N_3332,N_1091,N_1726);
nand U3333 (N_3333,N_2164,N_1797);
nand U3334 (N_3334,N_1425,N_1645);
or U3335 (N_3335,N_914,N_795);
nand U3336 (N_3336,N_17,N_1238);
nand U3337 (N_3337,N_1304,N_1641);
and U3338 (N_3338,N_2087,N_1873);
or U3339 (N_3339,N_1212,N_2356);
and U3340 (N_3340,N_1121,N_941);
and U3341 (N_3341,N_549,N_1850);
nor U3342 (N_3342,N_1152,N_2220);
xnor U3343 (N_3343,N_1633,N_2466);
nand U3344 (N_3344,N_2057,N_1069);
and U3345 (N_3345,N_389,N_651);
xor U3346 (N_3346,N_734,N_1559);
nor U3347 (N_3347,N_33,N_1314);
xnor U3348 (N_3348,N_509,N_437);
xor U3349 (N_3349,N_1701,N_134);
or U3350 (N_3350,N_2165,N_1160);
and U3351 (N_3351,N_1999,N_1976);
or U3352 (N_3352,N_175,N_1955);
nand U3353 (N_3353,N_1606,N_1893);
nand U3354 (N_3354,N_1441,N_1601);
or U3355 (N_3355,N_2408,N_2170);
nor U3356 (N_3356,N_2124,N_722);
nand U3357 (N_3357,N_935,N_1827);
nor U3358 (N_3358,N_1119,N_2314);
nand U3359 (N_3359,N_311,N_1704);
nor U3360 (N_3360,N_152,N_2195);
or U3361 (N_3361,N_1667,N_1032);
nand U3362 (N_3362,N_862,N_792);
or U3363 (N_3363,N_1669,N_1105);
and U3364 (N_3364,N_1380,N_1115);
nand U3365 (N_3365,N_1610,N_353);
nor U3366 (N_3366,N_1432,N_325);
or U3367 (N_3367,N_1423,N_1499);
nand U3368 (N_3368,N_2030,N_297);
xor U3369 (N_3369,N_364,N_2159);
or U3370 (N_3370,N_1849,N_1308);
nor U3371 (N_3371,N_241,N_1162);
nor U3372 (N_3372,N_680,N_2080);
nor U3373 (N_3373,N_2021,N_2136);
nand U3374 (N_3374,N_659,N_1928);
and U3375 (N_3375,N_1002,N_1816);
or U3376 (N_3376,N_668,N_184);
xnor U3377 (N_3377,N_2024,N_598);
or U3378 (N_3378,N_2465,N_973);
and U3379 (N_3379,N_820,N_2261);
nand U3380 (N_3380,N_894,N_1790);
xnor U3381 (N_3381,N_484,N_1427);
nor U3382 (N_3382,N_1346,N_1253);
and U3383 (N_3383,N_1406,N_918);
nor U3384 (N_3384,N_2214,N_866);
or U3385 (N_3385,N_1698,N_958);
xnor U3386 (N_3386,N_1369,N_422);
and U3387 (N_3387,N_1114,N_886);
nand U3388 (N_3388,N_1973,N_255);
or U3389 (N_3389,N_2032,N_1595);
and U3390 (N_3390,N_604,N_358);
and U3391 (N_3391,N_693,N_2258);
nor U3392 (N_3392,N_966,N_704);
or U3393 (N_3393,N_907,N_2225);
xor U3394 (N_3394,N_1328,N_1611);
and U3395 (N_3395,N_559,N_1307);
nand U3396 (N_3396,N_326,N_2410);
xor U3397 (N_3397,N_1297,N_1516);
nor U3398 (N_3398,N_1510,N_317);
nor U3399 (N_3399,N_176,N_652);
and U3400 (N_3400,N_168,N_275);
nand U3401 (N_3401,N_2076,N_1366);
nand U3402 (N_3402,N_15,N_355);
and U3403 (N_3403,N_812,N_1113);
xnor U3404 (N_3404,N_993,N_370);
xnor U3405 (N_3405,N_2456,N_2226);
nor U3406 (N_3406,N_736,N_1203);
xnor U3407 (N_3407,N_2302,N_1575);
and U3408 (N_3408,N_86,N_401);
xor U3409 (N_3409,N_129,N_2231);
and U3410 (N_3410,N_166,N_2499);
nand U3411 (N_3411,N_1294,N_584);
nand U3412 (N_3412,N_489,N_415);
nand U3413 (N_3413,N_156,N_1270);
nand U3414 (N_3414,N_950,N_2103);
and U3415 (N_3415,N_1596,N_1155);
and U3416 (N_3416,N_638,N_449);
nor U3417 (N_3417,N_2364,N_2091);
nand U3418 (N_3418,N_878,N_1148);
xor U3419 (N_3419,N_1538,N_2155);
and U3420 (N_3420,N_2430,N_593);
and U3421 (N_3421,N_2339,N_29);
nor U3422 (N_3422,N_2394,N_529);
nor U3423 (N_3423,N_552,N_1400);
nand U3424 (N_3424,N_318,N_46);
nand U3425 (N_3425,N_1330,N_664);
nor U3426 (N_3426,N_2423,N_1670);
or U3427 (N_3427,N_1066,N_1544);
nor U3428 (N_3428,N_2341,N_626);
and U3429 (N_3429,N_1384,N_2060);
or U3430 (N_3430,N_2005,N_694);
nand U3431 (N_3431,N_1572,N_1745);
or U3432 (N_3432,N_2424,N_287);
xor U3433 (N_3433,N_1239,N_160);
nor U3434 (N_3434,N_2329,N_1631);
nand U3435 (N_3435,N_13,N_2090);
nor U3436 (N_3436,N_2400,N_1707);
nand U3437 (N_3437,N_919,N_920);
nor U3438 (N_3438,N_428,N_905);
or U3439 (N_3439,N_898,N_1841);
nand U3440 (N_3440,N_1254,N_1638);
nor U3441 (N_3441,N_1936,N_1623);
and U3442 (N_3442,N_163,N_960);
nand U3443 (N_3443,N_1686,N_1039);
xor U3444 (N_3444,N_2392,N_2285);
nand U3445 (N_3445,N_2459,N_1773);
and U3446 (N_3446,N_1789,N_1859);
nor U3447 (N_3447,N_1938,N_1802);
or U3448 (N_3448,N_591,N_332);
nand U3449 (N_3449,N_1872,N_1421);
or U3450 (N_3450,N_602,N_2004);
or U3451 (N_3451,N_620,N_874);
nor U3452 (N_3452,N_227,N_1821);
and U3453 (N_3453,N_1470,N_2050);
xor U3454 (N_3454,N_1904,N_220);
and U3455 (N_3455,N_235,N_2281);
xnor U3456 (N_3456,N_453,N_1132);
nor U3457 (N_3457,N_1163,N_677);
or U3458 (N_3458,N_1129,N_407);
nand U3459 (N_3459,N_443,N_2061);
and U3460 (N_3460,N_200,N_2496);
nand U3461 (N_3461,N_2446,N_2197);
nor U3462 (N_3462,N_247,N_1240);
xnor U3463 (N_3463,N_725,N_1097);
nor U3464 (N_3464,N_582,N_2477);
nand U3465 (N_3465,N_2272,N_1460);
xor U3466 (N_3466,N_2200,N_1793);
nor U3467 (N_3467,N_819,N_1680);
xnor U3468 (N_3468,N_1389,N_639);
nand U3469 (N_3469,N_1815,N_697);
or U3470 (N_3470,N_379,N_63);
nor U3471 (N_3471,N_421,N_2062);
or U3472 (N_3472,N_1604,N_2330);
xor U3473 (N_3473,N_2409,N_2365);
xnor U3474 (N_3474,N_207,N_2407);
and U3475 (N_3475,N_1452,N_2328);
nand U3476 (N_3476,N_1901,N_1757);
or U3477 (N_3477,N_1347,N_34);
nand U3478 (N_3478,N_2417,N_1287);
nor U3479 (N_3479,N_733,N_1989);
nand U3480 (N_3480,N_245,N_2391);
xnor U3481 (N_3481,N_1193,N_1632);
nand U3482 (N_3482,N_1761,N_1250);
nor U3483 (N_3483,N_1943,N_1197);
nand U3484 (N_3484,N_298,N_1120);
and U3485 (N_3485,N_495,N_2395);
and U3486 (N_3486,N_439,N_1950);
and U3487 (N_3487,N_1316,N_18);
and U3488 (N_3488,N_105,N_2169);
nor U3489 (N_3489,N_464,N_462);
xnor U3490 (N_3490,N_926,N_2433);
or U3491 (N_3491,N_1891,N_2114);
nand U3492 (N_3492,N_576,N_2401);
or U3493 (N_3493,N_1970,N_1814);
nand U3494 (N_3494,N_1718,N_1232);
nand U3495 (N_3495,N_1133,N_1907);
or U3496 (N_3496,N_1562,N_1556);
and U3497 (N_3497,N_999,N_1715);
nand U3498 (N_3498,N_1958,N_165);
xor U3499 (N_3499,N_1581,N_1993);
and U3500 (N_3500,N_517,N_1774);
xnor U3501 (N_3501,N_1101,N_853);
or U3502 (N_3502,N_418,N_1405);
xnor U3503 (N_3503,N_1276,N_573);
nand U3504 (N_3504,N_459,N_2382);
or U3505 (N_3505,N_848,N_2405);
nand U3506 (N_3506,N_2116,N_968);
or U3507 (N_3507,N_292,N_869);
and U3508 (N_3508,N_615,N_2318);
nand U3509 (N_3509,N_2006,N_873);
nor U3510 (N_3510,N_2234,N_1526);
nand U3511 (N_3511,N_1962,N_686);
xnor U3512 (N_3512,N_1769,N_585);
xor U3513 (N_3513,N_516,N_257);
nand U3514 (N_3514,N_728,N_1534);
nand U3515 (N_3515,N_1402,N_1442);
or U3516 (N_3516,N_1433,N_233);
or U3517 (N_3517,N_2027,N_889);
and U3518 (N_3518,N_1853,N_2311);
or U3519 (N_3519,N_1969,N_1691);
xnor U3520 (N_3520,N_2126,N_856);
nand U3521 (N_3521,N_1224,N_2110);
nor U3522 (N_3522,N_2001,N_98);
and U3523 (N_3523,N_334,N_259);
nand U3524 (N_3524,N_2191,N_1877);
or U3525 (N_3525,N_427,N_2178);
nor U3526 (N_3526,N_288,N_1995);
nor U3527 (N_3527,N_1403,N_743);
and U3528 (N_3528,N_2115,N_2360);
or U3529 (N_3529,N_1317,N_104);
nand U3530 (N_3530,N_1211,N_1204);
or U3531 (N_3531,N_1835,N_1202);
xor U3532 (N_3532,N_1058,N_1925);
nand U3533 (N_3533,N_225,N_1244);
nor U3534 (N_3534,N_1561,N_2415);
nor U3535 (N_3535,N_1574,N_762);
and U3536 (N_3536,N_2323,N_2252);
nor U3537 (N_3537,N_1104,N_1622);
xor U3538 (N_3538,N_731,N_347);
or U3539 (N_3539,N_1921,N_675);
nor U3540 (N_3540,N_1279,N_2419);
xnor U3541 (N_3541,N_1932,N_726);
and U3542 (N_3542,N_2397,N_963);
nor U3543 (N_3543,N_981,N_782);
nor U3544 (N_3544,N_191,N_998);
nand U3545 (N_3545,N_2121,N_2484);
or U3546 (N_3546,N_286,N_1954);
nor U3547 (N_3547,N_1809,N_226);
xnor U3548 (N_3548,N_707,N_1586);
xor U3549 (N_3549,N_1846,N_1991);
nand U3550 (N_3550,N_2196,N_336);
xnor U3551 (N_3551,N_835,N_238);
or U3552 (N_3552,N_2023,N_1391);
xnor U3553 (N_3553,N_829,N_2390);
xnor U3554 (N_3554,N_1514,N_1894);
nand U3555 (N_3555,N_2352,N_1952);
and U3556 (N_3556,N_1657,N_60);
nand U3557 (N_3557,N_375,N_1179);
nor U3558 (N_3558,N_1077,N_2321);
xor U3559 (N_3559,N_2263,N_1263);
and U3560 (N_3560,N_1408,N_477);
nor U3561 (N_3561,N_2112,N_2089);
or U3562 (N_3562,N_2166,N_2325);
nand U3563 (N_3563,N_955,N_1988);
and U3564 (N_3564,N_996,N_1331);
nor U3565 (N_3565,N_583,N_2275);
xnor U3566 (N_3566,N_2452,N_831);
xnor U3567 (N_3567,N_540,N_813);
xnor U3568 (N_3568,N_1199,N_1356);
nand U3569 (N_3569,N_1642,N_1687);
nand U3570 (N_3570,N_1848,N_2183);
and U3571 (N_3571,N_1918,N_2439);
nand U3572 (N_3572,N_1124,N_469);
nand U3573 (N_3573,N_663,N_1481);
or U3574 (N_3574,N_1643,N_1064);
nor U3575 (N_3575,N_933,N_882);
or U3576 (N_3576,N_985,N_783);
nor U3577 (N_3577,N_1727,N_997);
nand U3578 (N_3578,N_2442,N_120);
nor U3579 (N_3579,N_769,N_650);
xnor U3580 (N_3580,N_508,N_119);
nand U3581 (N_3581,N_1258,N_1150);
nor U3582 (N_3582,N_327,N_627);
nor U3583 (N_3583,N_565,N_1147);
xor U3584 (N_3584,N_772,N_1771);
nand U3585 (N_3585,N_380,N_1739);
nor U3586 (N_3586,N_632,N_458);
xor U3587 (N_3587,N_545,N_1377);
nor U3588 (N_3588,N_868,N_564);
and U3589 (N_3589,N_954,N_1535);
xnor U3590 (N_3590,N_1381,N_2295);
and U3591 (N_3591,N_1630,N_1363);
or U3592 (N_3592,N_2438,N_1164);
or U3593 (N_3593,N_1094,N_1050);
nor U3594 (N_3594,N_1998,N_1456);
or U3595 (N_3595,N_1883,N_452);
or U3596 (N_3596,N_2358,N_631);
and U3597 (N_3597,N_947,N_1621);
nand U3598 (N_3598,N_2421,N_1178);
nand U3599 (N_3599,N_1011,N_1029);
or U3600 (N_3600,N_2411,N_1905);
or U3601 (N_3601,N_1351,N_838);
xnor U3602 (N_3602,N_1303,N_419);
and U3603 (N_3603,N_682,N_2413);
xnor U3604 (N_3604,N_310,N_1583);
or U3605 (N_3605,N_189,N_642);
nand U3606 (N_3606,N_2388,N_1822);
xor U3607 (N_3607,N_2469,N_219);
xnor U3608 (N_3608,N_959,N_488);
and U3609 (N_3609,N_1176,N_1497);
and U3610 (N_3610,N_1142,N_863);
nand U3611 (N_3611,N_1489,N_551);
xor U3612 (N_3612,N_614,N_1439);
nand U3613 (N_3613,N_2274,N_1043);
nand U3614 (N_3614,N_850,N_1917);
nand U3615 (N_3615,N_2398,N_1374);
xor U3616 (N_3616,N_987,N_2194);
nor U3617 (N_3617,N_1788,N_2461);
xor U3618 (N_3618,N_1466,N_2486);
nor U3619 (N_3619,N_2240,N_2029);
xnor U3620 (N_3620,N_590,N_335);
and U3621 (N_3621,N_1579,N_1994);
nor U3622 (N_3622,N_836,N_1483);
and U3623 (N_3623,N_1283,N_1755);
or U3624 (N_3624,N_1207,N_2011);
and U3625 (N_3625,N_1237,N_1390);
nor U3626 (N_3626,N_486,N_1748);
nand U3627 (N_3627,N_630,N_1733);
and U3628 (N_3628,N_1690,N_1759);
nor U3629 (N_3629,N_788,N_1046);
nor U3630 (N_3630,N_1018,N_179);
nor U3631 (N_3631,N_1382,N_303);
nor U3632 (N_3632,N_1379,N_1650);
nor U3633 (N_3633,N_2109,N_1388);
nand U3634 (N_3634,N_1868,N_1023);
xnor U3635 (N_3635,N_989,N_1428);
or U3636 (N_3636,N_1990,N_1578);
and U3637 (N_3637,N_1889,N_1266);
and U3638 (N_3638,N_897,N_2483);
xnor U3639 (N_3639,N_1736,N_1184);
or U3640 (N_3640,N_162,N_1265);
nor U3641 (N_3641,N_1471,N_1437);
and U3642 (N_3642,N_24,N_2096);
nand U3643 (N_3643,N_1444,N_1177);
xor U3644 (N_3644,N_988,N_1668);
nor U3645 (N_3645,N_671,N_1231);
and U3646 (N_3646,N_77,N_1420);
nor U3647 (N_3647,N_538,N_976);
or U3648 (N_3648,N_1171,N_2108);
xor U3649 (N_3649,N_629,N_88);
nand U3650 (N_3650,N_1333,N_2233);
nor U3651 (N_3651,N_308,N_875);
or U3652 (N_3652,N_2127,N_206);
nor U3653 (N_3653,N_2142,N_1706);
nand U3654 (N_3654,N_2216,N_2054);
nor U3655 (N_3655,N_504,N_994);
xor U3656 (N_3656,N_1223,N_2303);
or U3657 (N_3657,N_2497,N_1385);
and U3658 (N_3658,N_441,N_1646);
nor U3659 (N_3659,N_1144,N_472);
and U3660 (N_3660,N_2022,N_185);
nor U3661 (N_3661,N_892,N_911);
nor U3662 (N_3662,N_571,N_2213);
nand U3663 (N_3663,N_1806,N_2187);
nand U3664 (N_3664,N_1967,N_1364);
nor U3665 (N_3665,N_1985,N_1838);
xnor U3666 (N_3666,N_1298,N_1376);
or U3667 (N_3667,N_69,N_809);
and U3668 (N_3668,N_1464,N_215);
and U3669 (N_3669,N_1799,N_167);
and U3670 (N_3670,N_1664,N_2055);
nor U3671 (N_3671,N_1782,N_957);
xor U3672 (N_3672,N_536,N_1463);
and U3673 (N_3673,N_752,N_2000);
nor U3674 (N_3674,N_2326,N_893);
xnor U3675 (N_3675,N_967,N_1758);
xnor U3676 (N_3676,N_2338,N_1654);
and U3677 (N_3677,N_21,N_352);
nand U3678 (N_3678,N_216,N_646);
xor U3679 (N_3679,N_1518,N_2141);
xor U3680 (N_3680,N_2462,N_1626);
xor U3681 (N_3681,N_1709,N_1136);
nand U3682 (N_3682,N_390,N_173);
nand U3683 (N_3683,N_1358,N_2283);
xnor U3684 (N_3684,N_709,N_1309);
nand U3685 (N_3685,N_66,N_603);
nand U3686 (N_3686,N_2332,N_815);
or U3687 (N_3687,N_130,N_1537);
and U3688 (N_3688,N_96,N_143);
and U3689 (N_3689,N_1010,N_14);
xor U3690 (N_3690,N_2460,N_243);
xnor U3691 (N_3691,N_1052,N_392);
xor U3692 (N_3692,N_2451,N_587);
nand U3693 (N_3693,N_1909,N_118);
or U3694 (N_3694,N_622,N_1290);
xor U3695 (N_3695,N_633,N_1235);
nand U3696 (N_3696,N_228,N_1161);
or U3697 (N_3697,N_1074,N_922);
nor U3698 (N_3698,N_1187,N_2052);
nand U3699 (N_3699,N_687,N_242);
or U3700 (N_3700,N_912,N_2133);
xnor U3701 (N_3701,N_1716,N_2180);
nor U3702 (N_3702,N_2260,N_1134);
nand U3703 (N_3703,N_270,N_1800);
or U3704 (N_3704,N_2361,N_1784);
or U3705 (N_3705,N_2162,N_236);
nand U3706 (N_3706,N_739,N_2123);
or U3707 (N_3707,N_2010,N_1886);
xor U3708 (N_3708,N_201,N_1695);
and U3709 (N_3709,N_883,N_1840);
xor U3710 (N_3710,N_23,N_1332);
nor U3711 (N_3711,N_2335,N_1245);
xor U3712 (N_3712,N_1241,N_1221);
nor U3713 (N_3713,N_641,N_213);
xor U3714 (N_3714,N_267,N_1852);
nand U3715 (N_3715,N_157,N_42);
nor U3716 (N_3716,N_1415,N_781);
or U3717 (N_3717,N_1725,N_2349);
or U3718 (N_3718,N_2327,N_810);
and U3719 (N_3719,N_101,N_1049);
and U3720 (N_3720,N_1409,N_1059);
nand U3721 (N_3721,N_1569,N_1919);
and U3722 (N_3722,N_262,N_656);
nor U3723 (N_3723,N_1468,N_1107);
xor U3724 (N_3724,N_19,N_2134);
and U3725 (N_3725,N_770,N_1678);
nor U3726 (N_3726,N_2012,N_1961);
nand U3727 (N_3727,N_1900,N_1634);
nand U3728 (N_3728,N_1431,N_2137);
nand U3729 (N_3729,N_1615,N_842);
or U3730 (N_3730,N_1334,N_385);
or U3731 (N_3731,N_828,N_1383);
or U3732 (N_3732,N_759,N_1220);
xnor U3733 (N_3733,N_2457,N_2117);
nand U3734 (N_3734,N_1717,N_500);
xor U3735 (N_3735,N_1540,N_864);
and U3736 (N_3736,N_1222,N_2441);
and U3737 (N_3737,N_1504,N_2348);
xor U3738 (N_3738,N_221,N_417);
and U3739 (N_3739,N_1786,N_1767);
or U3740 (N_3740,N_1273,N_1350);
nor U3741 (N_3741,N_756,N_1965);
nand U3742 (N_3742,N_1196,N_322);
and U3743 (N_3743,N_356,N_580);
nand U3744 (N_3744,N_811,N_373);
nor U3745 (N_3745,N_929,N_2073);
and U3746 (N_3746,N_2215,N_2139);
nand U3747 (N_3747,N_2393,N_2145);
nor U3748 (N_3748,N_1357,N_942);
xnor U3749 (N_3749,N_2047,N_1061);
nor U3750 (N_3750,N_2264,N_290);
nand U3751 (N_3751,N_9,N_1152);
nor U3752 (N_3752,N_1148,N_1684);
xnor U3753 (N_3753,N_1348,N_813);
nand U3754 (N_3754,N_1407,N_1221);
and U3755 (N_3755,N_567,N_40);
nor U3756 (N_3756,N_312,N_515);
and U3757 (N_3757,N_676,N_1512);
nor U3758 (N_3758,N_95,N_2404);
or U3759 (N_3759,N_1144,N_1985);
and U3760 (N_3760,N_113,N_2476);
or U3761 (N_3761,N_1144,N_724);
xor U3762 (N_3762,N_2356,N_2040);
and U3763 (N_3763,N_443,N_1980);
nand U3764 (N_3764,N_2386,N_92);
nand U3765 (N_3765,N_1155,N_2412);
nand U3766 (N_3766,N_1835,N_1707);
nor U3767 (N_3767,N_2340,N_1330);
or U3768 (N_3768,N_2348,N_1240);
nand U3769 (N_3769,N_791,N_1431);
xor U3770 (N_3770,N_131,N_2183);
nand U3771 (N_3771,N_229,N_1525);
or U3772 (N_3772,N_745,N_1663);
xnor U3773 (N_3773,N_1282,N_670);
xnor U3774 (N_3774,N_712,N_61);
or U3775 (N_3775,N_1825,N_243);
xnor U3776 (N_3776,N_262,N_1950);
nand U3777 (N_3777,N_1905,N_1483);
or U3778 (N_3778,N_326,N_504);
xor U3779 (N_3779,N_278,N_233);
nand U3780 (N_3780,N_1334,N_1591);
xnor U3781 (N_3781,N_1709,N_1856);
xor U3782 (N_3782,N_1956,N_1497);
and U3783 (N_3783,N_1809,N_1262);
nand U3784 (N_3784,N_588,N_1344);
or U3785 (N_3785,N_2400,N_2212);
or U3786 (N_3786,N_2487,N_326);
and U3787 (N_3787,N_1748,N_195);
and U3788 (N_3788,N_2053,N_968);
and U3789 (N_3789,N_1590,N_467);
nor U3790 (N_3790,N_977,N_1997);
and U3791 (N_3791,N_2327,N_1965);
nor U3792 (N_3792,N_1586,N_1392);
and U3793 (N_3793,N_2250,N_749);
nor U3794 (N_3794,N_1132,N_2382);
nor U3795 (N_3795,N_65,N_2009);
nand U3796 (N_3796,N_1736,N_1113);
nand U3797 (N_3797,N_1968,N_984);
xor U3798 (N_3798,N_259,N_2170);
xor U3799 (N_3799,N_997,N_924);
xnor U3800 (N_3800,N_1438,N_1870);
nand U3801 (N_3801,N_674,N_501);
and U3802 (N_3802,N_1166,N_2143);
or U3803 (N_3803,N_101,N_1722);
nand U3804 (N_3804,N_3,N_1281);
nand U3805 (N_3805,N_65,N_1321);
nand U3806 (N_3806,N_1659,N_576);
xnor U3807 (N_3807,N_1533,N_2364);
or U3808 (N_3808,N_1180,N_490);
and U3809 (N_3809,N_1984,N_1049);
and U3810 (N_3810,N_35,N_300);
xnor U3811 (N_3811,N_2393,N_697);
xor U3812 (N_3812,N_1604,N_1506);
nand U3813 (N_3813,N_2272,N_644);
xor U3814 (N_3814,N_300,N_928);
xor U3815 (N_3815,N_2263,N_1475);
or U3816 (N_3816,N_2312,N_2157);
nor U3817 (N_3817,N_483,N_2412);
nand U3818 (N_3818,N_2049,N_226);
or U3819 (N_3819,N_2292,N_2340);
nor U3820 (N_3820,N_174,N_1880);
nand U3821 (N_3821,N_1352,N_228);
nand U3822 (N_3822,N_1173,N_2313);
and U3823 (N_3823,N_859,N_965);
nand U3824 (N_3824,N_8,N_18);
or U3825 (N_3825,N_575,N_2378);
or U3826 (N_3826,N_988,N_674);
xnor U3827 (N_3827,N_1092,N_698);
xor U3828 (N_3828,N_712,N_779);
and U3829 (N_3829,N_2119,N_989);
or U3830 (N_3830,N_795,N_1808);
or U3831 (N_3831,N_954,N_1423);
nand U3832 (N_3832,N_2254,N_1612);
xnor U3833 (N_3833,N_829,N_91);
or U3834 (N_3834,N_1103,N_2187);
and U3835 (N_3835,N_549,N_2466);
nor U3836 (N_3836,N_536,N_2288);
and U3837 (N_3837,N_788,N_1534);
nor U3838 (N_3838,N_1949,N_648);
or U3839 (N_3839,N_182,N_662);
xnor U3840 (N_3840,N_1329,N_400);
nand U3841 (N_3841,N_2174,N_2127);
nor U3842 (N_3842,N_2377,N_989);
nand U3843 (N_3843,N_1197,N_756);
and U3844 (N_3844,N_1483,N_2301);
xnor U3845 (N_3845,N_1870,N_793);
nand U3846 (N_3846,N_851,N_283);
xor U3847 (N_3847,N_616,N_1148);
xnor U3848 (N_3848,N_2053,N_2448);
and U3849 (N_3849,N_2460,N_419);
nor U3850 (N_3850,N_1959,N_2099);
nand U3851 (N_3851,N_1872,N_2435);
and U3852 (N_3852,N_2477,N_567);
and U3853 (N_3853,N_1633,N_2035);
nor U3854 (N_3854,N_429,N_1763);
nor U3855 (N_3855,N_1188,N_1397);
nor U3856 (N_3856,N_86,N_512);
and U3857 (N_3857,N_1263,N_1892);
nand U3858 (N_3858,N_1300,N_1358);
nand U3859 (N_3859,N_461,N_896);
or U3860 (N_3860,N_970,N_2082);
and U3861 (N_3861,N_387,N_1886);
xnor U3862 (N_3862,N_129,N_1832);
nand U3863 (N_3863,N_381,N_571);
and U3864 (N_3864,N_2339,N_1033);
or U3865 (N_3865,N_1923,N_173);
xor U3866 (N_3866,N_11,N_2457);
xnor U3867 (N_3867,N_1983,N_1563);
nor U3868 (N_3868,N_80,N_840);
nor U3869 (N_3869,N_2026,N_60);
xor U3870 (N_3870,N_184,N_1750);
nand U3871 (N_3871,N_1079,N_359);
or U3872 (N_3872,N_80,N_772);
nand U3873 (N_3873,N_158,N_179);
nand U3874 (N_3874,N_478,N_923);
or U3875 (N_3875,N_2063,N_1959);
xor U3876 (N_3876,N_1475,N_1029);
or U3877 (N_3877,N_799,N_802);
or U3878 (N_3878,N_191,N_393);
xor U3879 (N_3879,N_1853,N_1777);
nor U3880 (N_3880,N_127,N_775);
nand U3881 (N_3881,N_469,N_375);
nand U3882 (N_3882,N_675,N_2057);
nand U3883 (N_3883,N_617,N_377);
or U3884 (N_3884,N_482,N_2192);
or U3885 (N_3885,N_249,N_1788);
or U3886 (N_3886,N_909,N_1472);
nand U3887 (N_3887,N_532,N_617);
xnor U3888 (N_3888,N_2308,N_1769);
or U3889 (N_3889,N_1117,N_748);
and U3890 (N_3890,N_286,N_1463);
nor U3891 (N_3891,N_1561,N_1446);
and U3892 (N_3892,N_1766,N_2231);
or U3893 (N_3893,N_1201,N_2185);
nor U3894 (N_3894,N_2322,N_1419);
nand U3895 (N_3895,N_484,N_2203);
nor U3896 (N_3896,N_864,N_2136);
and U3897 (N_3897,N_1331,N_1795);
or U3898 (N_3898,N_126,N_648);
xor U3899 (N_3899,N_1633,N_1865);
or U3900 (N_3900,N_1380,N_1245);
nand U3901 (N_3901,N_814,N_2045);
nand U3902 (N_3902,N_1826,N_2154);
nand U3903 (N_3903,N_677,N_2388);
nor U3904 (N_3904,N_454,N_2282);
and U3905 (N_3905,N_1442,N_193);
or U3906 (N_3906,N_360,N_1682);
xnor U3907 (N_3907,N_474,N_1750);
or U3908 (N_3908,N_1667,N_1228);
nand U3909 (N_3909,N_805,N_696);
or U3910 (N_3910,N_1339,N_280);
nand U3911 (N_3911,N_2344,N_827);
xnor U3912 (N_3912,N_59,N_822);
or U3913 (N_3913,N_354,N_969);
or U3914 (N_3914,N_1936,N_1192);
or U3915 (N_3915,N_1358,N_2475);
xor U3916 (N_3916,N_2229,N_814);
nor U3917 (N_3917,N_1896,N_1813);
or U3918 (N_3918,N_608,N_1285);
nand U3919 (N_3919,N_774,N_1262);
nor U3920 (N_3920,N_1790,N_317);
xnor U3921 (N_3921,N_886,N_573);
or U3922 (N_3922,N_1895,N_116);
xnor U3923 (N_3923,N_407,N_1332);
nor U3924 (N_3924,N_1866,N_1088);
xnor U3925 (N_3925,N_1718,N_527);
xnor U3926 (N_3926,N_703,N_1404);
or U3927 (N_3927,N_951,N_239);
xnor U3928 (N_3928,N_1931,N_1234);
nand U3929 (N_3929,N_220,N_1870);
and U3930 (N_3930,N_781,N_1861);
nand U3931 (N_3931,N_397,N_910);
xor U3932 (N_3932,N_933,N_199);
nand U3933 (N_3933,N_288,N_442);
xor U3934 (N_3934,N_221,N_2328);
or U3935 (N_3935,N_616,N_1482);
and U3936 (N_3936,N_888,N_1159);
and U3937 (N_3937,N_1499,N_1952);
or U3938 (N_3938,N_1410,N_1031);
or U3939 (N_3939,N_674,N_2019);
or U3940 (N_3940,N_553,N_2232);
xor U3941 (N_3941,N_2422,N_1316);
nand U3942 (N_3942,N_1623,N_1027);
xor U3943 (N_3943,N_2101,N_2303);
or U3944 (N_3944,N_1821,N_2231);
nor U3945 (N_3945,N_561,N_2322);
xor U3946 (N_3946,N_459,N_1767);
nor U3947 (N_3947,N_98,N_1231);
or U3948 (N_3948,N_1394,N_1067);
xor U3949 (N_3949,N_1696,N_2440);
xor U3950 (N_3950,N_209,N_1608);
or U3951 (N_3951,N_1504,N_1823);
nor U3952 (N_3952,N_1986,N_36);
nor U3953 (N_3953,N_417,N_1153);
and U3954 (N_3954,N_1031,N_788);
nor U3955 (N_3955,N_2450,N_321);
nand U3956 (N_3956,N_639,N_1182);
or U3957 (N_3957,N_1894,N_1023);
xor U3958 (N_3958,N_1181,N_2273);
or U3959 (N_3959,N_1914,N_2046);
nor U3960 (N_3960,N_1610,N_409);
or U3961 (N_3961,N_885,N_1795);
nor U3962 (N_3962,N_508,N_1085);
xor U3963 (N_3963,N_1684,N_1835);
nand U3964 (N_3964,N_1213,N_1534);
xnor U3965 (N_3965,N_2091,N_178);
xnor U3966 (N_3966,N_890,N_660);
or U3967 (N_3967,N_906,N_377);
nor U3968 (N_3968,N_1246,N_1670);
nand U3969 (N_3969,N_1693,N_1043);
or U3970 (N_3970,N_2271,N_540);
xnor U3971 (N_3971,N_1716,N_2302);
nor U3972 (N_3972,N_398,N_230);
and U3973 (N_3973,N_2382,N_319);
nor U3974 (N_3974,N_1294,N_1002);
nand U3975 (N_3975,N_1612,N_520);
xor U3976 (N_3976,N_732,N_581);
and U3977 (N_3977,N_464,N_2416);
or U3978 (N_3978,N_1938,N_516);
or U3979 (N_3979,N_2358,N_66);
nor U3980 (N_3980,N_551,N_1818);
xor U3981 (N_3981,N_861,N_1811);
nor U3982 (N_3982,N_691,N_724);
or U3983 (N_3983,N_1921,N_990);
and U3984 (N_3984,N_2305,N_308);
and U3985 (N_3985,N_1520,N_1102);
or U3986 (N_3986,N_1344,N_1176);
or U3987 (N_3987,N_801,N_2298);
or U3988 (N_3988,N_964,N_1822);
nor U3989 (N_3989,N_726,N_1899);
nor U3990 (N_3990,N_907,N_1991);
and U3991 (N_3991,N_1594,N_520);
nand U3992 (N_3992,N_17,N_1631);
nand U3993 (N_3993,N_2371,N_140);
and U3994 (N_3994,N_1570,N_2301);
xor U3995 (N_3995,N_1981,N_1420);
nor U3996 (N_3996,N_146,N_232);
or U3997 (N_3997,N_1827,N_1174);
and U3998 (N_3998,N_1119,N_2377);
or U3999 (N_3999,N_349,N_52);
nand U4000 (N_4000,N_580,N_2432);
nor U4001 (N_4001,N_2489,N_1752);
and U4002 (N_4002,N_2221,N_92);
nand U4003 (N_4003,N_2105,N_1818);
and U4004 (N_4004,N_1755,N_1152);
and U4005 (N_4005,N_1244,N_1721);
or U4006 (N_4006,N_2279,N_1832);
and U4007 (N_4007,N_1729,N_2480);
nand U4008 (N_4008,N_792,N_2433);
and U4009 (N_4009,N_2016,N_2283);
and U4010 (N_4010,N_524,N_1666);
nand U4011 (N_4011,N_2429,N_2302);
xor U4012 (N_4012,N_1599,N_281);
and U4013 (N_4013,N_1802,N_516);
xor U4014 (N_4014,N_2215,N_1660);
nor U4015 (N_4015,N_196,N_1368);
nand U4016 (N_4016,N_2131,N_591);
nand U4017 (N_4017,N_1736,N_2459);
nand U4018 (N_4018,N_352,N_2352);
xor U4019 (N_4019,N_817,N_1897);
nor U4020 (N_4020,N_2401,N_27);
xor U4021 (N_4021,N_548,N_2178);
and U4022 (N_4022,N_2398,N_2093);
nor U4023 (N_4023,N_2407,N_1968);
and U4024 (N_4024,N_735,N_387);
xnor U4025 (N_4025,N_1699,N_911);
nor U4026 (N_4026,N_1331,N_635);
nor U4027 (N_4027,N_419,N_610);
nand U4028 (N_4028,N_373,N_1127);
and U4029 (N_4029,N_1939,N_110);
or U4030 (N_4030,N_1961,N_503);
xnor U4031 (N_4031,N_1868,N_592);
or U4032 (N_4032,N_699,N_461);
nand U4033 (N_4033,N_725,N_1446);
nand U4034 (N_4034,N_1971,N_1609);
or U4035 (N_4035,N_1056,N_1978);
or U4036 (N_4036,N_1487,N_531);
xor U4037 (N_4037,N_655,N_1148);
and U4038 (N_4038,N_316,N_695);
and U4039 (N_4039,N_19,N_670);
nand U4040 (N_4040,N_1888,N_1792);
xnor U4041 (N_4041,N_839,N_306);
nor U4042 (N_4042,N_744,N_70);
nand U4043 (N_4043,N_2325,N_735);
nand U4044 (N_4044,N_2134,N_2348);
xor U4045 (N_4045,N_1525,N_1392);
nand U4046 (N_4046,N_1216,N_300);
and U4047 (N_4047,N_1065,N_1255);
and U4048 (N_4048,N_1972,N_1534);
nor U4049 (N_4049,N_103,N_1100);
or U4050 (N_4050,N_1967,N_604);
xor U4051 (N_4051,N_2072,N_119);
or U4052 (N_4052,N_1492,N_438);
nand U4053 (N_4053,N_620,N_2258);
nor U4054 (N_4054,N_368,N_521);
or U4055 (N_4055,N_547,N_1765);
and U4056 (N_4056,N_1857,N_331);
xor U4057 (N_4057,N_1964,N_1230);
and U4058 (N_4058,N_1007,N_2079);
or U4059 (N_4059,N_1677,N_1753);
and U4060 (N_4060,N_376,N_2265);
xnor U4061 (N_4061,N_70,N_27);
and U4062 (N_4062,N_162,N_2386);
nand U4063 (N_4063,N_1523,N_964);
nand U4064 (N_4064,N_2499,N_1906);
nand U4065 (N_4065,N_29,N_1452);
and U4066 (N_4066,N_1893,N_109);
nand U4067 (N_4067,N_1215,N_124);
xor U4068 (N_4068,N_19,N_1857);
or U4069 (N_4069,N_258,N_1719);
nor U4070 (N_4070,N_2354,N_986);
and U4071 (N_4071,N_637,N_2498);
nor U4072 (N_4072,N_36,N_898);
nor U4073 (N_4073,N_2091,N_885);
nand U4074 (N_4074,N_759,N_189);
or U4075 (N_4075,N_731,N_2124);
or U4076 (N_4076,N_2072,N_1307);
and U4077 (N_4077,N_1468,N_2150);
xnor U4078 (N_4078,N_14,N_196);
nor U4079 (N_4079,N_2077,N_1378);
xor U4080 (N_4080,N_1140,N_175);
xnor U4081 (N_4081,N_97,N_1753);
xnor U4082 (N_4082,N_2009,N_2359);
xnor U4083 (N_4083,N_1461,N_995);
or U4084 (N_4084,N_1708,N_1317);
or U4085 (N_4085,N_686,N_935);
and U4086 (N_4086,N_533,N_448);
nor U4087 (N_4087,N_1202,N_2182);
nand U4088 (N_4088,N_2428,N_401);
nor U4089 (N_4089,N_1025,N_1726);
or U4090 (N_4090,N_1594,N_17);
nand U4091 (N_4091,N_1344,N_335);
xnor U4092 (N_4092,N_1028,N_320);
or U4093 (N_4093,N_246,N_2135);
xnor U4094 (N_4094,N_403,N_1346);
xor U4095 (N_4095,N_605,N_1867);
nand U4096 (N_4096,N_1390,N_1361);
or U4097 (N_4097,N_417,N_219);
xnor U4098 (N_4098,N_2342,N_5);
or U4099 (N_4099,N_303,N_1350);
or U4100 (N_4100,N_585,N_1844);
nand U4101 (N_4101,N_2436,N_1457);
xnor U4102 (N_4102,N_384,N_1606);
and U4103 (N_4103,N_2473,N_2025);
nor U4104 (N_4104,N_1562,N_1750);
and U4105 (N_4105,N_751,N_1319);
and U4106 (N_4106,N_1624,N_1447);
nor U4107 (N_4107,N_1955,N_463);
and U4108 (N_4108,N_1464,N_1165);
nand U4109 (N_4109,N_66,N_19);
nand U4110 (N_4110,N_499,N_529);
nor U4111 (N_4111,N_687,N_1385);
and U4112 (N_4112,N_1476,N_2009);
or U4113 (N_4113,N_1240,N_166);
nor U4114 (N_4114,N_1095,N_1923);
nand U4115 (N_4115,N_2129,N_1031);
xnor U4116 (N_4116,N_1220,N_1328);
nor U4117 (N_4117,N_2215,N_2412);
and U4118 (N_4118,N_855,N_1113);
or U4119 (N_4119,N_2380,N_1463);
nand U4120 (N_4120,N_538,N_1025);
nand U4121 (N_4121,N_1532,N_345);
nor U4122 (N_4122,N_2488,N_2151);
or U4123 (N_4123,N_364,N_508);
xor U4124 (N_4124,N_671,N_381);
nor U4125 (N_4125,N_532,N_1606);
nand U4126 (N_4126,N_2098,N_2395);
and U4127 (N_4127,N_1462,N_902);
and U4128 (N_4128,N_2180,N_1187);
nor U4129 (N_4129,N_143,N_2401);
nand U4130 (N_4130,N_444,N_971);
and U4131 (N_4131,N_1406,N_2328);
or U4132 (N_4132,N_1876,N_344);
xor U4133 (N_4133,N_1014,N_41);
xor U4134 (N_4134,N_997,N_1663);
and U4135 (N_4135,N_1363,N_2412);
xor U4136 (N_4136,N_1643,N_1120);
and U4137 (N_4137,N_1108,N_2265);
nor U4138 (N_4138,N_2121,N_2388);
xor U4139 (N_4139,N_2490,N_1914);
nor U4140 (N_4140,N_446,N_1303);
nor U4141 (N_4141,N_988,N_2390);
nor U4142 (N_4142,N_307,N_1724);
xor U4143 (N_4143,N_2311,N_1811);
or U4144 (N_4144,N_253,N_2449);
and U4145 (N_4145,N_1529,N_1055);
and U4146 (N_4146,N_607,N_97);
xnor U4147 (N_4147,N_368,N_469);
nor U4148 (N_4148,N_906,N_977);
or U4149 (N_4149,N_218,N_1261);
xnor U4150 (N_4150,N_117,N_92);
nor U4151 (N_4151,N_2421,N_1880);
nor U4152 (N_4152,N_1402,N_2349);
xor U4153 (N_4153,N_2497,N_353);
or U4154 (N_4154,N_2471,N_546);
nand U4155 (N_4155,N_208,N_487);
and U4156 (N_4156,N_1925,N_649);
nor U4157 (N_4157,N_237,N_2021);
xnor U4158 (N_4158,N_1348,N_657);
xnor U4159 (N_4159,N_1974,N_136);
or U4160 (N_4160,N_1910,N_1055);
and U4161 (N_4161,N_1194,N_446);
nand U4162 (N_4162,N_804,N_1729);
and U4163 (N_4163,N_2378,N_1344);
and U4164 (N_4164,N_1479,N_114);
xnor U4165 (N_4165,N_2459,N_1047);
or U4166 (N_4166,N_2098,N_2183);
xnor U4167 (N_4167,N_456,N_1476);
nand U4168 (N_4168,N_979,N_223);
nand U4169 (N_4169,N_405,N_87);
nor U4170 (N_4170,N_527,N_832);
nor U4171 (N_4171,N_2172,N_705);
and U4172 (N_4172,N_231,N_1707);
or U4173 (N_4173,N_112,N_290);
xor U4174 (N_4174,N_2374,N_2497);
or U4175 (N_4175,N_1961,N_231);
or U4176 (N_4176,N_2279,N_251);
xor U4177 (N_4177,N_263,N_453);
nor U4178 (N_4178,N_1585,N_1011);
nor U4179 (N_4179,N_1742,N_1406);
nor U4180 (N_4180,N_658,N_956);
nand U4181 (N_4181,N_1464,N_1258);
xnor U4182 (N_4182,N_814,N_677);
or U4183 (N_4183,N_900,N_1111);
xnor U4184 (N_4184,N_266,N_1990);
xor U4185 (N_4185,N_1978,N_640);
and U4186 (N_4186,N_1768,N_320);
or U4187 (N_4187,N_2103,N_1248);
or U4188 (N_4188,N_560,N_650);
and U4189 (N_4189,N_2199,N_834);
nor U4190 (N_4190,N_296,N_1080);
xor U4191 (N_4191,N_1376,N_1872);
xnor U4192 (N_4192,N_1784,N_1073);
xnor U4193 (N_4193,N_2314,N_2128);
nand U4194 (N_4194,N_2095,N_171);
nand U4195 (N_4195,N_2379,N_1309);
nand U4196 (N_4196,N_2191,N_1495);
or U4197 (N_4197,N_683,N_1800);
or U4198 (N_4198,N_2332,N_314);
xnor U4199 (N_4199,N_440,N_2380);
nand U4200 (N_4200,N_1806,N_444);
or U4201 (N_4201,N_1234,N_494);
xor U4202 (N_4202,N_475,N_180);
and U4203 (N_4203,N_1487,N_1814);
xor U4204 (N_4204,N_938,N_2403);
nor U4205 (N_4205,N_1422,N_1894);
or U4206 (N_4206,N_896,N_983);
or U4207 (N_4207,N_1975,N_457);
or U4208 (N_4208,N_1272,N_2149);
nor U4209 (N_4209,N_1153,N_2495);
nand U4210 (N_4210,N_1147,N_1957);
and U4211 (N_4211,N_104,N_1378);
and U4212 (N_4212,N_1775,N_2033);
nor U4213 (N_4213,N_1064,N_1545);
and U4214 (N_4214,N_1487,N_878);
xnor U4215 (N_4215,N_1180,N_2497);
xor U4216 (N_4216,N_758,N_225);
and U4217 (N_4217,N_638,N_151);
nor U4218 (N_4218,N_1194,N_1616);
nand U4219 (N_4219,N_438,N_1039);
nor U4220 (N_4220,N_2123,N_972);
and U4221 (N_4221,N_2375,N_251);
xnor U4222 (N_4222,N_192,N_1979);
and U4223 (N_4223,N_933,N_2400);
and U4224 (N_4224,N_1624,N_781);
xor U4225 (N_4225,N_1685,N_560);
and U4226 (N_4226,N_1623,N_165);
nand U4227 (N_4227,N_1029,N_1457);
nor U4228 (N_4228,N_1054,N_668);
and U4229 (N_4229,N_1222,N_320);
and U4230 (N_4230,N_712,N_138);
nor U4231 (N_4231,N_114,N_1337);
and U4232 (N_4232,N_1453,N_36);
nand U4233 (N_4233,N_834,N_1801);
and U4234 (N_4234,N_1666,N_1113);
xnor U4235 (N_4235,N_1824,N_356);
nand U4236 (N_4236,N_1836,N_846);
xor U4237 (N_4237,N_562,N_1008);
xor U4238 (N_4238,N_1908,N_1253);
xnor U4239 (N_4239,N_1515,N_686);
nor U4240 (N_4240,N_1597,N_425);
and U4241 (N_4241,N_208,N_394);
nand U4242 (N_4242,N_403,N_582);
nor U4243 (N_4243,N_1726,N_2051);
nand U4244 (N_4244,N_1741,N_515);
nor U4245 (N_4245,N_2326,N_1524);
nor U4246 (N_4246,N_2132,N_938);
nor U4247 (N_4247,N_2124,N_1308);
xor U4248 (N_4248,N_1489,N_673);
and U4249 (N_4249,N_452,N_2196);
nand U4250 (N_4250,N_1418,N_457);
xnor U4251 (N_4251,N_583,N_188);
nand U4252 (N_4252,N_1186,N_46);
xnor U4253 (N_4253,N_557,N_653);
or U4254 (N_4254,N_2283,N_1665);
or U4255 (N_4255,N_124,N_2225);
nor U4256 (N_4256,N_1180,N_1197);
or U4257 (N_4257,N_2003,N_707);
xnor U4258 (N_4258,N_1734,N_2352);
nand U4259 (N_4259,N_207,N_1593);
or U4260 (N_4260,N_1014,N_1250);
nand U4261 (N_4261,N_1674,N_1233);
xnor U4262 (N_4262,N_504,N_1128);
nor U4263 (N_4263,N_1324,N_4);
or U4264 (N_4264,N_988,N_978);
and U4265 (N_4265,N_1280,N_661);
nor U4266 (N_4266,N_148,N_2261);
nor U4267 (N_4267,N_639,N_129);
or U4268 (N_4268,N_1147,N_1490);
nor U4269 (N_4269,N_441,N_34);
xnor U4270 (N_4270,N_1660,N_1653);
or U4271 (N_4271,N_2399,N_333);
nor U4272 (N_4272,N_301,N_457);
or U4273 (N_4273,N_293,N_2302);
xnor U4274 (N_4274,N_439,N_2301);
nor U4275 (N_4275,N_1161,N_1353);
and U4276 (N_4276,N_764,N_2034);
and U4277 (N_4277,N_1927,N_1216);
xor U4278 (N_4278,N_379,N_223);
xnor U4279 (N_4279,N_826,N_2101);
or U4280 (N_4280,N_605,N_1170);
nand U4281 (N_4281,N_1218,N_1418);
nand U4282 (N_4282,N_1866,N_349);
or U4283 (N_4283,N_1299,N_1116);
nor U4284 (N_4284,N_2173,N_355);
xor U4285 (N_4285,N_232,N_913);
nand U4286 (N_4286,N_2280,N_1936);
or U4287 (N_4287,N_1111,N_722);
nor U4288 (N_4288,N_1444,N_12);
nor U4289 (N_4289,N_1962,N_659);
nand U4290 (N_4290,N_2225,N_1319);
nor U4291 (N_4291,N_2487,N_590);
and U4292 (N_4292,N_1026,N_1772);
nand U4293 (N_4293,N_244,N_38);
or U4294 (N_4294,N_657,N_806);
nor U4295 (N_4295,N_2109,N_2078);
nor U4296 (N_4296,N_1739,N_1205);
xor U4297 (N_4297,N_1763,N_2311);
nor U4298 (N_4298,N_2308,N_823);
or U4299 (N_4299,N_451,N_997);
nor U4300 (N_4300,N_1937,N_517);
nor U4301 (N_4301,N_931,N_1564);
xor U4302 (N_4302,N_1511,N_978);
xor U4303 (N_4303,N_791,N_1190);
nand U4304 (N_4304,N_1352,N_238);
xor U4305 (N_4305,N_113,N_284);
nand U4306 (N_4306,N_2349,N_2285);
nor U4307 (N_4307,N_2392,N_2159);
nor U4308 (N_4308,N_554,N_1105);
nand U4309 (N_4309,N_2348,N_1979);
xor U4310 (N_4310,N_1817,N_2478);
nand U4311 (N_4311,N_1248,N_1763);
or U4312 (N_4312,N_976,N_1751);
nor U4313 (N_4313,N_2282,N_328);
xnor U4314 (N_4314,N_712,N_1223);
xor U4315 (N_4315,N_202,N_950);
nor U4316 (N_4316,N_1262,N_397);
nor U4317 (N_4317,N_875,N_972);
or U4318 (N_4318,N_136,N_1561);
nor U4319 (N_4319,N_633,N_478);
or U4320 (N_4320,N_463,N_1705);
or U4321 (N_4321,N_950,N_1076);
and U4322 (N_4322,N_1659,N_728);
or U4323 (N_4323,N_452,N_2029);
nor U4324 (N_4324,N_1037,N_2166);
xor U4325 (N_4325,N_1183,N_1850);
xnor U4326 (N_4326,N_837,N_1324);
and U4327 (N_4327,N_590,N_1795);
or U4328 (N_4328,N_1628,N_2331);
and U4329 (N_4329,N_2316,N_1989);
xor U4330 (N_4330,N_591,N_652);
or U4331 (N_4331,N_180,N_649);
nor U4332 (N_4332,N_1865,N_316);
xnor U4333 (N_4333,N_2430,N_1816);
or U4334 (N_4334,N_957,N_856);
and U4335 (N_4335,N_597,N_2400);
xnor U4336 (N_4336,N_2076,N_1955);
nor U4337 (N_4337,N_2235,N_1937);
nand U4338 (N_4338,N_2134,N_1997);
xor U4339 (N_4339,N_1195,N_1839);
nand U4340 (N_4340,N_2121,N_1030);
nor U4341 (N_4341,N_1926,N_1809);
xor U4342 (N_4342,N_904,N_1008);
nand U4343 (N_4343,N_361,N_1515);
or U4344 (N_4344,N_1840,N_2099);
xnor U4345 (N_4345,N_2110,N_2385);
xnor U4346 (N_4346,N_1125,N_1966);
and U4347 (N_4347,N_1678,N_200);
xor U4348 (N_4348,N_1873,N_719);
or U4349 (N_4349,N_1116,N_1506);
nor U4350 (N_4350,N_1526,N_1970);
nand U4351 (N_4351,N_475,N_2084);
or U4352 (N_4352,N_63,N_1249);
xor U4353 (N_4353,N_1632,N_630);
and U4354 (N_4354,N_102,N_707);
xor U4355 (N_4355,N_1253,N_1762);
nor U4356 (N_4356,N_315,N_1092);
and U4357 (N_4357,N_1811,N_1563);
xnor U4358 (N_4358,N_1433,N_1762);
and U4359 (N_4359,N_1798,N_1838);
nor U4360 (N_4360,N_217,N_2394);
and U4361 (N_4361,N_2459,N_970);
or U4362 (N_4362,N_2351,N_2131);
xnor U4363 (N_4363,N_1089,N_1772);
xor U4364 (N_4364,N_772,N_1291);
nor U4365 (N_4365,N_2157,N_1138);
nand U4366 (N_4366,N_2463,N_646);
xnor U4367 (N_4367,N_2019,N_2437);
nor U4368 (N_4368,N_806,N_2034);
and U4369 (N_4369,N_1325,N_2201);
and U4370 (N_4370,N_415,N_1404);
or U4371 (N_4371,N_1296,N_1458);
and U4372 (N_4372,N_814,N_1743);
or U4373 (N_4373,N_2019,N_1632);
nand U4374 (N_4374,N_1201,N_866);
nand U4375 (N_4375,N_1234,N_788);
and U4376 (N_4376,N_2491,N_1495);
nand U4377 (N_4377,N_957,N_893);
nand U4378 (N_4378,N_2355,N_760);
and U4379 (N_4379,N_1722,N_1187);
nand U4380 (N_4380,N_958,N_476);
and U4381 (N_4381,N_1566,N_2384);
nor U4382 (N_4382,N_2388,N_2285);
nor U4383 (N_4383,N_120,N_787);
nand U4384 (N_4384,N_885,N_888);
nor U4385 (N_4385,N_711,N_1606);
xor U4386 (N_4386,N_1765,N_2305);
nand U4387 (N_4387,N_223,N_1806);
xor U4388 (N_4388,N_472,N_1612);
and U4389 (N_4389,N_995,N_2155);
or U4390 (N_4390,N_611,N_97);
or U4391 (N_4391,N_1541,N_2258);
or U4392 (N_4392,N_284,N_2113);
or U4393 (N_4393,N_404,N_2019);
xnor U4394 (N_4394,N_554,N_2372);
xor U4395 (N_4395,N_1982,N_1168);
xnor U4396 (N_4396,N_948,N_1810);
and U4397 (N_4397,N_1507,N_2241);
nand U4398 (N_4398,N_688,N_745);
nor U4399 (N_4399,N_81,N_1193);
nand U4400 (N_4400,N_2113,N_1127);
or U4401 (N_4401,N_495,N_1811);
and U4402 (N_4402,N_1957,N_746);
nor U4403 (N_4403,N_13,N_2172);
nor U4404 (N_4404,N_1581,N_465);
nand U4405 (N_4405,N_1228,N_1759);
nand U4406 (N_4406,N_2018,N_413);
or U4407 (N_4407,N_894,N_2061);
nor U4408 (N_4408,N_1580,N_1317);
and U4409 (N_4409,N_1973,N_713);
or U4410 (N_4410,N_152,N_2281);
and U4411 (N_4411,N_1147,N_323);
nor U4412 (N_4412,N_1797,N_1863);
xnor U4413 (N_4413,N_1108,N_1178);
or U4414 (N_4414,N_2445,N_1517);
and U4415 (N_4415,N_896,N_1365);
nand U4416 (N_4416,N_1450,N_1456);
nor U4417 (N_4417,N_878,N_692);
and U4418 (N_4418,N_1013,N_321);
nand U4419 (N_4419,N_753,N_777);
xnor U4420 (N_4420,N_549,N_1181);
xnor U4421 (N_4421,N_261,N_881);
xnor U4422 (N_4422,N_2171,N_83);
xor U4423 (N_4423,N_1219,N_961);
nand U4424 (N_4424,N_368,N_257);
or U4425 (N_4425,N_2327,N_1235);
nor U4426 (N_4426,N_2189,N_1367);
and U4427 (N_4427,N_919,N_2363);
or U4428 (N_4428,N_2387,N_1776);
xnor U4429 (N_4429,N_1963,N_262);
nand U4430 (N_4430,N_1894,N_136);
or U4431 (N_4431,N_2165,N_517);
nor U4432 (N_4432,N_464,N_1921);
or U4433 (N_4433,N_279,N_294);
or U4434 (N_4434,N_408,N_2377);
xnor U4435 (N_4435,N_571,N_1606);
and U4436 (N_4436,N_2167,N_1177);
and U4437 (N_4437,N_688,N_183);
xnor U4438 (N_4438,N_1864,N_758);
xor U4439 (N_4439,N_1056,N_715);
and U4440 (N_4440,N_1555,N_967);
xnor U4441 (N_4441,N_1650,N_2020);
xor U4442 (N_4442,N_2452,N_1375);
nand U4443 (N_4443,N_905,N_1401);
nor U4444 (N_4444,N_780,N_970);
and U4445 (N_4445,N_1063,N_260);
nor U4446 (N_4446,N_2066,N_1345);
or U4447 (N_4447,N_2323,N_1396);
nor U4448 (N_4448,N_1397,N_2188);
and U4449 (N_4449,N_1667,N_2392);
nand U4450 (N_4450,N_547,N_1389);
or U4451 (N_4451,N_805,N_731);
or U4452 (N_4452,N_1921,N_1834);
or U4453 (N_4453,N_1975,N_2035);
or U4454 (N_4454,N_14,N_2491);
xnor U4455 (N_4455,N_922,N_640);
xor U4456 (N_4456,N_1414,N_1364);
nor U4457 (N_4457,N_126,N_398);
and U4458 (N_4458,N_1640,N_1617);
or U4459 (N_4459,N_154,N_1862);
or U4460 (N_4460,N_2193,N_133);
xnor U4461 (N_4461,N_1952,N_112);
xor U4462 (N_4462,N_196,N_2162);
xnor U4463 (N_4463,N_1031,N_86);
and U4464 (N_4464,N_1507,N_1122);
or U4465 (N_4465,N_169,N_604);
xor U4466 (N_4466,N_68,N_1684);
nor U4467 (N_4467,N_1858,N_721);
and U4468 (N_4468,N_533,N_2084);
and U4469 (N_4469,N_936,N_2078);
and U4470 (N_4470,N_2256,N_499);
xnor U4471 (N_4471,N_47,N_1434);
nor U4472 (N_4472,N_980,N_309);
nor U4473 (N_4473,N_1851,N_313);
xnor U4474 (N_4474,N_1225,N_1322);
nand U4475 (N_4475,N_1936,N_1994);
nor U4476 (N_4476,N_455,N_2136);
or U4477 (N_4477,N_793,N_1035);
or U4478 (N_4478,N_2443,N_1514);
xnor U4479 (N_4479,N_1137,N_1258);
or U4480 (N_4480,N_1959,N_1130);
xnor U4481 (N_4481,N_2469,N_1815);
xnor U4482 (N_4482,N_2233,N_1164);
or U4483 (N_4483,N_1497,N_2301);
xnor U4484 (N_4484,N_33,N_331);
nand U4485 (N_4485,N_1093,N_2319);
and U4486 (N_4486,N_1961,N_1872);
xor U4487 (N_4487,N_913,N_1550);
xnor U4488 (N_4488,N_1665,N_1416);
nand U4489 (N_4489,N_2269,N_65);
and U4490 (N_4490,N_2343,N_844);
nand U4491 (N_4491,N_738,N_183);
xor U4492 (N_4492,N_1494,N_2069);
and U4493 (N_4493,N_2237,N_1450);
or U4494 (N_4494,N_743,N_1065);
or U4495 (N_4495,N_128,N_859);
nand U4496 (N_4496,N_1880,N_2427);
nor U4497 (N_4497,N_871,N_193);
and U4498 (N_4498,N_2068,N_448);
or U4499 (N_4499,N_1333,N_870);
xnor U4500 (N_4500,N_2486,N_1194);
or U4501 (N_4501,N_1072,N_1611);
nand U4502 (N_4502,N_1771,N_1737);
nor U4503 (N_4503,N_1250,N_214);
or U4504 (N_4504,N_673,N_479);
nand U4505 (N_4505,N_2373,N_1222);
and U4506 (N_4506,N_2450,N_1259);
or U4507 (N_4507,N_1168,N_313);
or U4508 (N_4508,N_1645,N_317);
xor U4509 (N_4509,N_2207,N_476);
and U4510 (N_4510,N_2316,N_1527);
nor U4511 (N_4511,N_1216,N_942);
nor U4512 (N_4512,N_1185,N_843);
nand U4513 (N_4513,N_2404,N_370);
and U4514 (N_4514,N_1625,N_521);
and U4515 (N_4515,N_315,N_861);
xor U4516 (N_4516,N_405,N_937);
nand U4517 (N_4517,N_1301,N_1935);
nor U4518 (N_4518,N_62,N_598);
and U4519 (N_4519,N_330,N_2362);
and U4520 (N_4520,N_1540,N_944);
or U4521 (N_4521,N_390,N_1141);
or U4522 (N_4522,N_874,N_305);
xor U4523 (N_4523,N_697,N_127);
and U4524 (N_4524,N_22,N_993);
nand U4525 (N_4525,N_1220,N_473);
xnor U4526 (N_4526,N_86,N_1220);
nor U4527 (N_4527,N_1078,N_1487);
xor U4528 (N_4528,N_51,N_46);
and U4529 (N_4529,N_849,N_345);
xnor U4530 (N_4530,N_316,N_2086);
nor U4531 (N_4531,N_161,N_1939);
and U4532 (N_4532,N_819,N_2168);
nor U4533 (N_4533,N_2180,N_2410);
xor U4534 (N_4534,N_2013,N_1463);
nor U4535 (N_4535,N_288,N_1888);
nand U4536 (N_4536,N_1347,N_2296);
xor U4537 (N_4537,N_2175,N_1812);
nand U4538 (N_4538,N_1654,N_1362);
and U4539 (N_4539,N_632,N_2094);
or U4540 (N_4540,N_945,N_7);
or U4541 (N_4541,N_509,N_2397);
xor U4542 (N_4542,N_2042,N_535);
xor U4543 (N_4543,N_1314,N_1829);
and U4544 (N_4544,N_51,N_1701);
nor U4545 (N_4545,N_976,N_703);
nand U4546 (N_4546,N_1021,N_261);
or U4547 (N_4547,N_1880,N_382);
nor U4548 (N_4548,N_1462,N_2016);
and U4549 (N_4549,N_1583,N_608);
or U4550 (N_4550,N_1371,N_497);
nand U4551 (N_4551,N_1300,N_2259);
nor U4552 (N_4552,N_1616,N_664);
or U4553 (N_4553,N_344,N_1570);
nor U4554 (N_4554,N_1937,N_243);
nor U4555 (N_4555,N_620,N_770);
nor U4556 (N_4556,N_2009,N_1423);
nand U4557 (N_4557,N_1089,N_489);
nand U4558 (N_4558,N_870,N_2493);
nor U4559 (N_4559,N_826,N_1644);
nor U4560 (N_4560,N_1867,N_1349);
xnor U4561 (N_4561,N_664,N_697);
or U4562 (N_4562,N_2097,N_1044);
nor U4563 (N_4563,N_2057,N_904);
xor U4564 (N_4564,N_1554,N_333);
nand U4565 (N_4565,N_1028,N_1347);
and U4566 (N_4566,N_1980,N_2490);
and U4567 (N_4567,N_36,N_1312);
nand U4568 (N_4568,N_1432,N_2242);
and U4569 (N_4569,N_1474,N_1176);
nand U4570 (N_4570,N_502,N_665);
or U4571 (N_4571,N_1667,N_832);
and U4572 (N_4572,N_2435,N_1263);
nand U4573 (N_4573,N_80,N_1730);
xor U4574 (N_4574,N_481,N_337);
and U4575 (N_4575,N_844,N_79);
nand U4576 (N_4576,N_286,N_375);
xnor U4577 (N_4577,N_1448,N_499);
nand U4578 (N_4578,N_1301,N_270);
and U4579 (N_4579,N_636,N_1731);
xnor U4580 (N_4580,N_1601,N_2012);
and U4581 (N_4581,N_127,N_1812);
nand U4582 (N_4582,N_407,N_2488);
and U4583 (N_4583,N_1324,N_1706);
or U4584 (N_4584,N_121,N_1037);
and U4585 (N_4585,N_1265,N_956);
xnor U4586 (N_4586,N_407,N_2009);
or U4587 (N_4587,N_308,N_2119);
or U4588 (N_4588,N_1294,N_980);
xor U4589 (N_4589,N_1260,N_1999);
or U4590 (N_4590,N_1783,N_2231);
and U4591 (N_4591,N_672,N_1248);
and U4592 (N_4592,N_1259,N_436);
nor U4593 (N_4593,N_2431,N_635);
xnor U4594 (N_4594,N_91,N_1214);
nor U4595 (N_4595,N_2091,N_1750);
or U4596 (N_4596,N_656,N_198);
and U4597 (N_4597,N_1457,N_752);
xnor U4598 (N_4598,N_2345,N_148);
xnor U4599 (N_4599,N_1227,N_1776);
xnor U4600 (N_4600,N_731,N_618);
or U4601 (N_4601,N_1344,N_1789);
nor U4602 (N_4602,N_582,N_2067);
nor U4603 (N_4603,N_2052,N_389);
nor U4604 (N_4604,N_2410,N_603);
nand U4605 (N_4605,N_1173,N_941);
nand U4606 (N_4606,N_387,N_2231);
nand U4607 (N_4607,N_1250,N_425);
nand U4608 (N_4608,N_326,N_333);
nand U4609 (N_4609,N_1395,N_1105);
nor U4610 (N_4610,N_738,N_495);
nand U4611 (N_4611,N_867,N_2223);
nand U4612 (N_4612,N_872,N_1004);
nor U4613 (N_4613,N_1171,N_88);
nand U4614 (N_4614,N_2370,N_1985);
nand U4615 (N_4615,N_1723,N_716);
xnor U4616 (N_4616,N_1382,N_1210);
and U4617 (N_4617,N_142,N_2498);
nand U4618 (N_4618,N_572,N_583);
or U4619 (N_4619,N_1466,N_53);
nand U4620 (N_4620,N_1599,N_2466);
or U4621 (N_4621,N_269,N_484);
nand U4622 (N_4622,N_274,N_341);
nor U4623 (N_4623,N_362,N_820);
xor U4624 (N_4624,N_976,N_1832);
xnor U4625 (N_4625,N_898,N_727);
or U4626 (N_4626,N_1522,N_1770);
or U4627 (N_4627,N_1100,N_2162);
and U4628 (N_4628,N_1813,N_1673);
and U4629 (N_4629,N_2193,N_1707);
or U4630 (N_4630,N_1393,N_1245);
xnor U4631 (N_4631,N_15,N_1156);
or U4632 (N_4632,N_846,N_2344);
nand U4633 (N_4633,N_336,N_1951);
nor U4634 (N_4634,N_672,N_2208);
nand U4635 (N_4635,N_1450,N_1419);
and U4636 (N_4636,N_894,N_1230);
nand U4637 (N_4637,N_1582,N_800);
or U4638 (N_4638,N_360,N_306);
nor U4639 (N_4639,N_1420,N_1069);
or U4640 (N_4640,N_2444,N_2197);
and U4641 (N_4641,N_1120,N_388);
and U4642 (N_4642,N_1670,N_1514);
nand U4643 (N_4643,N_2023,N_2340);
and U4644 (N_4644,N_1981,N_1067);
and U4645 (N_4645,N_747,N_1003);
or U4646 (N_4646,N_2439,N_251);
and U4647 (N_4647,N_2479,N_245);
nor U4648 (N_4648,N_2024,N_1332);
and U4649 (N_4649,N_2080,N_1591);
or U4650 (N_4650,N_1132,N_1211);
and U4651 (N_4651,N_2358,N_2234);
nand U4652 (N_4652,N_82,N_1695);
nor U4653 (N_4653,N_221,N_145);
and U4654 (N_4654,N_2382,N_368);
nor U4655 (N_4655,N_1894,N_1374);
or U4656 (N_4656,N_1424,N_192);
nand U4657 (N_4657,N_1238,N_1273);
nor U4658 (N_4658,N_965,N_824);
or U4659 (N_4659,N_1432,N_398);
xnor U4660 (N_4660,N_2293,N_1160);
nand U4661 (N_4661,N_289,N_2257);
nand U4662 (N_4662,N_2298,N_1605);
or U4663 (N_4663,N_38,N_585);
or U4664 (N_4664,N_1834,N_1970);
nor U4665 (N_4665,N_67,N_1657);
xor U4666 (N_4666,N_443,N_2154);
or U4667 (N_4667,N_2011,N_705);
nor U4668 (N_4668,N_1327,N_1355);
and U4669 (N_4669,N_172,N_318);
nor U4670 (N_4670,N_1436,N_267);
and U4671 (N_4671,N_917,N_1450);
xnor U4672 (N_4672,N_222,N_2197);
nor U4673 (N_4673,N_378,N_2130);
xnor U4674 (N_4674,N_285,N_598);
nor U4675 (N_4675,N_2217,N_2475);
nor U4676 (N_4676,N_2229,N_2014);
xnor U4677 (N_4677,N_2375,N_1962);
and U4678 (N_4678,N_221,N_1604);
xor U4679 (N_4679,N_2199,N_323);
and U4680 (N_4680,N_1476,N_1617);
or U4681 (N_4681,N_1633,N_918);
xor U4682 (N_4682,N_56,N_65);
nor U4683 (N_4683,N_1461,N_503);
or U4684 (N_4684,N_165,N_1651);
nor U4685 (N_4685,N_2080,N_689);
nand U4686 (N_4686,N_2366,N_664);
nand U4687 (N_4687,N_1647,N_409);
or U4688 (N_4688,N_1116,N_4);
nor U4689 (N_4689,N_548,N_1807);
nand U4690 (N_4690,N_732,N_2283);
nor U4691 (N_4691,N_1200,N_122);
xnor U4692 (N_4692,N_1498,N_939);
or U4693 (N_4693,N_466,N_1756);
xnor U4694 (N_4694,N_536,N_1210);
nand U4695 (N_4695,N_392,N_2271);
xnor U4696 (N_4696,N_143,N_2459);
nand U4697 (N_4697,N_1623,N_1970);
or U4698 (N_4698,N_1175,N_2199);
or U4699 (N_4699,N_2102,N_226);
or U4700 (N_4700,N_2453,N_2245);
nor U4701 (N_4701,N_830,N_1212);
and U4702 (N_4702,N_290,N_2166);
nor U4703 (N_4703,N_46,N_1893);
nor U4704 (N_4704,N_946,N_1963);
nand U4705 (N_4705,N_1305,N_680);
nor U4706 (N_4706,N_1555,N_508);
xnor U4707 (N_4707,N_1166,N_1562);
nor U4708 (N_4708,N_874,N_248);
nor U4709 (N_4709,N_1679,N_1040);
and U4710 (N_4710,N_284,N_1710);
nor U4711 (N_4711,N_2229,N_1432);
and U4712 (N_4712,N_1740,N_570);
xor U4713 (N_4713,N_204,N_367);
nor U4714 (N_4714,N_2388,N_2007);
and U4715 (N_4715,N_1664,N_665);
and U4716 (N_4716,N_995,N_1366);
nand U4717 (N_4717,N_350,N_2476);
nor U4718 (N_4718,N_818,N_185);
and U4719 (N_4719,N_1403,N_38);
or U4720 (N_4720,N_920,N_219);
or U4721 (N_4721,N_2174,N_2078);
or U4722 (N_4722,N_31,N_2440);
xnor U4723 (N_4723,N_1461,N_1974);
nor U4724 (N_4724,N_971,N_133);
nand U4725 (N_4725,N_1583,N_122);
nand U4726 (N_4726,N_2323,N_547);
nand U4727 (N_4727,N_1092,N_723);
and U4728 (N_4728,N_1232,N_290);
nor U4729 (N_4729,N_2010,N_2095);
nor U4730 (N_4730,N_1344,N_1917);
nor U4731 (N_4731,N_881,N_2460);
xnor U4732 (N_4732,N_395,N_1109);
and U4733 (N_4733,N_786,N_2338);
and U4734 (N_4734,N_2470,N_1623);
or U4735 (N_4735,N_1541,N_1129);
nor U4736 (N_4736,N_1293,N_352);
nand U4737 (N_4737,N_1955,N_445);
nor U4738 (N_4738,N_887,N_1860);
and U4739 (N_4739,N_813,N_457);
xor U4740 (N_4740,N_2187,N_2310);
or U4741 (N_4741,N_2340,N_2326);
or U4742 (N_4742,N_2474,N_1692);
xnor U4743 (N_4743,N_383,N_1757);
or U4744 (N_4744,N_437,N_1854);
nor U4745 (N_4745,N_1266,N_659);
nor U4746 (N_4746,N_1281,N_542);
or U4747 (N_4747,N_841,N_1326);
nand U4748 (N_4748,N_1682,N_59);
or U4749 (N_4749,N_228,N_339);
and U4750 (N_4750,N_1111,N_557);
or U4751 (N_4751,N_1626,N_1009);
nand U4752 (N_4752,N_1592,N_2313);
nor U4753 (N_4753,N_2347,N_1718);
nor U4754 (N_4754,N_1397,N_997);
nor U4755 (N_4755,N_1655,N_2384);
nor U4756 (N_4756,N_223,N_457);
nand U4757 (N_4757,N_46,N_1762);
and U4758 (N_4758,N_231,N_156);
or U4759 (N_4759,N_920,N_1506);
nor U4760 (N_4760,N_290,N_2480);
nor U4761 (N_4761,N_1411,N_1108);
and U4762 (N_4762,N_2218,N_1604);
xor U4763 (N_4763,N_1416,N_2177);
nand U4764 (N_4764,N_2286,N_1344);
nor U4765 (N_4765,N_784,N_1170);
nand U4766 (N_4766,N_573,N_895);
xor U4767 (N_4767,N_1254,N_2393);
or U4768 (N_4768,N_2371,N_1262);
and U4769 (N_4769,N_461,N_1770);
and U4770 (N_4770,N_982,N_531);
nor U4771 (N_4771,N_943,N_1494);
nand U4772 (N_4772,N_1145,N_1213);
or U4773 (N_4773,N_1402,N_510);
and U4774 (N_4774,N_2085,N_1908);
and U4775 (N_4775,N_1215,N_947);
or U4776 (N_4776,N_1664,N_599);
and U4777 (N_4777,N_1378,N_1092);
and U4778 (N_4778,N_2436,N_684);
xor U4779 (N_4779,N_1316,N_2191);
nor U4780 (N_4780,N_1353,N_575);
and U4781 (N_4781,N_882,N_2060);
nor U4782 (N_4782,N_1047,N_741);
or U4783 (N_4783,N_1870,N_578);
nor U4784 (N_4784,N_1834,N_671);
nand U4785 (N_4785,N_2372,N_711);
and U4786 (N_4786,N_514,N_2458);
nand U4787 (N_4787,N_171,N_1197);
and U4788 (N_4788,N_415,N_1569);
nand U4789 (N_4789,N_1976,N_1903);
nor U4790 (N_4790,N_823,N_463);
and U4791 (N_4791,N_420,N_1579);
nor U4792 (N_4792,N_930,N_1854);
nand U4793 (N_4793,N_716,N_2374);
xor U4794 (N_4794,N_2298,N_2312);
xor U4795 (N_4795,N_1147,N_832);
and U4796 (N_4796,N_266,N_2150);
or U4797 (N_4797,N_2140,N_177);
or U4798 (N_4798,N_1493,N_840);
and U4799 (N_4799,N_1091,N_369);
nand U4800 (N_4800,N_255,N_939);
or U4801 (N_4801,N_1897,N_2173);
xnor U4802 (N_4802,N_1588,N_455);
xnor U4803 (N_4803,N_923,N_1278);
nand U4804 (N_4804,N_826,N_1079);
nand U4805 (N_4805,N_172,N_152);
nand U4806 (N_4806,N_1731,N_2272);
or U4807 (N_4807,N_59,N_691);
or U4808 (N_4808,N_1204,N_1538);
or U4809 (N_4809,N_1706,N_2255);
or U4810 (N_4810,N_851,N_266);
xnor U4811 (N_4811,N_1421,N_1160);
nor U4812 (N_4812,N_1051,N_1292);
and U4813 (N_4813,N_2220,N_1297);
xnor U4814 (N_4814,N_869,N_539);
or U4815 (N_4815,N_1265,N_871);
nand U4816 (N_4816,N_1520,N_1917);
and U4817 (N_4817,N_726,N_1239);
nor U4818 (N_4818,N_1148,N_1222);
or U4819 (N_4819,N_1081,N_1857);
nor U4820 (N_4820,N_513,N_2493);
xnor U4821 (N_4821,N_680,N_1466);
or U4822 (N_4822,N_397,N_1478);
and U4823 (N_4823,N_1754,N_1721);
or U4824 (N_4824,N_1111,N_294);
or U4825 (N_4825,N_794,N_954);
nand U4826 (N_4826,N_2061,N_1141);
or U4827 (N_4827,N_2180,N_689);
and U4828 (N_4828,N_1858,N_52);
nor U4829 (N_4829,N_434,N_2209);
and U4830 (N_4830,N_265,N_1785);
or U4831 (N_4831,N_1873,N_1638);
and U4832 (N_4832,N_1702,N_1291);
nor U4833 (N_4833,N_1096,N_1330);
or U4834 (N_4834,N_1486,N_401);
xor U4835 (N_4835,N_189,N_2476);
or U4836 (N_4836,N_653,N_67);
and U4837 (N_4837,N_1963,N_353);
or U4838 (N_4838,N_100,N_309);
and U4839 (N_4839,N_482,N_791);
or U4840 (N_4840,N_1138,N_309);
nand U4841 (N_4841,N_1947,N_2091);
and U4842 (N_4842,N_313,N_337);
or U4843 (N_4843,N_102,N_2449);
and U4844 (N_4844,N_1329,N_2005);
or U4845 (N_4845,N_1595,N_2315);
nor U4846 (N_4846,N_1425,N_2051);
and U4847 (N_4847,N_1658,N_1508);
and U4848 (N_4848,N_1844,N_1933);
nand U4849 (N_4849,N_2114,N_1022);
or U4850 (N_4850,N_113,N_115);
xnor U4851 (N_4851,N_1366,N_1385);
xnor U4852 (N_4852,N_2235,N_2037);
or U4853 (N_4853,N_609,N_425);
and U4854 (N_4854,N_1860,N_1951);
xor U4855 (N_4855,N_607,N_429);
nor U4856 (N_4856,N_1201,N_971);
or U4857 (N_4857,N_2074,N_1954);
xor U4858 (N_4858,N_2044,N_1811);
nor U4859 (N_4859,N_2115,N_1523);
and U4860 (N_4860,N_1793,N_1406);
and U4861 (N_4861,N_2298,N_235);
xor U4862 (N_4862,N_1952,N_874);
xnor U4863 (N_4863,N_1572,N_734);
or U4864 (N_4864,N_959,N_2071);
nor U4865 (N_4865,N_962,N_1371);
nor U4866 (N_4866,N_10,N_1285);
or U4867 (N_4867,N_1363,N_157);
and U4868 (N_4868,N_765,N_2337);
nor U4869 (N_4869,N_1023,N_2171);
nor U4870 (N_4870,N_112,N_1269);
nor U4871 (N_4871,N_1760,N_1473);
nand U4872 (N_4872,N_2425,N_173);
and U4873 (N_4873,N_1972,N_456);
xor U4874 (N_4874,N_1232,N_371);
xor U4875 (N_4875,N_12,N_1967);
nor U4876 (N_4876,N_1626,N_2328);
xor U4877 (N_4877,N_212,N_536);
nor U4878 (N_4878,N_1276,N_1935);
xnor U4879 (N_4879,N_2213,N_2360);
xor U4880 (N_4880,N_1224,N_1928);
and U4881 (N_4881,N_904,N_2348);
xor U4882 (N_4882,N_1348,N_1176);
or U4883 (N_4883,N_1986,N_253);
and U4884 (N_4884,N_2328,N_2321);
and U4885 (N_4885,N_1624,N_48);
xnor U4886 (N_4886,N_2307,N_360);
xor U4887 (N_4887,N_1153,N_375);
nor U4888 (N_4888,N_1064,N_2466);
nor U4889 (N_4889,N_603,N_1297);
and U4890 (N_4890,N_679,N_1287);
xnor U4891 (N_4891,N_2495,N_993);
xor U4892 (N_4892,N_253,N_625);
xnor U4893 (N_4893,N_943,N_1334);
or U4894 (N_4894,N_1294,N_608);
nand U4895 (N_4895,N_1304,N_2420);
and U4896 (N_4896,N_1883,N_827);
xnor U4897 (N_4897,N_2040,N_1296);
and U4898 (N_4898,N_2361,N_969);
xnor U4899 (N_4899,N_1344,N_495);
and U4900 (N_4900,N_713,N_247);
or U4901 (N_4901,N_2461,N_475);
nand U4902 (N_4902,N_148,N_938);
nand U4903 (N_4903,N_2211,N_149);
nor U4904 (N_4904,N_1020,N_2062);
and U4905 (N_4905,N_1306,N_699);
xnor U4906 (N_4906,N_550,N_1894);
or U4907 (N_4907,N_2495,N_1429);
or U4908 (N_4908,N_1753,N_522);
nand U4909 (N_4909,N_1022,N_1589);
xnor U4910 (N_4910,N_1904,N_63);
nand U4911 (N_4911,N_1772,N_2149);
or U4912 (N_4912,N_622,N_337);
xor U4913 (N_4913,N_1123,N_2457);
xnor U4914 (N_4914,N_582,N_780);
nor U4915 (N_4915,N_15,N_484);
or U4916 (N_4916,N_2205,N_2142);
nand U4917 (N_4917,N_529,N_2361);
nor U4918 (N_4918,N_803,N_1417);
and U4919 (N_4919,N_656,N_2078);
nor U4920 (N_4920,N_2047,N_818);
and U4921 (N_4921,N_114,N_907);
nor U4922 (N_4922,N_808,N_876);
nand U4923 (N_4923,N_896,N_326);
xnor U4924 (N_4924,N_2271,N_1276);
nand U4925 (N_4925,N_164,N_1263);
and U4926 (N_4926,N_1607,N_828);
nor U4927 (N_4927,N_1592,N_466);
nand U4928 (N_4928,N_1690,N_1404);
xnor U4929 (N_4929,N_2308,N_213);
and U4930 (N_4930,N_1814,N_1918);
or U4931 (N_4931,N_2243,N_642);
nor U4932 (N_4932,N_526,N_455);
xor U4933 (N_4933,N_1441,N_640);
or U4934 (N_4934,N_285,N_2450);
xor U4935 (N_4935,N_1516,N_2038);
nand U4936 (N_4936,N_1254,N_1182);
and U4937 (N_4937,N_237,N_340);
xnor U4938 (N_4938,N_1157,N_39);
or U4939 (N_4939,N_966,N_1267);
or U4940 (N_4940,N_508,N_481);
xor U4941 (N_4941,N_640,N_1899);
or U4942 (N_4942,N_684,N_1193);
or U4943 (N_4943,N_2494,N_1480);
nor U4944 (N_4944,N_683,N_475);
or U4945 (N_4945,N_1317,N_1087);
nand U4946 (N_4946,N_428,N_510);
or U4947 (N_4947,N_132,N_1953);
nand U4948 (N_4948,N_113,N_1343);
xnor U4949 (N_4949,N_1588,N_2280);
nand U4950 (N_4950,N_1728,N_2310);
or U4951 (N_4951,N_1889,N_402);
xor U4952 (N_4952,N_1715,N_1528);
or U4953 (N_4953,N_505,N_2207);
nand U4954 (N_4954,N_2004,N_1283);
or U4955 (N_4955,N_639,N_785);
or U4956 (N_4956,N_2167,N_1381);
nand U4957 (N_4957,N_944,N_1144);
or U4958 (N_4958,N_905,N_66);
or U4959 (N_4959,N_742,N_968);
nor U4960 (N_4960,N_2366,N_2129);
or U4961 (N_4961,N_675,N_570);
nor U4962 (N_4962,N_529,N_1887);
or U4963 (N_4963,N_343,N_64);
nand U4964 (N_4964,N_1896,N_278);
nor U4965 (N_4965,N_1129,N_1783);
or U4966 (N_4966,N_826,N_69);
nor U4967 (N_4967,N_927,N_108);
or U4968 (N_4968,N_1607,N_1875);
nand U4969 (N_4969,N_1016,N_2281);
nor U4970 (N_4970,N_2149,N_1849);
nand U4971 (N_4971,N_306,N_69);
xor U4972 (N_4972,N_72,N_1843);
xor U4973 (N_4973,N_1267,N_619);
and U4974 (N_4974,N_2374,N_2326);
nand U4975 (N_4975,N_2333,N_869);
and U4976 (N_4976,N_56,N_1805);
and U4977 (N_4977,N_353,N_1439);
nor U4978 (N_4978,N_569,N_1241);
and U4979 (N_4979,N_1460,N_1976);
nand U4980 (N_4980,N_1194,N_470);
and U4981 (N_4981,N_995,N_137);
xnor U4982 (N_4982,N_1986,N_2227);
nor U4983 (N_4983,N_1391,N_1523);
xor U4984 (N_4984,N_1608,N_1820);
xnor U4985 (N_4985,N_898,N_1542);
nand U4986 (N_4986,N_2090,N_67);
or U4987 (N_4987,N_1964,N_490);
nand U4988 (N_4988,N_2476,N_1923);
nand U4989 (N_4989,N_1281,N_1270);
nand U4990 (N_4990,N_1862,N_330);
or U4991 (N_4991,N_1814,N_1738);
nor U4992 (N_4992,N_121,N_2259);
or U4993 (N_4993,N_2351,N_1483);
nand U4994 (N_4994,N_968,N_1634);
nor U4995 (N_4995,N_1136,N_2481);
or U4996 (N_4996,N_281,N_1925);
and U4997 (N_4997,N_65,N_912);
nor U4998 (N_4998,N_1695,N_1076);
xor U4999 (N_4999,N_1402,N_1085);
or U5000 (N_5000,N_2742,N_2836);
xnor U5001 (N_5001,N_4481,N_4350);
nor U5002 (N_5002,N_3315,N_4302);
xor U5003 (N_5003,N_3504,N_3835);
and U5004 (N_5004,N_2515,N_2745);
xor U5005 (N_5005,N_3673,N_4138);
or U5006 (N_5006,N_3245,N_3678);
nor U5007 (N_5007,N_4849,N_3507);
nor U5008 (N_5008,N_2577,N_3262);
or U5009 (N_5009,N_3544,N_4415);
nand U5010 (N_5010,N_4386,N_4485);
nand U5011 (N_5011,N_3374,N_3200);
and U5012 (N_5012,N_3923,N_3853);
xor U5013 (N_5013,N_3759,N_3751);
or U5014 (N_5014,N_2623,N_3893);
nor U5015 (N_5015,N_2739,N_4439);
nor U5016 (N_5016,N_2806,N_4269);
and U5017 (N_5017,N_4100,N_4846);
xor U5018 (N_5018,N_4772,N_4999);
nor U5019 (N_5019,N_3359,N_4600);
xnor U5020 (N_5020,N_3159,N_2644);
or U5021 (N_5021,N_4303,N_4002);
nor U5022 (N_5022,N_2611,N_4933);
nor U5023 (N_5023,N_4437,N_3513);
xnor U5024 (N_5024,N_2821,N_4893);
and U5025 (N_5025,N_2951,N_4165);
xnor U5026 (N_5026,N_3945,N_3051);
and U5027 (N_5027,N_4839,N_2506);
nor U5028 (N_5028,N_3278,N_2677);
xor U5029 (N_5029,N_4878,N_3270);
or U5030 (N_5030,N_4831,N_4022);
nand U5031 (N_5031,N_4382,N_3367);
xor U5032 (N_5032,N_4595,N_4273);
xor U5033 (N_5033,N_3495,N_4234);
xor U5034 (N_5034,N_4363,N_4869);
xnor U5035 (N_5035,N_2659,N_4690);
nor U5036 (N_5036,N_3439,N_3774);
and U5037 (N_5037,N_3994,N_4913);
xnor U5038 (N_5038,N_2561,N_2875);
and U5039 (N_5039,N_3191,N_3968);
or U5040 (N_5040,N_4498,N_2798);
nor U5041 (N_5041,N_4187,N_4209);
and U5042 (N_5042,N_3209,N_4291);
xor U5043 (N_5043,N_4531,N_3559);
nand U5044 (N_5044,N_4333,N_2637);
xor U5045 (N_5045,N_3413,N_3955);
xor U5046 (N_5046,N_3466,N_4671);
and U5047 (N_5047,N_2887,N_3970);
or U5048 (N_5048,N_3587,N_3857);
nor U5049 (N_5049,N_3060,N_2549);
nand U5050 (N_5050,N_2691,N_3907);
or U5051 (N_5051,N_2928,N_3908);
and U5052 (N_5052,N_4254,N_4072);
nand U5053 (N_5053,N_3609,N_4031);
xnor U5054 (N_5054,N_2630,N_3233);
or U5055 (N_5055,N_4293,N_2733);
nand U5056 (N_5056,N_4385,N_3280);
nor U5057 (N_5057,N_2993,N_2926);
nor U5058 (N_5058,N_3383,N_3515);
and U5059 (N_5059,N_3824,N_3497);
and U5060 (N_5060,N_2564,N_2930);
or U5061 (N_5061,N_3025,N_4968);
xnor U5062 (N_5062,N_3873,N_3339);
and U5063 (N_5063,N_2729,N_3640);
or U5064 (N_5064,N_2925,N_4570);
nand U5065 (N_5065,N_4155,N_3172);
and U5066 (N_5066,N_4411,N_4397);
nor U5067 (N_5067,N_4802,N_3127);
nor U5068 (N_5068,N_3210,N_2563);
or U5069 (N_5069,N_4368,N_3643);
xnor U5070 (N_5070,N_3176,N_3454);
and U5071 (N_5071,N_4815,N_3808);
and U5072 (N_5072,N_4680,N_4109);
and U5073 (N_5073,N_3114,N_3900);
nand U5074 (N_5074,N_2958,N_3153);
xnor U5075 (N_5075,N_4745,N_2698);
and U5076 (N_5076,N_2957,N_3805);
nor U5077 (N_5077,N_4722,N_4843);
nor U5078 (N_5078,N_4617,N_4612);
or U5079 (N_5079,N_3899,N_3163);
nor U5080 (N_5080,N_2812,N_4230);
xnor U5081 (N_5081,N_3211,N_4080);
nand U5082 (N_5082,N_4715,N_3676);
or U5083 (N_5083,N_3485,N_2852);
nand U5084 (N_5084,N_3097,N_4227);
nor U5085 (N_5085,N_3498,N_3998);
nor U5086 (N_5086,N_2789,N_4013);
and U5087 (N_5087,N_4300,N_3831);
nand U5088 (N_5088,N_3425,N_3343);
xnor U5089 (N_5089,N_2913,N_4925);
and U5090 (N_5090,N_3294,N_2646);
nor U5091 (N_5091,N_3275,N_2710);
nand U5092 (N_5092,N_3380,N_3796);
nor U5093 (N_5093,N_3412,N_3442);
nand U5094 (N_5094,N_3563,N_2971);
nor U5095 (N_5095,N_2676,N_2790);
nand U5096 (N_5096,N_3251,N_3444);
and U5097 (N_5097,N_4009,N_3479);
nor U5098 (N_5098,N_4006,N_2865);
nand U5099 (N_5099,N_3397,N_2603);
and U5100 (N_5100,N_2936,N_2756);
xor U5101 (N_5101,N_4692,N_3880);
xnor U5102 (N_5102,N_3946,N_4391);
xnor U5103 (N_5103,N_4944,N_4226);
and U5104 (N_5104,N_3224,N_4725);
nor U5105 (N_5105,N_3776,N_4463);
nor U5106 (N_5106,N_3128,N_4988);
and U5107 (N_5107,N_4528,N_3866);
nand U5108 (N_5108,N_3166,N_3287);
and U5109 (N_5109,N_2979,N_3576);
nor U5110 (N_5110,N_3213,N_3897);
xnor U5111 (N_5111,N_3617,N_4643);
xnor U5112 (N_5112,N_3811,N_2586);
or U5113 (N_5113,N_4267,N_3373);
nand U5114 (N_5114,N_3874,N_2560);
nand U5115 (N_5115,N_2902,N_3394);
xnor U5116 (N_5116,N_2767,N_4535);
and U5117 (N_5117,N_2638,N_4036);
nor U5118 (N_5118,N_2885,N_4129);
xor U5119 (N_5119,N_4532,N_3292);
nand U5120 (N_5120,N_2805,N_3615);
nor U5121 (N_5121,N_3445,N_4395);
nor U5122 (N_5122,N_4121,N_2660);
nand U5123 (N_5123,N_4844,N_4568);
nand U5124 (N_5124,N_4794,N_4214);
nand U5125 (N_5125,N_2968,N_3016);
and U5126 (N_5126,N_3989,N_3987);
nand U5127 (N_5127,N_2932,N_3732);
nand U5128 (N_5128,N_4076,N_3117);
xnor U5129 (N_5129,N_2788,N_3288);
nand U5130 (N_5130,N_3584,N_4943);
or U5131 (N_5131,N_4879,N_3596);
or U5132 (N_5132,N_4963,N_4610);
nand U5133 (N_5133,N_4343,N_4171);
nand U5134 (N_5134,N_2690,N_2686);
nand U5135 (N_5135,N_3271,N_3652);
nand U5136 (N_5136,N_4655,N_3942);
nand U5137 (N_5137,N_4496,N_2682);
or U5138 (N_5138,N_2656,N_3856);
xnor U5139 (N_5139,N_4635,N_2544);
nand U5140 (N_5140,N_4270,N_4593);
xnor U5141 (N_5141,N_4818,N_2622);
xor U5142 (N_5142,N_2599,N_4200);
xnor U5143 (N_5143,N_3341,N_4663);
or U5144 (N_5144,N_2948,N_3527);
nor U5145 (N_5145,N_2985,N_3736);
nand U5146 (N_5146,N_3250,N_2769);
xnor U5147 (N_5147,N_3407,N_2662);
nor U5148 (N_5148,N_3591,N_4912);
or U5149 (N_5149,N_4704,N_3142);
or U5150 (N_5150,N_2990,N_2940);
and U5151 (N_5151,N_3557,N_4452);
xnor U5152 (N_5152,N_4266,N_3523);
xor U5153 (N_5153,N_4618,N_4057);
nand U5154 (N_5154,N_3928,N_4323);
nor U5155 (N_5155,N_2912,N_4140);
or U5156 (N_5156,N_2719,N_3937);
and U5157 (N_5157,N_4739,N_3168);
and U5158 (N_5158,N_2956,N_4661);
and U5159 (N_5159,N_2681,N_4317);
and U5160 (N_5160,N_4744,N_3846);
nor U5161 (N_5161,N_4465,N_3252);
nor U5162 (N_5162,N_4901,N_4763);
or U5163 (N_5163,N_3565,N_3305);
or U5164 (N_5164,N_3657,N_3129);
or U5165 (N_5165,N_3603,N_3653);
or U5166 (N_5166,N_4734,N_3954);
and U5167 (N_5167,N_4630,N_2614);
nor U5168 (N_5168,N_2640,N_4938);
or U5169 (N_5169,N_3423,N_3944);
nand U5170 (N_5170,N_3951,N_3966);
nor U5171 (N_5171,N_3530,N_2752);
nor U5172 (N_5172,N_3018,N_2896);
nand U5173 (N_5173,N_3849,N_3369);
and U5174 (N_5174,N_4217,N_4244);
xor U5175 (N_5175,N_3671,N_2914);
xnor U5176 (N_5176,N_2541,N_4945);
xnor U5177 (N_5177,N_3253,N_3242);
xnor U5178 (N_5178,N_3405,N_2813);
and U5179 (N_5179,N_2619,N_3722);
nand U5180 (N_5180,N_2987,N_4037);
nand U5181 (N_5181,N_4365,N_3894);
or U5182 (N_5182,N_4807,N_4039);
or U5183 (N_5183,N_3206,N_3030);
or U5184 (N_5184,N_2618,N_4426);
and U5185 (N_5185,N_3660,N_4873);
xnor U5186 (N_5186,N_3589,N_4880);
nor U5187 (N_5187,N_4128,N_3758);
nand U5188 (N_5188,N_4205,N_3094);
nor U5189 (N_5189,N_4297,N_2744);
xor U5190 (N_5190,N_3139,N_2811);
nor U5191 (N_5191,N_4554,N_4978);
nand U5192 (N_5192,N_4045,N_3500);
nor U5193 (N_5193,N_3223,N_3570);
or U5194 (N_5194,N_2859,N_3199);
nor U5195 (N_5195,N_3600,N_4316);
or U5196 (N_5196,N_3308,N_3698);
or U5197 (N_5197,N_4709,N_3834);
nor U5198 (N_5198,N_4942,N_4832);
xnor U5199 (N_5199,N_2799,N_3302);
or U5200 (N_5200,N_4821,N_3791);
nand U5201 (N_5201,N_4918,N_3043);
xnor U5202 (N_5202,N_4579,N_3022);
xnor U5203 (N_5203,N_3529,N_4969);
and U5204 (N_5204,N_4399,N_3586);
nor U5205 (N_5205,N_3289,N_3099);
nor U5206 (N_5206,N_3408,N_4202);
nor U5207 (N_5207,N_3389,N_4971);
nor U5208 (N_5208,N_2553,N_4759);
nor U5209 (N_5209,N_4791,N_3390);
and U5210 (N_5210,N_4688,N_4823);
nand U5211 (N_5211,N_3110,N_3474);
nor U5212 (N_5212,N_4046,N_3183);
nor U5213 (N_5213,N_3642,N_3710);
nor U5214 (N_5214,N_4923,N_4207);
xnor U5215 (N_5215,N_4376,N_4471);
xnor U5216 (N_5216,N_2507,N_4338);
and U5217 (N_5217,N_4929,N_3912);
xor U5218 (N_5218,N_4814,N_3592);
nor U5219 (N_5219,N_3410,N_3649);
nand U5220 (N_5220,N_3685,N_3203);
nand U5221 (N_5221,N_3311,N_4433);
xnor U5222 (N_5222,N_3562,N_4594);
nor U5223 (N_5223,N_4352,N_3182);
nand U5224 (N_5224,N_2610,N_4985);
xor U5225 (N_5225,N_2703,N_4288);
or U5226 (N_5226,N_4626,N_2757);
nand U5227 (N_5227,N_3489,N_3066);
nand U5228 (N_5228,N_3990,N_3887);
xor U5229 (N_5229,N_3050,N_2701);
nor U5230 (N_5230,N_2702,N_4636);
and U5231 (N_5231,N_2959,N_3450);
nand U5232 (N_5232,N_2688,N_4907);
xor U5233 (N_5233,N_4049,N_3137);
and U5234 (N_5234,N_3606,N_4418);
nand U5235 (N_5235,N_4114,N_4872);
nor U5236 (N_5236,N_3962,N_4061);
and U5237 (N_5237,N_3622,N_3919);
nand U5238 (N_5238,N_3088,N_4224);
or U5239 (N_5239,N_4565,N_2751);
and U5240 (N_5240,N_4975,N_4694);
and U5241 (N_5241,N_2998,N_3391);
nand U5242 (N_5242,N_4665,N_2607);
xor U5243 (N_5243,N_4658,N_3612);
and U5244 (N_5244,N_3680,N_4569);
nor U5245 (N_5245,N_2888,N_3301);
xor U5246 (N_5246,N_3664,N_4909);
nor U5247 (N_5247,N_2548,N_2793);
or U5248 (N_5248,N_3169,N_4998);
nor U5249 (N_5249,N_4346,N_3334);
nand U5250 (N_5250,N_4522,N_4572);
xnor U5251 (N_5251,N_4356,N_3635);
or U5252 (N_5252,N_3859,N_4748);
nand U5253 (N_5253,N_3516,N_3136);
xor U5254 (N_5254,N_4474,N_2890);
nand U5255 (N_5255,N_3690,N_4774);
nor U5256 (N_5256,N_2886,N_3734);
and U5257 (N_5257,N_4125,N_2546);
nand U5258 (N_5258,N_2654,N_4713);
nand U5259 (N_5259,N_2641,N_2721);
nand U5260 (N_5260,N_3800,N_4870);
and U5261 (N_5261,N_4149,N_3038);
and U5262 (N_5262,N_4034,N_3692);
xnor U5263 (N_5263,N_2786,N_3167);
and U5264 (N_5264,N_4364,N_3468);
nor U5265 (N_5265,N_3478,N_4811);
xnor U5266 (N_5266,N_4592,N_3991);
nand U5267 (N_5267,N_3430,N_4897);
and U5268 (N_5268,N_4495,N_3514);
or U5269 (N_5269,N_4476,N_4615);
nand U5270 (N_5270,N_2804,N_4296);
and U5271 (N_5271,N_4074,N_3309);
or U5272 (N_5272,N_2608,N_2976);
nand U5273 (N_5273,N_2587,N_4351);
nand U5274 (N_5274,N_2725,N_2864);
and U5275 (N_5275,N_4597,N_3855);
xor U5276 (N_5276,N_3327,N_4740);
nor U5277 (N_5277,N_3451,N_4252);
nand U5278 (N_5278,N_2679,N_4856);
and U5279 (N_5279,N_2632,N_4706);
and U5280 (N_5280,N_3348,N_3215);
and U5281 (N_5281,N_4979,N_4687);
nor U5282 (N_5282,N_3668,N_3701);
and U5283 (N_5283,N_2601,N_4805);
nor U5284 (N_5284,N_4780,N_2685);
nand U5285 (N_5285,N_3027,N_4258);
nor U5286 (N_5286,N_3487,N_3464);
xnor U5287 (N_5287,N_3401,N_2901);
and U5288 (N_5288,N_3865,N_3971);
or U5289 (N_5289,N_2652,N_4097);
xnor U5290 (N_5290,N_2861,N_3350);
or U5291 (N_5291,N_4124,N_4429);
nand U5292 (N_5292,N_3845,N_4369);
nor U5293 (N_5293,N_4840,N_3786);
and U5294 (N_5294,N_4287,N_2689);
xnor U5295 (N_5295,N_3775,N_4871);
and U5296 (N_5296,N_3452,N_3618);
nand U5297 (N_5297,N_2770,N_4460);
nand U5298 (N_5298,N_4198,N_3669);
xnor U5299 (N_5299,N_2731,N_2715);
xnor U5300 (N_5300,N_4776,N_3357);
xor U5301 (N_5301,N_4512,N_2768);
and U5302 (N_5302,N_3074,N_2747);
and U5303 (N_5303,N_2938,N_3465);
nor U5304 (N_5304,N_4679,N_4102);
and U5305 (N_5305,N_3844,N_4141);
nor U5306 (N_5306,N_4054,N_4444);
nand U5307 (N_5307,N_4019,N_4403);
nand U5308 (N_5308,N_3627,N_3847);
or U5309 (N_5309,N_2916,N_4987);
nor U5310 (N_5310,N_4573,N_2700);
and U5311 (N_5311,N_3065,N_4885);
xor U5312 (N_5312,N_3716,N_3240);
and U5313 (N_5313,N_3696,N_3010);
and U5314 (N_5314,N_4084,N_3354);
xor U5315 (N_5315,N_4319,N_3816);
nor U5316 (N_5316,N_3230,N_3014);
nand U5317 (N_5317,N_4803,N_3982);
xor U5318 (N_5318,N_4221,N_4308);
and U5319 (N_5319,N_4070,N_4150);
xor U5320 (N_5320,N_3699,N_3614);
and U5321 (N_5321,N_3267,N_3143);
nor U5322 (N_5322,N_3693,N_2856);
and U5323 (N_5323,N_2754,N_2693);
or U5324 (N_5324,N_3554,N_2829);
and U5325 (N_5325,N_3475,N_4672);
nor U5326 (N_5326,N_3938,N_2919);
and U5327 (N_5327,N_4769,N_3019);
or U5328 (N_5328,N_2808,N_4179);
nand U5329 (N_5329,N_4854,N_2933);
or U5330 (N_5330,N_4746,N_3814);
nor U5331 (N_5331,N_3123,N_3798);
nand U5332 (N_5332,N_3870,N_4717);
nor U5333 (N_5333,N_4211,N_3007);
nand U5334 (N_5334,N_4459,N_4309);
xor U5335 (N_5335,N_3787,N_4265);
or U5336 (N_5336,N_4268,N_4766);
nand U5337 (N_5337,N_3891,N_4334);
and U5338 (N_5338,N_2697,N_3477);
or U5339 (N_5339,N_3682,N_4799);
xor U5340 (N_5340,N_3707,N_3871);
or U5341 (N_5341,N_2523,N_2514);
nor U5342 (N_5342,N_4223,N_2605);
xnor U5343 (N_5343,N_4700,N_2639);
or U5344 (N_5344,N_4174,N_4372);
xnor U5345 (N_5345,N_4208,N_3349);
and U5346 (N_5346,N_4147,N_4405);
and U5347 (N_5347,N_3882,N_4098);
and U5348 (N_5348,N_3783,N_4447);
nor U5349 (N_5349,N_4081,N_3534);
nand U5350 (N_5350,N_2532,N_3631);
nand U5351 (N_5351,N_4004,N_2962);
nand U5352 (N_5352,N_3598,N_4542);
and U5353 (N_5353,N_4176,N_2503);
nor U5354 (N_5354,N_4219,N_4957);
or U5355 (N_5355,N_3620,N_3906);
nor U5356 (N_5356,N_4540,N_2723);
xor U5357 (N_5357,N_3109,N_3216);
and U5358 (N_5358,N_3539,N_3039);
or U5359 (N_5359,N_4563,N_4282);
nor U5360 (N_5360,N_4062,N_3806);
or U5361 (N_5361,N_2991,N_2822);
and U5362 (N_5362,N_2807,N_4727);
xor U5363 (N_5363,N_3836,N_3009);
and U5364 (N_5364,N_2761,N_3306);
nor U5365 (N_5365,N_3769,N_3090);
nand U5366 (N_5366,N_3372,N_3636);
xnor U5367 (N_5367,N_3358,N_2785);
nor U5368 (N_5368,N_2955,N_2866);
nand U5369 (N_5369,N_3869,N_4065);
nand U5370 (N_5370,N_3089,N_3034);
or U5371 (N_5371,N_4862,N_4470);
and U5372 (N_5372,N_2802,N_3960);
nor U5373 (N_5373,N_3629,N_3731);
xnor U5374 (N_5374,N_4030,N_3608);
and U5375 (N_5375,N_3616,N_3428);
nand U5376 (N_5376,N_4035,N_3054);
or U5377 (N_5377,N_2997,N_4956);
nand U5378 (N_5378,N_4464,N_4261);
or U5379 (N_5379,N_4392,N_3611);
nor U5380 (N_5380,N_4702,N_3543);
or U5381 (N_5381,N_3102,N_2647);
nand U5382 (N_5382,N_4851,N_3188);
nor U5383 (N_5383,N_4161,N_4132);
nor U5384 (N_5384,N_4668,N_4043);
and U5385 (N_5385,N_2884,N_4172);
and U5386 (N_5386,N_3406,N_2550);
nor U5387 (N_5387,N_2722,N_2830);
or U5388 (N_5388,N_4591,N_4402);
nand U5389 (N_5389,N_3247,N_3469);
nor U5390 (N_5390,N_2571,N_2664);
and U5391 (N_5391,N_3307,N_4071);
or U5392 (N_5392,N_4624,N_4770);
nand U5393 (N_5393,N_3265,N_4083);
nand U5394 (N_5394,N_4075,N_2635);
nor U5395 (N_5395,N_4064,N_4167);
nor U5396 (N_5396,N_2661,N_3901);
xnor U5397 (N_5397,N_4277,N_4497);
or U5398 (N_5398,N_4197,N_4018);
xnor U5399 (N_5399,N_3402,N_3761);
and U5400 (N_5400,N_4755,N_3795);
nand U5401 (N_5401,N_4499,N_3093);
and U5402 (N_5402,N_2600,N_2848);
xor U5403 (N_5403,N_4456,N_4613);
nor U5404 (N_5404,N_4449,N_3839);
xor U5405 (N_5405,N_3863,N_4242);
nand U5406 (N_5406,N_4325,N_4530);
or U5407 (N_5407,N_4714,N_4432);
nand U5408 (N_5408,N_3750,N_2582);
and U5409 (N_5409,N_3967,N_4571);
xor U5410 (N_5410,N_4414,N_4358);
nand U5411 (N_5411,N_4934,N_4094);
or U5412 (N_5412,N_3936,N_2972);
xor U5413 (N_5413,N_2684,N_3197);
xnor U5414 (N_5414,N_2568,N_4785);
or U5415 (N_5415,N_3067,N_4162);
xnor U5416 (N_5416,N_4357,N_3910);
nor U5417 (N_5417,N_4513,N_4027);
and U5418 (N_5418,N_3322,N_3132);
and U5419 (N_5419,N_3953,N_4866);
and U5420 (N_5420,N_2512,N_2839);
xnor U5421 (N_5421,N_3850,N_3858);
and U5422 (N_5422,N_4504,N_3903);
nand U5423 (N_5423,N_3665,N_4848);
and U5424 (N_5424,N_3453,N_4603);
nor U5425 (N_5425,N_3319,N_3221);
nand U5426 (N_5426,N_2915,N_3675);
and U5427 (N_5427,N_4651,N_4000);
nand U5428 (N_5428,N_3386,N_3983);
nand U5429 (N_5429,N_4604,N_2595);
or U5430 (N_5430,N_3313,N_2778);
or U5431 (N_5431,N_3918,N_3145);
nor U5432 (N_5432,N_3473,N_3239);
xnor U5433 (N_5433,N_4322,N_4292);
xor U5434 (N_5434,N_4960,N_3104);
xor U5435 (N_5435,N_4231,N_3377);
xor U5436 (N_5436,N_2704,N_4586);
or U5437 (N_5437,N_3877,N_2565);
or U5438 (N_5438,N_3108,N_4516);
or U5439 (N_5439,N_4650,N_3610);
nor U5440 (N_5440,N_3630,N_4684);
and U5441 (N_5441,N_3916,N_4251);
nand U5442 (N_5442,N_3318,N_2773);
xor U5443 (N_5443,N_2783,N_3355);
or U5444 (N_5444,N_4890,N_4825);
and U5445 (N_5445,N_4646,N_3533);
nor U5446 (N_5446,N_2847,N_3830);
and U5447 (N_5447,N_3053,N_4367);
nand U5448 (N_5448,N_3493,N_3602);
or U5449 (N_5449,N_3291,N_2855);
or U5450 (N_5450,N_4331,N_3929);
nand U5451 (N_5451,N_3257,N_2537);
and U5452 (N_5452,N_3661,N_4020);
xor U5453 (N_5453,N_4777,N_3184);
nor U5454 (N_5454,N_3781,N_3162);
or U5455 (N_5455,N_4567,N_3148);
or U5456 (N_5456,N_4294,N_2837);
and U5457 (N_5457,N_3999,N_4339);
nor U5458 (N_5458,N_3152,N_3809);
and U5459 (N_5459,N_4099,N_4360);
and U5460 (N_5460,N_3555,N_3772);
or U5461 (N_5461,N_4115,N_4883);
or U5462 (N_5462,N_4991,N_3540);
nand U5463 (N_5463,N_3446,N_2777);
nand U5464 (N_5464,N_2892,N_4738);
or U5465 (N_5465,N_4666,N_3512);
xnor U5466 (N_5466,N_3532,N_4921);
and U5467 (N_5467,N_3235,N_3368);
or U5468 (N_5468,N_4067,N_4683);
nand U5469 (N_5469,N_3726,N_4492);
and U5470 (N_5470,N_3155,N_3645);
xnor U5471 (N_5471,N_3101,N_3330);
nand U5472 (N_5472,N_4253,N_2853);
nor U5473 (N_5473,N_3467,N_3185);
nor U5474 (N_5474,N_2909,N_3517);
xor U5475 (N_5475,N_4861,N_2621);
and U5476 (N_5476,N_2517,N_3757);
xor U5477 (N_5477,N_2509,N_2738);
xnor U5478 (N_5478,N_4246,N_3788);
and U5479 (N_5479,N_3496,N_3963);
or U5480 (N_5480,N_4550,N_3528);
xor U5481 (N_5481,N_3531,N_3626);
or U5482 (N_5482,N_3848,N_3040);
xnor U5483 (N_5483,N_4574,N_3655);
nor U5484 (N_5484,N_3773,N_3822);
nor U5485 (N_5485,N_4750,N_4577);
nand U5486 (N_5486,N_4935,N_3069);
xor U5487 (N_5487,N_3713,N_4274);
nor U5488 (N_5488,N_4410,N_4424);
and U5489 (N_5489,N_4324,N_3161);
or U5490 (N_5490,N_4381,N_3739);
or U5491 (N_5491,N_3058,N_2883);
nand U5492 (N_5492,N_2960,N_3896);
nor U5493 (N_5493,N_2917,N_4157);
and U5494 (N_5494,N_3552,N_2889);
xor U5495 (N_5495,N_4536,N_2502);
xor U5496 (N_5496,N_3098,N_3258);
or U5497 (N_5497,N_3650,N_3956);
or U5498 (N_5498,N_4089,N_2727);
and U5499 (N_5499,N_4290,N_2593);
xor U5500 (N_5500,N_3457,N_2743);
nand U5501 (N_5501,N_4373,N_4517);
or U5502 (N_5502,N_2570,N_4491);
or U5503 (N_5503,N_3792,N_2764);
nand U5504 (N_5504,N_3285,N_4733);
xor U5505 (N_5505,N_2653,N_4606);
nand U5506 (N_5506,N_4557,N_4900);
or U5507 (N_5507,N_2562,N_2583);
xor U5508 (N_5508,N_3599,N_2575);
and U5509 (N_5509,N_3208,N_3006);
and U5510 (N_5510,N_3861,N_3421);
nand U5511 (N_5511,N_4250,N_4436);
xnor U5512 (N_5512,N_3441,N_4916);
nor U5513 (N_5513,N_4078,N_2657);
nor U5514 (N_5514,N_3363,N_3597);
or U5515 (N_5515,N_3116,N_3566);
nand U5516 (N_5516,N_3949,N_4473);
xnor U5517 (N_5517,N_3337,N_3674);
or U5518 (N_5518,N_3977,N_3976);
and U5519 (N_5519,N_4068,N_2740);
xnor U5520 (N_5520,N_4503,N_4335);
or U5521 (N_5521,N_3904,N_3965);
nor U5522 (N_5522,N_4272,N_3826);
xnor U5523 (N_5523,N_4556,N_3973);
nor U5524 (N_5524,N_4249,N_4857);
nor U5525 (N_5525,N_4620,N_4438);
xnor U5526 (N_5526,N_2629,N_3813);
or U5527 (N_5527,N_4298,N_3393);
nand U5528 (N_5528,N_4301,N_3249);
xor U5529 (N_5529,N_4884,N_3304);
nand U5530 (N_5530,N_2881,N_2774);
nand U5531 (N_5531,N_4581,N_2921);
or U5532 (N_5532,N_3458,N_4012);
and U5533 (N_5533,N_3324,N_4675);
and U5534 (N_5534,N_3841,N_4631);
or U5535 (N_5535,N_3958,N_2908);
and U5536 (N_5536,N_4344,N_4629);
and U5537 (N_5537,N_3141,N_2964);
or U5538 (N_5538,N_4218,N_3422);
or U5539 (N_5539,N_3243,N_2590);
and U5540 (N_5540,N_2649,N_4326);
xor U5541 (N_5541,N_2678,N_2809);
or U5542 (N_5542,N_3794,N_4674);
and U5543 (N_5543,N_2540,N_3062);
and U5544 (N_5544,N_4017,N_3248);
nand U5545 (N_5545,N_3911,N_2900);
nor U5546 (N_5546,N_2787,N_4511);
nand U5547 (N_5547,N_4789,N_4887);
or U5548 (N_5548,N_4657,N_4056);
or U5549 (N_5549,N_2597,N_2555);
and U5550 (N_5550,N_3714,N_3071);
xnor U5551 (N_5551,N_3020,N_4116);
xor U5552 (N_5552,N_2992,N_4166);
xnor U5553 (N_5553,N_3659,N_4833);
nor U5554 (N_5554,N_3825,N_4228);
or U5555 (N_5555,N_2999,N_3174);
xor U5556 (N_5556,N_4307,N_4984);
nor U5557 (N_5557,N_3864,N_3480);
nor U5558 (N_5558,N_4448,N_4091);
nand U5559 (N_5559,N_4553,N_2927);
nand U5560 (N_5560,N_3332,N_2937);
xor U5561 (N_5561,N_3063,N_4723);
nor U5562 (N_5562,N_4962,N_4086);
or U5563 (N_5563,N_3588,N_4201);
nor U5564 (N_5564,N_3579,N_4007);
nor U5565 (N_5565,N_4830,N_4705);
nand U5566 (N_5566,N_4989,N_4278);
nand U5567 (N_5567,N_4434,N_4525);
or U5568 (N_5568,N_2573,N_4137);
and U5569 (N_5569,N_4678,N_2734);
and U5570 (N_5570,N_3100,N_4010);
or U5571 (N_5571,N_4954,N_3447);
or U5572 (N_5572,N_4183,N_2531);
xor U5573 (N_5573,N_3684,N_4611);
xnor U5574 (N_5574,N_4173,N_4152);
nor U5575 (N_5575,N_3745,N_2850);
nor U5576 (N_5576,N_2862,N_2530);
or U5577 (N_5577,N_3688,N_4412);
nor U5578 (N_5578,N_4315,N_4669);
xnor U5579 (N_5579,N_4732,N_3506);
nor U5580 (N_5580,N_4271,N_3961);
or U5581 (N_5581,N_4716,N_4256);
and U5582 (N_5582,N_4820,N_3264);
nor U5583 (N_5583,N_2772,N_4451);
nand U5584 (N_5584,N_2935,N_3472);
or U5585 (N_5585,N_3765,N_4028);
and U5586 (N_5586,N_3234,N_3028);
or U5587 (N_5587,N_4764,N_4685);
xor U5588 (N_5588,N_4127,N_3077);
nand U5589 (N_5589,N_4151,N_4106);
nand U5590 (N_5590,N_3205,N_4387);
nand U5591 (N_5591,N_4865,N_2663);
and U5592 (N_5592,N_4941,N_3689);
or U5593 (N_5593,N_4107,N_3178);
nor U5594 (N_5594,N_2670,N_2818);
nand U5595 (N_5595,N_3399,N_2929);
and U5596 (N_5596,N_4730,N_2834);
or U5597 (N_5597,N_4383,N_3733);
nand U5598 (N_5598,N_3201,N_4859);
and U5599 (N_5599,N_3677,N_3255);
and U5600 (N_5600,N_4995,N_3420);
or U5601 (N_5601,N_4765,N_3819);
or U5602 (N_5602,N_4564,N_2795);
xor U5603 (N_5603,N_2920,N_4354);
xnor U5604 (N_5604,N_2980,N_3719);
nand U5605 (N_5605,N_3842,N_4838);
xor U5606 (N_5606,N_2882,N_4523);
xor U5607 (N_5607,N_4509,N_2878);
and U5608 (N_5608,N_3639,N_3491);
nand U5609 (N_5609,N_4576,N_2762);
nand U5610 (N_5610,N_4038,N_4144);
and U5611 (N_5611,N_2714,N_4953);
nand U5612 (N_5612,N_4640,N_4394);
and U5613 (N_5613,N_4195,N_4313);
nand U5614 (N_5614,N_4264,N_4544);
nor U5615 (N_5615,N_4654,N_3338);
xor U5616 (N_5616,N_3283,N_4431);
xor U5617 (N_5617,N_4048,N_4919);
and U5618 (N_5618,N_3913,N_4972);
nor U5619 (N_5619,N_3687,N_4980);
nor U5620 (N_5620,N_3840,N_2628);
or U5621 (N_5621,N_3187,N_2975);
and U5622 (N_5622,N_4461,N_4413);
xor U5623 (N_5623,N_4607,N_4286);
and U5624 (N_5624,N_2539,N_4578);
and U5625 (N_5625,N_4676,N_4736);
nand U5626 (N_5626,N_4822,N_3175);
or U5627 (N_5627,N_2504,N_2591);
nor U5628 (N_5628,N_2776,N_3741);
nor U5629 (N_5629,N_2569,N_4609);
and U5630 (N_5630,N_3933,N_3959);
nor U5631 (N_5631,N_2846,N_3111);
xnor U5632 (N_5632,N_3728,N_2626);
xnor U5633 (N_5633,N_4915,N_3564);
and U5634 (N_5634,N_2741,N_4926);
xor U5635 (N_5635,N_3648,N_4614);
nor U5636 (N_5636,N_3134,N_3604);
or U5637 (N_5637,N_3414,N_4757);
xor U5638 (N_5638,N_3437,N_3130);
nand U5639 (N_5639,N_2843,N_2650);
xnor U5640 (N_5640,N_3073,N_4786);
or U5641 (N_5641,N_4904,N_3290);
xor U5642 (N_5642,N_3885,N_4454);
nand U5643 (N_5643,N_4063,N_4735);
and U5644 (N_5644,N_3095,N_3632);
nand U5645 (N_5645,N_3268,N_3193);
xor U5646 (N_5646,N_4059,N_3755);
or U5647 (N_5647,N_4508,N_3867);
nand U5648 (N_5648,N_4605,N_3084);
or U5649 (N_5649,N_2748,N_2858);
or U5650 (N_5650,N_3151,N_4981);
nand U5651 (N_5651,N_4959,N_3427);
nor U5652 (N_5652,N_4380,N_3228);
or U5653 (N_5653,N_2589,N_2825);
nor U5654 (N_5654,N_4024,N_3790);
and U5655 (N_5655,N_4066,N_4260);
or U5656 (N_5656,N_3121,N_2823);
and U5657 (N_5657,N_4077,N_4526);
nand U5658 (N_5658,N_4518,N_2784);
xnor U5659 (N_5659,N_4180,N_3729);
xnor U5660 (N_5660,N_3670,N_3323);
or U5661 (N_5661,N_2840,N_3388);
and U5662 (N_5662,N_2898,N_4585);
and U5663 (N_5663,N_2775,N_3526);
or U5664 (N_5664,N_2907,N_4239);
xnor U5665 (N_5665,N_4608,N_4082);
and U5666 (N_5666,N_3416,N_4784);
or U5667 (N_5667,N_4262,N_2718);
xnor U5668 (N_5668,N_4533,N_4112);
or U5669 (N_5669,N_3061,N_3415);
and U5670 (N_5670,N_3336,N_2965);
xnor U5671 (N_5671,N_3613,N_4908);
nand U5672 (N_5672,N_3012,N_4951);
nor U5673 (N_5673,N_4961,N_2547);
xnor U5674 (N_5674,N_4236,N_3538);
nand U5675 (N_5675,N_3872,N_2596);
nor U5676 (N_5676,N_3260,N_4582);
or U5677 (N_5677,N_3371,N_2746);
nand U5678 (N_5678,N_4375,N_4483);
xor U5679 (N_5679,N_3832,N_3411);
xor U5680 (N_5680,N_3984,N_2973);
and U5681 (N_5681,N_2950,N_4502);
xor U5682 (N_5682,N_4182,N_3551);
xnor U5683 (N_5683,N_2574,N_3106);
xor U5684 (N_5684,N_3501,N_3471);
xnor U5685 (N_5685,N_3036,N_2513);
nand U5686 (N_5686,N_4628,N_2984);
xor U5687 (N_5687,N_4955,N_2872);
nand U5688 (N_5688,N_3715,N_4892);
xnor U5689 (N_5689,N_4924,N_4754);
nor U5690 (N_5690,N_2771,N_3827);
and U5691 (N_5691,N_3691,N_3549);
or U5692 (N_5692,N_3078,N_4850);
xnor U5693 (N_5693,N_3764,N_3400);
nand U5694 (N_5694,N_3567,N_2556);
or U5695 (N_5695,N_4320,N_3560);
xnor U5696 (N_5696,N_3641,N_3059);
nor U5697 (N_5697,N_4104,N_3002);
xor U5698 (N_5698,N_4281,N_3149);
nor U5699 (N_5699,N_2801,N_4469);
xnor U5700 (N_5700,N_4965,N_2755);
or U5701 (N_5701,N_3920,N_2665);
or U5702 (N_5702,N_3883,N_2713);
xnor U5703 (N_5703,N_3746,N_4135);
nor U5704 (N_5704,N_3561,N_4466);
nand U5705 (N_5705,N_4922,N_2522);
or U5706 (N_5706,N_4642,N_4798);
nor U5707 (N_5707,N_2934,N_3569);
nand U5708 (N_5708,N_4510,N_4703);
or U5709 (N_5709,N_4105,N_4560);
or U5710 (N_5710,N_4472,N_3536);
xor U5711 (N_5711,N_3218,N_4824);
nor U5712 (N_5712,N_3023,N_3192);
nand U5713 (N_5713,N_3431,N_4185);
xnor U5714 (N_5714,N_4336,N_3052);
and U5715 (N_5715,N_2500,N_3724);
xor U5716 (N_5716,N_2726,N_4450);
or U5717 (N_5717,N_3799,N_2737);
nand U5718 (N_5718,N_4627,N_3625);
and U5719 (N_5719,N_3521,N_3647);
nor U5720 (N_5720,N_4342,N_3385);
nand U5721 (N_5721,N_3194,N_4976);
nor U5722 (N_5722,N_2753,N_3777);
nand U5723 (N_5723,N_4939,N_3418);
nor U5724 (N_5724,N_4808,N_4967);
nor U5725 (N_5725,N_3658,N_2559);
or U5726 (N_5726,N_2501,N_4992);
and U5727 (N_5727,N_4015,N_3802);
nand U5728 (N_5728,N_4095,N_2508);
xnor U5729 (N_5729,N_4026,N_4524);
xnor U5730 (N_5730,N_4482,N_4804);
xor U5731 (N_5731,N_3426,N_4222);
or U5732 (N_5732,N_2717,N_4930);
xnor U5733 (N_5733,N_3236,N_2869);
xnor U5734 (N_5734,N_3057,N_3637);
xor U5735 (N_5735,N_3886,N_3005);
xor U5736 (N_5736,N_3940,N_3981);
xor U5737 (N_5737,N_3607,N_3654);
xnor U5738 (N_5738,N_4889,N_4697);
and U5739 (N_5739,N_3927,N_3312);
xnor U5740 (N_5740,N_2525,N_4506);
and U5741 (N_5741,N_4193,N_2543);
and U5742 (N_5742,N_3993,N_4599);
or U5743 (N_5743,N_3720,N_3181);
and U5744 (N_5744,N_4158,N_3524);
nand U5745 (N_5745,N_4551,N_2533);
or U5746 (N_5746,N_3771,N_3281);
and U5747 (N_5747,N_3072,N_2669);
xor U5748 (N_5748,N_4816,N_3525);
or U5749 (N_5749,N_3943,N_4795);
xor U5750 (N_5750,N_4927,N_3438);
or U5751 (N_5751,N_3828,N_4379);
xnor U5752 (N_5752,N_2794,N_4559);
or U5753 (N_5753,N_2831,N_3941);
and U5754 (N_5754,N_3683,N_3656);
or U5755 (N_5755,N_3709,N_4787);
and U5756 (N_5756,N_2796,N_2579);
nor U5757 (N_5757,N_3644,N_4729);
or U5758 (N_5758,N_2797,N_4113);
nand U5759 (N_5759,N_4731,N_2552);
nor U5760 (N_5760,N_3378,N_4042);
and U5761 (N_5761,N_2732,N_3226);
and U5762 (N_5762,N_4353,N_3344);
or U5763 (N_5763,N_4101,N_3449);
xor U5764 (N_5764,N_3932,N_2838);
xnor U5765 (N_5765,N_3681,N_2627);
xnor U5766 (N_5766,N_2988,N_2880);
nor U5767 (N_5767,N_4053,N_2526);
xor U5768 (N_5768,N_2643,N_2906);
xor U5769 (N_5769,N_3293,N_2584);
and U5770 (N_5770,N_4484,N_4345);
nor U5771 (N_5771,N_3577,N_3518);
or U5772 (N_5772,N_3760,N_3212);
nor U5773 (N_5773,N_2879,N_3122);
xnor U5774 (N_5774,N_4189,N_3351);
nor U5775 (N_5775,N_3881,N_3398);
nor U5776 (N_5776,N_3124,N_4561);
and U5777 (N_5777,N_3952,N_3204);
nand U5778 (N_5778,N_3817,N_2598);
xnor U5779 (N_5779,N_4902,N_4023);
nor U5780 (N_5780,N_3860,N_4812);
nand U5781 (N_5781,N_2994,N_3700);
and U5782 (N_5782,N_2580,N_4088);
or U5783 (N_5783,N_2545,N_3370);
nand U5784 (N_5784,N_3269,N_3256);
xnor U5785 (N_5785,N_2824,N_3138);
and U5786 (N_5786,N_2708,N_3379);
and U5787 (N_5787,N_2841,N_4275);
nand U5788 (N_5788,N_4837,N_4698);
and U5789 (N_5789,N_3793,N_3737);
or U5790 (N_5790,N_4384,N_4656);
xnor U5791 (N_5791,N_4659,N_3026);
xor U5792 (N_5792,N_4660,N_4276);
and U5793 (N_5793,N_2953,N_4139);
xnor U5794 (N_5794,N_4168,N_4903);
nand U5795 (N_5795,N_2578,N_3905);
nor U5796 (N_5796,N_3580,N_4191);
nand U5797 (N_5797,N_3346,N_2518);
xor U5798 (N_5798,N_3807,N_3997);
nor U5799 (N_5799,N_4541,N_4986);
nand U5800 (N_5800,N_4069,N_2576);
and U5801 (N_5801,N_2781,N_2893);
nor U5802 (N_5802,N_2905,N_2633);
nor U5803 (N_5803,N_3049,N_2827);
xnor U5804 (N_5804,N_4455,N_3667);
nor U5805 (N_5805,N_3092,N_3041);
or U5806 (N_5806,N_4964,N_3171);
nor U5807 (N_5807,N_4055,N_4468);
nor U5808 (N_5808,N_4225,N_4829);
nor U5809 (N_5809,N_4192,N_4408);
xnor U5810 (N_5810,N_2674,N_3623);
xnor U5811 (N_5811,N_4809,N_4906);
xnor U5812 (N_5812,N_2996,N_2696);
nand U5813 (N_5813,N_4245,N_4737);
and U5814 (N_5814,N_4788,N_2828);
xnor U5815 (N_5815,N_4050,N_4355);
and U5816 (N_5816,N_3436,N_2554);
or U5817 (N_5817,N_3803,N_4430);
nor U5818 (N_5818,N_4489,N_3666);
nand U5819 (N_5819,N_3705,N_4589);
and U5820 (N_5820,N_4751,N_4210);
or U5821 (N_5821,N_3702,N_4670);
and U5822 (N_5822,N_3590,N_3986);
nand U5823 (N_5823,N_4806,N_4775);
or U5824 (N_5824,N_4858,N_3922);
nor U5825 (N_5825,N_3196,N_3915);
nor U5826 (N_5826,N_3502,N_3170);
nand U5827 (N_5827,N_3768,N_3545);
nor U5828 (N_5828,N_2989,N_2792);
or U5829 (N_5829,N_2918,N_4111);
and U5830 (N_5830,N_3076,N_3244);
xnor U5831 (N_5831,N_2868,N_4406);
nand U5832 (N_5832,N_4505,N_2899);
nand U5833 (N_5833,N_3140,N_4284);
nand U5834 (N_5834,N_4548,N_4490);
or U5835 (N_5835,N_3279,N_3969);
nand U5836 (N_5836,N_3829,N_2712);
and U5837 (N_5837,N_3924,N_4673);
nor U5838 (N_5838,N_3582,N_4021);
xnor U5839 (N_5839,N_4813,N_2791);
and U5840 (N_5840,N_4741,N_3766);
xor U5841 (N_5841,N_3695,N_4310);
xnor U5842 (N_5842,N_4073,N_4566);
nand U5843 (N_5843,N_3878,N_4817);
nand U5844 (N_5844,N_3080,N_4936);
xnor U5845 (N_5845,N_3934,N_3056);
xor U5846 (N_5846,N_4304,N_3229);
or U5847 (N_5847,N_3325,N_3382);
and U5848 (N_5848,N_2857,N_3812);
or U5849 (N_5849,N_4695,N_4241);
nor U5850 (N_5850,N_4895,N_3000);
xor U5851 (N_5851,N_4875,N_4756);
or U5852 (N_5852,N_4910,N_3125);
xor U5853 (N_5853,N_4982,N_3112);
and U5854 (N_5854,N_4721,N_4558);
xor U5855 (N_5855,N_4760,N_4797);
nand U5856 (N_5856,N_4853,N_3556);
nor U5857 (N_5857,N_4952,N_4771);
or U5858 (N_5858,N_2995,N_4882);
or U5859 (N_5859,N_4682,N_3068);
xnor U5860 (N_5860,N_4652,N_3455);
nor U5861 (N_5861,N_4958,N_4602);
or U5862 (N_5862,N_3387,N_2876);
nand U5863 (N_5863,N_2894,N_4819);
nand U5864 (N_5864,N_4330,N_3708);
and U5865 (N_5865,N_4994,N_3541);
or U5866 (N_5866,N_4194,N_4701);
and U5867 (N_5867,N_2671,N_4488);
xor U5868 (N_5868,N_4029,N_3086);
nor U5869 (N_5869,N_4493,N_3747);
xnor U5870 (N_5870,N_4543,N_4761);
and U5871 (N_5871,N_2820,N_2779);
and U5872 (N_5872,N_2765,N_3158);
nand U5873 (N_5873,N_2606,N_3595);
or U5874 (N_5874,N_4285,N_4044);
nor U5875 (N_5875,N_3890,N_2977);
xnor U5876 (N_5876,N_4622,N_4691);
or U5877 (N_5877,N_3917,N_3403);
and U5878 (N_5878,N_3490,N_3133);
or U5879 (N_5879,N_3120,N_4842);
nor U5880 (N_5880,N_2842,N_3672);
nand U5881 (N_5881,N_3756,N_2970);
nand U5882 (N_5882,N_3364,N_4724);
xnor U5883 (N_5883,N_4881,N_2810);
xnor U5884 (N_5884,N_2724,N_4462);
and U5885 (N_5885,N_3553,N_3217);
or U5886 (N_5886,N_4280,N_2592);
and U5887 (N_5887,N_4362,N_4545);
nand U5888 (N_5888,N_3992,N_4052);
and U5889 (N_5889,N_4696,N_4790);
nor U5890 (N_5890,N_3721,N_3173);
nand U5891 (N_5891,N_4487,N_4625);
nand U5892 (N_5892,N_3519,N_2944);
xor U5893 (N_5893,N_4868,N_3284);
and U5894 (N_5894,N_2585,N_2588);
or U5895 (N_5895,N_4108,N_4118);
xnor U5896 (N_5896,N_4398,N_4966);
xnor U5897 (N_5897,N_4393,N_4479);
nor U5898 (N_5898,N_3898,N_4864);
or U5899 (N_5899,N_4590,N_2524);
and U5900 (N_5900,N_4421,N_2766);
or U5901 (N_5901,N_4133,N_3980);
and U5902 (N_5902,N_4990,N_3033);
and U5903 (N_5903,N_3375,N_4347);
nand U5904 (N_5904,N_3360,N_3876);
or U5905 (N_5905,N_2897,N_3663);
xnor U5906 (N_5906,N_3926,N_4170);
nand U5907 (N_5907,N_4621,N_4235);
nand U5908 (N_5908,N_4928,N_2720);
nand U5909 (N_5909,N_3520,N_4196);
nand U5910 (N_5910,N_3537,N_3091);
xor U5911 (N_5911,N_3272,N_3147);
and U5912 (N_5912,N_3254,N_3619);
nor U5913 (N_5913,N_3198,N_3046);
and U5914 (N_5914,N_3711,N_4388);
nor U5915 (N_5915,N_3939,N_4937);
nand U5916 (N_5916,N_3045,N_4299);
nor U5917 (N_5917,N_2542,N_3352);
nor U5918 (N_5918,N_4163,N_2683);
nand U5919 (N_5919,N_4247,N_3037);
xnor U5920 (N_5920,N_2758,N_2903);
nand U5921 (N_5921,N_4828,N_4093);
nor U5922 (N_5922,N_3113,N_4110);
nand U5923 (N_5923,N_4143,N_3432);
and U5924 (N_5924,N_3833,N_4159);
or U5925 (N_5925,N_3024,N_2527);
nor U5926 (N_5926,N_4529,N_4860);
or U5927 (N_5927,N_3237,N_3286);
xor U5928 (N_5928,N_2680,N_2672);
and U5929 (N_5929,N_3202,N_3064);
nand U5930 (N_5930,N_4623,N_3361);
and U5931 (N_5931,N_2961,N_4122);
nand U5932 (N_5932,N_3435,N_3972);
xor U5933 (N_5933,N_3365,N_3190);
and U5934 (N_5934,N_4216,N_4644);
nor U5935 (N_5935,N_4060,N_4707);
nor U5936 (N_5936,N_3510,N_4711);
and U5937 (N_5937,N_2521,N_4126);
xnor U5938 (N_5938,N_4442,N_3328);
nand U5939 (N_5939,N_4283,N_4914);
nand U5940 (N_5940,N_3494,N_4983);
xor U5941 (N_5941,N_4949,N_3456);
and U5942 (N_5942,N_3585,N_4475);
nor U5943 (N_5943,N_3417,N_3463);
nand U5944 (N_5944,N_4164,N_4874);
xnor U5945 (N_5945,N_3633,N_2624);
and U5946 (N_5946,N_4047,N_4632);
or U5947 (N_5947,N_2615,N_4359);
or U5948 (N_5948,N_4229,N_3778);
or U5949 (N_5949,N_3575,N_4743);
or U5950 (N_5950,N_3165,N_3222);
nor U5951 (N_5951,N_2536,N_3017);
and U5952 (N_5952,N_3031,N_3356);
and U5953 (N_5953,N_3055,N_2817);
and U5954 (N_5954,N_3914,N_3396);
nand U5955 (N_5955,N_3340,N_4087);
and U5956 (N_5956,N_4598,N_2634);
xor U5957 (N_5957,N_4793,N_4233);
xor U5958 (N_5958,N_3274,N_4134);
nor U5959 (N_5959,N_3838,N_3297);
nand U5960 (N_5960,N_4896,N_3679);
nand U5961 (N_5961,N_3499,N_4932);
nand U5962 (N_5962,N_4855,N_3044);
nor U5963 (N_5963,N_4549,N_4686);
or U5964 (N_5964,N_3704,N_2952);
nor U5965 (N_5965,N_3725,N_3931);
nand U5966 (N_5966,N_3770,N_4090);
or U5967 (N_5967,N_2602,N_4480);
nor U5968 (N_5968,N_4160,N_2943);
nand U5969 (N_5969,N_2736,N_3837);
or U5970 (N_5970,N_2505,N_3424);
nand U5971 (N_5971,N_3909,N_3957);
and U5972 (N_5972,N_4834,N_4835);
and U5973 (N_5973,N_2760,N_4177);
or U5974 (N_5974,N_4407,N_3988);
nor U5975 (N_5975,N_3317,N_3329);
xnor U5976 (N_5976,N_2612,N_3740);
or U5977 (N_5977,N_4973,N_3347);
or U5978 (N_5978,N_4378,N_2694);
and U5979 (N_5979,N_3752,N_4058);
xor U5980 (N_5980,N_3047,N_4546);
xnor U5981 (N_5981,N_2844,N_4016);
nand U5982 (N_5982,N_3131,N_3697);
nand U5983 (N_5983,N_2819,N_2939);
or U5984 (N_5984,N_3277,N_2815);
and U5985 (N_5985,N_4289,N_2981);
or U5986 (N_5986,N_2877,N_3889);
xor U5987 (N_5987,N_4340,N_3246);
nand U5988 (N_5988,N_4240,N_4458);
and U5989 (N_5989,N_3601,N_4190);
and U5990 (N_5990,N_3115,N_4148);
and U5991 (N_5991,N_2969,N_3392);
and U5992 (N_5992,N_3964,N_3409);
or U5993 (N_5993,N_3547,N_4888);
or U5994 (N_5994,N_4538,N_3335);
nor U5995 (N_5995,N_2945,N_3550);
nand U5996 (N_5996,N_3995,N_3851);
nand U5997 (N_5997,N_4041,N_3742);
nand U5998 (N_5998,N_3310,N_3079);
or U5999 (N_5999,N_3321,N_2716);
nor U6000 (N_6000,N_3146,N_3021);
or U6001 (N_6001,N_3320,N_4616);
or U6002 (N_6002,N_4014,N_3081);
nor U6003 (N_6003,N_3947,N_4153);
nand U6004 (N_6004,N_3785,N_4898);
and U6005 (N_6005,N_3593,N_3748);
nor U6006 (N_6006,N_4996,N_4401);
or U6007 (N_6007,N_4993,N_2922);
and U6008 (N_6008,N_4547,N_2668);
nor U6009 (N_6009,N_2687,N_4747);
nor U6010 (N_6010,N_4847,N_3331);
nor U6011 (N_6011,N_2923,N_4719);
xor U6012 (N_6012,N_2730,N_3727);
nor U6013 (N_6013,N_3978,N_2636);
nand U6014 (N_6014,N_3333,N_3621);
and U6015 (N_6015,N_3316,N_4575);
and U6016 (N_6016,N_3381,N_4708);
xnor U6017 (N_6017,N_4188,N_4348);
and U6018 (N_6018,N_2871,N_4514);
or U6019 (N_6019,N_4534,N_3821);
xor U6020 (N_6020,N_3001,N_4341);
nor U6021 (N_6021,N_4521,N_4130);
or U6022 (N_6022,N_3419,N_4445);
and U6023 (N_6023,N_2528,N_3476);
nor U6024 (N_6024,N_3295,N_4596);
or U6025 (N_6025,N_4894,N_3366);
and U6026 (N_6026,N_3083,N_2816);
nand U6027 (N_6027,N_4767,N_3126);
nand U6028 (N_6028,N_3105,N_4169);
xor U6029 (N_6029,N_3266,N_3888);
or U6030 (N_6030,N_4681,N_4588);
or U6031 (N_6031,N_3895,N_2617);
nor U6032 (N_6032,N_2699,N_2711);
xnor U6033 (N_6033,N_3763,N_3434);
nand U6034 (N_6034,N_2924,N_3263);
and U6035 (N_6035,N_2519,N_2581);
nand U6036 (N_6036,N_4467,N_4826);
and U6037 (N_6037,N_4580,N_4321);
nor U6038 (N_6038,N_3107,N_4950);
xnor U6039 (N_6039,N_2904,N_3429);
or U6040 (N_6040,N_4051,N_3150);
nand U6041 (N_6041,N_3628,N_3433);
and U6042 (N_6042,N_4184,N_3085);
nor U6043 (N_6043,N_4486,N_3326);
nand U6044 (N_6044,N_3177,N_2566);
xor U6045 (N_6045,N_3571,N_2631);
xor U6046 (N_6046,N_3574,N_4863);
nand U6047 (N_6047,N_3029,N_4801);
or U6048 (N_6048,N_3508,N_3638);
nor U6049 (N_6049,N_4601,N_4940);
and U6050 (N_6050,N_4377,N_4123);
or U6051 (N_6051,N_4361,N_3395);
xor U6052 (N_6052,N_4145,N_3789);
and U6053 (N_6053,N_4371,N_2707);
xor U6054 (N_6054,N_2616,N_4477);
nor U6055 (N_6055,N_3930,N_3207);
and U6056 (N_6056,N_4478,N_3749);
nor U6057 (N_6057,N_4782,N_4810);
or U6058 (N_6058,N_3004,N_2675);
nand U6059 (N_6059,N_3902,N_2558);
or U6060 (N_6060,N_2803,N_2870);
xor U6061 (N_6061,N_3219,N_2966);
nand U6062 (N_6062,N_4425,N_3744);
nor U6063 (N_6063,N_3008,N_3011);
and U6064 (N_6064,N_4917,N_3303);
xnor U6065 (N_6065,N_2863,N_4370);
xor U6066 (N_6066,N_4079,N_2511);
or U6067 (N_6067,N_4327,N_2982);
nor U6068 (N_6068,N_2604,N_2814);
nor U6069 (N_6069,N_3314,N_4947);
nand U6070 (N_6070,N_4443,N_4257);
nor U6071 (N_6071,N_2705,N_4131);
or U6072 (N_6072,N_4238,N_2709);
nor U6073 (N_6073,N_3735,N_3179);
and U6074 (N_6074,N_4136,N_4552);
nand U6075 (N_6075,N_3884,N_4349);
xnor U6076 (N_6076,N_4305,N_4416);
and U6077 (N_6077,N_4427,N_3509);
or U6078 (N_6078,N_3797,N_2845);
xnor U6079 (N_6079,N_4025,N_2534);
or U6080 (N_6080,N_4648,N_3404);
xnor U6081 (N_6081,N_2800,N_4641);
xnor U6082 (N_6082,N_4259,N_4040);
nor U6083 (N_6083,N_4970,N_2692);
xor U6084 (N_6084,N_4507,N_2849);
or U6085 (N_6085,N_3723,N_3985);
xnor U6086 (N_6086,N_3180,N_3483);
or U6087 (N_6087,N_4712,N_3259);
and U6088 (N_6088,N_3461,N_4905);
nor U6089 (N_6089,N_4899,N_4146);
nand U6090 (N_6090,N_4948,N_3384);
nand U6091 (N_6091,N_3738,N_3070);
xnor U6092 (N_6092,N_2867,N_2645);
or U6093 (N_6093,N_4186,N_3624);
xnor U6094 (N_6094,N_3015,N_4852);
nor U6095 (N_6095,N_4085,N_4728);
nor U6096 (N_6096,N_3470,N_2873);
nand U6097 (N_6097,N_3892,N_4800);
nand U6098 (N_6098,N_3342,N_3103);
nand U6099 (N_6099,N_3300,N_4758);
xor U6100 (N_6100,N_4876,N_2947);
or U6101 (N_6101,N_4255,N_2651);
and U6102 (N_6102,N_3443,N_4877);
and U6103 (N_6103,N_3353,N_2832);
xnor U6104 (N_6104,N_3921,N_3522);
or U6105 (N_6105,N_3779,N_4423);
nand U6106 (N_6106,N_3118,N_2954);
nand U6107 (N_6107,N_4033,N_3823);
xnor U6108 (N_6108,N_4867,N_4997);
or U6109 (N_6109,N_4762,N_4836);
nor U6110 (N_6110,N_4537,N_4435);
nand U6111 (N_6111,N_3782,N_2666);
nand U6112 (N_6112,N_3974,N_4753);
nor U6113 (N_6113,N_4011,N_3925);
xor U6114 (N_6114,N_3484,N_4662);
nand U6115 (N_6115,N_3854,N_3979);
nand U6116 (N_6116,N_3362,N_2613);
and U6117 (N_6117,N_3220,N_2941);
and U6118 (N_6118,N_4120,N_3784);
xor U6119 (N_6119,N_2728,N_3753);
nand U6120 (N_6120,N_3195,N_3276);
xor U6121 (N_6121,N_4206,N_3482);
xnor U6122 (N_6122,N_3003,N_2735);
or U6123 (N_6123,N_4638,N_2983);
and U6124 (N_6124,N_3013,N_3345);
or U6125 (N_6125,N_2516,N_3815);
or U6126 (N_6126,N_3282,N_3164);
or U6127 (N_6127,N_4400,N_3583);
nand U6128 (N_6128,N_4845,N_3546);
nand U6129 (N_6129,N_4742,N_3214);
nand U6130 (N_6130,N_4562,N_4374);
or U6131 (N_6131,N_4689,N_4886);
nor U6132 (N_6132,N_3503,N_2706);
or U6133 (N_6133,N_4441,N_4422);
and U6134 (N_6134,N_2594,N_3572);
or U6135 (N_6135,N_3227,N_2946);
nand U6136 (N_6136,N_4539,N_4500);
nand U6137 (N_6137,N_2851,N_3804);
or U6138 (N_6138,N_3376,N_4213);
and U6139 (N_6139,N_2567,N_3780);
and U6140 (N_6140,N_3578,N_4156);
nand U6141 (N_6141,N_3717,N_3486);
xnor U6142 (N_6142,N_4718,N_4667);
nand U6143 (N_6143,N_4032,N_4653);
nor U6144 (N_6144,N_3462,N_3558);
or U6145 (N_6145,N_4645,N_4279);
nand U6146 (N_6146,N_4783,N_4119);
xnor U6147 (N_6147,N_2854,N_2763);
nor U6148 (N_6148,N_3743,N_3160);
nand U6149 (N_6149,N_2759,N_2978);
nand U6150 (N_6150,N_2835,N_4584);
nor U6151 (N_6151,N_3048,N_3843);
nand U6152 (N_6152,N_3686,N_2673);
or U6153 (N_6153,N_3862,N_2911);
xnor U6154 (N_6154,N_4204,N_4389);
and U6155 (N_6155,N_4587,N_4647);
nand U6156 (N_6156,N_4634,N_3868);
and U6157 (N_6157,N_2667,N_3488);
or U6158 (N_6158,N_3032,N_3492);
xnor U6159 (N_6159,N_2931,N_4220);
xnor U6160 (N_6160,N_4318,N_4404);
or U6161 (N_6161,N_3581,N_4312);
nor U6162 (N_6162,N_2974,N_3144);
nor U6163 (N_6163,N_2538,N_3950);
or U6164 (N_6164,N_3241,N_3505);
or U6165 (N_6165,N_3154,N_3730);
and U6166 (N_6166,N_4920,N_4519);
or U6167 (N_6167,N_3299,N_4792);
or U6168 (N_6168,N_2891,N_3189);
nand U6169 (N_6169,N_3948,N_3818);
xor U6170 (N_6170,N_2833,N_4366);
and U6171 (N_6171,N_3298,N_4008);
nor U6172 (N_6172,N_3231,N_4440);
nand U6173 (N_6173,N_4329,N_2655);
or U6174 (N_6174,N_3157,N_4778);
xnor U6175 (N_6175,N_4178,N_4314);
nand U6176 (N_6176,N_2510,N_3460);
or U6177 (N_6177,N_4096,N_4001);
and U6178 (N_6178,N_2967,N_4420);
and U6179 (N_6179,N_4796,N_4494);
nand U6180 (N_6180,N_3440,N_2949);
and U6181 (N_6181,N_4649,N_3273);
and U6182 (N_6182,N_4677,N_2910);
and U6183 (N_6183,N_3762,N_4409);
and U6184 (N_6184,N_4946,N_3232);
xor U6185 (N_6185,N_2963,N_4749);
or U6186 (N_6186,N_4619,N_4419);
nor U6187 (N_6187,N_4555,N_4637);
or U6188 (N_6188,N_3767,N_4974);
and U6189 (N_6189,N_4693,N_3156);
xnor U6190 (N_6190,N_2557,N_4911);
xnor U6191 (N_6191,N_3075,N_3511);
nor U6192 (N_6192,N_4827,N_3706);
xnor U6193 (N_6193,N_4417,N_4175);
or U6194 (N_6194,N_4092,N_4752);
and U6195 (N_6195,N_4773,N_3535);
xnor U6196 (N_6196,N_3810,N_4215);
xor U6197 (N_6197,N_4664,N_3875);
nand U6198 (N_6198,N_4891,N_4720);
nor U6199 (N_6199,N_3225,N_3605);
nor U6200 (N_6200,N_4212,N_4977);
or U6201 (N_6201,N_2780,N_2695);
and U6202 (N_6202,N_4243,N_4263);
and U6203 (N_6203,N_4117,N_3261);
or U6204 (N_6204,N_3573,N_4457);
and U6205 (N_6205,N_4199,N_4501);
nor U6206 (N_6206,N_4203,N_2529);
or U6207 (N_6207,N_3042,N_3296);
nor U6208 (N_6208,N_4337,N_3548);
nor U6209 (N_6209,N_4699,N_4639);
and U6210 (N_6210,N_4311,N_3646);
xor U6211 (N_6211,N_2782,N_4779);
nand U6212 (N_6212,N_2535,N_2750);
nand U6213 (N_6213,N_4005,N_3035);
or U6214 (N_6214,N_2895,N_4181);
or U6215 (N_6215,N_3935,N_2749);
or U6216 (N_6216,N_4295,N_2874);
nand U6217 (N_6217,N_3481,N_4306);
nor U6218 (N_6218,N_4248,N_3087);
xnor U6219 (N_6219,N_3718,N_4390);
and U6220 (N_6220,N_2860,N_3694);
xnor U6221 (N_6221,N_4515,N_2625);
nor U6222 (N_6222,N_3703,N_4003);
nor U6223 (N_6223,N_4453,N_3542);
nor U6224 (N_6224,N_4781,N_4527);
nand U6225 (N_6225,N_4633,N_3568);
nor U6226 (N_6226,N_4446,N_3186);
or U6227 (N_6227,N_2942,N_4726);
nor U6228 (N_6228,N_2551,N_4931);
nor U6229 (N_6229,N_3801,N_3996);
nand U6230 (N_6230,N_3096,N_2648);
nor U6231 (N_6231,N_2520,N_3135);
and U6232 (N_6232,N_4768,N_4154);
xor U6233 (N_6233,N_3879,N_3712);
and U6234 (N_6234,N_4142,N_4237);
and U6235 (N_6235,N_3594,N_2609);
nor U6236 (N_6236,N_4332,N_4710);
nand U6237 (N_6237,N_4328,N_2572);
xor U6238 (N_6238,N_3238,N_3651);
xnor U6239 (N_6239,N_3754,N_4232);
or U6240 (N_6240,N_2658,N_4428);
nand U6241 (N_6241,N_2620,N_3119);
nand U6242 (N_6242,N_3852,N_4103);
and U6243 (N_6243,N_3634,N_3459);
and U6244 (N_6244,N_2986,N_2826);
nand U6245 (N_6245,N_4396,N_3820);
nand U6246 (N_6246,N_4583,N_2642);
and U6247 (N_6247,N_3975,N_3662);
nor U6248 (N_6248,N_3448,N_4520);
or U6249 (N_6249,N_3082,N_4841);
nand U6250 (N_6250,N_3099,N_3972);
and U6251 (N_6251,N_4695,N_2743);
nand U6252 (N_6252,N_4342,N_3442);
and U6253 (N_6253,N_3186,N_3396);
xnor U6254 (N_6254,N_2500,N_4257);
nor U6255 (N_6255,N_3182,N_2722);
xor U6256 (N_6256,N_3155,N_2697);
nand U6257 (N_6257,N_4444,N_3270);
nand U6258 (N_6258,N_4015,N_2955);
nor U6259 (N_6259,N_3754,N_4905);
xnor U6260 (N_6260,N_3455,N_3321);
or U6261 (N_6261,N_4514,N_4033);
xor U6262 (N_6262,N_2741,N_3591);
nand U6263 (N_6263,N_3550,N_4852);
nor U6264 (N_6264,N_3881,N_2923);
or U6265 (N_6265,N_4039,N_4383);
xnor U6266 (N_6266,N_3641,N_2861);
nand U6267 (N_6267,N_3900,N_4628);
or U6268 (N_6268,N_2531,N_4170);
and U6269 (N_6269,N_3554,N_3707);
nand U6270 (N_6270,N_4818,N_3669);
nand U6271 (N_6271,N_2841,N_2927);
xor U6272 (N_6272,N_2920,N_2927);
nand U6273 (N_6273,N_4462,N_4194);
or U6274 (N_6274,N_2690,N_4041);
or U6275 (N_6275,N_4164,N_4446);
nand U6276 (N_6276,N_3849,N_3476);
xnor U6277 (N_6277,N_3199,N_4966);
nand U6278 (N_6278,N_4837,N_3731);
nor U6279 (N_6279,N_4694,N_2544);
or U6280 (N_6280,N_4630,N_3886);
nand U6281 (N_6281,N_3430,N_2511);
and U6282 (N_6282,N_3113,N_4596);
xnor U6283 (N_6283,N_4695,N_3386);
nand U6284 (N_6284,N_4467,N_4517);
or U6285 (N_6285,N_4911,N_4755);
or U6286 (N_6286,N_4915,N_2833);
nor U6287 (N_6287,N_3899,N_3785);
nand U6288 (N_6288,N_2520,N_3013);
nor U6289 (N_6289,N_2888,N_4169);
nand U6290 (N_6290,N_3149,N_4817);
or U6291 (N_6291,N_3344,N_4247);
nor U6292 (N_6292,N_4589,N_3698);
or U6293 (N_6293,N_3590,N_4238);
or U6294 (N_6294,N_3935,N_4062);
xnor U6295 (N_6295,N_3767,N_2997);
nand U6296 (N_6296,N_2807,N_4525);
nor U6297 (N_6297,N_4223,N_4819);
nor U6298 (N_6298,N_3945,N_4163);
nor U6299 (N_6299,N_4751,N_4902);
xnor U6300 (N_6300,N_2725,N_2520);
or U6301 (N_6301,N_4246,N_2654);
nor U6302 (N_6302,N_4761,N_4934);
or U6303 (N_6303,N_4210,N_2713);
nor U6304 (N_6304,N_4444,N_3300);
nor U6305 (N_6305,N_2675,N_3009);
xnor U6306 (N_6306,N_3019,N_3130);
nand U6307 (N_6307,N_3365,N_2923);
and U6308 (N_6308,N_2857,N_3868);
or U6309 (N_6309,N_4658,N_3653);
or U6310 (N_6310,N_3566,N_3928);
or U6311 (N_6311,N_4774,N_3486);
nand U6312 (N_6312,N_2919,N_3600);
or U6313 (N_6313,N_2515,N_4750);
and U6314 (N_6314,N_3741,N_3180);
xor U6315 (N_6315,N_4806,N_3781);
nand U6316 (N_6316,N_3635,N_4159);
and U6317 (N_6317,N_2765,N_4052);
xnor U6318 (N_6318,N_3830,N_4959);
xor U6319 (N_6319,N_3517,N_3694);
nor U6320 (N_6320,N_3942,N_3856);
nand U6321 (N_6321,N_3828,N_4328);
and U6322 (N_6322,N_4655,N_2546);
or U6323 (N_6323,N_4110,N_4760);
xor U6324 (N_6324,N_2950,N_4065);
nand U6325 (N_6325,N_3331,N_3541);
or U6326 (N_6326,N_3795,N_4407);
or U6327 (N_6327,N_3930,N_2652);
and U6328 (N_6328,N_3779,N_4834);
nand U6329 (N_6329,N_4651,N_3821);
or U6330 (N_6330,N_3572,N_4014);
nand U6331 (N_6331,N_4024,N_3414);
or U6332 (N_6332,N_3911,N_3350);
xor U6333 (N_6333,N_3063,N_4312);
xor U6334 (N_6334,N_4917,N_2874);
nor U6335 (N_6335,N_2865,N_2864);
xor U6336 (N_6336,N_2904,N_2970);
or U6337 (N_6337,N_3454,N_2520);
nand U6338 (N_6338,N_3086,N_3162);
xor U6339 (N_6339,N_4703,N_3454);
xnor U6340 (N_6340,N_4238,N_4677);
xor U6341 (N_6341,N_3047,N_3933);
or U6342 (N_6342,N_3623,N_4126);
or U6343 (N_6343,N_3218,N_3764);
nor U6344 (N_6344,N_2895,N_2507);
nand U6345 (N_6345,N_4444,N_2904);
nand U6346 (N_6346,N_4775,N_4383);
or U6347 (N_6347,N_3415,N_3450);
nor U6348 (N_6348,N_3243,N_3054);
nand U6349 (N_6349,N_2896,N_3746);
xor U6350 (N_6350,N_3139,N_3409);
nand U6351 (N_6351,N_3486,N_3805);
nand U6352 (N_6352,N_2708,N_4478);
nand U6353 (N_6353,N_4231,N_3579);
nor U6354 (N_6354,N_4082,N_4801);
or U6355 (N_6355,N_3247,N_2678);
nand U6356 (N_6356,N_4715,N_3179);
and U6357 (N_6357,N_4040,N_3475);
nor U6358 (N_6358,N_4534,N_2702);
nor U6359 (N_6359,N_3411,N_3615);
nor U6360 (N_6360,N_3793,N_4771);
and U6361 (N_6361,N_2577,N_3016);
nand U6362 (N_6362,N_3873,N_4643);
nor U6363 (N_6363,N_4254,N_3717);
and U6364 (N_6364,N_4965,N_4801);
or U6365 (N_6365,N_2641,N_4622);
or U6366 (N_6366,N_3584,N_3277);
nor U6367 (N_6367,N_4000,N_3928);
and U6368 (N_6368,N_2535,N_2715);
nand U6369 (N_6369,N_4506,N_3110);
or U6370 (N_6370,N_2621,N_3057);
and U6371 (N_6371,N_2962,N_2614);
nor U6372 (N_6372,N_4198,N_3936);
and U6373 (N_6373,N_4531,N_4935);
xor U6374 (N_6374,N_3078,N_3588);
nand U6375 (N_6375,N_3023,N_3883);
nand U6376 (N_6376,N_3204,N_3858);
xor U6377 (N_6377,N_4143,N_4327);
nand U6378 (N_6378,N_3187,N_3336);
or U6379 (N_6379,N_4475,N_4334);
nor U6380 (N_6380,N_3660,N_2718);
xnor U6381 (N_6381,N_3648,N_4238);
and U6382 (N_6382,N_3252,N_4426);
and U6383 (N_6383,N_4463,N_3564);
nand U6384 (N_6384,N_3699,N_3750);
nor U6385 (N_6385,N_3448,N_4339);
and U6386 (N_6386,N_4719,N_4896);
nand U6387 (N_6387,N_2561,N_3659);
xnor U6388 (N_6388,N_3959,N_2607);
or U6389 (N_6389,N_2965,N_3161);
nand U6390 (N_6390,N_4376,N_3862);
nor U6391 (N_6391,N_4198,N_4980);
or U6392 (N_6392,N_4742,N_4444);
xnor U6393 (N_6393,N_3781,N_4060);
nor U6394 (N_6394,N_2789,N_3953);
nor U6395 (N_6395,N_3387,N_2712);
nand U6396 (N_6396,N_3489,N_3160);
nand U6397 (N_6397,N_4770,N_3969);
or U6398 (N_6398,N_4684,N_3740);
and U6399 (N_6399,N_4495,N_3919);
nor U6400 (N_6400,N_3818,N_3554);
and U6401 (N_6401,N_4690,N_4022);
nand U6402 (N_6402,N_4398,N_2792);
and U6403 (N_6403,N_4678,N_4084);
nand U6404 (N_6404,N_4231,N_2806);
nor U6405 (N_6405,N_4733,N_4019);
and U6406 (N_6406,N_4848,N_3532);
nand U6407 (N_6407,N_3938,N_4646);
xor U6408 (N_6408,N_4352,N_3320);
nand U6409 (N_6409,N_3614,N_2761);
xor U6410 (N_6410,N_3673,N_2939);
or U6411 (N_6411,N_4631,N_4741);
xnor U6412 (N_6412,N_3887,N_4535);
and U6413 (N_6413,N_4999,N_3652);
nor U6414 (N_6414,N_3385,N_4908);
nor U6415 (N_6415,N_3535,N_4014);
xor U6416 (N_6416,N_2636,N_3308);
or U6417 (N_6417,N_3403,N_4083);
nand U6418 (N_6418,N_3462,N_2841);
and U6419 (N_6419,N_4417,N_2736);
nand U6420 (N_6420,N_3269,N_3982);
nor U6421 (N_6421,N_4589,N_2684);
xor U6422 (N_6422,N_3432,N_3499);
nor U6423 (N_6423,N_3567,N_3806);
nor U6424 (N_6424,N_3391,N_2667);
xnor U6425 (N_6425,N_3419,N_2981);
or U6426 (N_6426,N_3267,N_4856);
or U6427 (N_6427,N_4009,N_3625);
nor U6428 (N_6428,N_2825,N_3021);
or U6429 (N_6429,N_3389,N_3588);
xor U6430 (N_6430,N_3001,N_3845);
xnor U6431 (N_6431,N_3043,N_4558);
and U6432 (N_6432,N_3167,N_4294);
and U6433 (N_6433,N_3936,N_4655);
and U6434 (N_6434,N_3891,N_4391);
or U6435 (N_6435,N_3754,N_3121);
nand U6436 (N_6436,N_4930,N_4842);
xor U6437 (N_6437,N_3301,N_3432);
nor U6438 (N_6438,N_4022,N_3187);
xor U6439 (N_6439,N_4399,N_3905);
and U6440 (N_6440,N_3574,N_3756);
and U6441 (N_6441,N_3256,N_3786);
nand U6442 (N_6442,N_4648,N_2860);
or U6443 (N_6443,N_4663,N_2733);
nand U6444 (N_6444,N_3436,N_4540);
xnor U6445 (N_6445,N_4278,N_2502);
and U6446 (N_6446,N_3616,N_2695);
or U6447 (N_6447,N_4714,N_2584);
or U6448 (N_6448,N_4750,N_4428);
xor U6449 (N_6449,N_3782,N_3401);
xnor U6450 (N_6450,N_4723,N_3941);
and U6451 (N_6451,N_4035,N_3143);
xnor U6452 (N_6452,N_2914,N_3972);
nand U6453 (N_6453,N_3329,N_4684);
or U6454 (N_6454,N_2992,N_4026);
nand U6455 (N_6455,N_4237,N_2999);
nor U6456 (N_6456,N_4088,N_4494);
and U6457 (N_6457,N_3757,N_3025);
and U6458 (N_6458,N_4824,N_2847);
nand U6459 (N_6459,N_4494,N_4625);
nand U6460 (N_6460,N_4911,N_4062);
xor U6461 (N_6461,N_4712,N_3507);
or U6462 (N_6462,N_3125,N_2642);
xnor U6463 (N_6463,N_4591,N_4489);
nor U6464 (N_6464,N_4900,N_2578);
nand U6465 (N_6465,N_3472,N_3822);
xor U6466 (N_6466,N_4658,N_2817);
nand U6467 (N_6467,N_3579,N_4298);
and U6468 (N_6468,N_3868,N_4125);
xor U6469 (N_6469,N_3902,N_4976);
xnor U6470 (N_6470,N_4767,N_2702);
nand U6471 (N_6471,N_4657,N_3969);
and U6472 (N_6472,N_2880,N_4292);
nor U6473 (N_6473,N_2806,N_4896);
nor U6474 (N_6474,N_3525,N_3594);
and U6475 (N_6475,N_2925,N_3633);
nand U6476 (N_6476,N_3067,N_4532);
xor U6477 (N_6477,N_4549,N_4141);
and U6478 (N_6478,N_4427,N_2982);
or U6479 (N_6479,N_2800,N_2952);
nor U6480 (N_6480,N_3904,N_4506);
or U6481 (N_6481,N_4749,N_3632);
nand U6482 (N_6482,N_3675,N_3302);
xnor U6483 (N_6483,N_3732,N_3266);
nand U6484 (N_6484,N_4268,N_4273);
xor U6485 (N_6485,N_3474,N_2798);
or U6486 (N_6486,N_2520,N_3626);
nand U6487 (N_6487,N_4618,N_2958);
nand U6488 (N_6488,N_2989,N_4090);
xnor U6489 (N_6489,N_3019,N_3084);
nor U6490 (N_6490,N_3834,N_2610);
nand U6491 (N_6491,N_3877,N_4892);
xnor U6492 (N_6492,N_4107,N_3187);
or U6493 (N_6493,N_3562,N_3577);
and U6494 (N_6494,N_4690,N_3101);
or U6495 (N_6495,N_4594,N_2676);
nor U6496 (N_6496,N_4301,N_4551);
or U6497 (N_6497,N_3250,N_3749);
and U6498 (N_6498,N_3037,N_4224);
and U6499 (N_6499,N_3378,N_2715);
nand U6500 (N_6500,N_4317,N_2860);
or U6501 (N_6501,N_4798,N_3995);
xnor U6502 (N_6502,N_3618,N_4335);
nor U6503 (N_6503,N_3664,N_3401);
and U6504 (N_6504,N_3072,N_2989);
xor U6505 (N_6505,N_4660,N_2630);
and U6506 (N_6506,N_4991,N_2854);
nor U6507 (N_6507,N_2661,N_3020);
xnor U6508 (N_6508,N_4867,N_4754);
nand U6509 (N_6509,N_3053,N_4352);
and U6510 (N_6510,N_3002,N_3823);
xor U6511 (N_6511,N_4640,N_4529);
nor U6512 (N_6512,N_4644,N_4374);
or U6513 (N_6513,N_4176,N_3832);
nor U6514 (N_6514,N_4281,N_3225);
nor U6515 (N_6515,N_3771,N_2673);
or U6516 (N_6516,N_4344,N_4258);
nor U6517 (N_6517,N_2566,N_3801);
and U6518 (N_6518,N_3814,N_3056);
and U6519 (N_6519,N_3442,N_3559);
and U6520 (N_6520,N_2562,N_3778);
nand U6521 (N_6521,N_3367,N_4761);
nor U6522 (N_6522,N_3679,N_4184);
or U6523 (N_6523,N_3946,N_3486);
or U6524 (N_6524,N_4912,N_3213);
and U6525 (N_6525,N_4730,N_3402);
xor U6526 (N_6526,N_4629,N_3724);
xnor U6527 (N_6527,N_3183,N_3285);
nand U6528 (N_6528,N_3811,N_3370);
or U6529 (N_6529,N_3839,N_3937);
and U6530 (N_6530,N_2864,N_3836);
and U6531 (N_6531,N_3474,N_3749);
and U6532 (N_6532,N_3165,N_3144);
nor U6533 (N_6533,N_3866,N_3960);
nor U6534 (N_6534,N_4024,N_4693);
nor U6535 (N_6535,N_4909,N_4000);
nand U6536 (N_6536,N_2798,N_3248);
xnor U6537 (N_6537,N_2819,N_3040);
or U6538 (N_6538,N_3442,N_4076);
and U6539 (N_6539,N_3448,N_3902);
and U6540 (N_6540,N_3554,N_3512);
xnor U6541 (N_6541,N_4498,N_3359);
and U6542 (N_6542,N_3748,N_4634);
xor U6543 (N_6543,N_3298,N_4277);
or U6544 (N_6544,N_3370,N_3443);
and U6545 (N_6545,N_4389,N_2535);
xor U6546 (N_6546,N_4048,N_3901);
nand U6547 (N_6547,N_2805,N_2822);
nand U6548 (N_6548,N_3058,N_2922);
or U6549 (N_6549,N_2507,N_4211);
xnor U6550 (N_6550,N_3443,N_3480);
or U6551 (N_6551,N_2517,N_3113);
nand U6552 (N_6552,N_4165,N_4420);
or U6553 (N_6553,N_3608,N_3386);
nor U6554 (N_6554,N_3226,N_3669);
and U6555 (N_6555,N_3882,N_3920);
nand U6556 (N_6556,N_3127,N_4632);
xnor U6557 (N_6557,N_4557,N_4741);
and U6558 (N_6558,N_3369,N_3340);
xnor U6559 (N_6559,N_4593,N_3998);
xnor U6560 (N_6560,N_3789,N_2549);
or U6561 (N_6561,N_4677,N_2659);
xnor U6562 (N_6562,N_4968,N_2759);
or U6563 (N_6563,N_3631,N_3626);
xnor U6564 (N_6564,N_4079,N_4649);
or U6565 (N_6565,N_3946,N_3420);
and U6566 (N_6566,N_4345,N_2881);
nor U6567 (N_6567,N_3025,N_2928);
and U6568 (N_6568,N_3299,N_3643);
nand U6569 (N_6569,N_4944,N_4628);
or U6570 (N_6570,N_2808,N_4223);
nor U6571 (N_6571,N_3258,N_4672);
or U6572 (N_6572,N_4624,N_3357);
xnor U6573 (N_6573,N_2628,N_3657);
and U6574 (N_6574,N_2847,N_4697);
nor U6575 (N_6575,N_3192,N_4204);
xnor U6576 (N_6576,N_4316,N_3884);
or U6577 (N_6577,N_4563,N_4820);
or U6578 (N_6578,N_4855,N_4853);
nor U6579 (N_6579,N_4405,N_4989);
and U6580 (N_6580,N_3977,N_3553);
nand U6581 (N_6581,N_2520,N_4096);
or U6582 (N_6582,N_3663,N_4879);
nand U6583 (N_6583,N_4653,N_4417);
xor U6584 (N_6584,N_3350,N_4692);
nor U6585 (N_6585,N_2906,N_4241);
xnor U6586 (N_6586,N_3859,N_2754);
nand U6587 (N_6587,N_4942,N_2677);
nor U6588 (N_6588,N_2770,N_3648);
nand U6589 (N_6589,N_4723,N_4022);
or U6590 (N_6590,N_3764,N_4898);
nor U6591 (N_6591,N_3207,N_2895);
or U6592 (N_6592,N_4870,N_2606);
nand U6593 (N_6593,N_4659,N_2956);
and U6594 (N_6594,N_4628,N_3691);
nor U6595 (N_6595,N_2649,N_4981);
and U6596 (N_6596,N_2573,N_4465);
xor U6597 (N_6597,N_3961,N_2637);
or U6598 (N_6598,N_4173,N_4203);
nand U6599 (N_6599,N_4486,N_4946);
nor U6600 (N_6600,N_2662,N_4163);
or U6601 (N_6601,N_4927,N_3408);
nand U6602 (N_6602,N_2916,N_3408);
or U6603 (N_6603,N_3318,N_4028);
nand U6604 (N_6604,N_4820,N_3926);
or U6605 (N_6605,N_4589,N_4299);
nand U6606 (N_6606,N_4511,N_2680);
nor U6607 (N_6607,N_3363,N_3037);
xnor U6608 (N_6608,N_2523,N_4862);
nor U6609 (N_6609,N_3660,N_3545);
nand U6610 (N_6610,N_2564,N_2772);
xor U6611 (N_6611,N_4324,N_3869);
nand U6612 (N_6612,N_4141,N_4689);
or U6613 (N_6613,N_4916,N_4747);
or U6614 (N_6614,N_4777,N_4311);
and U6615 (N_6615,N_3640,N_3667);
xnor U6616 (N_6616,N_4493,N_3351);
nor U6617 (N_6617,N_4021,N_4490);
or U6618 (N_6618,N_3931,N_4888);
and U6619 (N_6619,N_3309,N_2910);
nand U6620 (N_6620,N_4147,N_4130);
xor U6621 (N_6621,N_4161,N_4406);
or U6622 (N_6622,N_3087,N_4444);
or U6623 (N_6623,N_4339,N_3869);
and U6624 (N_6624,N_2632,N_3590);
xor U6625 (N_6625,N_3648,N_2985);
nor U6626 (N_6626,N_3788,N_2830);
nor U6627 (N_6627,N_3898,N_3431);
xnor U6628 (N_6628,N_3701,N_3475);
or U6629 (N_6629,N_3755,N_2659);
nor U6630 (N_6630,N_3079,N_3534);
or U6631 (N_6631,N_3272,N_2558);
xor U6632 (N_6632,N_2648,N_4652);
or U6633 (N_6633,N_3933,N_3384);
or U6634 (N_6634,N_4681,N_4867);
and U6635 (N_6635,N_4145,N_4510);
and U6636 (N_6636,N_3013,N_3305);
or U6637 (N_6637,N_2820,N_4964);
nand U6638 (N_6638,N_4501,N_3761);
nand U6639 (N_6639,N_4830,N_3841);
or U6640 (N_6640,N_3317,N_3583);
or U6641 (N_6641,N_4555,N_4715);
nor U6642 (N_6642,N_4579,N_3943);
nor U6643 (N_6643,N_2745,N_4174);
nand U6644 (N_6644,N_3282,N_3583);
and U6645 (N_6645,N_4290,N_3921);
nand U6646 (N_6646,N_4138,N_4346);
nor U6647 (N_6647,N_3137,N_3984);
nand U6648 (N_6648,N_2721,N_4848);
nand U6649 (N_6649,N_2533,N_2542);
and U6650 (N_6650,N_3231,N_3653);
nor U6651 (N_6651,N_3915,N_2528);
or U6652 (N_6652,N_2679,N_3544);
nor U6653 (N_6653,N_3373,N_3929);
or U6654 (N_6654,N_3233,N_4579);
nor U6655 (N_6655,N_4660,N_4383);
or U6656 (N_6656,N_4447,N_3541);
nor U6657 (N_6657,N_4342,N_2629);
xor U6658 (N_6658,N_4909,N_4651);
xnor U6659 (N_6659,N_3022,N_2788);
nor U6660 (N_6660,N_3782,N_3082);
nand U6661 (N_6661,N_4448,N_3090);
xor U6662 (N_6662,N_3761,N_4261);
nand U6663 (N_6663,N_4537,N_4979);
and U6664 (N_6664,N_3301,N_4999);
nor U6665 (N_6665,N_3208,N_2743);
nor U6666 (N_6666,N_4875,N_3176);
and U6667 (N_6667,N_4262,N_2813);
nand U6668 (N_6668,N_3008,N_3324);
xnor U6669 (N_6669,N_4695,N_3206);
nor U6670 (N_6670,N_3720,N_3196);
nor U6671 (N_6671,N_4515,N_3894);
nand U6672 (N_6672,N_2672,N_4800);
xnor U6673 (N_6673,N_3422,N_2551);
and U6674 (N_6674,N_3316,N_3584);
and U6675 (N_6675,N_3029,N_4601);
and U6676 (N_6676,N_4625,N_3918);
nor U6677 (N_6677,N_3523,N_4520);
xnor U6678 (N_6678,N_4150,N_4414);
nor U6679 (N_6679,N_3443,N_3976);
nand U6680 (N_6680,N_4140,N_2970);
or U6681 (N_6681,N_2829,N_4328);
or U6682 (N_6682,N_3366,N_4308);
or U6683 (N_6683,N_3921,N_4252);
or U6684 (N_6684,N_4254,N_4941);
nor U6685 (N_6685,N_4642,N_3333);
or U6686 (N_6686,N_3609,N_4017);
or U6687 (N_6687,N_3422,N_3855);
nand U6688 (N_6688,N_2918,N_2795);
and U6689 (N_6689,N_2833,N_3988);
nand U6690 (N_6690,N_4402,N_3619);
nor U6691 (N_6691,N_3617,N_3972);
xor U6692 (N_6692,N_3032,N_3293);
or U6693 (N_6693,N_3995,N_4254);
nor U6694 (N_6694,N_3427,N_3106);
and U6695 (N_6695,N_4689,N_4979);
and U6696 (N_6696,N_3334,N_4353);
nor U6697 (N_6697,N_2680,N_3698);
nor U6698 (N_6698,N_3554,N_4670);
xnor U6699 (N_6699,N_3079,N_2501);
nor U6700 (N_6700,N_4683,N_3639);
or U6701 (N_6701,N_4707,N_4228);
and U6702 (N_6702,N_3702,N_4560);
and U6703 (N_6703,N_3491,N_3432);
and U6704 (N_6704,N_3911,N_4324);
and U6705 (N_6705,N_4230,N_3597);
or U6706 (N_6706,N_2743,N_4681);
or U6707 (N_6707,N_3196,N_3570);
nand U6708 (N_6708,N_4345,N_3360);
nor U6709 (N_6709,N_4712,N_2571);
xor U6710 (N_6710,N_3388,N_4483);
nor U6711 (N_6711,N_3719,N_4971);
or U6712 (N_6712,N_4397,N_3172);
and U6713 (N_6713,N_3538,N_3324);
or U6714 (N_6714,N_3548,N_4942);
and U6715 (N_6715,N_4913,N_4348);
and U6716 (N_6716,N_4082,N_3713);
nor U6717 (N_6717,N_2597,N_4842);
nor U6718 (N_6718,N_2981,N_4576);
xnor U6719 (N_6719,N_4033,N_3494);
nand U6720 (N_6720,N_3691,N_3081);
nor U6721 (N_6721,N_2637,N_2765);
nor U6722 (N_6722,N_4515,N_4977);
nand U6723 (N_6723,N_2574,N_3750);
and U6724 (N_6724,N_3911,N_3715);
or U6725 (N_6725,N_3533,N_2537);
nand U6726 (N_6726,N_4991,N_3726);
xor U6727 (N_6727,N_4431,N_2588);
xor U6728 (N_6728,N_4729,N_4997);
and U6729 (N_6729,N_3091,N_2866);
nand U6730 (N_6730,N_3626,N_2880);
xnor U6731 (N_6731,N_2741,N_4806);
nor U6732 (N_6732,N_3495,N_3040);
xor U6733 (N_6733,N_3891,N_4445);
nor U6734 (N_6734,N_4663,N_4095);
or U6735 (N_6735,N_3735,N_3955);
nand U6736 (N_6736,N_2531,N_2749);
or U6737 (N_6737,N_4764,N_3518);
or U6738 (N_6738,N_4611,N_3496);
nor U6739 (N_6739,N_4780,N_2553);
nand U6740 (N_6740,N_3584,N_4250);
nor U6741 (N_6741,N_2906,N_4354);
xnor U6742 (N_6742,N_4242,N_2516);
nand U6743 (N_6743,N_4274,N_3327);
or U6744 (N_6744,N_3201,N_3985);
nand U6745 (N_6745,N_4248,N_4316);
nand U6746 (N_6746,N_3465,N_3039);
xor U6747 (N_6747,N_3176,N_3761);
and U6748 (N_6748,N_3682,N_4369);
xor U6749 (N_6749,N_3027,N_3070);
nor U6750 (N_6750,N_3086,N_3739);
nor U6751 (N_6751,N_2874,N_3824);
xor U6752 (N_6752,N_2554,N_4170);
nand U6753 (N_6753,N_3900,N_2648);
and U6754 (N_6754,N_4999,N_4577);
or U6755 (N_6755,N_3169,N_2945);
and U6756 (N_6756,N_3717,N_3185);
nor U6757 (N_6757,N_2713,N_3972);
xor U6758 (N_6758,N_4931,N_4395);
nor U6759 (N_6759,N_3101,N_4483);
xnor U6760 (N_6760,N_4169,N_4978);
nor U6761 (N_6761,N_2860,N_4217);
or U6762 (N_6762,N_4706,N_3573);
xnor U6763 (N_6763,N_2558,N_3134);
xor U6764 (N_6764,N_4537,N_3358);
and U6765 (N_6765,N_3048,N_2708);
or U6766 (N_6766,N_3204,N_4068);
or U6767 (N_6767,N_4625,N_4195);
nor U6768 (N_6768,N_2857,N_3741);
and U6769 (N_6769,N_4202,N_2811);
nor U6770 (N_6770,N_3237,N_4609);
or U6771 (N_6771,N_3400,N_4886);
xor U6772 (N_6772,N_3125,N_2602);
or U6773 (N_6773,N_3775,N_3406);
nand U6774 (N_6774,N_4508,N_3865);
and U6775 (N_6775,N_4577,N_3042);
and U6776 (N_6776,N_2866,N_4815);
nor U6777 (N_6777,N_3825,N_3984);
nand U6778 (N_6778,N_3122,N_2568);
nor U6779 (N_6779,N_4939,N_3892);
xor U6780 (N_6780,N_3477,N_4957);
nand U6781 (N_6781,N_3846,N_3500);
or U6782 (N_6782,N_3040,N_4737);
and U6783 (N_6783,N_3030,N_2815);
or U6784 (N_6784,N_3721,N_2509);
or U6785 (N_6785,N_3887,N_3014);
nand U6786 (N_6786,N_2832,N_2587);
xnor U6787 (N_6787,N_4844,N_4760);
nor U6788 (N_6788,N_3086,N_2621);
or U6789 (N_6789,N_2816,N_3081);
nor U6790 (N_6790,N_4620,N_3303);
nand U6791 (N_6791,N_3957,N_4307);
or U6792 (N_6792,N_3046,N_4216);
and U6793 (N_6793,N_3580,N_4930);
nor U6794 (N_6794,N_2583,N_3551);
xor U6795 (N_6795,N_4209,N_2689);
xnor U6796 (N_6796,N_3725,N_3822);
nor U6797 (N_6797,N_3126,N_4795);
and U6798 (N_6798,N_3439,N_4557);
and U6799 (N_6799,N_2848,N_4223);
xnor U6800 (N_6800,N_2792,N_4166);
or U6801 (N_6801,N_4432,N_2651);
or U6802 (N_6802,N_2951,N_4892);
nand U6803 (N_6803,N_3072,N_3985);
nand U6804 (N_6804,N_4932,N_4672);
xnor U6805 (N_6805,N_4411,N_3002);
or U6806 (N_6806,N_3360,N_3975);
and U6807 (N_6807,N_3840,N_4407);
or U6808 (N_6808,N_2900,N_4131);
or U6809 (N_6809,N_4855,N_4232);
and U6810 (N_6810,N_4454,N_3035);
nor U6811 (N_6811,N_3895,N_2920);
nand U6812 (N_6812,N_4982,N_3932);
nand U6813 (N_6813,N_4951,N_2749);
xnor U6814 (N_6814,N_3813,N_3581);
or U6815 (N_6815,N_2763,N_4070);
xnor U6816 (N_6816,N_3978,N_4676);
and U6817 (N_6817,N_4123,N_4744);
xnor U6818 (N_6818,N_2821,N_3995);
or U6819 (N_6819,N_4115,N_2531);
or U6820 (N_6820,N_2804,N_2551);
nand U6821 (N_6821,N_2886,N_4070);
xnor U6822 (N_6822,N_4890,N_3697);
nand U6823 (N_6823,N_4795,N_2611);
or U6824 (N_6824,N_3010,N_4431);
or U6825 (N_6825,N_3289,N_2749);
and U6826 (N_6826,N_2540,N_4813);
nor U6827 (N_6827,N_3953,N_3525);
or U6828 (N_6828,N_2501,N_4293);
nor U6829 (N_6829,N_3964,N_4952);
and U6830 (N_6830,N_3333,N_2683);
nand U6831 (N_6831,N_3765,N_4544);
or U6832 (N_6832,N_2687,N_2834);
nand U6833 (N_6833,N_4575,N_4045);
nor U6834 (N_6834,N_4668,N_2808);
and U6835 (N_6835,N_4206,N_3758);
or U6836 (N_6836,N_3301,N_4640);
nand U6837 (N_6837,N_3201,N_4747);
nand U6838 (N_6838,N_4107,N_4478);
and U6839 (N_6839,N_4422,N_2649);
and U6840 (N_6840,N_4093,N_4082);
nand U6841 (N_6841,N_3560,N_4245);
or U6842 (N_6842,N_4072,N_3525);
xnor U6843 (N_6843,N_4439,N_3635);
or U6844 (N_6844,N_3239,N_3803);
and U6845 (N_6845,N_2983,N_4453);
nor U6846 (N_6846,N_4402,N_4542);
nand U6847 (N_6847,N_2910,N_4148);
xor U6848 (N_6848,N_4926,N_4170);
xnor U6849 (N_6849,N_3246,N_4345);
xor U6850 (N_6850,N_4224,N_4847);
and U6851 (N_6851,N_3392,N_2966);
and U6852 (N_6852,N_2943,N_3076);
nor U6853 (N_6853,N_2599,N_3892);
nor U6854 (N_6854,N_3854,N_4264);
xor U6855 (N_6855,N_4892,N_3560);
nor U6856 (N_6856,N_3821,N_4892);
or U6857 (N_6857,N_3909,N_3989);
and U6858 (N_6858,N_3413,N_3562);
nor U6859 (N_6859,N_3430,N_3451);
xnor U6860 (N_6860,N_4142,N_3049);
nor U6861 (N_6861,N_4927,N_3981);
and U6862 (N_6862,N_3978,N_4256);
and U6863 (N_6863,N_3715,N_4659);
or U6864 (N_6864,N_3412,N_3071);
or U6865 (N_6865,N_3184,N_4713);
nor U6866 (N_6866,N_3096,N_4308);
nand U6867 (N_6867,N_2836,N_4078);
xor U6868 (N_6868,N_4136,N_3619);
and U6869 (N_6869,N_4731,N_3276);
nor U6870 (N_6870,N_4871,N_3548);
xnor U6871 (N_6871,N_4812,N_3770);
nor U6872 (N_6872,N_2778,N_4056);
and U6873 (N_6873,N_4050,N_3514);
nor U6874 (N_6874,N_3081,N_4492);
xnor U6875 (N_6875,N_3742,N_4587);
nand U6876 (N_6876,N_4248,N_2543);
xnor U6877 (N_6877,N_4348,N_4102);
or U6878 (N_6878,N_3179,N_3471);
nor U6879 (N_6879,N_4263,N_4541);
and U6880 (N_6880,N_4775,N_2556);
or U6881 (N_6881,N_3122,N_4265);
nor U6882 (N_6882,N_3853,N_4667);
and U6883 (N_6883,N_4589,N_3713);
or U6884 (N_6884,N_4767,N_4639);
nor U6885 (N_6885,N_4205,N_4852);
nor U6886 (N_6886,N_4853,N_2813);
nand U6887 (N_6887,N_4711,N_4425);
nor U6888 (N_6888,N_3807,N_3087);
nand U6889 (N_6889,N_4184,N_4104);
nand U6890 (N_6890,N_2539,N_3406);
nor U6891 (N_6891,N_3448,N_4064);
nand U6892 (N_6892,N_3623,N_4468);
or U6893 (N_6893,N_3331,N_4074);
or U6894 (N_6894,N_3582,N_4158);
or U6895 (N_6895,N_3914,N_3403);
and U6896 (N_6896,N_3500,N_3892);
nand U6897 (N_6897,N_3653,N_2896);
or U6898 (N_6898,N_3412,N_3851);
or U6899 (N_6899,N_3367,N_4362);
xor U6900 (N_6900,N_3378,N_3571);
or U6901 (N_6901,N_4027,N_4778);
nand U6902 (N_6902,N_4846,N_2799);
or U6903 (N_6903,N_4455,N_4388);
xnor U6904 (N_6904,N_4276,N_4093);
nor U6905 (N_6905,N_4592,N_2964);
nor U6906 (N_6906,N_4740,N_4590);
nand U6907 (N_6907,N_2783,N_2774);
nor U6908 (N_6908,N_3415,N_3163);
nand U6909 (N_6909,N_4541,N_3256);
and U6910 (N_6910,N_2748,N_4608);
nor U6911 (N_6911,N_4348,N_4111);
xor U6912 (N_6912,N_3896,N_2765);
and U6913 (N_6913,N_2532,N_3233);
nand U6914 (N_6914,N_3046,N_3809);
and U6915 (N_6915,N_4506,N_3864);
or U6916 (N_6916,N_3053,N_4141);
or U6917 (N_6917,N_3445,N_4154);
nand U6918 (N_6918,N_4438,N_2990);
xnor U6919 (N_6919,N_3539,N_3593);
nand U6920 (N_6920,N_4112,N_4508);
nor U6921 (N_6921,N_4387,N_4965);
xnor U6922 (N_6922,N_4397,N_4561);
nand U6923 (N_6923,N_4218,N_2923);
nand U6924 (N_6924,N_4592,N_3113);
and U6925 (N_6925,N_4551,N_4316);
nand U6926 (N_6926,N_3026,N_3551);
nand U6927 (N_6927,N_4483,N_2525);
nand U6928 (N_6928,N_4640,N_3019);
xnor U6929 (N_6929,N_2506,N_3916);
nor U6930 (N_6930,N_2891,N_4715);
nand U6931 (N_6931,N_4144,N_4707);
nand U6932 (N_6932,N_3120,N_2562);
xnor U6933 (N_6933,N_3764,N_4923);
nor U6934 (N_6934,N_4880,N_4273);
and U6935 (N_6935,N_4417,N_3757);
or U6936 (N_6936,N_3134,N_2817);
and U6937 (N_6937,N_3348,N_3932);
nor U6938 (N_6938,N_4845,N_4274);
nand U6939 (N_6939,N_3928,N_4869);
and U6940 (N_6940,N_4209,N_3311);
and U6941 (N_6941,N_3662,N_4886);
nand U6942 (N_6942,N_2849,N_4040);
nor U6943 (N_6943,N_4634,N_4973);
and U6944 (N_6944,N_3284,N_3070);
nor U6945 (N_6945,N_4665,N_4758);
nor U6946 (N_6946,N_4478,N_3077);
and U6947 (N_6947,N_4731,N_3868);
and U6948 (N_6948,N_3437,N_3306);
xnor U6949 (N_6949,N_2563,N_4753);
or U6950 (N_6950,N_2933,N_4965);
nor U6951 (N_6951,N_4729,N_2703);
xnor U6952 (N_6952,N_4789,N_2745);
or U6953 (N_6953,N_3400,N_2522);
and U6954 (N_6954,N_2815,N_4041);
xor U6955 (N_6955,N_4868,N_4654);
nor U6956 (N_6956,N_4483,N_3769);
or U6957 (N_6957,N_3972,N_4498);
or U6958 (N_6958,N_4708,N_4720);
and U6959 (N_6959,N_4065,N_2757);
and U6960 (N_6960,N_4067,N_3452);
nor U6961 (N_6961,N_4195,N_4075);
and U6962 (N_6962,N_3214,N_3560);
or U6963 (N_6963,N_4874,N_4050);
nand U6964 (N_6964,N_2895,N_3639);
xor U6965 (N_6965,N_2889,N_4117);
nand U6966 (N_6966,N_4801,N_4755);
nand U6967 (N_6967,N_4883,N_3956);
xor U6968 (N_6968,N_4222,N_3355);
nor U6969 (N_6969,N_4489,N_3405);
nor U6970 (N_6970,N_4633,N_3859);
xor U6971 (N_6971,N_3046,N_3715);
xor U6972 (N_6972,N_2534,N_4438);
nor U6973 (N_6973,N_4146,N_4750);
nand U6974 (N_6974,N_3573,N_4657);
or U6975 (N_6975,N_4673,N_4379);
or U6976 (N_6976,N_3808,N_4580);
xnor U6977 (N_6977,N_4138,N_2747);
xnor U6978 (N_6978,N_4530,N_4510);
and U6979 (N_6979,N_4043,N_3670);
nand U6980 (N_6980,N_4626,N_3970);
xnor U6981 (N_6981,N_4028,N_3496);
and U6982 (N_6982,N_3289,N_3537);
or U6983 (N_6983,N_3395,N_3595);
nor U6984 (N_6984,N_3660,N_3925);
xnor U6985 (N_6985,N_2631,N_3589);
nor U6986 (N_6986,N_3360,N_3350);
or U6987 (N_6987,N_3129,N_4353);
and U6988 (N_6988,N_4671,N_4839);
nor U6989 (N_6989,N_3764,N_3783);
xor U6990 (N_6990,N_4615,N_3239);
nand U6991 (N_6991,N_4377,N_4384);
or U6992 (N_6992,N_3622,N_2915);
xor U6993 (N_6993,N_3477,N_2944);
or U6994 (N_6994,N_3539,N_4630);
nor U6995 (N_6995,N_4101,N_2910);
nor U6996 (N_6996,N_4369,N_3880);
or U6997 (N_6997,N_2898,N_2975);
nor U6998 (N_6998,N_2575,N_3862);
nor U6999 (N_6999,N_3902,N_4590);
nand U7000 (N_7000,N_4377,N_3731);
and U7001 (N_7001,N_4668,N_4415);
nand U7002 (N_7002,N_4919,N_2783);
xnor U7003 (N_7003,N_3491,N_3380);
nand U7004 (N_7004,N_3930,N_2978);
and U7005 (N_7005,N_3849,N_3474);
nand U7006 (N_7006,N_4177,N_4015);
nand U7007 (N_7007,N_4437,N_4541);
and U7008 (N_7008,N_2726,N_3860);
or U7009 (N_7009,N_2747,N_3636);
nor U7010 (N_7010,N_4977,N_4857);
or U7011 (N_7011,N_3304,N_4439);
or U7012 (N_7012,N_4850,N_4346);
and U7013 (N_7013,N_3151,N_4649);
or U7014 (N_7014,N_3381,N_4014);
xor U7015 (N_7015,N_2604,N_3526);
xnor U7016 (N_7016,N_4031,N_4976);
nor U7017 (N_7017,N_4210,N_4850);
and U7018 (N_7018,N_3104,N_3125);
or U7019 (N_7019,N_4258,N_2699);
nand U7020 (N_7020,N_2509,N_4415);
or U7021 (N_7021,N_4257,N_3699);
nand U7022 (N_7022,N_3002,N_2635);
and U7023 (N_7023,N_2602,N_2784);
nor U7024 (N_7024,N_3828,N_4957);
nand U7025 (N_7025,N_3420,N_4659);
xor U7026 (N_7026,N_2597,N_3810);
or U7027 (N_7027,N_4742,N_3590);
nand U7028 (N_7028,N_3834,N_3682);
nand U7029 (N_7029,N_2789,N_3304);
or U7030 (N_7030,N_4269,N_3885);
nor U7031 (N_7031,N_3637,N_3764);
nor U7032 (N_7032,N_4979,N_4856);
or U7033 (N_7033,N_2768,N_4623);
xnor U7034 (N_7034,N_3924,N_2958);
or U7035 (N_7035,N_4305,N_4282);
or U7036 (N_7036,N_3061,N_4203);
and U7037 (N_7037,N_4193,N_3048);
xor U7038 (N_7038,N_3678,N_3991);
nand U7039 (N_7039,N_3292,N_4057);
nand U7040 (N_7040,N_3810,N_2796);
nor U7041 (N_7041,N_2685,N_4519);
nand U7042 (N_7042,N_2640,N_4812);
xnor U7043 (N_7043,N_3488,N_4293);
nor U7044 (N_7044,N_3339,N_3200);
xnor U7045 (N_7045,N_4960,N_4419);
xnor U7046 (N_7046,N_3945,N_4169);
or U7047 (N_7047,N_4572,N_4999);
or U7048 (N_7048,N_3926,N_2695);
nor U7049 (N_7049,N_2622,N_2636);
nand U7050 (N_7050,N_3612,N_4587);
nand U7051 (N_7051,N_3569,N_2745);
nand U7052 (N_7052,N_4385,N_2747);
or U7053 (N_7053,N_4837,N_4510);
and U7054 (N_7054,N_4460,N_3564);
and U7055 (N_7055,N_4990,N_4246);
or U7056 (N_7056,N_3919,N_4728);
xor U7057 (N_7057,N_4032,N_4108);
nand U7058 (N_7058,N_4424,N_4103);
or U7059 (N_7059,N_4856,N_4553);
or U7060 (N_7060,N_4467,N_4669);
nor U7061 (N_7061,N_3807,N_3879);
or U7062 (N_7062,N_2980,N_4729);
xnor U7063 (N_7063,N_3614,N_4698);
or U7064 (N_7064,N_2590,N_2847);
xnor U7065 (N_7065,N_4961,N_4972);
or U7066 (N_7066,N_4921,N_4818);
xnor U7067 (N_7067,N_4849,N_2955);
xor U7068 (N_7068,N_3678,N_3516);
nor U7069 (N_7069,N_4302,N_2711);
nor U7070 (N_7070,N_3694,N_4908);
nand U7071 (N_7071,N_3328,N_2511);
and U7072 (N_7072,N_3792,N_4080);
nand U7073 (N_7073,N_3548,N_4515);
or U7074 (N_7074,N_2847,N_2929);
and U7075 (N_7075,N_4157,N_3318);
and U7076 (N_7076,N_3917,N_4586);
and U7077 (N_7077,N_3021,N_4305);
and U7078 (N_7078,N_2591,N_4074);
or U7079 (N_7079,N_3139,N_3369);
or U7080 (N_7080,N_3598,N_3202);
xor U7081 (N_7081,N_3199,N_2744);
nand U7082 (N_7082,N_2883,N_3483);
and U7083 (N_7083,N_3483,N_2905);
nand U7084 (N_7084,N_4782,N_3466);
nand U7085 (N_7085,N_4308,N_2788);
nor U7086 (N_7086,N_3718,N_3733);
nor U7087 (N_7087,N_4673,N_4479);
nor U7088 (N_7088,N_2973,N_4527);
and U7089 (N_7089,N_4615,N_3849);
xor U7090 (N_7090,N_4390,N_2503);
nor U7091 (N_7091,N_4351,N_3445);
or U7092 (N_7092,N_4097,N_4886);
nor U7093 (N_7093,N_3535,N_2677);
nand U7094 (N_7094,N_4367,N_3003);
xor U7095 (N_7095,N_4455,N_3137);
and U7096 (N_7096,N_2726,N_4051);
xnor U7097 (N_7097,N_4078,N_4498);
nand U7098 (N_7098,N_4258,N_3794);
or U7099 (N_7099,N_4830,N_3917);
xnor U7100 (N_7100,N_4107,N_3109);
xnor U7101 (N_7101,N_4270,N_4224);
or U7102 (N_7102,N_2667,N_2844);
and U7103 (N_7103,N_3168,N_4455);
or U7104 (N_7104,N_4502,N_3200);
nand U7105 (N_7105,N_3775,N_4596);
xnor U7106 (N_7106,N_4303,N_4213);
or U7107 (N_7107,N_2857,N_4049);
nand U7108 (N_7108,N_3549,N_3061);
nand U7109 (N_7109,N_3022,N_3030);
nor U7110 (N_7110,N_4742,N_4825);
or U7111 (N_7111,N_2959,N_4859);
and U7112 (N_7112,N_2779,N_3095);
and U7113 (N_7113,N_4776,N_2531);
nor U7114 (N_7114,N_4089,N_2791);
nand U7115 (N_7115,N_3662,N_4210);
nor U7116 (N_7116,N_3487,N_4553);
nor U7117 (N_7117,N_3098,N_4623);
xor U7118 (N_7118,N_3013,N_4872);
nor U7119 (N_7119,N_3934,N_4485);
or U7120 (N_7120,N_3854,N_4777);
nor U7121 (N_7121,N_2510,N_4800);
and U7122 (N_7122,N_3594,N_4915);
or U7123 (N_7123,N_4647,N_3073);
and U7124 (N_7124,N_4656,N_4661);
xor U7125 (N_7125,N_4701,N_3974);
nand U7126 (N_7126,N_4266,N_2632);
nor U7127 (N_7127,N_4396,N_3635);
nand U7128 (N_7128,N_3213,N_2863);
or U7129 (N_7129,N_3107,N_2711);
or U7130 (N_7130,N_4406,N_4334);
nand U7131 (N_7131,N_2710,N_2969);
or U7132 (N_7132,N_3206,N_3742);
nor U7133 (N_7133,N_4426,N_2856);
nand U7134 (N_7134,N_2509,N_3470);
nand U7135 (N_7135,N_4520,N_2795);
and U7136 (N_7136,N_3276,N_2990);
nand U7137 (N_7137,N_3007,N_4421);
nand U7138 (N_7138,N_3373,N_2857);
nand U7139 (N_7139,N_3899,N_3339);
nor U7140 (N_7140,N_4977,N_4108);
xnor U7141 (N_7141,N_4784,N_4516);
and U7142 (N_7142,N_3410,N_3251);
or U7143 (N_7143,N_3615,N_2530);
nor U7144 (N_7144,N_4274,N_2836);
and U7145 (N_7145,N_3672,N_3985);
nor U7146 (N_7146,N_3392,N_4230);
nand U7147 (N_7147,N_3465,N_4779);
nand U7148 (N_7148,N_4759,N_4187);
and U7149 (N_7149,N_4447,N_4486);
nor U7150 (N_7150,N_4532,N_4215);
or U7151 (N_7151,N_4946,N_4554);
and U7152 (N_7152,N_4576,N_4978);
nand U7153 (N_7153,N_3612,N_3171);
or U7154 (N_7154,N_2582,N_2519);
and U7155 (N_7155,N_4519,N_3921);
xnor U7156 (N_7156,N_4174,N_3607);
and U7157 (N_7157,N_2933,N_3916);
and U7158 (N_7158,N_2750,N_3830);
nor U7159 (N_7159,N_4301,N_3656);
nor U7160 (N_7160,N_2633,N_3984);
nor U7161 (N_7161,N_2791,N_2954);
nand U7162 (N_7162,N_4631,N_2643);
nor U7163 (N_7163,N_4751,N_3483);
or U7164 (N_7164,N_4316,N_3300);
nand U7165 (N_7165,N_4874,N_3047);
and U7166 (N_7166,N_4576,N_4991);
and U7167 (N_7167,N_4065,N_4400);
xnor U7168 (N_7168,N_3201,N_3082);
nor U7169 (N_7169,N_4120,N_4310);
and U7170 (N_7170,N_3914,N_4131);
nor U7171 (N_7171,N_2997,N_4768);
xor U7172 (N_7172,N_2829,N_3262);
or U7173 (N_7173,N_4895,N_3136);
xor U7174 (N_7174,N_2656,N_3371);
or U7175 (N_7175,N_2657,N_2769);
and U7176 (N_7176,N_4687,N_4587);
nand U7177 (N_7177,N_2696,N_4738);
nand U7178 (N_7178,N_4443,N_2713);
and U7179 (N_7179,N_4439,N_4333);
and U7180 (N_7180,N_2749,N_2694);
or U7181 (N_7181,N_3540,N_4546);
xnor U7182 (N_7182,N_4652,N_2562);
nand U7183 (N_7183,N_3625,N_3476);
xnor U7184 (N_7184,N_3977,N_4081);
xnor U7185 (N_7185,N_4901,N_3608);
and U7186 (N_7186,N_4974,N_4925);
xnor U7187 (N_7187,N_4429,N_4455);
nor U7188 (N_7188,N_4743,N_3480);
nor U7189 (N_7189,N_4622,N_4086);
and U7190 (N_7190,N_4387,N_3264);
nand U7191 (N_7191,N_4673,N_4894);
nor U7192 (N_7192,N_3910,N_4874);
nor U7193 (N_7193,N_4532,N_3776);
and U7194 (N_7194,N_4387,N_3386);
xnor U7195 (N_7195,N_2896,N_4511);
nand U7196 (N_7196,N_3513,N_4516);
nor U7197 (N_7197,N_4123,N_4519);
or U7198 (N_7198,N_4837,N_3954);
nand U7199 (N_7199,N_2792,N_2638);
nand U7200 (N_7200,N_4532,N_3229);
or U7201 (N_7201,N_4658,N_4135);
and U7202 (N_7202,N_3156,N_4550);
and U7203 (N_7203,N_3528,N_4692);
nand U7204 (N_7204,N_4096,N_4424);
and U7205 (N_7205,N_3670,N_4782);
and U7206 (N_7206,N_3625,N_3456);
and U7207 (N_7207,N_3503,N_2521);
nand U7208 (N_7208,N_4804,N_3675);
nor U7209 (N_7209,N_3179,N_3546);
nand U7210 (N_7210,N_3806,N_2834);
nand U7211 (N_7211,N_3408,N_2520);
and U7212 (N_7212,N_3483,N_3324);
nand U7213 (N_7213,N_3976,N_4312);
nand U7214 (N_7214,N_4470,N_4522);
nand U7215 (N_7215,N_2540,N_2597);
or U7216 (N_7216,N_3449,N_2874);
nand U7217 (N_7217,N_4684,N_4607);
nor U7218 (N_7218,N_4452,N_4993);
or U7219 (N_7219,N_4926,N_3995);
xor U7220 (N_7220,N_4915,N_2752);
xnor U7221 (N_7221,N_3648,N_3021);
nand U7222 (N_7222,N_3293,N_3323);
nor U7223 (N_7223,N_4993,N_4827);
and U7224 (N_7224,N_2873,N_3013);
xnor U7225 (N_7225,N_4573,N_4176);
nor U7226 (N_7226,N_3572,N_2996);
or U7227 (N_7227,N_3482,N_3170);
nand U7228 (N_7228,N_4057,N_3542);
nor U7229 (N_7229,N_3552,N_2708);
xor U7230 (N_7230,N_3644,N_4062);
nand U7231 (N_7231,N_3427,N_4191);
nor U7232 (N_7232,N_3061,N_2788);
or U7233 (N_7233,N_4766,N_2589);
and U7234 (N_7234,N_3347,N_4369);
xor U7235 (N_7235,N_4275,N_4099);
nand U7236 (N_7236,N_2557,N_3215);
and U7237 (N_7237,N_2790,N_4316);
nand U7238 (N_7238,N_2880,N_3865);
and U7239 (N_7239,N_4569,N_3786);
nand U7240 (N_7240,N_2752,N_2626);
and U7241 (N_7241,N_3250,N_3507);
nand U7242 (N_7242,N_4684,N_4579);
nand U7243 (N_7243,N_3274,N_4808);
or U7244 (N_7244,N_4884,N_3165);
and U7245 (N_7245,N_2996,N_2659);
xor U7246 (N_7246,N_4121,N_3133);
xnor U7247 (N_7247,N_3400,N_3750);
xor U7248 (N_7248,N_3199,N_3687);
xnor U7249 (N_7249,N_2874,N_3559);
xor U7250 (N_7250,N_4262,N_3736);
or U7251 (N_7251,N_2920,N_2939);
nand U7252 (N_7252,N_3472,N_3622);
nor U7253 (N_7253,N_2983,N_2633);
xor U7254 (N_7254,N_3830,N_2993);
or U7255 (N_7255,N_3749,N_3168);
nor U7256 (N_7256,N_3644,N_3035);
nand U7257 (N_7257,N_3792,N_4531);
xor U7258 (N_7258,N_4888,N_3379);
nor U7259 (N_7259,N_4464,N_3095);
nand U7260 (N_7260,N_4515,N_2655);
xor U7261 (N_7261,N_3522,N_4866);
xor U7262 (N_7262,N_4966,N_4244);
and U7263 (N_7263,N_3785,N_2977);
and U7264 (N_7264,N_3740,N_4678);
nor U7265 (N_7265,N_4206,N_2534);
nor U7266 (N_7266,N_3587,N_4763);
or U7267 (N_7267,N_4295,N_4801);
nor U7268 (N_7268,N_4617,N_2701);
xor U7269 (N_7269,N_4696,N_2589);
nor U7270 (N_7270,N_4727,N_4134);
and U7271 (N_7271,N_3100,N_4104);
and U7272 (N_7272,N_3167,N_3089);
and U7273 (N_7273,N_3864,N_4887);
or U7274 (N_7274,N_4487,N_4840);
nand U7275 (N_7275,N_4010,N_2914);
nor U7276 (N_7276,N_4944,N_2603);
nand U7277 (N_7277,N_3074,N_2734);
and U7278 (N_7278,N_3135,N_4103);
xor U7279 (N_7279,N_4410,N_4203);
or U7280 (N_7280,N_3911,N_3806);
and U7281 (N_7281,N_2932,N_4258);
nor U7282 (N_7282,N_3983,N_3131);
nand U7283 (N_7283,N_3836,N_2917);
and U7284 (N_7284,N_4980,N_3610);
nand U7285 (N_7285,N_4224,N_3784);
and U7286 (N_7286,N_4656,N_3176);
nand U7287 (N_7287,N_4895,N_2627);
or U7288 (N_7288,N_2762,N_3053);
and U7289 (N_7289,N_3424,N_4992);
nand U7290 (N_7290,N_4792,N_4381);
xor U7291 (N_7291,N_4951,N_3805);
or U7292 (N_7292,N_4072,N_4441);
nand U7293 (N_7293,N_4517,N_3272);
nor U7294 (N_7294,N_4824,N_4252);
and U7295 (N_7295,N_3240,N_4645);
nand U7296 (N_7296,N_3216,N_4388);
or U7297 (N_7297,N_4573,N_4253);
and U7298 (N_7298,N_3443,N_4292);
nor U7299 (N_7299,N_4918,N_3860);
nand U7300 (N_7300,N_3698,N_2972);
nor U7301 (N_7301,N_3417,N_3697);
nor U7302 (N_7302,N_3178,N_4267);
nor U7303 (N_7303,N_2681,N_3204);
nand U7304 (N_7304,N_4403,N_3024);
nand U7305 (N_7305,N_3122,N_4834);
or U7306 (N_7306,N_4916,N_3355);
and U7307 (N_7307,N_4062,N_3896);
nand U7308 (N_7308,N_4823,N_3764);
nor U7309 (N_7309,N_3524,N_3120);
or U7310 (N_7310,N_4977,N_4571);
or U7311 (N_7311,N_2894,N_2609);
and U7312 (N_7312,N_2957,N_4713);
nand U7313 (N_7313,N_2951,N_4494);
nor U7314 (N_7314,N_3615,N_3908);
and U7315 (N_7315,N_3182,N_4224);
nand U7316 (N_7316,N_4672,N_3071);
xnor U7317 (N_7317,N_2650,N_4943);
xor U7318 (N_7318,N_3113,N_3796);
and U7319 (N_7319,N_3090,N_3152);
and U7320 (N_7320,N_4347,N_3080);
nor U7321 (N_7321,N_3959,N_4151);
or U7322 (N_7322,N_2891,N_3839);
nor U7323 (N_7323,N_4025,N_4451);
and U7324 (N_7324,N_3632,N_3199);
or U7325 (N_7325,N_2630,N_2818);
nor U7326 (N_7326,N_2955,N_3305);
nor U7327 (N_7327,N_3781,N_2689);
or U7328 (N_7328,N_3863,N_4111);
nand U7329 (N_7329,N_2503,N_3376);
and U7330 (N_7330,N_3429,N_4675);
or U7331 (N_7331,N_4297,N_4601);
or U7332 (N_7332,N_4039,N_3672);
nor U7333 (N_7333,N_3049,N_3091);
xor U7334 (N_7334,N_3401,N_2905);
nand U7335 (N_7335,N_4169,N_4985);
xor U7336 (N_7336,N_3060,N_3307);
and U7337 (N_7337,N_3504,N_4864);
and U7338 (N_7338,N_3516,N_3300);
or U7339 (N_7339,N_3303,N_4767);
xnor U7340 (N_7340,N_4655,N_4385);
and U7341 (N_7341,N_2502,N_3587);
nor U7342 (N_7342,N_3859,N_4161);
nor U7343 (N_7343,N_4568,N_4075);
and U7344 (N_7344,N_3327,N_3804);
xnor U7345 (N_7345,N_3645,N_2536);
or U7346 (N_7346,N_4244,N_3534);
nor U7347 (N_7347,N_3420,N_4459);
nor U7348 (N_7348,N_3709,N_3628);
nor U7349 (N_7349,N_3613,N_4392);
nor U7350 (N_7350,N_3148,N_2629);
xor U7351 (N_7351,N_4932,N_3630);
or U7352 (N_7352,N_3339,N_4110);
xnor U7353 (N_7353,N_2826,N_2847);
nor U7354 (N_7354,N_3583,N_2782);
nor U7355 (N_7355,N_4097,N_3479);
nand U7356 (N_7356,N_4787,N_3358);
or U7357 (N_7357,N_2975,N_3796);
nand U7358 (N_7358,N_3838,N_4611);
and U7359 (N_7359,N_3619,N_4274);
or U7360 (N_7360,N_3806,N_2675);
xnor U7361 (N_7361,N_3684,N_4444);
nor U7362 (N_7362,N_3239,N_4498);
xor U7363 (N_7363,N_3474,N_4532);
or U7364 (N_7364,N_4889,N_4091);
nor U7365 (N_7365,N_4515,N_3181);
nand U7366 (N_7366,N_4133,N_2906);
or U7367 (N_7367,N_3248,N_4865);
or U7368 (N_7368,N_3042,N_2861);
xor U7369 (N_7369,N_4377,N_4434);
nor U7370 (N_7370,N_4168,N_2859);
nor U7371 (N_7371,N_4902,N_2818);
xor U7372 (N_7372,N_4244,N_4137);
nand U7373 (N_7373,N_3795,N_3011);
or U7374 (N_7374,N_4418,N_3406);
xor U7375 (N_7375,N_3326,N_4809);
or U7376 (N_7376,N_3604,N_3219);
or U7377 (N_7377,N_4671,N_2816);
nor U7378 (N_7378,N_2566,N_3167);
and U7379 (N_7379,N_3645,N_3726);
or U7380 (N_7380,N_4644,N_2637);
nand U7381 (N_7381,N_3181,N_4737);
or U7382 (N_7382,N_3001,N_3617);
and U7383 (N_7383,N_3372,N_3785);
nand U7384 (N_7384,N_2586,N_3207);
nor U7385 (N_7385,N_2935,N_3898);
and U7386 (N_7386,N_3400,N_3730);
xnor U7387 (N_7387,N_4498,N_3989);
nand U7388 (N_7388,N_4010,N_4074);
nor U7389 (N_7389,N_3692,N_3752);
or U7390 (N_7390,N_4533,N_3261);
xor U7391 (N_7391,N_2769,N_3678);
nand U7392 (N_7392,N_3346,N_3617);
and U7393 (N_7393,N_4053,N_4402);
nor U7394 (N_7394,N_3787,N_4638);
and U7395 (N_7395,N_4890,N_3785);
nor U7396 (N_7396,N_4153,N_3616);
xnor U7397 (N_7397,N_3683,N_4010);
and U7398 (N_7398,N_3608,N_3420);
nor U7399 (N_7399,N_2821,N_2720);
nor U7400 (N_7400,N_3833,N_2932);
nor U7401 (N_7401,N_2940,N_2794);
nor U7402 (N_7402,N_3900,N_3448);
xor U7403 (N_7403,N_4375,N_2586);
nand U7404 (N_7404,N_3458,N_4394);
or U7405 (N_7405,N_4189,N_4527);
xnor U7406 (N_7406,N_4771,N_2644);
nor U7407 (N_7407,N_4907,N_4407);
nor U7408 (N_7408,N_2905,N_3276);
or U7409 (N_7409,N_2556,N_3929);
or U7410 (N_7410,N_2906,N_3381);
xnor U7411 (N_7411,N_4393,N_4242);
or U7412 (N_7412,N_4276,N_3262);
and U7413 (N_7413,N_4328,N_4024);
or U7414 (N_7414,N_2621,N_4725);
nor U7415 (N_7415,N_4467,N_4278);
or U7416 (N_7416,N_3397,N_3780);
nand U7417 (N_7417,N_4089,N_4227);
xor U7418 (N_7418,N_2518,N_4484);
xnor U7419 (N_7419,N_4661,N_3787);
nor U7420 (N_7420,N_3440,N_2686);
nor U7421 (N_7421,N_2784,N_4757);
nor U7422 (N_7422,N_3860,N_3461);
or U7423 (N_7423,N_2939,N_3002);
nand U7424 (N_7424,N_4067,N_4954);
nor U7425 (N_7425,N_4426,N_2632);
nor U7426 (N_7426,N_3634,N_2979);
and U7427 (N_7427,N_4764,N_3565);
xor U7428 (N_7428,N_3623,N_4019);
and U7429 (N_7429,N_3907,N_2868);
nand U7430 (N_7430,N_4435,N_3329);
nand U7431 (N_7431,N_3224,N_4803);
and U7432 (N_7432,N_4701,N_4733);
or U7433 (N_7433,N_3151,N_4038);
and U7434 (N_7434,N_3313,N_3915);
nand U7435 (N_7435,N_4147,N_2878);
or U7436 (N_7436,N_4481,N_4459);
and U7437 (N_7437,N_4014,N_3939);
and U7438 (N_7438,N_3183,N_4258);
nand U7439 (N_7439,N_4687,N_3230);
or U7440 (N_7440,N_3810,N_4468);
and U7441 (N_7441,N_3113,N_4929);
and U7442 (N_7442,N_4428,N_3487);
xnor U7443 (N_7443,N_2698,N_3474);
or U7444 (N_7444,N_2952,N_3763);
nor U7445 (N_7445,N_3515,N_3815);
xnor U7446 (N_7446,N_3174,N_2752);
or U7447 (N_7447,N_3350,N_4085);
nor U7448 (N_7448,N_4724,N_3924);
xnor U7449 (N_7449,N_4669,N_4106);
nand U7450 (N_7450,N_4114,N_3040);
nand U7451 (N_7451,N_4333,N_3006);
and U7452 (N_7452,N_3613,N_2638);
xor U7453 (N_7453,N_4490,N_4003);
xnor U7454 (N_7454,N_4609,N_4173);
nand U7455 (N_7455,N_4691,N_2940);
nand U7456 (N_7456,N_2542,N_2630);
nand U7457 (N_7457,N_2689,N_4237);
xor U7458 (N_7458,N_3445,N_4880);
nand U7459 (N_7459,N_3700,N_3093);
xnor U7460 (N_7460,N_2689,N_2748);
xnor U7461 (N_7461,N_4315,N_4508);
and U7462 (N_7462,N_4020,N_2633);
nor U7463 (N_7463,N_2852,N_2782);
and U7464 (N_7464,N_2809,N_3831);
nor U7465 (N_7465,N_3037,N_4182);
nor U7466 (N_7466,N_3576,N_2756);
nand U7467 (N_7467,N_2534,N_3086);
nand U7468 (N_7468,N_4461,N_3082);
nand U7469 (N_7469,N_4096,N_3720);
or U7470 (N_7470,N_2714,N_2835);
or U7471 (N_7471,N_4418,N_4839);
and U7472 (N_7472,N_4644,N_4189);
and U7473 (N_7473,N_3130,N_4411);
and U7474 (N_7474,N_3053,N_4902);
xnor U7475 (N_7475,N_4293,N_3103);
nor U7476 (N_7476,N_3719,N_2733);
and U7477 (N_7477,N_3197,N_4931);
and U7478 (N_7478,N_3977,N_4296);
nor U7479 (N_7479,N_3567,N_3451);
xnor U7480 (N_7480,N_4652,N_4821);
or U7481 (N_7481,N_4349,N_3599);
and U7482 (N_7482,N_4661,N_3693);
xor U7483 (N_7483,N_2862,N_3742);
nand U7484 (N_7484,N_3161,N_4941);
xnor U7485 (N_7485,N_4117,N_2674);
xnor U7486 (N_7486,N_4640,N_4454);
or U7487 (N_7487,N_4151,N_4895);
and U7488 (N_7488,N_4901,N_4062);
or U7489 (N_7489,N_3551,N_2927);
nor U7490 (N_7490,N_2517,N_3686);
and U7491 (N_7491,N_3667,N_3526);
or U7492 (N_7492,N_3230,N_3958);
nand U7493 (N_7493,N_3026,N_4800);
nor U7494 (N_7494,N_3315,N_4269);
nand U7495 (N_7495,N_3548,N_4339);
nand U7496 (N_7496,N_3908,N_4471);
nand U7497 (N_7497,N_3102,N_3515);
nor U7498 (N_7498,N_2500,N_2590);
nand U7499 (N_7499,N_3570,N_3712);
and U7500 (N_7500,N_5240,N_5078);
or U7501 (N_7501,N_5480,N_6178);
and U7502 (N_7502,N_6078,N_6597);
nor U7503 (N_7503,N_6799,N_7334);
and U7504 (N_7504,N_6658,N_7364);
xnor U7505 (N_7505,N_6687,N_5247);
nand U7506 (N_7506,N_6720,N_6361);
and U7507 (N_7507,N_5146,N_5826);
or U7508 (N_7508,N_6647,N_5032);
nor U7509 (N_7509,N_5459,N_5035);
or U7510 (N_7510,N_6853,N_5984);
or U7511 (N_7511,N_5603,N_5132);
nor U7512 (N_7512,N_5847,N_6869);
and U7513 (N_7513,N_5817,N_6014);
nand U7514 (N_7514,N_7474,N_6313);
nand U7515 (N_7515,N_5675,N_6623);
nand U7516 (N_7516,N_6311,N_5574);
and U7517 (N_7517,N_6444,N_5181);
xnor U7518 (N_7518,N_7018,N_6914);
xnor U7519 (N_7519,N_6061,N_6490);
and U7520 (N_7520,N_5891,N_6447);
or U7521 (N_7521,N_6828,N_5430);
xor U7522 (N_7522,N_6166,N_6754);
xor U7523 (N_7523,N_5721,N_5207);
and U7524 (N_7524,N_6471,N_5183);
and U7525 (N_7525,N_6579,N_5606);
nand U7526 (N_7526,N_5732,N_6011);
nand U7527 (N_7527,N_6648,N_7313);
and U7528 (N_7528,N_6945,N_5698);
and U7529 (N_7529,N_6614,N_5338);
xnor U7530 (N_7530,N_7198,N_5953);
nor U7531 (N_7531,N_5941,N_5112);
nand U7532 (N_7532,N_5622,N_6775);
nand U7533 (N_7533,N_7010,N_5086);
xor U7534 (N_7534,N_5014,N_7082);
or U7535 (N_7535,N_5440,N_6719);
xnor U7536 (N_7536,N_5541,N_6610);
nor U7537 (N_7537,N_6947,N_6776);
nand U7538 (N_7538,N_6736,N_6628);
and U7539 (N_7539,N_5185,N_6894);
and U7540 (N_7540,N_6810,N_5040);
nand U7541 (N_7541,N_7051,N_5141);
or U7542 (N_7542,N_7077,N_7420);
nand U7543 (N_7543,N_5515,N_6511);
and U7544 (N_7544,N_6424,N_5643);
or U7545 (N_7545,N_6862,N_5798);
nor U7546 (N_7546,N_6352,N_7447);
and U7547 (N_7547,N_5224,N_6578);
xnor U7548 (N_7548,N_6861,N_6482);
xnor U7549 (N_7549,N_6452,N_5288);
nor U7550 (N_7550,N_5790,N_5463);
and U7551 (N_7551,N_6060,N_5432);
nor U7552 (N_7552,N_6333,N_5437);
xor U7553 (N_7553,N_5104,N_5627);
nand U7554 (N_7554,N_7112,N_5038);
nand U7555 (N_7555,N_5850,N_6065);
xnor U7556 (N_7556,N_6600,N_6241);
and U7557 (N_7557,N_6394,N_5692);
or U7558 (N_7558,N_6770,N_5951);
and U7559 (N_7559,N_5490,N_5879);
nor U7560 (N_7560,N_5514,N_5502);
xnor U7561 (N_7561,N_7205,N_6325);
and U7562 (N_7562,N_5042,N_5007);
or U7563 (N_7563,N_6027,N_5198);
nand U7564 (N_7564,N_7401,N_7029);
xor U7565 (N_7565,N_6278,N_5690);
or U7566 (N_7566,N_5592,N_6133);
nor U7567 (N_7567,N_6935,N_7282);
and U7568 (N_7568,N_5292,N_5378);
or U7569 (N_7569,N_6539,N_6239);
nor U7570 (N_7570,N_5680,N_5917);
and U7571 (N_7571,N_5899,N_5345);
nand U7572 (N_7572,N_5862,N_6070);
or U7573 (N_7573,N_5701,N_5749);
or U7574 (N_7574,N_6167,N_5666);
nand U7575 (N_7575,N_5838,N_5967);
and U7576 (N_7576,N_6906,N_5520);
nand U7577 (N_7577,N_7480,N_6707);
or U7578 (N_7578,N_5106,N_5272);
xor U7579 (N_7579,N_5614,N_5800);
xor U7580 (N_7580,N_7078,N_6415);
nor U7581 (N_7581,N_6972,N_7215);
and U7582 (N_7582,N_6222,N_7286);
and U7583 (N_7583,N_5852,N_5392);
and U7584 (N_7584,N_5560,N_5579);
xnor U7585 (N_7585,N_5725,N_6905);
nor U7586 (N_7586,N_6301,N_5221);
and U7587 (N_7587,N_6104,N_5789);
nand U7588 (N_7588,N_5179,N_5791);
and U7589 (N_7589,N_5889,N_7045);
nand U7590 (N_7590,N_7002,N_6435);
nand U7591 (N_7591,N_7415,N_6498);
nand U7592 (N_7592,N_7161,N_6635);
and U7593 (N_7593,N_6542,N_5534);
and U7594 (N_7594,N_6686,N_6083);
and U7595 (N_7595,N_6473,N_5408);
xnor U7596 (N_7596,N_5155,N_7394);
nand U7597 (N_7597,N_5704,N_7322);
nand U7598 (N_7598,N_7389,N_6870);
nor U7599 (N_7599,N_6378,N_6018);
xor U7600 (N_7600,N_5575,N_6981);
or U7601 (N_7601,N_5091,N_6533);
xor U7602 (N_7602,N_6187,N_5924);
nor U7603 (N_7603,N_6817,N_6238);
or U7604 (N_7604,N_5944,N_6149);
xnor U7605 (N_7605,N_7383,N_7009);
and U7606 (N_7606,N_5685,N_6886);
xnor U7607 (N_7607,N_5825,N_6348);
xnor U7608 (N_7608,N_5263,N_6266);
and U7609 (N_7609,N_7342,N_6345);
nor U7610 (N_7610,N_6038,N_7165);
xnor U7611 (N_7611,N_6946,N_6681);
xor U7612 (N_7612,N_5448,N_6064);
nor U7613 (N_7613,N_5878,N_6470);
nand U7614 (N_7614,N_6001,N_5369);
nand U7615 (N_7615,N_5312,N_7084);
nand U7616 (N_7616,N_7418,N_6331);
xor U7617 (N_7617,N_7092,N_6657);
or U7618 (N_7618,N_6612,N_6580);
and U7619 (N_7619,N_5943,N_7316);
nor U7620 (N_7620,N_6012,N_5691);
nand U7621 (N_7621,N_5773,N_6085);
or U7622 (N_7622,N_7042,N_5588);
nand U7623 (N_7623,N_6299,N_5180);
and U7624 (N_7624,N_5381,N_6552);
xnor U7625 (N_7625,N_5499,N_6044);
nand U7626 (N_7626,N_6765,N_5567);
xnor U7627 (N_7627,N_6440,N_6419);
xor U7628 (N_7628,N_5543,N_5730);
xnor U7629 (N_7629,N_5449,N_5111);
nor U7630 (N_7630,N_6743,N_6651);
and U7631 (N_7631,N_7168,N_6196);
nand U7632 (N_7632,N_5154,N_5920);
and U7633 (N_7633,N_5897,N_5079);
nand U7634 (N_7634,N_5297,N_6875);
xor U7635 (N_7635,N_5255,N_6640);
nand U7636 (N_7636,N_7232,N_7167);
xor U7637 (N_7637,N_6461,N_6901);
or U7638 (N_7638,N_6215,N_5200);
nand U7639 (N_7639,N_5022,N_5009);
or U7640 (N_7640,N_7169,N_6492);
nor U7641 (N_7641,N_7061,N_6460);
xnor U7642 (N_7642,N_6164,N_6667);
xnor U7643 (N_7643,N_6709,N_6092);
and U7644 (N_7644,N_7477,N_6293);
and U7645 (N_7645,N_6739,N_6129);
and U7646 (N_7646,N_5919,N_5768);
and U7647 (N_7647,N_6260,N_5625);
nand U7648 (N_7648,N_7271,N_6992);
nand U7649 (N_7649,N_5929,N_6317);
nand U7650 (N_7650,N_5143,N_5488);
nor U7651 (N_7651,N_5905,N_6087);
nor U7652 (N_7652,N_6140,N_6409);
and U7653 (N_7653,N_7210,N_5674);
nor U7654 (N_7654,N_5846,N_5815);
nor U7655 (N_7655,N_6637,N_7201);
nand U7656 (N_7656,N_6483,N_7291);
or U7657 (N_7657,N_5849,N_7347);
and U7658 (N_7658,N_5393,N_5568);
xnor U7659 (N_7659,N_7498,N_6514);
or U7660 (N_7660,N_5248,N_6661);
nor U7661 (N_7661,N_6206,N_5452);
and U7662 (N_7662,N_5192,N_5736);
or U7663 (N_7663,N_5638,N_5851);
xnor U7664 (N_7664,N_6662,N_6019);
xor U7665 (N_7665,N_7369,N_5976);
and U7666 (N_7666,N_6631,N_7425);
xor U7667 (N_7667,N_6268,N_5257);
xor U7668 (N_7668,N_6724,N_6632);
xnor U7669 (N_7669,N_7093,N_6646);
or U7670 (N_7670,N_6931,N_6588);
nor U7671 (N_7671,N_5828,N_5202);
nor U7672 (N_7672,N_6226,N_7435);
or U7673 (N_7673,N_5306,N_6867);
xor U7674 (N_7674,N_7280,N_6969);
or U7675 (N_7675,N_5571,N_5716);
or U7676 (N_7676,N_7359,N_6571);
nor U7677 (N_7677,N_7381,N_7158);
or U7678 (N_7678,N_5114,N_5793);
nor U7679 (N_7679,N_5241,N_6798);
or U7680 (N_7680,N_5404,N_7059);
and U7681 (N_7681,N_7295,N_5819);
nor U7682 (N_7682,N_5486,N_6172);
nand U7683 (N_7683,N_5900,N_7033);
and U7684 (N_7684,N_6704,N_5485);
nand U7685 (N_7685,N_7008,N_6303);
and U7686 (N_7686,N_6948,N_6652);
or U7687 (N_7687,N_5761,N_5434);
or U7688 (N_7688,N_6357,N_7004);
xnor U7689 (N_7689,N_7318,N_6537);
nand U7690 (N_7690,N_7130,N_5478);
nor U7691 (N_7691,N_6413,N_5352);
and U7692 (N_7692,N_7106,N_5710);
nor U7693 (N_7693,N_5228,N_5150);
or U7694 (N_7694,N_5282,N_6634);
and U7695 (N_7695,N_5886,N_6996);
or U7696 (N_7696,N_5264,N_6041);
nor U7697 (N_7697,N_7341,N_5960);
and U7698 (N_7698,N_7235,N_6198);
nor U7699 (N_7699,N_5855,N_5890);
xor U7700 (N_7700,N_6699,N_5479);
xor U7701 (N_7701,N_6550,N_7174);
nor U7702 (N_7702,N_6145,N_5649);
nor U7703 (N_7703,N_5333,N_7413);
nor U7704 (N_7704,N_5232,N_6814);
or U7705 (N_7705,N_7240,N_6718);
nor U7706 (N_7706,N_6581,N_5363);
xor U7707 (N_7707,N_7258,N_5623);
and U7708 (N_7708,N_5617,N_6385);
nor U7709 (N_7709,N_5885,N_6845);
and U7710 (N_7710,N_6941,N_6095);
and U7711 (N_7711,N_6319,N_6355);
nor U7712 (N_7712,N_5682,N_5677);
or U7713 (N_7713,N_6146,N_5137);
xnor U7714 (N_7714,N_6349,N_6998);
xnor U7715 (N_7715,N_5597,N_7265);
xor U7716 (N_7716,N_5291,N_5027);
nor U7717 (N_7717,N_7261,N_6072);
and U7718 (N_7718,N_6157,N_6747);
or U7719 (N_7719,N_5555,N_6836);
or U7720 (N_7720,N_5050,N_5006);
xor U7721 (N_7721,N_6639,N_6389);
xnor U7722 (N_7722,N_7197,N_6118);
or U7723 (N_7723,N_5407,N_5085);
or U7724 (N_7724,N_6520,N_7113);
xor U7725 (N_7725,N_5750,N_7285);
nand U7726 (N_7726,N_6541,N_5746);
xor U7727 (N_7727,N_6984,N_6208);
and U7728 (N_7728,N_6150,N_6749);
nand U7729 (N_7729,N_6857,N_6493);
nand U7730 (N_7730,N_6567,N_6315);
or U7731 (N_7731,N_5536,N_6242);
nand U7732 (N_7732,N_5005,N_5896);
and U7733 (N_7733,N_5071,N_6171);
xor U7734 (N_7734,N_5045,N_6259);
nor U7735 (N_7735,N_7151,N_6621);
nor U7736 (N_7736,N_5503,N_6456);
and U7737 (N_7737,N_6575,N_5498);
or U7738 (N_7738,N_6964,N_6427);
or U7739 (N_7739,N_5388,N_5330);
nand U7740 (N_7740,N_6577,N_6695);
nand U7741 (N_7741,N_5599,N_7283);
or U7742 (N_7742,N_5636,N_5344);
xor U7743 (N_7743,N_5375,N_6841);
nand U7744 (N_7744,N_5081,N_6730);
or U7745 (N_7745,N_5445,N_5537);
nand U7746 (N_7746,N_7214,N_6391);
or U7747 (N_7747,N_5476,N_5783);
xor U7748 (N_7748,N_5218,N_6199);
nand U7749 (N_7749,N_5780,N_5804);
or U7750 (N_7750,N_7392,N_5201);
xnor U7751 (N_7751,N_6101,N_6849);
nand U7752 (N_7752,N_5808,N_7148);
xnor U7753 (N_7753,N_7387,N_6457);
or U7754 (N_7754,N_5493,N_5546);
xnor U7755 (N_7755,N_5915,N_5420);
nor U7756 (N_7756,N_5892,N_6446);
and U7757 (N_7757,N_6590,N_7350);
nand U7758 (N_7758,N_7136,N_6740);
xor U7759 (N_7759,N_5837,N_7451);
xor U7760 (N_7760,N_5424,N_5191);
xnor U7761 (N_7761,N_5147,N_6844);
nor U7762 (N_7762,N_6365,N_6069);
nor U7763 (N_7763,N_5940,N_5661);
or U7764 (N_7764,N_6077,N_5170);
and U7765 (N_7765,N_6891,N_5428);
nand U7766 (N_7766,N_6183,N_5733);
nor U7767 (N_7767,N_5065,N_6053);
nor U7768 (N_7768,N_6054,N_6030);
nor U7769 (N_7769,N_5051,N_6497);
and U7770 (N_7770,N_5914,N_5694);
or U7771 (N_7771,N_6816,N_5765);
nand U7772 (N_7772,N_5993,N_5932);
nor U7773 (N_7773,N_6418,N_6887);
or U7774 (N_7774,N_6965,N_6910);
and U7775 (N_7775,N_5261,N_6000);
xnor U7776 (N_7776,N_7453,N_7122);
nand U7777 (N_7777,N_5021,N_6458);
nor U7778 (N_7778,N_6063,N_6442);
nor U7779 (N_7779,N_5665,N_6881);
and U7780 (N_7780,N_6915,N_5570);
nand U7781 (N_7781,N_7249,N_5922);
xnor U7782 (N_7782,N_5801,N_5830);
nand U7783 (N_7783,N_6341,N_7123);
nor U7784 (N_7784,N_6494,N_6024);
xor U7785 (N_7785,N_6288,N_7360);
and U7786 (N_7786,N_5296,N_5545);
or U7787 (N_7787,N_7058,N_5087);
nand U7788 (N_7788,N_5167,N_5707);
and U7789 (N_7789,N_7098,N_5620);
xnor U7790 (N_7790,N_5171,N_7175);
nand U7791 (N_7791,N_7468,N_5279);
and U7792 (N_7792,N_7200,N_5672);
and U7793 (N_7793,N_5758,N_6032);
or U7794 (N_7794,N_5057,N_5662);
or U7795 (N_7795,N_6245,N_6067);
nand U7796 (N_7796,N_5702,N_6263);
nand U7797 (N_7797,N_6475,N_6777);
nor U7798 (N_7798,N_5429,N_6512);
xor U7799 (N_7799,N_7353,N_5512);
or U7800 (N_7800,N_5466,N_6694);
nor U7801 (N_7801,N_6793,N_5398);
nor U7802 (N_7802,N_6269,N_7374);
nor U7803 (N_7803,N_7053,N_6322);
and U7804 (N_7804,N_5641,N_5196);
and U7805 (N_7805,N_6161,N_5874);
nand U7806 (N_7806,N_6256,N_6821);
nand U7807 (N_7807,N_5958,N_7020);
or U7808 (N_7808,N_6794,N_6144);
nand U7809 (N_7809,N_5797,N_6752);
nor U7810 (N_7810,N_6273,N_5551);
xor U7811 (N_7811,N_6109,N_6673);
and U7812 (N_7812,N_6679,N_6976);
nand U7813 (N_7813,N_6139,N_7340);
xor U7814 (N_7814,N_5645,N_6827);
xnor U7815 (N_7815,N_7223,N_6207);
and U7816 (N_7816,N_5305,N_5002);
nand U7817 (N_7817,N_7162,N_5860);
nor U7818 (N_7818,N_6243,N_6688);
or U7819 (N_7819,N_6383,N_6464);
or U7820 (N_7820,N_7372,N_6582);
or U7821 (N_7821,N_6509,N_6429);
nor U7822 (N_7822,N_6443,N_5177);
or U7823 (N_7823,N_5577,N_7027);
and U7824 (N_7824,N_6832,N_5562);
nand U7825 (N_7825,N_6526,N_5843);
nor U7826 (N_7826,N_6717,N_7022);
nand U7827 (N_7827,N_5640,N_6500);
and U7828 (N_7828,N_6570,N_5903);
nand U7829 (N_7829,N_7450,N_6059);
xnor U7830 (N_7830,N_5446,N_6592);
nor U7831 (N_7831,N_7041,N_6626);
or U7832 (N_7832,N_6264,N_6643);
and U7833 (N_7833,N_5161,N_6280);
nand U7834 (N_7834,N_5921,N_6835);
and U7835 (N_7835,N_5911,N_7190);
xor U7836 (N_7836,N_6585,N_5794);
xnor U7837 (N_7837,N_5611,N_6936);
or U7838 (N_7838,N_5098,N_6463);
nand U7839 (N_7839,N_7408,N_5217);
or U7840 (N_7840,N_6223,N_6422);
xnor U7841 (N_7841,N_5506,N_6017);
nand U7842 (N_7842,N_7325,N_5313);
nor U7843 (N_7843,N_6123,N_5744);
or U7844 (N_7844,N_5723,N_5916);
nor U7845 (N_7845,N_6397,N_6221);
nand U7846 (N_7846,N_6091,N_5714);
nand U7847 (N_7847,N_6818,N_5162);
nor U7848 (N_7848,N_6733,N_6979);
nand U7849 (N_7849,N_6831,N_6057);
nand U7850 (N_7850,N_7289,N_5693);
or U7851 (N_7851,N_7245,N_6854);
nor U7852 (N_7852,N_7102,N_7469);
nor U7853 (N_7853,N_7129,N_5739);
nor U7854 (N_7854,N_5280,N_6281);
nand U7855 (N_7855,N_5013,N_7107);
nor U7856 (N_7856,N_5148,N_6698);
and U7857 (N_7857,N_5365,N_5912);
or U7858 (N_7858,N_6165,N_6455);
nand U7859 (N_7859,N_6186,N_5678);
and U7860 (N_7860,N_6339,N_5947);
or U7861 (N_7861,N_6439,N_7090);
nand U7862 (N_7862,N_6741,N_5766);
xnor U7863 (N_7863,N_7308,N_5259);
or U7864 (N_7864,N_5602,N_6374);
nor U7865 (N_7865,N_5632,N_7026);
nand U7866 (N_7866,N_5304,N_7319);
nand U7867 (N_7867,N_5358,N_6154);
xor U7868 (N_7868,N_5708,N_6750);
or U7869 (N_7869,N_5600,N_5073);
or U7870 (N_7870,N_6595,N_5274);
or U7871 (N_7871,N_5067,N_6576);
or U7872 (N_7872,N_6748,N_5936);
nor U7873 (N_7873,N_6666,N_7448);
nand U7874 (N_7874,N_7035,N_6230);
or U7875 (N_7875,N_6672,N_6134);
nor U7876 (N_7876,N_5220,N_6195);
or U7877 (N_7877,N_7075,N_5684);
xnor U7878 (N_7878,N_5105,N_6504);
and U7879 (N_7879,N_7356,N_5556);
nor U7880 (N_7880,N_6400,N_7236);
and U7881 (N_7881,N_6217,N_7478);
or U7882 (N_7882,N_7095,N_6534);
nor U7883 (N_7883,N_7296,N_6346);
nand U7884 (N_7884,N_5120,N_5935);
nand U7885 (N_7885,N_5133,N_5583);
nand U7886 (N_7886,N_7428,N_5487);
and U7887 (N_7887,N_5858,N_6093);
nor U7888 (N_7888,N_6283,N_5028);
nor U7889 (N_7889,N_5511,N_6745);
nand U7890 (N_7890,N_6068,N_6035);
xor U7891 (N_7891,N_6958,N_7094);
and U7892 (N_7892,N_5368,N_5281);
or U7893 (N_7893,N_5841,N_5743);
or U7894 (N_7894,N_5954,N_5735);
or U7895 (N_7895,N_6220,N_7013);
and U7896 (N_7896,N_6496,N_5117);
nor U7897 (N_7897,N_5391,N_5656);
xor U7898 (N_7898,N_5380,N_7177);
nor U7899 (N_7899,N_5894,N_6908);
nand U7900 (N_7900,N_7231,N_5152);
and U7901 (N_7901,N_7463,N_6603);
nor U7902 (N_7902,N_5153,N_5979);
xor U7903 (N_7903,N_6432,N_6796);
nand U7904 (N_7904,N_6107,N_5811);
nand U7905 (N_7905,N_5823,N_6684);
or U7906 (N_7906,N_5456,N_7324);
or U7907 (N_7907,N_6983,N_7373);
and U7908 (N_7908,N_6729,N_5458);
xnor U7909 (N_7909,N_5945,N_6522);
xor U7910 (N_7910,N_6872,N_5003);
nor U7911 (N_7911,N_5024,N_5598);
and U7912 (N_7912,N_6434,N_5718);
nand U7913 (N_7913,N_7103,N_6602);
or U7914 (N_7914,N_7348,N_7088);
or U7915 (N_7915,N_5530,N_7157);
xor U7916 (N_7916,N_6121,N_6287);
nand U7917 (N_7917,N_6677,N_5670);
and U7918 (N_7918,N_6320,N_7208);
xor U7919 (N_7919,N_6994,N_7248);
or U7920 (N_7920,N_5531,N_6332);
or U7921 (N_7921,N_6433,N_7273);
nand U7922 (N_7922,N_7398,N_5564);
xor U7923 (N_7923,N_5354,N_7030);
xnor U7924 (N_7924,N_6888,N_6766);
nor U7925 (N_7925,N_6148,N_7142);
or U7926 (N_7926,N_7457,N_6188);
and U7927 (N_7927,N_5031,N_5273);
and U7928 (N_7928,N_6115,N_5854);
nand U7929 (N_7929,N_6804,N_5001);
or U7930 (N_7930,N_5245,N_5631);
nor U7931 (N_7931,N_5930,N_5887);
xor U7932 (N_7932,N_5127,N_5184);
and U7933 (N_7933,N_6555,N_6721);
nor U7934 (N_7934,N_5527,N_6561);
and U7935 (N_7935,N_5820,N_7386);
and U7936 (N_7936,N_6013,N_5433);
or U7937 (N_7937,N_5307,N_7227);
and U7938 (N_7938,N_6644,N_6386);
or U7939 (N_7939,N_5321,N_6535);
xnor U7940 (N_7940,N_5484,N_5438);
nand U7941 (N_7941,N_6760,N_6089);
and U7942 (N_7942,N_6650,N_5342);
nor U7943 (N_7943,N_6898,N_6584);
nor U7944 (N_7944,N_6531,N_7409);
or U7945 (N_7945,N_7105,N_5399);
or U7946 (N_7946,N_5635,N_6645);
xnor U7947 (N_7947,N_7349,N_7263);
nand U7948 (N_7948,N_5955,N_6402);
or U7949 (N_7949,N_7426,N_7109);
xor U7950 (N_7950,N_5443,N_6495);
nand U7951 (N_7951,N_7462,N_6384);
xnor U7952 (N_7952,N_5848,N_7040);
or U7953 (N_7953,N_7351,N_5346);
or U7954 (N_7954,N_6056,N_6523);
nor U7955 (N_7955,N_5151,N_5046);
nor U7956 (N_7956,N_5489,N_5060);
nor U7957 (N_7957,N_7065,N_6554);
nor U7958 (N_7958,N_7253,N_6708);
and U7959 (N_7959,N_5235,N_6949);
or U7960 (N_7960,N_5594,N_6978);
or U7961 (N_7961,N_5178,N_6237);
or U7962 (N_7962,N_7147,N_5083);
nor U7963 (N_7963,N_5999,N_7329);
or U7964 (N_7964,N_7133,N_5806);
and U7965 (N_7965,N_7320,N_6548);
nand U7966 (N_7966,N_6620,N_7001);
xnor U7967 (N_7967,N_5362,N_5927);
or U7968 (N_7968,N_6757,N_7417);
nor U7969 (N_7969,N_5318,N_7202);
xor U7970 (N_7970,N_6538,N_5351);
xnor U7971 (N_7971,N_5034,N_6885);
nand U7972 (N_7972,N_6758,N_6696);
or U7973 (N_7973,N_6131,N_6487);
nand U7974 (N_7974,N_5370,N_5441);
nand U7975 (N_7975,N_6850,N_5777);
or U7976 (N_7976,N_5576,N_5722);
xnor U7977 (N_7977,N_6606,N_6956);
nand U7978 (N_7978,N_5876,N_7073);
nand U7979 (N_7979,N_5019,N_5390);
nor U7980 (N_7980,N_6569,N_6051);
nor U7981 (N_7981,N_6848,N_5757);
nand U7982 (N_7982,N_7390,N_7070);
nand U7983 (N_7983,N_6290,N_5467);
nor U7984 (N_7984,N_6191,N_7276);
xor U7985 (N_7985,N_7052,N_7083);
or U7986 (N_7986,N_5518,N_5135);
xnor U7987 (N_7987,N_6182,N_5122);
and U7988 (N_7988,N_6480,N_7455);
nand U7989 (N_7989,N_6342,N_6501);
xor U7990 (N_7990,N_6882,N_6682);
and U7991 (N_7991,N_5158,N_6725);
nand U7992 (N_7992,N_5077,N_7309);
nand U7993 (N_7993,N_7327,N_7363);
or U7994 (N_7994,N_5172,N_6046);
nand U7995 (N_7995,N_7229,N_5047);
or U7996 (N_7996,N_6174,N_7159);
and U7997 (N_7997,N_5671,N_5497);
nor U7998 (N_7998,N_5738,N_5347);
xnor U7999 (N_7999,N_7191,N_6937);
nor U8000 (N_8000,N_5495,N_6006);
xor U8001 (N_8001,N_5108,N_5319);
nor U8002 (N_8002,N_5573,N_6358);
and U8003 (N_8003,N_5964,N_5910);
or U8004 (N_8004,N_6153,N_5267);
nor U8005 (N_8005,N_5422,N_5118);
nor U8006 (N_8006,N_5861,N_6021);
xor U8007 (N_8007,N_6627,N_6811);
xor U8008 (N_8008,N_7345,N_7422);
xnor U8009 (N_8009,N_5290,N_7126);
xor U8010 (N_8010,N_7330,N_5018);
and U8011 (N_8011,N_5471,N_6528);
nand U8012 (N_8012,N_5973,N_6876);
and U8013 (N_8013,N_6291,N_5096);
xor U8014 (N_8014,N_7486,N_5136);
or U8015 (N_8015,N_5295,N_6484);
or U8016 (N_8016,N_7423,N_5190);
or U8017 (N_8017,N_6669,N_5754);
and U8018 (N_8018,N_6363,N_6156);
xor U8019 (N_8019,N_6653,N_6170);
nand U8020 (N_8020,N_6852,N_6312);
or U8021 (N_8021,N_5385,N_6353);
nor U8022 (N_8022,N_5859,N_5097);
nor U8023 (N_8023,N_6993,N_7181);
and U8024 (N_8024,N_7185,N_6767);
nand U8025 (N_8025,N_7302,N_5772);
xnor U8026 (N_8026,N_6911,N_7139);
nand U8027 (N_8027,N_7049,N_6727);
nand U8028 (N_8028,N_5262,N_5074);
nor U8029 (N_8029,N_6202,N_6406);
xnor U8030 (N_8030,N_6343,N_5926);
or U8031 (N_8031,N_6874,N_6593);
or U8032 (N_8032,N_5873,N_7024);
nand U8033 (N_8033,N_6009,N_6200);
xnor U8034 (N_8034,N_7436,N_5011);
or U8035 (N_8035,N_5023,N_5881);
xor U8036 (N_8036,N_6184,N_6379);
nor U8037 (N_8037,N_5776,N_5872);
nand U8038 (N_8038,N_5030,N_6405);
nand U8039 (N_8039,N_7481,N_6556);
nor U8040 (N_8040,N_6102,N_5753);
nor U8041 (N_8041,N_6753,N_5308);
nor U8042 (N_8042,N_6448,N_6641);
nor U8043 (N_8043,N_5283,N_5668);
and U8044 (N_8044,N_5123,N_5769);
xnor U8045 (N_8045,N_5834,N_5316);
and U8046 (N_8046,N_5402,N_7449);
nand U8047 (N_8047,N_6809,N_7354);
xor U8048 (N_8048,N_7406,N_5453);
and U8049 (N_8049,N_6864,N_6671);
nand U8050 (N_8050,N_6205,N_7032);
xor U8051 (N_8051,N_5700,N_7252);
nand U8052 (N_8052,N_6713,N_6934);
nand U8053 (N_8053,N_6583,N_6163);
nor U8054 (N_8054,N_7267,N_6820);
nor U8055 (N_8055,N_5337,N_5286);
or U8056 (N_8056,N_7187,N_6963);
nor U8057 (N_8057,N_6968,N_6336);
and U8058 (N_8058,N_6604,N_5853);
nand U8059 (N_8059,N_5015,N_5741);
xnor U8060 (N_8060,N_6376,N_6565);
nand U8061 (N_8061,N_6568,N_6573);
or U8062 (N_8062,N_5566,N_5327);
xor U8063 (N_8063,N_6430,N_6834);
nor U8064 (N_8064,N_6950,N_6955);
nor U8065 (N_8065,N_7014,N_5687);
xor U8066 (N_8066,N_6801,N_6396);
and U8067 (N_8067,N_6168,N_5189);
or U8068 (N_8068,N_5893,N_5360);
or U8069 (N_8069,N_6253,N_6377);
and U8070 (N_8070,N_5957,N_5713);
nor U8071 (N_8071,N_5904,N_5813);
nor U8072 (N_8072,N_7300,N_7303);
or U8073 (N_8073,N_7414,N_6084);
and U8074 (N_8074,N_7338,N_7305);
xor U8075 (N_8075,N_6116,N_6476);
xnor U8076 (N_8076,N_7489,N_6823);
nor U8077 (N_8077,N_7424,N_7101);
or U8078 (N_8078,N_6633,N_5475);
xnor U8079 (N_8079,N_7421,N_6939);
nand U8080 (N_8080,N_6611,N_5372);
xnor U8081 (N_8081,N_6421,N_6249);
nand U8082 (N_8082,N_5004,N_5269);
nor U8083 (N_8083,N_7081,N_5651);
and U8084 (N_8084,N_5349,N_6197);
and U8085 (N_8085,N_6126,N_6251);
or U8086 (N_8086,N_6962,N_7301);
nor U8087 (N_8087,N_5516,N_6088);
nor U8088 (N_8088,N_5865,N_7079);
xnor U8089 (N_8089,N_6909,N_6926);
nor U8090 (N_8090,N_7054,N_5839);
or U8091 (N_8091,N_6052,N_6613);
xnor U8092 (N_8092,N_6925,N_5835);
nor U8093 (N_8093,N_6097,N_6960);
nand U8094 (N_8094,N_5985,N_6366);
and U8095 (N_8095,N_5238,N_6530);
nand U8096 (N_8096,N_6598,N_6007);
and U8097 (N_8097,N_5840,N_6833);
and U8098 (N_8098,N_6216,N_5986);
nor U8099 (N_8099,N_5130,N_5901);
and U8100 (N_8100,N_5165,N_7493);
nand U8101 (N_8101,N_5483,N_7396);
nand U8102 (N_8102,N_6381,N_5781);
nor U8103 (N_8103,N_6663,N_5863);
and U8104 (N_8104,N_5650,N_6340);
or U8105 (N_8105,N_7278,N_6545);
and U8106 (N_8106,N_5301,N_6773);
nor U8107 (N_8107,N_6927,N_6967);
nand U8108 (N_8108,N_6179,N_5585);
or U8109 (N_8109,N_5144,N_6112);
nand U8110 (N_8110,N_7256,N_6227);
nand U8111 (N_8111,N_6591,N_6023);
and U8112 (N_8112,N_7388,N_6108);
nor U8113 (N_8113,N_7459,N_7044);
or U8114 (N_8114,N_5175,N_6923);
or U8115 (N_8115,N_7180,N_5669);
nand U8116 (N_8116,N_5907,N_6791);
or U8117 (N_8117,N_6277,N_7172);
xnor U8118 (N_8118,N_7495,N_5523);
xnor U8119 (N_8119,N_6697,N_5582);
nor U8120 (N_8120,N_6670,N_5664);
and U8121 (N_8121,N_5084,N_5048);
or U8122 (N_8122,N_6270,N_6327);
nand U8123 (N_8123,N_7056,N_5580);
xnor U8124 (N_8124,N_6151,N_5663);
and U8125 (N_8125,N_7166,N_7404);
nand U8126 (N_8126,N_7154,N_6474);
xnor U8127 (N_8127,N_6090,N_7446);
and U8128 (N_8128,N_5204,N_7160);
or U8129 (N_8129,N_7357,N_5619);
xor U8130 (N_8130,N_7321,N_6615);
nand U8131 (N_8131,N_6587,N_6359);
nand U8132 (N_8132,N_7213,N_6125);
xor U8133 (N_8133,N_6877,N_7005);
xor U8134 (N_8134,N_6436,N_5717);
nor U8135 (N_8135,N_6505,N_6459);
or U8136 (N_8136,N_5983,N_6917);
and U8137 (N_8137,N_6491,N_5052);
or U8138 (N_8138,N_6176,N_6462);
nand U8139 (N_8139,N_7218,N_6654);
or U8140 (N_8140,N_6778,N_5090);
and U8141 (N_8141,N_7234,N_6141);
nor U8142 (N_8142,N_5187,N_6244);
or U8143 (N_8143,N_6020,N_6081);
nand U8144 (N_8144,N_6438,N_6629);
nor U8145 (N_8145,N_5616,N_5975);
and U8146 (N_8146,N_6307,N_6073);
or U8147 (N_8147,N_5212,N_5596);
or U8148 (N_8148,N_6408,N_5252);
and U8149 (N_8149,N_5223,N_6525);
xor U8150 (N_8150,N_5374,N_7186);
xnor U8151 (N_8151,N_7346,N_6944);
nor U8152 (N_8152,N_5246,N_6989);
nand U8153 (N_8153,N_6524,N_7437);
xor U8154 (N_8154,N_5549,N_5436);
xnor U8155 (N_8155,N_5822,N_6354);
nand U8156 (N_8156,N_5624,N_6536);
nand U8157 (N_8157,N_6656,N_6557);
nor U8158 (N_8158,N_5036,N_6508);
and U8159 (N_8159,N_7000,N_5626);
and U8160 (N_8160,N_5933,N_5550);
xor U8161 (N_8161,N_5720,N_6478);
or U8162 (N_8162,N_5630,N_5383);
nand U8163 (N_8163,N_6735,N_6812);
nor U8164 (N_8164,N_7391,N_7438);
and U8165 (N_8165,N_5044,N_7337);
xnor U8166 (N_8166,N_5419,N_5504);
nor U8167 (N_8167,N_5856,N_6272);
and U8168 (N_8168,N_6813,N_7494);
and U8169 (N_8169,N_6224,N_5329);
and U8170 (N_8170,N_7003,N_6417);
and U8171 (N_8171,N_6031,N_5734);
xnor U8172 (N_8172,N_5978,N_6761);
xnor U8173 (N_8173,N_7237,N_6544);
xnor U8174 (N_8174,N_5268,N_6043);
and U8175 (N_8175,N_7310,N_6294);
xnor U8176 (N_8176,N_6285,N_7226);
or U8177 (N_8177,N_6247,N_6840);
nand U8178 (N_8178,N_5188,N_5332);
xor U8179 (N_8179,N_7104,N_5561);
nand U8180 (N_8180,N_5379,N_6532);
nand U8181 (N_8181,N_5884,N_6305);
or U8182 (N_8182,N_7150,N_5174);
nor U8183 (N_8183,N_7471,N_6211);
nor U8184 (N_8184,N_5528,N_5948);
and U8185 (N_8185,N_6098,N_6399);
nor U8186 (N_8186,N_6586,N_5173);
nor U8187 (N_8187,N_6454,N_5965);
nand U8188 (N_8188,N_5145,N_7118);
nand U8189 (N_8189,N_6540,N_5140);
and U8190 (N_8190,N_6338,N_5206);
xor U8191 (N_8191,N_5870,N_7143);
nor U8192 (N_8192,N_5361,N_5075);
or U8193 (N_8193,N_6966,N_6130);
and U8194 (N_8194,N_5470,N_6004);
and U8195 (N_8195,N_6074,N_6971);
nand U8196 (N_8196,N_6010,N_7299);
nor U8197 (N_8197,N_6466,N_7488);
nor U8198 (N_8198,N_6806,N_6152);
nor U8199 (N_8199,N_5763,N_6372);
nand U8200 (N_8200,N_6080,N_7230);
and U8201 (N_8201,N_7272,N_5000);
nor U8202 (N_8202,N_5350,N_5389);
nand U8203 (N_8203,N_5737,N_5457);
nor U8204 (N_8204,N_7483,N_6257);
xor U8205 (N_8205,N_7221,N_7242);
or U8206 (N_8206,N_5938,N_5542);
nand U8207 (N_8207,N_5997,N_6795);
and U8208 (N_8208,N_7366,N_5230);
nor U8209 (N_8209,N_7343,N_5548);
xor U8210 (N_8210,N_6477,N_6860);
nor U8211 (N_8211,N_6797,N_7339);
or U8212 (N_8212,N_5505,N_7066);
and U8213 (N_8213,N_7490,N_5501);
and U8214 (N_8214,N_5110,N_5277);
xnor U8215 (N_8215,N_7097,N_7099);
and U8216 (N_8216,N_6425,N_5644);
xnor U8217 (N_8217,N_6467,N_6192);
nand U8218 (N_8218,N_6479,N_5877);
and U8219 (N_8219,N_5634,N_5256);
and U8220 (N_8220,N_5474,N_5186);
xor U8221 (N_8221,N_5807,N_5335);
nor U8222 (N_8222,N_7086,N_5121);
or U8223 (N_8223,N_5166,N_5234);
and U8224 (N_8224,N_6100,N_5655);
or U8225 (N_8225,N_5928,N_6660);
xnor U8226 (N_8226,N_6037,N_6529);
nand U8227 (N_8227,N_6298,N_7326);
or U8228 (N_8228,N_7377,N_6889);
nor U8229 (N_8229,N_5169,N_7456);
nor U8230 (N_8230,N_5119,N_5056);
xnor U8231 (N_8231,N_7336,N_6124);
or U8232 (N_8232,N_5082,N_6710);
and U8233 (N_8233,N_5591,N_5525);
nor U8234 (N_8234,N_7292,N_6481);
and U8235 (N_8235,N_5017,N_7491);
and U8236 (N_8236,N_7149,N_5454);
xor U8237 (N_8237,N_6772,N_7378);
nand U8238 (N_8238,N_6468,N_6572);
and U8239 (N_8239,N_5317,N_6465);
or U8240 (N_8240,N_6407,N_7277);
xnor U8241 (N_8241,N_5857,N_5227);
nor U8242 (N_8242,N_7188,N_7444);
nor U8243 (N_8243,N_6204,N_5260);
xor U8244 (N_8244,N_6275,N_7199);
or U8245 (N_8245,N_6132,N_6880);
or U8246 (N_8246,N_6049,N_6506);
xor U8247 (N_8247,N_6235,N_5088);
or U8248 (N_8248,N_5314,N_7011);
nand U8249 (N_8249,N_5689,N_5326);
nand U8250 (N_8250,N_7220,N_7379);
and U8251 (N_8251,N_6789,N_5522);
nand U8252 (N_8252,N_7071,N_5728);
or U8253 (N_8253,N_5996,N_7131);
xor U8254 (N_8254,N_6103,N_6856);
nand U8255 (N_8255,N_5831,N_5683);
nor U8256 (N_8256,N_5774,N_5779);
or U8257 (N_8257,N_5400,N_7304);
or U8258 (N_8258,N_7432,N_7499);
nand U8259 (N_8259,N_5214,N_6330);
nand U8260 (N_8260,N_6169,N_6304);
nor U8261 (N_8261,N_6712,N_5866);
nand U8262 (N_8262,N_5080,N_7487);
and U8263 (N_8263,N_5906,N_5987);
or U8264 (N_8264,N_7442,N_5657);
and U8265 (N_8265,N_5646,N_7087);
and U8266 (N_8266,N_5925,N_5258);
nand U8267 (N_8267,N_6560,N_6824);
nor U8268 (N_8268,N_5810,N_6624);
or U8269 (N_8269,N_5593,N_5331);
nor U8270 (N_8270,N_5756,N_6075);
and U8271 (N_8271,N_7333,N_6488);
or U8272 (N_8272,N_7194,N_7067);
nor U8273 (N_8273,N_7461,N_5293);
or U8274 (N_8274,N_5062,N_6071);
xnor U8275 (N_8275,N_7482,N_5195);
and U8276 (N_8276,N_5679,N_6693);
nor U8277 (N_8277,N_5557,N_7115);
nand U8278 (N_8278,N_5465,N_7247);
xnor U8279 (N_8279,N_6781,N_6426);
xor U8280 (N_8280,N_6904,N_5992);
nor U8281 (N_8281,N_7465,N_5210);
xnor U8282 (N_8282,N_5590,N_5845);
nor U8283 (N_8283,N_6016,N_7370);
and U8284 (N_8284,N_6158,N_7416);
and U8285 (N_8285,N_5395,N_5126);
and U8286 (N_8286,N_5029,N_6680);
nor U8287 (N_8287,N_6117,N_7120);
nand U8288 (N_8288,N_6472,N_7472);
nand U8289 (N_8289,N_7317,N_6147);
nand U8290 (N_8290,N_5160,N_5742);
nor U8291 (N_8291,N_5061,N_5802);
nand U8292 (N_8292,N_6995,N_7132);
xnor U8293 (N_8293,N_6261,N_5394);
nor U8294 (N_8294,N_5500,N_7192);
xnor U8295 (N_8295,N_5751,N_6838);
xor U8296 (N_8296,N_5752,N_5341);
xor U8297 (N_8297,N_6676,N_6751);
and U8298 (N_8298,N_5010,N_5770);
nor U8299 (N_8299,N_5068,N_5020);
nand U8300 (N_8300,N_7385,N_5219);
or U8301 (N_8301,N_5931,N_5468);
xor U8302 (N_8302,N_6918,N_5956);
xor U8303 (N_8303,N_5621,N_7266);
nand U8304 (N_8304,N_7074,N_7117);
nand U8305 (N_8305,N_6924,N_5524);
and U8306 (N_8306,N_7038,N_6047);
xnor U8307 (N_8307,N_6617,N_6212);
nor U8308 (N_8308,N_6855,N_5320);
xor U8309 (N_8309,N_7397,N_6279);
nand U8310 (N_8310,N_5159,N_6826);
and U8311 (N_8311,N_5427,N_6414);
nand U8312 (N_8312,N_7433,N_6382);
xnor U8313 (N_8313,N_5762,N_6066);
and U8314 (N_8314,N_5508,N_7100);
and U8315 (N_8315,N_6246,N_5788);
xnor U8316 (N_8316,N_7358,N_6871);
or U8317 (N_8317,N_5712,N_6829);
or U8318 (N_8318,N_6193,N_6289);
nor U8319 (N_8319,N_5197,N_6388);
nor U8320 (N_8320,N_6441,N_6058);
nand U8321 (N_8321,N_6691,N_6042);
nand U8322 (N_8322,N_6618,N_5637);
nor U8323 (N_8323,N_5315,N_7145);
nor U8324 (N_8324,N_5785,N_7312);
xnor U8325 (N_8325,N_6702,N_5517);
nand U8326 (N_8326,N_5658,N_6784);
or U8327 (N_8327,N_5008,N_5991);
nand U8328 (N_8328,N_5033,N_5942);
nor U8329 (N_8329,N_6563,N_7328);
xnor U8330 (N_8330,N_5667,N_5633);
or U8331 (N_8331,N_6449,N_6819);
or U8332 (N_8332,N_5719,N_6316);
or U8333 (N_8333,N_5431,N_6866);
and U8334 (N_8334,N_5760,N_6665);
or U8335 (N_8335,N_6254,N_6453);
nor U8336 (N_8336,N_7257,N_5653);
nor U8337 (N_8337,N_5055,N_5253);
nor U8338 (N_8338,N_7476,N_6907);
nand U8339 (N_8339,N_5792,N_5157);
xor U8340 (N_8340,N_5581,N_6689);
and U8341 (N_8341,N_7250,N_6685);
nor U8342 (N_8342,N_6711,N_7062);
nand U8343 (N_8343,N_5289,N_6203);
and U8344 (N_8344,N_5251,N_5447);
or U8345 (N_8345,N_5211,N_7050);
nor U8346 (N_8346,N_5284,N_7209);
and U8347 (N_8347,N_5799,N_5966);
nand U8348 (N_8348,N_6233,N_6683);
xor U8349 (N_8349,N_7176,N_5194);
and U8350 (N_8350,N_6997,N_5642);
xor U8351 (N_8351,N_6896,N_6344);
nor U8352 (N_8352,N_6609,N_6822);
nand U8353 (N_8353,N_5481,N_6973);
nand U8354 (N_8354,N_6040,N_5902);
xnor U8355 (N_8355,N_5908,N_6922);
and U8356 (N_8356,N_6335,N_6062);
nor U8357 (N_8357,N_5072,N_6589);
xor U8358 (N_8358,N_6744,N_5299);
nor U8359 (N_8359,N_5455,N_5242);
and U8360 (N_8360,N_7243,N_5748);
nand U8361 (N_8361,N_7270,N_7128);
or U8362 (N_8362,N_6553,N_6916);
xnor U8363 (N_8363,N_6034,N_5294);
or U8364 (N_8364,N_6786,N_5328);
nand U8365 (N_8365,N_6286,N_5139);
nor U8366 (N_8366,N_5923,N_6785);
nand U8367 (N_8367,N_5559,N_6005);
xor U8368 (N_8368,N_5376,N_5450);
nor U8369 (N_8369,N_6549,N_5521);
and U8370 (N_8370,N_6328,N_6362);
nor U8371 (N_8371,N_5439,N_6258);
nor U8372 (N_8372,N_6194,N_6334);
xnor U8373 (N_8373,N_7025,N_5101);
nor U8374 (N_8374,N_6029,N_5025);
nand U8375 (N_8375,N_6974,N_7344);
nand U8376 (N_8376,N_5681,N_7268);
and U8377 (N_8377,N_5589,N_5778);
xor U8378 (N_8378,N_6630,N_5477);
nor U8379 (N_8379,N_5939,N_6111);
nand U8380 (N_8380,N_5934,N_5364);
xnor U8381 (N_8381,N_5418,N_5974);
or U8382 (N_8382,N_7069,N_7043);
nor U8383 (N_8383,N_7055,N_6723);
or U8384 (N_8384,N_6985,N_5442);
nor U8385 (N_8385,N_7063,N_6390);
and U8386 (N_8386,N_5417,N_5544);
nand U8387 (N_8387,N_7259,N_5138);
and U8388 (N_8388,N_6306,N_5604);
and U8389 (N_8389,N_5715,N_7239);
xnor U8390 (N_8390,N_5586,N_5100);
or U8391 (N_8391,N_5384,N_5309);
nor U8392 (N_8392,N_6607,N_7238);
or U8393 (N_8393,N_6267,N_6879);
or U8394 (N_8394,N_6360,N_6039);
xor U8395 (N_8395,N_6295,N_6959);
or U8396 (N_8396,N_6201,N_7315);
nand U8397 (N_8397,N_7207,N_6351);
nor U8398 (N_8398,N_7367,N_5805);
xnor U8399 (N_8399,N_6510,N_7284);
and U8400 (N_8400,N_5982,N_5569);
xor U8401 (N_8401,N_5601,N_6137);
nor U8402 (N_8402,N_6551,N_6128);
nand U8403 (N_8403,N_6210,N_5287);
or U8404 (N_8404,N_5652,N_5740);
or U8405 (N_8405,N_5357,N_5883);
and U8406 (N_8406,N_5727,N_5969);
or U8407 (N_8407,N_7443,N_7125);
xnor U8408 (N_8408,N_5412,N_5089);
nor U8409 (N_8409,N_5539,N_6469);
nor U8410 (N_8410,N_5867,N_6250);
xnor U8411 (N_8411,N_7431,N_6746);
nand U8412 (N_8412,N_5659,N_6055);
xor U8413 (N_8413,N_6920,N_7173);
nor U8414 (N_8414,N_6213,N_6892);
nor U8415 (N_8415,N_5367,N_5697);
nand U8416 (N_8416,N_5012,N_6143);
nor U8417 (N_8417,N_6961,N_5711);
and U8418 (N_8418,N_5336,N_5970);
nor U8419 (N_8419,N_5968,N_6451);
xor U8420 (N_8420,N_7068,N_7048);
xnor U8421 (N_8421,N_6048,N_5509);
nand U8422 (N_8422,N_5216,N_6300);
or U8423 (N_8423,N_5871,N_6094);
or U8424 (N_8424,N_5994,N_7137);
nand U8425 (N_8425,N_6393,N_6282);
nand U8426 (N_8426,N_5037,N_5444);
xor U8427 (N_8427,N_7064,N_5724);
xnor U8428 (N_8428,N_5435,N_5298);
nor U8429 (N_8429,N_7110,N_5565);
nand U8430 (N_8430,N_6768,N_5472);
nand U8431 (N_8431,N_5998,N_7403);
and U8432 (N_8432,N_5249,N_6485);
nor U8433 (N_8433,N_5182,N_7430);
nand U8434 (N_8434,N_5699,N_6700);
nor U8435 (N_8435,N_7475,N_6218);
nor U8436 (N_8436,N_5377,N_7140);
xnor U8437 (N_8437,N_6705,N_5981);
and U8438 (N_8438,N_6297,N_7089);
xor U8439 (N_8439,N_5587,N_5386);
xnor U8440 (N_8440,N_5125,N_5213);
xnor U8441 (N_8441,N_5275,N_5824);
xnor U8442 (N_8442,N_6731,N_5116);
and U8443 (N_8443,N_7127,N_5821);
or U8444 (N_8444,N_5959,N_6347);
nor U8445 (N_8445,N_5696,N_5695);
xnor U8446 (N_8446,N_6050,N_6403);
or U8447 (N_8447,N_7178,N_5063);
xnor U8448 (N_8448,N_6815,N_5208);
nand U8449 (N_8449,N_5688,N_6987);
or U8450 (N_8450,N_7331,N_6232);
or U8451 (N_8451,N_5832,N_7323);
or U8452 (N_8452,N_6655,N_6574);
xor U8453 (N_8453,N_5913,N_7466);
or U8454 (N_8454,N_6392,N_6756);
xnor U8455 (N_8455,N_5254,N_5882);
nand U8456 (N_8456,N_5767,N_6373);
nor U8457 (N_8457,N_6225,N_6980);
nand U8458 (N_8458,N_5492,N_5946);
xnor U8459 (N_8459,N_7375,N_7204);
xnor U8460 (N_8460,N_5371,N_6701);
or U8461 (N_8461,N_5898,N_6437);
nor U8462 (N_8462,N_6977,N_7233);
nand U8463 (N_8463,N_5093,N_6431);
xnor U8464 (N_8464,N_5209,N_7380);
nor U8465 (N_8465,N_5199,N_6883);
nand U8466 (N_8466,N_7228,N_6113);
nand U8467 (N_8467,N_5413,N_6502);
and U8468 (N_8468,N_6732,N_7244);
and U8469 (N_8469,N_5836,N_7212);
xor U8470 (N_8470,N_5961,N_5373);
or U8471 (N_8471,N_5552,N_6668);
nor U8472 (N_8472,N_5532,N_6234);
nor U8473 (N_8473,N_6162,N_7384);
and U8474 (N_8474,N_6308,N_5405);
and U8475 (N_8475,N_5115,N_7407);
nand U8476 (N_8476,N_6755,N_7395);
xnor U8477 (N_8477,N_6942,N_6209);
nor U8478 (N_8478,N_5971,N_7287);
nor U8479 (N_8479,N_5237,N_5533);
xor U8480 (N_8480,N_6248,N_6715);
nand U8481 (N_8481,N_6897,N_6028);
nor U8482 (N_8482,N_6387,N_7179);
or U8483 (N_8483,N_5387,N_6240);
xnor U8484 (N_8484,N_5963,N_5425);
xor U8485 (N_8485,N_5782,N_7352);
xnor U8486 (N_8486,N_6564,N_6160);
xor U8487 (N_8487,N_7458,N_5977);
nand U8488 (N_8488,N_6830,N_5648);
or U8489 (N_8489,N_7307,N_5403);
and U8490 (N_8490,N_6728,N_6231);
and U8491 (N_8491,N_6135,N_5989);
nand U8492 (N_8492,N_6858,N_7402);
nand U8493 (N_8493,N_5990,N_7031);
nor U8494 (N_8494,N_6738,N_5787);
and U8495 (N_8495,N_6364,N_7023);
xnor U8496 (N_8496,N_6177,N_6136);
xnor U8497 (N_8497,N_6847,N_7060);
or U8498 (N_8498,N_5613,N_6499);
or U8499 (N_8499,N_5415,N_5039);
nand U8500 (N_8500,N_6703,N_5323);
xor U8501 (N_8501,N_5705,N_7368);
xnor U8502 (N_8502,N_7217,N_7410);
or U8503 (N_8503,N_7473,N_6086);
or U8504 (N_8504,N_6369,N_5410);
and U8505 (N_8505,N_6276,N_5382);
or U8506 (N_8506,N_6486,N_7189);
nand U8507 (N_8507,N_5066,N_7269);
or U8508 (N_8508,N_7015,N_6022);
and U8509 (N_8509,N_5124,N_6675);
or U8510 (N_8510,N_5473,N_6716);
nor U8511 (N_8511,N_6159,N_5610);
nand U8512 (N_8512,N_6846,N_5628);
and U8513 (N_8513,N_6236,N_6842);
or U8514 (N_8514,N_6787,N_5134);
or U8515 (N_8515,N_6106,N_5747);
xor U8516 (N_8516,N_6622,N_5880);
xnor U8517 (N_8517,N_7108,N_7057);
and U8518 (N_8518,N_6843,N_7091);
or U8519 (N_8519,N_7144,N_5554);
nor U8520 (N_8520,N_5193,N_7124);
and U8521 (N_8521,N_6082,N_5168);
nor U8522 (N_8522,N_6214,N_5771);
xor U8523 (N_8523,N_5236,N_5812);
xnor U8524 (N_8524,N_5396,N_7193);
xnor U8525 (N_8525,N_7464,N_7222);
and U8526 (N_8526,N_5461,N_5513);
and U8527 (N_8527,N_6008,N_6642);
or U8528 (N_8528,N_6180,N_6370);
nand U8529 (N_8529,N_7182,N_7016);
nand U8530 (N_8530,N_6527,N_6428);
xnor U8531 (N_8531,N_6356,N_5355);
and U8532 (N_8532,N_6033,N_7211);
or U8533 (N_8533,N_5359,N_7134);
or U8534 (N_8534,N_7412,N_7076);
xnor U8535 (N_8535,N_6863,N_5482);
or U8536 (N_8536,N_6943,N_6957);
or U8537 (N_8537,N_5605,N_6762);
or U8538 (N_8538,N_5092,N_6420);
xnor U8539 (N_8539,N_6274,N_7116);
xor U8540 (N_8540,N_5795,N_7382);
or U8541 (N_8541,N_5233,N_5339);
or U8542 (N_8542,N_7034,N_7114);
xor U8543 (N_8543,N_6521,N_5496);
nor U8544 (N_8544,N_7496,N_6265);
nor U8545 (N_8545,N_5595,N_6489);
and U8546 (N_8546,N_7365,N_5829);
or U8547 (N_8547,N_7163,N_6803);
nor U8548 (N_8548,N_6003,N_6930);
xor U8549 (N_8549,N_6401,N_6722);
nor U8550 (N_8550,N_5842,N_5366);
xor U8551 (N_8551,N_6002,N_5709);
and U8552 (N_8552,N_5142,N_7255);
or U8553 (N_8553,N_5888,N_7262);
xnor U8554 (N_8554,N_6368,N_5451);
and U8555 (N_8555,N_7135,N_6674);
nor U8556 (N_8556,N_6938,N_5553);
and U8557 (N_8557,N_5131,N_6138);
nor U8558 (N_8558,N_6890,N_6292);
nand U8559 (N_8559,N_6175,N_7039);
xor U8560 (N_8560,N_5409,N_7260);
or U8561 (N_8561,N_7019,N_5755);
nor U8562 (N_8562,N_7046,N_6851);
xnor U8563 (N_8563,N_6503,N_6792);
or U8564 (N_8564,N_5676,N_5164);
nor U8565 (N_8565,N_5411,N_6900);
xnor U8566 (N_8566,N_6982,N_5519);
nor U8567 (N_8567,N_5043,N_6507);
xnor U8568 (N_8568,N_5406,N_5814);
nand U8569 (N_8569,N_7371,N_7246);
and U8570 (N_8570,N_5076,N_5311);
nand U8571 (N_8571,N_6839,N_6566);
nor U8572 (N_8572,N_5041,N_5266);
nand U8573 (N_8573,N_7445,N_6692);
and U8574 (N_8574,N_7203,N_6371);
or U8575 (N_8575,N_6990,N_7080);
nand U8576 (N_8576,N_7293,N_7298);
xnor U8577 (N_8577,N_6219,N_6513);
or U8578 (N_8578,N_6142,N_7146);
xnor U8579 (N_8579,N_6181,N_5156);
and U8580 (N_8580,N_5660,N_7021);
nand U8581 (N_8581,N_7224,N_7467);
or U8582 (N_8582,N_6913,N_5469);
xor U8583 (N_8583,N_6296,N_5731);
xnor U8584 (N_8584,N_6929,N_6970);
nor U8585 (N_8585,N_6114,N_6547);
nand U8586 (N_8586,N_7439,N_6873);
nor U8587 (N_8587,N_7012,N_6079);
xnor U8588 (N_8588,N_5572,N_5064);
or U8589 (N_8589,N_6252,N_5726);
xor U8590 (N_8590,N_7006,N_5163);
or U8591 (N_8591,N_5054,N_6337);
nand U8592 (N_8592,N_5962,N_7017);
nor U8593 (N_8593,N_7297,N_6255);
nand U8594 (N_8594,N_5538,N_6594);
or U8595 (N_8595,N_6309,N_5540);
nand U8596 (N_8596,N_5107,N_7007);
nor U8597 (N_8597,N_5421,N_7156);
or U8598 (N_8598,N_5786,N_5058);
or U8599 (N_8599,N_5510,N_6999);
or U8600 (N_8600,N_7170,N_7096);
nor U8601 (N_8601,N_5426,N_6122);
nor U8602 (N_8602,N_5639,N_5069);
and U8603 (N_8603,N_6690,N_5239);
nand U8604 (N_8604,N_5285,N_6764);
xor U8605 (N_8605,N_5972,N_6608);
nor U8606 (N_8606,N_5300,N_5340);
or U8607 (N_8607,N_5507,N_5128);
xnor U8608 (N_8608,N_6988,N_5995);
nand U8609 (N_8609,N_6800,N_5535);
nor U8610 (N_8610,N_6616,N_5324);
or U8611 (N_8611,N_5706,N_7434);
xor U8612 (N_8612,N_5026,N_6605);
xnor U8613 (N_8613,N_6375,N_6808);
nand U8614 (N_8614,N_6318,N_5563);
nand U8615 (N_8615,N_6763,N_5203);
nor U8616 (N_8616,N_6314,N_6310);
xnor U8617 (N_8617,N_6155,N_6173);
xor U8618 (N_8618,N_7047,N_6714);
xor U8619 (N_8619,N_5094,N_5703);
xnor U8620 (N_8620,N_5460,N_7470);
nor U8621 (N_8621,N_6329,N_7440);
or U8622 (N_8622,N_6805,N_5059);
or U8623 (N_8623,N_5250,N_6951);
or U8624 (N_8624,N_7362,N_5827);
nand U8625 (N_8625,N_5491,N_5334);
nand U8626 (N_8626,N_7241,N_7119);
nand U8627 (N_8627,N_6302,N_7400);
or U8628 (N_8628,N_6769,N_5547);
and U8629 (N_8629,N_6884,N_6262);
or U8630 (N_8630,N_6865,N_5745);
xnor U8631 (N_8631,N_6423,N_5397);
or U8632 (N_8632,N_5875,N_7251);
nand U8633 (N_8633,N_5816,N_5607);
and U8634 (N_8634,N_6110,N_6185);
or U8635 (N_8635,N_7314,N_7195);
and U8636 (N_8636,N_6726,N_6664);
and U8637 (N_8637,N_5278,N_7361);
nor U8638 (N_8638,N_6228,N_6562);
and U8639 (N_8639,N_7028,N_5462);
and U8640 (N_8640,N_5949,N_6954);
nor U8641 (N_8641,N_6543,N_5215);
and U8642 (N_8642,N_7452,N_6099);
or U8643 (N_8643,N_6519,N_6782);
nor U8644 (N_8644,N_6928,N_6025);
xnor U8645 (N_8645,N_7254,N_6742);
xor U8646 (N_8646,N_6619,N_5764);
nand U8647 (N_8647,N_6559,N_6912);
xnor U8648 (N_8648,N_7153,N_6788);
and U8649 (N_8649,N_7479,N_5558);
nor U8650 (N_8650,N_6380,N_7072);
nand U8651 (N_8651,N_5686,N_6706);
and U8652 (N_8652,N_7037,N_6771);
nor U8653 (N_8653,N_5988,N_5864);
xor U8654 (N_8654,N_6659,N_7275);
nand U8655 (N_8655,N_6953,N_6450);
xor U8656 (N_8656,N_7164,N_6189);
nor U8657 (N_8657,N_5578,N_7497);
or U8658 (N_8658,N_7376,N_5803);
or U8659 (N_8659,N_7085,N_5895);
or U8660 (N_8660,N_5270,N_6780);
and U8661 (N_8661,N_6398,N_5276);
nor U8662 (N_8662,N_7288,N_5102);
xor U8663 (N_8663,N_7216,N_6350);
or U8664 (N_8664,N_6893,N_6940);
nand U8665 (N_8665,N_6271,N_5265);
and U8666 (N_8666,N_7427,N_5729);
nand U8667 (N_8667,N_6599,N_6636);
xor U8668 (N_8668,N_6807,N_5099);
or U8669 (N_8669,N_6991,N_7138);
nor U8670 (N_8670,N_6759,N_5937);
and U8671 (N_8671,N_5615,N_6558);
xor U8672 (N_8672,N_7306,N_7219);
nor U8673 (N_8673,N_5113,N_6412);
xor U8674 (N_8674,N_6868,N_6825);
or U8675 (N_8675,N_6076,N_5103);
nand U8676 (N_8676,N_7411,N_5950);
or U8677 (N_8677,N_7184,N_7279);
xor U8678 (N_8678,N_5229,N_7335);
nor U8679 (N_8679,N_6790,N_5243);
nand U8680 (N_8680,N_5918,N_6625);
nor U8681 (N_8681,N_6324,N_7141);
and U8682 (N_8682,N_5464,N_5818);
nand U8683 (N_8683,N_5053,N_6323);
nor U8684 (N_8684,N_7441,N_5423);
nor U8685 (N_8685,N_6395,N_5325);
and U8686 (N_8686,N_6975,N_6638);
and U8687 (N_8687,N_6015,N_6783);
xor U8688 (N_8688,N_6932,N_5647);
or U8689 (N_8689,N_6045,N_7290);
nor U8690 (N_8690,N_6774,N_6410);
or U8691 (N_8691,N_6933,N_7393);
and U8692 (N_8692,N_7460,N_6802);
or U8693 (N_8693,N_7405,N_6321);
nor U8694 (N_8694,N_6921,N_5909);
and U8695 (N_8695,N_7355,N_6518);
nor U8696 (N_8696,N_6837,N_7454);
nand U8697 (N_8697,N_5176,N_5673);
nand U8698 (N_8698,N_7111,N_6596);
nand U8699 (N_8699,N_5205,N_7429);
and U8700 (N_8700,N_7419,N_5070);
nand U8701 (N_8701,N_5231,N_5310);
xnor U8702 (N_8702,N_6515,N_6127);
or U8703 (N_8703,N_6445,N_5401);
or U8704 (N_8704,N_5618,N_5654);
nor U8705 (N_8705,N_6416,N_5149);
nor U8706 (N_8706,N_6899,N_5129);
xor U8707 (N_8707,N_7171,N_5775);
nor U8708 (N_8708,N_7206,N_5609);
xor U8709 (N_8709,N_5356,N_5784);
nand U8710 (N_8710,N_5869,N_6119);
xnor U8711 (N_8711,N_5529,N_5809);
xnor U8712 (N_8712,N_5416,N_7225);
xor U8713 (N_8713,N_6859,N_5494);
nor U8714 (N_8714,N_5095,N_7485);
nor U8715 (N_8715,N_6737,N_6026);
and U8716 (N_8716,N_6649,N_5844);
nor U8717 (N_8717,N_7196,N_5833);
nor U8718 (N_8718,N_7492,N_6411);
nor U8719 (N_8719,N_6517,N_7036);
nand U8720 (N_8720,N_6190,N_6105);
or U8721 (N_8721,N_7332,N_5016);
nor U8722 (N_8722,N_7484,N_5343);
or U8723 (N_8723,N_7183,N_5302);
nor U8724 (N_8724,N_7264,N_6902);
nor U8725 (N_8725,N_5353,N_5612);
xor U8726 (N_8726,N_6678,N_6284);
and U8727 (N_8727,N_5222,N_5608);
nor U8728 (N_8728,N_5629,N_5225);
or U8729 (N_8729,N_6878,N_6096);
or U8730 (N_8730,N_5109,N_5584);
and U8731 (N_8731,N_5414,N_6895);
nand U8732 (N_8732,N_5303,N_6903);
and U8733 (N_8733,N_6036,N_6326);
nand U8734 (N_8734,N_6986,N_7294);
or U8735 (N_8735,N_7121,N_5049);
nor U8736 (N_8736,N_5759,N_6367);
and U8737 (N_8737,N_6546,N_5980);
nand U8738 (N_8738,N_6779,N_5322);
or U8739 (N_8739,N_6404,N_6516);
and U8740 (N_8740,N_7152,N_5271);
nand U8741 (N_8741,N_5348,N_5526);
xor U8742 (N_8742,N_7311,N_7281);
xnor U8743 (N_8743,N_5226,N_5868);
nand U8744 (N_8744,N_6229,N_6120);
nor U8745 (N_8745,N_6734,N_5952);
nor U8746 (N_8746,N_7274,N_6919);
xor U8747 (N_8747,N_7399,N_5796);
nand U8748 (N_8748,N_6601,N_7155);
nand U8749 (N_8749,N_5244,N_6952);
or U8750 (N_8750,N_5932,N_6689);
nand U8751 (N_8751,N_6563,N_6540);
or U8752 (N_8752,N_7061,N_7303);
nor U8753 (N_8753,N_7080,N_5239);
xor U8754 (N_8754,N_6556,N_7193);
or U8755 (N_8755,N_7272,N_6091);
nor U8756 (N_8756,N_6983,N_6860);
nand U8757 (N_8757,N_6975,N_5374);
xor U8758 (N_8758,N_6706,N_5757);
xnor U8759 (N_8759,N_5601,N_5362);
or U8760 (N_8760,N_6972,N_5560);
or U8761 (N_8761,N_5099,N_5830);
and U8762 (N_8762,N_6859,N_6749);
nand U8763 (N_8763,N_6450,N_7162);
nor U8764 (N_8764,N_5506,N_5337);
and U8765 (N_8765,N_6495,N_5010);
and U8766 (N_8766,N_6563,N_7267);
nand U8767 (N_8767,N_5522,N_5816);
nor U8768 (N_8768,N_7253,N_5780);
nor U8769 (N_8769,N_5716,N_5679);
nor U8770 (N_8770,N_7010,N_5225);
and U8771 (N_8771,N_6739,N_6237);
and U8772 (N_8772,N_7316,N_5942);
xnor U8773 (N_8773,N_5580,N_6806);
nand U8774 (N_8774,N_5817,N_7432);
and U8775 (N_8775,N_5724,N_5182);
nor U8776 (N_8776,N_5819,N_6889);
xor U8777 (N_8777,N_7236,N_5991);
or U8778 (N_8778,N_5356,N_6310);
and U8779 (N_8779,N_5497,N_7145);
and U8780 (N_8780,N_5736,N_6081);
nor U8781 (N_8781,N_6820,N_7082);
or U8782 (N_8782,N_5265,N_6178);
xor U8783 (N_8783,N_6032,N_5166);
nand U8784 (N_8784,N_6780,N_6728);
or U8785 (N_8785,N_5159,N_5986);
and U8786 (N_8786,N_5907,N_5383);
nor U8787 (N_8787,N_6733,N_6536);
and U8788 (N_8788,N_6347,N_5605);
and U8789 (N_8789,N_5862,N_5073);
and U8790 (N_8790,N_6569,N_5973);
nand U8791 (N_8791,N_7382,N_7022);
xnor U8792 (N_8792,N_6979,N_5874);
and U8793 (N_8793,N_5037,N_5032);
or U8794 (N_8794,N_5518,N_5211);
nor U8795 (N_8795,N_5136,N_6238);
nor U8796 (N_8796,N_5336,N_5117);
and U8797 (N_8797,N_6322,N_7384);
nor U8798 (N_8798,N_5102,N_6052);
and U8799 (N_8799,N_5241,N_5467);
nand U8800 (N_8800,N_5930,N_6046);
or U8801 (N_8801,N_7344,N_7129);
nor U8802 (N_8802,N_5864,N_7327);
and U8803 (N_8803,N_6398,N_7063);
xor U8804 (N_8804,N_7333,N_5340);
nand U8805 (N_8805,N_6333,N_7255);
nand U8806 (N_8806,N_7041,N_5405);
nor U8807 (N_8807,N_5405,N_6595);
nor U8808 (N_8808,N_7116,N_6874);
nor U8809 (N_8809,N_6122,N_5798);
xor U8810 (N_8810,N_6465,N_7409);
xnor U8811 (N_8811,N_7262,N_6296);
nand U8812 (N_8812,N_5280,N_6006);
or U8813 (N_8813,N_5421,N_5993);
or U8814 (N_8814,N_5587,N_5124);
nor U8815 (N_8815,N_5207,N_6937);
nand U8816 (N_8816,N_5475,N_5157);
or U8817 (N_8817,N_5597,N_5743);
or U8818 (N_8818,N_7121,N_5147);
nor U8819 (N_8819,N_6647,N_5926);
nor U8820 (N_8820,N_5089,N_6145);
or U8821 (N_8821,N_5454,N_6527);
or U8822 (N_8822,N_5109,N_5230);
or U8823 (N_8823,N_6137,N_6049);
nor U8824 (N_8824,N_7003,N_6792);
nand U8825 (N_8825,N_6723,N_5654);
or U8826 (N_8826,N_6275,N_5081);
xor U8827 (N_8827,N_5122,N_5585);
or U8828 (N_8828,N_5598,N_5641);
and U8829 (N_8829,N_6321,N_7175);
or U8830 (N_8830,N_6683,N_5210);
or U8831 (N_8831,N_5920,N_7328);
xor U8832 (N_8832,N_5391,N_6391);
nor U8833 (N_8833,N_5446,N_6688);
and U8834 (N_8834,N_6735,N_5740);
nand U8835 (N_8835,N_7268,N_5515);
xor U8836 (N_8836,N_6869,N_5706);
xnor U8837 (N_8837,N_5290,N_5610);
or U8838 (N_8838,N_7240,N_5840);
and U8839 (N_8839,N_6505,N_6889);
and U8840 (N_8840,N_6944,N_6508);
nor U8841 (N_8841,N_6449,N_7226);
nor U8842 (N_8842,N_7120,N_7249);
and U8843 (N_8843,N_7494,N_6580);
nand U8844 (N_8844,N_7421,N_5838);
nor U8845 (N_8845,N_6931,N_6522);
and U8846 (N_8846,N_6616,N_5909);
and U8847 (N_8847,N_5530,N_7391);
nor U8848 (N_8848,N_5044,N_6406);
nor U8849 (N_8849,N_7412,N_5907);
nand U8850 (N_8850,N_5270,N_6108);
or U8851 (N_8851,N_6691,N_5647);
xor U8852 (N_8852,N_5824,N_7109);
and U8853 (N_8853,N_6998,N_6200);
nand U8854 (N_8854,N_7248,N_7138);
nand U8855 (N_8855,N_6555,N_7482);
and U8856 (N_8856,N_7086,N_7300);
nand U8857 (N_8857,N_6573,N_7317);
nor U8858 (N_8858,N_6816,N_6096);
and U8859 (N_8859,N_6999,N_5843);
nor U8860 (N_8860,N_5074,N_5369);
or U8861 (N_8861,N_6134,N_5697);
xnor U8862 (N_8862,N_6159,N_5550);
or U8863 (N_8863,N_5917,N_5425);
xnor U8864 (N_8864,N_6284,N_5351);
xnor U8865 (N_8865,N_7350,N_7074);
nand U8866 (N_8866,N_6864,N_6609);
xor U8867 (N_8867,N_6589,N_7067);
nor U8868 (N_8868,N_5742,N_5920);
xor U8869 (N_8869,N_5257,N_6091);
nor U8870 (N_8870,N_7178,N_6387);
or U8871 (N_8871,N_5844,N_6472);
nor U8872 (N_8872,N_7432,N_5954);
xor U8873 (N_8873,N_6937,N_6019);
or U8874 (N_8874,N_6389,N_6059);
nor U8875 (N_8875,N_5952,N_7311);
nand U8876 (N_8876,N_7037,N_5187);
and U8877 (N_8877,N_5797,N_6962);
xnor U8878 (N_8878,N_7023,N_5965);
or U8879 (N_8879,N_6510,N_6003);
nand U8880 (N_8880,N_5645,N_6090);
nor U8881 (N_8881,N_6849,N_5150);
xor U8882 (N_8882,N_6610,N_5515);
nor U8883 (N_8883,N_7026,N_5684);
xor U8884 (N_8884,N_6224,N_5144);
nand U8885 (N_8885,N_6023,N_6458);
and U8886 (N_8886,N_7345,N_7113);
nand U8887 (N_8887,N_5747,N_6652);
nor U8888 (N_8888,N_6443,N_7207);
xnor U8889 (N_8889,N_7216,N_7045);
nor U8890 (N_8890,N_7008,N_7487);
nand U8891 (N_8891,N_5915,N_6391);
nand U8892 (N_8892,N_6387,N_5139);
xor U8893 (N_8893,N_7147,N_5072);
nor U8894 (N_8894,N_7243,N_5012);
nor U8895 (N_8895,N_5959,N_5636);
nor U8896 (N_8896,N_5075,N_6930);
xor U8897 (N_8897,N_5739,N_5927);
xnor U8898 (N_8898,N_6495,N_5412);
and U8899 (N_8899,N_6037,N_7328);
and U8900 (N_8900,N_5355,N_6017);
xnor U8901 (N_8901,N_5572,N_5353);
and U8902 (N_8902,N_7010,N_5563);
or U8903 (N_8903,N_7099,N_7206);
nor U8904 (N_8904,N_7125,N_5661);
xnor U8905 (N_8905,N_5398,N_7034);
or U8906 (N_8906,N_5113,N_6614);
xnor U8907 (N_8907,N_5613,N_6178);
and U8908 (N_8908,N_6918,N_6767);
or U8909 (N_8909,N_6945,N_6948);
nand U8910 (N_8910,N_6029,N_5417);
nand U8911 (N_8911,N_6720,N_6682);
and U8912 (N_8912,N_7049,N_5590);
nor U8913 (N_8913,N_5056,N_5499);
nand U8914 (N_8914,N_7465,N_6181);
nor U8915 (N_8915,N_6899,N_5763);
nor U8916 (N_8916,N_6100,N_5501);
nand U8917 (N_8917,N_6320,N_5037);
nor U8918 (N_8918,N_5301,N_7128);
nand U8919 (N_8919,N_6707,N_5622);
xor U8920 (N_8920,N_6339,N_7252);
and U8921 (N_8921,N_5905,N_6503);
nand U8922 (N_8922,N_6782,N_5211);
xor U8923 (N_8923,N_7459,N_6042);
xnor U8924 (N_8924,N_6442,N_5194);
and U8925 (N_8925,N_7054,N_5694);
xnor U8926 (N_8926,N_7250,N_5031);
nor U8927 (N_8927,N_6988,N_5796);
or U8928 (N_8928,N_6006,N_5126);
nand U8929 (N_8929,N_5968,N_6750);
xor U8930 (N_8930,N_6774,N_7356);
and U8931 (N_8931,N_7292,N_6167);
or U8932 (N_8932,N_7066,N_6569);
nand U8933 (N_8933,N_7217,N_6450);
nor U8934 (N_8934,N_5488,N_5908);
nor U8935 (N_8935,N_6281,N_5790);
and U8936 (N_8936,N_7274,N_5544);
nor U8937 (N_8937,N_5784,N_5414);
xor U8938 (N_8938,N_7116,N_6179);
xnor U8939 (N_8939,N_6724,N_7487);
nand U8940 (N_8940,N_5113,N_5186);
and U8941 (N_8941,N_5343,N_7375);
or U8942 (N_8942,N_5868,N_5914);
nor U8943 (N_8943,N_5049,N_6019);
nor U8944 (N_8944,N_7345,N_5750);
or U8945 (N_8945,N_5589,N_6953);
and U8946 (N_8946,N_5081,N_6407);
nand U8947 (N_8947,N_6327,N_7462);
xnor U8948 (N_8948,N_5894,N_7408);
nand U8949 (N_8949,N_6394,N_5852);
nor U8950 (N_8950,N_5322,N_5251);
nand U8951 (N_8951,N_7449,N_5593);
nand U8952 (N_8952,N_6289,N_7288);
xnor U8953 (N_8953,N_6982,N_6901);
nor U8954 (N_8954,N_5809,N_6458);
xor U8955 (N_8955,N_5926,N_6005);
or U8956 (N_8956,N_5227,N_5085);
or U8957 (N_8957,N_5328,N_5846);
nand U8958 (N_8958,N_7079,N_7499);
xor U8959 (N_8959,N_5687,N_5777);
xor U8960 (N_8960,N_5136,N_6014);
xor U8961 (N_8961,N_7024,N_6628);
xor U8962 (N_8962,N_5049,N_5399);
and U8963 (N_8963,N_6493,N_5108);
or U8964 (N_8964,N_5123,N_7121);
or U8965 (N_8965,N_6535,N_5586);
and U8966 (N_8966,N_5554,N_7256);
nand U8967 (N_8967,N_5575,N_5119);
nand U8968 (N_8968,N_6096,N_6123);
nand U8969 (N_8969,N_6378,N_5703);
or U8970 (N_8970,N_5937,N_5701);
nand U8971 (N_8971,N_5394,N_5212);
nand U8972 (N_8972,N_6664,N_6013);
and U8973 (N_8973,N_5121,N_7287);
nor U8974 (N_8974,N_5051,N_7243);
or U8975 (N_8975,N_7405,N_5298);
and U8976 (N_8976,N_7139,N_5967);
or U8977 (N_8977,N_7370,N_6660);
or U8978 (N_8978,N_5875,N_6777);
xnor U8979 (N_8979,N_5645,N_7189);
and U8980 (N_8980,N_7267,N_5490);
and U8981 (N_8981,N_6807,N_5180);
or U8982 (N_8982,N_5661,N_5142);
or U8983 (N_8983,N_5023,N_5876);
nor U8984 (N_8984,N_5339,N_7264);
nor U8985 (N_8985,N_5257,N_5786);
and U8986 (N_8986,N_5462,N_5421);
nand U8987 (N_8987,N_6609,N_5641);
nor U8988 (N_8988,N_7399,N_7282);
and U8989 (N_8989,N_5587,N_6493);
nor U8990 (N_8990,N_6179,N_5796);
nand U8991 (N_8991,N_7123,N_7404);
and U8992 (N_8992,N_6120,N_6967);
and U8993 (N_8993,N_5495,N_6470);
xnor U8994 (N_8994,N_5854,N_7388);
nand U8995 (N_8995,N_6986,N_7040);
nand U8996 (N_8996,N_6517,N_5750);
xnor U8997 (N_8997,N_5494,N_5918);
nor U8998 (N_8998,N_5543,N_6065);
nand U8999 (N_8999,N_5819,N_6250);
or U9000 (N_9000,N_5153,N_6035);
and U9001 (N_9001,N_5854,N_5817);
xnor U9002 (N_9002,N_6972,N_6711);
and U9003 (N_9003,N_7483,N_5986);
or U9004 (N_9004,N_5798,N_6816);
or U9005 (N_9005,N_5051,N_7169);
xnor U9006 (N_9006,N_6752,N_5631);
nand U9007 (N_9007,N_6067,N_7164);
nor U9008 (N_9008,N_5841,N_5062);
nand U9009 (N_9009,N_6031,N_6016);
xor U9010 (N_9010,N_5902,N_5647);
and U9011 (N_9011,N_5281,N_5463);
and U9012 (N_9012,N_6130,N_6132);
xnor U9013 (N_9013,N_5157,N_6363);
and U9014 (N_9014,N_7151,N_5570);
xnor U9015 (N_9015,N_5249,N_7417);
nand U9016 (N_9016,N_6321,N_7494);
and U9017 (N_9017,N_5029,N_7016);
or U9018 (N_9018,N_5994,N_6881);
nor U9019 (N_9019,N_6396,N_6924);
nor U9020 (N_9020,N_7138,N_7147);
xnor U9021 (N_9021,N_5963,N_5464);
and U9022 (N_9022,N_7193,N_6201);
nor U9023 (N_9023,N_5281,N_5887);
xor U9024 (N_9024,N_5962,N_6369);
and U9025 (N_9025,N_5507,N_5947);
and U9026 (N_9026,N_5623,N_5795);
nand U9027 (N_9027,N_6425,N_5034);
nor U9028 (N_9028,N_5183,N_5348);
and U9029 (N_9029,N_7016,N_6049);
nor U9030 (N_9030,N_5532,N_5382);
nor U9031 (N_9031,N_5593,N_6176);
nand U9032 (N_9032,N_5307,N_5565);
nor U9033 (N_9033,N_6287,N_5641);
and U9034 (N_9034,N_6061,N_6590);
or U9035 (N_9035,N_5598,N_7015);
nor U9036 (N_9036,N_6948,N_7397);
and U9037 (N_9037,N_6600,N_7341);
xnor U9038 (N_9038,N_5412,N_7240);
nand U9039 (N_9039,N_6042,N_5204);
nor U9040 (N_9040,N_7382,N_7479);
xor U9041 (N_9041,N_6206,N_6032);
nand U9042 (N_9042,N_6607,N_5949);
nand U9043 (N_9043,N_6680,N_5184);
nor U9044 (N_9044,N_6958,N_6956);
xnor U9045 (N_9045,N_6203,N_5322);
nor U9046 (N_9046,N_6492,N_5293);
nor U9047 (N_9047,N_6467,N_6400);
nor U9048 (N_9048,N_7012,N_6233);
or U9049 (N_9049,N_6680,N_7215);
nor U9050 (N_9050,N_6655,N_7396);
xor U9051 (N_9051,N_6424,N_6348);
nand U9052 (N_9052,N_7148,N_6054);
and U9053 (N_9053,N_5328,N_6516);
and U9054 (N_9054,N_6116,N_5544);
nand U9055 (N_9055,N_6930,N_5137);
nor U9056 (N_9056,N_7339,N_6220);
and U9057 (N_9057,N_5163,N_5976);
xnor U9058 (N_9058,N_7060,N_6887);
and U9059 (N_9059,N_6693,N_6183);
xnor U9060 (N_9060,N_7159,N_7223);
and U9061 (N_9061,N_7335,N_6606);
xor U9062 (N_9062,N_6236,N_6704);
nor U9063 (N_9063,N_7027,N_5239);
xnor U9064 (N_9064,N_5793,N_7036);
nor U9065 (N_9065,N_6178,N_5536);
or U9066 (N_9066,N_6500,N_7050);
or U9067 (N_9067,N_5337,N_5881);
nand U9068 (N_9068,N_5019,N_5795);
xor U9069 (N_9069,N_7035,N_5577);
and U9070 (N_9070,N_6991,N_7064);
nor U9071 (N_9071,N_7160,N_6138);
nor U9072 (N_9072,N_5167,N_5895);
and U9073 (N_9073,N_5785,N_6211);
nor U9074 (N_9074,N_5264,N_5895);
nand U9075 (N_9075,N_6129,N_5631);
nand U9076 (N_9076,N_5997,N_7335);
xor U9077 (N_9077,N_7181,N_5117);
or U9078 (N_9078,N_5175,N_6306);
nor U9079 (N_9079,N_6999,N_7426);
and U9080 (N_9080,N_7130,N_5190);
and U9081 (N_9081,N_6753,N_6079);
nand U9082 (N_9082,N_6104,N_5027);
nand U9083 (N_9083,N_5470,N_6178);
or U9084 (N_9084,N_6770,N_7172);
nand U9085 (N_9085,N_5078,N_5975);
nand U9086 (N_9086,N_6753,N_7227);
or U9087 (N_9087,N_7471,N_5644);
or U9088 (N_9088,N_6015,N_6157);
nand U9089 (N_9089,N_5521,N_5663);
xor U9090 (N_9090,N_5461,N_5174);
or U9091 (N_9091,N_6110,N_6730);
and U9092 (N_9092,N_7321,N_7335);
or U9093 (N_9093,N_5905,N_6482);
nand U9094 (N_9094,N_5328,N_6090);
or U9095 (N_9095,N_7471,N_5075);
or U9096 (N_9096,N_5147,N_6575);
nand U9097 (N_9097,N_6856,N_7332);
nor U9098 (N_9098,N_5269,N_7012);
or U9099 (N_9099,N_5291,N_7470);
nand U9100 (N_9100,N_6208,N_6636);
nand U9101 (N_9101,N_5323,N_5726);
or U9102 (N_9102,N_6344,N_5634);
or U9103 (N_9103,N_5377,N_5469);
xnor U9104 (N_9104,N_6652,N_6318);
or U9105 (N_9105,N_5288,N_7031);
and U9106 (N_9106,N_5909,N_5513);
nand U9107 (N_9107,N_5625,N_7402);
nor U9108 (N_9108,N_5940,N_5833);
nor U9109 (N_9109,N_5221,N_5223);
nor U9110 (N_9110,N_6078,N_6335);
xor U9111 (N_9111,N_6508,N_6733);
or U9112 (N_9112,N_7431,N_6091);
and U9113 (N_9113,N_6663,N_6407);
and U9114 (N_9114,N_6371,N_6038);
nand U9115 (N_9115,N_7034,N_7105);
nor U9116 (N_9116,N_6827,N_5429);
or U9117 (N_9117,N_6709,N_6621);
and U9118 (N_9118,N_6680,N_6030);
xnor U9119 (N_9119,N_5254,N_7032);
nor U9120 (N_9120,N_5001,N_6417);
nand U9121 (N_9121,N_6812,N_6378);
nor U9122 (N_9122,N_7342,N_5363);
nor U9123 (N_9123,N_7065,N_5461);
or U9124 (N_9124,N_5461,N_6394);
xnor U9125 (N_9125,N_7471,N_6748);
nor U9126 (N_9126,N_6684,N_5859);
xnor U9127 (N_9127,N_6880,N_5133);
xnor U9128 (N_9128,N_5780,N_5545);
xor U9129 (N_9129,N_5181,N_6870);
nand U9130 (N_9130,N_6288,N_7408);
and U9131 (N_9131,N_5729,N_5841);
xnor U9132 (N_9132,N_5535,N_5364);
or U9133 (N_9133,N_6653,N_5531);
or U9134 (N_9134,N_6757,N_5237);
or U9135 (N_9135,N_5276,N_7067);
nor U9136 (N_9136,N_6360,N_5838);
and U9137 (N_9137,N_6182,N_5162);
nand U9138 (N_9138,N_6268,N_5651);
nor U9139 (N_9139,N_6616,N_6784);
xor U9140 (N_9140,N_7455,N_5530);
nand U9141 (N_9141,N_7418,N_6360);
nand U9142 (N_9142,N_6518,N_5253);
nor U9143 (N_9143,N_5734,N_6939);
or U9144 (N_9144,N_5473,N_5515);
and U9145 (N_9145,N_6466,N_6297);
and U9146 (N_9146,N_5966,N_5971);
or U9147 (N_9147,N_6308,N_5223);
nand U9148 (N_9148,N_5530,N_6444);
nor U9149 (N_9149,N_7318,N_6481);
nand U9150 (N_9150,N_6467,N_6915);
nand U9151 (N_9151,N_7288,N_6006);
or U9152 (N_9152,N_6329,N_7326);
xor U9153 (N_9153,N_6606,N_6980);
xor U9154 (N_9154,N_6738,N_7257);
or U9155 (N_9155,N_5760,N_6072);
nand U9156 (N_9156,N_6113,N_7462);
or U9157 (N_9157,N_6245,N_6320);
nor U9158 (N_9158,N_7299,N_7306);
nor U9159 (N_9159,N_5501,N_6767);
and U9160 (N_9160,N_5173,N_6506);
or U9161 (N_9161,N_6546,N_6373);
xnor U9162 (N_9162,N_6927,N_6926);
or U9163 (N_9163,N_6424,N_7165);
xor U9164 (N_9164,N_6437,N_7387);
or U9165 (N_9165,N_6836,N_5199);
and U9166 (N_9166,N_6427,N_6839);
or U9167 (N_9167,N_5865,N_6284);
or U9168 (N_9168,N_6095,N_7151);
nand U9169 (N_9169,N_6784,N_6259);
or U9170 (N_9170,N_6122,N_5930);
xnor U9171 (N_9171,N_7458,N_7109);
nand U9172 (N_9172,N_5221,N_6146);
xor U9173 (N_9173,N_6136,N_6533);
xor U9174 (N_9174,N_5655,N_7451);
nand U9175 (N_9175,N_7237,N_5542);
xnor U9176 (N_9176,N_6497,N_6478);
nand U9177 (N_9177,N_5941,N_7289);
xnor U9178 (N_9178,N_6570,N_6283);
nand U9179 (N_9179,N_7456,N_5284);
xnor U9180 (N_9180,N_7338,N_6094);
and U9181 (N_9181,N_6076,N_6211);
and U9182 (N_9182,N_7324,N_7471);
and U9183 (N_9183,N_5509,N_7087);
and U9184 (N_9184,N_7023,N_5073);
and U9185 (N_9185,N_5588,N_7404);
xor U9186 (N_9186,N_5590,N_6898);
and U9187 (N_9187,N_5062,N_6900);
and U9188 (N_9188,N_6549,N_5204);
or U9189 (N_9189,N_5419,N_6852);
nand U9190 (N_9190,N_6734,N_7384);
nand U9191 (N_9191,N_7109,N_6357);
xor U9192 (N_9192,N_6476,N_5731);
nand U9193 (N_9193,N_5293,N_6280);
nand U9194 (N_9194,N_6235,N_7030);
and U9195 (N_9195,N_6302,N_6203);
nor U9196 (N_9196,N_6800,N_5941);
nor U9197 (N_9197,N_7003,N_5151);
or U9198 (N_9198,N_5827,N_5654);
xor U9199 (N_9199,N_5077,N_5750);
and U9200 (N_9200,N_6444,N_5067);
or U9201 (N_9201,N_6783,N_5901);
nand U9202 (N_9202,N_6499,N_5846);
nor U9203 (N_9203,N_7446,N_5238);
nand U9204 (N_9204,N_5520,N_6106);
or U9205 (N_9205,N_5325,N_6896);
nor U9206 (N_9206,N_7128,N_6074);
and U9207 (N_9207,N_5083,N_7148);
and U9208 (N_9208,N_6892,N_6425);
or U9209 (N_9209,N_7163,N_5269);
and U9210 (N_9210,N_6327,N_5205);
nand U9211 (N_9211,N_6705,N_5977);
nor U9212 (N_9212,N_5073,N_6042);
xnor U9213 (N_9213,N_6763,N_6486);
nand U9214 (N_9214,N_6235,N_7421);
or U9215 (N_9215,N_6670,N_7421);
xnor U9216 (N_9216,N_5613,N_7265);
nand U9217 (N_9217,N_5605,N_5403);
xnor U9218 (N_9218,N_5082,N_6356);
nor U9219 (N_9219,N_5504,N_6467);
nand U9220 (N_9220,N_7180,N_6303);
xnor U9221 (N_9221,N_6106,N_5473);
nand U9222 (N_9222,N_5554,N_6072);
and U9223 (N_9223,N_6690,N_7481);
or U9224 (N_9224,N_5311,N_6962);
xnor U9225 (N_9225,N_6687,N_6737);
nand U9226 (N_9226,N_5453,N_6521);
nand U9227 (N_9227,N_5451,N_7277);
nand U9228 (N_9228,N_5101,N_6479);
xor U9229 (N_9229,N_5038,N_5720);
nand U9230 (N_9230,N_7220,N_5521);
and U9231 (N_9231,N_5867,N_6793);
xor U9232 (N_9232,N_5317,N_7165);
xor U9233 (N_9233,N_6642,N_5972);
xor U9234 (N_9234,N_6777,N_5777);
xor U9235 (N_9235,N_6528,N_5870);
and U9236 (N_9236,N_5670,N_7253);
nand U9237 (N_9237,N_5469,N_5907);
xnor U9238 (N_9238,N_7178,N_5729);
nand U9239 (N_9239,N_5823,N_6627);
xor U9240 (N_9240,N_6970,N_6087);
nor U9241 (N_9241,N_7320,N_5676);
and U9242 (N_9242,N_7271,N_6980);
or U9243 (N_9243,N_5607,N_5450);
xnor U9244 (N_9244,N_6322,N_5500);
or U9245 (N_9245,N_5483,N_7241);
or U9246 (N_9246,N_6868,N_7469);
and U9247 (N_9247,N_6750,N_6320);
xor U9248 (N_9248,N_6958,N_5268);
xor U9249 (N_9249,N_5269,N_5943);
or U9250 (N_9250,N_6673,N_7282);
or U9251 (N_9251,N_5572,N_6041);
or U9252 (N_9252,N_5213,N_5835);
nand U9253 (N_9253,N_5854,N_5425);
nor U9254 (N_9254,N_7069,N_6366);
and U9255 (N_9255,N_5540,N_7081);
xnor U9256 (N_9256,N_6472,N_6032);
nor U9257 (N_9257,N_7121,N_5885);
xnor U9258 (N_9258,N_5853,N_7183);
and U9259 (N_9259,N_5590,N_7354);
xnor U9260 (N_9260,N_5482,N_5392);
nor U9261 (N_9261,N_6639,N_7191);
nand U9262 (N_9262,N_7464,N_6060);
nand U9263 (N_9263,N_5058,N_5080);
nor U9264 (N_9264,N_5019,N_5092);
xor U9265 (N_9265,N_6160,N_7036);
xnor U9266 (N_9266,N_6112,N_6811);
nor U9267 (N_9267,N_5563,N_6492);
or U9268 (N_9268,N_5433,N_5075);
xor U9269 (N_9269,N_5864,N_6390);
or U9270 (N_9270,N_6820,N_7123);
and U9271 (N_9271,N_7132,N_6404);
nand U9272 (N_9272,N_5990,N_6901);
nand U9273 (N_9273,N_7392,N_6223);
nor U9274 (N_9274,N_6028,N_5526);
nor U9275 (N_9275,N_5130,N_5512);
and U9276 (N_9276,N_6034,N_6329);
and U9277 (N_9277,N_5094,N_6199);
or U9278 (N_9278,N_5554,N_6869);
xor U9279 (N_9279,N_7354,N_6709);
and U9280 (N_9280,N_6987,N_6170);
nand U9281 (N_9281,N_6275,N_5779);
nor U9282 (N_9282,N_5057,N_6050);
or U9283 (N_9283,N_5547,N_6488);
or U9284 (N_9284,N_6778,N_5729);
and U9285 (N_9285,N_7036,N_6180);
and U9286 (N_9286,N_6696,N_6169);
and U9287 (N_9287,N_7041,N_5650);
or U9288 (N_9288,N_6753,N_7106);
and U9289 (N_9289,N_6379,N_6437);
or U9290 (N_9290,N_5354,N_5311);
nor U9291 (N_9291,N_6469,N_6249);
xnor U9292 (N_9292,N_5065,N_5112);
nand U9293 (N_9293,N_6592,N_6894);
and U9294 (N_9294,N_6657,N_7317);
nor U9295 (N_9295,N_5609,N_6564);
or U9296 (N_9296,N_6350,N_5148);
xnor U9297 (N_9297,N_5392,N_6083);
nand U9298 (N_9298,N_6457,N_5118);
nor U9299 (N_9299,N_5685,N_6224);
and U9300 (N_9300,N_6963,N_7278);
nand U9301 (N_9301,N_7084,N_5058);
xor U9302 (N_9302,N_5200,N_5549);
nor U9303 (N_9303,N_7105,N_6477);
xnor U9304 (N_9304,N_6684,N_6168);
nand U9305 (N_9305,N_5082,N_5875);
nor U9306 (N_9306,N_6918,N_5252);
xnor U9307 (N_9307,N_5030,N_6410);
xnor U9308 (N_9308,N_5178,N_7297);
nand U9309 (N_9309,N_6085,N_5630);
nor U9310 (N_9310,N_7124,N_6185);
nand U9311 (N_9311,N_6117,N_6106);
or U9312 (N_9312,N_5731,N_5708);
nor U9313 (N_9313,N_5062,N_6497);
xnor U9314 (N_9314,N_5218,N_7047);
xnor U9315 (N_9315,N_5998,N_5519);
nand U9316 (N_9316,N_6033,N_6010);
xor U9317 (N_9317,N_6872,N_5320);
nor U9318 (N_9318,N_6960,N_5212);
nand U9319 (N_9319,N_6512,N_5431);
nand U9320 (N_9320,N_5376,N_5810);
and U9321 (N_9321,N_7252,N_7475);
or U9322 (N_9322,N_5014,N_6845);
or U9323 (N_9323,N_5056,N_5513);
and U9324 (N_9324,N_5180,N_5428);
xnor U9325 (N_9325,N_6948,N_5275);
or U9326 (N_9326,N_5273,N_7176);
and U9327 (N_9327,N_5337,N_6443);
or U9328 (N_9328,N_6881,N_6115);
and U9329 (N_9329,N_7149,N_6638);
or U9330 (N_9330,N_6606,N_5262);
and U9331 (N_9331,N_6998,N_5650);
nor U9332 (N_9332,N_6466,N_6149);
or U9333 (N_9333,N_5994,N_7417);
nand U9334 (N_9334,N_6594,N_5395);
nor U9335 (N_9335,N_6643,N_6721);
nand U9336 (N_9336,N_6694,N_6788);
nand U9337 (N_9337,N_6099,N_6322);
and U9338 (N_9338,N_6720,N_6604);
nor U9339 (N_9339,N_6746,N_6568);
and U9340 (N_9340,N_5694,N_7285);
xor U9341 (N_9341,N_6235,N_5048);
nand U9342 (N_9342,N_7327,N_7419);
nand U9343 (N_9343,N_6813,N_5538);
nor U9344 (N_9344,N_5564,N_6598);
nor U9345 (N_9345,N_5568,N_6616);
or U9346 (N_9346,N_6987,N_7005);
nand U9347 (N_9347,N_5255,N_6455);
and U9348 (N_9348,N_5580,N_7108);
xor U9349 (N_9349,N_7452,N_7273);
or U9350 (N_9350,N_5574,N_6710);
and U9351 (N_9351,N_6167,N_5201);
xnor U9352 (N_9352,N_6532,N_6843);
xnor U9353 (N_9353,N_6515,N_5521);
nor U9354 (N_9354,N_5445,N_7446);
nor U9355 (N_9355,N_5794,N_6685);
and U9356 (N_9356,N_6303,N_5944);
xor U9357 (N_9357,N_6752,N_6467);
nor U9358 (N_9358,N_5477,N_7491);
nand U9359 (N_9359,N_5748,N_5746);
or U9360 (N_9360,N_5543,N_5242);
and U9361 (N_9361,N_6253,N_6469);
xor U9362 (N_9362,N_5965,N_6144);
nand U9363 (N_9363,N_6652,N_5017);
or U9364 (N_9364,N_6228,N_5270);
or U9365 (N_9365,N_5139,N_5526);
or U9366 (N_9366,N_6042,N_5640);
nand U9367 (N_9367,N_7381,N_6060);
or U9368 (N_9368,N_6860,N_5298);
nand U9369 (N_9369,N_5263,N_7148);
xor U9370 (N_9370,N_7463,N_5157);
xnor U9371 (N_9371,N_7445,N_5091);
xor U9372 (N_9372,N_5079,N_5428);
nand U9373 (N_9373,N_6992,N_6401);
and U9374 (N_9374,N_5719,N_5929);
nor U9375 (N_9375,N_5676,N_5377);
xor U9376 (N_9376,N_6515,N_5726);
and U9377 (N_9377,N_7231,N_7331);
and U9378 (N_9378,N_6885,N_6355);
nand U9379 (N_9379,N_7211,N_7206);
nor U9380 (N_9380,N_5958,N_6692);
nand U9381 (N_9381,N_6249,N_7399);
or U9382 (N_9382,N_5239,N_6911);
xnor U9383 (N_9383,N_5351,N_5902);
and U9384 (N_9384,N_7460,N_7127);
and U9385 (N_9385,N_6854,N_5507);
xnor U9386 (N_9386,N_5851,N_5904);
and U9387 (N_9387,N_7168,N_5764);
nand U9388 (N_9388,N_5457,N_7466);
xnor U9389 (N_9389,N_6211,N_7339);
nor U9390 (N_9390,N_5622,N_6581);
xnor U9391 (N_9391,N_6634,N_5587);
nor U9392 (N_9392,N_5461,N_5175);
and U9393 (N_9393,N_5173,N_6097);
and U9394 (N_9394,N_5363,N_6527);
xnor U9395 (N_9395,N_6082,N_6447);
and U9396 (N_9396,N_6524,N_6266);
and U9397 (N_9397,N_6362,N_5773);
and U9398 (N_9398,N_6623,N_6120);
nand U9399 (N_9399,N_7172,N_7082);
xor U9400 (N_9400,N_7254,N_5227);
and U9401 (N_9401,N_5964,N_5645);
or U9402 (N_9402,N_6779,N_6754);
and U9403 (N_9403,N_5849,N_6049);
and U9404 (N_9404,N_5665,N_5569);
and U9405 (N_9405,N_5768,N_6118);
or U9406 (N_9406,N_5048,N_7225);
xnor U9407 (N_9407,N_5462,N_7014);
nor U9408 (N_9408,N_7349,N_5099);
or U9409 (N_9409,N_6170,N_6000);
nor U9410 (N_9410,N_5207,N_6454);
nor U9411 (N_9411,N_7216,N_6001);
and U9412 (N_9412,N_5236,N_5655);
nor U9413 (N_9413,N_5650,N_5839);
xor U9414 (N_9414,N_5962,N_6830);
nor U9415 (N_9415,N_5169,N_5460);
and U9416 (N_9416,N_5408,N_5174);
nor U9417 (N_9417,N_6192,N_5376);
or U9418 (N_9418,N_7013,N_6607);
xnor U9419 (N_9419,N_5917,N_7046);
nand U9420 (N_9420,N_6449,N_6930);
or U9421 (N_9421,N_6139,N_6720);
nand U9422 (N_9422,N_7129,N_6436);
nor U9423 (N_9423,N_6236,N_7201);
nand U9424 (N_9424,N_6599,N_7311);
or U9425 (N_9425,N_7464,N_7103);
nor U9426 (N_9426,N_5946,N_6852);
xnor U9427 (N_9427,N_7151,N_6474);
or U9428 (N_9428,N_6538,N_5024);
or U9429 (N_9429,N_6364,N_5969);
or U9430 (N_9430,N_5717,N_5599);
nor U9431 (N_9431,N_5804,N_5592);
nor U9432 (N_9432,N_7440,N_5785);
nand U9433 (N_9433,N_6654,N_5790);
and U9434 (N_9434,N_6345,N_6092);
or U9435 (N_9435,N_5489,N_6800);
xnor U9436 (N_9436,N_6961,N_5324);
or U9437 (N_9437,N_7460,N_6971);
nand U9438 (N_9438,N_5064,N_7001);
xor U9439 (N_9439,N_6719,N_6931);
or U9440 (N_9440,N_7328,N_6723);
and U9441 (N_9441,N_6167,N_5972);
and U9442 (N_9442,N_6181,N_7052);
nand U9443 (N_9443,N_7064,N_6728);
nor U9444 (N_9444,N_5666,N_6892);
nand U9445 (N_9445,N_6474,N_6534);
and U9446 (N_9446,N_7034,N_5829);
xor U9447 (N_9447,N_7147,N_5104);
nor U9448 (N_9448,N_6077,N_7312);
nand U9449 (N_9449,N_7072,N_6599);
xor U9450 (N_9450,N_5903,N_5822);
xnor U9451 (N_9451,N_6072,N_5149);
and U9452 (N_9452,N_7432,N_6976);
nand U9453 (N_9453,N_7487,N_6487);
or U9454 (N_9454,N_6039,N_5091);
nand U9455 (N_9455,N_7330,N_6394);
or U9456 (N_9456,N_5742,N_7469);
nand U9457 (N_9457,N_5471,N_6248);
or U9458 (N_9458,N_5736,N_6885);
xor U9459 (N_9459,N_5602,N_5484);
xnor U9460 (N_9460,N_6647,N_7029);
xor U9461 (N_9461,N_7445,N_6025);
xor U9462 (N_9462,N_5138,N_5114);
nor U9463 (N_9463,N_7034,N_5119);
nand U9464 (N_9464,N_6632,N_5498);
nand U9465 (N_9465,N_7296,N_5001);
nand U9466 (N_9466,N_5203,N_6780);
or U9467 (N_9467,N_6834,N_6554);
and U9468 (N_9468,N_7419,N_5964);
nand U9469 (N_9469,N_5457,N_5356);
nor U9470 (N_9470,N_5440,N_5974);
nor U9471 (N_9471,N_6126,N_5379);
nor U9472 (N_9472,N_7453,N_6286);
nor U9473 (N_9473,N_6710,N_5367);
nor U9474 (N_9474,N_6639,N_5765);
nor U9475 (N_9475,N_5093,N_6562);
nor U9476 (N_9476,N_5231,N_5940);
and U9477 (N_9477,N_5607,N_5127);
nand U9478 (N_9478,N_5883,N_5315);
nor U9479 (N_9479,N_6667,N_5625);
and U9480 (N_9480,N_6418,N_6964);
xor U9481 (N_9481,N_5900,N_7027);
nor U9482 (N_9482,N_6090,N_6395);
xor U9483 (N_9483,N_5085,N_6699);
or U9484 (N_9484,N_5001,N_5819);
or U9485 (N_9485,N_5465,N_6570);
nor U9486 (N_9486,N_5751,N_6742);
and U9487 (N_9487,N_5889,N_7116);
or U9488 (N_9488,N_6416,N_5661);
or U9489 (N_9489,N_7172,N_7068);
or U9490 (N_9490,N_6463,N_6867);
nor U9491 (N_9491,N_5524,N_5717);
or U9492 (N_9492,N_6970,N_5200);
or U9493 (N_9493,N_6702,N_5768);
xnor U9494 (N_9494,N_7423,N_5928);
and U9495 (N_9495,N_5810,N_7496);
xor U9496 (N_9496,N_6742,N_7135);
nand U9497 (N_9497,N_7177,N_7096);
nand U9498 (N_9498,N_7478,N_6268);
nand U9499 (N_9499,N_6953,N_7000);
xnor U9500 (N_9500,N_5527,N_5947);
or U9501 (N_9501,N_6762,N_7079);
nor U9502 (N_9502,N_5531,N_5727);
and U9503 (N_9503,N_6953,N_6015);
nand U9504 (N_9504,N_5554,N_5939);
xnor U9505 (N_9505,N_5025,N_5298);
xor U9506 (N_9506,N_6923,N_7276);
and U9507 (N_9507,N_5011,N_7280);
and U9508 (N_9508,N_5887,N_5809);
nand U9509 (N_9509,N_5182,N_7225);
and U9510 (N_9510,N_7454,N_7251);
or U9511 (N_9511,N_5848,N_6721);
and U9512 (N_9512,N_7487,N_5369);
nand U9513 (N_9513,N_6497,N_6193);
nand U9514 (N_9514,N_5737,N_6947);
or U9515 (N_9515,N_6946,N_6496);
nand U9516 (N_9516,N_6840,N_7254);
and U9517 (N_9517,N_6074,N_6343);
nand U9518 (N_9518,N_7358,N_6689);
nand U9519 (N_9519,N_6042,N_7261);
or U9520 (N_9520,N_5816,N_7404);
or U9521 (N_9521,N_7081,N_6492);
nand U9522 (N_9522,N_5229,N_5469);
nand U9523 (N_9523,N_5967,N_5553);
xnor U9524 (N_9524,N_5268,N_5270);
nand U9525 (N_9525,N_6379,N_6214);
nor U9526 (N_9526,N_5259,N_5735);
or U9527 (N_9527,N_5744,N_5110);
and U9528 (N_9528,N_5546,N_6365);
nand U9529 (N_9529,N_6092,N_6251);
and U9530 (N_9530,N_5151,N_6008);
xnor U9531 (N_9531,N_6935,N_6218);
nor U9532 (N_9532,N_6655,N_7409);
xnor U9533 (N_9533,N_7110,N_6801);
and U9534 (N_9534,N_6101,N_5056);
or U9535 (N_9535,N_5595,N_5025);
xor U9536 (N_9536,N_6866,N_5100);
or U9537 (N_9537,N_6842,N_6128);
xnor U9538 (N_9538,N_6886,N_7443);
or U9539 (N_9539,N_5639,N_5894);
nor U9540 (N_9540,N_6980,N_6222);
xnor U9541 (N_9541,N_5949,N_5107);
and U9542 (N_9542,N_5775,N_7458);
and U9543 (N_9543,N_5190,N_5566);
nor U9544 (N_9544,N_7470,N_5815);
nand U9545 (N_9545,N_6535,N_5726);
nor U9546 (N_9546,N_6113,N_6188);
nand U9547 (N_9547,N_5798,N_5575);
or U9548 (N_9548,N_6659,N_6716);
nor U9549 (N_9549,N_7281,N_6228);
nand U9550 (N_9550,N_5760,N_7276);
or U9551 (N_9551,N_6327,N_5118);
nor U9552 (N_9552,N_7164,N_5727);
nand U9553 (N_9553,N_6210,N_6675);
and U9554 (N_9554,N_5762,N_7478);
xor U9555 (N_9555,N_5339,N_6137);
or U9556 (N_9556,N_6490,N_7483);
or U9557 (N_9557,N_5616,N_5411);
nand U9558 (N_9558,N_7042,N_6080);
or U9559 (N_9559,N_5308,N_5246);
and U9560 (N_9560,N_6753,N_5599);
xnor U9561 (N_9561,N_6772,N_7143);
or U9562 (N_9562,N_5646,N_5227);
xor U9563 (N_9563,N_6544,N_5276);
or U9564 (N_9564,N_5585,N_6684);
xor U9565 (N_9565,N_7262,N_6843);
and U9566 (N_9566,N_7117,N_5896);
or U9567 (N_9567,N_6750,N_6306);
or U9568 (N_9568,N_6224,N_6598);
nand U9569 (N_9569,N_5222,N_5399);
or U9570 (N_9570,N_5494,N_6141);
and U9571 (N_9571,N_5123,N_6721);
xor U9572 (N_9572,N_7082,N_5446);
xnor U9573 (N_9573,N_5234,N_5683);
nand U9574 (N_9574,N_5651,N_7468);
and U9575 (N_9575,N_6197,N_5097);
nor U9576 (N_9576,N_6921,N_5783);
nor U9577 (N_9577,N_7145,N_6296);
and U9578 (N_9578,N_5450,N_6833);
or U9579 (N_9579,N_5137,N_6720);
or U9580 (N_9580,N_7133,N_7273);
nor U9581 (N_9581,N_5595,N_5336);
nor U9582 (N_9582,N_5808,N_5390);
or U9583 (N_9583,N_6288,N_5274);
nor U9584 (N_9584,N_7153,N_6568);
nand U9585 (N_9585,N_6197,N_5130);
and U9586 (N_9586,N_6723,N_6841);
and U9587 (N_9587,N_6617,N_5753);
xnor U9588 (N_9588,N_7365,N_5848);
and U9589 (N_9589,N_6116,N_7402);
and U9590 (N_9590,N_5594,N_7034);
and U9591 (N_9591,N_5203,N_5035);
and U9592 (N_9592,N_6245,N_6402);
nand U9593 (N_9593,N_5303,N_6320);
nand U9594 (N_9594,N_5347,N_5696);
nor U9595 (N_9595,N_5658,N_6822);
and U9596 (N_9596,N_7420,N_7205);
or U9597 (N_9597,N_5401,N_7481);
xor U9598 (N_9598,N_6734,N_6261);
nor U9599 (N_9599,N_5364,N_5638);
and U9600 (N_9600,N_5727,N_6569);
or U9601 (N_9601,N_5455,N_5056);
nand U9602 (N_9602,N_5455,N_6976);
nand U9603 (N_9603,N_6968,N_6600);
nor U9604 (N_9604,N_5494,N_7364);
nand U9605 (N_9605,N_5941,N_6840);
nand U9606 (N_9606,N_5853,N_6345);
xnor U9607 (N_9607,N_5363,N_6163);
nand U9608 (N_9608,N_7160,N_7013);
and U9609 (N_9609,N_5286,N_5832);
and U9610 (N_9610,N_5476,N_6501);
or U9611 (N_9611,N_5942,N_6276);
nor U9612 (N_9612,N_7064,N_7340);
xor U9613 (N_9613,N_5149,N_6638);
nand U9614 (N_9614,N_5333,N_5305);
nand U9615 (N_9615,N_5479,N_5596);
and U9616 (N_9616,N_7395,N_5995);
nor U9617 (N_9617,N_5876,N_5433);
or U9618 (N_9618,N_5943,N_5447);
and U9619 (N_9619,N_6440,N_7146);
nand U9620 (N_9620,N_6918,N_6488);
nor U9621 (N_9621,N_6766,N_6986);
nand U9622 (N_9622,N_6437,N_6238);
xor U9623 (N_9623,N_5009,N_5420);
nand U9624 (N_9624,N_6349,N_5371);
nand U9625 (N_9625,N_6662,N_6993);
xnor U9626 (N_9626,N_5910,N_7229);
xnor U9627 (N_9627,N_6875,N_6211);
nor U9628 (N_9628,N_5715,N_7262);
or U9629 (N_9629,N_5219,N_6040);
nand U9630 (N_9630,N_6292,N_5600);
xnor U9631 (N_9631,N_5588,N_6260);
and U9632 (N_9632,N_6464,N_7303);
or U9633 (N_9633,N_5010,N_5620);
nor U9634 (N_9634,N_5714,N_5555);
or U9635 (N_9635,N_7330,N_7025);
nor U9636 (N_9636,N_6287,N_6494);
nand U9637 (N_9637,N_6685,N_6119);
and U9638 (N_9638,N_6306,N_5468);
nor U9639 (N_9639,N_7386,N_6716);
xor U9640 (N_9640,N_6408,N_6756);
nor U9641 (N_9641,N_5819,N_7112);
and U9642 (N_9642,N_5155,N_6230);
or U9643 (N_9643,N_7258,N_6075);
nor U9644 (N_9644,N_5544,N_6753);
nand U9645 (N_9645,N_5130,N_6299);
or U9646 (N_9646,N_7083,N_5373);
nor U9647 (N_9647,N_6028,N_5166);
nand U9648 (N_9648,N_7014,N_6893);
xor U9649 (N_9649,N_5996,N_5534);
and U9650 (N_9650,N_5455,N_5523);
nand U9651 (N_9651,N_5372,N_5739);
nor U9652 (N_9652,N_5454,N_6213);
xor U9653 (N_9653,N_5594,N_7114);
xor U9654 (N_9654,N_6507,N_6406);
nor U9655 (N_9655,N_5418,N_7372);
xnor U9656 (N_9656,N_7021,N_5499);
nand U9657 (N_9657,N_6789,N_5692);
and U9658 (N_9658,N_6835,N_6959);
nor U9659 (N_9659,N_5582,N_6464);
nand U9660 (N_9660,N_7032,N_5914);
nor U9661 (N_9661,N_5572,N_5549);
and U9662 (N_9662,N_7483,N_6420);
and U9663 (N_9663,N_6337,N_7188);
nand U9664 (N_9664,N_6071,N_5190);
nand U9665 (N_9665,N_5854,N_7356);
xnor U9666 (N_9666,N_7359,N_5457);
nor U9667 (N_9667,N_6486,N_5822);
or U9668 (N_9668,N_5124,N_6299);
or U9669 (N_9669,N_5172,N_5541);
xor U9670 (N_9670,N_6719,N_6683);
nor U9671 (N_9671,N_5833,N_6648);
nand U9672 (N_9672,N_6362,N_5393);
nor U9673 (N_9673,N_5871,N_6044);
nor U9674 (N_9674,N_5388,N_6004);
nand U9675 (N_9675,N_6628,N_6697);
or U9676 (N_9676,N_7118,N_5631);
xor U9677 (N_9677,N_6140,N_7235);
nand U9678 (N_9678,N_7006,N_6854);
nor U9679 (N_9679,N_6302,N_7158);
or U9680 (N_9680,N_5939,N_6488);
and U9681 (N_9681,N_5885,N_6326);
nand U9682 (N_9682,N_6105,N_7211);
nand U9683 (N_9683,N_6681,N_6043);
xnor U9684 (N_9684,N_7320,N_5379);
xor U9685 (N_9685,N_6804,N_6749);
and U9686 (N_9686,N_7397,N_7267);
xnor U9687 (N_9687,N_6796,N_5408);
nand U9688 (N_9688,N_6026,N_7472);
nand U9689 (N_9689,N_6991,N_6323);
and U9690 (N_9690,N_5118,N_7462);
and U9691 (N_9691,N_6269,N_6268);
and U9692 (N_9692,N_6368,N_7010);
or U9693 (N_9693,N_6731,N_7469);
nor U9694 (N_9694,N_6705,N_5349);
and U9695 (N_9695,N_5163,N_7274);
nand U9696 (N_9696,N_6746,N_6357);
or U9697 (N_9697,N_5894,N_7433);
nand U9698 (N_9698,N_6349,N_5355);
nor U9699 (N_9699,N_5089,N_5714);
nor U9700 (N_9700,N_6723,N_5366);
nand U9701 (N_9701,N_7341,N_6380);
and U9702 (N_9702,N_7003,N_5022);
nor U9703 (N_9703,N_6239,N_6306);
nand U9704 (N_9704,N_5932,N_5070);
nand U9705 (N_9705,N_7231,N_6615);
xor U9706 (N_9706,N_6491,N_5308);
xnor U9707 (N_9707,N_5722,N_5583);
or U9708 (N_9708,N_6993,N_5705);
or U9709 (N_9709,N_5061,N_6828);
or U9710 (N_9710,N_5489,N_6016);
and U9711 (N_9711,N_5440,N_5201);
nor U9712 (N_9712,N_7443,N_5212);
nand U9713 (N_9713,N_5514,N_6024);
nor U9714 (N_9714,N_6974,N_5110);
nor U9715 (N_9715,N_6353,N_5393);
or U9716 (N_9716,N_6285,N_6910);
nand U9717 (N_9717,N_6933,N_5056);
and U9718 (N_9718,N_5865,N_5657);
nand U9719 (N_9719,N_5643,N_7110);
nand U9720 (N_9720,N_5599,N_5014);
or U9721 (N_9721,N_5696,N_7357);
nor U9722 (N_9722,N_6049,N_5547);
nand U9723 (N_9723,N_6312,N_5064);
xnor U9724 (N_9724,N_6326,N_5613);
nor U9725 (N_9725,N_5999,N_5615);
nand U9726 (N_9726,N_6508,N_5984);
xnor U9727 (N_9727,N_6283,N_6792);
and U9728 (N_9728,N_5251,N_5363);
or U9729 (N_9729,N_6826,N_5606);
and U9730 (N_9730,N_6489,N_5877);
or U9731 (N_9731,N_7211,N_6725);
nor U9732 (N_9732,N_5886,N_6330);
and U9733 (N_9733,N_5646,N_5201);
xor U9734 (N_9734,N_5418,N_7135);
nand U9735 (N_9735,N_5108,N_5121);
nand U9736 (N_9736,N_6556,N_5567);
nand U9737 (N_9737,N_7487,N_6387);
nor U9738 (N_9738,N_5375,N_6812);
xor U9739 (N_9739,N_5926,N_7281);
nor U9740 (N_9740,N_5586,N_6969);
xor U9741 (N_9741,N_6645,N_5046);
or U9742 (N_9742,N_6864,N_6195);
nand U9743 (N_9743,N_5022,N_5773);
xor U9744 (N_9744,N_6041,N_6972);
xnor U9745 (N_9745,N_5435,N_5218);
nand U9746 (N_9746,N_6956,N_7083);
and U9747 (N_9747,N_7346,N_7448);
xnor U9748 (N_9748,N_5997,N_6644);
or U9749 (N_9749,N_5526,N_6075);
xnor U9750 (N_9750,N_5692,N_5547);
xor U9751 (N_9751,N_6182,N_5386);
or U9752 (N_9752,N_5546,N_6614);
or U9753 (N_9753,N_5776,N_6276);
and U9754 (N_9754,N_6530,N_6966);
or U9755 (N_9755,N_5915,N_6396);
nor U9756 (N_9756,N_6411,N_5530);
nand U9757 (N_9757,N_5788,N_7193);
xnor U9758 (N_9758,N_6156,N_5822);
or U9759 (N_9759,N_6002,N_5190);
nand U9760 (N_9760,N_6082,N_6578);
nand U9761 (N_9761,N_7284,N_5404);
and U9762 (N_9762,N_6674,N_5039);
xnor U9763 (N_9763,N_5819,N_7066);
and U9764 (N_9764,N_6664,N_5217);
nor U9765 (N_9765,N_5508,N_5915);
xnor U9766 (N_9766,N_5323,N_6457);
nand U9767 (N_9767,N_5052,N_5138);
or U9768 (N_9768,N_5915,N_5291);
or U9769 (N_9769,N_5514,N_6057);
nor U9770 (N_9770,N_6468,N_6176);
and U9771 (N_9771,N_5944,N_5916);
nand U9772 (N_9772,N_7192,N_7041);
and U9773 (N_9773,N_7112,N_5652);
nor U9774 (N_9774,N_6702,N_5999);
nand U9775 (N_9775,N_6759,N_5281);
nand U9776 (N_9776,N_7182,N_6735);
xnor U9777 (N_9777,N_7209,N_6587);
nand U9778 (N_9778,N_5679,N_6865);
xnor U9779 (N_9779,N_6783,N_7285);
and U9780 (N_9780,N_5938,N_5802);
nor U9781 (N_9781,N_6980,N_7462);
nor U9782 (N_9782,N_6614,N_5267);
and U9783 (N_9783,N_5172,N_6587);
nand U9784 (N_9784,N_5150,N_6504);
nand U9785 (N_9785,N_5480,N_7276);
or U9786 (N_9786,N_6633,N_7357);
nand U9787 (N_9787,N_5526,N_6703);
and U9788 (N_9788,N_5790,N_6089);
and U9789 (N_9789,N_5569,N_7042);
or U9790 (N_9790,N_7364,N_5745);
or U9791 (N_9791,N_5009,N_7150);
or U9792 (N_9792,N_5164,N_5313);
nor U9793 (N_9793,N_7258,N_6660);
or U9794 (N_9794,N_6318,N_5512);
xnor U9795 (N_9795,N_6826,N_6523);
nand U9796 (N_9796,N_7009,N_5733);
nand U9797 (N_9797,N_5376,N_5150);
or U9798 (N_9798,N_5508,N_6673);
nor U9799 (N_9799,N_6338,N_6989);
nand U9800 (N_9800,N_7443,N_5686);
or U9801 (N_9801,N_6049,N_7167);
and U9802 (N_9802,N_6061,N_6615);
nor U9803 (N_9803,N_5593,N_6758);
or U9804 (N_9804,N_6557,N_5281);
nand U9805 (N_9805,N_5408,N_5132);
and U9806 (N_9806,N_5760,N_6112);
and U9807 (N_9807,N_7312,N_7243);
or U9808 (N_9808,N_7495,N_6345);
and U9809 (N_9809,N_5112,N_5555);
nand U9810 (N_9810,N_5897,N_5811);
nor U9811 (N_9811,N_6911,N_5098);
and U9812 (N_9812,N_5044,N_6934);
nand U9813 (N_9813,N_7089,N_6178);
nor U9814 (N_9814,N_6590,N_6230);
nand U9815 (N_9815,N_6214,N_7262);
nor U9816 (N_9816,N_7011,N_5853);
nor U9817 (N_9817,N_5571,N_6563);
and U9818 (N_9818,N_7131,N_5878);
and U9819 (N_9819,N_6740,N_6105);
or U9820 (N_9820,N_5039,N_6316);
nor U9821 (N_9821,N_5249,N_6845);
and U9822 (N_9822,N_6113,N_7305);
nor U9823 (N_9823,N_7251,N_5268);
and U9824 (N_9824,N_6090,N_6059);
xor U9825 (N_9825,N_5579,N_5750);
or U9826 (N_9826,N_7494,N_5774);
nor U9827 (N_9827,N_7037,N_6142);
nand U9828 (N_9828,N_7005,N_5263);
xor U9829 (N_9829,N_6106,N_7188);
nor U9830 (N_9830,N_6229,N_6614);
or U9831 (N_9831,N_5006,N_7116);
or U9832 (N_9832,N_6518,N_7293);
xnor U9833 (N_9833,N_7395,N_6044);
xnor U9834 (N_9834,N_5606,N_5459);
nor U9835 (N_9835,N_5785,N_6831);
nand U9836 (N_9836,N_7097,N_5492);
nor U9837 (N_9837,N_7200,N_6848);
xnor U9838 (N_9838,N_6998,N_7320);
nand U9839 (N_9839,N_5795,N_5727);
or U9840 (N_9840,N_5130,N_7463);
nand U9841 (N_9841,N_6355,N_5360);
nand U9842 (N_9842,N_5925,N_6339);
or U9843 (N_9843,N_6305,N_5399);
nand U9844 (N_9844,N_5563,N_6663);
xor U9845 (N_9845,N_7258,N_5314);
nor U9846 (N_9846,N_5190,N_7464);
nor U9847 (N_9847,N_5099,N_5109);
and U9848 (N_9848,N_6289,N_5430);
and U9849 (N_9849,N_6530,N_5505);
nand U9850 (N_9850,N_7324,N_7328);
or U9851 (N_9851,N_5483,N_7073);
and U9852 (N_9852,N_6918,N_6626);
and U9853 (N_9853,N_6083,N_6637);
xor U9854 (N_9854,N_5151,N_6189);
or U9855 (N_9855,N_6021,N_5578);
or U9856 (N_9856,N_5726,N_5277);
nor U9857 (N_9857,N_7110,N_7460);
xnor U9858 (N_9858,N_6536,N_5479);
or U9859 (N_9859,N_5402,N_5251);
nand U9860 (N_9860,N_5402,N_6217);
xnor U9861 (N_9861,N_7071,N_7213);
or U9862 (N_9862,N_7047,N_6388);
or U9863 (N_9863,N_7125,N_5888);
or U9864 (N_9864,N_7200,N_6123);
nand U9865 (N_9865,N_5830,N_7435);
nand U9866 (N_9866,N_7464,N_5497);
and U9867 (N_9867,N_6015,N_6520);
and U9868 (N_9868,N_5482,N_6658);
and U9869 (N_9869,N_7071,N_5024);
xnor U9870 (N_9870,N_6787,N_5063);
nor U9871 (N_9871,N_7188,N_5034);
nor U9872 (N_9872,N_5926,N_6267);
and U9873 (N_9873,N_6366,N_6924);
nand U9874 (N_9874,N_5603,N_5590);
and U9875 (N_9875,N_6865,N_5755);
nor U9876 (N_9876,N_5054,N_6391);
xor U9877 (N_9877,N_5761,N_5253);
xor U9878 (N_9878,N_5187,N_7393);
xnor U9879 (N_9879,N_5302,N_6516);
nand U9880 (N_9880,N_5590,N_5213);
or U9881 (N_9881,N_6932,N_6209);
and U9882 (N_9882,N_6130,N_6084);
nand U9883 (N_9883,N_7022,N_5101);
xnor U9884 (N_9884,N_6835,N_7153);
nor U9885 (N_9885,N_6974,N_6075);
xor U9886 (N_9886,N_5174,N_5989);
xnor U9887 (N_9887,N_5067,N_6713);
xnor U9888 (N_9888,N_7440,N_5156);
or U9889 (N_9889,N_7094,N_5849);
xnor U9890 (N_9890,N_6591,N_7351);
nand U9891 (N_9891,N_6135,N_5699);
nor U9892 (N_9892,N_6392,N_6183);
and U9893 (N_9893,N_6416,N_5829);
and U9894 (N_9894,N_5231,N_5230);
and U9895 (N_9895,N_6565,N_5591);
or U9896 (N_9896,N_5653,N_5394);
nor U9897 (N_9897,N_5438,N_5068);
and U9898 (N_9898,N_5508,N_6217);
or U9899 (N_9899,N_6911,N_5954);
nor U9900 (N_9900,N_5081,N_6799);
xnor U9901 (N_9901,N_5627,N_5049);
xnor U9902 (N_9902,N_7265,N_6834);
xnor U9903 (N_9903,N_7437,N_5298);
and U9904 (N_9904,N_7388,N_6405);
and U9905 (N_9905,N_5823,N_6043);
or U9906 (N_9906,N_7471,N_6606);
or U9907 (N_9907,N_6193,N_5818);
or U9908 (N_9908,N_5117,N_6567);
nand U9909 (N_9909,N_5536,N_7294);
and U9910 (N_9910,N_5858,N_6262);
nand U9911 (N_9911,N_6701,N_5574);
and U9912 (N_9912,N_6470,N_5160);
nand U9913 (N_9913,N_6848,N_6473);
xnor U9914 (N_9914,N_6942,N_5122);
nand U9915 (N_9915,N_7059,N_6667);
or U9916 (N_9916,N_6579,N_5950);
or U9917 (N_9917,N_6278,N_5194);
nand U9918 (N_9918,N_5734,N_5217);
nand U9919 (N_9919,N_6935,N_5434);
xnor U9920 (N_9920,N_6413,N_5681);
and U9921 (N_9921,N_6725,N_6014);
or U9922 (N_9922,N_6687,N_5197);
nand U9923 (N_9923,N_5441,N_6518);
or U9924 (N_9924,N_6510,N_7334);
and U9925 (N_9925,N_5342,N_5693);
nand U9926 (N_9926,N_5875,N_6404);
xor U9927 (N_9927,N_6150,N_6045);
xor U9928 (N_9928,N_6932,N_5700);
and U9929 (N_9929,N_7282,N_5950);
nand U9930 (N_9930,N_6545,N_6315);
or U9931 (N_9931,N_6741,N_6026);
xor U9932 (N_9932,N_5232,N_5913);
nand U9933 (N_9933,N_6296,N_7354);
or U9934 (N_9934,N_7009,N_5429);
xnor U9935 (N_9935,N_5390,N_7438);
and U9936 (N_9936,N_5560,N_5646);
nand U9937 (N_9937,N_7240,N_6450);
and U9938 (N_9938,N_5804,N_7321);
nor U9939 (N_9939,N_6241,N_5730);
nor U9940 (N_9940,N_6930,N_5363);
or U9941 (N_9941,N_5284,N_5857);
and U9942 (N_9942,N_6755,N_7334);
or U9943 (N_9943,N_5491,N_7168);
nand U9944 (N_9944,N_7283,N_5674);
nand U9945 (N_9945,N_6087,N_5357);
nor U9946 (N_9946,N_5881,N_6778);
nand U9947 (N_9947,N_6269,N_6091);
nor U9948 (N_9948,N_5986,N_6243);
and U9949 (N_9949,N_5366,N_6380);
xnor U9950 (N_9950,N_7480,N_5064);
or U9951 (N_9951,N_5708,N_6619);
or U9952 (N_9952,N_5806,N_6113);
and U9953 (N_9953,N_5396,N_5422);
or U9954 (N_9954,N_7004,N_5301);
and U9955 (N_9955,N_5627,N_5864);
and U9956 (N_9956,N_5828,N_6334);
and U9957 (N_9957,N_6801,N_6558);
nand U9958 (N_9958,N_5484,N_5643);
or U9959 (N_9959,N_7388,N_5289);
or U9960 (N_9960,N_7450,N_6039);
nor U9961 (N_9961,N_6337,N_5367);
and U9962 (N_9962,N_6572,N_6221);
and U9963 (N_9963,N_7183,N_5604);
xnor U9964 (N_9964,N_7400,N_7106);
nand U9965 (N_9965,N_5331,N_6121);
or U9966 (N_9966,N_5154,N_5094);
nor U9967 (N_9967,N_7041,N_7412);
xnor U9968 (N_9968,N_6900,N_5636);
or U9969 (N_9969,N_6232,N_5332);
nand U9970 (N_9970,N_7126,N_7392);
nand U9971 (N_9971,N_6711,N_6952);
nand U9972 (N_9972,N_5747,N_5949);
nand U9973 (N_9973,N_5091,N_5536);
xor U9974 (N_9974,N_7267,N_6203);
and U9975 (N_9975,N_7088,N_5315);
and U9976 (N_9976,N_5312,N_6884);
nor U9977 (N_9977,N_5329,N_5650);
xnor U9978 (N_9978,N_6959,N_6146);
nand U9979 (N_9979,N_5480,N_6793);
xnor U9980 (N_9980,N_5228,N_5949);
nand U9981 (N_9981,N_6537,N_6116);
nand U9982 (N_9982,N_6630,N_6795);
nand U9983 (N_9983,N_5862,N_5273);
xor U9984 (N_9984,N_5245,N_6557);
and U9985 (N_9985,N_6872,N_6212);
and U9986 (N_9986,N_5308,N_7181);
or U9987 (N_9987,N_5585,N_6079);
and U9988 (N_9988,N_7318,N_6434);
nand U9989 (N_9989,N_6618,N_6383);
xor U9990 (N_9990,N_6510,N_7303);
nor U9991 (N_9991,N_5054,N_6029);
nor U9992 (N_9992,N_6537,N_5086);
and U9993 (N_9993,N_6302,N_6775);
or U9994 (N_9994,N_5793,N_5805);
or U9995 (N_9995,N_5721,N_6453);
or U9996 (N_9996,N_5297,N_6834);
xor U9997 (N_9997,N_7090,N_7189);
xnor U9998 (N_9998,N_7286,N_5043);
xor U9999 (N_9999,N_5314,N_5707);
or U10000 (N_10000,N_9048,N_8286);
nor U10001 (N_10001,N_9266,N_8580);
nor U10002 (N_10002,N_8787,N_8987);
nor U10003 (N_10003,N_8860,N_7678);
and U10004 (N_10004,N_8422,N_7972);
or U10005 (N_10005,N_7845,N_9739);
and U10006 (N_10006,N_8471,N_8125);
and U10007 (N_10007,N_7979,N_9433);
nand U10008 (N_10008,N_8674,N_7648);
and U10009 (N_10009,N_7987,N_9638);
xor U10010 (N_10010,N_9170,N_9618);
xor U10011 (N_10011,N_9846,N_9591);
xor U10012 (N_10012,N_8963,N_9222);
and U10013 (N_10013,N_7771,N_9627);
and U10014 (N_10014,N_8306,N_9341);
xnor U10015 (N_10015,N_9430,N_9242);
nand U10016 (N_10016,N_7581,N_7576);
xnor U10017 (N_10017,N_9223,N_9611);
and U10018 (N_10018,N_9181,N_8549);
and U10019 (N_10019,N_7900,N_9561);
nand U10020 (N_10020,N_8999,N_7811);
or U10021 (N_10021,N_9677,N_8486);
or U10022 (N_10022,N_9533,N_8344);
or U10023 (N_10023,N_8560,N_9473);
or U10024 (N_10024,N_8161,N_9752);
nand U10025 (N_10025,N_8059,N_8098);
nor U10026 (N_10026,N_9052,N_9687);
and U10027 (N_10027,N_9096,N_8715);
or U10028 (N_10028,N_8440,N_8666);
nor U10029 (N_10029,N_9393,N_8792);
nand U10030 (N_10030,N_8983,N_9570);
or U10031 (N_10031,N_8158,N_8922);
nor U10032 (N_10032,N_8193,N_8940);
and U10033 (N_10033,N_8510,N_8022);
and U10034 (N_10034,N_9690,N_8961);
and U10035 (N_10035,N_7695,N_8620);
or U10036 (N_10036,N_8200,N_8701);
xor U10037 (N_10037,N_8507,N_9523);
nor U10038 (N_10038,N_9244,N_8959);
or U10039 (N_10039,N_9005,N_7716);
nor U10040 (N_10040,N_9596,N_9312);
nor U10041 (N_10041,N_8622,N_8968);
and U10042 (N_10042,N_8206,N_8250);
nand U10043 (N_10043,N_8449,N_9708);
or U10044 (N_10044,N_9858,N_8530);
and U10045 (N_10045,N_9108,N_7999);
and U10046 (N_10046,N_7705,N_8166);
nor U10047 (N_10047,N_8347,N_8085);
and U10048 (N_10048,N_9094,N_9289);
and U10049 (N_10049,N_9324,N_8176);
or U10050 (N_10050,N_8266,N_8757);
or U10051 (N_10051,N_7502,N_8242);
nor U10052 (N_10052,N_8838,N_8769);
and U10053 (N_10053,N_9540,N_8577);
xor U10054 (N_10054,N_9162,N_8993);
and U10055 (N_10055,N_9435,N_8481);
xor U10056 (N_10056,N_7674,N_7807);
xor U10057 (N_10057,N_9432,N_9890);
and U10058 (N_10058,N_8677,N_8755);
and U10059 (N_10059,N_8177,N_9123);
nand U10060 (N_10060,N_7616,N_8590);
or U10061 (N_10061,N_9977,N_9097);
nor U10062 (N_10062,N_9002,N_9198);
or U10063 (N_10063,N_8205,N_9179);
nand U10064 (N_10064,N_7608,N_8061);
xor U10065 (N_10065,N_8776,N_7518);
xor U10066 (N_10066,N_9817,N_8605);
or U10067 (N_10067,N_7967,N_8474);
or U10068 (N_10068,N_9125,N_7683);
or U10069 (N_10069,N_8942,N_9200);
nand U10070 (N_10070,N_9345,N_9558);
xnor U10071 (N_10071,N_9325,N_7762);
nand U10072 (N_10072,N_9499,N_9417);
and U10073 (N_10073,N_7927,N_9042);
and U10074 (N_10074,N_8941,N_8339);
xnor U10075 (N_10075,N_8844,N_9806);
nor U10076 (N_10076,N_9247,N_8656);
nand U10077 (N_10077,N_9751,N_8662);
nor U10078 (N_10078,N_8433,N_9330);
or U10079 (N_10079,N_7799,N_7692);
xor U10080 (N_10080,N_8456,N_9472);
or U10081 (N_10081,N_7739,N_9762);
nand U10082 (N_10082,N_9347,N_7530);
or U10083 (N_10083,N_7968,N_9518);
nor U10084 (N_10084,N_8178,N_7991);
xor U10085 (N_10085,N_7669,N_9950);
nor U10086 (N_10086,N_8635,N_7862);
or U10087 (N_10087,N_8774,N_8589);
nor U10088 (N_10088,N_8964,N_8824);
nor U10089 (N_10089,N_9655,N_9623);
or U10090 (N_10090,N_7889,N_8329);
and U10091 (N_10091,N_9863,N_9144);
and U10092 (N_10092,N_8257,N_9311);
or U10093 (N_10093,N_9342,N_8670);
or U10094 (N_10094,N_8739,N_8434);
nor U10095 (N_10095,N_9254,N_9470);
or U10096 (N_10096,N_9485,N_9383);
nand U10097 (N_10097,N_9018,N_8529);
nand U10098 (N_10098,N_9665,N_8279);
nand U10099 (N_10099,N_7569,N_9530);
and U10100 (N_10100,N_8508,N_8187);
or U10101 (N_10101,N_7788,N_9861);
nand U10102 (N_10102,N_9423,N_8336);
nand U10103 (N_10103,N_7687,N_8626);
nand U10104 (N_10104,N_9166,N_7712);
nand U10105 (N_10105,N_9625,N_8520);
nor U10106 (N_10106,N_9074,N_8249);
xor U10107 (N_10107,N_7601,N_7599);
nor U10108 (N_10108,N_9446,N_7522);
xor U10109 (N_10109,N_8730,N_9425);
xor U10110 (N_10110,N_7745,N_7540);
and U10111 (N_10111,N_9562,N_9259);
or U10112 (N_10112,N_8684,N_9700);
xor U10113 (N_10113,N_8986,N_9648);
nand U10114 (N_10114,N_9673,N_9698);
nor U10115 (N_10115,N_9497,N_9974);
xnor U10116 (N_10116,N_7768,N_8174);
nand U10117 (N_10117,N_9969,N_9990);
xor U10118 (N_10118,N_8621,N_9051);
xor U10119 (N_10119,N_8858,N_8136);
nand U10120 (N_10120,N_9337,N_7717);
nor U10121 (N_10121,N_9501,N_8705);
nand U10122 (N_10122,N_8687,N_9017);
or U10123 (N_10123,N_8394,N_7864);
or U10124 (N_10124,N_8293,N_9185);
and U10125 (N_10125,N_8618,N_7930);
nand U10126 (N_10126,N_8221,N_8021);
nor U10127 (N_10127,N_9122,N_8294);
nand U10128 (N_10128,N_9458,N_8568);
nor U10129 (N_10129,N_8540,N_9882);
nand U10130 (N_10130,N_9091,N_9686);
nor U10131 (N_10131,N_9927,N_8606);
and U10132 (N_10132,N_8832,N_8634);
xor U10133 (N_10133,N_8199,N_9715);
or U10134 (N_10134,N_7849,N_9934);
or U10135 (N_10135,N_9394,N_9864);
and U10136 (N_10136,N_9609,N_7587);
or U10137 (N_10137,N_9055,N_8823);
or U10138 (N_10138,N_9025,N_7758);
nor U10139 (N_10139,N_9692,N_8132);
nand U10140 (N_10140,N_8967,N_7760);
xnor U10141 (N_10141,N_9366,N_8041);
and U10142 (N_10142,N_9845,N_7996);
and U10143 (N_10143,N_8298,N_8804);
nand U10144 (N_10144,N_9954,N_9187);
or U10145 (N_10145,N_8040,N_8361);
or U10146 (N_10146,N_9824,N_7598);
xor U10147 (N_10147,N_9046,N_8383);
xor U10148 (N_10148,N_9675,N_7664);
xnor U10149 (N_10149,N_9488,N_8359);
and U10150 (N_10150,N_7945,N_7812);
nor U10151 (N_10151,N_8420,N_8430);
nor U10152 (N_10152,N_9389,N_8454);
nand U10153 (N_10153,N_9422,N_9288);
or U10154 (N_10154,N_8495,N_8297);
nand U10155 (N_10155,N_7868,N_9644);
xor U10156 (N_10156,N_8090,N_8794);
or U10157 (N_10157,N_9742,N_9361);
nor U10158 (N_10158,N_8065,N_8853);
nand U10159 (N_10159,N_9968,N_8018);
nor U10160 (N_10160,N_7986,N_8623);
nand U10161 (N_10161,N_8747,N_9953);
or U10162 (N_10162,N_9998,N_8204);
xnor U10163 (N_10163,N_8013,N_9886);
nand U10164 (N_10164,N_9993,N_9997);
nor U10165 (N_10165,N_8107,N_7850);
nor U10166 (N_10166,N_8489,N_8732);
nand U10167 (N_10167,N_9822,N_8720);
xnor U10168 (N_10168,N_8355,N_9286);
or U10169 (N_10169,N_8324,N_8814);
and U10170 (N_10170,N_9117,N_7854);
xor U10171 (N_10171,N_7858,N_8783);
and U10172 (N_10172,N_7514,N_9201);
nor U10173 (N_10173,N_9032,N_9368);
nor U10174 (N_10174,N_8856,N_9078);
or U10175 (N_10175,N_9028,N_7702);
nand U10176 (N_10176,N_7617,N_7652);
and U10177 (N_10177,N_7912,N_7506);
nand U10178 (N_10178,N_9169,N_9320);
and U10179 (N_10179,N_9981,N_8005);
or U10180 (N_10180,N_9976,N_9471);
and U10181 (N_10181,N_9722,N_9946);
nand U10182 (N_10182,N_8716,N_8464);
nor U10183 (N_10183,N_9474,N_8068);
nor U10184 (N_10184,N_8307,N_8810);
nor U10185 (N_10185,N_8570,N_7528);
nand U10186 (N_10186,N_9679,N_8503);
xnor U10187 (N_10187,N_9702,N_8937);
or U10188 (N_10188,N_8772,N_9328);
and U10189 (N_10189,N_7763,N_8582);
xnor U10190 (N_10190,N_7538,N_8323);
xor U10191 (N_10191,N_9711,N_9348);
xnor U10192 (N_10192,N_7672,N_7846);
nor U10193 (N_10193,N_7646,N_8110);
or U10194 (N_10194,N_8567,N_8170);
xnor U10195 (N_10195,N_9036,N_9230);
nor U10196 (N_10196,N_8271,N_8548);
xnor U10197 (N_10197,N_8609,N_9957);
or U10198 (N_10198,N_7696,N_9888);
and U10199 (N_10199,N_9691,N_9826);
nand U10200 (N_10200,N_8402,N_9402);
and U10201 (N_10201,N_9867,N_7657);
nand U10202 (N_10202,N_8375,N_7767);
nand U10203 (N_10203,N_9588,N_8809);
or U10204 (N_10204,N_9447,N_9418);
nand U10205 (N_10205,N_7611,N_8534);
xor U10206 (N_10206,N_8863,N_9829);
nand U10207 (N_10207,N_8706,N_7837);
or U10208 (N_10208,N_9904,N_8699);
xor U10209 (N_10209,N_8074,N_9924);
or U10210 (N_10210,N_7690,N_9479);
or U10211 (N_10211,N_7805,N_9140);
nor U10212 (N_10212,N_8274,N_8815);
nand U10213 (N_10213,N_8943,N_8697);
or U10214 (N_10214,N_8921,N_8997);
nand U10215 (N_10215,N_8789,N_8139);
and U10216 (N_10216,N_9725,N_7531);
nand U10217 (N_10217,N_9965,N_7755);
nand U10218 (N_10218,N_8953,N_9830);
xnor U10219 (N_10219,N_9438,N_9131);
nor U10220 (N_10220,N_8599,N_9955);
nand U10221 (N_10221,N_7627,N_9597);
and U10222 (N_10222,N_9630,N_9468);
nor U10223 (N_10223,N_9874,N_7764);
xor U10224 (N_10224,N_9548,N_8015);
xor U10225 (N_10225,N_9941,N_8835);
and U10226 (N_10226,N_8436,N_7951);
and U10227 (N_10227,N_9825,N_9719);
xor U10228 (N_10228,N_9424,N_9916);
nor U10229 (N_10229,N_9411,N_9039);
and U10230 (N_10230,N_8254,N_8868);
and U10231 (N_10231,N_8321,N_8962);
and U10232 (N_10232,N_7824,N_9378);
nor U10233 (N_10233,N_9478,N_9788);
or U10234 (N_10234,N_7668,N_9121);
nor U10235 (N_10235,N_9219,N_9569);
and U10236 (N_10236,N_8252,N_9631);
and U10237 (N_10237,N_7644,N_9521);
nand U10238 (N_10238,N_9452,N_9847);
and U10239 (N_10239,N_8553,N_8437);
xor U10240 (N_10240,N_9188,N_8255);
xor U10241 (N_10241,N_8358,N_8591);
xor U10242 (N_10242,N_7981,N_9186);
xnor U10243 (N_10243,N_9009,N_7711);
nor U10244 (N_10244,N_7728,N_8100);
nand U10245 (N_10245,N_8401,N_9126);
and U10246 (N_10246,N_8105,N_9582);
or U10247 (N_10247,N_8146,N_8979);
or U10248 (N_10248,N_8388,N_9877);
nor U10249 (N_10249,N_8588,N_9544);
and U10250 (N_10250,N_9619,N_9915);
or U10251 (N_10251,N_7628,N_8082);
or U10252 (N_10252,N_8412,N_8104);
nor U10253 (N_10253,N_8494,N_9607);
nand U10254 (N_10254,N_8632,N_8882);
or U10255 (N_10255,N_9054,N_9833);
nor U10256 (N_10256,N_8496,N_8506);
nand U10257 (N_10257,N_8539,N_8444);
and U10258 (N_10258,N_7806,N_9217);
or U10259 (N_10259,N_8688,N_9111);
and U10260 (N_10260,N_8598,N_8554);
and U10261 (N_10261,N_8122,N_8314);
xnor U10262 (N_10262,N_9891,N_8129);
xnor U10263 (N_10263,N_8463,N_9620);
xnor U10264 (N_10264,N_8010,N_8583);
and U10265 (N_10265,N_7567,N_8169);
or U10266 (N_10266,N_9212,N_8807);
nor U10267 (N_10267,N_8517,N_9081);
or U10268 (N_10268,N_8859,N_9705);
nand U10269 (N_10269,N_7590,N_7777);
or U10270 (N_10270,N_7833,N_7719);
or U10271 (N_10271,N_9395,N_9158);
or U10272 (N_10272,N_9937,N_8043);
nor U10273 (N_10273,N_8285,N_8846);
nor U10274 (N_10274,N_7978,N_8754);
xnor U10275 (N_10275,N_9871,N_8528);
and U10276 (N_10276,N_9792,N_9130);
nor U10277 (N_10277,N_8902,N_8681);
nand U10278 (N_10278,N_9203,N_9405);
xor U10279 (N_10279,N_8818,N_8400);
xnor U10280 (N_10280,N_9109,N_9962);
nor U10281 (N_10281,N_9783,N_8502);
xor U10282 (N_10282,N_9951,N_7625);
xor U10283 (N_10283,N_8133,N_9717);
or U10284 (N_10284,N_8011,N_8111);
nor U10285 (N_10285,N_9593,N_9355);
and U10286 (N_10286,N_7899,N_9085);
nand U10287 (N_10287,N_7896,N_9994);
and U10288 (N_10288,N_9214,N_9309);
xnor U10289 (N_10289,N_8864,N_9336);
nor U10290 (N_10290,N_8320,N_8470);
nor U10291 (N_10291,N_8201,N_7752);
and U10292 (N_10292,N_7722,N_9106);
or U10293 (N_10293,N_7640,N_9145);
and U10294 (N_10294,N_9746,N_9240);
xor U10295 (N_10295,N_7675,N_8908);
and U10296 (N_10296,N_8511,N_7756);
nor U10297 (N_10297,N_8417,N_7516);
nand U10298 (N_10298,N_7781,N_9089);
nand U10299 (N_10299,N_9606,N_8340);
xnor U10300 (N_10300,N_8092,N_9498);
or U10301 (N_10301,N_9728,N_8322);
nand U10302 (N_10302,N_9989,N_8647);
or U10303 (N_10303,N_8801,N_9160);
or U10304 (N_10304,N_8871,N_9495);
nor U10305 (N_10305,N_9584,N_9730);
xnor U10306 (N_10306,N_9409,N_9876);
xor U10307 (N_10307,N_9204,N_7857);
nor U10308 (N_10308,N_9386,N_7708);
nand U10309 (N_10309,N_7609,N_9729);
nor U10310 (N_10310,N_9525,N_9813);
nor U10311 (N_10311,N_9503,N_8270);
and U10312 (N_10312,N_9800,N_9734);
and U10313 (N_10313,N_8207,N_8602);
nand U10314 (N_10314,N_8172,N_9044);
nor U10315 (N_10315,N_7524,N_8382);
nand U10316 (N_10316,N_9804,N_9765);
or U10317 (N_10317,N_9727,N_8991);
or U10318 (N_10318,N_8876,N_9269);
and U10319 (N_10319,N_8645,N_7888);
nand U10320 (N_10320,N_9547,N_8160);
and U10321 (N_10321,N_9546,N_9972);
or U10322 (N_10322,N_9587,N_8042);
or U10323 (N_10323,N_9785,N_9413);
nand U10324 (N_10324,N_9092,N_8728);
xor U10325 (N_10325,N_9477,N_9577);
xnor U10326 (N_10326,N_7691,N_9150);
nor U10327 (N_10327,N_9480,N_9694);
and U10328 (N_10328,N_9787,N_8096);
and U10329 (N_10329,N_8938,N_7729);
or U10330 (N_10330,N_8182,N_8406);
xor U10331 (N_10331,N_7950,N_8302);
or U10332 (N_10332,N_8998,N_8989);
nand U10333 (N_10333,N_8350,N_8793);
and U10334 (N_10334,N_8753,N_8919);
and U10335 (N_10335,N_8235,N_9881);
or U10336 (N_10336,N_9322,N_7940);
xor U10337 (N_10337,N_7926,N_9724);
xnor U10338 (N_10338,N_7801,N_8779);
xnor U10339 (N_10339,N_8897,N_9592);
nor U10340 (N_10340,N_8183,N_8453);
nor U10341 (N_10341,N_8229,N_9349);
nor U10342 (N_10342,N_9563,N_9878);
xor U10343 (N_10343,N_8230,N_9772);
or U10344 (N_10344,N_8156,N_9559);
xnor U10345 (N_10345,N_9918,N_8037);
and U10346 (N_10346,N_7882,N_8671);
xor U10347 (N_10347,N_8682,N_7544);
and U10348 (N_10348,N_9731,N_9098);
and U10349 (N_10349,N_8181,N_8368);
nand U10350 (N_10350,N_7875,N_9766);
and U10351 (N_10351,N_8218,N_8773);
nor U10352 (N_10352,N_9683,N_9524);
xnor U10353 (N_10353,N_8708,N_8016);
nand U10354 (N_10354,N_8265,N_8084);
nand U10355 (N_10355,N_8829,N_7580);
nand U10356 (N_10356,N_7543,N_9791);
nor U10357 (N_10357,N_8912,N_9531);
xor U10358 (N_10358,N_7759,N_8544);
xnor U10359 (N_10359,N_8654,N_7953);
or U10360 (N_10360,N_8480,N_8364);
or U10361 (N_10361,N_8223,N_9670);
xor U10362 (N_10362,N_8492,N_8811);
nand U10363 (N_10363,N_9022,N_7954);
nor U10364 (N_10364,N_8079,N_9385);
xor U10365 (N_10365,N_9963,N_7521);
and U10366 (N_10366,N_9760,N_9526);
nand U10367 (N_10367,N_7554,N_7741);
nand U10368 (N_10368,N_9484,N_7552);
or U10369 (N_10369,N_8044,N_7592);
xnor U10370 (N_10370,N_9987,N_8131);
nor U10371 (N_10371,N_8929,N_8009);
and U10372 (N_10372,N_8001,N_7783);
nand U10373 (N_10373,N_8974,N_7971);
and U10374 (N_10374,N_8240,N_9398);
nand U10375 (N_10375,N_9504,N_9684);
nor U10376 (N_10376,N_9154,N_8328);
nor U10377 (N_10377,N_8873,N_8694);
nor U10378 (N_10378,N_8573,N_9663);
xnor U10379 (N_10379,N_8718,N_8816);
xnor U10380 (N_10380,N_8063,N_7634);
nand U10381 (N_10381,N_7526,N_8729);
and U10382 (N_10382,N_7802,N_7629);
nor U10383 (N_10383,N_8752,N_9929);
nor U10384 (N_10384,N_8109,N_8676);
nor U10385 (N_10385,N_9809,N_8806);
or U10386 (N_10386,N_9982,N_9029);
and U10387 (N_10387,N_9237,N_9651);
or U10388 (N_10388,N_9257,N_9369);
nor U10389 (N_10389,N_8756,N_9508);
or U10390 (N_10390,N_7842,N_9522);
nor U10391 (N_10391,N_8244,N_7892);
nor U10392 (N_10392,N_9701,N_8569);
nand U10393 (N_10393,N_8737,N_8035);
nand U10394 (N_10394,N_8124,N_8438);
and U10395 (N_10395,N_7931,N_9416);
or U10396 (N_10396,N_9986,N_9925);
and U10397 (N_10397,N_7872,N_8123);
and U10398 (N_10398,N_9454,N_9695);
nand U10399 (N_10399,N_8280,N_9828);
xor U10400 (N_10400,N_8241,N_8416);
and U10401 (N_10401,N_8854,N_8883);
xor U10402 (N_10402,N_9024,N_9090);
xor U10403 (N_10403,N_7797,N_8759);
xor U10404 (N_10404,N_7982,N_7757);
or U10405 (N_10405,N_9084,N_9448);
nand U10406 (N_10406,N_9236,N_8740);
and U10407 (N_10407,N_9453,N_8006);
xnor U10408 (N_10408,N_9952,N_9270);
nand U10409 (N_10409,N_8683,N_8958);
nor U10410 (N_10410,N_8414,N_8004);
nor U10411 (N_10411,N_9262,N_8469);
xor U10412 (N_10412,N_9307,N_8276);
xor U10413 (N_10413,N_8509,N_8309);
nor U10414 (N_10414,N_9983,N_9000);
or U10415 (N_10415,N_7831,N_9064);
and U10416 (N_10416,N_7558,N_9959);
nor U10417 (N_10417,N_9047,N_7963);
nor U10418 (N_10418,N_9775,N_9113);
nor U10419 (N_10419,N_8215,N_9505);
xnor U10420 (N_10420,N_7834,N_7561);
nand U10421 (N_10421,N_9370,N_8333);
nor U10422 (N_10422,N_9075,N_7694);
xor U10423 (N_10423,N_9988,N_9208);
or U10424 (N_10424,N_8319,N_8121);
xnor U10425 (N_10425,N_9793,N_8233);
or U10426 (N_10426,N_8366,N_9870);
and U10427 (N_10427,N_8791,N_9260);
nor U10428 (N_10428,N_9895,N_8499);
or U10429 (N_10429,N_8062,N_9143);
nand U10430 (N_10430,N_9440,N_9816);
and U10431 (N_10431,N_8984,N_9571);
and U10432 (N_10432,N_8945,N_9397);
or U10433 (N_10433,N_9104,N_7794);
nand U10434 (N_10434,N_8033,N_8028);
or U10435 (N_10435,N_8053,N_9726);
or U10436 (N_10436,N_9971,N_8140);
nor U10437 (N_10437,N_9153,N_8578);
xor U10438 (N_10438,N_8933,N_8613);
or U10439 (N_10439,N_9671,N_8867);
nor U10440 (N_10440,N_9033,N_7547);
and U10441 (N_10441,N_8106,N_9662);
xnor U10442 (N_10442,N_9602,N_9585);
xor U10443 (N_10443,N_7748,N_8435);
nand U10444 (N_10444,N_9382,N_9298);
and U10445 (N_10445,N_9502,N_9936);
and U10446 (N_10446,N_9105,N_9377);
or U10447 (N_10447,N_7740,N_9892);
nand U10448 (N_10448,N_9494,N_7605);
nor U10449 (N_10449,N_8163,N_8906);
xor U10450 (N_10450,N_8399,N_9960);
nor U10451 (N_10451,N_8977,N_8231);
or U10452 (N_10452,N_8624,N_8537);
and U10453 (N_10453,N_8915,N_7671);
and U10454 (N_10454,N_7765,N_8346);
and U10455 (N_10455,N_9794,N_9991);
or U10456 (N_10456,N_7920,N_8960);
nand U10457 (N_10457,N_8543,N_8790);
nor U10458 (N_10458,N_7637,N_9340);
xnor U10459 (N_10459,N_8576,N_7789);
and U10460 (N_10460,N_7723,N_8633);
xor U10461 (N_10461,N_8026,N_9475);
nor U10462 (N_10462,N_9650,N_7860);
nor U10463 (N_10463,N_7532,N_8812);
nor U10464 (N_10464,N_9486,N_9263);
xor U10465 (N_10465,N_9396,N_9512);
nor U10466 (N_10466,N_8839,N_8564);
or U10467 (N_10467,N_9948,N_8887);
nor U10468 (N_10468,N_9973,N_9672);
or U10469 (N_10469,N_8822,N_8426);
or U10470 (N_10470,N_9681,N_8550);
nand U10471 (N_10471,N_9391,N_8429);
nand U10472 (N_10472,N_9814,N_7790);
and U10473 (N_10473,N_8762,N_8808);
nand U10474 (N_10474,N_9689,N_9127);
xor U10475 (N_10475,N_8334,N_9832);
and U10476 (N_10476,N_8395,N_8965);
nor U10477 (N_10477,N_8880,N_9736);
nand U10478 (N_10478,N_7555,N_7918);
xnor U10479 (N_10479,N_9818,N_8890);
nor U10480 (N_10480,N_9088,N_8224);
nor U10481 (N_10481,N_9883,N_9461);
or U10482 (N_10482,N_7614,N_7635);
nor U10483 (N_10483,N_8248,N_8419);
nand U10484 (N_10484,N_8768,N_9834);
nor U10485 (N_10485,N_7693,N_7620);
nor U10486 (N_10486,N_8203,N_8152);
nand U10487 (N_10487,N_9057,N_9843);
nand U10488 (N_10488,N_8648,N_9329);
and U10489 (N_10489,N_7823,N_8619);
nor U10490 (N_10490,N_7673,N_9839);
xnor U10491 (N_10491,N_8735,N_7747);
nand U10492 (N_10492,N_9803,N_9060);
nor U10493 (N_10493,N_8381,N_8652);
and U10494 (N_10494,N_7861,N_8052);
or U10495 (N_10495,N_8243,N_8025);
nor U10496 (N_10496,N_8032,N_9155);
and U10497 (N_10497,N_9220,N_9066);
xor U10498 (N_10498,N_8896,N_9926);
nor U10499 (N_10499,N_8698,N_9364);
xor U10500 (N_10500,N_7653,N_9469);
nor U10501 (N_10501,N_8545,N_8038);
and U10502 (N_10502,N_8512,N_9680);
or U10503 (N_10503,N_7726,N_7776);
xnor U10504 (N_10504,N_9283,N_8423);
and U10505 (N_10505,N_8641,N_9733);
xor U10506 (N_10506,N_8234,N_9372);
nand U10507 (N_10507,N_9343,N_7937);
nand U10508 (N_10508,N_8194,N_9844);
xor U10509 (N_10509,N_7615,N_9253);
or U10510 (N_10510,N_8721,N_9810);
nor U10511 (N_10511,N_7816,N_9072);
nor U10512 (N_10512,N_7515,N_9482);
or U10513 (N_10513,N_8980,N_7980);
or U10514 (N_10514,N_9489,N_8878);
and U10515 (N_10515,N_8326,N_8841);
and U10516 (N_10516,N_8211,N_7984);
nand U10517 (N_10517,N_9493,N_8466);
nand U10518 (N_10518,N_9375,N_7713);
nor U10519 (N_10519,N_9579,N_9541);
nand U10520 (N_10520,N_9583,N_7737);
or U10521 (N_10521,N_8370,N_7700);
xor U10522 (N_10522,N_9157,N_8566);
xnor U10523 (N_10523,N_9517,N_7583);
and U10524 (N_10524,N_7856,N_9573);
or U10525 (N_10525,N_9062,N_8631);
nor U10526 (N_10526,N_9116,N_9908);
nor U10527 (N_10527,N_9038,N_7880);
and U10528 (N_10528,N_8722,N_7542);
nor U10529 (N_10529,N_7588,N_7786);
xnor U10530 (N_10530,N_8316,N_8519);
nand U10531 (N_10531,N_9399,N_8060);
and U10532 (N_10532,N_8421,N_8345);
nand U10533 (N_10533,N_8724,N_8102);
nor U10534 (N_10534,N_9100,N_8390);
or U10535 (N_10535,N_8646,N_7564);
xnor U10536 (N_10536,N_9193,N_8077);
xor U10537 (N_10537,N_8222,N_9985);
xor U10538 (N_10538,N_8487,N_8558);
and U10539 (N_10539,N_8711,N_8625);
and U10540 (N_10540,N_8027,N_9812);
xnor U10541 (N_10541,N_8712,N_7666);
nor U10542 (N_10542,N_9261,N_8596);
nor U10543 (N_10543,N_9568,N_7992);
nand U10544 (N_10544,N_8658,N_9647);
and U10545 (N_10545,N_8289,N_8115);
nand U10546 (N_10546,N_8155,N_9621);
and U10547 (N_10547,N_9352,N_8261);
and U10548 (N_10548,N_7559,N_9543);
and U10549 (N_10549,N_9012,N_9911);
nor U10550 (N_10550,N_9021,N_9400);
and U10551 (N_10551,N_8899,N_9906);
nand U10552 (N_10552,N_9640,N_9168);
and U10553 (N_10553,N_8245,N_9823);
nand U10554 (N_10554,N_9838,N_7969);
and U10555 (N_10555,N_7936,N_8869);
nand U10556 (N_10556,N_7698,N_9049);
nor U10557 (N_10557,N_7638,N_9857);
xnor U10558 (N_10558,N_7873,N_8017);
xnor U10559 (N_10559,N_8601,N_8180);
or U10560 (N_10560,N_7507,N_9566);
xor U10561 (N_10561,N_9964,N_7798);
or U10562 (N_10562,N_8073,N_8145);
or U10563 (N_10563,N_7822,N_7914);
and U10564 (N_10564,N_9666,N_7923);
and U10565 (N_10565,N_9646,N_7907);
nand U10566 (N_10566,N_9318,N_9001);
nand U10567 (N_10567,N_7651,N_9557);
xnor U10568 (N_10568,N_8008,N_7970);
or U10569 (N_10569,N_8055,N_9581);
xor U10570 (N_10570,N_8884,N_9710);
nor U10571 (N_10571,N_8640,N_7715);
nand U10572 (N_10572,N_8616,N_7562);
or U10573 (N_10573,N_7925,N_9313);
and U10574 (N_10574,N_7742,N_8600);
nor U10575 (N_10575,N_8278,N_8610);
xor U10576 (N_10576,N_8501,N_9893);
and U10577 (N_10577,N_9837,N_9850);
nand U10578 (N_10578,N_9575,N_8524);
and U10579 (N_10579,N_8817,N_7626);
or U10580 (N_10580,N_8523,N_8655);
nand U10581 (N_10581,N_8886,N_8374);
and U10582 (N_10582,N_8551,N_9519);
or U10583 (N_10583,N_7570,N_9949);
nor U10584 (N_10584,N_8263,N_8103);
xor U10585 (N_10585,N_8894,N_8723);
nand U10586 (N_10586,N_8069,N_7613);
or U10587 (N_10587,N_9528,N_9761);
and U10588 (N_10588,N_9750,N_9781);
or U10589 (N_10589,N_8981,N_7733);
and U10590 (N_10590,N_7942,N_8563);
nand U10591 (N_10591,N_7649,N_8749);
nor U10592 (N_10592,N_8483,N_8833);
xor U10593 (N_10593,N_9490,N_8455);
and U10594 (N_10594,N_8861,N_7766);
and U10595 (N_10595,N_7602,N_8467);
nand U10596 (N_10596,N_8608,N_8525);
and U10597 (N_10597,N_8559,N_9004);
nor U10598 (N_10598,N_7859,N_9082);
or U10599 (N_10599,N_9500,N_7815);
xor U10600 (N_10600,N_8473,N_8352);
nand U10601 (N_10601,N_8877,N_9586);
nor U10602 (N_10602,N_9159,N_9914);
xor U10603 (N_10603,N_8479,N_8587);
xnor U10604 (N_10604,N_7898,N_8581);
nand U10605 (N_10605,N_9617,N_9056);
xnor U10606 (N_10606,N_8056,N_7821);
or U10607 (N_10607,N_8113,N_9374);
or U10608 (N_10608,N_7539,N_9555);
xor U10609 (N_10609,N_8232,N_9273);
nor U10610 (N_10610,N_7510,N_9737);
nor U10611 (N_10611,N_9306,N_7782);
xor U10612 (N_10612,N_9599,N_9626);
or U10613 (N_10613,N_8836,N_8072);
and U10614 (N_10614,N_7594,N_9149);
nor U10615 (N_10615,N_8898,N_7624);
xor U10616 (N_10616,N_8491,N_7660);
nor U10617 (N_10617,N_8198,N_9552);
xor U10618 (N_10618,N_8657,N_8678);
xor U10619 (N_10619,N_8239,N_9408);
nor U10620 (N_10620,N_7894,N_9805);
xor U10621 (N_10621,N_7836,N_7622);
nand U10622 (N_10622,N_9709,N_8970);
nor U10623 (N_10623,N_8936,N_8710);
xnor U10624 (N_10624,N_9390,N_8407);
nor U10625 (N_10625,N_8287,N_9682);
nor U10626 (N_10626,N_9601,N_9770);
xor U10627 (N_10627,N_7639,N_7887);
xnor U10628 (N_10628,N_8947,N_7519);
nor U10629 (N_10629,N_8058,N_8852);
and U10630 (N_10630,N_8579,N_8259);
xnor U10631 (N_10631,N_9901,N_7650);
nand U10632 (N_10632,N_7878,N_9649);
or U10633 (N_10633,N_8134,N_8952);
xor U10634 (N_10634,N_9360,N_7938);
and U10635 (N_10635,N_9545,N_8262);
xnor U10636 (N_10636,N_8403,N_8088);
nand U10637 (N_10637,N_9854,N_8819);
nor U10638 (N_10638,N_7924,N_9462);
xnor U10639 (N_10639,N_9714,N_9604);
nand U10640 (N_10640,N_8389,N_7595);
nor U10641 (N_10641,N_8862,N_8465);
xnor U10642 (N_10642,N_8874,N_8148);
and U10643 (N_10643,N_9565,N_8630);
and U10644 (N_10644,N_7725,N_9381);
or U10645 (N_10645,N_7903,N_8191);
and U10646 (N_10646,N_9045,N_9401);
xnor U10647 (N_10647,N_9119,N_9301);
and U10648 (N_10648,N_8555,N_9063);
nor U10649 (N_10649,N_8442,N_9511);
nand U10650 (N_10650,N_7814,N_9798);
nor U10651 (N_10651,N_7688,N_9600);
xnor U10652 (N_10652,N_7784,N_9773);
and U10653 (N_10653,N_9860,N_9900);
or U10654 (N_10654,N_8607,N_9527);
xor U10655 (N_10655,N_7869,N_9206);
nand U10656 (N_10656,N_8653,N_7886);
nand U10657 (N_10657,N_8847,N_8925);
nor U10658 (N_10658,N_8994,N_9903);
or U10659 (N_10659,N_7685,N_8445);
xnor U10660 (N_10660,N_7840,N_8197);
and U10661 (N_10661,N_7647,N_9133);
and U10662 (N_10662,N_8317,N_7808);
and U10663 (N_10663,N_9654,N_9862);
nor U10664 (N_10664,N_9268,N_9932);
nand U10665 (N_10665,N_8335,N_7734);
nand U10666 (N_10666,N_8973,N_9189);
nand U10667 (N_10667,N_8179,N_9202);
nor U10668 (N_10668,N_9459,N_8951);
nand U10669 (N_10669,N_9849,N_8192);
nand U10670 (N_10670,N_8972,N_8458);
and U10671 (N_10671,N_7985,N_8150);
nor U10672 (N_10672,N_7645,N_9177);
or U10673 (N_10673,N_7670,N_7534);
nor U10674 (N_10674,N_7548,N_9898);
or U10675 (N_10675,N_7965,N_7568);
nor U10676 (N_10676,N_8932,N_9980);
or U10677 (N_10677,N_8717,N_9635);
xnor U10678 (N_10678,N_9706,N_8138);
and U10679 (N_10679,N_9629,N_9225);
or U10680 (N_10680,N_8380,N_9653);
or U10681 (N_10681,N_8700,N_9744);
xnor U10682 (N_10682,N_8303,N_8094);
nor U10683 (N_10683,N_9796,N_7557);
nor U10684 (N_10684,N_8743,N_8315);
nor U10685 (N_10685,N_9403,N_7727);
nor U10686 (N_10686,N_7935,N_7961);
or U10687 (N_10687,N_8725,N_8914);
and U10688 (N_10688,N_7904,N_9852);
xor U10689 (N_10689,N_9331,N_9956);
or U10690 (N_10690,N_8547,N_9099);
and U10691 (N_10691,N_8142,N_9151);
and U10692 (N_10692,N_8020,N_7704);
nand U10693 (N_10693,N_7659,N_8282);
or U10694 (N_10694,N_7843,N_9639);
nor U10695 (N_10695,N_8693,N_9134);
xnor U10696 (N_10696,N_9315,N_9842);
nor U10697 (N_10697,N_8837,N_9889);
nor U10698 (N_10698,N_8944,N_9282);
nor U10699 (N_10699,N_9836,N_8586);
nor U10700 (N_10700,N_9855,N_8195);
and U10701 (N_10701,N_7947,N_9248);
nor U10702 (N_10702,N_8343,N_7885);
and U10703 (N_10703,N_8450,N_8795);
or U10704 (N_10704,N_8975,N_7551);
xnor U10705 (N_10705,N_8692,N_8283);
xor U10706 (N_10706,N_8165,N_8650);
or U10707 (N_10707,N_8220,N_7939);
and U10708 (N_10708,N_8476,N_8522);
and U10709 (N_10709,N_8130,N_8695);
and U10710 (N_10710,N_9574,N_9218);
xnor U10711 (N_10711,N_7503,N_8760);
xor U10712 (N_10712,N_8014,N_9747);
nor U10713 (N_10713,N_9768,N_9632);
and U10714 (N_10714,N_8834,N_9554);
nor U10715 (N_10715,N_7565,N_9184);
and U10716 (N_10716,N_7560,N_9069);
nor U10717 (N_10717,N_8448,N_8341);
nor U10718 (N_10718,N_8418,N_9678);
nor U10719 (N_10719,N_8775,N_7710);
nor U10720 (N_10720,N_9128,N_7770);
or U10721 (N_10721,N_8093,N_8924);
xor U10722 (N_10722,N_9258,N_9840);
xnor U10723 (N_10723,N_9308,N_9738);
xor U10724 (N_10724,N_9356,N_9992);
or U10725 (N_10725,N_9174,N_8369);
or U10726 (N_10726,N_9608,N_8889);
and U10727 (N_10727,N_9040,N_7820);
or U10728 (N_10728,N_7731,N_9388);
or U10729 (N_10729,N_8500,N_8785);
or U10730 (N_10730,N_7959,N_9748);
nand U10731 (N_10731,N_8439,N_8149);
or U10732 (N_10732,N_9239,N_8482);
xnor U10733 (N_10733,N_8157,N_8029);
nor U10734 (N_10734,N_9071,N_7871);
nor U10735 (N_10735,N_9657,N_8813);
xor U10736 (N_10736,N_9841,N_9235);
nor U10737 (N_10737,N_9718,N_9226);
and U10738 (N_10738,N_9935,N_8217);
nand U10739 (N_10739,N_8595,N_9241);
or U10740 (N_10740,N_7874,N_9115);
nand U10741 (N_10741,N_9780,N_9873);
nand U10742 (N_10742,N_9182,N_7995);
nor U10743 (N_10743,N_7778,N_9821);
xnor U10744 (N_10744,N_8584,N_9358);
xor U10745 (N_10745,N_9869,N_9868);
or U10746 (N_10746,N_7579,N_7606);
or U10747 (N_10747,N_7701,N_9333);
and U10748 (N_10748,N_8227,N_9481);
nand U10749 (N_10749,N_8765,N_8668);
and U10750 (N_10750,N_8351,N_8497);
nand U10751 (N_10751,N_8802,N_7582);
or U10752 (N_10752,N_9008,N_9351);
nand U10753 (N_10753,N_7630,N_8190);
nand U10754 (N_10754,N_9132,N_8310);
xor U10755 (N_10755,N_9664,N_7876);
xnor U10756 (N_10756,N_8923,N_8057);
and U10757 (N_10757,N_9656,N_9668);
and U10758 (N_10758,N_7718,N_7932);
nor U10759 (N_10759,N_7736,N_8238);
and U10760 (N_10760,N_7636,N_9392);
nor U10761 (N_10761,N_8126,N_8446);
nand U10762 (N_10762,N_9290,N_8604);
or U10763 (N_10763,N_9335,N_8002);
nor U10764 (N_10764,N_8212,N_7913);
or U10765 (N_10765,N_9050,N_9293);
nor U10766 (N_10766,N_7988,N_8629);
nor U10767 (N_10767,N_8391,N_7593);
nor U10768 (N_10768,N_7844,N_8855);
or U10769 (N_10769,N_8651,N_9795);
xnor U10770 (N_10770,N_8260,N_8012);
xnor U10771 (N_10771,N_7689,N_9713);
or U10772 (N_10772,N_8939,N_9164);
or U10773 (N_10773,N_8373,N_9576);
nand U10774 (N_10774,N_8910,N_9279);
nor U10775 (N_10775,N_9658,N_9758);
nor U10776 (N_10776,N_8127,N_9087);
and U10777 (N_10777,N_8830,N_7721);
xnor U10778 (N_10778,N_8119,N_9578);
nor U10779 (N_10779,N_8935,N_9979);
nand U10780 (N_10780,N_8820,N_7976);
or U10781 (N_10781,N_7680,N_7960);
xnor U10782 (N_10782,N_9879,N_9614);
nor U10783 (N_10783,N_9802,N_8371);
or U10784 (N_10784,N_9443,N_8253);
and U10785 (N_10785,N_9872,N_9542);
xor U10786 (N_10786,N_8926,N_8562);
and U10787 (N_10787,N_9280,N_8081);
nor U10788 (N_10788,N_7901,N_8593);
xor U10789 (N_10789,N_7586,N_7848);
and U10790 (N_10790,N_8565,N_9323);
xor U10791 (N_10791,N_8475,N_9445);
and U10792 (N_10792,N_8378,N_9138);
nor U10793 (N_10793,N_8228,N_7571);
nand U10794 (N_10794,N_7772,N_8054);
nand U10795 (N_10795,N_8866,N_8848);
nor U10796 (N_10796,N_7709,N_7838);
nand U10797 (N_10797,N_9902,N_9819);
nor U10798 (N_10798,N_8097,N_8457);
and U10799 (N_10799,N_7870,N_8597);
and U10800 (N_10800,N_8000,N_8311);
or U10801 (N_10801,N_9299,N_9613);
and U10802 (N_10802,N_9238,N_9442);
and U10803 (N_10803,N_8304,N_8731);
nand U10804 (N_10804,N_8431,N_8571);
or U10805 (N_10805,N_8164,N_7654);
xor U10806 (N_10806,N_9232,N_8927);
and U10807 (N_10807,N_8413,N_9167);
or U10808 (N_10808,N_9827,N_8946);
nor U10809 (N_10809,N_9720,N_8049);
or U10810 (N_10810,N_8901,N_8118);
nand U10811 (N_10811,N_8349,N_9093);
or U10812 (N_10812,N_9321,N_9907);
xor U10813 (N_10813,N_9190,N_9173);
or U10814 (N_10814,N_8663,N_8185);
nand U10815 (N_10815,N_7891,N_9799);
or U10816 (N_10816,N_7993,N_8362);
xor U10817 (N_10817,N_8526,N_9622);
or U10818 (N_10818,N_9835,N_7911);
xor U10819 (N_10819,N_9641,N_9848);
nor U10820 (N_10820,N_8209,N_8154);
nor U10821 (N_10821,N_9139,N_7610);
or U10822 (N_10822,N_9227,N_9897);
nor U10823 (N_10823,N_9415,N_8247);
nor U10824 (N_10824,N_8982,N_8272);
xor U10825 (N_10825,N_9536,N_7525);
nand U10826 (N_10826,N_9271,N_9427);
nor U10827 (N_10827,N_7631,N_9961);
or U10828 (N_10828,N_9716,N_7703);
or U10829 (N_10829,N_8857,N_9102);
or U10830 (N_10830,N_8556,N_7852);
nand U10831 (N_10831,N_9199,N_8425);
nor U10832 (N_10832,N_9137,N_8246);
nor U10833 (N_10833,N_9297,N_9410);
and U10834 (N_10834,N_9013,N_9676);
or U10835 (N_10835,N_9114,N_8143);
or U10836 (N_10836,N_9851,N_8066);
nor U10837 (N_10837,N_9107,N_9880);
and U10838 (N_10838,N_7511,N_8954);
nand U10839 (N_10839,N_7746,N_8680);
and U10840 (N_10840,N_9930,N_9978);
xnor U10841 (N_10841,N_8210,N_8050);
nand U10842 (N_10842,N_9275,N_7964);
nand U10843 (N_10843,N_9195,N_9379);
and U10844 (N_10844,N_7877,N_8101);
nor U10845 (N_10845,N_8292,N_9589);
nor U10846 (N_10846,N_9550,N_8766);
and U10847 (N_10847,N_9068,N_9755);
and U10848 (N_10848,N_7773,N_8397);
or U10849 (N_10849,N_8461,N_8117);
xor U10850 (N_10850,N_7535,N_9492);
or U10851 (N_10851,N_8917,N_7676);
xor U10852 (N_10852,N_9539,N_7919);
or U10853 (N_10853,N_9231,N_8269);
xor U10854 (N_10854,N_9633,N_8086);
or U10855 (N_10855,N_9233,N_8367);
xor U10856 (N_10856,N_7826,N_8673);
xnor U10857 (N_10857,N_8726,N_7574);
xnor U10858 (N_10858,N_8213,N_8514);
nand U10859 (N_10859,N_9532,N_9745);
xor U10860 (N_10860,N_9373,N_8318);
xor U10861 (N_10861,N_8661,N_8202);
and U10862 (N_10862,N_8064,N_7504);
or U10863 (N_10863,N_9327,N_8405);
xnor U10864 (N_10864,N_8805,N_8850);
and U10865 (N_10865,N_7523,N_8909);
nand U10866 (N_10866,N_9624,N_8851);
and U10867 (N_10867,N_8331,N_9917);
and U10868 (N_10868,N_8827,N_9350);
and U10869 (N_10869,N_8572,N_8734);
xor U10870 (N_10870,N_8782,N_8071);
xnor U10871 (N_10871,N_8763,N_9124);
nor U10872 (N_10872,N_9634,N_8777);
or U10873 (N_10873,N_9743,N_8376);
or U10874 (N_10874,N_8821,N_7841);
nand U10875 (N_10875,N_9491,N_7966);
nand U10876 (N_10876,N_9939,N_9246);
xnor U10877 (N_10877,N_9894,N_8300);
nor U10878 (N_10878,N_7642,N_8411);
or U10879 (N_10879,N_7623,N_9205);
xor U10880 (N_10880,N_9707,N_9006);
or U10881 (N_10881,N_8295,N_9277);
nor U10882 (N_10882,N_7827,N_7735);
nor U10883 (N_10883,N_8490,N_8796);
nand U10884 (N_10884,N_9011,N_8781);
xnor U10885 (N_10885,N_8393,N_7819);
xor U10886 (N_10886,N_7730,N_9912);
nand U10887 (N_10887,N_9264,N_8893);
and U10888 (N_10888,N_7686,N_8301);
nor U10889 (N_10889,N_8575,N_9213);
nand U10890 (N_10890,N_9016,N_7916);
and U10891 (N_10891,N_7556,N_9789);
and U10892 (N_10892,N_9224,N_8427);
or U10893 (N_10893,N_9359,N_8338);
nand U10894 (N_10894,N_9065,N_7897);
or U10895 (N_10895,N_8332,N_9487);
and U10896 (N_10896,N_7929,N_9652);
or U10897 (N_10897,N_7754,N_8707);
nand U10898 (N_10898,N_7893,N_8907);
nor U10899 (N_10899,N_9590,N_8114);
and U10900 (N_10900,N_9175,N_9234);
or U10901 (N_10901,N_8911,N_9741);
nor U10902 (N_10902,N_9196,N_7501);
and U10903 (N_10903,N_9669,N_7973);
nor U10904 (N_10904,N_9464,N_9910);
nor U10905 (N_10905,N_9152,N_8686);
nand U10906 (N_10906,N_8542,N_8424);
nand U10907 (N_10907,N_9007,N_7955);
and U10908 (N_10908,N_9967,N_7909);
nor U10909 (N_10909,N_8736,N_9221);
or U10910 (N_10910,N_9387,N_9767);
xor U10911 (N_10911,N_8849,N_7744);
nor U10912 (N_10912,N_9027,N_7738);
or U10913 (N_10913,N_9194,N_8313);
nand U10914 (N_10914,N_9229,N_8881);
nand U10915 (N_10915,N_9086,N_8432);
nor U10916 (N_10916,N_8803,N_9010);
xnor U10917 (N_10917,N_8521,N_9161);
xor U10918 (N_10918,N_8356,N_8459);
xnor U10919 (N_10919,N_9688,N_8019);
nand U10920 (N_10920,N_9334,N_9256);
or U10921 (N_10921,N_9572,N_9674);
nand U10922 (N_10922,N_7905,N_9703);
nor U10923 (N_10923,N_8237,N_9070);
nand U10924 (N_10924,N_9922,N_9693);
or U10925 (N_10925,N_7751,N_9460);
or U10926 (N_10926,N_8428,N_9749);
nor U10927 (N_10927,N_9610,N_9786);
or U10928 (N_10928,N_8168,N_9171);
nor U10929 (N_10929,N_8083,N_9782);
xnor U10930 (N_10930,N_7563,N_9274);
or U10931 (N_10931,N_7600,N_9685);
nor U10932 (N_10932,N_8216,N_8080);
or U10933 (N_10933,N_8034,N_7661);
xor U10934 (N_10934,N_9302,N_8978);
xnor U10935 (N_10935,N_8360,N_8642);
or U10936 (N_10936,N_8679,N_9753);
nand U10937 (N_10937,N_7663,N_7573);
nand U10938 (N_10938,N_7883,N_7908);
nor U10939 (N_10939,N_8264,N_8644);
or U10940 (N_10940,N_9300,N_8685);
nor U10941 (N_10941,N_7682,N_7792);
or U10942 (N_10942,N_9759,N_8745);
and U10943 (N_10943,N_8536,N_9141);
nor U10944 (N_10944,N_9165,N_8727);
or U10945 (N_10945,N_7508,N_8636);
nor U10946 (N_10946,N_8036,N_9058);
and U10947 (N_10947,N_9790,N_9580);
nor U10948 (N_10948,N_9567,N_8903);
and U10949 (N_10949,N_9984,N_8159);
nor U10950 (N_10950,N_7825,N_9384);
or U10951 (N_10951,N_7800,N_7743);
and U10952 (N_10952,N_9905,N_7948);
or U10953 (N_10953,N_8410,N_9450);
or U10954 (N_10954,N_8664,N_9887);
or U10955 (N_10955,N_9135,N_8024);
or U10956 (N_10956,N_7795,N_7549);
or U10957 (N_10957,N_9243,N_9778);
xor U10958 (N_10958,N_8236,N_7780);
or U10959 (N_10959,N_9076,N_9899);
nor U10960 (N_10960,N_9537,N_8904);
xnor U10961 (N_10961,N_8515,N_9061);
and U10962 (N_10962,N_8460,N_8048);
xor U10963 (N_10963,N_7612,N_9250);
nand U10964 (N_10964,N_8895,N_9732);
nor U10965 (N_10965,N_9249,N_8535);
xor U10966 (N_10966,N_7665,N_9712);
and U10967 (N_10967,N_8527,N_9659);
or U10968 (N_10968,N_9455,N_8291);
nor U10969 (N_10969,N_8363,N_8971);
nor U10970 (N_10970,N_8870,N_9875);
xor U10971 (N_10971,N_9067,N_8051);
and U10972 (N_10972,N_7933,N_9363);
nand U10973 (N_10973,N_7553,N_8900);
or U10974 (N_10974,N_8251,N_8225);
and U10975 (N_10975,N_9465,N_7774);
xnor U10976 (N_10976,N_7910,N_7796);
nor U10977 (N_10977,N_7779,N_8219);
nand U10978 (N_10978,N_7853,N_8186);
or U10979 (N_10979,N_9251,N_9295);
or U10980 (N_10980,N_9764,N_8277);
and U10981 (N_10981,N_8594,N_8913);
nand U10982 (N_10982,N_8865,N_7509);
nand U10983 (N_10983,N_9211,N_8451);
nand U10984 (N_10984,N_9429,N_8557);
or U10985 (N_10985,N_9520,N_9210);
and U10986 (N_10986,N_9538,N_9721);
xor U10987 (N_10987,N_8175,N_8744);
nor U10988 (N_10988,N_8342,N_9970);
nor U10989 (N_10989,N_9483,N_8875);
xor U10990 (N_10990,N_9316,N_8327);
or U10991 (N_10991,N_8538,N_8533);
xnor U10992 (N_10992,N_8047,N_8738);
or U10993 (N_10993,N_8843,N_8546);
nor U10994 (N_10994,N_8513,N_7952);
and U10995 (N_10995,N_9943,N_7707);
nor U10996 (N_10996,N_7750,N_7537);
xnor U10997 (N_10997,N_7589,N_9615);
nor U10998 (N_10998,N_9146,N_7633);
xor U10999 (N_10999,N_8447,N_9820);
xor U11000 (N_11000,N_9938,N_7835);
nand U11001 (N_11001,N_7917,N_7962);
xor U11002 (N_11002,N_9603,N_8498);
or U11003 (N_11003,N_8357,N_9346);
nor U11004 (N_11004,N_9496,N_8516);
xor U11005 (N_11005,N_8485,N_7998);
and U11006 (N_11006,N_9110,N_9815);
nor U11007 (N_11007,N_8966,N_8039);
nand U11008 (N_11008,N_7550,N_7791);
and U11009 (N_11009,N_7597,N_8330);
or U11010 (N_11010,N_7830,N_7769);
nand U11011 (N_11011,N_9757,N_8950);
nand U11012 (N_11012,N_8404,N_8949);
and U11013 (N_11013,N_7847,N_7958);
xnor U11014 (N_11014,N_9041,N_8691);
nand U11015 (N_11015,N_9947,N_8628);
xor U11016 (N_11016,N_8305,N_8256);
nand U11017 (N_11017,N_8045,N_9885);
xnor U11018 (N_11018,N_8675,N_9771);
nor U11019 (N_11019,N_8828,N_8128);
nor U11020 (N_11020,N_9856,N_8415);
or U11021 (N_11021,N_9866,N_8798);
and U11022 (N_11022,N_9354,N_9095);
xor U11023 (N_11023,N_9053,N_8468);
nand U11024 (N_11024,N_8386,N_9365);
and U11025 (N_11025,N_8258,N_8784);
and U11026 (N_11026,N_9426,N_7641);
nor U11027 (N_11027,N_8372,N_8188);
nand U11028 (N_11028,N_9353,N_7915);
or U11029 (N_11029,N_7879,N_9913);
xnor U11030 (N_11030,N_7655,N_8484);
nor U11031 (N_11031,N_9697,N_8532);
or U11032 (N_11032,N_8778,N_8770);
xor U11033 (N_11033,N_7732,N_8354);
nand U11034 (N_11034,N_8799,N_9966);
xor U11035 (N_11035,N_8167,N_9436);
or U11036 (N_11036,N_8299,N_8462);
or U11037 (N_11037,N_8443,N_8504);
and U11038 (N_11038,N_9291,N_9754);
xor U11039 (N_11039,N_9933,N_7505);
xor U11040 (N_11040,N_8934,N_7865);
nand U11041 (N_11041,N_9457,N_7753);
nor U11042 (N_11042,N_9944,N_9549);
xnor U11043 (N_11043,N_9439,N_8141);
or U11044 (N_11044,N_8585,N_7596);
or U11045 (N_11045,N_8696,N_8312);
nand U11046 (N_11046,N_9735,N_9476);
and U11047 (N_11047,N_9660,N_9118);
nand U11048 (N_11048,N_7577,N_9367);
xor U11049 (N_11049,N_9207,N_9419);
xor U11050 (N_11050,N_8452,N_7607);
and U11051 (N_11051,N_9120,N_8750);
nor U11052 (N_11052,N_8771,N_7566);
and U11053 (N_11053,N_8992,N_9406);
or U11054 (N_11054,N_8611,N_9272);
nand U11055 (N_11055,N_9801,N_9304);
or U11056 (N_11056,N_7944,N_8046);
nand U11057 (N_11057,N_8472,N_7990);
xnor U11058 (N_11058,N_8800,N_9317);
nand U11059 (N_11059,N_7813,N_9456);
nand U11060 (N_11060,N_7803,N_7839);
or U11061 (N_11061,N_9628,N_9428);
nand U11062 (N_11062,N_9945,N_9197);
xor U11063 (N_11063,N_8969,N_9919);
or U11064 (N_11064,N_7684,N_8493);
nand U11065 (N_11065,N_9940,N_9294);
xor U11066 (N_11066,N_8659,N_9995);
nor U11067 (N_11067,N_9344,N_7761);
nor U11068 (N_11068,N_9594,N_7677);
and U11069 (N_11069,N_9163,N_7720);
nand U11070 (N_11070,N_8746,N_8365);
xnor U11071 (N_11071,N_8976,N_9101);
nand U11072 (N_11072,N_9612,N_8003);
xor U11073 (N_11073,N_9616,N_9362);
and U11074 (N_11074,N_7584,N_8120);
and U11075 (N_11075,N_7603,N_9035);
nand U11076 (N_11076,N_7829,N_8741);
and U11077 (N_11077,N_8541,N_9564);
xor U11078 (N_11078,N_9215,N_9216);
and U11079 (N_11079,N_9191,N_8385);
xnor U11080 (N_11080,N_8518,N_7572);
nand U11081 (N_11081,N_7828,N_8826);
and U11082 (N_11082,N_9605,N_7667);
or U11083 (N_11083,N_9763,N_9928);
nor U11084 (N_11084,N_9278,N_9310);
or U11085 (N_11085,N_8184,N_7934);
and U11086 (N_11086,N_7749,N_9642);
nor U11087 (N_11087,N_9636,N_8920);
xor U11088 (N_11088,N_9534,N_8273);
nor U11089 (N_11089,N_9999,N_9515);
xor U11090 (N_11090,N_9811,N_7714);
or U11091 (N_11091,N_9192,N_8842);
xor U11092 (N_11092,N_8957,N_9326);
nand U11093 (N_11093,N_9147,N_7697);
xor U11094 (N_11094,N_8719,N_9696);
nor U11095 (N_11095,N_7810,N_7591);
and U11096 (N_11096,N_8665,N_9529);
xor U11097 (N_11097,N_9339,N_7867);
nand U11098 (N_11098,N_8353,N_7632);
and U11099 (N_11099,N_8931,N_9136);
and U11100 (N_11100,N_8733,N_8135);
nor U11101 (N_11101,N_8384,N_9853);
nor U11102 (N_11102,N_9797,N_9643);
and U11103 (N_11103,N_7785,N_8087);
and U11104 (N_11104,N_8173,N_7946);
nor U11105 (N_11105,N_9014,N_9265);
nand U11106 (N_11106,N_9556,N_8099);
nor U11107 (N_11107,N_7832,N_8928);
nor U11108 (N_11108,N_8189,N_8392);
xnor U11109 (N_11109,N_9287,N_9451);
and U11110 (N_11110,N_9831,N_9079);
xnor U11111 (N_11111,N_9444,N_9404);
nand U11112 (N_11112,N_9437,N_8879);
and U11113 (N_11113,N_9172,N_9865);
nand U11114 (N_11114,N_9704,N_7533);
or U11115 (N_11115,N_9463,N_8308);
and U11116 (N_11116,N_8892,N_9083);
or U11117 (N_11117,N_9296,N_8742);
xor U11118 (N_11118,N_9414,N_8614);
nand U11119 (N_11119,N_7890,N_8713);
and U11120 (N_11120,N_8786,N_8398);
or U11121 (N_11121,N_7656,N_7575);
or U11122 (N_11122,N_9507,N_9281);
and U11123 (N_11123,N_7974,N_7855);
and U11124 (N_11124,N_8956,N_8788);
xnor U11125 (N_11125,N_9449,N_8268);
nor U11126 (N_11126,N_9551,N_8639);
or U11127 (N_11127,N_9080,N_7541);
and U11128 (N_11128,N_8930,N_7881);
and U11129 (N_11129,N_9740,N_7809);
or U11130 (N_11130,N_9178,N_8574);
xor U11131 (N_11131,N_7658,N_8070);
or U11132 (N_11132,N_9276,N_8617);
nand U11133 (N_11133,N_8751,N_9421);
and U11134 (N_11134,N_8995,N_8689);
nand U11135 (N_11135,N_9923,N_7956);
xor U11136 (N_11136,N_9920,N_8845);
and U11137 (N_11137,N_9015,N_8091);
xor U11138 (N_11138,N_8076,N_8714);
or U11139 (N_11139,N_9514,N_8396);
nor U11140 (N_11140,N_8478,N_8764);
nand U11141 (N_11141,N_9292,N_7921);
xor U11142 (N_11142,N_9180,N_9023);
and U11143 (N_11143,N_8690,N_7529);
xnor U11144 (N_11144,N_9255,N_7621);
and U11145 (N_11145,N_8916,N_9467);
nor U11146 (N_11146,N_8488,N_7787);
or U11147 (N_11147,N_7545,N_8918);
nor U11148 (N_11148,N_7997,N_9896);
and U11149 (N_11149,N_9252,N_8108);
and U11150 (N_11150,N_9699,N_7699);
nor U11151 (N_11151,N_8153,N_8089);
xor U11152 (N_11152,N_9183,N_9020);
or U11153 (N_11153,N_8669,N_8031);
xnor U11154 (N_11154,N_9319,N_8872);
xor U11155 (N_11155,N_8095,N_8891);
and U11156 (N_11156,N_9156,N_7817);
xnor U11157 (N_11157,N_8325,N_7500);
nand U11158 (N_11158,N_8409,N_8441);
xor U11159 (N_11159,N_9466,N_8281);
nor U11160 (N_11160,N_7513,N_9332);
nand U11161 (N_11161,N_8592,N_9357);
nor U11162 (N_11162,N_8284,N_9441);
or U11163 (N_11163,N_9003,N_8078);
nor U11164 (N_11164,N_9942,N_8780);
and U11165 (N_11165,N_9598,N_8948);
xor U11166 (N_11166,N_8275,N_8348);
xnor U11167 (N_11167,N_9148,N_7949);
or U11168 (N_11168,N_8748,N_7851);
or U11169 (N_11169,N_9510,N_9129);
xnor U11170 (N_11170,N_8761,N_7618);
nand U11171 (N_11171,N_8162,N_9661);
nor U11172 (N_11172,N_7546,N_8505);
nor U11173 (N_11173,N_8704,N_8825);
nor U11174 (N_11174,N_9975,N_9103);
or U11175 (N_11175,N_9784,N_7895);
nand U11176 (N_11176,N_7863,N_9779);
nor U11177 (N_11177,N_8667,N_9412);
nand U11178 (N_11178,N_7941,N_9884);
or U11179 (N_11179,N_9176,N_7619);
and U11180 (N_11180,N_8990,N_9560);
or U11181 (N_11181,N_8147,N_8267);
xor U11182 (N_11182,N_8905,N_7681);
and U11183 (N_11183,N_8408,N_9209);
nand U11184 (N_11184,N_8643,N_7902);
or U11185 (N_11185,N_7706,N_9245);
nand U11186 (N_11186,N_9645,N_8552);
nor U11187 (N_11187,N_9037,N_8672);
or U11188 (N_11188,N_8296,N_7975);
and U11189 (N_11189,N_8840,N_7512);
nand U11190 (N_11190,N_8137,N_9776);
nor U11191 (N_11191,N_9756,N_8758);
nor U11192 (N_11192,N_7922,N_8660);
or U11193 (N_11193,N_9059,N_8116);
nor U11194 (N_11194,N_8885,N_8955);
nand U11195 (N_11195,N_7585,N_9303);
and U11196 (N_11196,N_8612,N_7643);
nand U11197 (N_11197,N_8637,N_9030);
and U11198 (N_11198,N_7679,N_9073);
nand U11199 (N_11199,N_8151,N_9769);
or U11200 (N_11200,N_9506,N_9314);
nor U11201 (N_11201,N_7977,N_9112);
nand U11202 (N_11202,N_8377,N_7604);
or U11203 (N_11203,N_9420,N_8531);
nand U11204 (N_11204,N_9034,N_8603);
or U11205 (N_11205,N_7793,N_8112);
nand U11206 (N_11206,N_7804,N_8702);
xnor U11207 (N_11207,N_8023,N_8196);
xor U11208 (N_11208,N_8337,N_9553);
nand U11209 (N_11209,N_7994,N_8030);
nand U11210 (N_11210,N_9996,N_9807);
and U11211 (N_11211,N_7520,N_8638);
or U11212 (N_11212,N_7818,N_8075);
and U11213 (N_11213,N_8290,N_7724);
xnor U11214 (N_11214,N_9958,N_8985);
xnor U11215 (N_11215,N_7983,N_9376);
xnor U11216 (N_11216,N_8477,N_8988);
and U11217 (N_11217,N_8561,N_9305);
nand U11218 (N_11218,N_7866,N_9043);
nand U11219 (N_11219,N_9516,N_8208);
and U11220 (N_11220,N_9434,N_8387);
or U11221 (N_11221,N_9019,N_9777);
nor U11222 (N_11222,N_7517,N_7957);
and U11223 (N_11223,N_7989,N_9338);
nor U11224 (N_11224,N_8767,N_8007);
and U11225 (N_11225,N_9774,N_9284);
and U11226 (N_11226,N_9667,N_8996);
xor U11227 (N_11227,N_8797,N_9431);
xnor U11228 (N_11228,N_9380,N_7578);
and U11229 (N_11229,N_8627,N_7906);
or U11230 (N_11230,N_9931,N_9859);
nand U11231 (N_11231,N_8288,N_9371);
xor U11232 (N_11232,N_9285,N_9723);
and U11233 (N_11233,N_8649,N_9808);
xor U11234 (N_11234,N_8709,N_8067);
xnor U11235 (N_11235,N_8888,N_8144);
nor U11236 (N_11236,N_9921,N_9026);
xnor U11237 (N_11237,N_8703,N_7884);
nor U11238 (N_11238,N_8831,N_9267);
or U11239 (N_11239,N_8615,N_8171);
nor U11240 (N_11240,N_7775,N_9228);
nor U11241 (N_11241,N_9535,N_9031);
and U11242 (N_11242,N_7943,N_7527);
nor U11243 (N_11243,N_7928,N_7662);
xor U11244 (N_11244,N_8214,N_9509);
nor U11245 (N_11245,N_9513,N_8226);
xor U11246 (N_11246,N_9142,N_9407);
nor U11247 (N_11247,N_9595,N_9077);
nor U11248 (N_11248,N_9909,N_9637);
xor U11249 (N_11249,N_7536,N_8379);
nand U11250 (N_11250,N_9538,N_8534);
xnor U11251 (N_11251,N_7762,N_9437);
nor U11252 (N_11252,N_8061,N_8022);
xnor U11253 (N_11253,N_7587,N_8392);
xnor U11254 (N_11254,N_9155,N_8235);
xnor U11255 (N_11255,N_8894,N_8439);
nand U11256 (N_11256,N_8294,N_7652);
and U11257 (N_11257,N_8585,N_8102);
xor U11258 (N_11258,N_8917,N_8572);
or U11259 (N_11259,N_8763,N_8821);
nor U11260 (N_11260,N_8999,N_8807);
nor U11261 (N_11261,N_8345,N_8318);
xnor U11262 (N_11262,N_8724,N_8591);
and U11263 (N_11263,N_8441,N_9130);
and U11264 (N_11264,N_8504,N_9712);
nor U11265 (N_11265,N_7889,N_8135);
and U11266 (N_11266,N_9744,N_9668);
xor U11267 (N_11267,N_7894,N_7658);
or U11268 (N_11268,N_8860,N_7839);
and U11269 (N_11269,N_9525,N_7627);
xnor U11270 (N_11270,N_8084,N_9076);
and U11271 (N_11271,N_8027,N_9926);
nor U11272 (N_11272,N_9721,N_9924);
nor U11273 (N_11273,N_7951,N_9603);
and U11274 (N_11274,N_7997,N_8861);
and U11275 (N_11275,N_8942,N_8872);
xor U11276 (N_11276,N_7871,N_8599);
and U11277 (N_11277,N_7711,N_9927);
xnor U11278 (N_11278,N_9735,N_9267);
and U11279 (N_11279,N_7863,N_9367);
nor U11280 (N_11280,N_9145,N_9339);
xnor U11281 (N_11281,N_8195,N_7593);
and U11282 (N_11282,N_8598,N_8381);
or U11283 (N_11283,N_8165,N_8568);
nand U11284 (N_11284,N_7724,N_7527);
nand U11285 (N_11285,N_8821,N_9834);
xor U11286 (N_11286,N_8694,N_9653);
nand U11287 (N_11287,N_8873,N_9608);
nor U11288 (N_11288,N_9107,N_8501);
and U11289 (N_11289,N_9559,N_8689);
nor U11290 (N_11290,N_8189,N_8238);
xnor U11291 (N_11291,N_8613,N_8753);
and U11292 (N_11292,N_8937,N_7878);
nor U11293 (N_11293,N_9454,N_7875);
and U11294 (N_11294,N_9465,N_8069);
xnor U11295 (N_11295,N_7623,N_8085);
or U11296 (N_11296,N_8724,N_9180);
nor U11297 (N_11297,N_7580,N_7714);
nor U11298 (N_11298,N_9259,N_9981);
or U11299 (N_11299,N_8413,N_7829);
xnor U11300 (N_11300,N_8011,N_7622);
and U11301 (N_11301,N_8950,N_9315);
nor U11302 (N_11302,N_8917,N_8333);
nor U11303 (N_11303,N_8088,N_9993);
nor U11304 (N_11304,N_8616,N_7545);
or U11305 (N_11305,N_9773,N_8462);
nand U11306 (N_11306,N_8284,N_9570);
xor U11307 (N_11307,N_7849,N_7759);
nand U11308 (N_11308,N_8311,N_8305);
nand U11309 (N_11309,N_9131,N_7884);
nand U11310 (N_11310,N_8295,N_7697);
and U11311 (N_11311,N_8333,N_7765);
nor U11312 (N_11312,N_7543,N_9137);
nor U11313 (N_11313,N_7792,N_7921);
xnor U11314 (N_11314,N_8192,N_7822);
or U11315 (N_11315,N_8538,N_8623);
nor U11316 (N_11316,N_9460,N_9271);
or U11317 (N_11317,N_9968,N_9636);
or U11318 (N_11318,N_8452,N_8137);
nand U11319 (N_11319,N_9193,N_9696);
nor U11320 (N_11320,N_8154,N_9693);
or U11321 (N_11321,N_7577,N_7780);
nand U11322 (N_11322,N_8942,N_8519);
nand U11323 (N_11323,N_8667,N_8305);
nor U11324 (N_11324,N_8193,N_9431);
xor U11325 (N_11325,N_9291,N_8191);
or U11326 (N_11326,N_8999,N_7767);
or U11327 (N_11327,N_7745,N_9432);
nand U11328 (N_11328,N_9502,N_9334);
nand U11329 (N_11329,N_8239,N_8437);
or U11330 (N_11330,N_8839,N_7870);
nor U11331 (N_11331,N_9288,N_9863);
or U11332 (N_11332,N_8888,N_9269);
or U11333 (N_11333,N_8629,N_8847);
nor U11334 (N_11334,N_9161,N_8659);
nor U11335 (N_11335,N_9622,N_9035);
nor U11336 (N_11336,N_8516,N_8057);
and U11337 (N_11337,N_7650,N_8051);
xnor U11338 (N_11338,N_9357,N_8402);
or U11339 (N_11339,N_8179,N_9622);
or U11340 (N_11340,N_7653,N_7750);
or U11341 (N_11341,N_9321,N_9828);
nor U11342 (N_11342,N_9817,N_9261);
nand U11343 (N_11343,N_9862,N_9885);
nor U11344 (N_11344,N_7589,N_7633);
or U11345 (N_11345,N_8338,N_9819);
nand U11346 (N_11346,N_7812,N_7773);
and U11347 (N_11347,N_8842,N_9707);
or U11348 (N_11348,N_7933,N_8036);
nor U11349 (N_11349,N_7563,N_9046);
and U11350 (N_11350,N_9534,N_8960);
or U11351 (N_11351,N_7895,N_8712);
xor U11352 (N_11352,N_7778,N_8244);
nand U11353 (N_11353,N_8527,N_9963);
xor U11354 (N_11354,N_9759,N_9752);
or U11355 (N_11355,N_7712,N_9038);
nand U11356 (N_11356,N_8030,N_8078);
nor U11357 (N_11357,N_7575,N_7674);
nor U11358 (N_11358,N_9009,N_9429);
and U11359 (N_11359,N_9590,N_8380);
or U11360 (N_11360,N_7572,N_8428);
or U11361 (N_11361,N_8828,N_9653);
nand U11362 (N_11362,N_7927,N_7998);
or U11363 (N_11363,N_8786,N_9966);
or U11364 (N_11364,N_8904,N_9254);
or U11365 (N_11365,N_9180,N_8585);
or U11366 (N_11366,N_8301,N_9366);
or U11367 (N_11367,N_8656,N_9946);
or U11368 (N_11368,N_7991,N_8370);
nand U11369 (N_11369,N_9500,N_9754);
and U11370 (N_11370,N_9407,N_9538);
or U11371 (N_11371,N_8134,N_9197);
xor U11372 (N_11372,N_8539,N_7865);
nand U11373 (N_11373,N_9788,N_9118);
and U11374 (N_11374,N_8391,N_9758);
and U11375 (N_11375,N_9307,N_9661);
nor U11376 (N_11376,N_9685,N_7636);
nand U11377 (N_11377,N_8585,N_8148);
and U11378 (N_11378,N_7534,N_8133);
or U11379 (N_11379,N_9373,N_8368);
xnor U11380 (N_11380,N_9603,N_8886);
or U11381 (N_11381,N_7538,N_8313);
and U11382 (N_11382,N_8185,N_7848);
nand U11383 (N_11383,N_7959,N_8756);
or U11384 (N_11384,N_8179,N_8184);
or U11385 (N_11385,N_9837,N_8529);
nand U11386 (N_11386,N_7549,N_8345);
xor U11387 (N_11387,N_9745,N_8978);
xor U11388 (N_11388,N_8531,N_8267);
nand U11389 (N_11389,N_8234,N_8170);
or U11390 (N_11390,N_9038,N_9258);
or U11391 (N_11391,N_8033,N_9616);
nand U11392 (N_11392,N_7731,N_9940);
nor U11393 (N_11393,N_8743,N_7649);
or U11394 (N_11394,N_8811,N_9436);
and U11395 (N_11395,N_7951,N_9759);
xnor U11396 (N_11396,N_8490,N_9837);
or U11397 (N_11397,N_9236,N_8499);
xnor U11398 (N_11398,N_7804,N_9946);
xor U11399 (N_11399,N_8454,N_9206);
xnor U11400 (N_11400,N_7657,N_9170);
and U11401 (N_11401,N_7877,N_9354);
and U11402 (N_11402,N_8004,N_9960);
nor U11403 (N_11403,N_9313,N_9042);
nor U11404 (N_11404,N_9342,N_8413);
or U11405 (N_11405,N_9081,N_9834);
or U11406 (N_11406,N_8210,N_9806);
or U11407 (N_11407,N_8183,N_7641);
or U11408 (N_11408,N_8907,N_8856);
and U11409 (N_11409,N_8748,N_9509);
xnor U11410 (N_11410,N_8210,N_9037);
or U11411 (N_11411,N_8431,N_8959);
or U11412 (N_11412,N_8219,N_8986);
nor U11413 (N_11413,N_9111,N_9545);
or U11414 (N_11414,N_9298,N_8070);
nand U11415 (N_11415,N_9258,N_8478);
and U11416 (N_11416,N_9764,N_8532);
nand U11417 (N_11417,N_8580,N_9234);
nand U11418 (N_11418,N_7520,N_8903);
or U11419 (N_11419,N_9674,N_7632);
nor U11420 (N_11420,N_7987,N_9944);
and U11421 (N_11421,N_7750,N_7639);
xnor U11422 (N_11422,N_8708,N_8958);
or U11423 (N_11423,N_7982,N_7687);
nand U11424 (N_11424,N_8646,N_9908);
nand U11425 (N_11425,N_8230,N_7592);
xnor U11426 (N_11426,N_7750,N_7640);
nand U11427 (N_11427,N_7749,N_8391);
and U11428 (N_11428,N_8693,N_8986);
and U11429 (N_11429,N_8412,N_9377);
and U11430 (N_11430,N_8618,N_9234);
nand U11431 (N_11431,N_9064,N_9898);
nor U11432 (N_11432,N_9161,N_7704);
and U11433 (N_11433,N_8998,N_7574);
nor U11434 (N_11434,N_7924,N_9790);
nor U11435 (N_11435,N_9686,N_8333);
nor U11436 (N_11436,N_8658,N_7904);
xor U11437 (N_11437,N_8009,N_8319);
nand U11438 (N_11438,N_9940,N_9801);
or U11439 (N_11439,N_8628,N_8633);
xnor U11440 (N_11440,N_9300,N_7665);
nor U11441 (N_11441,N_9997,N_8044);
nor U11442 (N_11442,N_9729,N_9934);
and U11443 (N_11443,N_8482,N_7772);
nand U11444 (N_11444,N_8347,N_9825);
xor U11445 (N_11445,N_9034,N_9183);
or U11446 (N_11446,N_7808,N_7753);
and U11447 (N_11447,N_9641,N_9532);
nand U11448 (N_11448,N_7502,N_7990);
nor U11449 (N_11449,N_9320,N_8716);
xnor U11450 (N_11450,N_7927,N_9433);
xor U11451 (N_11451,N_8153,N_9156);
or U11452 (N_11452,N_8569,N_9233);
nor U11453 (N_11453,N_7923,N_7628);
nor U11454 (N_11454,N_9065,N_8159);
nor U11455 (N_11455,N_9964,N_9833);
nand U11456 (N_11456,N_9028,N_7774);
and U11457 (N_11457,N_8691,N_9357);
and U11458 (N_11458,N_8726,N_9035);
or U11459 (N_11459,N_8179,N_9979);
nand U11460 (N_11460,N_7817,N_7578);
or U11461 (N_11461,N_7713,N_8685);
or U11462 (N_11462,N_9703,N_9175);
xor U11463 (N_11463,N_9096,N_9037);
nand U11464 (N_11464,N_9738,N_8434);
nand U11465 (N_11465,N_8972,N_7977);
and U11466 (N_11466,N_9497,N_7619);
or U11467 (N_11467,N_9731,N_8313);
xnor U11468 (N_11468,N_9314,N_9643);
nand U11469 (N_11469,N_9842,N_8012);
nand U11470 (N_11470,N_8841,N_8221);
or U11471 (N_11471,N_8478,N_9862);
nor U11472 (N_11472,N_9390,N_9324);
and U11473 (N_11473,N_8594,N_8345);
or U11474 (N_11474,N_8644,N_9506);
xor U11475 (N_11475,N_9261,N_9026);
nand U11476 (N_11476,N_7884,N_9695);
and U11477 (N_11477,N_9675,N_7877);
or U11478 (N_11478,N_8866,N_9124);
and U11479 (N_11479,N_8224,N_9644);
xnor U11480 (N_11480,N_8524,N_8265);
or U11481 (N_11481,N_7731,N_8796);
nand U11482 (N_11482,N_7954,N_9598);
or U11483 (N_11483,N_9851,N_9677);
and U11484 (N_11484,N_7648,N_9245);
nand U11485 (N_11485,N_9990,N_9016);
and U11486 (N_11486,N_8981,N_8441);
or U11487 (N_11487,N_7965,N_9807);
xor U11488 (N_11488,N_8618,N_9046);
nand U11489 (N_11489,N_9650,N_7854);
or U11490 (N_11490,N_9130,N_9186);
nor U11491 (N_11491,N_7606,N_9292);
nor U11492 (N_11492,N_9974,N_7533);
nor U11493 (N_11493,N_8931,N_7964);
xnor U11494 (N_11494,N_8555,N_7835);
xnor U11495 (N_11495,N_9647,N_9972);
nor U11496 (N_11496,N_8343,N_7793);
nor U11497 (N_11497,N_9467,N_8637);
xnor U11498 (N_11498,N_8144,N_7687);
and U11499 (N_11499,N_9831,N_8927);
nand U11500 (N_11500,N_8958,N_7832);
and U11501 (N_11501,N_8880,N_8048);
nand U11502 (N_11502,N_8384,N_9517);
or U11503 (N_11503,N_8927,N_8954);
xor U11504 (N_11504,N_8491,N_9228);
nor U11505 (N_11505,N_9112,N_8377);
and U11506 (N_11506,N_7911,N_9269);
nor U11507 (N_11507,N_9662,N_9844);
xor U11508 (N_11508,N_7716,N_9567);
or U11509 (N_11509,N_9783,N_8924);
nor U11510 (N_11510,N_8278,N_9111);
nand U11511 (N_11511,N_8073,N_8277);
nand U11512 (N_11512,N_9701,N_7794);
or U11513 (N_11513,N_8425,N_8820);
nand U11514 (N_11514,N_7851,N_9774);
nand U11515 (N_11515,N_9444,N_8641);
xnor U11516 (N_11516,N_9874,N_9309);
xnor U11517 (N_11517,N_9318,N_9968);
xnor U11518 (N_11518,N_9019,N_7670);
and U11519 (N_11519,N_8530,N_9348);
nand U11520 (N_11520,N_8889,N_7962);
xnor U11521 (N_11521,N_9717,N_7918);
nor U11522 (N_11522,N_8602,N_7915);
nor U11523 (N_11523,N_9052,N_9022);
xnor U11524 (N_11524,N_9681,N_9030);
and U11525 (N_11525,N_8443,N_8011);
nor U11526 (N_11526,N_7692,N_9682);
and U11527 (N_11527,N_8870,N_9495);
nor U11528 (N_11528,N_8359,N_9819);
xnor U11529 (N_11529,N_8699,N_9282);
or U11530 (N_11530,N_8227,N_9359);
nor U11531 (N_11531,N_7510,N_8999);
and U11532 (N_11532,N_7696,N_7939);
nor U11533 (N_11533,N_8905,N_7518);
xor U11534 (N_11534,N_8834,N_9269);
nand U11535 (N_11535,N_8273,N_9473);
nor U11536 (N_11536,N_8157,N_9479);
nor U11537 (N_11537,N_9984,N_8631);
xnor U11538 (N_11538,N_8368,N_9680);
xor U11539 (N_11539,N_9963,N_9238);
xnor U11540 (N_11540,N_9509,N_7637);
or U11541 (N_11541,N_9696,N_7975);
nor U11542 (N_11542,N_7934,N_9782);
nor U11543 (N_11543,N_8579,N_9709);
nor U11544 (N_11544,N_8986,N_9354);
and U11545 (N_11545,N_8067,N_9963);
or U11546 (N_11546,N_9044,N_8995);
or U11547 (N_11547,N_7654,N_9015);
and U11548 (N_11548,N_8697,N_7563);
or U11549 (N_11549,N_7835,N_9457);
and U11550 (N_11550,N_7657,N_8389);
nand U11551 (N_11551,N_9217,N_8619);
or U11552 (N_11552,N_9073,N_8879);
nor U11553 (N_11553,N_8960,N_9749);
and U11554 (N_11554,N_9074,N_7755);
or U11555 (N_11555,N_7520,N_9572);
or U11556 (N_11556,N_8672,N_7703);
nor U11557 (N_11557,N_8455,N_9894);
and U11558 (N_11558,N_9636,N_9164);
nor U11559 (N_11559,N_8696,N_9892);
and U11560 (N_11560,N_8017,N_9499);
nand U11561 (N_11561,N_7842,N_8512);
xnor U11562 (N_11562,N_9242,N_9160);
nor U11563 (N_11563,N_8363,N_9989);
nor U11564 (N_11564,N_7903,N_9923);
nand U11565 (N_11565,N_8063,N_8120);
or U11566 (N_11566,N_8346,N_8688);
nor U11567 (N_11567,N_8940,N_9491);
xnor U11568 (N_11568,N_9883,N_9620);
and U11569 (N_11569,N_9384,N_8816);
xor U11570 (N_11570,N_8237,N_8083);
nor U11571 (N_11571,N_8959,N_9598);
nand U11572 (N_11572,N_7519,N_8618);
xor U11573 (N_11573,N_8486,N_9547);
nand U11574 (N_11574,N_7820,N_9946);
or U11575 (N_11575,N_8889,N_9781);
nor U11576 (N_11576,N_8717,N_8169);
nor U11577 (N_11577,N_9107,N_8554);
xnor U11578 (N_11578,N_7563,N_8427);
or U11579 (N_11579,N_9922,N_8155);
xnor U11580 (N_11580,N_7620,N_8111);
nand U11581 (N_11581,N_8988,N_9674);
xor U11582 (N_11582,N_9739,N_8486);
nand U11583 (N_11583,N_9696,N_7629);
nor U11584 (N_11584,N_8779,N_7919);
or U11585 (N_11585,N_9237,N_9356);
nor U11586 (N_11586,N_7951,N_8364);
nor U11587 (N_11587,N_9313,N_9341);
nand U11588 (N_11588,N_7583,N_8323);
xnor U11589 (N_11589,N_8108,N_8482);
nor U11590 (N_11590,N_7728,N_7666);
or U11591 (N_11591,N_8312,N_8925);
xnor U11592 (N_11592,N_8430,N_7533);
and U11593 (N_11593,N_8848,N_8980);
or U11594 (N_11594,N_9966,N_8574);
nand U11595 (N_11595,N_8882,N_9622);
xor U11596 (N_11596,N_7865,N_9797);
xnor U11597 (N_11597,N_7731,N_8995);
xor U11598 (N_11598,N_7920,N_9386);
xor U11599 (N_11599,N_9740,N_9356);
xnor U11600 (N_11600,N_8103,N_7870);
nand U11601 (N_11601,N_9936,N_9346);
or U11602 (N_11602,N_8864,N_8054);
or U11603 (N_11603,N_9322,N_7942);
and U11604 (N_11604,N_9799,N_9899);
nor U11605 (N_11605,N_8327,N_8930);
xnor U11606 (N_11606,N_7850,N_7638);
nor U11607 (N_11607,N_8109,N_7534);
nor U11608 (N_11608,N_8080,N_8309);
xor U11609 (N_11609,N_8106,N_9443);
xnor U11610 (N_11610,N_9833,N_9099);
xor U11611 (N_11611,N_7777,N_8141);
nor U11612 (N_11612,N_8868,N_8308);
xor U11613 (N_11613,N_9085,N_8046);
xor U11614 (N_11614,N_9524,N_8991);
and U11615 (N_11615,N_7598,N_8329);
and U11616 (N_11616,N_7928,N_9608);
or U11617 (N_11617,N_8566,N_9211);
nor U11618 (N_11618,N_7742,N_9924);
or U11619 (N_11619,N_9488,N_9019);
nor U11620 (N_11620,N_8916,N_9403);
nand U11621 (N_11621,N_9458,N_7724);
or U11622 (N_11622,N_8540,N_8788);
and U11623 (N_11623,N_7991,N_8112);
and U11624 (N_11624,N_8192,N_7845);
or U11625 (N_11625,N_9822,N_7621);
or U11626 (N_11626,N_9857,N_9675);
or U11627 (N_11627,N_9244,N_7585);
xnor U11628 (N_11628,N_9065,N_8184);
nor U11629 (N_11629,N_8558,N_8291);
or U11630 (N_11630,N_9447,N_9087);
nand U11631 (N_11631,N_9996,N_9596);
nand U11632 (N_11632,N_8512,N_8773);
or U11633 (N_11633,N_7620,N_9365);
xor U11634 (N_11634,N_9573,N_9210);
or U11635 (N_11635,N_8426,N_8500);
or U11636 (N_11636,N_8125,N_8078);
or U11637 (N_11637,N_9193,N_9431);
nand U11638 (N_11638,N_9096,N_8260);
xnor U11639 (N_11639,N_9380,N_8038);
xor U11640 (N_11640,N_9977,N_9128);
nor U11641 (N_11641,N_8233,N_9811);
xor U11642 (N_11642,N_9483,N_8433);
or U11643 (N_11643,N_8875,N_9199);
nor U11644 (N_11644,N_8978,N_9264);
xnor U11645 (N_11645,N_9884,N_7570);
xnor U11646 (N_11646,N_8973,N_7631);
xnor U11647 (N_11647,N_8921,N_8295);
xor U11648 (N_11648,N_8107,N_8266);
xnor U11649 (N_11649,N_8364,N_8023);
xnor U11650 (N_11650,N_7706,N_8720);
nor U11651 (N_11651,N_8418,N_7743);
or U11652 (N_11652,N_8648,N_9365);
nand U11653 (N_11653,N_7876,N_8567);
nor U11654 (N_11654,N_7583,N_9516);
or U11655 (N_11655,N_8965,N_9269);
nor U11656 (N_11656,N_8052,N_7901);
and U11657 (N_11657,N_9189,N_9015);
nand U11658 (N_11658,N_8797,N_7922);
xnor U11659 (N_11659,N_9966,N_7558);
nor U11660 (N_11660,N_8633,N_8318);
xnor U11661 (N_11661,N_9415,N_9773);
nand U11662 (N_11662,N_7644,N_9656);
or U11663 (N_11663,N_9475,N_7853);
xnor U11664 (N_11664,N_8770,N_9529);
or U11665 (N_11665,N_8794,N_9857);
nor U11666 (N_11666,N_9154,N_8116);
nand U11667 (N_11667,N_7815,N_8998);
nor U11668 (N_11668,N_8351,N_9171);
and U11669 (N_11669,N_8785,N_7907);
nand U11670 (N_11670,N_9645,N_7851);
nand U11671 (N_11671,N_8265,N_9090);
or U11672 (N_11672,N_7784,N_8817);
nor U11673 (N_11673,N_8030,N_7875);
nor U11674 (N_11674,N_7524,N_8516);
or U11675 (N_11675,N_9859,N_9841);
xnor U11676 (N_11676,N_9977,N_9703);
and U11677 (N_11677,N_9711,N_7932);
or U11678 (N_11678,N_8339,N_8609);
nor U11679 (N_11679,N_8526,N_8018);
nand U11680 (N_11680,N_7919,N_9601);
xor U11681 (N_11681,N_7678,N_9554);
xor U11682 (N_11682,N_7685,N_8271);
or U11683 (N_11683,N_9941,N_7529);
nand U11684 (N_11684,N_9846,N_9742);
nor U11685 (N_11685,N_9418,N_9429);
nor U11686 (N_11686,N_9673,N_9513);
nand U11687 (N_11687,N_9901,N_8364);
and U11688 (N_11688,N_9773,N_7735);
nor U11689 (N_11689,N_8361,N_9547);
nor U11690 (N_11690,N_9100,N_9140);
or U11691 (N_11691,N_8527,N_9875);
or U11692 (N_11692,N_9439,N_8369);
or U11693 (N_11693,N_7501,N_8977);
nor U11694 (N_11694,N_9503,N_8018);
xor U11695 (N_11695,N_9416,N_7667);
and U11696 (N_11696,N_9655,N_9747);
xnor U11697 (N_11697,N_9733,N_9672);
and U11698 (N_11698,N_9052,N_7635);
or U11699 (N_11699,N_8996,N_9496);
nor U11700 (N_11700,N_9991,N_7641);
xor U11701 (N_11701,N_8922,N_8405);
nor U11702 (N_11702,N_7884,N_8655);
or U11703 (N_11703,N_8975,N_9983);
nand U11704 (N_11704,N_9653,N_7574);
nand U11705 (N_11705,N_8475,N_8532);
nor U11706 (N_11706,N_9862,N_9725);
nand U11707 (N_11707,N_9347,N_8677);
and U11708 (N_11708,N_8937,N_9076);
xnor U11709 (N_11709,N_8972,N_8581);
and U11710 (N_11710,N_9808,N_8804);
and U11711 (N_11711,N_9304,N_8221);
xor U11712 (N_11712,N_7766,N_9525);
or U11713 (N_11713,N_9564,N_8852);
xnor U11714 (N_11714,N_7586,N_7648);
nor U11715 (N_11715,N_8494,N_9540);
nand U11716 (N_11716,N_8332,N_9777);
nor U11717 (N_11717,N_8278,N_8877);
nor U11718 (N_11718,N_8124,N_9210);
nor U11719 (N_11719,N_7650,N_8542);
nor U11720 (N_11720,N_7617,N_7540);
nand U11721 (N_11721,N_7782,N_8815);
nand U11722 (N_11722,N_7675,N_8840);
or U11723 (N_11723,N_7746,N_9073);
and U11724 (N_11724,N_9663,N_9931);
xor U11725 (N_11725,N_8393,N_9721);
nand U11726 (N_11726,N_8441,N_7537);
xor U11727 (N_11727,N_8384,N_9958);
and U11728 (N_11728,N_7902,N_7610);
and U11729 (N_11729,N_8884,N_7772);
xnor U11730 (N_11730,N_8298,N_8600);
or U11731 (N_11731,N_8521,N_7749);
nand U11732 (N_11732,N_9393,N_8561);
xor U11733 (N_11733,N_7884,N_8145);
nor U11734 (N_11734,N_8617,N_8773);
or U11735 (N_11735,N_8159,N_7865);
xnor U11736 (N_11736,N_7942,N_8815);
nor U11737 (N_11737,N_7532,N_8977);
nand U11738 (N_11738,N_8672,N_8489);
or U11739 (N_11739,N_9766,N_8852);
or U11740 (N_11740,N_8254,N_7628);
and U11741 (N_11741,N_9361,N_9288);
or U11742 (N_11742,N_9643,N_9157);
xnor U11743 (N_11743,N_9314,N_7514);
xor U11744 (N_11744,N_8567,N_9940);
or U11745 (N_11745,N_8029,N_9294);
or U11746 (N_11746,N_8263,N_7669);
and U11747 (N_11747,N_8317,N_7695);
nand U11748 (N_11748,N_8637,N_8786);
nor U11749 (N_11749,N_8412,N_7933);
nor U11750 (N_11750,N_7959,N_9074);
xnor U11751 (N_11751,N_9954,N_7723);
and U11752 (N_11752,N_9854,N_8969);
and U11753 (N_11753,N_9603,N_8927);
nand U11754 (N_11754,N_8270,N_9547);
xor U11755 (N_11755,N_8841,N_9265);
and U11756 (N_11756,N_8043,N_9153);
nand U11757 (N_11757,N_9956,N_7842);
or U11758 (N_11758,N_9148,N_8817);
nand U11759 (N_11759,N_9181,N_8368);
nor U11760 (N_11760,N_9781,N_8092);
xnor U11761 (N_11761,N_9385,N_9046);
and U11762 (N_11762,N_9114,N_8303);
xnor U11763 (N_11763,N_7804,N_9744);
nand U11764 (N_11764,N_8998,N_8176);
nor U11765 (N_11765,N_8290,N_9581);
and U11766 (N_11766,N_8541,N_8434);
or U11767 (N_11767,N_9641,N_9050);
nor U11768 (N_11768,N_7601,N_9175);
xnor U11769 (N_11769,N_9327,N_9419);
xnor U11770 (N_11770,N_9775,N_7699);
xnor U11771 (N_11771,N_9363,N_9218);
or U11772 (N_11772,N_9463,N_8812);
or U11773 (N_11773,N_9401,N_9808);
nor U11774 (N_11774,N_9696,N_8872);
nor U11775 (N_11775,N_9710,N_9698);
or U11776 (N_11776,N_9718,N_8384);
and U11777 (N_11777,N_7545,N_8456);
xnor U11778 (N_11778,N_7810,N_7701);
nor U11779 (N_11779,N_8543,N_8195);
nor U11780 (N_11780,N_9858,N_9388);
or U11781 (N_11781,N_9208,N_9506);
nand U11782 (N_11782,N_9910,N_9159);
xnor U11783 (N_11783,N_9537,N_9518);
and U11784 (N_11784,N_9889,N_8868);
nor U11785 (N_11785,N_8951,N_9855);
xnor U11786 (N_11786,N_8938,N_7711);
nor U11787 (N_11787,N_8435,N_7871);
nand U11788 (N_11788,N_7848,N_7695);
and U11789 (N_11789,N_7871,N_7502);
nor U11790 (N_11790,N_7802,N_9283);
or U11791 (N_11791,N_9399,N_8547);
nor U11792 (N_11792,N_8779,N_9598);
nor U11793 (N_11793,N_9466,N_7941);
nand U11794 (N_11794,N_9616,N_7893);
nor U11795 (N_11795,N_7578,N_8461);
or U11796 (N_11796,N_9256,N_9336);
nand U11797 (N_11797,N_8704,N_9629);
nor U11798 (N_11798,N_9047,N_8923);
nor U11799 (N_11799,N_7787,N_9868);
nor U11800 (N_11800,N_8067,N_9343);
or U11801 (N_11801,N_7983,N_9289);
and U11802 (N_11802,N_9546,N_9628);
nor U11803 (N_11803,N_9034,N_7653);
nand U11804 (N_11804,N_8471,N_9617);
nor U11805 (N_11805,N_9608,N_7507);
nand U11806 (N_11806,N_7750,N_9503);
nand U11807 (N_11807,N_8313,N_7836);
nand U11808 (N_11808,N_8770,N_9412);
nor U11809 (N_11809,N_9584,N_8509);
xor U11810 (N_11810,N_9832,N_9926);
or U11811 (N_11811,N_7929,N_8311);
nor U11812 (N_11812,N_7714,N_9504);
xnor U11813 (N_11813,N_8462,N_8439);
nor U11814 (N_11814,N_9601,N_8765);
and U11815 (N_11815,N_8302,N_8745);
nand U11816 (N_11816,N_7906,N_7687);
and U11817 (N_11817,N_8899,N_8521);
nor U11818 (N_11818,N_8466,N_8685);
nand U11819 (N_11819,N_7820,N_7861);
and U11820 (N_11820,N_9854,N_8321);
and U11821 (N_11821,N_8520,N_9533);
xor U11822 (N_11822,N_9710,N_8440);
xnor U11823 (N_11823,N_8301,N_8050);
nor U11824 (N_11824,N_9427,N_8822);
xnor U11825 (N_11825,N_8048,N_9632);
and U11826 (N_11826,N_9532,N_8271);
nand U11827 (N_11827,N_9990,N_8361);
nor U11828 (N_11828,N_8091,N_8536);
and U11829 (N_11829,N_9686,N_9758);
or U11830 (N_11830,N_9870,N_9379);
xor U11831 (N_11831,N_8423,N_8844);
nand U11832 (N_11832,N_7617,N_7794);
or U11833 (N_11833,N_7796,N_9846);
or U11834 (N_11834,N_8837,N_8266);
nor U11835 (N_11835,N_8677,N_8440);
xnor U11836 (N_11836,N_9261,N_8231);
nor U11837 (N_11837,N_9627,N_7919);
or U11838 (N_11838,N_8883,N_8259);
nor U11839 (N_11839,N_9888,N_7563);
nor U11840 (N_11840,N_9252,N_9631);
xnor U11841 (N_11841,N_8592,N_9846);
nor U11842 (N_11842,N_9174,N_9429);
xor U11843 (N_11843,N_9407,N_8124);
nand U11844 (N_11844,N_9863,N_8141);
and U11845 (N_11845,N_9824,N_9224);
nand U11846 (N_11846,N_8400,N_9011);
xor U11847 (N_11847,N_8410,N_9094);
xor U11848 (N_11848,N_7903,N_9673);
xor U11849 (N_11849,N_8683,N_9282);
nor U11850 (N_11850,N_9575,N_9474);
nand U11851 (N_11851,N_8164,N_8436);
or U11852 (N_11852,N_9001,N_8490);
nand U11853 (N_11853,N_9530,N_9806);
or U11854 (N_11854,N_9902,N_9573);
nor U11855 (N_11855,N_7613,N_9176);
nor U11856 (N_11856,N_8400,N_8324);
xor U11857 (N_11857,N_9400,N_8821);
nand U11858 (N_11858,N_8038,N_8210);
and U11859 (N_11859,N_8443,N_9643);
xor U11860 (N_11860,N_7800,N_8146);
or U11861 (N_11861,N_7748,N_7889);
and U11862 (N_11862,N_9429,N_8009);
nand U11863 (N_11863,N_8423,N_9101);
and U11864 (N_11864,N_7976,N_8642);
nor U11865 (N_11865,N_7715,N_9645);
nand U11866 (N_11866,N_8380,N_9033);
xnor U11867 (N_11867,N_9523,N_8204);
nor U11868 (N_11868,N_9952,N_9747);
xnor U11869 (N_11869,N_8694,N_8781);
and U11870 (N_11870,N_9819,N_9439);
nor U11871 (N_11871,N_8834,N_7758);
or U11872 (N_11872,N_7511,N_8008);
or U11873 (N_11873,N_9750,N_8790);
nor U11874 (N_11874,N_8125,N_9958);
nand U11875 (N_11875,N_8279,N_7908);
or U11876 (N_11876,N_9668,N_9938);
nand U11877 (N_11877,N_7951,N_8187);
xnor U11878 (N_11878,N_9590,N_8243);
nand U11879 (N_11879,N_7828,N_8240);
or U11880 (N_11880,N_9365,N_7608);
xor U11881 (N_11881,N_7974,N_9885);
and U11882 (N_11882,N_9140,N_9171);
and U11883 (N_11883,N_9701,N_9250);
xnor U11884 (N_11884,N_7746,N_8340);
or U11885 (N_11885,N_8234,N_9349);
or U11886 (N_11886,N_9542,N_8793);
nand U11887 (N_11887,N_8702,N_9596);
or U11888 (N_11888,N_7732,N_9307);
xnor U11889 (N_11889,N_7801,N_9918);
and U11890 (N_11890,N_8436,N_8538);
or U11891 (N_11891,N_8055,N_9313);
or U11892 (N_11892,N_8705,N_9858);
xor U11893 (N_11893,N_7689,N_8858);
and U11894 (N_11894,N_8877,N_8890);
nor U11895 (N_11895,N_8049,N_8593);
and U11896 (N_11896,N_9844,N_9075);
or U11897 (N_11897,N_8929,N_9661);
nor U11898 (N_11898,N_9552,N_7790);
xnor U11899 (N_11899,N_8802,N_9883);
or U11900 (N_11900,N_8324,N_9373);
or U11901 (N_11901,N_9729,N_8990);
and U11902 (N_11902,N_9091,N_8925);
xnor U11903 (N_11903,N_8491,N_7625);
nand U11904 (N_11904,N_8954,N_9144);
xnor U11905 (N_11905,N_9808,N_8689);
nand U11906 (N_11906,N_9267,N_8541);
or U11907 (N_11907,N_8507,N_9712);
nor U11908 (N_11908,N_8324,N_8605);
nor U11909 (N_11909,N_9831,N_8148);
or U11910 (N_11910,N_7631,N_8171);
and U11911 (N_11911,N_9162,N_9278);
xor U11912 (N_11912,N_9892,N_8621);
or U11913 (N_11913,N_8585,N_7650);
nand U11914 (N_11914,N_9411,N_9694);
nand U11915 (N_11915,N_9380,N_9744);
nor U11916 (N_11916,N_8523,N_9449);
or U11917 (N_11917,N_9172,N_9003);
nand U11918 (N_11918,N_7652,N_9137);
nand U11919 (N_11919,N_9031,N_7773);
and U11920 (N_11920,N_9449,N_9989);
nor U11921 (N_11921,N_9503,N_9602);
nand U11922 (N_11922,N_9196,N_8665);
and U11923 (N_11923,N_7548,N_8336);
nand U11924 (N_11924,N_9080,N_9885);
or U11925 (N_11925,N_9833,N_7878);
and U11926 (N_11926,N_9387,N_7914);
and U11927 (N_11927,N_9131,N_7521);
or U11928 (N_11928,N_9939,N_9370);
nand U11929 (N_11929,N_8059,N_9636);
or U11930 (N_11930,N_8416,N_8169);
nand U11931 (N_11931,N_9534,N_9524);
nor U11932 (N_11932,N_9542,N_9767);
nand U11933 (N_11933,N_7528,N_8130);
nand U11934 (N_11934,N_8545,N_9204);
or U11935 (N_11935,N_8187,N_8233);
nand U11936 (N_11936,N_7897,N_9357);
or U11937 (N_11937,N_9580,N_9608);
nor U11938 (N_11938,N_9000,N_8223);
nand U11939 (N_11939,N_9030,N_8436);
and U11940 (N_11940,N_9909,N_9949);
nor U11941 (N_11941,N_8614,N_8626);
and U11942 (N_11942,N_9775,N_8958);
nand U11943 (N_11943,N_8743,N_9389);
nand U11944 (N_11944,N_9713,N_8341);
and U11945 (N_11945,N_7936,N_7957);
xnor U11946 (N_11946,N_9732,N_8163);
nand U11947 (N_11947,N_9047,N_7851);
or U11948 (N_11948,N_8968,N_9996);
and U11949 (N_11949,N_8374,N_9517);
nand U11950 (N_11950,N_9450,N_7743);
xor U11951 (N_11951,N_7578,N_9491);
nand U11952 (N_11952,N_9430,N_7807);
and U11953 (N_11953,N_9872,N_8651);
or U11954 (N_11954,N_8140,N_8036);
and U11955 (N_11955,N_9290,N_9945);
xor U11956 (N_11956,N_9811,N_9184);
nand U11957 (N_11957,N_9190,N_7877);
nand U11958 (N_11958,N_8655,N_7627);
nor U11959 (N_11959,N_8736,N_8080);
and U11960 (N_11960,N_8932,N_8320);
and U11961 (N_11961,N_7804,N_8533);
and U11962 (N_11962,N_7585,N_7847);
nand U11963 (N_11963,N_9512,N_8722);
and U11964 (N_11964,N_8874,N_7514);
nand U11965 (N_11965,N_9356,N_9551);
nand U11966 (N_11966,N_8784,N_8724);
nor U11967 (N_11967,N_8500,N_8110);
and U11968 (N_11968,N_9837,N_8851);
nor U11969 (N_11969,N_9589,N_9545);
and U11970 (N_11970,N_8033,N_8767);
and U11971 (N_11971,N_8710,N_8940);
and U11972 (N_11972,N_7568,N_7604);
and U11973 (N_11973,N_9599,N_9503);
nand U11974 (N_11974,N_8064,N_9381);
nand U11975 (N_11975,N_9824,N_8582);
nor U11976 (N_11976,N_7582,N_9713);
xnor U11977 (N_11977,N_7819,N_7928);
and U11978 (N_11978,N_8903,N_8841);
nand U11979 (N_11979,N_8556,N_8309);
nor U11980 (N_11980,N_9802,N_8499);
nor U11981 (N_11981,N_8478,N_9176);
or U11982 (N_11982,N_9843,N_9572);
or U11983 (N_11983,N_8652,N_9258);
nand U11984 (N_11984,N_9517,N_7532);
and U11985 (N_11985,N_7729,N_9396);
or U11986 (N_11986,N_9251,N_8525);
nor U11987 (N_11987,N_7809,N_9113);
or U11988 (N_11988,N_8124,N_9634);
or U11989 (N_11989,N_9824,N_8161);
and U11990 (N_11990,N_9298,N_9593);
and U11991 (N_11991,N_8087,N_8005);
nor U11992 (N_11992,N_7612,N_9372);
nand U11993 (N_11993,N_9961,N_9280);
nand U11994 (N_11994,N_7949,N_7711);
xor U11995 (N_11995,N_8469,N_8982);
or U11996 (N_11996,N_9716,N_9319);
xnor U11997 (N_11997,N_8159,N_7714);
nor U11998 (N_11998,N_9578,N_7657);
or U11999 (N_11999,N_8239,N_8901);
nor U12000 (N_12000,N_7940,N_8898);
or U12001 (N_12001,N_9419,N_8864);
and U12002 (N_12002,N_7785,N_8103);
and U12003 (N_12003,N_8211,N_9603);
or U12004 (N_12004,N_8559,N_8099);
nor U12005 (N_12005,N_7882,N_9658);
or U12006 (N_12006,N_9545,N_7500);
nand U12007 (N_12007,N_8856,N_7612);
or U12008 (N_12008,N_8216,N_8888);
xnor U12009 (N_12009,N_9213,N_8620);
nor U12010 (N_12010,N_8328,N_7674);
nor U12011 (N_12011,N_7991,N_8919);
nand U12012 (N_12012,N_9891,N_9079);
and U12013 (N_12013,N_8083,N_8971);
nand U12014 (N_12014,N_7797,N_9923);
xnor U12015 (N_12015,N_8065,N_8175);
nor U12016 (N_12016,N_8055,N_8145);
nor U12017 (N_12017,N_9413,N_7544);
nor U12018 (N_12018,N_8517,N_9983);
and U12019 (N_12019,N_8740,N_7602);
nor U12020 (N_12020,N_8268,N_8147);
nand U12021 (N_12021,N_9664,N_8373);
nand U12022 (N_12022,N_9350,N_8141);
and U12023 (N_12023,N_9043,N_7843);
xnor U12024 (N_12024,N_9135,N_7623);
nand U12025 (N_12025,N_8078,N_8828);
and U12026 (N_12026,N_7858,N_8342);
nor U12027 (N_12027,N_8263,N_9628);
or U12028 (N_12028,N_8558,N_8972);
nand U12029 (N_12029,N_7860,N_7559);
xor U12030 (N_12030,N_8291,N_9383);
and U12031 (N_12031,N_8989,N_9202);
xor U12032 (N_12032,N_9733,N_8694);
or U12033 (N_12033,N_9869,N_8800);
and U12034 (N_12034,N_8328,N_9862);
xor U12035 (N_12035,N_8103,N_8689);
xnor U12036 (N_12036,N_8935,N_9274);
xor U12037 (N_12037,N_8161,N_9804);
xnor U12038 (N_12038,N_8861,N_8627);
or U12039 (N_12039,N_7957,N_9102);
nand U12040 (N_12040,N_9768,N_9989);
nand U12041 (N_12041,N_8921,N_8047);
nand U12042 (N_12042,N_8420,N_9037);
nor U12043 (N_12043,N_8747,N_9367);
or U12044 (N_12044,N_8053,N_9215);
xor U12045 (N_12045,N_8187,N_8931);
and U12046 (N_12046,N_8656,N_8232);
xnor U12047 (N_12047,N_9844,N_9439);
and U12048 (N_12048,N_9565,N_7622);
xnor U12049 (N_12049,N_9450,N_9052);
and U12050 (N_12050,N_9294,N_9277);
or U12051 (N_12051,N_9350,N_7786);
or U12052 (N_12052,N_8359,N_9450);
or U12053 (N_12053,N_8296,N_9953);
nand U12054 (N_12054,N_7539,N_9449);
or U12055 (N_12055,N_9112,N_7565);
xnor U12056 (N_12056,N_8322,N_7791);
nand U12057 (N_12057,N_8738,N_7644);
or U12058 (N_12058,N_7707,N_8980);
nand U12059 (N_12059,N_8480,N_7895);
nand U12060 (N_12060,N_8926,N_8944);
xor U12061 (N_12061,N_9458,N_9449);
and U12062 (N_12062,N_7804,N_8713);
xor U12063 (N_12063,N_8869,N_7509);
nor U12064 (N_12064,N_7951,N_8288);
and U12065 (N_12065,N_8494,N_9104);
or U12066 (N_12066,N_8116,N_9756);
or U12067 (N_12067,N_8621,N_9642);
or U12068 (N_12068,N_8744,N_9557);
nor U12069 (N_12069,N_9502,N_7594);
nor U12070 (N_12070,N_7635,N_8617);
or U12071 (N_12071,N_7676,N_8930);
or U12072 (N_12072,N_7515,N_8618);
nand U12073 (N_12073,N_9880,N_8822);
or U12074 (N_12074,N_9610,N_7754);
nand U12075 (N_12075,N_8026,N_8245);
and U12076 (N_12076,N_9056,N_7688);
nand U12077 (N_12077,N_7787,N_8539);
and U12078 (N_12078,N_7578,N_8451);
and U12079 (N_12079,N_9304,N_9227);
nand U12080 (N_12080,N_8325,N_9811);
xor U12081 (N_12081,N_9636,N_8331);
xor U12082 (N_12082,N_9002,N_8908);
and U12083 (N_12083,N_9599,N_8107);
and U12084 (N_12084,N_8450,N_8166);
nand U12085 (N_12085,N_7615,N_8721);
xnor U12086 (N_12086,N_8699,N_9555);
and U12087 (N_12087,N_9102,N_9710);
xor U12088 (N_12088,N_8089,N_8568);
and U12089 (N_12089,N_8861,N_9946);
nand U12090 (N_12090,N_9424,N_9331);
or U12091 (N_12091,N_9850,N_9309);
xor U12092 (N_12092,N_8257,N_9645);
or U12093 (N_12093,N_9089,N_8277);
nand U12094 (N_12094,N_8714,N_7540);
nand U12095 (N_12095,N_8320,N_8735);
nand U12096 (N_12096,N_8557,N_8457);
nor U12097 (N_12097,N_7615,N_7559);
xor U12098 (N_12098,N_9950,N_8974);
nor U12099 (N_12099,N_9595,N_9903);
nand U12100 (N_12100,N_9061,N_8698);
or U12101 (N_12101,N_8302,N_8442);
nor U12102 (N_12102,N_7765,N_9591);
nand U12103 (N_12103,N_8743,N_7793);
nor U12104 (N_12104,N_9154,N_7968);
xor U12105 (N_12105,N_8481,N_7625);
nand U12106 (N_12106,N_9194,N_7837);
or U12107 (N_12107,N_7660,N_9949);
and U12108 (N_12108,N_9593,N_8134);
nand U12109 (N_12109,N_8661,N_8649);
nor U12110 (N_12110,N_7694,N_8250);
xnor U12111 (N_12111,N_9911,N_7542);
or U12112 (N_12112,N_7776,N_7604);
nor U12113 (N_12113,N_7661,N_9865);
nor U12114 (N_12114,N_7804,N_9127);
or U12115 (N_12115,N_7673,N_9380);
or U12116 (N_12116,N_7517,N_7886);
nand U12117 (N_12117,N_8580,N_9604);
nor U12118 (N_12118,N_8545,N_8536);
or U12119 (N_12119,N_8663,N_7923);
xnor U12120 (N_12120,N_9183,N_8303);
and U12121 (N_12121,N_7765,N_8445);
nand U12122 (N_12122,N_9767,N_8433);
and U12123 (N_12123,N_7558,N_9373);
or U12124 (N_12124,N_8237,N_9230);
nor U12125 (N_12125,N_9018,N_9155);
and U12126 (N_12126,N_8409,N_9107);
xnor U12127 (N_12127,N_8957,N_7829);
or U12128 (N_12128,N_9557,N_8372);
or U12129 (N_12129,N_8370,N_8981);
nand U12130 (N_12130,N_9863,N_9506);
nand U12131 (N_12131,N_8852,N_9632);
nor U12132 (N_12132,N_9631,N_8263);
and U12133 (N_12133,N_9244,N_9346);
nor U12134 (N_12134,N_7796,N_8936);
and U12135 (N_12135,N_7563,N_8159);
nand U12136 (N_12136,N_9658,N_9621);
and U12137 (N_12137,N_8454,N_9835);
and U12138 (N_12138,N_8127,N_7690);
nor U12139 (N_12139,N_9502,N_7740);
nor U12140 (N_12140,N_8352,N_8074);
nand U12141 (N_12141,N_8573,N_7682);
or U12142 (N_12142,N_8531,N_8559);
nand U12143 (N_12143,N_9509,N_8085);
xnor U12144 (N_12144,N_9403,N_8884);
or U12145 (N_12145,N_9982,N_9438);
nand U12146 (N_12146,N_8547,N_7526);
and U12147 (N_12147,N_9563,N_9939);
nand U12148 (N_12148,N_8337,N_8159);
nor U12149 (N_12149,N_9691,N_9276);
xor U12150 (N_12150,N_9315,N_9494);
nor U12151 (N_12151,N_9645,N_8360);
or U12152 (N_12152,N_8802,N_8886);
nor U12153 (N_12153,N_8987,N_8664);
or U12154 (N_12154,N_9039,N_9143);
or U12155 (N_12155,N_9767,N_7684);
and U12156 (N_12156,N_9503,N_7519);
or U12157 (N_12157,N_8991,N_7796);
nand U12158 (N_12158,N_7890,N_8259);
and U12159 (N_12159,N_8934,N_9810);
xor U12160 (N_12160,N_8986,N_8238);
or U12161 (N_12161,N_8136,N_8926);
or U12162 (N_12162,N_9130,N_8317);
nand U12163 (N_12163,N_8705,N_8914);
xor U12164 (N_12164,N_9946,N_8137);
and U12165 (N_12165,N_8858,N_9863);
or U12166 (N_12166,N_9555,N_8460);
and U12167 (N_12167,N_8842,N_8021);
xnor U12168 (N_12168,N_8403,N_7564);
or U12169 (N_12169,N_8081,N_9061);
and U12170 (N_12170,N_8773,N_9048);
nor U12171 (N_12171,N_9761,N_8037);
or U12172 (N_12172,N_7531,N_9427);
or U12173 (N_12173,N_8444,N_9195);
and U12174 (N_12174,N_9138,N_8752);
xor U12175 (N_12175,N_8664,N_7787);
and U12176 (N_12176,N_8288,N_9897);
or U12177 (N_12177,N_7690,N_9699);
xor U12178 (N_12178,N_8660,N_9168);
or U12179 (N_12179,N_8456,N_7679);
xor U12180 (N_12180,N_8967,N_9508);
or U12181 (N_12181,N_8374,N_8016);
nand U12182 (N_12182,N_8922,N_9997);
or U12183 (N_12183,N_9124,N_7810);
or U12184 (N_12184,N_7643,N_8412);
or U12185 (N_12185,N_9334,N_9378);
xor U12186 (N_12186,N_7946,N_7636);
or U12187 (N_12187,N_9715,N_7825);
xor U12188 (N_12188,N_9196,N_9671);
and U12189 (N_12189,N_9871,N_9077);
nand U12190 (N_12190,N_8131,N_8102);
nor U12191 (N_12191,N_8046,N_9762);
and U12192 (N_12192,N_8559,N_9484);
or U12193 (N_12193,N_8232,N_7884);
or U12194 (N_12194,N_9770,N_9723);
and U12195 (N_12195,N_9547,N_9703);
nor U12196 (N_12196,N_9877,N_8961);
nor U12197 (N_12197,N_8231,N_8310);
and U12198 (N_12198,N_9983,N_7878);
nor U12199 (N_12199,N_7934,N_9569);
nor U12200 (N_12200,N_8916,N_8625);
or U12201 (N_12201,N_8874,N_7874);
and U12202 (N_12202,N_8902,N_8951);
and U12203 (N_12203,N_7775,N_8313);
and U12204 (N_12204,N_8286,N_9890);
xor U12205 (N_12205,N_8354,N_8762);
xnor U12206 (N_12206,N_8970,N_7871);
nand U12207 (N_12207,N_7819,N_9264);
nand U12208 (N_12208,N_8466,N_8273);
and U12209 (N_12209,N_8222,N_9856);
or U12210 (N_12210,N_8257,N_8244);
nor U12211 (N_12211,N_7658,N_8097);
xnor U12212 (N_12212,N_7744,N_7790);
nand U12213 (N_12213,N_9642,N_8577);
or U12214 (N_12214,N_8818,N_9955);
nand U12215 (N_12215,N_8191,N_9371);
and U12216 (N_12216,N_8214,N_7947);
and U12217 (N_12217,N_9975,N_9372);
xnor U12218 (N_12218,N_8488,N_9436);
and U12219 (N_12219,N_9771,N_9855);
or U12220 (N_12220,N_7918,N_7501);
xor U12221 (N_12221,N_8057,N_9533);
nand U12222 (N_12222,N_9902,N_8351);
nor U12223 (N_12223,N_7607,N_8651);
or U12224 (N_12224,N_8110,N_9618);
or U12225 (N_12225,N_7603,N_9997);
and U12226 (N_12226,N_7610,N_7769);
nor U12227 (N_12227,N_7989,N_9945);
and U12228 (N_12228,N_7876,N_8653);
and U12229 (N_12229,N_9429,N_8065);
or U12230 (N_12230,N_8341,N_9523);
or U12231 (N_12231,N_9645,N_9662);
nor U12232 (N_12232,N_7523,N_9946);
or U12233 (N_12233,N_8627,N_7526);
xnor U12234 (N_12234,N_8400,N_7831);
and U12235 (N_12235,N_8865,N_9913);
nor U12236 (N_12236,N_9119,N_7717);
xnor U12237 (N_12237,N_8336,N_9168);
nor U12238 (N_12238,N_8983,N_8643);
nand U12239 (N_12239,N_8040,N_8971);
nor U12240 (N_12240,N_8948,N_9135);
and U12241 (N_12241,N_8953,N_9527);
xnor U12242 (N_12242,N_7698,N_9349);
and U12243 (N_12243,N_8695,N_7842);
nor U12244 (N_12244,N_9342,N_9828);
or U12245 (N_12245,N_8492,N_7647);
nand U12246 (N_12246,N_8421,N_9852);
nor U12247 (N_12247,N_9947,N_8660);
xor U12248 (N_12248,N_7617,N_7989);
or U12249 (N_12249,N_8621,N_8252);
or U12250 (N_12250,N_9590,N_9722);
or U12251 (N_12251,N_9768,N_9743);
xnor U12252 (N_12252,N_8985,N_9008);
xor U12253 (N_12253,N_8023,N_8938);
or U12254 (N_12254,N_9210,N_9396);
or U12255 (N_12255,N_7819,N_8154);
or U12256 (N_12256,N_7760,N_8341);
nor U12257 (N_12257,N_8731,N_7956);
and U12258 (N_12258,N_7538,N_7766);
xor U12259 (N_12259,N_8463,N_9898);
nand U12260 (N_12260,N_8752,N_8703);
nor U12261 (N_12261,N_8546,N_7939);
and U12262 (N_12262,N_8338,N_9903);
xnor U12263 (N_12263,N_7663,N_8754);
xor U12264 (N_12264,N_8146,N_8628);
and U12265 (N_12265,N_9177,N_8241);
nor U12266 (N_12266,N_8977,N_7715);
nand U12267 (N_12267,N_8996,N_8204);
xor U12268 (N_12268,N_7560,N_7880);
nand U12269 (N_12269,N_7627,N_8036);
or U12270 (N_12270,N_7636,N_8369);
or U12271 (N_12271,N_8002,N_9855);
nor U12272 (N_12272,N_8131,N_9339);
and U12273 (N_12273,N_7640,N_8463);
xnor U12274 (N_12274,N_9978,N_8741);
and U12275 (N_12275,N_7590,N_7820);
or U12276 (N_12276,N_8766,N_9875);
or U12277 (N_12277,N_9199,N_9705);
and U12278 (N_12278,N_9792,N_8253);
and U12279 (N_12279,N_8925,N_9935);
nor U12280 (N_12280,N_9383,N_7859);
or U12281 (N_12281,N_9089,N_7856);
nand U12282 (N_12282,N_7553,N_9760);
nor U12283 (N_12283,N_7960,N_9601);
and U12284 (N_12284,N_7963,N_9267);
nand U12285 (N_12285,N_9677,N_8072);
and U12286 (N_12286,N_8828,N_8169);
xor U12287 (N_12287,N_8950,N_7597);
xnor U12288 (N_12288,N_8477,N_8393);
and U12289 (N_12289,N_9982,N_8786);
and U12290 (N_12290,N_8650,N_8892);
nand U12291 (N_12291,N_8433,N_8697);
and U12292 (N_12292,N_8079,N_8470);
xor U12293 (N_12293,N_7719,N_9269);
and U12294 (N_12294,N_8635,N_9605);
nor U12295 (N_12295,N_8531,N_7776);
xor U12296 (N_12296,N_8973,N_9268);
xnor U12297 (N_12297,N_9030,N_8064);
or U12298 (N_12298,N_8438,N_9458);
xor U12299 (N_12299,N_8806,N_9513);
nand U12300 (N_12300,N_8015,N_7553);
nor U12301 (N_12301,N_8165,N_9923);
or U12302 (N_12302,N_9015,N_7562);
nor U12303 (N_12303,N_9923,N_8943);
and U12304 (N_12304,N_8822,N_9070);
and U12305 (N_12305,N_9748,N_9455);
xnor U12306 (N_12306,N_9354,N_7777);
nand U12307 (N_12307,N_9607,N_9422);
xor U12308 (N_12308,N_8453,N_8982);
and U12309 (N_12309,N_7593,N_9554);
nor U12310 (N_12310,N_7974,N_7916);
xnor U12311 (N_12311,N_8763,N_8706);
nand U12312 (N_12312,N_9348,N_9024);
and U12313 (N_12313,N_8118,N_7891);
and U12314 (N_12314,N_9846,N_9294);
xor U12315 (N_12315,N_7516,N_9926);
nor U12316 (N_12316,N_8818,N_7727);
xor U12317 (N_12317,N_9195,N_7561);
or U12318 (N_12318,N_8283,N_9489);
xnor U12319 (N_12319,N_9899,N_7883);
and U12320 (N_12320,N_8223,N_7946);
nor U12321 (N_12321,N_8687,N_8165);
nand U12322 (N_12322,N_9777,N_8073);
or U12323 (N_12323,N_8847,N_7500);
and U12324 (N_12324,N_9809,N_8866);
and U12325 (N_12325,N_7961,N_8754);
or U12326 (N_12326,N_9107,N_7913);
nand U12327 (N_12327,N_9139,N_9907);
nand U12328 (N_12328,N_9528,N_7937);
xnor U12329 (N_12329,N_8264,N_9060);
and U12330 (N_12330,N_8300,N_8470);
or U12331 (N_12331,N_7821,N_8158);
xnor U12332 (N_12332,N_7981,N_8880);
xnor U12333 (N_12333,N_9816,N_7932);
or U12334 (N_12334,N_7810,N_9067);
nor U12335 (N_12335,N_9607,N_9926);
xnor U12336 (N_12336,N_7633,N_8972);
nor U12337 (N_12337,N_9655,N_8303);
nor U12338 (N_12338,N_7724,N_9494);
xor U12339 (N_12339,N_8634,N_8114);
or U12340 (N_12340,N_7891,N_8927);
nor U12341 (N_12341,N_7608,N_7761);
or U12342 (N_12342,N_8932,N_9847);
or U12343 (N_12343,N_8771,N_8563);
nor U12344 (N_12344,N_8663,N_8644);
xor U12345 (N_12345,N_8207,N_9286);
xnor U12346 (N_12346,N_9990,N_8350);
and U12347 (N_12347,N_9998,N_9190);
nand U12348 (N_12348,N_9404,N_8334);
xor U12349 (N_12349,N_8615,N_9628);
nand U12350 (N_12350,N_8292,N_9339);
nand U12351 (N_12351,N_7701,N_8485);
xnor U12352 (N_12352,N_8106,N_8390);
nor U12353 (N_12353,N_7984,N_9540);
and U12354 (N_12354,N_8187,N_8242);
or U12355 (N_12355,N_8421,N_9433);
nor U12356 (N_12356,N_9489,N_8204);
or U12357 (N_12357,N_8095,N_8392);
or U12358 (N_12358,N_9423,N_9926);
and U12359 (N_12359,N_9563,N_7898);
or U12360 (N_12360,N_9689,N_7963);
or U12361 (N_12361,N_8241,N_8408);
nand U12362 (N_12362,N_7674,N_7857);
and U12363 (N_12363,N_8475,N_9264);
or U12364 (N_12364,N_7833,N_9839);
xor U12365 (N_12365,N_7560,N_9722);
nand U12366 (N_12366,N_7585,N_7867);
nand U12367 (N_12367,N_8222,N_8881);
or U12368 (N_12368,N_8988,N_8308);
or U12369 (N_12369,N_9221,N_9417);
nand U12370 (N_12370,N_8608,N_9300);
xnor U12371 (N_12371,N_7578,N_7870);
or U12372 (N_12372,N_9588,N_9328);
nor U12373 (N_12373,N_7629,N_7830);
nor U12374 (N_12374,N_7897,N_7726);
xnor U12375 (N_12375,N_7657,N_8015);
nor U12376 (N_12376,N_8618,N_9328);
nand U12377 (N_12377,N_9118,N_9506);
nand U12378 (N_12378,N_8324,N_8700);
nor U12379 (N_12379,N_8245,N_9621);
xor U12380 (N_12380,N_9521,N_7744);
xor U12381 (N_12381,N_9563,N_8269);
and U12382 (N_12382,N_9152,N_9480);
and U12383 (N_12383,N_7935,N_8206);
and U12384 (N_12384,N_7715,N_8991);
or U12385 (N_12385,N_8189,N_8233);
or U12386 (N_12386,N_9747,N_9688);
and U12387 (N_12387,N_9098,N_7646);
and U12388 (N_12388,N_7933,N_9397);
nand U12389 (N_12389,N_9110,N_8884);
and U12390 (N_12390,N_8353,N_9530);
and U12391 (N_12391,N_8872,N_7992);
nand U12392 (N_12392,N_9707,N_9663);
xnor U12393 (N_12393,N_7813,N_9452);
and U12394 (N_12394,N_9528,N_8044);
xnor U12395 (N_12395,N_8663,N_9384);
and U12396 (N_12396,N_8227,N_9147);
and U12397 (N_12397,N_9485,N_9640);
nor U12398 (N_12398,N_8959,N_9495);
nor U12399 (N_12399,N_9387,N_7717);
nand U12400 (N_12400,N_8162,N_8724);
and U12401 (N_12401,N_9685,N_8516);
nand U12402 (N_12402,N_9117,N_8852);
nand U12403 (N_12403,N_8838,N_8418);
xor U12404 (N_12404,N_8762,N_8604);
nor U12405 (N_12405,N_7683,N_9243);
or U12406 (N_12406,N_9385,N_9212);
or U12407 (N_12407,N_9523,N_9444);
nand U12408 (N_12408,N_8266,N_8080);
nand U12409 (N_12409,N_8025,N_7937);
and U12410 (N_12410,N_7507,N_9897);
or U12411 (N_12411,N_8099,N_9716);
and U12412 (N_12412,N_9846,N_8298);
and U12413 (N_12413,N_7935,N_8844);
nor U12414 (N_12414,N_7745,N_9741);
nor U12415 (N_12415,N_9858,N_9535);
xor U12416 (N_12416,N_7845,N_7682);
nand U12417 (N_12417,N_9081,N_9948);
nor U12418 (N_12418,N_9151,N_7716);
or U12419 (N_12419,N_8985,N_8355);
xnor U12420 (N_12420,N_8721,N_9333);
nand U12421 (N_12421,N_8110,N_9123);
nor U12422 (N_12422,N_8635,N_7698);
xnor U12423 (N_12423,N_9408,N_9963);
nand U12424 (N_12424,N_9440,N_8548);
nand U12425 (N_12425,N_9700,N_9766);
xnor U12426 (N_12426,N_8494,N_8352);
nor U12427 (N_12427,N_8347,N_9283);
and U12428 (N_12428,N_9801,N_9300);
nor U12429 (N_12429,N_9660,N_8461);
and U12430 (N_12430,N_9769,N_8397);
xor U12431 (N_12431,N_9161,N_9603);
nor U12432 (N_12432,N_9097,N_7626);
nand U12433 (N_12433,N_8775,N_8677);
nor U12434 (N_12434,N_9992,N_8305);
or U12435 (N_12435,N_8678,N_9769);
or U12436 (N_12436,N_9335,N_8707);
nor U12437 (N_12437,N_8223,N_7635);
nand U12438 (N_12438,N_8376,N_9119);
and U12439 (N_12439,N_9072,N_8706);
and U12440 (N_12440,N_7746,N_8064);
and U12441 (N_12441,N_9803,N_9597);
and U12442 (N_12442,N_9843,N_8271);
or U12443 (N_12443,N_7589,N_9338);
and U12444 (N_12444,N_9554,N_8439);
nand U12445 (N_12445,N_9549,N_7857);
nand U12446 (N_12446,N_9163,N_8427);
nor U12447 (N_12447,N_8305,N_9083);
and U12448 (N_12448,N_7924,N_9699);
or U12449 (N_12449,N_8866,N_7681);
nand U12450 (N_12450,N_9320,N_9077);
nand U12451 (N_12451,N_9391,N_9210);
or U12452 (N_12452,N_8229,N_9722);
nand U12453 (N_12453,N_8450,N_9309);
and U12454 (N_12454,N_8661,N_8421);
xnor U12455 (N_12455,N_9279,N_9473);
nand U12456 (N_12456,N_7850,N_9640);
xnor U12457 (N_12457,N_9491,N_8714);
or U12458 (N_12458,N_9161,N_7823);
or U12459 (N_12459,N_8929,N_9545);
nand U12460 (N_12460,N_8538,N_9939);
nor U12461 (N_12461,N_8569,N_9536);
or U12462 (N_12462,N_7511,N_9429);
or U12463 (N_12463,N_8084,N_9709);
or U12464 (N_12464,N_8238,N_9784);
nand U12465 (N_12465,N_9546,N_8052);
nand U12466 (N_12466,N_8564,N_8684);
nand U12467 (N_12467,N_7675,N_7531);
nor U12468 (N_12468,N_8282,N_8827);
nor U12469 (N_12469,N_9330,N_7575);
or U12470 (N_12470,N_7825,N_8985);
nand U12471 (N_12471,N_8758,N_8485);
and U12472 (N_12472,N_9032,N_7553);
or U12473 (N_12473,N_8929,N_7541);
nand U12474 (N_12474,N_9356,N_9372);
and U12475 (N_12475,N_8845,N_7810);
nor U12476 (N_12476,N_9329,N_8064);
nor U12477 (N_12477,N_7710,N_7654);
xor U12478 (N_12478,N_9799,N_8891);
or U12479 (N_12479,N_9410,N_7695);
or U12480 (N_12480,N_8318,N_9675);
nor U12481 (N_12481,N_9448,N_7557);
or U12482 (N_12482,N_8814,N_8880);
and U12483 (N_12483,N_8723,N_9441);
and U12484 (N_12484,N_7648,N_9015);
nand U12485 (N_12485,N_8744,N_9503);
nor U12486 (N_12486,N_9200,N_7637);
nand U12487 (N_12487,N_9081,N_8529);
xnor U12488 (N_12488,N_8625,N_8720);
or U12489 (N_12489,N_9721,N_8081);
and U12490 (N_12490,N_9815,N_8616);
nand U12491 (N_12491,N_8802,N_9237);
and U12492 (N_12492,N_9712,N_7688);
or U12493 (N_12493,N_9285,N_8520);
xnor U12494 (N_12494,N_7774,N_9080);
nand U12495 (N_12495,N_7624,N_9450);
xor U12496 (N_12496,N_7504,N_9544);
or U12497 (N_12497,N_8178,N_9227);
or U12498 (N_12498,N_7591,N_7576);
xnor U12499 (N_12499,N_9943,N_8351);
nand U12500 (N_12500,N_10007,N_11186);
nor U12501 (N_12501,N_10788,N_11751);
xnor U12502 (N_12502,N_11307,N_11424);
or U12503 (N_12503,N_12166,N_11438);
and U12504 (N_12504,N_11855,N_12274);
xnor U12505 (N_12505,N_12457,N_10423);
or U12506 (N_12506,N_11390,N_10187);
xor U12507 (N_12507,N_11471,N_11052);
nand U12508 (N_12508,N_12219,N_10198);
nand U12509 (N_12509,N_11662,N_10195);
nand U12510 (N_12510,N_10605,N_10400);
and U12511 (N_12511,N_11548,N_11122);
nand U12512 (N_12512,N_11554,N_11739);
and U12513 (N_12513,N_10524,N_10740);
nand U12514 (N_12514,N_11126,N_11901);
or U12515 (N_12515,N_10263,N_11860);
and U12516 (N_12516,N_11789,N_11773);
or U12517 (N_12517,N_11892,N_11513);
nor U12518 (N_12518,N_11946,N_11346);
nor U12519 (N_12519,N_10657,N_10579);
nor U12520 (N_12520,N_12084,N_10927);
or U12521 (N_12521,N_11388,N_10877);
xnor U12522 (N_12522,N_10250,N_12351);
nor U12523 (N_12523,N_12299,N_10905);
nor U12524 (N_12524,N_10399,N_10582);
and U12525 (N_12525,N_10414,N_10247);
or U12526 (N_12526,N_11960,N_10826);
xor U12527 (N_12527,N_11366,N_10088);
nor U12528 (N_12528,N_11680,N_11454);
nand U12529 (N_12529,N_10833,N_12370);
xnor U12530 (N_12530,N_10120,N_11130);
nor U12531 (N_12531,N_12443,N_10189);
or U12532 (N_12532,N_10346,N_11357);
and U12533 (N_12533,N_12026,N_10327);
nor U12534 (N_12534,N_11531,N_10434);
nor U12535 (N_12535,N_10946,N_12101);
xor U12536 (N_12536,N_12319,N_12478);
or U12537 (N_12537,N_10589,N_10661);
xnor U12538 (N_12538,N_11313,N_12305);
or U12539 (N_12539,N_10167,N_10588);
and U12540 (N_12540,N_10968,N_11004);
or U12541 (N_12541,N_10259,N_10337);
or U12542 (N_12542,N_10306,N_11393);
xnor U12543 (N_12543,N_10026,N_10966);
and U12544 (N_12544,N_11279,N_11128);
xnor U12545 (N_12545,N_12364,N_12056);
xor U12546 (N_12546,N_10666,N_11633);
nand U12547 (N_12547,N_10301,N_11582);
and U12548 (N_12548,N_10769,N_10834);
nor U12549 (N_12549,N_10385,N_11895);
and U12550 (N_12550,N_12117,N_11087);
or U12551 (N_12551,N_11288,N_11578);
nand U12552 (N_12552,N_11885,N_10068);
nor U12553 (N_12553,N_12151,N_10479);
nor U12554 (N_12554,N_11194,N_10778);
nor U12555 (N_12555,N_11301,N_11422);
and U12556 (N_12556,N_11080,N_11841);
nand U12557 (N_12557,N_11423,N_12418);
or U12558 (N_12558,N_10892,N_10736);
nor U12559 (N_12559,N_10454,N_10133);
and U12560 (N_12560,N_10389,N_10768);
nand U12561 (N_12561,N_12204,N_12196);
and U12562 (N_12562,N_12013,N_10531);
or U12563 (N_12563,N_11172,N_10832);
xnor U12564 (N_12564,N_12498,N_12137);
xnor U12565 (N_12565,N_11356,N_11803);
nor U12566 (N_12566,N_10274,N_11026);
nand U12567 (N_12567,N_11312,N_10160);
nand U12568 (N_12568,N_12349,N_10997);
xor U12569 (N_12569,N_10475,N_10251);
or U12570 (N_12570,N_10271,N_10295);
xor U12571 (N_12571,N_10325,N_11107);
nand U12572 (N_12572,N_12255,N_10842);
xor U12573 (N_12573,N_11378,N_12469);
and U12574 (N_12574,N_10101,N_12023);
nor U12575 (N_12575,N_11403,N_10446);
or U12576 (N_12576,N_10302,N_11459);
nand U12577 (N_12577,N_10790,N_10585);
xnor U12578 (N_12578,N_12479,N_10720);
nor U12579 (N_12579,N_11408,N_11826);
nand U12580 (N_12580,N_10581,N_12165);
nor U12581 (N_12581,N_11854,N_11386);
and U12582 (N_12582,N_11251,N_10921);
nor U12583 (N_12583,N_10128,N_11639);
or U12584 (N_12584,N_12156,N_10759);
xor U12585 (N_12585,N_11266,N_10982);
nor U12586 (N_12586,N_10038,N_11023);
and U12587 (N_12587,N_10313,N_12053);
and U12588 (N_12588,N_10627,N_11838);
nor U12589 (N_12589,N_11853,N_10083);
and U12590 (N_12590,N_10872,N_10806);
xnor U12591 (N_12591,N_10859,N_10967);
or U12592 (N_12592,N_10548,N_12292);
nand U12593 (N_12593,N_10932,N_12231);
xor U12594 (N_12594,N_10122,N_12163);
nor U12595 (N_12595,N_10800,N_11289);
nand U12596 (N_12596,N_11064,N_11444);
nor U12597 (N_12597,N_11059,N_11482);
and U12598 (N_12598,N_11687,N_11652);
xnor U12599 (N_12599,N_10724,N_12400);
and U12600 (N_12600,N_11098,N_11238);
nand U12601 (N_12601,N_10489,N_10347);
xor U12602 (N_12602,N_10836,N_11961);
or U12603 (N_12603,N_11956,N_12143);
and U12604 (N_12604,N_11807,N_11399);
or U12605 (N_12605,N_11074,N_11906);
or U12606 (N_12606,N_12437,N_11959);
or U12607 (N_12607,N_11463,N_11686);
or U12608 (N_12608,N_11001,N_11040);
xor U12609 (N_12609,N_12040,N_10474);
and U12610 (N_12610,N_10119,N_11630);
xnor U12611 (N_12611,N_10121,N_10591);
nor U12612 (N_12612,N_12359,N_10344);
or U12613 (N_12613,N_11611,N_12054);
and U12614 (N_12614,N_12035,N_12241);
and U12615 (N_12615,N_11066,N_11569);
xor U12616 (N_12616,N_11748,N_12366);
nand U12617 (N_12617,N_11450,N_10342);
nor U12618 (N_12618,N_11006,N_11614);
xor U12619 (N_12619,N_12417,N_12218);
and U12620 (N_12620,N_11371,N_12394);
and U12621 (N_12621,N_10017,N_10248);
or U12622 (N_12622,N_11617,N_11310);
nor U12623 (N_12623,N_11579,N_11615);
xor U12624 (N_12624,N_12230,N_12111);
xnor U12625 (N_12625,N_11747,N_11110);
xnor U12626 (N_12626,N_12452,N_12461);
nand U12627 (N_12627,N_10380,N_12289);
nor U12628 (N_12628,N_11760,N_11114);
nand U12629 (N_12629,N_12310,N_11705);
or U12630 (N_12630,N_11264,N_12285);
xor U12631 (N_12631,N_11129,N_10178);
xnor U12632 (N_12632,N_10291,N_12181);
nor U12633 (N_12633,N_10062,N_11102);
xnor U12634 (N_12634,N_12318,N_12290);
nor U12635 (N_12635,N_10654,N_11836);
or U12636 (N_12636,N_10047,N_10791);
nor U12637 (N_12637,N_11037,N_12159);
and U12638 (N_12638,N_10883,N_10359);
nand U12639 (N_12639,N_11239,N_10223);
xnor U12640 (N_12640,N_10786,N_11494);
nor U12641 (N_12641,N_11862,N_10757);
nand U12642 (N_12642,N_11411,N_11175);
nor U12643 (N_12643,N_11586,N_11512);
and U12644 (N_12644,N_11592,N_11690);
and U12645 (N_12645,N_11036,N_11360);
xor U12646 (N_12646,N_11204,N_10236);
xor U12647 (N_12647,N_10435,N_12264);
xnor U12648 (N_12648,N_11635,N_10050);
and U12649 (N_12649,N_10387,N_12293);
or U12650 (N_12650,N_12254,N_12427);
nor U12651 (N_12651,N_11088,N_11092);
nand U12652 (N_12652,N_12209,N_12182);
or U12653 (N_12653,N_10429,N_12295);
xnor U12654 (N_12654,N_11456,N_11453);
and U12655 (N_12655,N_12393,N_11071);
and U12656 (N_12656,N_10484,N_12078);
or U12657 (N_12657,N_10099,N_11035);
and U12658 (N_12658,N_12051,N_11299);
and U12659 (N_12659,N_10199,N_10957);
xnor U12660 (N_12660,N_10881,N_10290);
nand U12661 (N_12661,N_10461,N_12010);
nor U12662 (N_12662,N_10087,N_12031);
nand U12663 (N_12663,N_11764,N_10360);
nor U12664 (N_12664,N_10221,N_10526);
nor U12665 (N_12665,N_10981,N_10143);
xnor U12666 (N_12666,N_11246,N_12385);
nand U12667 (N_12667,N_10234,N_10563);
xor U12668 (N_12668,N_11947,N_10642);
nand U12669 (N_12669,N_10130,N_11332);
xnor U12670 (N_12670,N_11145,N_10293);
nand U12671 (N_12671,N_10055,N_12388);
nand U12672 (N_12672,N_12017,N_11234);
nand U12673 (N_12673,N_12138,N_10470);
and U12674 (N_12674,N_12186,N_10712);
nor U12675 (N_12675,N_11044,N_11774);
or U12676 (N_12676,N_12201,N_11989);
xnor U12677 (N_12677,N_12162,N_10862);
nand U12678 (N_12678,N_11945,N_10555);
nand U12679 (N_12679,N_12025,N_11762);
and U12680 (N_12680,N_11149,N_10752);
nor U12681 (N_12681,N_11277,N_11201);
xnor U12682 (N_12682,N_11955,N_12036);
nor U12683 (N_12683,N_11089,N_11858);
nor U12684 (N_12684,N_11560,N_10770);
and U12685 (N_12685,N_10540,N_11840);
and U12686 (N_12686,N_11417,N_11708);
and U12687 (N_12687,N_10730,N_10218);
nand U12688 (N_12688,N_12337,N_12381);
and U12689 (N_12689,N_11118,N_10255);
nor U12690 (N_12690,N_10108,N_12046);
and U12691 (N_12691,N_11124,N_12249);
or U12692 (N_12692,N_10443,N_10084);
nor U12693 (N_12693,N_11030,N_10970);
xor U12694 (N_12694,N_11191,N_10878);
or U12695 (N_12695,N_11406,N_10985);
nor U12696 (N_12696,N_10940,N_12161);
and U12697 (N_12697,N_11551,N_10317);
and U12698 (N_12698,N_10956,N_10487);
and U12699 (N_12699,N_11768,N_11663);
nor U12700 (N_12700,N_12014,N_11908);
nor U12701 (N_12701,N_11187,N_10018);
and U12702 (N_12702,N_10969,N_12379);
nor U12703 (N_12703,N_11100,N_12077);
or U12704 (N_12704,N_10508,N_10311);
nand U12705 (N_12705,N_10809,N_10145);
xnor U12706 (N_12706,N_11488,N_11013);
or U12707 (N_12707,N_10609,N_11738);
and U12708 (N_12708,N_11500,N_10362);
and U12709 (N_12709,N_11568,N_11309);
nand U12710 (N_12710,N_11799,N_10460);
xor U12711 (N_12711,N_12407,N_10869);
xor U12712 (N_12712,N_11625,N_11948);
nand U12713 (N_12713,N_10185,N_11090);
nor U12714 (N_12714,N_10449,N_10158);
nor U12715 (N_12715,N_12405,N_11469);
nand U12716 (N_12716,N_11156,N_12043);
nand U12717 (N_12717,N_10888,N_10624);
and U12718 (N_12718,N_12470,N_11075);
or U12719 (N_12719,N_11584,N_10655);
and U12720 (N_12720,N_11606,N_10534);
or U12721 (N_12721,N_12211,N_10278);
and U12722 (N_12722,N_10267,N_12376);
or U12723 (N_12723,N_11376,N_10012);
and U12724 (N_12724,N_11015,N_11628);
xor U12725 (N_12725,N_12496,N_12140);
and U12726 (N_12726,N_12399,N_10637);
and U12727 (N_12727,N_10377,N_10530);
or U12728 (N_12728,N_10929,N_11334);
or U12729 (N_12729,N_10965,N_11632);
nand U12730 (N_12730,N_12173,N_10544);
nor U12731 (N_12731,N_11601,N_11538);
xnor U12732 (N_12732,N_10639,N_10758);
xor U12733 (N_12733,N_10726,N_10407);
nor U12734 (N_12734,N_12476,N_11924);
nand U12735 (N_12735,N_10804,N_12065);
and U12736 (N_12736,N_12474,N_10008);
nor U12737 (N_12737,N_11268,N_11389);
or U12738 (N_12738,N_11340,N_12224);
or U12739 (N_12739,N_10920,N_10139);
nor U12740 (N_12740,N_12093,N_11884);
xnor U12741 (N_12741,N_11249,N_11027);
and U12742 (N_12742,N_12180,N_11957);
nand U12743 (N_12743,N_11867,N_12425);
xnor U12744 (N_12744,N_11783,N_10751);
nor U12745 (N_12745,N_11910,N_12451);
nor U12746 (N_12746,N_10095,N_12118);
nand U12747 (N_12747,N_12397,N_11281);
and U12748 (N_12748,N_10252,N_10977);
and U12749 (N_12749,N_10628,N_10871);
xor U12750 (N_12750,N_10527,N_12480);
xor U12751 (N_12751,N_10256,N_12263);
nand U12752 (N_12752,N_10496,N_10091);
nand U12753 (N_12753,N_10636,N_10989);
nand U12754 (N_12754,N_11295,N_10704);
xnor U12755 (N_12755,N_11969,N_11219);
and U12756 (N_12756,N_10687,N_11881);
nor U12757 (N_12757,N_11121,N_10276);
nand U12758 (N_12758,N_11458,N_10885);
and U12759 (N_12759,N_11303,N_11882);
or U12760 (N_12760,N_11155,N_11396);
nand U12761 (N_12761,N_10264,N_12448);
xor U12762 (N_12762,N_10607,N_12052);
and U12763 (N_12763,N_11692,N_12481);
xor U12764 (N_12764,N_11688,N_10756);
nor U12765 (N_12765,N_10701,N_12416);
nand U12766 (N_12766,N_10512,N_12340);
xor U12767 (N_12767,N_12175,N_11041);
and U12768 (N_12768,N_11518,N_12298);
nand U12769 (N_12769,N_10580,N_12383);
nor U12770 (N_12770,N_11527,N_11963);
nand U12771 (N_12771,N_11224,N_10115);
nor U12772 (N_12772,N_10835,N_12123);
xor U12773 (N_12773,N_11880,N_11174);
and U12774 (N_12774,N_10378,N_11368);
xor U12775 (N_12775,N_12042,N_10963);
nor U12776 (N_12776,N_10695,N_10780);
or U12777 (N_12777,N_11819,N_10292);
and U12778 (N_12778,N_11998,N_11173);
nor U12779 (N_12779,N_10324,N_10598);
and U12780 (N_12780,N_10352,N_10254);
nor U12781 (N_12781,N_10974,N_12371);
xor U12782 (N_12782,N_11225,N_11432);
nand U12783 (N_12783,N_12357,N_10914);
and U12784 (N_12784,N_11651,N_11917);
nor U12785 (N_12785,N_12253,N_10450);
nand U12786 (N_12786,N_12311,N_10764);
and U12787 (N_12787,N_11631,N_12495);
xnor U12788 (N_12788,N_12092,N_10688);
or U12789 (N_12789,N_11811,N_10995);
and U12790 (N_12790,N_11232,N_10357);
xor U12791 (N_12791,N_11675,N_10441);
or U12792 (N_12792,N_12472,N_10622);
nand U12793 (N_12793,N_12436,N_11053);
xnor U12794 (N_12794,N_10909,N_12170);
nand U12795 (N_12795,N_12287,N_11550);
or U12796 (N_12796,N_10147,N_10610);
nor U12797 (N_12797,N_10789,N_11929);
nand U12798 (N_12798,N_11095,N_11328);
xnor U12799 (N_12799,N_11532,N_10922);
or U12800 (N_12800,N_12473,N_11868);
nor U12801 (N_12801,N_11039,N_11434);
nand U12802 (N_12802,N_12200,N_11865);
xor U12803 (N_12803,N_11123,N_11361);
and U12804 (N_12804,N_12217,N_10287);
or U12805 (N_12805,N_11655,N_10427);
nor U12806 (N_12806,N_10558,N_10795);
xor U12807 (N_12807,N_10054,N_12426);
and U12808 (N_12808,N_10950,N_10802);
nor U12809 (N_12809,N_11978,N_11805);
nand U12810 (N_12810,N_10100,N_11641);
xnor U12811 (N_12811,N_12235,N_10358);
nand U12812 (N_12812,N_11698,N_12061);
or U12813 (N_12813,N_12157,N_11427);
nor U12814 (N_12814,N_10281,N_11715);
or U12815 (N_12815,N_12435,N_11079);
and U12816 (N_12816,N_12185,N_12491);
nor U12817 (N_12817,N_11380,N_10113);
nand U12818 (N_12818,N_10741,N_12072);
or U12819 (N_12819,N_11517,N_11391);
and U12820 (N_12820,N_11971,N_10210);
and U12821 (N_12821,N_12361,N_11869);
or U12822 (N_12822,N_12341,N_11503);
xor U12823 (N_12823,N_10801,N_11740);
xnor U12824 (N_12824,N_11545,N_11852);
nand U12825 (N_12825,N_10188,N_11117);
nor U12826 (N_12826,N_12389,N_11888);
and U12827 (N_12827,N_10825,N_10253);
and U12828 (N_12828,N_11324,N_10201);
nor U12829 (N_12829,N_11374,N_11185);
and U12830 (N_12830,N_10338,N_11681);
or U12831 (N_12831,N_10107,N_12355);
nand U12832 (N_12832,N_12074,N_12281);
or U12833 (N_12833,N_10529,N_11283);
xnor U12834 (N_12834,N_10608,N_11804);
or U12835 (N_12835,N_10953,N_11778);
nor U12836 (N_12836,N_11139,N_10009);
nand U12837 (N_12837,N_11684,N_10612);
xnor U12838 (N_12838,N_10493,N_10296);
xor U12839 (N_12839,N_12304,N_11083);
nor U12840 (N_12840,N_10678,N_10345);
nor U12841 (N_12841,N_12432,N_11497);
nand U12842 (N_12842,N_10803,N_12213);
nand U12843 (N_12843,N_12222,N_10984);
nor U12844 (N_12844,N_10964,N_11430);
nand U12845 (N_12845,N_10240,N_11097);
or U12846 (N_12846,N_10320,N_11877);
xor U12847 (N_12847,N_12490,N_11610);
xor U12848 (N_12848,N_11997,N_10978);
and U12849 (N_12849,N_10163,N_11700);
and U12850 (N_12850,N_12420,N_12107);
or U12851 (N_12851,N_11954,N_10551);
nand U12852 (N_12852,N_11190,N_12167);
or U12853 (N_12853,N_10299,N_11580);
nor U12854 (N_12854,N_12234,N_11942);
and U12855 (N_12855,N_12477,N_10282);
xnor U12856 (N_12856,N_11790,N_10438);
and U12857 (N_12857,N_10601,N_11984);
or U12858 (N_12858,N_10469,N_11563);
xor U12859 (N_12859,N_11810,N_11542);
and U12860 (N_12860,N_11546,N_10615);
or U12861 (N_12861,N_12353,N_11833);
or U12862 (N_12862,N_11253,N_11570);
nor U12863 (N_12863,N_10224,N_11609);
or U12864 (N_12864,N_11055,N_10595);
nand U12865 (N_12865,N_10517,N_11195);
and U12866 (N_12866,N_12326,N_12021);
or U12867 (N_12867,N_11189,N_10890);
xnor U12868 (N_12868,N_11069,N_11333);
or U12869 (N_12869,N_11757,N_11321);
or U12870 (N_12870,N_10785,N_11337);
nor U12871 (N_12871,N_12335,N_11448);
nand U12872 (N_12872,N_10379,N_12243);
and U12873 (N_12873,N_11769,N_12037);
and U12874 (N_12874,N_10706,N_10599);
nand U12875 (N_12875,N_11891,N_10072);
or U12876 (N_12876,N_11649,N_12467);
or U12877 (N_12877,N_11086,N_11874);
and U12878 (N_12878,N_12450,N_10542);
xor U12879 (N_12879,N_11802,N_11590);
nand U12880 (N_12880,N_10403,N_12019);
or U12881 (N_12881,N_12286,N_10866);
nand U12882 (N_12882,N_10354,N_10369);
xor U12883 (N_12883,N_10754,N_10716);
or U12884 (N_12884,N_12041,N_12282);
xnor U12885 (N_12885,N_12422,N_10048);
or U12886 (N_12886,N_12060,N_11723);
and U12887 (N_12887,N_10880,N_10215);
nand U12888 (N_12888,N_11750,N_11850);
nor U12889 (N_12889,N_11153,N_10341);
xor U12890 (N_12890,N_12483,N_11857);
and U12891 (N_12891,N_11166,N_11808);
nand U12892 (N_12892,N_11017,N_10904);
nand U12893 (N_12893,N_11327,N_10284);
and U12894 (N_12894,N_12328,N_12176);
nand U12895 (N_12895,N_11367,N_10478);
or U12896 (N_12896,N_11325,N_11094);
xor U12897 (N_12897,N_11046,N_11377);
nor U12898 (N_12898,N_12252,N_11033);
and U12899 (N_12899,N_11207,N_10175);
and U12900 (N_12900,N_10670,N_10040);
nor U12901 (N_12901,N_10660,N_10053);
xor U12902 (N_12902,N_11477,N_12245);
nand U12903 (N_12903,N_12172,N_10578);
and U12904 (N_12904,N_10902,N_10089);
nor U12905 (N_12905,N_10186,N_10954);
xor U12906 (N_12906,N_10822,N_10014);
and U12907 (N_12907,N_11620,N_10584);
xor U12908 (N_12908,N_11177,N_11714);
or U12909 (N_12909,N_10694,N_10235);
xor U12910 (N_12910,N_10691,N_11395);
xnor U12911 (N_12911,N_12102,N_10041);
nand U12912 (N_12912,N_12272,N_11668);
and U12913 (N_12913,N_12131,N_10465);
and U12914 (N_12914,N_11976,N_11983);
xnor U12915 (N_12915,N_10838,N_11161);
and U12916 (N_12916,N_11659,N_10674);
xor U12917 (N_12917,N_11029,N_10705);
nor U12918 (N_12918,N_10260,N_11435);
or U12919 (N_12919,N_10721,N_10958);
nand U12920 (N_12920,N_11719,N_11467);
or U12921 (N_12921,N_12112,N_11958);
xor U12922 (N_12922,N_12446,N_12334);
xor U12923 (N_12923,N_11878,N_11515);
nand U12924 (N_12924,N_11180,N_10368);
or U12925 (N_12925,N_11392,N_12312);
or U12926 (N_12926,N_10028,N_10168);
and U12927 (N_12927,N_10525,N_11661);
nand U12928 (N_12928,N_10515,N_12346);
nor U12929 (N_12929,N_11599,N_11058);
or U12930 (N_12930,N_11887,N_12221);
or U12931 (N_12931,N_10837,N_12086);
nor U12932 (N_12932,N_12369,N_11082);
nor U12933 (N_12933,N_10374,N_11685);
and U12934 (N_12934,N_10870,N_12171);
and U12935 (N_12935,N_10351,N_11144);
and U12936 (N_12936,N_12007,N_12266);
nor U12937 (N_12937,N_10522,N_12459);
and U12938 (N_12938,N_10340,N_12352);
or U12939 (N_12939,N_12475,N_11975);
xor U12940 (N_12940,N_11428,N_11441);
nand U12941 (N_12941,N_11486,N_12442);
or U12942 (N_12942,N_11644,N_10209);
nand U12943 (N_12943,N_11056,N_10568);
nand U12944 (N_12944,N_10861,N_10696);
nand U12945 (N_12945,N_12148,N_10629);
xnor U12946 (N_12946,N_10532,N_11593);
or U12947 (N_12947,N_12142,N_10169);
nand U12948 (N_12948,N_10082,N_12278);
and U12949 (N_12949,N_12147,N_11616);
or U12950 (N_12950,N_10882,N_12244);
xnor U12951 (N_12951,N_11188,N_11717);
xnor U12952 (N_12952,N_10002,N_10390);
nor U12953 (N_12953,N_10738,N_10973);
and U12954 (N_12954,N_12073,N_11991);
nand U12955 (N_12955,N_10850,N_10535);
nor U12956 (N_12956,N_11148,N_10875);
nor U12957 (N_12957,N_10876,N_10216);
or U12958 (N_12958,N_10986,N_11049);
and U12959 (N_12959,N_11168,N_10572);
nand U12960 (N_12960,N_10440,N_11111);
nor U12961 (N_12961,N_11743,N_10899);
nor U12962 (N_12962,N_11311,N_11861);
and U12963 (N_12963,N_10110,N_12485);
or U12964 (N_12964,N_11536,N_10635);
or U12965 (N_12965,N_11873,N_10396);
or U12966 (N_12966,N_10242,N_10370);
and U12967 (N_12967,N_12223,N_10466);
nor U12968 (N_12968,N_11091,N_11382);
or U12969 (N_12969,N_12133,N_11243);
nor U12970 (N_12970,N_11231,N_10990);
xnor U12971 (N_12971,N_10680,N_11523);
xor U12972 (N_12972,N_11605,N_12152);
nor U12973 (N_12973,N_11795,N_11741);
nand U12974 (N_12974,N_11561,N_11256);
nand U12975 (N_12975,N_10777,N_10630);
or U12976 (N_12976,N_12199,N_11970);
nor U12977 (N_12977,N_10463,N_12232);
nor U12978 (N_12978,N_11559,N_10560);
or U12979 (N_12979,N_11839,N_10024);
and U12980 (N_12980,N_11255,N_10105);
and U12981 (N_12981,N_11784,N_10428);
nand U12982 (N_12982,N_11047,N_11372);
xor U12983 (N_12983,N_11541,N_10810);
or U12984 (N_12984,N_10505,N_12374);
nor U12985 (N_12985,N_11673,N_11431);
xor U12986 (N_12986,N_12090,N_11950);
or U12987 (N_12987,N_10845,N_11414);
nor U12988 (N_12988,N_12308,N_10782);
nand U12989 (N_12989,N_12158,N_11791);
nor U12990 (N_12990,N_11544,N_10137);
nor U12991 (N_12991,N_12115,N_11786);
and U12992 (N_12992,N_10853,N_11216);
nand U12993 (N_12993,N_10180,N_11856);
xor U12994 (N_12994,N_10910,N_12297);
and U12995 (N_12995,N_11755,N_10184);
nand U12996 (N_12996,N_12039,N_11761);
or U12997 (N_12997,N_11703,N_11205);
xnor U12998 (N_12998,N_10148,N_11939);
and U12999 (N_12999,N_11654,N_11835);
nand U13000 (N_13000,N_10413,N_10005);
xnor U13001 (N_13001,N_10994,N_11247);
or U13002 (N_13002,N_10992,N_11412);
nor U13003 (N_13003,N_10732,N_10926);
nand U13004 (N_13004,N_12391,N_11398);
and U13005 (N_13005,N_11511,N_10776);
or U13006 (N_13006,N_11109,N_11355);
or U13007 (N_13007,N_10857,N_11996);
nand U13008 (N_13008,N_11101,N_11733);
xor U13009 (N_13009,N_10506,N_10065);
xor U13010 (N_13010,N_11830,N_10503);
xnor U13011 (N_13011,N_11447,N_12070);
xnor U13012 (N_13012,N_11481,N_12484);
or U13013 (N_13013,N_12248,N_10270);
or U13014 (N_13014,N_11846,N_11042);
and U13015 (N_13015,N_11208,N_11782);
nor U13016 (N_13016,N_12120,N_10207);
or U13017 (N_13017,N_12434,N_11728);
or U13018 (N_13018,N_10931,N_10388);
and U13019 (N_13019,N_10722,N_10381);
or U13020 (N_13020,N_10520,N_11018);
nand U13021 (N_13021,N_10150,N_12225);
xor U13022 (N_13022,N_12493,N_10052);
nor U13023 (N_13023,N_11455,N_12382);
xor U13024 (N_13024,N_11930,N_10852);
xnor U13025 (N_13025,N_12114,N_11163);
and U13026 (N_13026,N_11445,N_11812);
nor U13027 (N_13027,N_11549,N_12377);
and U13028 (N_13028,N_10979,N_10102);
or U13029 (N_13029,N_11016,N_11057);
or U13030 (N_13030,N_11009,N_11300);
nand U13031 (N_13031,N_11753,N_11449);
xnor U13032 (N_13032,N_11522,N_11749);
nand U13033 (N_13033,N_11952,N_10363);
or U13034 (N_13034,N_11540,N_10739);
nand U13035 (N_13035,N_11359,N_11151);
nand U13036 (N_13036,N_11461,N_10060);
nor U13037 (N_13037,N_10562,N_10049);
or U13038 (N_13038,N_11076,N_11509);
or U13039 (N_13039,N_10718,N_11660);
or U13040 (N_13040,N_10001,N_10708);
and U13041 (N_13041,N_10590,N_10439);
nand U13042 (N_13042,N_11716,N_10571);
nor U13043 (N_13043,N_12464,N_12089);
and U13044 (N_13044,N_10152,N_11524);
and U13045 (N_13045,N_10815,N_10498);
nand U13046 (N_13046,N_10889,N_11282);
xnor U13047 (N_13047,N_10417,N_10907);
or U13048 (N_13048,N_10860,N_10509);
nor U13049 (N_13049,N_12002,N_10261);
nor U13050 (N_13050,N_11972,N_12020);
nand U13051 (N_13051,N_10194,N_11214);
and U13052 (N_13052,N_10576,N_11604);
nor U13053 (N_13053,N_12113,N_10561);
and U13054 (N_13054,N_11520,N_10649);
xor U13055 (N_13055,N_12375,N_12329);
nor U13056 (N_13056,N_10425,N_10677);
xnor U13057 (N_13057,N_10021,N_11045);
or U13058 (N_13058,N_10539,N_10165);
xnor U13059 (N_13059,N_11702,N_12082);
or U13060 (N_13060,N_10366,N_11154);
nor U13061 (N_13061,N_10081,N_11510);
xor U13062 (N_13062,N_10142,N_12256);
nor U13063 (N_13063,N_12058,N_11112);
xor U13064 (N_13064,N_12205,N_11815);
nand U13065 (N_13065,N_11127,N_12402);
xnor U13066 (N_13066,N_11480,N_11038);
or U13067 (N_13067,N_10076,N_10510);
nor U13068 (N_13068,N_11171,N_10546);
xnor U13069 (N_13069,N_11387,N_11667);
nor U13070 (N_13070,N_11160,N_10015);
xor U13071 (N_13071,N_10945,N_10027);
nand U13072 (N_13072,N_11931,N_10376);
nor U13073 (N_13073,N_11727,N_10383);
nand U13074 (N_13074,N_11823,N_12273);
nor U13075 (N_13075,N_11407,N_10225);
xnor U13076 (N_13076,N_10442,N_11451);
nor U13077 (N_13077,N_10821,N_12108);
nor U13078 (N_13078,N_11893,N_11566);
and U13079 (N_13079,N_11227,N_10536);
nand U13080 (N_13080,N_11936,N_11270);
nand U13081 (N_13081,N_10901,N_10737);
nand U13082 (N_13082,N_12421,N_10771);
nand U13083 (N_13083,N_12076,N_10886);
nand U13084 (N_13084,N_12067,N_10538);
nand U13085 (N_13085,N_12198,N_10200);
or U13086 (N_13086,N_10071,N_10051);
or U13087 (N_13087,N_11697,N_12195);
nor U13088 (N_13088,N_11974,N_10204);
nor U13089 (N_13089,N_10314,N_10318);
nor U13090 (N_13090,N_11212,N_12438);
nand U13091 (N_13091,N_12368,N_10693);
xor U13092 (N_13092,N_12424,N_10455);
nand U13093 (N_13093,N_11331,N_10734);
or U13094 (N_13094,N_11263,N_11354);
nor U13095 (N_13095,N_10723,N_12358);
xnor U13096 (N_13096,N_11794,N_11696);
nor U13097 (N_13097,N_12261,N_11221);
nor U13098 (N_13098,N_11294,N_11063);
and U13099 (N_13099,N_11982,N_11233);
nand U13100 (N_13100,N_10300,N_12307);
nor U13101 (N_13101,N_10840,N_12343);
xnor U13102 (N_13102,N_11831,N_11257);
and U13103 (N_13103,N_10066,N_12411);
and U13104 (N_13104,N_11647,N_10944);
nand U13105 (N_13105,N_11870,N_12099);
xor U13106 (N_13106,N_11199,N_11521);
and U13107 (N_13107,N_12033,N_10507);
or U13108 (N_13108,N_11514,N_10781);
and U13109 (N_13109,N_10213,N_10653);
and U13110 (N_13110,N_10552,N_11636);
or U13111 (N_13111,N_10500,N_11024);
nand U13112 (N_13112,N_12395,N_11608);
and U13113 (N_13113,N_11665,N_10433);
nor U13114 (N_13114,N_10208,N_10939);
nand U13115 (N_13115,N_10025,N_12348);
nand U13116 (N_13116,N_10171,N_11993);
and U13117 (N_13117,N_12242,N_10398);
xnor U13118 (N_13118,N_10013,N_11650);
nand U13119 (N_13119,N_10710,N_10634);
xnor U13120 (N_13120,N_11344,N_11588);
nand U13121 (N_13121,N_11973,N_11923);
and U13122 (N_13122,N_11261,N_10230);
and U13123 (N_13123,N_11275,N_12237);
xor U13124 (N_13124,N_11701,N_11581);
nand U13125 (N_13125,N_10792,N_12022);
xor U13126 (N_13126,N_11022,N_12440);
or U13127 (N_13127,N_11285,N_11922);
and U13128 (N_13128,N_11134,N_10772);
or U13129 (N_13129,N_10323,N_10042);
nor U13130 (N_13130,N_12468,N_10633);
or U13131 (N_13131,N_11011,N_10495);
and U13132 (N_13132,N_11081,N_10893);
or U13133 (N_13133,N_11265,N_10212);
nand U13134 (N_13134,N_10268,N_11785);
and U13135 (N_13135,N_11162,N_11280);
nand U13136 (N_13136,N_11600,N_11215);
and U13137 (N_13137,N_11505,N_10416);
xnor U13138 (N_13138,N_10067,N_10231);
xor U13139 (N_13139,N_11426,N_11140);
and U13140 (N_13140,N_11742,N_10382);
nor U13141 (N_13141,N_10728,N_11345);
nor U13142 (N_13142,N_11875,N_12069);
and U13143 (N_13143,N_11746,N_11832);
and U13144 (N_13144,N_10233,N_10279);
and U13145 (N_13145,N_11914,N_10090);
nor U13146 (N_13146,N_10085,N_11051);
xnor U13147 (N_13147,N_11383,N_10011);
or U13148 (N_13148,N_12153,N_10448);
nor U13149 (N_13149,N_10126,N_11597);
xor U13150 (N_13150,N_11602,N_11756);
xnor U13151 (N_13151,N_10063,N_10326);
xnor U13152 (N_13152,N_11478,N_10330);
nor U13153 (N_13153,N_11896,N_10597);
nor U13154 (N_13154,N_10074,N_12063);
xor U13155 (N_13155,N_11000,N_10333);
or U13156 (N_13156,N_12270,N_10412);
nor U13157 (N_13157,N_11131,N_11779);
nand U13158 (N_13158,N_12338,N_10851);
nand U13159 (N_13159,N_11788,N_11664);
and U13160 (N_13160,N_10858,N_10136);
nor U13161 (N_13161,N_12210,N_12049);
xnor U13162 (N_13162,N_10131,N_11859);
xor U13163 (N_13163,N_11193,N_10916);
and U13164 (N_13164,N_11889,N_11902);
xnor U13165 (N_13165,N_11462,N_12106);
nor U13166 (N_13166,N_12497,N_10229);
or U13167 (N_13167,N_12229,N_10034);
nor U13168 (N_13168,N_12071,N_11907);
or U13169 (N_13169,N_10672,N_10915);
nand U13170 (N_13170,N_11607,N_10000);
nor U13171 (N_13171,N_11990,N_11470);
nand U13172 (N_13172,N_10683,N_11898);
nand U13173 (N_13173,N_11104,N_10371);
and U13174 (N_13174,N_10426,N_10887);
or U13175 (N_13175,N_10232,N_11731);
xor U13176 (N_13176,N_10227,N_10557);
and U13177 (N_13177,N_10733,N_10488);
nor U13178 (N_13178,N_11646,N_10632);
nand U13179 (N_13179,N_10164,N_10686);
and U13180 (N_13180,N_12404,N_10436);
or U13181 (N_13181,N_11484,N_11329);
and U13182 (N_13182,N_10865,N_10692);
or U13183 (N_13183,N_12098,N_11125);
or U13184 (N_13184,N_10127,N_11585);
or U13185 (N_13185,N_10244,N_11565);
and U13186 (N_13186,N_11485,N_10149);
xor U13187 (N_13187,N_10698,N_10983);
nand U13188 (N_13188,N_10375,N_11988);
and U13189 (N_13189,N_10742,N_10820);
or U13190 (N_13190,N_11864,N_11465);
nand U13191 (N_13191,N_11416,N_11113);
xnor U13192 (N_13192,N_10663,N_11925);
nand U13193 (N_13193,N_11085,N_10166);
nor U13194 (N_13194,N_12460,N_11932);
nand U13195 (N_13195,N_12197,N_11273);
nor U13196 (N_13196,N_11828,N_11994);
and U13197 (N_13197,N_12189,N_10243);
xor U13198 (N_13198,N_10174,N_11381);
xnor U13199 (N_13199,N_10991,N_11433);
xnor U13200 (N_13200,N_11365,N_11583);
and U13201 (N_13201,N_11206,N_11916);
nand U13202 (N_13202,N_11209,N_10746);
nand U13203 (N_13203,N_12095,N_10135);
or U13204 (N_13204,N_10714,N_11567);
nand U13205 (N_13205,N_11508,N_10298);
and U13206 (N_13206,N_10613,N_11315);
and U13207 (N_13207,N_10125,N_12414);
nand U13208 (N_13208,N_10335,N_11676);
and U13209 (N_13209,N_10594,N_12045);
nand U13210 (N_13210,N_11226,N_12322);
and U13211 (N_13211,N_12300,N_10482);
or U13212 (N_13212,N_12233,N_10702);
nor U13213 (N_13213,N_11547,N_10154);
nor U13214 (N_13214,N_10205,N_11474);
xnor U13215 (N_13215,N_12431,N_11787);
and U13216 (N_13216,N_12350,N_11629);
xor U13217 (N_13217,N_11351,N_11218);
nor U13218 (N_13218,N_12463,N_10277);
or U13219 (N_13219,N_11780,N_11073);
xor U13220 (N_13220,N_10863,N_11845);
or U13221 (N_13221,N_11236,N_11736);
and U13222 (N_13222,N_12239,N_10808);
xor U13223 (N_13223,N_10193,N_12193);
xor U13224 (N_13224,N_12184,N_10421);
nand U13225 (N_13225,N_12083,N_11577);
nor U13226 (N_13226,N_10492,N_10156);
xor U13227 (N_13227,N_10092,N_10938);
xor U13228 (N_13228,N_10394,N_11777);
or U13229 (N_13229,N_11405,N_12064);
nor U13230 (N_13230,N_10671,N_11370);
or U13231 (N_13231,N_11834,N_10491);
nand U13232 (N_13232,N_10499,N_11694);
nor U13233 (N_13233,N_11169,N_10554);
xor U13234 (N_13234,N_12342,N_10673);
nand U13235 (N_13235,N_11574,N_12226);
and U13236 (N_13236,N_11718,N_12081);
and U13237 (N_13237,N_11872,N_10350);
xnor U13238 (N_13238,N_10976,N_12354);
xnor U13239 (N_13239,N_12408,N_12302);
or U13240 (N_13240,N_11178,N_10685);
or U13241 (N_13241,N_11883,N_11305);
and U13242 (N_13242,N_12325,N_11297);
or U13243 (N_13243,N_10502,N_12214);
or U13244 (N_13244,N_10019,N_11707);
nand U13245 (N_13245,N_10395,N_11648);
xnor U13246 (N_13246,N_11339,N_10124);
nor U13247 (N_13247,N_11420,N_11375);
xnor U13248 (N_13248,N_12179,N_11670);
and U13249 (N_13249,N_11589,N_12356);
or U13250 (N_13250,N_10807,N_10811);
or U13251 (N_13251,N_10864,N_10078);
and U13252 (N_13252,N_12367,N_10519);
or U13253 (N_13253,N_10715,N_11242);
or U13254 (N_13254,N_12127,N_11133);
and U13255 (N_13255,N_12456,N_12303);
or U13256 (N_13256,N_10823,N_11072);
nand U13257 (N_13257,N_11235,N_10747);
nor U13258 (N_13258,N_12317,N_12441);
and U13259 (N_13259,N_10182,N_10550);
xnor U13260 (N_13260,N_10727,N_10308);
or U13261 (N_13261,N_11116,N_10134);
nand U13262 (N_13262,N_11772,N_12145);
nand U13263 (N_13263,N_11248,N_10748);
and U13264 (N_13264,N_10043,N_11060);
or U13265 (N_13265,N_11899,N_12339);
or U13266 (N_13266,N_10942,N_10104);
nor U13267 (N_13267,N_11240,N_11489);
xor U13268 (N_13268,N_10817,N_11847);
xnor U13269 (N_13269,N_10444,N_11062);
xor U13270 (N_13270,N_10729,N_10356);
nor U13271 (N_13271,N_11781,N_12250);
and U13272 (N_13272,N_12315,N_11418);
xnor U13273 (N_13273,N_10056,N_12396);
or U13274 (N_13274,N_11320,N_11526);
xnor U13275 (N_13275,N_11276,N_12194);
nand U13276 (N_13276,N_11758,N_11941);
nor U13277 (N_13277,N_12212,N_10574);
or U13278 (N_13278,N_12372,N_10873);
and U13279 (N_13279,N_10980,N_10528);
nand U13280 (N_13280,N_11622,N_11135);
and U13281 (N_13281,N_10310,N_10410);
xor U13282 (N_13282,N_12149,N_11197);
xor U13283 (N_13283,N_11228,N_10570);
xnor U13284 (N_13284,N_11944,N_11394);
xor U13285 (N_13285,N_12240,N_11621);
nand U13286 (N_13286,N_11278,N_11229);
nand U13287 (N_13287,N_12066,N_10682);
or U13288 (N_13288,N_10044,N_10022);
xor U13289 (N_13289,N_10906,N_10431);
and U13290 (N_13290,N_11410,N_11010);
xor U13291 (N_13291,N_12409,N_10573);
and U13292 (N_13292,N_10181,N_11306);
or U13293 (N_13293,N_11792,N_11385);
xor U13294 (N_13294,N_10173,N_10567);
and U13295 (N_13295,N_12257,N_10824);
nand U13296 (N_13296,N_10117,N_11439);
nand U13297 (N_13297,N_10003,N_12097);
nand U13298 (N_13298,N_10564,N_11842);
and U13299 (N_13299,N_10023,N_10912);
or U13300 (N_13300,N_12110,N_11890);
or U13301 (N_13301,N_11977,N_11587);
nand U13302 (N_13302,N_11050,N_10566);
or U13303 (N_13303,N_11363,N_10895);
xor U13304 (N_13304,N_10462,N_10948);
and U13305 (N_13305,N_11304,N_10257);
nor U13306 (N_13306,N_10619,N_11318);
nand U13307 (N_13307,N_12000,N_10464);
or U13308 (N_13308,N_11643,N_11025);
xor U13309 (N_13309,N_12392,N_10336);
nand U13310 (N_13310,N_11642,N_10897);
and U13311 (N_13311,N_11262,N_10220);
nand U13312 (N_13312,N_11008,N_10504);
or U13313 (N_13313,N_11220,N_10445);
or U13314 (N_13314,N_12386,N_10891);
or U13315 (N_13315,N_10404,N_10451);
and U13316 (N_13316,N_11070,N_12100);
and U13317 (N_13317,N_11250,N_11157);
xnor U13318 (N_13318,N_10109,N_12288);
xnor U13319 (N_13319,N_10405,N_10775);
and U13320 (N_13320,N_11937,N_10828);
and U13321 (N_13321,N_12378,N_10773);
nand U13322 (N_13322,N_12294,N_11028);
and U13323 (N_13323,N_12203,N_12458);
and U13324 (N_13324,N_10432,N_12057);
xnor U13325 (N_13325,N_12259,N_12454);
nor U13326 (N_13326,N_10668,N_10575);
nor U13327 (N_13327,N_10675,N_11572);
or U13328 (N_13328,N_11797,N_11640);
or U13329 (N_13329,N_11093,N_10667);
or U13330 (N_13330,N_11965,N_12492);
or U13331 (N_13331,N_11691,N_10266);
nand U13332 (N_13332,N_10283,N_11308);
and U13333 (N_13333,N_10035,N_11077);
and U13334 (N_13334,N_10943,N_11796);
and U13335 (N_13335,N_12428,N_11666);
xnor U13336 (N_13336,N_10069,N_10397);
or U13337 (N_13337,N_11400,N_11065);
xnor U13338 (N_13338,N_11343,N_12314);
and U13339 (N_13339,N_10925,N_12306);
nor U13340 (N_13340,N_10709,N_11745);
and U13341 (N_13341,N_11254,N_12068);
and U13342 (N_13342,N_12050,N_11909);
nand U13343 (N_13343,N_10321,N_11837);
xnor U13344 (N_13344,N_12471,N_11876);
nand U13345 (N_13345,N_12316,N_12465);
nand U13346 (N_13346,N_11985,N_10577);
or U13347 (N_13347,N_11106,N_11737);
and U13348 (N_13348,N_12365,N_11724);
nand U13349 (N_13349,N_10596,N_12403);
nor U13350 (N_13350,N_11034,N_11271);
xnor U13351 (N_13351,N_11709,N_12192);
or U13352 (N_13352,N_11949,N_11825);
nor U13353 (N_13353,N_10349,N_12177);
nand U13354 (N_13354,N_12160,N_12006);
xor U13355 (N_13355,N_12265,N_10602);
or U13356 (N_13356,N_10650,N_11533);
nor U13357 (N_13357,N_12206,N_10249);
xor U13358 (N_13358,N_12009,N_12301);
and U13359 (N_13359,N_11979,N_11591);
or U13360 (N_13360,N_11844,N_10418);
and U13361 (N_13361,N_10625,N_11183);
nand U13362 (N_13362,N_10241,N_11291);
and U13363 (N_13363,N_10547,N_11904);
nand U13364 (N_13364,N_10355,N_12183);
and U13365 (N_13365,N_11543,N_10700);
or U13366 (N_13366,N_10844,N_10294);
nand U13367 (N_13367,N_11537,N_12220);
nand U13368 (N_13368,N_10206,N_11713);
or U13369 (N_13369,N_11986,N_10080);
nand U13370 (N_13370,N_10176,N_12178);
nand U13371 (N_13371,N_11817,N_11244);
xor U13372 (N_13372,N_11078,N_10245);
nor U13373 (N_13373,N_11335,N_10631);
or U13374 (N_13374,N_11564,N_11598);
and U13375 (N_13375,N_12044,N_10146);
nand U13376 (N_13376,N_10309,N_11793);
nand U13377 (N_13377,N_12028,N_12236);
and U13378 (N_13378,N_10760,N_10998);
nand U13379 (N_13379,N_10217,N_10616);
or U13380 (N_13380,N_10197,N_12047);
and U13381 (N_13381,N_12146,N_12168);
nand U13382 (N_13382,N_10353,N_10621);
nand U13383 (N_13383,N_11460,N_11928);
or U13384 (N_13384,N_10819,N_12333);
and U13385 (N_13385,N_11302,N_11021);
nand U13386 (N_13386,N_12136,N_12001);
nand U13387 (N_13387,N_12238,N_11138);
and U13388 (N_13388,N_11362,N_10059);
nor U13389 (N_13389,N_10480,N_11669);
or U13390 (N_13390,N_10911,N_11814);
nor U13391 (N_13391,N_11170,N_12380);
nand U13392 (N_13392,N_11142,N_10816);
nor U13393 (N_13393,N_12258,N_11911);
xnor U13394 (N_13394,N_12430,N_11951);
nand U13395 (N_13395,N_11323,N_10010);
xor U13396 (N_13396,N_12271,N_10315);
nor U13397 (N_13397,N_10079,N_12345);
and U13398 (N_13398,N_12268,N_11409);
nor U13399 (N_13399,N_11657,N_11866);
nand U13400 (N_13400,N_12444,N_12320);
and U13401 (N_13401,N_11987,N_10203);
and U13402 (N_13402,N_10923,N_10334);
xor U13403 (N_13403,N_11352,N_10467);
xor U13404 (N_13404,N_10196,N_11818);
or U13405 (N_13405,N_11672,N_12494);
nor U13406 (N_13406,N_10459,N_11806);
xnor U13407 (N_13407,N_11618,N_11272);
and U13408 (N_13408,N_11506,N_11576);
and U13409 (N_13409,N_11712,N_10490);
xor U13410 (N_13410,N_12401,N_12139);
nand U13411 (N_13411,N_10924,N_11516);
or U13412 (N_13412,N_12415,N_11031);
nor U13413 (N_13413,N_11003,N_10928);
xnor U13414 (N_13414,N_11490,N_10537);
or U13415 (N_13415,N_11813,N_12280);
and U13416 (N_13416,N_10191,N_11933);
xor U13417 (N_13417,N_10626,N_11286);
and U13418 (N_13418,N_10959,N_10903);
and U13419 (N_13419,N_10793,N_10848);
and U13420 (N_13420,N_11539,N_11693);
xnor U13421 (N_13421,N_10214,N_10839);
nand U13422 (N_13422,N_10651,N_11284);
or U13423 (N_13423,N_11496,N_11457);
xnor U13424 (N_13424,N_10045,N_10549);
nor U13425 (N_13425,N_10159,N_10365);
nand U13426 (N_13426,N_11108,N_10697);
nor U13427 (N_13427,N_11338,N_11594);
nor U13428 (N_13428,N_10393,N_11401);
xor U13429 (N_13429,N_10960,N_10643);
or U13430 (N_13430,N_12482,N_12187);
or U13431 (N_13431,N_11919,N_12129);
and U13432 (N_13432,N_11759,N_10269);
or U13433 (N_13433,N_10918,N_11237);
nand U13434 (N_13434,N_10719,N_12466);
xnor U13435 (N_13435,N_11754,N_12433);
nand U13436 (N_13436,N_10103,N_10361);
or U13437 (N_13437,N_10057,N_10228);
nand U13438 (N_13438,N_12005,N_11210);
xnor U13439 (N_13439,N_12096,N_11176);
and U13440 (N_13440,N_11619,N_11962);
nand U13441 (N_13441,N_11440,N_12331);
nor U13442 (N_13442,N_12055,N_12362);
xor U13443 (N_13443,N_12449,N_10162);
xnor U13444 (N_13444,N_10592,N_10485);
xor U13445 (N_13445,N_10569,N_12016);
and U13446 (N_13446,N_10798,N_11596);
nand U13447 (N_13447,N_11442,N_10155);
nor U13448 (N_13448,N_11348,N_10511);
xor U13449 (N_13449,N_11905,N_12174);
nor U13450 (N_13450,N_10391,N_11734);
or U13451 (N_13451,N_12154,N_10975);
and U13452 (N_13452,N_12445,N_12094);
nor U13453 (N_13453,N_11801,N_12276);
xnor U13454 (N_13454,N_11595,N_10339);
xnor U13455 (N_13455,N_12412,N_12313);
xnor U13456 (N_13456,N_10118,N_12447);
or U13457 (N_13457,N_11775,N_11558);
and U13458 (N_13458,N_10606,N_12453);
and U13459 (N_13459,N_11314,N_11143);
xor U13460 (N_13460,N_11479,N_10061);
or U13461 (N_13461,N_11181,N_11626);
or U13462 (N_13462,N_11269,N_10611);
or U13463 (N_13463,N_11966,N_12251);
or U13464 (N_13464,N_10408,N_11940);
nor U13465 (N_13465,N_10304,N_10961);
nand U13466 (N_13466,N_12284,N_12164);
nor U13467 (N_13467,N_10999,N_10468);
nand U13468 (N_13468,N_10659,N_11921);
and U13469 (N_13469,N_10501,N_11623);
xor U13470 (N_13470,N_11634,N_11350);
xor U13471 (N_13471,N_11897,N_11437);
and U13472 (N_13472,N_10447,N_10935);
or U13473 (N_13473,N_10033,N_10971);
xnor U13474 (N_13474,N_10843,N_10471);
or U13475 (N_13475,N_11499,N_12109);
or U13476 (N_13476,N_12062,N_11682);
nor U13477 (N_13477,N_11863,N_10211);
or U13478 (N_13478,N_10799,N_11934);
xor U13479 (N_13479,N_11322,N_11918);
xnor U13480 (N_13480,N_10093,N_10319);
nor U13481 (N_13481,N_10422,N_10258);
or U13482 (N_13482,N_12012,N_10401);
nor U13483 (N_13483,N_11182,N_10472);
or U13484 (N_13484,N_10424,N_11358);
nand U13485 (N_13485,N_10794,N_11767);
xnor U13486 (N_13486,N_12103,N_11507);
nor U13487 (N_13487,N_10238,N_11259);
xor U13488 (N_13488,N_10689,N_10516);
xnor U13489 (N_13489,N_11152,N_11504);
or U13490 (N_13490,N_12105,N_10419);
nand U13491 (N_13491,N_10586,N_11677);
nor U13492 (N_13492,N_10652,N_10409);
xor U13493 (N_13493,N_10151,N_11492);
and U13494 (N_13494,N_11258,N_11084);
and U13495 (N_13495,N_11223,N_11552);
xnor U13496 (N_13496,N_11821,N_12246);
xor U13497 (N_13497,N_11711,N_10111);
nand U13498 (N_13498,N_11658,N_12169);
or U13499 (N_13499,N_10640,N_11849);
xnor U13500 (N_13500,N_10641,N_11732);
xnor U13501 (N_13501,N_11099,N_10097);
nor U13502 (N_13502,N_10614,N_11992);
or U13503 (N_13503,N_11241,N_10761);
xor U13504 (N_13504,N_11472,N_12003);
nand U13505 (N_13505,N_10874,N_10064);
and U13506 (N_13506,N_11824,N_11330);
nand U13507 (N_13507,N_10486,N_11007);
xnor U13508 (N_13508,N_12321,N_12208);
nand U13509 (N_13509,N_12398,N_12486);
nand U13510 (N_13510,N_10289,N_12216);
or U13511 (N_13511,N_11637,N_11483);
nand U13512 (N_13512,N_10996,N_11203);
and U13513 (N_13513,N_12128,N_11816);
nor U13514 (N_13514,N_10648,N_10553);
or U13515 (N_13515,N_11342,N_11132);
xnor U13516 (N_13516,N_12347,N_11829);
xor U13517 (N_13517,N_10656,N_12499);
and U13518 (N_13518,N_11534,N_10077);
and U13519 (N_13519,N_11695,N_11141);
xnor U13520 (N_13520,N_10936,N_11336);
nor U13521 (N_13521,N_11404,N_12260);
xor U13522 (N_13522,N_11425,N_11776);
nor U13523 (N_13523,N_11943,N_10941);
nand U13524 (N_13524,N_11200,N_10031);
nand U13525 (N_13525,N_12360,N_11562);
or U13526 (N_13526,N_10141,N_11468);
nand U13527 (N_13527,N_10016,N_10937);
and U13528 (N_13528,N_10312,N_11179);
or U13529 (N_13529,N_11012,N_10900);
and U13530 (N_13530,N_10457,N_10411);
nand U13531 (N_13531,N_12413,N_11196);
nor U13532 (N_13532,N_12079,N_10593);
or U13533 (N_13533,N_10947,N_11105);
xnor U13534 (N_13534,N_11553,N_10556);
and U13535 (N_13535,N_10272,N_10545);
nand U13536 (N_13536,N_11436,N_11054);
or U13537 (N_13537,N_10006,N_11466);
xnor U13538 (N_13538,N_10600,N_12048);
or U13539 (N_13539,N_11926,N_10541);
nand U13540 (N_13540,N_10058,N_11296);
and U13541 (N_13541,N_11556,N_11213);
or U13542 (N_13542,N_10725,N_11726);
and U13543 (N_13543,N_11528,N_10646);
xnor U13544 (N_13544,N_12332,N_10847);
nor U13545 (N_13545,N_11347,N_10430);
or U13546 (N_13546,N_10116,N_11167);
nand U13547 (N_13547,N_10172,N_10762);
nand U13548 (N_13548,N_10774,N_10841);
xor U13549 (N_13549,N_12439,N_10855);
nor U13550 (N_13550,N_10587,N_12390);
nand U13551 (N_13551,N_12150,N_12406);
nand U13552 (N_13552,N_10543,N_10559);
nor U13553 (N_13553,N_12202,N_12134);
nand U13554 (N_13554,N_11735,N_12488);
or U13555 (N_13555,N_10094,N_10004);
nand U13556 (N_13556,N_11638,N_11555);
and U13557 (N_13557,N_11827,N_10898);
nor U13558 (N_13558,N_10665,N_11252);
xnor U13559 (N_13559,N_12363,N_12124);
xor U13560 (N_13560,N_11851,N_11211);
and U13561 (N_13561,N_11699,N_10183);
xnor U13562 (N_13562,N_10779,N_10699);
and U13563 (N_13563,N_11032,N_10179);
and U13564 (N_13564,N_10676,N_11487);
xnor U13565 (N_13565,N_10813,N_11019);
nor U13566 (N_13566,N_10831,N_10222);
and U13567 (N_13567,N_10856,N_11822);
and U13568 (N_13568,N_11002,N_10030);
or U13569 (N_13569,N_11953,N_11353);
and U13570 (N_13570,N_12191,N_12215);
or U13571 (N_13571,N_11575,N_10020);
or U13572 (N_13572,N_10908,N_10521);
nor U13573 (N_13573,N_12018,N_10303);
and U13574 (N_13574,N_11364,N_12087);
nand U13575 (N_13575,N_10617,N_10518);
nand U13576 (N_13576,N_10402,N_11710);
nor U13577 (N_13577,N_11501,N_12429);
nand U13578 (N_13578,N_10477,N_12027);
and U13579 (N_13579,N_11421,N_11886);
nor U13580 (N_13580,N_12227,N_10952);
nor U13581 (N_13581,N_10812,N_11557);
or U13582 (N_13582,N_10745,N_10140);
nor U13583 (N_13583,N_11725,N_10114);
and U13584 (N_13584,N_11165,N_10713);
xnor U13585 (N_13585,N_10073,N_10032);
xor U13586 (N_13586,N_11502,N_12088);
or U13587 (N_13587,N_11683,N_11653);
nand U13588 (N_13588,N_11429,N_12384);
xor U13589 (N_13589,N_10753,N_11384);
nand U13590 (N_13590,N_11529,N_10046);
nor U13591 (N_13591,N_10679,N_12030);
and U13592 (N_13592,N_12487,N_12135);
xor U13593 (N_13593,N_11820,N_10744);
and U13594 (N_13594,N_10039,N_10735);
xnor U13595 (N_13595,N_10483,N_10796);
xnor U13596 (N_13596,N_11980,N_12228);
xor U13597 (N_13597,N_10913,N_10153);
xnor U13598 (N_13598,N_11476,N_10681);
or U13599 (N_13599,N_12330,N_11446);
xnor U13600 (N_13600,N_11765,N_12410);
xnor U13601 (N_13601,N_10112,N_10638);
nor U13602 (N_13602,N_10161,N_11146);
xor U13603 (N_13603,N_10962,N_10384);
nor U13604 (N_13604,N_10372,N_10684);
xnor U13605 (N_13605,N_10854,N_12085);
and U13606 (N_13606,N_11115,N_11809);
and U13607 (N_13607,N_12279,N_11103);
and U13608 (N_13608,N_11150,N_11349);
nand U13609 (N_13609,N_11903,N_11981);
or U13610 (N_13610,N_12327,N_11706);
nor U13611 (N_13611,N_10750,N_11192);
nand U13612 (N_13612,N_12029,N_11290);
and U13613 (N_13613,N_12489,N_11627);
or U13614 (N_13614,N_10458,N_12155);
xor U13615 (N_13615,N_11292,N_12455);
nor U13616 (N_13616,N_11068,N_10513);
or U13617 (N_13617,N_11493,N_10367);
nand U13618 (N_13618,N_11217,N_10364);
or U13619 (N_13619,N_11147,N_10933);
or U13620 (N_13620,N_11671,N_11198);
xor U13621 (N_13621,N_10129,N_11927);
or U13622 (N_13622,N_11995,N_10138);
or U13623 (N_13623,N_11798,N_11571);
or U13624 (N_13624,N_11525,N_10703);
xor U13625 (N_13625,N_10157,N_10618);
and U13626 (N_13626,N_11222,N_11120);
nand U13627 (N_13627,N_11415,N_11014);
or U13628 (N_13628,N_10437,N_11498);
xnor U13629 (N_13629,N_11530,N_11164);
and U13630 (N_13630,N_12419,N_12034);
nand U13631 (N_13631,N_10086,N_10288);
nor U13632 (N_13632,N_11679,N_11770);
xor U13633 (N_13633,N_12141,N_10452);
nor U13634 (N_13634,N_11729,N_12032);
nand U13635 (N_13635,N_12207,N_12423);
or U13636 (N_13636,N_11316,N_11202);
nor U13637 (N_13637,N_10285,N_11573);
nand U13638 (N_13638,N_11879,N_11744);
xor U13639 (N_13639,N_10645,N_10879);
nor U13640 (N_13640,N_11645,N_10286);
nand U13641 (N_13641,N_11912,N_12080);
nor U13642 (N_13642,N_10481,N_10192);
nor U13643 (N_13643,N_11319,N_10784);
and U13644 (N_13644,N_10988,N_12011);
nand U13645 (N_13645,N_10765,N_11678);
nand U13646 (N_13646,N_12126,N_10328);
xor U13647 (N_13647,N_10036,N_11612);
nor U13648 (N_13648,N_11260,N_10930);
nand U13649 (N_13649,N_10343,N_10202);
xor U13650 (N_13650,N_10993,N_10305);
or U13651 (N_13651,N_12323,N_10669);
nand U13652 (N_13652,N_10867,N_10476);
or U13653 (N_13653,N_11184,N_10494);
and U13654 (N_13654,N_11274,N_10767);
nor U13655 (N_13655,N_11341,N_10316);
and U13656 (N_13656,N_12024,N_10075);
and U13657 (N_13657,N_12132,N_10972);
xor U13658 (N_13658,N_12119,N_12291);
xnor U13659 (N_13659,N_10297,N_10731);
nor U13660 (N_13660,N_11379,N_11871);
nand U13661 (N_13661,N_10884,N_11005);
nor U13662 (N_13662,N_12275,N_12283);
and U13663 (N_13663,N_11915,N_11419);
and U13664 (N_13664,N_10386,N_10331);
nor U13665 (N_13665,N_10896,N_10919);
and U13666 (N_13666,N_10533,N_11491);
nand U13667 (N_13667,N_12015,N_10707);
or U13668 (N_13668,N_11061,N_10583);
or U13669 (N_13669,N_11722,N_10265);
nor U13670 (N_13670,N_10787,N_10951);
nor U13671 (N_13671,N_11020,N_10717);
nor U13672 (N_13672,N_11043,N_10830);
or U13673 (N_13673,N_10514,N_10348);
and U13674 (N_13674,N_10322,N_11624);
nor U13675 (N_13675,N_10392,N_11900);
xnor U13676 (N_13676,N_10818,N_10917);
nand U13677 (N_13677,N_12075,N_12104);
or U13678 (N_13678,N_10473,N_10894);
nand U13679 (N_13679,N_11752,N_10805);
nand U13680 (N_13680,N_10226,N_10332);
xnor U13681 (N_13681,N_11397,N_12144);
and U13682 (N_13682,N_11326,N_11913);
nand U13683 (N_13683,N_10237,N_12059);
or U13684 (N_13684,N_10662,N_10934);
xor U13685 (N_13685,N_10846,N_10690);
and U13686 (N_13686,N_11843,N_11048);
nand U13687 (N_13687,N_12190,N_11720);
nor U13688 (N_13688,N_11938,N_10849);
and U13689 (N_13689,N_10623,N_10955);
nor U13690 (N_13690,N_10177,N_11096);
nand U13691 (N_13691,N_10098,N_10373);
and U13692 (N_13692,N_12008,N_11689);
nor U13693 (N_13693,N_12462,N_11848);
nor U13694 (N_13694,N_11920,N_11452);
nand U13695 (N_13695,N_12004,N_12324);
nand U13696 (N_13696,N_11721,N_11613);
and U13697 (N_13697,N_12122,N_11999);
nor U13698 (N_13698,N_10453,N_11763);
nand U13699 (N_13699,N_10814,N_10190);
nor U13700 (N_13700,N_10783,N_10123);
and U13701 (N_13701,N_11603,N_10949);
and U13702 (N_13702,N_11287,N_12277);
and U13703 (N_13703,N_10766,N_10106);
nor U13704 (N_13704,N_10246,N_12267);
nor U13705 (N_13705,N_11967,N_10262);
xor U13706 (N_13706,N_10647,N_10565);
nor U13707 (N_13707,N_11495,N_11245);
nor U13708 (N_13708,N_10620,N_11766);
nand U13709 (N_13709,N_11137,N_10307);
or U13710 (N_13710,N_12296,N_10329);
nand U13711 (N_13711,N_10797,N_10644);
nor U13712 (N_13712,N_10280,N_10749);
nor U13713 (N_13713,N_10827,N_10219);
or U13714 (N_13714,N_10868,N_10604);
xnor U13715 (N_13715,N_11119,N_11771);
nor U13716 (N_13716,N_11894,N_10132);
or U13717 (N_13717,N_11730,N_12373);
and U13718 (N_13718,N_11230,N_10096);
or U13719 (N_13719,N_12091,N_12038);
xnor U13720 (N_13720,N_10829,N_10711);
xnor U13721 (N_13721,N_12130,N_12125);
nand U13722 (N_13722,N_11475,N_10523);
nand U13723 (N_13723,N_10406,N_11298);
nand U13724 (N_13724,N_10273,N_12247);
nand U13725 (N_13725,N_11317,N_10170);
nand U13726 (N_13726,N_10987,N_11267);
xnor U13727 (N_13727,N_11158,N_11443);
nand U13728 (N_13728,N_10603,N_12336);
or U13729 (N_13729,N_11535,N_10456);
nor U13730 (N_13730,N_11369,N_11935);
and U13731 (N_13731,N_11674,N_12387);
xnor U13732 (N_13732,N_11136,N_11067);
or U13733 (N_13733,N_10144,N_10420);
or U13734 (N_13734,N_11159,N_11373);
and U13735 (N_13735,N_11473,N_12344);
xor U13736 (N_13736,N_11704,N_12188);
and U13737 (N_13737,N_10743,N_10239);
and U13738 (N_13738,N_12262,N_10415);
nand U13739 (N_13739,N_10497,N_12116);
nand U13740 (N_13740,N_10763,N_11800);
and U13741 (N_13741,N_11402,N_12309);
and U13742 (N_13742,N_11413,N_10029);
and U13743 (N_13743,N_10658,N_11293);
and U13744 (N_13744,N_10755,N_10070);
xor U13745 (N_13745,N_10275,N_11964);
nor U13746 (N_13746,N_10037,N_12121);
xnor U13747 (N_13747,N_11968,N_12269);
or U13748 (N_13748,N_10664,N_11656);
nand U13749 (N_13749,N_11519,N_11464);
and U13750 (N_13750,N_10097,N_10059);
nand U13751 (N_13751,N_10631,N_11468);
nand U13752 (N_13752,N_12399,N_12270);
xnor U13753 (N_13753,N_10176,N_10059);
or U13754 (N_13754,N_10256,N_11460);
nor U13755 (N_13755,N_12063,N_10142);
xnor U13756 (N_13756,N_10347,N_10344);
nor U13757 (N_13757,N_11113,N_12088);
and U13758 (N_13758,N_11898,N_11510);
xnor U13759 (N_13759,N_12331,N_11403);
nor U13760 (N_13760,N_10958,N_10093);
or U13761 (N_13761,N_11574,N_11590);
and U13762 (N_13762,N_11362,N_10633);
nor U13763 (N_13763,N_10974,N_10687);
nor U13764 (N_13764,N_11632,N_11064);
or U13765 (N_13765,N_10653,N_12213);
and U13766 (N_13766,N_12075,N_10932);
and U13767 (N_13767,N_11996,N_10735);
nor U13768 (N_13768,N_10671,N_11251);
or U13769 (N_13769,N_11524,N_10192);
xnor U13770 (N_13770,N_11617,N_11228);
or U13771 (N_13771,N_12167,N_10660);
and U13772 (N_13772,N_11706,N_11733);
nor U13773 (N_13773,N_11149,N_11289);
xor U13774 (N_13774,N_11784,N_12000);
and U13775 (N_13775,N_10247,N_10014);
xor U13776 (N_13776,N_11777,N_11078);
and U13777 (N_13777,N_10519,N_11224);
or U13778 (N_13778,N_11148,N_10468);
or U13779 (N_13779,N_11755,N_12390);
nand U13780 (N_13780,N_11919,N_10706);
xnor U13781 (N_13781,N_11803,N_11773);
nor U13782 (N_13782,N_11349,N_11465);
or U13783 (N_13783,N_11409,N_11327);
nand U13784 (N_13784,N_10991,N_10812);
nor U13785 (N_13785,N_10737,N_11427);
xnor U13786 (N_13786,N_10212,N_12395);
or U13787 (N_13787,N_11675,N_11416);
nand U13788 (N_13788,N_12004,N_12057);
or U13789 (N_13789,N_12224,N_10648);
xor U13790 (N_13790,N_12105,N_10874);
or U13791 (N_13791,N_10949,N_10116);
or U13792 (N_13792,N_10754,N_10297);
nor U13793 (N_13793,N_11055,N_12030);
xnor U13794 (N_13794,N_11224,N_12291);
nor U13795 (N_13795,N_11131,N_11023);
xor U13796 (N_13796,N_12257,N_10358);
nor U13797 (N_13797,N_12043,N_12417);
and U13798 (N_13798,N_11686,N_10451);
xor U13799 (N_13799,N_10308,N_10537);
nand U13800 (N_13800,N_10917,N_11719);
or U13801 (N_13801,N_11509,N_12029);
or U13802 (N_13802,N_10611,N_11505);
nor U13803 (N_13803,N_10840,N_10626);
xor U13804 (N_13804,N_10411,N_10623);
nand U13805 (N_13805,N_10823,N_10662);
xnor U13806 (N_13806,N_12336,N_11139);
and U13807 (N_13807,N_10749,N_10540);
nor U13808 (N_13808,N_11492,N_11904);
or U13809 (N_13809,N_10184,N_11359);
or U13810 (N_13810,N_10205,N_12164);
and U13811 (N_13811,N_10467,N_11779);
xor U13812 (N_13812,N_11838,N_10958);
and U13813 (N_13813,N_11257,N_10357);
xnor U13814 (N_13814,N_11284,N_10440);
nand U13815 (N_13815,N_11613,N_10815);
nor U13816 (N_13816,N_11695,N_11312);
xnor U13817 (N_13817,N_12274,N_11677);
xor U13818 (N_13818,N_12062,N_10255);
nand U13819 (N_13819,N_10453,N_12156);
and U13820 (N_13820,N_10025,N_10863);
or U13821 (N_13821,N_11766,N_11111);
nand U13822 (N_13822,N_11691,N_11130);
nand U13823 (N_13823,N_10296,N_10055);
xnor U13824 (N_13824,N_11607,N_12152);
nor U13825 (N_13825,N_11739,N_10684);
or U13826 (N_13826,N_12382,N_11802);
nor U13827 (N_13827,N_11415,N_10524);
and U13828 (N_13828,N_10652,N_12485);
nor U13829 (N_13829,N_12019,N_10159);
xnor U13830 (N_13830,N_11833,N_10040);
and U13831 (N_13831,N_10228,N_10078);
and U13832 (N_13832,N_11515,N_10739);
xor U13833 (N_13833,N_10663,N_10557);
nand U13834 (N_13834,N_11629,N_12319);
nor U13835 (N_13835,N_12375,N_10267);
nor U13836 (N_13836,N_12237,N_11364);
and U13837 (N_13837,N_12030,N_11087);
nand U13838 (N_13838,N_12448,N_10257);
or U13839 (N_13839,N_10015,N_10839);
nor U13840 (N_13840,N_10705,N_10183);
nand U13841 (N_13841,N_10146,N_12032);
xor U13842 (N_13842,N_12122,N_11149);
xor U13843 (N_13843,N_12223,N_10391);
xnor U13844 (N_13844,N_12080,N_12216);
nor U13845 (N_13845,N_12339,N_10819);
nand U13846 (N_13846,N_10727,N_11513);
and U13847 (N_13847,N_11120,N_11432);
and U13848 (N_13848,N_12337,N_12358);
or U13849 (N_13849,N_11223,N_11817);
nand U13850 (N_13850,N_11736,N_10206);
and U13851 (N_13851,N_10197,N_11142);
and U13852 (N_13852,N_11190,N_12246);
and U13853 (N_13853,N_10385,N_10462);
xnor U13854 (N_13854,N_11894,N_10901);
or U13855 (N_13855,N_12270,N_11654);
nor U13856 (N_13856,N_10062,N_12095);
nor U13857 (N_13857,N_11846,N_12457);
xor U13858 (N_13858,N_10609,N_10050);
or U13859 (N_13859,N_10376,N_10581);
nor U13860 (N_13860,N_12067,N_10951);
nor U13861 (N_13861,N_10092,N_10050);
nand U13862 (N_13862,N_10463,N_10133);
nand U13863 (N_13863,N_10489,N_10625);
nand U13864 (N_13864,N_12212,N_10568);
or U13865 (N_13865,N_11326,N_10277);
or U13866 (N_13866,N_11893,N_12482);
xnor U13867 (N_13867,N_12280,N_10794);
nor U13868 (N_13868,N_12201,N_11360);
and U13869 (N_13869,N_12006,N_12176);
or U13870 (N_13870,N_11679,N_12263);
xnor U13871 (N_13871,N_11830,N_11524);
and U13872 (N_13872,N_11501,N_10478);
xor U13873 (N_13873,N_12010,N_10408);
nor U13874 (N_13874,N_12441,N_10213);
nand U13875 (N_13875,N_11672,N_10430);
and U13876 (N_13876,N_11971,N_12347);
nor U13877 (N_13877,N_11084,N_11960);
xor U13878 (N_13878,N_11313,N_10794);
or U13879 (N_13879,N_12175,N_10683);
xnor U13880 (N_13880,N_11868,N_11222);
nor U13881 (N_13881,N_10117,N_10949);
nand U13882 (N_13882,N_10945,N_10656);
nand U13883 (N_13883,N_11233,N_11903);
xor U13884 (N_13884,N_11250,N_11830);
xnor U13885 (N_13885,N_11753,N_10378);
or U13886 (N_13886,N_10840,N_12499);
nand U13887 (N_13887,N_12450,N_11861);
nand U13888 (N_13888,N_10856,N_12366);
nor U13889 (N_13889,N_11803,N_12188);
xnor U13890 (N_13890,N_11082,N_11850);
nor U13891 (N_13891,N_10995,N_12166);
nor U13892 (N_13892,N_10706,N_10237);
nand U13893 (N_13893,N_10095,N_10472);
nand U13894 (N_13894,N_11892,N_10921);
xnor U13895 (N_13895,N_12021,N_11862);
xor U13896 (N_13896,N_10586,N_10108);
nand U13897 (N_13897,N_12062,N_11086);
nand U13898 (N_13898,N_12392,N_11717);
xnor U13899 (N_13899,N_11550,N_11400);
nand U13900 (N_13900,N_11163,N_10072);
and U13901 (N_13901,N_10854,N_11999);
and U13902 (N_13902,N_10839,N_11916);
nor U13903 (N_13903,N_11944,N_12174);
xor U13904 (N_13904,N_12497,N_11930);
nand U13905 (N_13905,N_10487,N_10159);
nand U13906 (N_13906,N_11897,N_11240);
xnor U13907 (N_13907,N_11080,N_11333);
and U13908 (N_13908,N_10430,N_11212);
and U13909 (N_13909,N_12285,N_10908);
nand U13910 (N_13910,N_10488,N_12186);
and U13911 (N_13911,N_10167,N_11178);
or U13912 (N_13912,N_10989,N_10694);
xor U13913 (N_13913,N_10938,N_10854);
nor U13914 (N_13914,N_10169,N_11292);
nor U13915 (N_13915,N_10390,N_12165);
nor U13916 (N_13916,N_11652,N_11275);
xor U13917 (N_13917,N_10029,N_11770);
or U13918 (N_13918,N_12280,N_11981);
xor U13919 (N_13919,N_11647,N_10738);
xnor U13920 (N_13920,N_11405,N_11717);
nand U13921 (N_13921,N_11098,N_11382);
xnor U13922 (N_13922,N_12258,N_10777);
or U13923 (N_13923,N_11077,N_10213);
and U13924 (N_13924,N_10600,N_11600);
nand U13925 (N_13925,N_11267,N_10874);
nor U13926 (N_13926,N_12497,N_10977);
nor U13927 (N_13927,N_10406,N_12171);
nand U13928 (N_13928,N_10164,N_10223);
xor U13929 (N_13929,N_12018,N_11963);
nor U13930 (N_13930,N_10742,N_10405);
nor U13931 (N_13931,N_12224,N_11100);
and U13932 (N_13932,N_11465,N_11038);
xnor U13933 (N_13933,N_10960,N_11431);
and U13934 (N_13934,N_10854,N_11087);
and U13935 (N_13935,N_12476,N_10016);
and U13936 (N_13936,N_10876,N_10438);
or U13937 (N_13937,N_11987,N_10741);
and U13938 (N_13938,N_12075,N_11070);
nand U13939 (N_13939,N_12271,N_11235);
or U13940 (N_13940,N_10045,N_12054);
nand U13941 (N_13941,N_11291,N_10318);
nand U13942 (N_13942,N_12286,N_12307);
xnor U13943 (N_13943,N_10988,N_12478);
or U13944 (N_13944,N_12450,N_10179);
and U13945 (N_13945,N_11312,N_10411);
xor U13946 (N_13946,N_10268,N_11724);
nand U13947 (N_13947,N_11928,N_10525);
xnor U13948 (N_13948,N_11755,N_10013);
or U13949 (N_13949,N_10527,N_12229);
or U13950 (N_13950,N_10506,N_10399);
and U13951 (N_13951,N_11409,N_10560);
and U13952 (N_13952,N_11593,N_10607);
and U13953 (N_13953,N_12400,N_12387);
or U13954 (N_13954,N_11528,N_10745);
nand U13955 (N_13955,N_10736,N_11661);
or U13956 (N_13956,N_10986,N_10670);
nand U13957 (N_13957,N_10637,N_10835);
and U13958 (N_13958,N_11928,N_10528);
xor U13959 (N_13959,N_12196,N_10870);
nand U13960 (N_13960,N_12028,N_11996);
and U13961 (N_13961,N_10530,N_11573);
nand U13962 (N_13962,N_12278,N_11169);
or U13963 (N_13963,N_11985,N_11647);
and U13964 (N_13964,N_11261,N_11252);
nand U13965 (N_13965,N_10807,N_10330);
nor U13966 (N_13966,N_12371,N_10905);
xnor U13967 (N_13967,N_11997,N_10845);
nand U13968 (N_13968,N_10613,N_11364);
nand U13969 (N_13969,N_11163,N_11007);
nor U13970 (N_13970,N_10584,N_10853);
nor U13971 (N_13971,N_11448,N_10147);
and U13972 (N_13972,N_10527,N_10787);
xnor U13973 (N_13973,N_10019,N_12005);
nor U13974 (N_13974,N_10970,N_10116);
and U13975 (N_13975,N_10912,N_10500);
or U13976 (N_13976,N_11593,N_10378);
or U13977 (N_13977,N_11471,N_11130);
xor U13978 (N_13978,N_11290,N_10719);
nor U13979 (N_13979,N_11259,N_11058);
nor U13980 (N_13980,N_11080,N_11442);
nor U13981 (N_13981,N_10864,N_11858);
nor U13982 (N_13982,N_12097,N_10884);
or U13983 (N_13983,N_11594,N_11670);
or U13984 (N_13984,N_11010,N_10528);
or U13985 (N_13985,N_12039,N_12311);
or U13986 (N_13986,N_10588,N_11265);
nand U13987 (N_13987,N_11403,N_11405);
nand U13988 (N_13988,N_10678,N_10894);
or U13989 (N_13989,N_10381,N_10940);
and U13990 (N_13990,N_12244,N_11892);
and U13991 (N_13991,N_10827,N_12161);
and U13992 (N_13992,N_11362,N_12369);
and U13993 (N_13993,N_10526,N_12300);
nor U13994 (N_13994,N_10092,N_11969);
xor U13995 (N_13995,N_12493,N_10634);
and U13996 (N_13996,N_12197,N_10517);
nor U13997 (N_13997,N_11876,N_10341);
or U13998 (N_13998,N_12083,N_12153);
or U13999 (N_13999,N_12141,N_10346);
xor U14000 (N_14000,N_11304,N_10944);
xor U14001 (N_14001,N_11873,N_11122);
nor U14002 (N_14002,N_11819,N_10986);
and U14003 (N_14003,N_12367,N_12388);
or U14004 (N_14004,N_11672,N_12306);
nand U14005 (N_14005,N_11534,N_10730);
and U14006 (N_14006,N_11842,N_11690);
nor U14007 (N_14007,N_10499,N_10226);
nand U14008 (N_14008,N_11251,N_11734);
and U14009 (N_14009,N_10192,N_10579);
or U14010 (N_14010,N_10337,N_10263);
and U14011 (N_14011,N_10076,N_10389);
xor U14012 (N_14012,N_11783,N_11325);
xnor U14013 (N_14013,N_11105,N_11452);
or U14014 (N_14014,N_12391,N_10142);
or U14015 (N_14015,N_11664,N_11656);
nand U14016 (N_14016,N_12279,N_11154);
or U14017 (N_14017,N_11416,N_11569);
and U14018 (N_14018,N_10951,N_10606);
or U14019 (N_14019,N_11930,N_10980);
nor U14020 (N_14020,N_10775,N_12318);
and U14021 (N_14021,N_10659,N_11531);
or U14022 (N_14022,N_11992,N_10530);
and U14023 (N_14023,N_11051,N_11242);
or U14024 (N_14024,N_10975,N_10532);
nand U14025 (N_14025,N_10939,N_10947);
xnor U14026 (N_14026,N_11709,N_12130);
or U14027 (N_14027,N_10121,N_10298);
xor U14028 (N_14028,N_11890,N_11701);
xnor U14029 (N_14029,N_10137,N_10962);
xnor U14030 (N_14030,N_10054,N_10874);
or U14031 (N_14031,N_12345,N_11044);
nor U14032 (N_14032,N_10470,N_11409);
nor U14033 (N_14033,N_10305,N_12382);
and U14034 (N_14034,N_10530,N_11844);
nand U14035 (N_14035,N_10841,N_10372);
xor U14036 (N_14036,N_12003,N_12428);
xnor U14037 (N_14037,N_10067,N_11532);
xnor U14038 (N_14038,N_12187,N_10471);
and U14039 (N_14039,N_10020,N_12181);
nor U14040 (N_14040,N_12461,N_11108);
or U14041 (N_14041,N_10283,N_12230);
and U14042 (N_14042,N_11848,N_11725);
nand U14043 (N_14043,N_10380,N_10849);
nor U14044 (N_14044,N_10220,N_12482);
nand U14045 (N_14045,N_10246,N_11609);
or U14046 (N_14046,N_12180,N_11129);
and U14047 (N_14047,N_10753,N_10403);
and U14048 (N_14048,N_10914,N_11073);
nor U14049 (N_14049,N_11612,N_12308);
xnor U14050 (N_14050,N_11140,N_12125);
nor U14051 (N_14051,N_10514,N_11620);
nor U14052 (N_14052,N_10837,N_10529);
and U14053 (N_14053,N_10426,N_12039);
and U14054 (N_14054,N_11347,N_11983);
or U14055 (N_14055,N_10899,N_12491);
nand U14056 (N_14056,N_11098,N_10519);
nor U14057 (N_14057,N_10012,N_11101);
or U14058 (N_14058,N_11305,N_12152);
nand U14059 (N_14059,N_11417,N_10626);
and U14060 (N_14060,N_11396,N_11960);
or U14061 (N_14061,N_12338,N_11853);
xnor U14062 (N_14062,N_12444,N_10745);
xnor U14063 (N_14063,N_12393,N_11942);
and U14064 (N_14064,N_10883,N_12258);
or U14065 (N_14065,N_10199,N_10427);
and U14066 (N_14066,N_10277,N_12316);
and U14067 (N_14067,N_11936,N_11847);
nand U14068 (N_14068,N_10356,N_10383);
xnor U14069 (N_14069,N_11092,N_11890);
or U14070 (N_14070,N_10559,N_11041);
nor U14071 (N_14071,N_11632,N_10803);
nor U14072 (N_14072,N_10152,N_11725);
or U14073 (N_14073,N_12165,N_12028);
or U14074 (N_14074,N_10041,N_12454);
xnor U14075 (N_14075,N_10557,N_11664);
and U14076 (N_14076,N_10095,N_10030);
xor U14077 (N_14077,N_10310,N_10460);
nor U14078 (N_14078,N_10537,N_11252);
xnor U14079 (N_14079,N_10376,N_10052);
xor U14080 (N_14080,N_10065,N_10409);
nor U14081 (N_14081,N_10803,N_10165);
or U14082 (N_14082,N_12066,N_12282);
nand U14083 (N_14083,N_10434,N_12088);
nor U14084 (N_14084,N_10638,N_11698);
and U14085 (N_14085,N_12280,N_11707);
nand U14086 (N_14086,N_11405,N_11106);
nor U14087 (N_14087,N_12470,N_10781);
and U14088 (N_14088,N_10360,N_11050);
nor U14089 (N_14089,N_11110,N_11209);
or U14090 (N_14090,N_11099,N_12035);
or U14091 (N_14091,N_10643,N_11210);
or U14092 (N_14092,N_12115,N_10738);
nand U14093 (N_14093,N_12334,N_10386);
xnor U14094 (N_14094,N_10338,N_11438);
nor U14095 (N_14095,N_11392,N_10255);
nor U14096 (N_14096,N_10605,N_10932);
or U14097 (N_14097,N_11422,N_11615);
or U14098 (N_14098,N_11515,N_11006);
or U14099 (N_14099,N_12363,N_11968);
xnor U14100 (N_14100,N_11400,N_11233);
nor U14101 (N_14101,N_10430,N_12152);
nand U14102 (N_14102,N_10755,N_10314);
or U14103 (N_14103,N_11650,N_10739);
nand U14104 (N_14104,N_10297,N_10753);
xor U14105 (N_14105,N_12145,N_10881);
or U14106 (N_14106,N_12367,N_10438);
xnor U14107 (N_14107,N_10436,N_10369);
and U14108 (N_14108,N_12250,N_10591);
and U14109 (N_14109,N_10455,N_10959);
xor U14110 (N_14110,N_11811,N_10694);
xor U14111 (N_14111,N_10217,N_11358);
nand U14112 (N_14112,N_11304,N_12127);
or U14113 (N_14113,N_12151,N_11281);
or U14114 (N_14114,N_12194,N_11977);
nor U14115 (N_14115,N_11789,N_11028);
and U14116 (N_14116,N_10761,N_11848);
xnor U14117 (N_14117,N_10226,N_12317);
xnor U14118 (N_14118,N_11091,N_10964);
or U14119 (N_14119,N_10178,N_10539);
or U14120 (N_14120,N_10139,N_11790);
or U14121 (N_14121,N_12022,N_11584);
or U14122 (N_14122,N_11755,N_11270);
xor U14123 (N_14123,N_12201,N_12178);
and U14124 (N_14124,N_12225,N_10846);
nand U14125 (N_14125,N_10889,N_11283);
and U14126 (N_14126,N_11803,N_11963);
or U14127 (N_14127,N_10031,N_10308);
xnor U14128 (N_14128,N_11945,N_10730);
nand U14129 (N_14129,N_11189,N_12313);
nand U14130 (N_14130,N_11224,N_10880);
xnor U14131 (N_14131,N_12493,N_10788);
nor U14132 (N_14132,N_10370,N_10626);
nor U14133 (N_14133,N_11319,N_12474);
nand U14134 (N_14134,N_10687,N_11492);
and U14135 (N_14135,N_12312,N_12420);
xor U14136 (N_14136,N_11172,N_10534);
nand U14137 (N_14137,N_11554,N_11172);
nand U14138 (N_14138,N_11268,N_12324);
nand U14139 (N_14139,N_11863,N_10011);
nand U14140 (N_14140,N_11005,N_11981);
xnor U14141 (N_14141,N_11547,N_10950);
or U14142 (N_14142,N_12423,N_10833);
xnor U14143 (N_14143,N_11766,N_11275);
xnor U14144 (N_14144,N_11885,N_11964);
xnor U14145 (N_14145,N_12394,N_10846);
or U14146 (N_14146,N_12236,N_11836);
xnor U14147 (N_14147,N_12431,N_10949);
or U14148 (N_14148,N_10322,N_12049);
xnor U14149 (N_14149,N_10282,N_10315);
xor U14150 (N_14150,N_10758,N_11718);
nand U14151 (N_14151,N_12100,N_10064);
nand U14152 (N_14152,N_10348,N_11653);
nand U14153 (N_14153,N_11333,N_10052);
nand U14154 (N_14154,N_11801,N_11661);
nor U14155 (N_14155,N_11417,N_11693);
or U14156 (N_14156,N_10438,N_11637);
or U14157 (N_14157,N_11750,N_12393);
and U14158 (N_14158,N_12319,N_12269);
nand U14159 (N_14159,N_11881,N_11222);
or U14160 (N_14160,N_10279,N_10653);
nand U14161 (N_14161,N_11207,N_11392);
and U14162 (N_14162,N_10624,N_10436);
or U14163 (N_14163,N_10783,N_10562);
nor U14164 (N_14164,N_11228,N_11923);
xnor U14165 (N_14165,N_11205,N_10364);
xnor U14166 (N_14166,N_10319,N_10505);
nor U14167 (N_14167,N_10652,N_11465);
or U14168 (N_14168,N_11431,N_11283);
nor U14169 (N_14169,N_11881,N_11050);
xnor U14170 (N_14170,N_11309,N_10790);
nor U14171 (N_14171,N_11021,N_10692);
or U14172 (N_14172,N_10651,N_11536);
nor U14173 (N_14173,N_10171,N_10201);
or U14174 (N_14174,N_10928,N_12047);
or U14175 (N_14175,N_10948,N_10017);
nor U14176 (N_14176,N_12327,N_12098);
or U14177 (N_14177,N_10222,N_10281);
nor U14178 (N_14178,N_11330,N_10425);
nand U14179 (N_14179,N_12273,N_11157);
nor U14180 (N_14180,N_11070,N_10268);
nor U14181 (N_14181,N_12380,N_10471);
and U14182 (N_14182,N_10738,N_11230);
or U14183 (N_14183,N_10950,N_11002);
and U14184 (N_14184,N_10046,N_11184);
nand U14185 (N_14185,N_10098,N_11249);
and U14186 (N_14186,N_11896,N_10334);
xnor U14187 (N_14187,N_11181,N_10399);
and U14188 (N_14188,N_11937,N_10832);
nor U14189 (N_14189,N_10529,N_11183);
or U14190 (N_14190,N_10600,N_10420);
xnor U14191 (N_14191,N_11313,N_10251);
nor U14192 (N_14192,N_12359,N_12429);
nor U14193 (N_14193,N_11600,N_12039);
nand U14194 (N_14194,N_10672,N_10067);
xor U14195 (N_14195,N_11737,N_10415);
or U14196 (N_14196,N_11778,N_11331);
xor U14197 (N_14197,N_11292,N_10057);
nand U14198 (N_14198,N_10503,N_10351);
xnor U14199 (N_14199,N_11570,N_12306);
nand U14200 (N_14200,N_11415,N_11546);
or U14201 (N_14201,N_10573,N_11019);
nand U14202 (N_14202,N_10803,N_11201);
or U14203 (N_14203,N_10365,N_10394);
nand U14204 (N_14204,N_12190,N_10974);
xnor U14205 (N_14205,N_11278,N_11031);
and U14206 (N_14206,N_11514,N_10788);
nand U14207 (N_14207,N_11389,N_11338);
xor U14208 (N_14208,N_10084,N_10527);
or U14209 (N_14209,N_11311,N_10717);
and U14210 (N_14210,N_11846,N_11099);
or U14211 (N_14211,N_12191,N_10162);
nor U14212 (N_14212,N_12413,N_11574);
nor U14213 (N_14213,N_11934,N_10268);
and U14214 (N_14214,N_12048,N_10101);
and U14215 (N_14215,N_12199,N_10908);
nor U14216 (N_14216,N_10693,N_11773);
or U14217 (N_14217,N_11092,N_10037);
and U14218 (N_14218,N_10834,N_10207);
or U14219 (N_14219,N_12203,N_10386);
xor U14220 (N_14220,N_10429,N_10324);
nor U14221 (N_14221,N_11645,N_11735);
nand U14222 (N_14222,N_11852,N_11259);
nor U14223 (N_14223,N_12119,N_12474);
xnor U14224 (N_14224,N_12331,N_12181);
xnor U14225 (N_14225,N_11572,N_11196);
nand U14226 (N_14226,N_11653,N_11397);
xnor U14227 (N_14227,N_12269,N_11402);
nor U14228 (N_14228,N_10783,N_10642);
nor U14229 (N_14229,N_11102,N_12315);
nor U14230 (N_14230,N_11772,N_11941);
nor U14231 (N_14231,N_11525,N_12332);
and U14232 (N_14232,N_11467,N_10836);
and U14233 (N_14233,N_11898,N_11742);
and U14234 (N_14234,N_12212,N_11865);
nor U14235 (N_14235,N_10345,N_11804);
xnor U14236 (N_14236,N_10401,N_11811);
xnor U14237 (N_14237,N_11202,N_10553);
xnor U14238 (N_14238,N_11397,N_12395);
nand U14239 (N_14239,N_10113,N_12332);
xnor U14240 (N_14240,N_10535,N_12076);
and U14241 (N_14241,N_10147,N_11025);
xnor U14242 (N_14242,N_11204,N_12070);
nand U14243 (N_14243,N_11374,N_12464);
nand U14244 (N_14244,N_10281,N_11096);
or U14245 (N_14245,N_11563,N_11949);
nor U14246 (N_14246,N_10879,N_10416);
and U14247 (N_14247,N_10742,N_11125);
or U14248 (N_14248,N_10247,N_10350);
and U14249 (N_14249,N_10823,N_11097);
nor U14250 (N_14250,N_10058,N_11609);
and U14251 (N_14251,N_11863,N_11633);
nand U14252 (N_14252,N_12063,N_12198);
nand U14253 (N_14253,N_11359,N_10323);
nor U14254 (N_14254,N_10482,N_11713);
nor U14255 (N_14255,N_10155,N_10087);
or U14256 (N_14256,N_10218,N_12209);
nand U14257 (N_14257,N_11270,N_11054);
nand U14258 (N_14258,N_11384,N_12230);
nor U14259 (N_14259,N_11886,N_11413);
nor U14260 (N_14260,N_12171,N_11358);
or U14261 (N_14261,N_10504,N_10192);
nor U14262 (N_14262,N_12145,N_10052);
or U14263 (N_14263,N_12339,N_11659);
or U14264 (N_14264,N_11098,N_10257);
nor U14265 (N_14265,N_10237,N_11152);
or U14266 (N_14266,N_11346,N_10910);
nand U14267 (N_14267,N_12330,N_10843);
and U14268 (N_14268,N_10980,N_10501);
or U14269 (N_14269,N_12072,N_10919);
nor U14270 (N_14270,N_11228,N_11045);
nor U14271 (N_14271,N_10469,N_11072);
nand U14272 (N_14272,N_10114,N_11291);
nor U14273 (N_14273,N_11442,N_12350);
xnor U14274 (N_14274,N_12273,N_12328);
nand U14275 (N_14275,N_11413,N_10680);
nor U14276 (N_14276,N_11851,N_12448);
and U14277 (N_14277,N_11093,N_10135);
or U14278 (N_14278,N_10811,N_10415);
and U14279 (N_14279,N_11825,N_11963);
xnor U14280 (N_14280,N_10183,N_11291);
or U14281 (N_14281,N_11535,N_10315);
nand U14282 (N_14282,N_11962,N_11492);
xor U14283 (N_14283,N_11207,N_10947);
or U14284 (N_14284,N_11132,N_12249);
nor U14285 (N_14285,N_10755,N_11595);
xor U14286 (N_14286,N_10124,N_11709);
nor U14287 (N_14287,N_11395,N_11520);
and U14288 (N_14288,N_10461,N_11214);
nand U14289 (N_14289,N_11798,N_11206);
or U14290 (N_14290,N_10737,N_11944);
and U14291 (N_14291,N_10901,N_12401);
nor U14292 (N_14292,N_11598,N_11051);
and U14293 (N_14293,N_10952,N_10777);
nor U14294 (N_14294,N_11371,N_10899);
nor U14295 (N_14295,N_11270,N_11047);
xnor U14296 (N_14296,N_11914,N_12413);
or U14297 (N_14297,N_12266,N_12312);
xnor U14298 (N_14298,N_10844,N_11656);
nor U14299 (N_14299,N_10306,N_10384);
xor U14300 (N_14300,N_12372,N_10273);
or U14301 (N_14301,N_10906,N_10417);
nand U14302 (N_14302,N_10706,N_12312);
nor U14303 (N_14303,N_12066,N_10001);
or U14304 (N_14304,N_12289,N_11089);
or U14305 (N_14305,N_10211,N_10731);
and U14306 (N_14306,N_11891,N_10728);
xor U14307 (N_14307,N_11800,N_10576);
nand U14308 (N_14308,N_10454,N_10347);
nor U14309 (N_14309,N_11947,N_12039);
xor U14310 (N_14310,N_10218,N_11419);
or U14311 (N_14311,N_10301,N_11573);
nand U14312 (N_14312,N_10039,N_10019);
and U14313 (N_14313,N_10147,N_11999);
xnor U14314 (N_14314,N_10847,N_11393);
or U14315 (N_14315,N_12139,N_11690);
nand U14316 (N_14316,N_11881,N_11215);
xnor U14317 (N_14317,N_10981,N_11742);
xor U14318 (N_14318,N_12317,N_10089);
nand U14319 (N_14319,N_10125,N_11738);
nor U14320 (N_14320,N_10347,N_12250);
xor U14321 (N_14321,N_11449,N_11606);
and U14322 (N_14322,N_10562,N_10622);
nor U14323 (N_14323,N_11113,N_10009);
xor U14324 (N_14324,N_12370,N_10045);
and U14325 (N_14325,N_11899,N_11532);
nand U14326 (N_14326,N_10610,N_12353);
nor U14327 (N_14327,N_11020,N_11039);
and U14328 (N_14328,N_10310,N_10969);
xnor U14329 (N_14329,N_11807,N_12038);
nor U14330 (N_14330,N_10598,N_12214);
xor U14331 (N_14331,N_10273,N_12412);
xor U14332 (N_14332,N_11546,N_11766);
nor U14333 (N_14333,N_12427,N_11758);
nor U14334 (N_14334,N_11336,N_11775);
nor U14335 (N_14335,N_11413,N_11595);
or U14336 (N_14336,N_10433,N_11358);
nor U14337 (N_14337,N_11332,N_12162);
xnor U14338 (N_14338,N_10318,N_10487);
nand U14339 (N_14339,N_11728,N_11138);
and U14340 (N_14340,N_12292,N_12237);
or U14341 (N_14341,N_11727,N_10100);
or U14342 (N_14342,N_10138,N_11204);
nand U14343 (N_14343,N_12306,N_12011);
and U14344 (N_14344,N_12407,N_11590);
nand U14345 (N_14345,N_12170,N_10372);
nor U14346 (N_14346,N_11182,N_11150);
nand U14347 (N_14347,N_10305,N_10736);
or U14348 (N_14348,N_10836,N_11024);
nor U14349 (N_14349,N_12330,N_10311);
nor U14350 (N_14350,N_10725,N_12163);
nand U14351 (N_14351,N_10477,N_11749);
nand U14352 (N_14352,N_11355,N_11870);
nor U14353 (N_14353,N_12400,N_10020);
nor U14354 (N_14354,N_10494,N_11855);
and U14355 (N_14355,N_11386,N_10176);
xnor U14356 (N_14356,N_11307,N_10678);
and U14357 (N_14357,N_10521,N_12065);
nor U14358 (N_14358,N_10838,N_11854);
or U14359 (N_14359,N_12391,N_12214);
or U14360 (N_14360,N_12096,N_12093);
nand U14361 (N_14361,N_10613,N_12015);
nand U14362 (N_14362,N_12363,N_10203);
xor U14363 (N_14363,N_11801,N_11937);
and U14364 (N_14364,N_12411,N_11907);
xor U14365 (N_14365,N_11758,N_12442);
nand U14366 (N_14366,N_11331,N_11643);
or U14367 (N_14367,N_11974,N_11610);
or U14368 (N_14368,N_10618,N_11647);
nand U14369 (N_14369,N_10110,N_10867);
nand U14370 (N_14370,N_10566,N_10066);
nand U14371 (N_14371,N_10176,N_11922);
and U14372 (N_14372,N_11655,N_11886);
nor U14373 (N_14373,N_10965,N_12269);
xor U14374 (N_14374,N_10710,N_12400);
nand U14375 (N_14375,N_11802,N_11981);
xnor U14376 (N_14376,N_10831,N_11966);
and U14377 (N_14377,N_11571,N_10155);
nand U14378 (N_14378,N_10584,N_11360);
or U14379 (N_14379,N_10480,N_11461);
nor U14380 (N_14380,N_12206,N_10111);
nand U14381 (N_14381,N_10598,N_10197);
xnor U14382 (N_14382,N_12214,N_12088);
or U14383 (N_14383,N_12302,N_10984);
and U14384 (N_14384,N_11941,N_10331);
or U14385 (N_14385,N_11752,N_11740);
and U14386 (N_14386,N_12299,N_11333);
and U14387 (N_14387,N_12479,N_11968);
nor U14388 (N_14388,N_10542,N_10204);
xor U14389 (N_14389,N_11262,N_10552);
or U14390 (N_14390,N_10256,N_10399);
xor U14391 (N_14391,N_11705,N_11632);
nor U14392 (N_14392,N_11762,N_11838);
nand U14393 (N_14393,N_12418,N_11460);
nand U14394 (N_14394,N_11365,N_11494);
or U14395 (N_14395,N_10436,N_12018);
or U14396 (N_14396,N_12457,N_10871);
nor U14397 (N_14397,N_10601,N_11991);
or U14398 (N_14398,N_10367,N_11352);
nor U14399 (N_14399,N_11745,N_12001);
nor U14400 (N_14400,N_11314,N_12062);
nor U14401 (N_14401,N_11619,N_10090);
xor U14402 (N_14402,N_11758,N_10026);
nand U14403 (N_14403,N_10367,N_10295);
or U14404 (N_14404,N_10522,N_12458);
nand U14405 (N_14405,N_11087,N_10205);
or U14406 (N_14406,N_11159,N_11072);
or U14407 (N_14407,N_10847,N_11424);
and U14408 (N_14408,N_11525,N_10886);
nand U14409 (N_14409,N_12343,N_11001);
or U14410 (N_14410,N_10287,N_12414);
xnor U14411 (N_14411,N_10708,N_11384);
and U14412 (N_14412,N_12165,N_10071);
and U14413 (N_14413,N_10555,N_11080);
nand U14414 (N_14414,N_11381,N_10299);
and U14415 (N_14415,N_11063,N_10272);
xor U14416 (N_14416,N_11495,N_11175);
nand U14417 (N_14417,N_11679,N_11618);
or U14418 (N_14418,N_12045,N_10263);
nand U14419 (N_14419,N_11545,N_10433);
or U14420 (N_14420,N_11778,N_11172);
and U14421 (N_14421,N_10899,N_10520);
nand U14422 (N_14422,N_10988,N_10708);
or U14423 (N_14423,N_10297,N_10894);
nand U14424 (N_14424,N_11522,N_11914);
or U14425 (N_14425,N_12307,N_11486);
or U14426 (N_14426,N_11700,N_11138);
and U14427 (N_14427,N_11824,N_10743);
nor U14428 (N_14428,N_11745,N_11177);
xnor U14429 (N_14429,N_11416,N_11215);
xor U14430 (N_14430,N_12118,N_10640);
xor U14431 (N_14431,N_12358,N_12480);
or U14432 (N_14432,N_10006,N_10654);
nor U14433 (N_14433,N_10595,N_11822);
nor U14434 (N_14434,N_11049,N_11191);
and U14435 (N_14435,N_10505,N_11472);
nand U14436 (N_14436,N_10517,N_11048);
nand U14437 (N_14437,N_10545,N_11307);
nand U14438 (N_14438,N_10858,N_10496);
or U14439 (N_14439,N_11347,N_11115);
or U14440 (N_14440,N_10449,N_10320);
xnor U14441 (N_14441,N_11524,N_12483);
xnor U14442 (N_14442,N_11437,N_12309);
nand U14443 (N_14443,N_11725,N_10910);
nand U14444 (N_14444,N_11191,N_11216);
and U14445 (N_14445,N_11582,N_11951);
nor U14446 (N_14446,N_10641,N_12036);
and U14447 (N_14447,N_11949,N_10336);
nor U14448 (N_14448,N_12330,N_11085);
and U14449 (N_14449,N_12246,N_10126);
and U14450 (N_14450,N_12464,N_11514);
nor U14451 (N_14451,N_10347,N_10467);
and U14452 (N_14452,N_10046,N_11941);
xnor U14453 (N_14453,N_11011,N_12349);
or U14454 (N_14454,N_11992,N_12445);
and U14455 (N_14455,N_10561,N_10129);
nand U14456 (N_14456,N_10978,N_10811);
or U14457 (N_14457,N_10980,N_12389);
or U14458 (N_14458,N_12075,N_11640);
nand U14459 (N_14459,N_11559,N_10529);
and U14460 (N_14460,N_10567,N_11149);
or U14461 (N_14461,N_10389,N_10362);
or U14462 (N_14462,N_11710,N_10862);
nor U14463 (N_14463,N_11287,N_10140);
or U14464 (N_14464,N_11832,N_11741);
or U14465 (N_14465,N_12495,N_12000);
nand U14466 (N_14466,N_11140,N_12069);
nand U14467 (N_14467,N_10628,N_10583);
xor U14468 (N_14468,N_11755,N_12488);
or U14469 (N_14469,N_10155,N_11508);
or U14470 (N_14470,N_12401,N_10430);
and U14471 (N_14471,N_11056,N_11152);
and U14472 (N_14472,N_12248,N_10548);
or U14473 (N_14473,N_10148,N_10629);
nor U14474 (N_14474,N_12392,N_10338);
or U14475 (N_14475,N_11886,N_12138);
nor U14476 (N_14476,N_11734,N_10592);
nor U14477 (N_14477,N_12059,N_10612);
xor U14478 (N_14478,N_10977,N_12106);
xnor U14479 (N_14479,N_11485,N_12148);
and U14480 (N_14480,N_10432,N_10966);
nor U14481 (N_14481,N_11396,N_11389);
nor U14482 (N_14482,N_11999,N_11055);
nor U14483 (N_14483,N_10514,N_10057);
or U14484 (N_14484,N_10825,N_10948);
or U14485 (N_14485,N_11523,N_11613);
nand U14486 (N_14486,N_10080,N_10751);
and U14487 (N_14487,N_11992,N_12039);
nand U14488 (N_14488,N_10386,N_11741);
xor U14489 (N_14489,N_10637,N_12218);
and U14490 (N_14490,N_12127,N_11225);
or U14491 (N_14491,N_10552,N_11202);
and U14492 (N_14492,N_10774,N_11131);
xor U14493 (N_14493,N_11440,N_10969);
and U14494 (N_14494,N_10394,N_11684);
and U14495 (N_14495,N_11990,N_11897);
nor U14496 (N_14496,N_11815,N_10693);
xor U14497 (N_14497,N_12376,N_11549);
nand U14498 (N_14498,N_10010,N_11145);
or U14499 (N_14499,N_10858,N_12113);
or U14500 (N_14500,N_12434,N_10420);
and U14501 (N_14501,N_10828,N_10971);
or U14502 (N_14502,N_10820,N_10506);
and U14503 (N_14503,N_10425,N_11169);
nand U14504 (N_14504,N_11472,N_11153);
and U14505 (N_14505,N_10811,N_10060);
xnor U14506 (N_14506,N_11851,N_11843);
nor U14507 (N_14507,N_11042,N_11021);
nand U14508 (N_14508,N_10582,N_11186);
and U14509 (N_14509,N_10350,N_12231);
and U14510 (N_14510,N_10342,N_12435);
and U14511 (N_14511,N_11832,N_10727);
nor U14512 (N_14512,N_12369,N_11466);
or U14513 (N_14513,N_12347,N_12273);
or U14514 (N_14514,N_10226,N_12274);
nand U14515 (N_14515,N_12155,N_11815);
and U14516 (N_14516,N_10483,N_10560);
or U14517 (N_14517,N_10849,N_11663);
xor U14518 (N_14518,N_10320,N_11244);
xnor U14519 (N_14519,N_11788,N_10056);
nand U14520 (N_14520,N_11733,N_10726);
and U14521 (N_14521,N_11013,N_11699);
nand U14522 (N_14522,N_11605,N_11597);
or U14523 (N_14523,N_10327,N_10073);
or U14524 (N_14524,N_10366,N_10072);
and U14525 (N_14525,N_11782,N_11316);
or U14526 (N_14526,N_11033,N_11315);
nand U14527 (N_14527,N_12459,N_12223);
nor U14528 (N_14528,N_10986,N_10657);
nand U14529 (N_14529,N_12170,N_11308);
and U14530 (N_14530,N_10484,N_10591);
or U14531 (N_14531,N_10483,N_11292);
and U14532 (N_14532,N_12071,N_12437);
nand U14533 (N_14533,N_10536,N_10730);
or U14534 (N_14534,N_11259,N_10658);
xor U14535 (N_14535,N_10474,N_11711);
nor U14536 (N_14536,N_11018,N_11867);
xnor U14537 (N_14537,N_10581,N_12408);
nand U14538 (N_14538,N_10025,N_11145);
xor U14539 (N_14539,N_10330,N_10167);
nand U14540 (N_14540,N_11524,N_12022);
nor U14541 (N_14541,N_11469,N_10621);
xor U14542 (N_14542,N_11852,N_12317);
and U14543 (N_14543,N_11170,N_10451);
nor U14544 (N_14544,N_10616,N_10071);
nand U14545 (N_14545,N_11488,N_11305);
xor U14546 (N_14546,N_10497,N_11224);
nor U14547 (N_14547,N_11859,N_11431);
and U14548 (N_14548,N_12358,N_11711);
nor U14549 (N_14549,N_10314,N_12471);
nor U14550 (N_14550,N_12049,N_11157);
and U14551 (N_14551,N_10584,N_12287);
nor U14552 (N_14552,N_12431,N_12412);
and U14553 (N_14553,N_10159,N_10503);
xor U14554 (N_14554,N_12366,N_10993);
xor U14555 (N_14555,N_11366,N_10038);
and U14556 (N_14556,N_11257,N_11942);
and U14557 (N_14557,N_10127,N_11592);
nor U14558 (N_14558,N_11326,N_10546);
or U14559 (N_14559,N_11429,N_11518);
xor U14560 (N_14560,N_11961,N_10549);
nand U14561 (N_14561,N_12207,N_10070);
nor U14562 (N_14562,N_10651,N_10683);
nand U14563 (N_14563,N_11642,N_11702);
nor U14564 (N_14564,N_11201,N_11859);
and U14565 (N_14565,N_12378,N_11858);
xnor U14566 (N_14566,N_12038,N_10140);
or U14567 (N_14567,N_10061,N_11156);
and U14568 (N_14568,N_10991,N_11097);
or U14569 (N_14569,N_11742,N_11737);
and U14570 (N_14570,N_12417,N_12386);
nor U14571 (N_14571,N_10385,N_12002);
nand U14572 (N_14572,N_12403,N_11795);
nor U14573 (N_14573,N_11756,N_11562);
or U14574 (N_14574,N_10519,N_11284);
nor U14575 (N_14575,N_12403,N_10623);
nand U14576 (N_14576,N_10690,N_11355);
xor U14577 (N_14577,N_12044,N_11902);
nand U14578 (N_14578,N_10380,N_11175);
and U14579 (N_14579,N_11641,N_11172);
and U14580 (N_14580,N_12054,N_11508);
or U14581 (N_14581,N_11874,N_12324);
or U14582 (N_14582,N_12271,N_11781);
xor U14583 (N_14583,N_10070,N_10167);
nand U14584 (N_14584,N_11225,N_11753);
and U14585 (N_14585,N_11231,N_11258);
or U14586 (N_14586,N_10064,N_11962);
xnor U14587 (N_14587,N_11508,N_10368);
and U14588 (N_14588,N_10548,N_10089);
or U14589 (N_14589,N_10887,N_11419);
nor U14590 (N_14590,N_11072,N_11507);
xor U14591 (N_14591,N_11624,N_12047);
and U14592 (N_14592,N_10179,N_12403);
nand U14593 (N_14593,N_11420,N_11408);
and U14594 (N_14594,N_11665,N_10824);
or U14595 (N_14595,N_11941,N_11448);
nand U14596 (N_14596,N_12129,N_10884);
or U14597 (N_14597,N_12322,N_11128);
nor U14598 (N_14598,N_10328,N_11312);
or U14599 (N_14599,N_10426,N_11067);
and U14600 (N_14600,N_11617,N_11815);
nand U14601 (N_14601,N_10042,N_11568);
xor U14602 (N_14602,N_10775,N_12368);
nand U14603 (N_14603,N_11360,N_12268);
nor U14604 (N_14604,N_11989,N_10027);
and U14605 (N_14605,N_12386,N_10292);
nand U14606 (N_14606,N_12440,N_12240);
and U14607 (N_14607,N_10753,N_11239);
nand U14608 (N_14608,N_10667,N_10368);
or U14609 (N_14609,N_11355,N_10419);
or U14610 (N_14610,N_11428,N_11099);
nor U14611 (N_14611,N_10198,N_12261);
nor U14612 (N_14612,N_11290,N_10281);
or U14613 (N_14613,N_10240,N_10773);
xnor U14614 (N_14614,N_11690,N_11158);
nand U14615 (N_14615,N_12250,N_11982);
and U14616 (N_14616,N_11096,N_11835);
and U14617 (N_14617,N_11867,N_12327);
nand U14618 (N_14618,N_11635,N_10724);
nor U14619 (N_14619,N_11285,N_10551);
nand U14620 (N_14620,N_10722,N_11522);
nor U14621 (N_14621,N_11245,N_11758);
or U14622 (N_14622,N_11529,N_11828);
and U14623 (N_14623,N_11930,N_12464);
nor U14624 (N_14624,N_11158,N_11520);
and U14625 (N_14625,N_10875,N_10793);
or U14626 (N_14626,N_10650,N_11506);
xor U14627 (N_14627,N_10639,N_10941);
nand U14628 (N_14628,N_12442,N_11046);
nand U14629 (N_14629,N_11526,N_10546);
and U14630 (N_14630,N_10255,N_12093);
xor U14631 (N_14631,N_10772,N_11928);
or U14632 (N_14632,N_10796,N_10062);
and U14633 (N_14633,N_10344,N_10778);
and U14634 (N_14634,N_11433,N_11560);
nand U14635 (N_14635,N_10198,N_11849);
or U14636 (N_14636,N_10019,N_11600);
and U14637 (N_14637,N_11813,N_12117);
nand U14638 (N_14638,N_10889,N_11936);
or U14639 (N_14639,N_11093,N_11492);
xnor U14640 (N_14640,N_12416,N_10984);
nand U14641 (N_14641,N_10293,N_11350);
xnor U14642 (N_14642,N_11164,N_10387);
nand U14643 (N_14643,N_12415,N_11697);
and U14644 (N_14644,N_11913,N_12472);
nand U14645 (N_14645,N_11979,N_10330);
nand U14646 (N_14646,N_12008,N_10378);
xor U14647 (N_14647,N_12343,N_11026);
nand U14648 (N_14648,N_10348,N_10337);
xor U14649 (N_14649,N_10555,N_11425);
nand U14650 (N_14650,N_10004,N_10236);
and U14651 (N_14651,N_10837,N_11407);
or U14652 (N_14652,N_11898,N_12015);
nor U14653 (N_14653,N_10619,N_11030);
nor U14654 (N_14654,N_10459,N_10728);
xnor U14655 (N_14655,N_12078,N_11609);
nor U14656 (N_14656,N_10345,N_10437);
xor U14657 (N_14657,N_10884,N_10874);
or U14658 (N_14658,N_10527,N_11190);
xnor U14659 (N_14659,N_12296,N_11358);
nor U14660 (N_14660,N_10472,N_11056);
nand U14661 (N_14661,N_12206,N_11439);
or U14662 (N_14662,N_12457,N_10296);
nand U14663 (N_14663,N_10773,N_11897);
and U14664 (N_14664,N_10252,N_11075);
or U14665 (N_14665,N_11044,N_12120);
xor U14666 (N_14666,N_11622,N_10025);
and U14667 (N_14667,N_11398,N_10262);
nand U14668 (N_14668,N_11901,N_11956);
nand U14669 (N_14669,N_11704,N_10040);
and U14670 (N_14670,N_10993,N_11369);
and U14671 (N_14671,N_11312,N_11356);
or U14672 (N_14672,N_10456,N_10918);
nor U14673 (N_14673,N_10917,N_10180);
xor U14674 (N_14674,N_10080,N_10354);
nor U14675 (N_14675,N_11803,N_10141);
and U14676 (N_14676,N_11827,N_12347);
or U14677 (N_14677,N_10633,N_10900);
nand U14678 (N_14678,N_10512,N_10736);
xnor U14679 (N_14679,N_11697,N_10225);
nor U14680 (N_14680,N_10630,N_10741);
nand U14681 (N_14681,N_12226,N_11307);
nand U14682 (N_14682,N_11943,N_10393);
or U14683 (N_14683,N_10769,N_10733);
nand U14684 (N_14684,N_10611,N_12430);
xnor U14685 (N_14685,N_12105,N_10505);
or U14686 (N_14686,N_10683,N_10894);
xnor U14687 (N_14687,N_12101,N_10752);
nand U14688 (N_14688,N_10142,N_10557);
nor U14689 (N_14689,N_10867,N_11690);
nor U14690 (N_14690,N_11331,N_10545);
or U14691 (N_14691,N_10002,N_12250);
nor U14692 (N_14692,N_11594,N_11221);
and U14693 (N_14693,N_10419,N_12353);
or U14694 (N_14694,N_10249,N_12169);
nand U14695 (N_14695,N_11424,N_12386);
nand U14696 (N_14696,N_12113,N_10666);
nand U14697 (N_14697,N_11000,N_11516);
nand U14698 (N_14698,N_10563,N_11712);
xor U14699 (N_14699,N_10548,N_11672);
or U14700 (N_14700,N_10954,N_12213);
or U14701 (N_14701,N_11853,N_10833);
xnor U14702 (N_14702,N_10598,N_10577);
and U14703 (N_14703,N_11553,N_11296);
and U14704 (N_14704,N_12358,N_12207);
nand U14705 (N_14705,N_10885,N_12230);
and U14706 (N_14706,N_11889,N_12239);
and U14707 (N_14707,N_10143,N_10795);
nor U14708 (N_14708,N_10427,N_11745);
and U14709 (N_14709,N_11371,N_10876);
xnor U14710 (N_14710,N_11453,N_11566);
nor U14711 (N_14711,N_11665,N_11157);
and U14712 (N_14712,N_11345,N_10932);
xnor U14713 (N_14713,N_10251,N_10953);
nand U14714 (N_14714,N_11313,N_11977);
or U14715 (N_14715,N_12249,N_10136);
nand U14716 (N_14716,N_10421,N_12215);
xnor U14717 (N_14717,N_12493,N_10173);
nand U14718 (N_14718,N_10113,N_11582);
xor U14719 (N_14719,N_11441,N_12380);
and U14720 (N_14720,N_10479,N_12120);
nor U14721 (N_14721,N_10160,N_10321);
xor U14722 (N_14722,N_10981,N_11146);
nand U14723 (N_14723,N_11030,N_11902);
and U14724 (N_14724,N_10280,N_11009);
nand U14725 (N_14725,N_11259,N_11284);
nor U14726 (N_14726,N_10357,N_10691);
nor U14727 (N_14727,N_11499,N_11221);
or U14728 (N_14728,N_10639,N_11785);
or U14729 (N_14729,N_11407,N_11812);
and U14730 (N_14730,N_12429,N_11008);
nor U14731 (N_14731,N_10432,N_12106);
nor U14732 (N_14732,N_11619,N_12283);
or U14733 (N_14733,N_10016,N_11775);
or U14734 (N_14734,N_10505,N_12116);
xnor U14735 (N_14735,N_11233,N_10240);
and U14736 (N_14736,N_10121,N_10262);
xor U14737 (N_14737,N_12433,N_12034);
nor U14738 (N_14738,N_11534,N_12021);
nand U14739 (N_14739,N_11171,N_11757);
or U14740 (N_14740,N_11275,N_12041);
and U14741 (N_14741,N_12015,N_12282);
nand U14742 (N_14742,N_10011,N_10774);
xnor U14743 (N_14743,N_10744,N_10748);
nand U14744 (N_14744,N_10966,N_10361);
nand U14745 (N_14745,N_11854,N_12266);
and U14746 (N_14746,N_12094,N_12424);
and U14747 (N_14747,N_10501,N_11487);
and U14748 (N_14748,N_10481,N_10385);
and U14749 (N_14749,N_11276,N_11381);
xnor U14750 (N_14750,N_10116,N_10767);
or U14751 (N_14751,N_12384,N_12216);
and U14752 (N_14752,N_11626,N_11160);
xnor U14753 (N_14753,N_10904,N_12233);
nor U14754 (N_14754,N_11715,N_10165);
and U14755 (N_14755,N_12118,N_11418);
xnor U14756 (N_14756,N_12147,N_10345);
nand U14757 (N_14757,N_11525,N_11826);
and U14758 (N_14758,N_10378,N_12225);
nand U14759 (N_14759,N_11002,N_10192);
or U14760 (N_14760,N_11258,N_12473);
or U14761 (N_14761,N_11363,N_11126);
or U14762 (N_14762,N_12022,N_10346);
nand U14763 (N_14763,N_10235,N_11128);
nand U14764 (N_14764,N_10691,N_10291);
xor U14765 (N_14765,N_11036,N_12003);
xor U14766 (N_14766,N_11044,N_11776);
nor U14767 (N_14767,N_11702,N_11019);
nor U14768 (N_14768,N_10882,N_11769);
nand U14769 (N_14769,N_11215,N_10928);
and U14770 (N_14770,N_11913,N_12018);
and U14771 (N_14771,N_11698,N_10794);
nor U14772 (N_14772,N_12230,N_11507);
nor U14773 (N_14773,N_10000,N_12300);
or U14774 (N_14774,N_12160,N_12333);
nand U14775 (N_14775,N_11189,N_10912);
or U14776 (N_14776,N_11902,N_11799);
xor U14777 (N_14777,N_11708,N_11133);
xnor U14778 (N_14778,N_11796,N_11093);
nor U14779 (N_14779,N_10791,N_11862);
nand U14780 (N_14780,N_10393,N_11283);
and U14781 (N_14781,N_10961,N_11577);
nor U14782 (N_14782,N_12300,N_11305);
and U14783 (N_14783,N_11564,N_10038);
xnor U14784 (N_14784,N_12314,N_11534);
or U14785 (N_14785,N_12460,N_12313);
nor U14786 (N_14786,N_11878,N_11200);
nand U14787 (N_14787,N_12076,N_12499);
nor U14788 (N_14788,N_10489,N_11612);
nand U14789 (N_14789,N_10706,N_12238);
nand U14790 (N_14790,N_10772,N_12239);
xor U14791 (N_14791,N_12260,N_11385);
or U14792 (N_14792,N_10590,N_10271);
xnor U14793 (N_14793,N_10340,N_10441);
nand U14794 (N_14794,N_11898,N_10754);
and U14795 (N_14795,N_11155,N_11878);
and U14796 (N_14796,N_10516,N_11698);
or U14797 (N_14797,N_11967,N_11617);
or U14798 (N_14798,N_10051,N_12236);
nor U14799 (N_14799,N_12133,N_10086);
and U14800 (N_14800,N_12442,N_10488);
nor U14801 (N_14801,N_11893,N_10196);
or U14802 (N_14802,N_10890,N_10777);
nand U14803 (N_14803,N_11334,N_12134);
and U14804 (N_14804,N_10750,N_12097);
xor U14805 (N_14805,N_11176,N_10224);
xor U14806 (N_14806,N_11603,N_11860);
xor U14807 (N_14807,N_11384,N_11679);
nand U14808 (N_14808,N_12245,N_10479);
nand U14809 (N_14809,N_10775,N_10281);
xnor U14810 (N_14810,N_11028,N_10732);
xor U14811 (N_14811,N_11439,N_11472);
xnor U14812 (N_14812,N_12321,N_10437);
nor U14813 (N_14813,N_12204,N_10787);
or U14814 (N_14814,N_11558,N_11655);
nand U14815 (N_14815,N_10879,N_12256);
nor U14816 (N_14816,N_11625,N_10647);
nand U14817 (N_14817,N_11218,N_12351);
and U14818 (N_14818,N_10709,N_10833);
nand U14819 (N_14819,N_10151,N_10800);
or U14820 (N_14820,N_12006,N_10174);
xor U14821 (N_14821,N_12081,N_11552);
and U14822 (N_14822,N_10388,N_11031);
or U14823 (N_14823,N_12108,N_11008);
and U14824 (N_14824,N_12425,N_11904);
or U14825 (N_14825,N_11052,N_10811);
or U14826 (N_14826,N_12380,N_10127);
nor U14827 (N_14827,N_11091,N_10542);
or U14828 (N_14828,N_10725,N_10064);
nor U14829 (N_14829,N_11014,N_12440);
nor U14830 (N_14830,N_11197,N_10145);
nor U14831 (N_14831,N_11126,N_10433);
nor U14832 (N_14832,N_10028,N_12238);
or U14833 (N_14833,N_10794,N_11598);
xnor U14834 (N_14834,N_11748,N_10308);
nand U14835 (N_14835,N_10696,N_11524);
xnor U14836 (N_14836,N_10481,N_11174);
xor U14837 (N_14837,N_10885,N_11978);
nor U14838 (N_14838,N_11392,N_11181);
nor U14839 (N_14839,N_10822,N_11838);
nor U14840 (N_14840,N_11267,N_12208);
xor U14841 (N_14841,N_11306,N_10754);
and U14842 (N_14842,N_12063,N_10691);
or U14843 (N_14843,N_11879,N_11247);
xnor U14844 (N_14844,N_11221,N_10481);
nor U14845 (N_14845,N_11257,N_11255);
nand U14846 (N_14846,N_10440,N_12169);
or U14847 (N_14847,N_10044,N_11890);
and U14848 (N_14848,N_12172,N_10081);
or U14849 (N_14849,N_11228,N_11803);
nand U14850 (N_14850,N_11272,N_10512);
xor U14851 (N_14851,N_11382,N_11818);
or U14852 (N_14852,N_11520,N_12434);
nand U14853 (N_14853,N_11522,N_11838);
and U14854 (N_14854,N_12296,N_11132);
and U14855 (N_14855,N_10640,N_10172);
nor U14856 (N_14856,N_10602,N_10429);
and U14857 (N_14857,N_11965,N_10216);
nand U14858 (N_14858,N_11648,N_10357);
nand U14859 (N_14859,N_11653,N_12046);
xnor U14860 (N_14860,N_10826,N_10494);
xor U14861 (N_14861,N_10461,N_10494);
or U14862 (N_14862,N_10016,N_11990);
and U14863 (N_14863,N_11336,N_12304);
or U14864 (N_14864,N_11230,N_11268);
xor U14865 (N_14865,N_12376,N_11047);
nor U14866 (N_14866,N_10932,N_10311);
nand U14867 (N_14867,N_10601,N_11809);
nand U14868 (N_14868,N_10501,N_11212);
nand U14869 (N_14869,N_10204,N_12157);
xor U14870 (N_14870,N_10190,N_10888);
and U14871 (N_14871,N_10535,N_12264);
nor U14872 (N_14872,N_10372,N_11274);
nor U14873 (N_14873,N_12007,N_11435);
and U14874 (N_14874,N_11060,N_10397);
xnor U14875 (N_14875,N_12336,N_10276);
or U14876 (N_14876,N_10016,N_11409);
xor U14877 (N_14877,N_11718,N_11945);
nor U14878 (N_14878,N_11434,N_11279);
nor U14879 (N_14879,N_11069,N_11275);
or U14880 (N_14880,N_11185,N_10743);
nand U14881 (N_14881,N_10752,N_10263);
and U14882 (N_14882,N_11566,N_12233);
or U14883 (N_14883,N_10241,N_11564);
or U14884 (N_14884,N_10038,N_12114);
xnor U14885 (N_14885,N_11328,N_10977);
and U14886 (N_14886,N_10031,N_11119);
xor U14887 (N_14887,N_11670,N_10404);
and U14888 (N_14888,N_10214,N_11970);
xor U14889 (N_14889,N_10286,N_10307);
nand U14890 (N_14890,N_10403,N_11570);
or U14891 (N_14891,N_10648,N_11340);
nor U14892 (N_14892,N_11047,N_11173);
nor U14893 (N_14893,N_10936,N_10840);
xnor U14894 (N_14894,N_10453,N_12287);
nand U14895 (N_14895,N_10347,N_11090);
or U14896 (N_14896,N_10642,N_10207);
or U14897 (N_14897,N_10906,N_10326);
or U14898 (N_14898,N_12186,N_10473);
and U14899 (N_14899,N_12434,N_11717);
or U14900 (N_14900,N_11716,N_11759);
nor U14901 (N_14901,N_10955,N_12308);
xor U14902 (N_14902,N_11506,N_10458);
xor U14903 (N_14903,N_11245,N_10551);
nor U14904 (N_14904,N_10814,N_11512);
and U14905 (N_14905,N_10313,N_11497);
xor U14906 (N_14906,N_10139,N_11431);
or U14907 (N_14907,N_11217,N_12379);
nand U14908 (N_14908,N_10324,N_10950);
xor U14909 (N_14909,N_11188,N_11879);
and U14910 (N_14910,N_10560,N_12288);
xor U14911 (N_14911,N_11266,N_11931);
nor U14912 (N_14912,N_10957,N_11005);
xor U14913 (N_14913,N_12003,N_12352);
xor U14914 (N_14914,N_10907,N_12342);
xor U14915 (N_14915,N_11274,N_11191);
and U14916 (N_14916,N_11657,N_12192);
xnor U14917 (N_14917,N_10648,N_11137);
nand U14918 (N_14918,N_11629,N_11528);
or U14919 (N_14919,N_11931,N_10711);
xnor U14920 (N_14920,N_11324,N_12195);
nor U14921 (N_14921,N_10091,N_12455);
or U14922 (N_14922,N_11845,N_10730);
nand U14923 (N_14923,N_11404,N_11553);
xor U14924 (N_14924,N_11092,N_11245);
and U14925 (N_14925,N_11376,N_12275);
nor U14926 (N_14926,N_10592,N_10023);
nor U14927 (N_14927,N_11268,N_12147);
nand U14928 (N_14928,N_11880,N_11125);
or U14929 (N_14929,N_12265,N_10764);
and U14930 (N_14930,N_11160,N_12241);
or U14931 (N_14931,N_12445,N_12303);
nand U14932 (N_14932,N_10989,N_10160);
nor U14933 (N_14933,N_10147,N_10012);
nand U14934 (N_14934,N_12240,N_11682);
xor U14935 (N_14935,N_10378,N_12180);
or U14936 (N_14936,N_11541,N_11686);
xnor U14937 (N_14937,N_12497,N_11459);
and U14938 (N_14938,N_12006,N_11097);
xor U14939 (N_14939,N_11932,N_10770);
nor U14940 (N_14940,N_10295,N_11402);
or U14941 (N_14941,N_10222,N_10668);
or U14942 (N_14942,N_10351,N_12129);
nor U14943 (N_14943,N_12477,N_10301);
nand U14944 (N_14944,N_11781,N_12165);
and U14945 (N_14945,N_11735,N_10721);
and U14946 (N_14946,N_10607,N_11409);
nor U14947 (N_14947,N_11312,N_12473);
nand U14948 (N_14948,N_11165,N_11139);
xor U14949 (N_14949,N_10327,N_10610);
nand U14950 (N_14950,N_10161,N_11660);
and U14951 (N_14951,N_12159,N_11487);
nand U14952 (N_14952,N_11804,N_10817);
or U14953 (N_14953,N_11993,N_11042);
xnor U14954 (N_14954,N_11652,N_10881);
or U14955 (N_14955,N_11635,N_11074);
and U14956 (N_14956,N_11111,N_11521);
and U14957 (N_14957,N_10667,N_10459);
xor U14958 (N_14958,N_10054,N_11033);
nor U14959 (N_14959,N_10623,N_10230);
xor U14960 (N_14960,N_12064,N_10903);
and U14961 (N_14961,N_10219,N_12126);
or U14962 (N_14962,N_12011,N_10547);
or U14963 (N_14963,N_10436,N_10334);
and U14964 (N_14964,N_12237,N_12130);
xnor U14965 (N_14965,N_12058,N_10401);
xnor U14966 (N_14966,N_10691,N_12014);
and U14967 (N_14967,N_12129,N_10304);
xor U14968 (N_14968,N_12384,N_10732);
xor U14969 (N_14969,N_11422,N_12169);
and U14970 (N_14970,N_12193,N_11330);
nor U14971 (N_14971,N_12489,N_12352);
or U14972 (N_14972,N_11197,N_11043);
or U14973 (N_14973,N_11436,N_10355);
and U14974 (N_14974,N_12010,N_10928);
or U14975 (N_14975,N_11541,N_10855);
nor U14976 (N_14976,N_10014,N_10641);
xor U14977 (N_14977,N_12474,N_11573);
nand U14978 (N_14978,N_12337,N_11258);
or U14979 (N_14979,N_11258,N_12351);
nand U14980 (N_14980,N_10025,N_11656);
nand U14981 (N_14981,N_11040,N_11211);
nor U14982 (N_14982,N_10846,N_11384);
nand U14983 (N_14983,N_10611,N_11639);
nand U14984 (N_14984,N_10903,N_11724);
nor U14985 (N_14985,N_11697,N_10181);
xor U14986 (N_14986,N_10999,N_10553);
nand U14987 (N_14987,N_10347,N_10505);
xor U14988 (N_14988,N_10516,N_12412);
or U14989 (N_14989,N_11294,N_10103);
and U14990 (N_14990,N_11836,N_11613);
and U14991 (N_14991,N_11240,N_12163);
xnor U14992 (N_14992,N_12282,N_10131);
nand U14993 (N_14993,N_11366,N_10218);
and U14994 (N_14994,N_11163,N_10256);
nor U14995 (N_14995,N_11226,N_11577);
nor U14996 (N_14996,N_11920,N_12290);
or U14997 (N_14997,N_11437,N_10055);
and U14998 (N_14998,N_11135,N_10158);
nor U14999 (N_14999,N_11689,N_10593);
or U15000 (N_15000,N_13933,N_14045);
nand U15001 (N_15001,N_14657,N_14990);
nor U15002 (N_15002,N_13668,N_14528);
xor U15003 (N_15003,N_13011,N_13206);
nand U15004 (N_15004,N_14531,N_13166);
xor U15005 (N_15005,N_13554,N_13303);
or U15006 (N_15006,N_12721,N_13158);
nor U15007 (N_15007,N_13106,N_14593);
xnor U15008 (N_15008,N_14444,N_14893);
and U15009 (N_15009,N_13133,N_14550);
and U15010 (N_15010,N_12867,N_13977);
nand U15011 (N_15011,N_14735,N_12583);
nor U15012 (N_15012,N_13810,N_13054);
nor U15013 (N_15013,N_13617,N_14062);
nor U15014 (N_15014,N_12668,N_14991);
nor U15015 (N_15015,N_14911,N_13837);
nor U15016 (N_15016,N_13586,N_14758);
nor U15017 (N_15017,N_14264,N_13545);
xnor U15018 (N_15018,N_13763,N_14136);
or U15019 (N_15019,N_14914,N_13299);
or U15020 (N_15020,N_14708,N_13563);
or U15021 (N_15021,N_13798,N_14071);
xnor U15022 (N_15022,N_13915,N_13677);
xnor U15023 (N_15023,N_14648,N_13832);
xnor U15024 (N_15024,N_14961,N_12679);
nor U15025 (N_15025,N_13698,N_14801);
nor U15026 (N_15026,N_13296,N_13318);
nor U15027 (N_15027,N_14395,N_13196);
or U15028 (N_15028,N_13795,N_13725);
and U15029 (N_15029,N_14995,N_12942);
nor U15030 (N_15030,N_12629,N_12945);
or U15031 (N_15031,N_13050,N_14554);
or U15032 (N_15032,N_13871,N_14213);
nand U15033 (N_15033,N_14085,N_13173);
nor U15034 (N_15034,N_13072,N_14372);
nand U15035 (N_15035,N_12961,N_14051);
xnor U15036 (N_15036,N_13530,N_13777);
or U15037 (N_15037,N_13649,N_14956);
and U15038 (N_15038,N_14788,N_12612);
xor U15039 (N_15039,N_12817,N_12968);
xor U15040 (N_15040,N_13778,N_13161);
nand U15041 (N_15041,N_13457,N_14289);
and U15042 (N_15042,N_13385,N_12815);
nor U15043 (N_15043,N_13217,N_12694);
and U15044 (N_15044,N_13227,N_13250);
xor U15045 (N_15045,N_14934,N_14259);
nand U15046 (N_15046,N_12518,N_14567);
and U15047 (N_15047,N_12785,N_14661);
or U15048 (N_15048,N_14111,N_13621);
or U15049 (N_15049,N_13201,N_13441);
nand U15050 (N_15050,N_13671,N_12911);
xor U15051 (N_15051,N_14297,N_14475);
and U15052 (N_15052,N_14844,N_12673);
nor U15053 (N_15053,N_13297,N_13988);
nand U15054 (N_15054,N_14469,N_14654);
nand U15055 (N_15055,N_14783,N_13784);
xor U15056 (N_15056,N_13485,N_12512);
nor U15057 (N_15057,N_12883,N_13560);
xnor U15058 (N_15058,N_14261,N_13374);
nor U15059 (N_15059,N_14534,N_12969);
xnor U15060 (N_15060,N_12756,N_14782);
nand U15061 (N_15061,N_13138,N_14899);
xor U15062 (N_15062,N_14124,N_14406);
nand U15063 (N_15063,N_12660,N_12597);
nand U15064 (N_15064,N_13680,N_12610);
or U15065 (N_15065,N_13464,N_14964);
or U15066 (N_15066,N_14920,N_12514);
or U15067 (N_15067,N_14631,N_14557);
xnor U15068 (N_15068,N_13010,N_14652);
and U15069 (N_15069,N_14919,N_13127);
or U15070 (N_15070,N_12702,N_14499);
xnor U15071 (N_15071,N_12764,N_14042);
and U15072 (N_15072,N_12591,N_14928);
and U15073 (N_15073,N_14526,N_13371);
nand U15074 (N_15074,N_13802,N_12651);
and U15075 (N_15075,N_14243,N_14702);
nor U15076 (N_15076,N_13404,N_12674);
nand U15077 (N_15077,N_13493,N_13547);
nor U15078 (N_15078,N_13996,N_13288);
or U15079 (N_15079,N_13618,N_13740);
nand U15080 (N_15080,N_12714,N_13867);
nor U15081 (N_15081,N_12749,N_13308);
nor U15082 (N_15082,N_14256,N_14588);
and U15083 (N_15083,N_14460,N_12823);
and U15084 (N_15084,N_13019,N_14755);
nand U15085 (N_15085,N_14330,N_14462);
or U15086 (N_15086,N_14089,N_13407);
xnor U15087 (N_15087,N_14232,N_13278);
nor U15088 (N_15088,N_13035,N_14542);
and U15089 (N_15089,N_14987,N_12520);
or U15090 (N_15090,N_13937,N_14113);
and U15091 (N_15091,N_13681,N_14574);
or U15092 (N_15092,N_14687,N_14388);
xor U15093 (N_15093,N_14457,N_12632);
nor U15094 (N_15094,N_14793,N_12645);
nor U15095 (N_15095,N_12923,N_13842);
nand U15096 (N_15096,N_13809,N_14034);
nor U15097 (N_15097,N_14228,N_13117);
or U15098 (N_15098,N_14117,N_12802);
or U15099 (N_15099,N_13110,N_14699);
xnor U15100 (N_15100,N_14487,N_13269);
nor U15101 (N_15101,N_14484,N_14293);
and U15102 (N_15102,N_13561,N_13350);
xor U15103 (N_15103,N_13957,N_13417);
xor U15104 (N_15104,N_12917,N_14456);
nor U15105 (N_15105,N_13815,N_13902);
or U15106 (N_15106,N_14267,N_12531);
or U15107 (N_15107,N_13116,N_12501);
xnor U15108 (N_15108,N_13222,N_13387);
nand U15109 (N_15109,N_13041,N_14323);
nand U15110 (N_15110,N_14020,N_13767);
nor U15111 (N_15111,N_13914,N_14674);
or U15112 (N_15112,N_13674,N_13616);
and U15113 (N_15113,N_12835,N_12821);
nor U15114 (N_15114,N_13048,N_14079);
nor U15115 (N_15115,N_14266,N_13347);
and U15116 (N_15116,N_13966,N_13532);
or U15117 (N_15117,N_12535,N_13109);
xor U15118 (N_15118,N_13970,N_13309);
xor U15119 (N_15119,N_14647,N_14032);
or U15120 (N_15120,N_13316,N_13372);
xor U15121 (N_15121,N_13263,N_12933);
xor U15122 (N_15122,N_14253,N_14922);
nor U15123 (N_15123,N_14892,N_14039);
or U15124 (N_15124,N_12984,N_13856);
nor U15125 (N_15125,N_12980,N_13277);
and U15126 (N_15126,N_12636,N_13008);
nor U15127 (N_15127,N_14828,N_13004);
nor U15128 (N_15128,N_14345,N_14143);
or U15129 (N_15129,N_14193,N_13433);
nor U15130 (N_15130,N_12809,N_14461);
xnor U15131 (N_15131,N_13678,N_14680);
and U15132 (N_15132,N_13564,N_13609);
nor U15133 (N_15133,N_14097,N_13862);
xor U15134 (N_15134,N_13195,N_14271);
or U15135 (N_15135,N_12831,N_14103);
nand U15136 (N_15136,N_14295,N_12508);
and U15137 (N_15137,N_14900,N_14001);
or U15138 (N_15138,N_12672,N_14751);
and U15139 (N_15139,N_13771,N_13952);
xnor U15140 (N_15140,N_12896,N_13453);
nand U15141 (N_15141,N_14500,N_12889);
nor U15142 (N_15142,N_13733,N_13722);
and U15143 (N_15143,N_13776,N_12919);
or U15144 (N_15144,N_13524,N_14018);
nor U15145 (N_15145,N_13180,N_13546);
xor U15146 (N_15146,N_13647,N_14616);
xor U15147 (N_15147,N_14564,N_13328);
nor U15148 (N_15148,N_14252,N_12539);
nor U15149 (N_15149,N_14343,N_13800);
and U15150 (N_15150,N_13307,N_13122);
or U15151 (N_15151,N_14239,N_13495);
nor U15152 (N_15152,N_13114,N_13604);
or U15153 (N_15153,N_14833,N_13521);
xor U15154 (N_15154,N_14960,N_14640);
xor U15155 (N_15155,N_14013,N_13220);
xnor U15156 (N_15156,N_13095,N_14337);
xor U15157 (N_15157,N_14689,N_14943);
and U15158 (N_15158,N_14764,N_14024);
or U15159 (N_15159,N_13852,N_13804);
nor U15160 (N_15160,N_12562,N_13973);
and U15161 (N_15161,N_14612,N_13215);
nand U15162 (N_15162,N_13285,N_13829);
nor U15163 (N_15163,N_13731,N_12774);
and U15164 (N_15164,N_13322,N_13213);
nor U15165 (N_15165,N_13934,N_14965);
nand U15166 (N_15166,N_13989,N_13388);
xor U15167 (N_15167,N_14161,N_14510);
nand U15168 (N_15168,N_13816,N_12976);
nor U15169 (N_15169,N_14507,N_14757);
xor U15170 (N_15170,N_14866,N_13568);
and U15171 (N_15171,N_12982,N_14794);
or U15172 (N_15172,N_14355,N_12738);
nand U15173 (N_15173,N_13504,N_12696);
nor U15174 (N_15174,N_12716,N_14579);
nor U15175 (N_15175,N_14873,N_14423);
and U15176 (N_15176,N_13790,N_13266);
nand U15177 (N_15177,N_12762,N_14332);
or U15178 (N_15178,N_13826,N_14549);
and U15179 (N_15179,N_14466,N_12997);
nor U15180 (N_15180,N_13182,N_14168);
or U15181 (N_15181,N_14971,N_14121);
nor U15182 (N_15182,N_13701,N_14731);
nand U15183 (N_15183,N_14320,N_13956);
or U15184 (N_15184,N_14150,N_13501);
xor U15185 (N_15185,N_13154,N_13936);
nor U15186 (N_15186,N_12907,N_14719);
or U15187 (N_15187,N_13788,N_14635);
xor U15188 (N_15188,N_14407,N_12665);
and U15189 (N_15189,N_13121,N_14497);
and U15190 (N_15190,N_13757,N_13469);
nor U15191 (N_15191,N_13199,N_14827);
xor U15192 (N_15192,N_14668,N_13141);
and U15193 (N_15193,N_14435,N_13378);
nand U15194 (N_15194,N_14352,N_14478);
or U15195 (N_15195,N_14182,N_12519);
xor U15196 (N_15196,N_13377,N_14712);
nand U15197 (N_15197,N_13500,N_14421);
nand U15198 (N_15198,N_14766,N_13555);
xnor U15199 (N_15199,N_13149,N_13014);
nand U15200 (N_15200,N_14063,N_12505);
xnor U15201 (N_15201,N_12647,N_14472);
or U15202 (N_15202,N_14932,N_14464);
and U15203 (N_15203,N_13926,N_14101);
and U15204 (N_15204,N_13750,N_13589);
nor U15205 (N_15205,N_14638,N_14225);
or U15206 (N_15206,N_13584,N_14592);
nor U15207 (N_15207,N_13931,N_14734);
or U15208 (N_15208,N_13093,N_12989);
and U15209 (N_15209,N_14524,N_12839);
nand U15210 (N_15210,N_14584,N_14147);
or U15211 (N_15211,N_13857,N_13713);
xor U15212 (N_15212,N_14037,N_13630);
and U15213 (N_15213,N_13900,N_12836);
nor U15214 (N_15214,N_12776,N_13174);
and U15215 (N_15215,N_13833,N_14587);
nand U15216 (N_15216,N_12953,N_14129);
nor U15217 (N_15217,N_13167,N_14011);
or U15218 (N_15218,N_13284,N_14781);
xor U15219 (N_15219,N_12656,N_14148);
and U15220 (N_15220,N_12916,N_12801);
xnor U15221 (N_15221,N_14308,N_13486);
xor U15222 (N_15222,N_14118,N_14302);
nor U15223 (N_15223,N_12676,N_13084);
and U15224 (N_15224,N_12548,N_13034);
nand U15225 (N_15225,N_13162,N_13484);
xnor U15226 (N_15226,N_12682,N_13695);
nor U15227 (N_15227,N_13030,N_14373);
nand U15228 (N_15228,N_14450,N_13801);
nand U15229 (N_15229,N_12654,N_14970);
or U15230 (N_15230,N_14727,N_12585);
and U15231 (N_15231,N_12791,N_14049);
or U15232 (N_15232,N_13410,N_13542);
or U15233 (N_15233,N_14262,N_13522);
nand U15234 (N_15234,N_13796,N_12937);
nor U15235 (N_15235,N_12579,N_14031);
or U15236 (N_15236,N_14921,N_13529);
nor U15237 (N_15237,N_13230,N_14572);
xnor U15238 (N_15238,N_13752,N_13036);
xnor U15239 (N_15239,N_14889,N_14325);
or U15240 (N_15240,N_13983,N_14931);
and U15241 (N_15241,N_14620,N_14359);
or U15242 (N_15242,N_14220,N_14966);
nor U15243 (N_15243,N_14152,N_12538);
nand U15244 (N_15244,N_13032,N_12534);
nand U15245 (N_15245,N_13155,N_14569);
or U15246 (N_15246,N_14997,N_12787);
and U15247 (N_15247,N_13979,N_14804);
nor U15248 (N_15248,N_13981,N_12759);
xnor U15249 (N_15249,N_14861,N_12955);
xnor U15250 (N_15250,N_12620,N_14980);
xnor U15251 (N_15251,N_14269,N_12901);
nand U15252 (N_15252,N_14184,N_13863);
and U15253 (N_15253,N_14468,N_13773);
nor U15254 (N_15254,N_12602,N_13716);
xnor U15255 (N_15255,N_14846,N_14802);
or U15256 (N_15256,N_13541,N_13961);
nand U15257 (N_15257,N_14930,N_12847);
or U15258 (N_15258,N_13016,N_12796);
and U15259 (N_15259,N_14068,N_13074);
and U15260 (N_15260,N_13982,N_13661);
xnor U15261 (N_15261,N_14436,N_13202);
and U15262 (N_15262,N_13163,N_13885);
xor U15263 (N_15263,N_14318,N_13039);
nand U15264 (N_15264,N_13125,N_13553);
xor U15265 (N_15265,N_13861,N_13444);
or U15266 (N_15266,N_13958,N_14690);
and U15267 (N_15267,N_12527,N_12580);
and U15268 (N_15268,N_13474,N_13634);
nand U15269 (N_15269,N_13502,N_13336);
nor U15270 (N_15270,N_13145,N_14603);
nand U15271 (N_15271,N_13534,N_13427);
or U15272 (N_15272,N_13909,N_12881);
nand U15273 (N_15273,N_14396,N_14397);
nor U15274 (N_15274,N_13459,N_12725);
nand U15275 (N_15275,N_12876,N_14026);
nor U15276 (N_15276,N_13452,N_12873);
nor U15277 (N_15277,N_13997,N_14730);
or U15278 (N_15278,N_14905,N_13419);
or U15279 (N_15279,N_13053,N_14547);
or U15280 (N_15280,N_14626,N_13253);
and U15281 (N_15281,N_13176,N_13324);
or U15282 (N_15282,N_13576,N_13972);
xnor U15283 (N_15283,N_12608,N_13381);
or U15284 (N_15284,N_13482,N_13274);
or U15285 (N_15285,N_14277,N_13256);
and U15286 (N_15286,N_13040,N_13276);
nand U15287 (N_15287,N_14958,N_12560);
or U15288 (N_15288,N_14649,N_13663);
and U15289 (N_15289,N_13005,N_14555);
or U15290 (N_15290,N_12992,N_12972);
xor U15291 (N_15291,N_13676,N_14093);
xor U15292 (N_15292,N_12543,N_14417);
nor U15293 (N_15293,N_12732,N_13779);
nor U15294 (N_15294,N_14055,N_14056);
nand U15295 (N_15295,N_13976,N_14183);
nand U15296 (N_15296,N_12515,N_13571);
and U15297 (N_15297,N_13775,N_13142);
and U15298 (N_15298,N_14177,N_13000);
xor U15299 (N_15299,N_14382,N_13831);
nor U15300 (N_15300,N_14733,N_12987);
and U15301 (N_15301,N_14951,N_14614);
nor U15302 (N_15302,N_12541,N_12913);
nor U15303 (N_15303,N_13919,N_12946);
or U15304 (N_15304,N_13646,N_14329);
nand U15305 (N_15305,N_14185,N_14301);
or U15306 (N_15306,N_13712,N_13238);
or U15307 (N_15307,N_14514,N_14254);
xor U15308 (N_15308,N_14453,N_14178);
nor U15309 (N_15309,N_13888,N_13940);
or U15310 (N_15310,N_14342,N_12596);
xor U15311 (N_15311,N_13843,N_14513);
and U15312 (N_15312,N_13056,N_12915);
or U15313 (N_15313,N_14632,N_14192);
or U15314 (N_15314,N_14140,N_13595);
and U15315 (N_15315,N_12736,N_14655);
xnor U15316 (N_15316,N_14545,N_13415);
nor U15317 (N_15317,N_12693,N_13334);
or U15318 (N_15318,N_13882,N_12808);
nand U15319 (N_15319,N_12536,N_14084);
nor U15320 (N_15320,N_14855,N_13448);
nand U15321 (N_15321,N_13792,N_14222);
or U15322 (N_15322,N_14044,N_14445);
xor U15323 (N_15323,N_12814,N_13283);
nand U15324 (N_15324,N_12530,N_12857);
nand U15325 (N_15325,N_13608,N_14105);
xor U15326 (N_15326,N_13437,N_14947);
xnor U15327 (N_15327,N_12573,N_14153);
and U15328 (N_15328,N_13366,N_13705);
nor U15329 (N_15329,N_14562,N_14999);
nand U15330 (N_15330,N_14282,N_13896);
or U15331 (N_15331,N_13910,N_14718);
and U15332 (N_15332,N_14621,N_14310);
and U15333 (N_15333,N_13839,N_13723);
or U15334 (N_15334,N_12793,N_12604);
xor U15335 (N_15335,N_13755,N_13537);
nand U15336 (N_15336,N_14984,N_14876);
or U15337 (N_15337,N_13246,N_13092);
or U15338 (N_15338,N_13252,N_13015);
or U15339 (N_15339,N_14146,N_14561);
and U15340 (N_15340,N_14328,N_14797);
or U15341 (N_15341,N_12792,N_13268);
nor U15342 (N_15342,N_13756,N_13013);
or U15343 (N_15343,N_13267,N_12581);
and U15344 (N_15344,N_13169,N_13642);
xor U15345 (N_15345,N_13549,N_13018);
nor U15346 (N_15346,N_13047,N_14741);
xnor U15347 (N_15347,N_14717,N_14949);
nand U15348 (N_15348,N_13251,N_13559);
xor U15349 (N_15349,N_12758,N_14772);
nor U15350 (N_15350,N_13239,N_12566);
and U15351 (N_15351,N_14072,N_13075);
nand U15352 (N_15352,N_13985,N_14795);
and U15353 (N_15353,N_14167,N_13416);
nand U15354 (N_15354,N_14636,N_12761);
or U15355 (N_15355,N_14347,N_12940);
nor U15356 (N_15356,N_14858,N_12564);
nand U15357 (N_15357,N_14877,N_14493);
nor U15358 (N_15358,N_13523,N_12936);
nor U15359 (N_15359,N_13999,N_14843);
and U15360 (N_15360,N_13128,N_13819);
nor U15361 (N_15361,N_13889,N_12746);
nor U15362 (N_15362,N_14618,N_12966);
xor U15363 (N_15363,N_13590,N_12698);
xor U15364 (N_15364,N_12576,N_13869);
nand U15365 (N_15365,N_14165,N_14145);
nand U15366 (N_15366,N_14685,N_12902);
nand U15367 (N_15367,N_12773,N_13746);
or U15368 (N_15368,N_13922,N_13944);
nor U15369 (N_15369,N_13629,N_14366);
and U15370 (N_15370,N_13480,N_13743);
nor U15371 (N_15371,N_13379,N_13622);
nor U15372 (N_15372,N_13411,N_14214);
nand U15373 (N_15373,N_12529,N_12798);
or U15374 (N_15374,N_14459,N_14314);
xor U15375 (N_15375,N_12775,N_14819);
and U15376 (N_15376,N_14869,N_14938);
nor U15377 (N_15377,N_14083,N_14371);
nor U15378 (N_15378,N_13157,N_12872);
nor U15379 (N_15379,N_14765,N_13744);
or U15380 (N_15380,N_13160,N_13515);
xor U15381 (N_15381,N_13812,N_13967);
and U15382 (N_15382,N_14599,N_14929);
nand U15383 (N_15383,N_12931,N_13305);
or U15384 (N_15384,N_14157,N_14291);
and U15385 (N_15385,N_14515,N_14172);
nand U15386 (N_15386,N_14059,N_12540);
xor U15387 (N_15387,N_13656,N_13353);
nor U15388 (N_15388,N_14280,N_12748);
xor U15389 (N_15389,N_12849,N_13467);
or U15390 (N_15390,N_14750,N_13209);
xnor U15391 (N_15391,N_13735,N_13129);
or U15392 (N_15392,N_12565,N_14512);
nor U15393 (N_15393,N_12545,N_12990);
nand U15394 (N_15394,N_13468,N_13886);
or U15395 (N_15395,N_14986,N_12544);
or U15396 (N_15396,N_12658,N_13478);
xnor U15397 (N_15397,N_12895,N_12552);
nand U15398 (N_15398,N_12615,N_12528);
nand U15399 (N_15399,N_12743,N_14309);
xnor U15400 (N_15400,N_13702,N_12879);
and U15401 (N_15401,N_14556,N_12810);
nand U15402 (N_15402,N_13099,N_14414);
nand U15403 (N_15403,N_13901,N_14927);
xnor U15404 (N_15404,N_14693,N_13064);
or U15405 (N_15405,N_13310,N_12719);
xnor U15406 (N_15406,N_13458,N_12670);
xor U15407 (N_15407,N_13741,N_14284);
nor U15408 (N_15408,N_14527,N_14054);
nor U15409 (N_15409,N_14380,N_13658);
xnor U15410 (N_15410,N_14810,N_14057);
or U15411 (N_15411,N_14304,N_12633);
or U15412 (N_15412,N_13420,N_13383);
or U15413 (N_15413,N_13631,N_13455);
nand U15414 (N_15414,N_14823,N_12906);
nor U15415 (N_15415,N_13300,N_13146);
nand U15416 (N_15416,N_13451,N_13949);
or U15417 (N_15417,N_14449,N_13082);
or U15418 (N_15418,N_14776,N_14189);
or U15419 (N_15419,N_13783,N_13980);
or U15420 (N_15420,N_13200,N_14033);
nand U15421 (N_15421,N_13893,N_12631);
nand U15422 (N_15422,N_14698,N_14822);
xor U15423 (N_15423,N_13548,N_13192);
or U15424 (N_15424,N_13587,N_14639);
xor U15425 (N_15425,N_13165,N_14541);
xor U15426 (N_15426,N_13248,N_14737);
nor U15427 (N_15427,N_14442,N_12991);
nor U15428 (N_15428,N_14073,N_13510);
or U15429 (N_15429,N_13850,N_14361);
or U15430 (N_15430,N_12888,N_12659);
or U15431 (N_15431,N_13598,N_14977);
nand U15432 (N_15432,N_13401,N_13052);
xnor U15433 (N_15433,N_13729,N_14455);
or U15434 (N_15434,N_13506,N_12828);
nor U15435 (N_15435,N_14230,N_13219);
nor U15436 (N_15436,N_12804,N_12753);
xnor U15437 (N_15437,N_14887,N_12840);
nand U15438 (N_15438,N_14009,N_13760);
or U15439 (N_15439,N_13593,N_13512);
or U15440 (N_15440,N_14306,N_14498);
xor U15441 (N_15441,N_13641,N_14155);
xnor U15442 (N_15442,N_14811,N_13083);
xnor U15443 (N_15443,N_13335,N_13096);
or U15444 (N_15444,N_14069,N_13139);
and U15445 (N_15445,N_13077,N_13186);
and U15446 (N_15446,N_14201,N_13320);
xnor U15447 (N_15447,N_13834,N_12819);
nand U15448 (N_15448,N_12996,N_13573);
or U15449 (N_15449,N_12533,N_14535);
nor U15450 (N_15450,N_13244,N_12558);
and U15451 (N_15451,N_13845,N_14944);
or U15452 (N_15452,N_13654,N_14882);
and U15453 (N_15453,N_14580,N_14135);
nand U15454 (N_15454,N_14563,N_14856);
or U15455 (N_15455,N_13577,N_13321);
nand U15456 (N_15456,N_14682,N_14215);
and U15457 (N_15457,N_13137,N_14785);
xnor U15458 (N_15458,N_13126,N_14326);
nor U15459 (N_15459,N_14962,N_13302);
nor U15460 (N_15460,N_13786,N_13187);
and U15461 (N_15461,N_12777,N_13751);
or U15462 (N_15462,N_13234,N_14906);
nor U15463 (N_15463,N_14094,N_14367);
nor U15464 (N_15464,N_14491,N_14433);
nand U15465 (N_15465,N_13435,N_13078);
nand U15466 (N_15466,N_13742,N_14862);
xor U15467 (N_15467,N_13643,N_13894);
or U15468 (N_15468,N_14067,N_12506);
and U15469 (N_15469,N_13876,N_14346);
nand U15470 (N_15470,N_14501,N_14275);
and U15471 (N_15471,N_12503,N_13503);
nor U15472 (N_15472,N_13289,N_14875);
nand U15473 (N_15473,N_14125,N_13517);
and U15474 (N_15474,N_14898,N_13009);
nand U15475 (N_15475,N_13208,N_12655);
nand U15476 (N_15476,N_14290,N_13575);
and U15477 (N_15477,N_14274,N_13446);
nand U15478 (N_15478,N_13023,N_14703);
and U15479 (N_15479,N_13373,N_12833);
xor U15480 (N_15480,N_14897,N_12878);
xor U15481 (N_15481,N_14369,N_14070);
or U15482 (N_15482,N_12877,N_14913);
and U15483 (N_15483,N_12695,N_12795);
and U15484 (N_15484,N_12854,N_14392);
nand U15485 (N_15485,N_12782,N_12747);
nor U15486 (N_15486,N_14176,N_14972);
nand U15487 (N_15487,N_13853,N_14247);
and U15488 (N_15488,N_12979,N_13405);
or U15489 (N_15489,N_13260,N_12897);
nand U15490 (N_15490,N_13607,N_13955);
and U15491 (N_15491,N_13665,N_14285);
xnor U15492 (N_15492,N_12850,N_13229);
and U15493 (N_15493,N_14348,N_12605);
xnor U15494 (N_15494,N_14470,N_12690);
nand U15495 (N_15495,N_14341,N_14821);
nand U15496 (N_15496,N_12772,N_13873);
nand U15497 (N_15497,N_12947,N_13397);
or U15498 (N_15498,N_12691,N_13060);
and U15499 (N_15499,N_14040,N_14761);
xor U15500 (N_15500,N_13904,N_13747);
nor U15501 (N_15501,N_13520,N_14803);
or U15502 (N_15502,N_12932,N_14231);
xor U15503 (N_15503,N_14204,N_13891);
or U15504 (N_15504,N_13103,N_13376);
xnor U15505 (N_15505,N_13807,N_14691);
or U15506 (N_15506,N_14360,N_13895);
nor U15507 (N_15507,N_14738,N_13963);
nor U15508 (N_15508,N_14319,N_12780);
nand U15509 (N_15509,N_14820,N_14186);
xor U15510 (N_15510,N_14678,N_13194);
xnor U15511 (N_15511,N_13235,N_14412);
and U15512 (N_15512,N_13518,N_13509);
nor U15513 (N_15513,N_14122,N_13986);
nand U15514 (N_15514,N_12806,N_13025);
nand U15515 (N_15515,N_12706,N_14065);
or U15516 (N_15516,N_14224,N_13536);
nand U15517 (N_15517,N_14142,N_14250);
or U15518 (N_15518,N_14611,N_12627);
or U15519 (N_15519,N_13650,N_13525);
and U15520 (N_15520,N_13068,N_14313);
nor U15521 (N_15521,N_13942,N_14430);
and U15522 (N_15522,N_13905,N_14173);
and U15523 (N_15523,N_13105,N_14763);
nor U15524 (N_15524,N_13423,N_13715);
nand U15525 (N_15525,N_13403,N_14210);
and U15526 (N_15526,N_12524,N_13667);
or U15527 (N_15527,N_13315,N_14842);
and U15528 (N_15528,N_13293,N_12869);
xnor U15529 (N_15529,N_13191,N_14060);
nor U15530 (N_15530,N_12511,N_13581);
or U15531 (N_15531,N_14663,N_14233);
or U15532 (N_15532,N_12884,N_13233);
xor U15533 (N_15533,N_14279,N_12848);
nor U15534 (N_15534,N_13421,N_13583);
or U15535 (N_15535,N_14700,N_14022);
nand U15536 (N_15536,N_13717,N_13456);
xnor U15537 (N_15537,N_13817,N_13319);
xnor U15538 (N_15538,N_13754,N_13090);
and U15539 (N_15539,N_14989,N_12813);
or U15540 (N_15540,N_14624,N_14081);
or U15541 (N_15541,N_12927,N_13070);
nand U15542 (N_15542,N_13247,N_13497);
nand U15543 (N_15543,N_13683,N_12705);
xnor U15544 (N_15544,N_14133,N_13171);
or U15545 (N_15545,N_14012,N_12500);
nand U15546 (N_15546,N_14518,N_12858);
or U15547 (N_15547,N_14749,N_13488);
xnor U15548 (N_15548,N_12790,N_12767);
xor U15549 (N_15549,N_13454,N_12752);
or U15550 (N_15550,N_13136,N_12960);
nand U15551 (N_15551,N_12588,N_14520);
and U15552 (N_15552,N_14851,N_14752);
nor U15553 (N_15553,N_14321,N_13306);
nand U15554 (N_15554,N_13431,N_14211);
nand U15555 (N_15555,N_14091,N_14881);
or U15556 (N_15556,N_14835,N_14714);
xnor U15557 (N_15557,N_13513,N_12568);
nor U15558 (N_15558,N_14798,N_14344);
and U15559 (N_15559,N_14092,N_14585);
nor U15560 (N_15560,N_14404,N_14601);
and U15561 (N_15561,N_14955,N_13507);
and U15562 (N_15562,N_13365,N_13880);
xnor U15563 (N_15563,N_14503,N_14760);
nor U15564 (N_15564,N_13814,N_14818);
nand U15565 (N_15565,N_13203,N_12771);
or U15566 (N_15566,N_12704,N_13838);
nand U15567 (N_15567,N_13279,N_12769);
or U15568 (N_15568,N_14939,N_14114);
and U15569 (N_15569,N_14149,N_14003);
nor U15570 (N_15570,N_14474,N_13612);
and U15571 (N_15571,N_14759,N_14870);
or U15572 (N_15572,N_14790,N_13912);
or U15573 (N_15573,N_13925,N_14123);
xor U15574 (N_15574,N_13721,N_13232);
nor U15575 (N_15575,N_13599,N_14036);
or U15576 (N_15576,N_14953,N_12822);
or U15577 (N_15577,N_13257,N_12794);
xnor U15578 (N_15578,N_14050,N_13362);
and U15579 (N_15579,N_14656,N_13566);
xor U15580 (N_15580,N_14653,N_14716);
or U15581 (N_15581,N_12920,N_14006);
nand U15582 (N_15582,N_12592,N_14586);
nand U15583 (N_15583,N_14721,N_13120);
or U15584 (N_15584,N_14998,N_13606);
or U15585 (N_15585,N_14273,N_13156);
nand U15586 (N_15586,N_14565,N_12619);
nor U15587 (N_15587,N_13425,N_13491);
and U15588 (N_15588,N_13923,N_14753);
nor U15589 (N_15589,N_13355,N_12890);
xor U15590 (N_15590,N_13291,N_13261);
nor U15591 (N_15591,N_12886,N_14747);
nand U15592 (N_15592,N_14800,N_13585);
xor U15593 (N_15593,N_13402,N_12859);
or U15594 (N_15594,N_13342,N_14043);
nor U15595 (N_15595,N_14241,N_14194);
or U15596 (N_15596,N_14625,N_13791);
nand U15597 (N_15597,N_14078,N_13363);
or U15598 (N_15598,N_13487,N_14768);
and U15599 (N_15599,N_13533,N_14130);
xnor U15600 (N_15600,N_12924,N_13361);
nor U15601 (N_15601,N_14029,N_13368);
or U15602 (N_15602,N_13657,N_12863);
or U15603 (N_15603,N_13704,N_13539);
or U15604 (N_15604,N_13978,N_13351);
and U15605 (N_15605,N_12550,N_13866);
and U15606 (N_15606,N_14251,N_14144);
nor U15607 (N_15607,N_14467,N_14451);
and U15608 (N_15608,N_13653,N_14560);
or U15609 (N_15609,N_14317,N_14316);
and U15610 (N_15610,N_14886,N_14940);
xnor U15611 (N_15611,N_12577,N_13153);
nand U15612 (N_15612,N_14868,N_14315);
nor U15613 (N_15613,N_14180,N_13728);
or U15614 (N_15614,N_13724,N_14568);
or U15615 (N_15615,N_13471,N_14664);
nor U15616 (N_15616,N_14744,N_14334);
xnor U15617 (N_15617,N_12635,N_13748);
xor U15618 (N_15618,N_12783,N_12521);
nor U15619 (N_15619,N_13175,N_13327);
nand U15620 (N_15620,N_12838,N_13911);
nand U15621 (N_15621,N_13820,N_13184);
xnor U15622 (N_15622,N_12846,N_14196);
or U15623 (N_15623,N_14265,N_14223);
nand U15624 (N_15624,N_13582,N_13929);
nand U15625 (N_15625,N_13144,N_12708);
and U15626 (N_15626,N_12871,N_12666);
xnor U15627 (N_15627,N_14099,N_14992);
nand U15628 (N_15628,N_12975,N_14901);
or U15629 (N_15629,N_13380,N_14762);
and U15630 (N_15630,N_14190,N_12523);
xnor U15631 (N_15631,N_12741,N_13394);
xnor U15632 (N_15632,N_13088,N_14061);
or U15633 (N_15633,N_13150,N_14826);
or U15634 (N_15634,N_14336,N_13494);
nand U15635 (N_15635,N_14390,N_12639);
and U15636 (N_15636,N_14857,N_14609);
xor U15637 (N_15637,N_14350,N_12880);
and U15638 (N_15638,N_14480,N_13811);
nand U15639 (N_15639,N_14619,N_13782);
xnor U15640 (N_15640,N_13172,N_12621);
xnor U15641 (N_15641,N_13107,N_12825);
nor U15642 (N_15642,N_14604,N_13700);
nor U15643 (N_15643,N_14377,N_14907);
nor U15644 (N_15644,N_12599,N_13442);
or U15645 (N_15645,N_12642,N_13189);
or U15646 (N_15646,N_14489,N_13406);
or U15647 (N_15647,N_13627,N_12513);
nor U15648 (N_15648,N_14354,N_14686);
and U15649 (N_15649,N_14854,N_12952);
nand U15650 (N_15650,N_13231,N_14375);
or U15651 (N_15651,N_12587,N_13868);
nor U15652 (N_15652,N_12618,N_14402);
nand U15653 (N_15653,N_13483,N_12663);
or U15654 (N_15654,N_14643,N_14025);
and U15655 (N_15655,N_13330,N_12755);
nor U15656 (N_15656,N_13830,N_13177);
and U15657 (N_15657,N_14669,N_13080);
or U15658 (N_15658,N_13516,N_13436);
nor U15659 (N_15659,N_12922,N_13921);
nand U15660 (N_15660,N_13567,N_12757);
and U15661 (N_15661,N_14742,N_14425);
xnor U15662 (N_15662,N_13398,N_12789);
nor U15663 (N_15663,N_14476,N_14107);
and U15664 (N_15664,N_14885,N_14226);
or U15665 (N_15665,N_14865,N_14871);
or U15666 (N_15666,N_14837,N_13221);
and U15667 (N_15667,N_12611,N_14387);
nand U15668 (N_15668,N_14198,N_13466);
xor U15669 (N_15669,N_14292,N_13389);
nand U15670 (N_15670,N_12827,N_12607);
and U15671 (N_15671,N_14975,N_13907);
or U15672 (N_15672,N_13135,N_13100);
xor U15673 (N_15673,N_13043,N_13051);
nor U15674 (N_15674,N_12797,N_13031);
nor U15675 (N_15675,N_14736,N_14902);
and U15676 (N_15676,N_12711,N_13489);
and U15677 (N_15677,N_14492,N_14728);
and U15678 (N_15678,N_13648,N_13588);
xor U15679 (N_15679,N_13367,N_14539);
or U15680 (N_15680,N_13111,N_13226);
nor U15681 (N_15681,N_13938,N_14353);
xnor U15682 (N_15682,N_13709,N_14769);
nand U15683 (N_15683,N_14447,N_14156);
and U15684 (N_15684,N_13439,N_14126);
nand U15685 (N_15685,N_14508,N_13346);
or U15686 (N_15686,N_13699,N_14945);
and U15687 (N_15687,N_14658,N_14509);
or U15688 (N_15688,N_12669,N_14634);
or U15689 (N_15689,N_14942,N_14335);
nor U15690 (N_15690,N_14771,N_14688);
and U15691 (N_15691,N_13770,N_14116);
xnor U15692 (N_15692,N_14959,N_13987);
xor U15693 (N_15693,N_14418,N_14950);
nor U15694 (N_15694,N_12553,N_12844);
or U15695 (N_15695,N_14683,N_13460);
or U15696 (N_15696,N_13119,N_14401);
xor U15697 (N_15697,N_13964,N_12561);
and U15698 (N_15698,N_14349,N_13364);
nand U15699 (N_15699,N_13951,N_13001);
and U15700 (N_15700,N_13210,N_13793);
xnor U15701 (N_15701,N_14729,N_12928);
nand U15702 (N_15702,N_13358,N_14884);
nand U15703 (N_15703,N_12834,N_12914);
nand U15704 (N_15704,N_13337,N_13562);
nand U15705 (N_15705,N_13594,N_12970);
and U15706 (N_15706,N_14517,N_12898);
nand U15707 (N_15707,N_14278,N_13848);
xnor U15708 (N_15708,N_12841,N_14365);
nand U15709 (N_15709,N_13044,N_12807);
and U15710 (N_15710,N_12909,N_12641);
nand U15711 (N_15711,N_14813,N_13438);
or U15712 (N_15712,N_12510,N_13835);
nand U15713 (N_15713,N_12981,N_14115);
nand U15714 (N_15714,N_12837,N_12572);
and U15715 (N_15715,N_14628,N_13029);
nand U15716 (N_15716,N_13827,N_12653);
xor U15717 (N_15717,N_14710,N_12677);
xnor U15718 (N_15718,N_14496,N_13759);
xnor U15719 (N_15719,N_14495,N_13148);
xor U15720 (N_15720,N_14504,N_14408);
or U15721 (N_15721,N_12595,N_12703);
xnor U15722 (N_15722,N_13994,N_12700);
or U15723 (N_15723,N_13295,N_12910);
nor U15724 (N_15724,N_12603,N_13939);
nand U15725 (N_15725,N_14591,N_14411);
and U15726 (N_15726,N_13159,N_14571);
or U15727 (N_15727,N_14651,N_13087);
or U15728 (N_15728,N_12930,N_13188);
and U15729 (N_15729,N_13479,N_14831);
xnor U15730 (N_15730,N_13613,N_12699);
xor U15731 (N_15731,N_12742,N_14602);
or U15732 (N_15732,N_12892,N_13275);
or U15733 (N_15733,N_13825,N_14429);
or U15734 (N_15734,N_13913,N_14824);
xor U15735 (N_15735,N_14711,N_13652);
xnor U15736 (N_15736,N_13890,N_14199);
and U15737 (N_15737,N_12870,N_13651);
and U15738 (N_15738,N_14454,N_13271);
or U15739 (N_15739,N_14217,N_14134);
and U15740 (N_15740,N_12686,N_12502);
xnor U15741 (N_15741,N_14327,N_14398);
and U15742 (N_15742,N_13340,N_14705);
nand U15743 (N_15743,N_13259,N_13124);
nand U15744 (N_15744,N_13946,N_14437);
xor U15745 (N_15745,N_13329,N_13860);
and U15746 (N_15746,N_14471,N_14007);
nand U15747 (N_15747,N_14276,N_13688);
nand U15748 (N_15748,N_14812,N_13112);
and U15749 (N_15749,N_12853,N_12594);
nor U15750 (N_15750,N_14829,N_12731);
nand U15751 (N_15751,N_14667,N_13745);
nor U15752 (N_15752,N_13726,N_14399);
or U15753 (N_15753,N_13430,N_13033);
nand U15754 (N_15754,N_13669,N_14158);
or U15755 (N_15755,N_14937,N_13694);
nor U15756 (N_15756,N_12965,N_13828);
xor U15757 (N_15757,N_14299,N_14058);
nand U15758 (N_15758,N_14912,N_13881);
nor U15759 (N_15759,N_13691,N_14860);
or U15760 (N_15760,N_13131,N_14212);
nand U15761 (N_15761,N_13734,N_14720);
and U15762 (N_15762,N_13635,N_13738);
nor U15763 (N_15763,N_12779,N_14351);
or U15764 (N_15764,N_14322,N_14166);
nand U15765 (N_15765,N_13059,N_13626);
nand U15766 (N_15766,N_13639,N_14888);
nand U15767 (N_15767,N_14370,N_14077);
nor U15768 (N_15768,N_14245,N_14709);
nand U15769 (N_15769,N_14573,N_14740);
nor U15770 (N_15770,N_14238,N_14203);
nor U15771 (N_15771,N_13574,N_14028);
xor U15772 (N_15772,N_12964,N_13655);
and U15773 (N_15773,N_14465,N_12584);
and U15774 (N_15774,N_13736,N_13969);
or U15775 (N_15775,N_13020,N_14627);
and U15776 (N_15776,N_14696,N_14008);
nand U15777 (N_15777,N_12662,N_14424);
and U15778 (N_15778,N_13408,N_13684);
nand U15779 (N_15779,N_13254,N_14623);
xnor U15780 (N_15780,N_14976,N_13102);
nand U15781 (N_15781,N_13498,N_14088);
nor U15782 (N_15782,N_14637,N_14494);
and U15783 (N_15783,N_14676,N_13384);
or U15784 (N_15784,N_14260,N_14041);
nor U15785 (N_15785,N_13356,N_13073);
nand U15786 (N_15786,N_13769,N_13344);
nand U15787 (N_15787,N_14806,N_14671);
nand U15788 (N_15788,N_13003,N_13535);
nand U15789 (N_15789,N_14724,N_13644);
and U15790 (N_15790,N_12832,N_14038);
and U15791 (N_15791,N_13780,N_14181);
and U15792 (N_15792,N_13865,N_14849);
xnor U15793 (N_15793,N_13265,N_13847);
and U15794 (N_15794,N_14543,N_13212);
and U15795 (N_15795,N_14413,N_12824);
xnor U15796 (N_15796,N_12582,N_13076);
nand U15797 (N_15797,N_14416,N_13370);
nor U15798 (N_15798,N_13556,N_14559);
xnor U15799 (N_15799,N_12707,N_14506);
or U15800 (N_15800,N_14695,N_14287);
xor U15801 (N_15801,N_14339,N_14074);
and U15802 (N_15802,N_13465,N_12803);
xnor U15803 (N_15803,N_14582,N_14780);
nor U15804 (N_15804,N_14532,N_14872);
and U15805 (N_15805,N_12935,N_13463);
or U15806 (N_15806,N_14452,N_13971);
xor U15807 (N_15807,N_12830,N_13006);
or U15808 (N_15808,N_12709,N_14814);
nand U15809 (N_15809,N_14848,N_12557);
and U15810 (N_15810,N_12590,N_13243);
nand U15811 (N_15811,N_14236,N_14540);
nor U15812 (N_15812,N_14064,N_13390);
nor U15813 (N_15813,N_14933,N_14394);
xor U15814 (N_15814,N_13341,N_12826);
nand U15815 (N_15815,N_14895,N_13708);
nor U15816 (N_15816,N_13620,N_13619);
nand U15817 (N_15817,N_13932,N_12985);
nor U15818 (N_15818,N_14926,N_12733);
or U15819 (N_15819,N_14880,N_14200);
nor U15820 (N_15820,N_12941,N_12986);
or U15821 (N_15821,N_13679,N_14288);
and U15822 (N_15822,N_13069,N_14847);
and U15823 (N_15823,N_14815,N_13193);
nand U15824 (N_15824,N_13998,N_12957);
nor U15825 (N_15825,N_14606,N_13822);
nand U15826 (N_15826,N_14641,N_14791);
nor U15827 (N_15827,N_14419,N_14529);
nor U15828 (N_15828,N_13965,N_14670);
or U15829 (N_15829,N_13789,N_13287);
nor U15830 (N_15830,N_12555,N_13026);
xnor U15831 (N_15831,N_13849,N_13764);
nor U15832 (N_15832,N_14486,N_13443);
and U15833 (N_15833,N_14324,N_14694);
or U15834 (N_15834,N_14405,N_14566);
and U15835 (N_15835,N_13130,N_13519);
nand U15836 (N_15836,N_13732,N_14257);
xnor U15837 (N_15837,N_13638,N_13270);
or U15838 (N_15838,N_14191,N_12763);
and U15839 (N_15839,N_14087,N_14374);
xnor U15840 (N_15840,N_13242,N_14596);
xor U15841 (N_15841,N_13086,N_14410);
xor U15842 (N_15842,N_13995,N_14595);
nor U15843 (N_15843,N_14948,N_13017);
nor U15844 (N_15844,N_13993,N_14598);
and U15845 (N_15845,N_14923,N_14234);
or U15846 (N_15846,N_13101,N_13579);
xnor U15847 (N_15847,N_14393,N_14935);
nor U15848 (N_15848,N_13924,N_14839);
nand U15849 (N_15849,N_12958,N_14659);
xnor U15850 (N_15850,N_13603,N_12556);
xnor U15851 (N_15851,N_14294,N_12739);
or U15852 (N_15852,N_13098,N_13531);
nor U15853 (N_15853,N_12887,N_12622);
nand U15854 (N_15854,N_13505,N_14896);
nor U15855 (N_15855,N_13286,N_13470);
or U15856 (N_15856,N_13935,N_14874);
nor U15857 (N_15857,N_14131,N_14502);
or U15858 (N_15858,N_12600,N_14076);
or U15859 (N_15859,N_14779,N_14098);
or U15860 (N_15860,N_13392,N_14622);
or U15861 (N_15861,N_14805,N_14745);
or U15862 (N_15862,N_14558,N_12865);
or U15863 (N_15863,N_12944,N_14446);
xnor U15864 (N_15864,N_14179,N_13313);
xnor U15865 (N_15865,N_14187,N_13737);
xnor U15866 (N_15866,N_12681,N_13081);
or U15867 (N_15867,N_14665,N_13803);
nor U15868 (N_15868,N_14832,N_13249);
nor U15869 (N_15869,N_13872,N_13718);
xor U15870 (N_15870,N_14605,N_12517);
and U15871 (N_15871,N_13241,N_13706);
nand U15872 (N_15872,N_13975,N_13434);
xnor U15873 (N_15873,N_12768,N_12570);
or U15874 (N_15874,N_14739,N_13903);
nor U15875 (N_15875,N_13508,N_14389);
nor U15876 (N_15876,N_13841,N_13216);
and U15877 (N_15877,N_14296,N_14551);
or U15878 (N_15878,N_13152,N_14538);
nand U15879 (N_15879,N_14021,N_14754);
nor U15880 (N_15880,N_14809,N_13424);
xnor U15881 (N_15881,N_12943,N_13908);
nor U15882 (N_15882,N_13920,N_14546);
nor U15883 (N_15883,N_14748,N_14830);
xor U15884 (N_15884,N_14867,N_13526);
or U15885 (N_15885,N_13391,N_12614);
and U15886 (N_15886,N_12509,N_12978);
nor U15887 (N_15887,N_14307,N_13892);
xnor U15888 (N_15888,N_14590,N_14046);
nand U15889 (N_15889,N_14715,N_14263);
nor U15890 (N_15890,N_13601,N_14778);
and U15891 (N_15891,N_13115,N_12805);
xor U15892 (N_15892,N_12766,N_13947);
nor U15893 (N_15893,N_13628,N_14679);
nand U15894 (N_15894,N_13514,N_12692);
and U15895 (N_15895,N_14681,N_12730);
and U15896 (N_15896,N_14090,N_12925);
nor U15897 (N_15897,N_14272,N_13447);
nand U15898 (N_15898,N_14963,N_13806);
nand U15899 (N_15899,N_14777,N_13762);
nand U15900 (N_15900,N_13079,N_14109);
nand U15901 (N_15901,N_12929,N_12860);
or U15902 (N_15902,N_12951,N_13846);
and U15903 (N_15903,N_13113,N_12899);
and U15904 (N_15904,N_14915,N_13462);
and U15905 (N_15905,N_13711,N_13185);
nand U15906 (N_15906,N_13787,N_14916);
and U15907 (N_15907,N_14525,N_12820);
and U15908 (N_15908,N_12974,N_13884);
and U15909 (N_15909,N_14607,N_14581);
and U15910 (N_15910,N_14075,N_12862);
and U15911 (N_15911,N_14575,N_13945);
or U15912 (N_15912,N_14583,N_13550);
xor U15913 (N_15913,N_13002,N_12675);
xnor U15914 (N_15914,N_13481,N_12900);
nand U15915 (N_15915,N_12722,N_13440);
xnor U15916 (N_15916,N_12770,N_14859);
xnor U15917 (N_15917,N_14675,N_12578);
and U15918 (N_15918,N_13569,N_14890);
xnor U15919 (N_15919,N_14973,N_14481);
and U15920 (N_15920,N_12983,N_14428);
or U15921 (N_15921,N_14505,N_12934);
and U15922 (N_15922,N_12678,N_12816);
nand U15923 (N_15923,N_13333,N_12650);
nand U15924 (N_15924,N_13797,N_13844);
or U15925 (N_15925,N_13343,N_12549);
nand U15926 (N_15926,N_13707,N_13858);
nor U15927 (N_15927,N_12551,N_13049);
xnor U15928 (N_15928,N_12684,N_13272);
xor U15929 (N_15929,N_13697,N_13211);
nand U15930 (N_15930,N_14364,N_14706);
nand U15931 (N_15931,N_12598,N_12751);
or U15932 (N_15932,N_13097,N_14248);
nand U15933 (N_15933,N_14286,N_14713);
or U15934 (N_15934,N_14311,N_13916);
xnor U15935 (N_15935,N_13918,N_13855);
and U15936 (N_15936,N_12683,N_12998);
or U15937 (N_15937,N_14386,N_14283);
nor U15938 (N_15938,N_13580,N_14677);
xor U15939 (N_15939,N_14894,N_12532);
xnor U15940 (N_15940,N_13851,N_14746);
or U15941 (N_15941,N_13761,N_12547);
nand U15942 (N_15942,N_13065,N_14015);
xnor U15943 (N_15943,N_13022,N_14594);
and U15944 (N_15944,N_13354,N_14666);
and U15945 (N_15945,N_12563,N_14521);
xor U15946 (N_15946,N_13666,N_14817);
nor U15947 (N_15947,N_14438,N_13071);
nand U15948 (N_15948,N_14941,N_12885);
nand U15949 (N_15949,N_13696,N_13941);
nor U15950 (N_15950,N_14458,N_14996);
xnor U15951 (N_15951,N_13887,N_13600);
nor U15952 (N_15952,N_13325,N_13294);
xnor U15953 (N_15953,N_13382,N_14792);
nor U15954 (N_15954,N_13511,N_13066);
xor U15955 (N_15955,N_14983,N_13134);
and U15956 (N_15956,N_13496,N_12856);
or U15957 (N_15957,N_13255,N_13689);
nor U15958 (N_15958,N_13314,N_13572);
nor U15959 (N_15959,N_12649,N_13281);
or U15960 (N_15960,N_12949,N_14246);
xnor U15961 (N_15961,N_13917,N_14169);
or U15962 (N_15962,N_12994,N_14552);
or U15963 (N_15963,N_14207,N_12893);
and U15964 (N_15964,N_14807,N_13170);
nor U15965 (N_15965,N_13874,N_12734);
and U15966 (N_15966,N_14082,N_13207);
or U15967 (N_15967,N_14633,N_12842);
or U15968 (N_15968,N_12737,N_13357);
and U15969 (N_15969,N_14104,N_14281);
nor U15970 (N_15970,N_13611,N_13714);
nor U15971 (N_15971,N_12977,N_13551);
or U15972 (N_15972,N_13927,N_14985);
and U15973 (N_15973,N_14171,N_13123);
nand U15974 (N_15974,N_14434,N_13610);
nor U15975 (N_15975,N_13058,N_13557);
nand U15976 (N_15976,N_13703,N_13450);
or U15977 (N_15977,N_13472,N_13490);
or U15978 (N_15978,N_14381,N_13067);
and U15979 (N_15979,N_12875,N_14139);
nor U15980 (N_15980,N_14047,N_13774);
xnor U15981 (N_15981,N_13326,N_14704);
nand U15982 (N_15982,N_14422,N_13824);
nor U15983 (N_15983,N_13565,N_12921);
nand U15984 (N_15984,N_14773,N_14376);
and U15985 (N_15985,N_12868,N_13426);
xnor U15986 (N_15986,N_13021,N_14732);
nor U15987 (N_15987,N_14100,N_13473);
nor U15988 (N_15988,N_12720,N_14229);
nor U15989 (N_15989,N_12601,N_14834);
nand U15990 (N_15990,N_14002,N_12939);
nor U15991 (N_15991,N_14333,N_13954);
and U15992 (N_15992,N_13223,N_14523);
nor U15993 (N_15993,N_14483,N_14650);
and U15994 (N_15994,N_13301,N_13236);
xnor U15995 (N_15995,N_13974,N_14816);
and U15996 (N_15996,N_13290,N_14356);
nor U15997 (N_15997,N_14170,N_13859);
or U15998 (N_15998,N_14312,N_12778);
or U15999 (N_15999,N_13794,N_13360);
and U16000 (N_16000,N_14237,N_13690);
nor U16001 (N_16001,N_12729,N_13968);
or U16002 (N_16002,N_14838,N_13960);
nand U16003 (N_16003,N_13879,N_13660);
nand U16004 (N_16004,N_14300,N_14775);
nor U16005 (N_16005,N_12554,N_14954);
or U16006 (N_16006,N_12754,N_12995);
and U16007 (N_16007,N_14255,N_14597);
nand U16008 (N_16008,N_12959,N_14052);
nand U16009 (N_16009,N_12971,N_14630);
and U16010 (N_16010,N_14864,N_13883);
xor U16011 (N_16011,N_12963,N_14615);
or U16012 (N_16012,N_12652,N_13686);
xor U16013 (N_16013,N_14610,N_13615);
and U16014 (N_16014,N_12648,N_14305);
or U16015 (N_16015,N_13089,N_12687);
nor U16016 (N_16016,N_14578,N_13959);
or U16017 (N_16017,N_13164,N_13659);
and U16018 (N_16018,N_14112,N_14110);
and U16019 (N_16019,N_13204,N_14608);
nor U16020 (N_16020,N_13877,N_14197);
xor U16021 (N_16021,N_13687,N_14799);
xnor U16022 (N_16022,N_13928,N_14672);
nand U16023 (N_16023,N_14485,N_14988);
or U16024 (N_16024,N_13399,N_12522);
nand U16025 (N_16025,N_13323,N_12617);
nand U16026 (N_16026,N_14743,N_12861);
nor U16027 (N_16027,N_12891,N_13637);
nand U16028 (N_16028,N_14415,N_14662);
nand U16029 (N_16029,N_13836,N_12882);
xor U16030 (N_16030,N_13906,N_14982);
or U16031 (N_16031,N_13875,N_13766);
nor U16032 (N_16032,N_14879,N_13592);
nand U16033 (N_16033,N_13984,N_12644);
nand U16034 (N_16034,N_14570,N_13664);
or U16035 (N_16035,N_12800,N_13823);
nor U16036 (N_16036,N_14403,N_13228);
nor U16037 (N_16037,N_12574,N_13375);
and U16038 (N_16038,N_12950,N_12542);
or U16039 (N_16039,N_13218,N_14440);
nand U16040 (N_16040,N_12715,N_14786);
nor U16041 (N_16041,N_12812,N_12894);
xnor U16042 (N_16042,N_13140,N_14479);
nor U16043 (N_16043,N_14080,N_14910);
nand U16044 (N_16044,N_14132,N_13476);
xnor U16045 (N_16045,N_14385,N_12864);
nor U16046 (N_16046,N_12664,N_13332);
nand U16047 (N_16047,N_12628,N_13445);
or U16048 (N_16048,N_13692,N_12799);
nor U16049 (N_16049,N_14235,N_14533);
xnor U16050 (N_16050,N_14432,N_13418);
nand U16051 (N_16051,N_14066,N_14427);
nor U16052 (N_16052,N_12559,N_12954);
and U16053 (N_16053,N_13672,N_14195);
xnor U16054 (N_16054,N_14174,N_12657);
nor U16055 (N_16055,N_14409,N_14936);
xor U16056 (N_16056,N_14787,N_14175);
xnor U16057 (N_16057,N_13720,N_14244);
or U16058 (N_16058,N_12784,N_12903);
and U16059 (N_16059,N_12717,N_14400);
xor U16060 (N_16060,N_14096,N_14726);
or U16061 (N_16061,N_14227,N_13414);
and U16062 (N_16062,N_13544,N_14697);
nand U16063 (N_16063,N_14770,N_12912);
and U16064 (N_16064,N_13062,N_13205);
nand U16065 (N_16065,N_13710,N_12667);
or U16066 (N_16066,N_13727,N_12606);
or U16067 (N_16067,N_13045,N_12640);
nand U16068 (N_16068,N_13821,N_12609);
nand U16069 (N_16069,N_12643,N_12571);
nor U16070 (N_16070,N_13400,N_14048);
or U16071 (N_16071,N_13878,N_12637);
and U16072 (N_16072,N_13499,N_14836);
and U16073 (N_16073,N_12718,N_13597);
and U16074 (N_16074,N_12999,N_14379);
nand U16075 (N_16075,N_13781,N_14208);
nand U16076 (N_16076,N_13990,N_13578);
or U16077 (N_16077,N_12626,N_14159);
nand U16078 (N_16078,N_12507,N_13632);
nand U16079 (N_16079,N_14338,N_14957);
nand U16080 (N_16080,N_12818,N_14163);
and U16081 (N_16081,N_13012,N_12852);
and U16082 (N_16082,N_14035,N_12866);
nand U16083 (N_16083,N_14249,N_13477);
xnor U16084 (N_16084,N_14298,N_14553);
nor U16085 (N_16085,N_14488,N_13685);
nor U16086 (N_16086,N_13898,N_14030);
nand U16087 (N_16087,N_12829,N_13596);
nor U16088 (N_16088,N_14431,N_14692);
xnor U16089 (N_16089,N_13492,N_13673);
nand U16090 (N_16090,N_14756,N_12710);
or U16091 (N_16091,N_13870,N_14918);
and U16092 (N_16092,N_14617,N_14808);
or U16093 (N_16093,N_14701,N_13682);
xnor U16094 (N_16094,N_14160,N_14268);
and U16095 (N_16095,N_14482,N_12625);
and U16096 (N_16096,N_12750,N_13179);
xnor U16097 (N_16097,N_14005,N_14979);
nor U16098 (N_16098,N_14825,N_13298);
nand U16099 (N_16099,N_14441,N_13264);
nand U16100 (N_16100,N_12962,N_14589);
nand U16101 (N_16101,N_13369,N_13758);
nor U16102 (N_16102,N_12855,N_14994);
nor U16103 (N_16103,N_12845,N_14904);
xor U16104 (N_16104,N_14850,N_14613);
xnor U16105 (N_16105,N_13359,N_13475);
nor U16106 (N_16106,N_12781,N_14128);
nand U16107 (N_16107,N_14443,N_14141);
and U16108 (N_16108,N_13273,N_13237);
xnor U16109 (N_16109,N_13753,N_13055);
nand U16110 (N_16110,N_12688,N_13772);
nand U16111 (N_16111,N_14138,N_13765);
xnor U16112 (N_16112,N_13151,N_12760);
nor U16113 (N_16113,N_14463,N_13591);
or U16114 (N_16114,N_14151,N_13552);
nand U16115 (N_16115,N_13317,N_12701);
or U16116 (N_16116,N_14840,N_14357);
nand U16117 (N_16117,N_14917,N_13429);
and U16118 (N_16118,N_13338,N_12967);
xor U16119 (N_16119,N_13412,N_12851);
and U16120 (N_16120,N_14789,N_14188);
or U16121 (N_16121,N_14004,N_13037);
or U16122 (N_16122,N_13007,N_13950);
nor U16123 (N_16123,N_13190,N_13962);
xnor U16124 (N_16124,N_13991,N_12918);
nor U16125 (N_16125,N_13108,N_12575);
xor U16126 (N_16126,N_13840,N_12735);
and U16127 (N_16127,N_13143,N_13558);
nor U16128 (N_16128,N_13214,N_13024);
nor U16129 (N_16129,N_13046,N_14206);
xor U16130 (N_16130,N_14137,N_13345);
nor U16131 (N_16131,N_13527,N_13409);
xor U16132 (N_16132,N_14883,N_13386);
xor U16133 (N_16133,N_12956,N_13240);
xnor U16134 (N_16134,N_13540,N_14086);
nor U16135 (N_16135,N_13168,N_12525);
nor U16136 (N_16136,N_12593,N_14362);
and U16137 (N_16137,N_14270,N_14516);
nand U16138 (N_16138,N_14767,N_14952);
and U16139 (N_16139,N_12786,N_12613);
nor U16140 (N_16140,N_13461,N_14027);
nand U16141 (N_16141,N_13393,N_14378);
or U16142 (N_16142,N_14723,N_12993);
nor U16143 (N_16143,N_13292,N_12537);
nor U16144 (N_16144,N_12744,N_14642);
nand U16145 (N_16145,N_12630,N_14216);
xor U16146 (N_16146,N_14853,N_13805);
or U16147 (N_16147,N_14331,N_13132);
xor U16148 (N_16148,N_12623,N_14725);
xnor U16149 (N_16149,N_13147,N_13118);
or U16150 (N_16150,N_13028,N_13449);
or U16151 (N_16151,N_14722,N_14522);
nand U16152 (N_16152,N_14784,N_13739);
or U16153 (N_16153,N_13730,N_13899);
xor U16154 (N_16154,N_13953,N_14841);
or U16155 (N_16155,N_13057,N_12546);
xnor U16156 (N_16156,N_14384,N_12504);
and U16157 (N_16157,N_14439,N_13258);
xnor U16158 (N_16158,N_13395,N_14908);
and U16159 (N_16159,N_14845,N_13422);
nor U16160 (N_16160,N_14205,N_14891);
or U16161 (N_16161,N_14221,N_13662);
and U16162 (N_16162,N_14383,N_14108);
xor U16163 (N_16163,N_13312,N_13625);
xor U16164 (N_16164,N_12745,N_13528);
nor U16165 (N_16165,N_14600,N_12712);
and U16166 (N_16166,N_12926,N_14473);
or U16167 (N_16167,N_12988,N_14629);
or U16168 (N_16168,N_12843,N_13224);
nor U16169 (N_16169,N_14968,N_14209);
nand U16170 (N_16170,N_14544,N_12616);
nand U16171 (N_16171,N_13027,N_13198);
and U16172 (N_16172,N_12634,N_12904);
xor U16173 (N_16173,N_12671,N_14646);
or U16174 (N_16174,N_14218,N_12973);
and U16175 (N_16175,N_14164,N_12516);
xor U16176 (N_16176,N_14363,N_13675);
nand U16177 (N_16177,N_13091,N_13094);
nor U16178 (N_16178,N_13943,N_14981);
nand U16179 (N_16179,N_14368,N_13670);
or U16180 (N_16180,N_13085,N_14420);
xor U16181 (N_16181,N_14946,N_14852);
nand U16182 (N_16182,N_13197,N_13178);
nor U16183 (N_16183,N_14023,N_12697);
xnor U16184 (N_16184,N_13749,N_14511);
nor U16185 (N_16185,N_14707,N_14016);
nor U16186 (N_16186,N_14119,N_14967);
nand U16187 (N_16187,N_13181,N_12728);
nand U16188 (N_16188,N_13038,N_12685);
or U16189 (N_16189,N_13785,N_12589);
and U16190 (N_16190,N_12569,N_13280);
or U16191 (N_16191,N_12638,N_13225);
and U16192 (N_16192,N_13349,N_14903);
or U16193 (N_16193,N_12726,N_13352);
nor U16194 (N_16194,N_13605,N_14774);
or U16195 (N_16195,N_12724,N_13042);
xor U16196 (N_16196,N_14644,N_14391);
nand U16197 (N_16197,N_13636,N_13808);
or U16198 (N_16198,N_12874,N_12908);
nor U16199 (N_16199,N_14978,N_13799);
xnor U16200 (N_16200,N_13543,N_13104);
nor U16201 (N_16201,N_14014,N_13854);
nor U16202 (N_16202,N_12788,N_13245);
and U16203 (N_16203,N_14258,N_14537);
xor U16204 (N_16204,N_14925,N_14660);
and U16205 (N_16205,N_14530,N_14154);
and U16206 (N_16206,N_12689,N_12905);
nor U16207 (N_16207,N_13602,N_14127);
xnor U16208 (N_16208,N_14053,N_12680);
or U16209 (N_16209,N_14102,N_13768);
nand U16210 (N_16210,N_14120,N_14426);
nand U16211 (N_16211,N_13311,N_13339);
and U16212 (N_16212,N_12646,N_13645);
nor U16213 (N_16213,N_13538,N_13633);
nor U16214 (N_16214,N_13818,N_14863);
xor U16215 (N_16215,N_14242,N_12727);
nor U16216 (N_16216,N_13348,N_14548);
nand U16217 (N_16217,N_12740,N_13930);
and U16218 (N_16218,N_12567,N_14340);
nand U16219 (N_16219,N_14240,N_13897);
xnor U16220 (N_16220,N_14974,N_12723);
xor U16221 (N_16221,N_13063,N_14576);
or U16222 (N_16222,N_14202,N_13282);
nor U16223 (N_16223,N_14969,N_13614);
nand U16224 (N_16224,N_13693,N_13183);
and U16225 (N_16225,N_14577,N_14490);
and U16226 (N_16226,N_13624,N_14645);
xor U16227 (N_16227,N_14477,N_13413);
or U16228 (N_16228,N_12586,N_14303);
and U16229 (N_16229,N_13992,N_14358);
and U16230 (N_16230,N_14219,N_13331);
xor U16231 (N_16231,N_14878,N_14993);
nor U16232 (N_16232,N_14684,N_14448);
nor U16233 (N_16233,N_14019,N_13428);
nand U16234 (N_16234,N_12624,N_13061);
xnor U16235 (N_16235,N_13304,N_13623);
or U16236 (N_16236,N_12661,N_13396);
or U16237 (N_16237,N_14536,N_14000);
or U16238 (N_16238,N_14909,N_13570);
nor U16239 (N_16239,N_14106,N_14673);
xnor U16240 (N_16240,N_14095,N_13864);
nand U16241 (N_16241,N_14162,N_12811);
and U16242 (N_16242,N_14017,N_13640);
xnor U16243 (N_16243,N_13262,N_13948);
nand U16244 (N_16244,N_12765,N_12713);
nor U16245 (N_16245,N_14796,N_13813);
xor U16246 (N_16246,N_13432,N_14924);
nand U16247 (N_16247,N_14519,N_12938);
nand U16248 (N_16248,N_14010,N_13719);
nand U16249 (N_16249,N_12526,N_12948);
nor U16250 (N_16250,N_13630,N_13907);
and U16251 (N_16251,N_13868,N_14823);
nand U16252 (N_16252,N_13318,N_13613);
or U16253 (N_16253,N_13977,N_13724);
or U16254 (N_16254,N_13120,N_13876);
and U16255 (N_16255,N_13865,N_13150);
and U16256 (N_16256,N_13476,N_12520);
and U16257 (N_16257,N_13588,N_13665);
and U16258 (N_16258,N_14941,N_13188);
nand U16259 (N_16259,N_12901,N_13898);
nor U16260 (N_16260,N_14421,N_12693);
or U16261 (N_16261,N_12880,N_12593);
and U16262 (N_16262,N_13992,N_13391);
nand U16263 (N_16263,N_14172,N_12686);
xnor U16264 (N_16264,N_13708,N_14984);
nor U16265 (N_16265,N_13133,N_12716);
and U16266 (N_16266,N_14743,N_14687);
or U16267 (N_16267,N_14101,N_13105);
and U16268 (N_16268,N_14119,N_14772);
or U16269 (N_16269,N_12579,N_13095);
or U16270 (N_16270,N_12897,N_14990);
nor U16271 (N_16271,N_13321,N_12710);
xor U16272 (N_16272,N_12666,N_13831);
and U16273 (N_16273,N_13345,N_13883);
nand U16274 (N_16274,N_14394,N_14791);
nand U16275 (N_16275,N_14310,N_13380);
xor U16276 (N_16276,N_12867,N_13760);
xnor U16277 (N_16277,N_14418,N_13092);
nor U16278 (N_16278,N_13478,N_13548);
and U16279 (N_16279,N_14225,N_14242);
nor U16280 (N_16280,N_12659,N_13948);
or U16281 (N_16281,N_14916,N_14002);
or U16282 (N_16282,N_14851,N_13356);
xnor U16283 (N_16283,N_13127,N_12725);
xnor U16284 (N_16284,N_13782,N_14409);
and U16285 (N_16285,N_13113,N_14325);
and U16286 (N_16286,N_13240,N_13992);
and U16287 (N_16287,N_14785,N_13375);
nand U16288 (N_16288,N_14177,N_14747);
xnor U16289 (N_16289,N_12628,N_14256);
nor U16290 (N_16290,N_14508,N_13427);
xor U16291 (N_16291,N_13439,N_13607);
nor U16292 (N_16292,N_14498,N_13975);
or U16293 (N_16293,N_13775,N_13831);
or U16294 (N_16294,N_14099,N_12659);
nor U16295 (N_16295,N_14839,N_14227);
nor U16296 (N_16296,N_12873,N_13380);
or U16297 (N_16297,N_13325,N_14590);
or U16298 (N_16298,N_12705,N_13392);
nand U16299 (N_16299,N_13259,N_14187);
xnor U16300 (N_16300,N_14129,N_12872);
nor U16301 (N_16301,N_13774,N_14345);
and U16302 (N_16302,N_13400,N_12919);
or U16303 (N_16303,N_12968,N_13174);
or U16304 (N_16304,N_14332,N_13227);
nand U16305 (N_16305,N_14327,N_13633);
xnor U16306 (N_16306,N_13146,N_13283);
nand U16307 (N_16307,N_14507,N_13006);
or U16308 (N_16308,N_14284,N_12943);
or U16309 (N_16309,N_13707,N_12663);
and U16310 (N_16310,N_13304,N_13751);
or U16311 (N_16311,N_14268,N_12668);
xor U16312 (N_16312,N_12605,N_13177);
and U16313 (N_16313,N_14223,N_14683);
nand U16314 (N_16314,N_13023,N_13772);
nor U16315 (N_16315,N_13501,N_13955);
xnor U16316 (N_16316,N_13612,N_13853);
and U16317 (N_16317,N_12842,N_13343);
nand U16318 (N_16318,N_12734,N_13642);
and U16319 (N_16319,N_14523,N_12641);
xor U16320 (N_16320,N_13205,N_13164);
and U16321 (N_16321,N_13425,N_14599);
and U16322 (N_16322,N_13828,N_14700);
or U16323 (N_16323,N_14481,N_12716);
xnor U16324 (N_16324,N_14196,N_14838);
and U16325 (N_16325,N_14259,N_12899);
nor U16326 (N_16326,N_14549,N_12667);
nor U16327 (N_16327,N_13691,N_14637);
and U16328 (N_16328,N_14702,N_13409);
nor U16329 (N_16329,N_13766,N_14513);
xnor U16330 (N_16330,N_13400,N_13582);
xor U16331 (N_16331,N_12729,N_14717);
xor U16332 (N_16332,N_14707,N_12989);
nand U16333 (N_16333,N_13082,N_14317);
xor U16334 (N_16334,N_13602,N_12985);
xor U16335 (N_16335,N_12801,N_14222);
or U16336 (N_16336,N_14684,N_13559);
nand U16337 (N_16337,N_14193,N_13978);
or U16338 (N_16338,N_14910,N_13196);
xnor U16339 (N_16339,N_13525,N_13749);
xor U16340 (N_16340,N_13693,N_14671);
xnor U16341 (N_16341,N_14369,N_14822);
nand U16342 (N_16342,N_12597,N_13269);
or U16343 (N_16343,N_13672,N_14660);
xnor U16344 (N_16344,N_12569,N_12632);
nand U16345 (N_16345,N_12744,N_13234);
nor U16346 (N_16346,N_13987,N_13651);
and U16347 (N_16347,N_14500,N_13416);
xor U16348 (N_16348,N_14079,N_12621);
and U16349 (N_16349,N_14375,N_14832);
or U16350 (N_16350,N_12861,N_12549);
nor U16351 (N_16351,N_12937,N_12651);
nor U16352 (N_16352,N_12746,N_13510);
or U16353 (N_16353,N_14470,N_13514);
nor U16354 (N_16354,N_14563,N_12970);
nand U16355 (N_16355,N_13986,N_12956);
nor U16356 (N_16356,N_12922,N_12866);
nand U16357 (N_16357,N_14574,N_12756);
xor U16358 (N_16358,N_14716,N_13628);
and U16359 (N_16359,N_13760,N_13375);
nor U16360 (N_16360,N_13468,N_12548);
nand U16361 (N_16361,N_13590,N_14409);
nand U16362 (N_16362,N_14077,N_13814);
nand U16363 (N_16363,N_13070,N_14676);
nand U16364 (N_16364,N_14277,N_12538);
nand U16365 (N_16365,N_12948,N_14329);
nor U16366 (N_16366,N_13024,N_13374);
and U16367 (N_16367,N_14001,N_12954);
nor U16368 (N_16368,N_14522,N_14711);
or U16369 (N_16369,N_14695,N_13002);
nand U16370 (N_16370,N_13578,N_13091);
and U16371 (N_16371,N_14876,N_14873);
nand U16372 (N_16372,N_12891,N_14267);
and U16373 (N_16373,N_14751,N_14414);
xnor U16374 (N_16374,N_14477,N_14561);
xor U16375 (N_16375,N_13838,N_13014);
nor U16376 (N_16376,N_13182,N_12662);
xor U16377 (N_16377,N_14035,N_12754);
nor U16378 (N_16378,N_14959,N_14925);
nor U16379 (N_16379,N_13361,N_13633);
nand U16380 (N_16380,N_14283,N_14844);
and U16381 (N_16381,N_12820,N_13000);
nand U16382 (N_16382,N_14813,N_14483);
nand U16383 (N_16383,N_13357,N_14641);
nor U16384 (N_16384,N_14082,N_12535);
or U16385 (N_16385,N_14413,N_14412);
nand U16386 (N_16386,N_14817,N_12628);
nor U16387 (N_16387,N_13682,N_13480);
nor U16388 (N_16388,N_13452,N_12621);
or U16389 (N_16389,N_14519,N_14597);
nor U16390 (N_16390,N_14383,N_13939);
and U16391 (N_16391,N_14685,N_13757);
xnor U16392 (N_16392,N_12583,N_12846);
xor U16393 (N_16393,N_12695,N_13093);
or U16394 (N_16394,N_12838,N_13450);
nand U16395 (N_16395,N_13929,N_12983);
nand U16396 (N_16396,N_14102,N_12799);
or U16397 (N_16397,N_13528,N_13258);
and U16398 (N_16398,N_13287,N_14655);
xnor U16399 (N_16399,N_12791,N_13792);
nand U16400 (N_16400,N_14565,N_12852);
nor U16401 (N_16401,N_13505,N_13803);
and U16402 (N_16402,N_14823,N_13382);
nor U16403 (N_16403,N_13254,N_14535);
and U16404 (N_16404,N_14037,N_12524);
or U16405 (N_16405,N_13928,N_12528);
or U16406 (N_16406,N_12545,N_13095);
nand U16407 (N_16407,N_14428,N_13451);
nor U16408 (N_16408,N_12858,N_13016);
xor U16409 (N_16409,N_12578,N_14116);
nand U16410 (N_16410,N_14922,N_12673);
nand U16411 (N_16411,N_14280,N_12659);
nor U16412 (N_16412,N_13159,N_13322);
and U16413 (N_16413,N_13289,N_13113);
nand U16414 (N_16414,N_13408,N_13946);
nor U16415 (N_16415,N_13197,N_13414);
and U16416 (N_16416,N_14242,N_13474);
nand U16417 (N_16417,N_14273,N_13157);
nand U16418 (N_16418,N_12561,N_12604);
xnor U16419 (N_16419,N_13938,N_14725);
xnor U16420 (N_16420,N_13489,N_13434);
or U16421 (N_16421,N_14209,N_12771);
xnor U16422 (N_16422,N_14206,N_13826);
nor U16423 (N_16423,N_13532,N_13734);
and U16424 (N_16424,N_12778,N_13400);
and U16425 (N_16425,N_14948,N_13489);
and U16426 (N_16426,N_13891,N_12862);
and U16427 (N_16427,N_12838,N_13798);
and U16428 (N_16428,N_13263,N_13196);
and U16429 (N_16429,N_13355,N_12564);
nand U16430 (N_16430,N_14980,N_12816);
nand U16431 (N_16431,N_14490,N_14695);
nor U16432 (N_16432,N_12610,N_12564);
and U16433 (N_16433,N_13796,N_13350);
or U16434 (N_16434,N_13052,N_13222);
and U16435 (N_16435,N_13454,N_12823);
and U16436 (N_16436,N_14768,N_12780);
xnor U16437 (N_16437,N_14609,N_13545);
nand U16438 (N_16438,N_13064,N_14118);
xor U16439 (N_16439,N_14306,N_13245);
xor U16440 (N_16440,N_12982,N_13135);
nand U16441 (N_16441,N_12790,N_13793);
or U16442 (N_16442,N_13508,N_13026);
or U16443 (N_16443,N_14566,N_14590);
nor U16444 (N_16444,N_14365,N_12517);
and U16445 (N_16445,N_14319,N_14390);
xnor U16446 (N_16446,N_14768,N_13326);
nand U16447 (N_16447,N_12839,N_13845);
nand U16448 (N_16448,N_14026,N_12750);
nor U16449 (N_16449,N_13732,N_13568);
and U16450 (N_16450,N_14649,N_12870);
nor U16451 (N_16451,N_14636,N_12663);
nor U16452 (N_16452,N_14757,N_14719);
nand U16453 (N_16453,N_14421,N_12561);
nor U16454 (N_16454,N_13232,N_12627);
or U16455 (N_16455,N_13913,N_13922);
nand U16456 (N_16456,N_12754,N_13124);
xnor U16457 (N_16457,N_14898,N_14875);
or U16458 (N_16458,N_14576,N_13844);
xor U16459 (N_16459,N_14063,N_14351);
nand U16460 (N_16460,N_14615,N_12735);
nand U16461 (N_16461,N_12938,N_12589);
nand U16462 (N_16462,N_14527,N_14210);
nor U16463 (N_16463,N_12538,N_14523);
nand U16464 (N_16464,N_14806,N_12680);
or U16465 (N_16465,N_14299,N_14958);
nor U16466 (N_16466,N_12651,N_12918);
or U16467 (N_16467,N_14844,N_12845);
or U16468 (N_16468,N_12993,N_14947);
nor U16469 (N_16469,N_13365,N_12719);
nand U16470 (N_16470,N_14325,N_13664);
xor U16471 (N_16471,N_14462,N_13348);
nand U16472 (N_16472,N_12648,N_13929);
or U16473 (N_16473,N_14975,N_13247);
or U16474 (N_16474,N_14218,N_14608);
nor U16475 (N_16475,N_12573,N_14441);
nand U16476 (N_16476,N_12532,N_12980);
xnor U16477 (N_16477,N_14588,N_12809);
nor U16478 (N_16478,N_13942,N_12916);
and U16479 (N_16479,N_14549,N_13126);
xor U16480 (N_16480,N_13689,N_12867);
and U16481 (N_16481,N_12517,N_13809);
xnor U16482 (N_16482,N_14370,N_14040);
and U16483 (N_16483,N_12695,N_13263);
or U16484 (N_16484,N_13071,N_12898);
nor U16485 (N_16485,N_13124,N_14850);
xnor U16486 (N_16486,N_14361,N_13964);
xor U16487 (N_16487,N_12501,N_13502);
nand U16488 (N_16488,N_12607,N_13338);
or U16489 (N_16489,N_14228,N_13490);
nor U16490 (N_16490,N_14143,N_13779);
nand U16491 (N_16491,N_13135,N_13518);
or U16492 (N_16492,N_12884,N_12886);
xor U16493 (N_16493,N_13604,N_14720);
xnor U16494 (N_16494,N_14866,N_14865);
nor U16495 (N_16495,N_13672,N_13393);
xnor U16496 (N_16496,N_14223,N_14229);
nor U16497 (N_16497,N_13219,N_14582);
or U16498 (N_16498,N_12982,N_13639);
and U16499 (N_16499,N_13958,N_13820);
xnor U16500 (N_16500,N_14689,N_13077);
and U16501 (N_16501,N_12983,N_14622);
nand U16502 (N_16502,N_14706,N_14980);
and U16503 (N_16503,N_14574,N_12607);
and U16504 (N_16504,N_13485,N_14879);
nand U16505 (N_16505,N_14849,N_12953);
xnor U16506 (N_16506,N_14599,N_14721);
xor U16507 (N_16507,N_14433,N_14642);
nand U16508 (N_16508,N_14522,N_13441);
xor U16509 (N_16509,N_13475,N_14736);
and U16510 (N_16510,N_14130,N_14473);
and U16511 (N_16511,N_14374,N_12803);
or U16512 (N_16512,N_12688,N_13046);
nor U16513 (N_16513,N_12941,N_13841);
or U16514 (N_16514,N_14708,N_13787);
or U16515 (N_16515,N_13916,N_13921);
or U16516 (N_16516,N_13324,N_13989);
nor U16517 (N_16517,N_13311,N_12807);
nand U16518 (N_16518,N_13214,N_13249);
xor U16519 (N_16519,N_12818,N_14815);
and U16520 (N_16520,N_13222,N_13119);
or U16521 (N_16521,N_12873,N_13213);
nand U16522 (N_16522,N_13191,N_13339);
nor U16523 (N_16523,N_14476,N_12891);
and U16524 (N_16524,N_14406,N_13849);
nand U16525 (N_16525,N_13710,N_12826);
nand U16526 (N_16526,N_12858,N_13960);
nand U16527 (N_16527,N_14053,N_13735);
and U16528 (N_16528,N_13951,N_12911);
and U16529 (N_16529,N_13709,N_13615);
nor U16530 (N_16530,N_13334,N_14040);
nor U16531 (N_16531,N_14978,N_13202);
xor U16532 (N_16532,N_13710,N_14804);
and U16533 (N_16533,N_14045,N_12992);
xnor U16534 (N_16534,N_13208,N_12924);
or U16535 (N_16535,N_14860,N_14880);
nand U16536 (N_16536,N_13107,N_13153);
nand U16537 (N_16537,N_14632,N_13996);
and U16538 (N_16538,N_14859,N_13211);
nand U16539 (N_16539,N_14862,N_13556);
nand U16540 (N_16540,N_14678,N_14147);
nand U16541 (N_16541,N_13158,N_13052);
nand U16542 (N_16542,N_12989,N_13542);
xor U16543 (N_16543,N_13206,N_13970);
and U16544 (N_16544,N_13980,N_13583);
xor U16545 (N_16545,N_13709,N_14726);
and U16546 (N_16546,N_12788,N_13347);
and U16547 (N_16547,N_12766,N_13214);
nor U16548 (N_16548,N_12695,N_14516);
and U16549 (N_16549,N_13086,N_14858);
nand U16550 (N_16550,N_13282,N_13255);
nor U16551 (N_16551,N_12625,N_14628);
nand U16552 (N_16552,N_13480,N_14191);
nand U16553 (N_16553,N_12548,N_13915);
xor U16554 (N_16554,N_14893,N_14834);
and U16555 (N_16555,N_14207,N_14655);
xnor U16556 (N_16556,N_13135,N_12763);
or U16557 (N_16557,N_13180,N_13909);
nor U16558 (N_16558,N_13696,N_12856);
xnor U16559 (N_16559,N_12874,N_14768);
or U16560 (N_16560,N_12724,N_13693);
nor U16561 (N_16561,N_14848,N_13039);
and U16562 (N_16562,N_14593,N_12690);
or U16563 (N_16563,N_13349,N_13630);
and U16564 (N_16564,N_14245,N_14074);
or U16565 (N_16565,N_13013,N_12756);
nand U16566 (N_16566,N_14979,N_14703);
and U16567 (N_16567,N_13684,N_12789);
nand U16568 (N_16568,N_14515,N_14290);
xor U16569 (N_16569,N_14944,N_12906);
xor U16570 (N_16570,N_12827,N_13203);
or U16571 (N_16571,N_14579,N_13255);
or U16572 (N_16572,N_14672,N_12756);
and U16573 (N_16573,N_14042,N_14185);
nor U16574 (N_16574,N_13592,N_12679);
nor U16575 (N_16575,N_14768,N_13966);
xor U16576 (N_16576,N_14371,N_13079);
and U16577 (N_16577,N_12962,N_14769);
or U16578 (N_16578,N_12964,N_14944);
nand U16579 (N_16579,N_14912,N_13598);
and U16580 (N_16580,N_13177,N_14163);
nand U16581 (N_16581,N_13018,N_14184);
xnor U16582 (N_16582,N_14273,N_13073);
or U16583 (N_16583,N_14603,N_13895);
nor U16584 (N_16584,N_14735,N_14671);
nor U16585 (N_16585,N_14460,N_12858);
xor U16586 (N_16586,N_12526,N_12866);
nor U16587 (N_16587,N_12703,N_13163);
and U16588 (N_16588,N_13640,N_14973);
or U16589 (N_16589,N_13625,N_12904);
or U16590 (N_16590,N_14835,N_14924);
or U16591 (N_16591,N_13004,N_14168);
xor U16592 (N_16592,N_13695,N_12930);
and U16593 (N_16593,N_14290,N_12578);
or U16594 (N_16594,N_14363,N_14102);
or U16595 (N_16595,N_13422,N_13104);
nand U16596 (N_16596,N_14611,N_14830);
xor U16597 (N_16597,N_13430,N_13514);
nand U16598 (N_16598,N_12826,N_14045);
nand U16599 (N_16599,N_14195,N_13490);
or U16600 (N_16600,N_13544,N_12501);
or U16601 (N_16601,N_12520,N_14907);
xor U16602 (N_16602,N_13368,N_13184);
or U16603 (N_16603,N_13247,N_13127);
and U16604 (N_16604,N_13646,N_14020);
or U16605 (N_16605,N_14446,N_12962);
nand U16606 (N_16606,N_13684,N_13999);
or U16607 (N_16607,N_14098,N_12760);
xor U16608 (N_16608,N_13336,N_13638);
or U16609 (N_16609,N_13377,N_14935);
or U16610 (N_16610,N_13118,N_13300);
nor U16611 (N_16611,N_14222,N_14359);
nor U16612 (N_16612,N_12639,N_14764);
xnor U16613 (N_16613,N_13076,N_14352);
or U16614 (N_16614,N_13228,N_14907);
nor U16615 (N_16615,N_12798,N_13658);
and U16616 (N_16616,N_13511,N_14908);
and U16617 (N_16617,N_12507,N_12912);
xnor U16618 (N_16618,N_14903,N_14105);
nor U16619 (N_16619,N_12862,N_13220);
nand U16620 (N_16620,N_12506,N_14632);
or U16621 (N_16621,N_13245,N_14069);
nand U16622 (N_16622,N_13759,N_14940);
or U16623 (N_16623,N_14622,N_12514);
or U16624 (N_16624,N_13282,N_13095);
nor U16625 (N_16625,N_14450,N_13263);
nor U16626 (N_16626,N_12909,N_14785);
nand U16627 (N_16627,N_13767,N_13035);
xnor U16628 (N_16628,N_14097,N_12809);
xnor U16629 (N_16629,N_14861,N_14216);
xor U16630 (N_16630,N_13382,N_13149);
or U16631 (N_16631,N_13676,N_14906);
nor U16632 (N_16632,N_14910,N_13975);
and U16633 (N_16633,N_14386,N_13746);
or U16634 (N_16634,N_13189,N_13101);
xor U16635 (N_16635,N_12736,N_14877);
nor U16636 (N_16636,N_14153,N_13233);
nand U16637 (N_16637,N_12928,N_13289);
nand U16638 (N_16638,N_13169,N_14605);
nor U16639 (N_16639,N_13120,N_12809);
and U16640 (N_16640,N_14490,N_14820);
or U16641 (N_16641,N_13417,N_14034);
xor U16642 (N_16642,N_14587,N_14623);
and U16643 (N_16643,N_14225,N_12941);
nor U16644 (N_16644,N_13183,N_13894);
nand U16645 (N_16645,N_14188,N_14518);
and U16646 (N_16646,N_13392,N_13427);
and U16647 (N_16647,N_13770,N_14711);
and U16648 (N_16648,N_12633,N_13331);
xnor U16649 (N_16649,N_13132,N_13121);
nor U16650 (N_16650,N_13326,N_12849);
xor U16651 (N_16651,N_14782,N_12772);
nand U16652 (N_16652,N_13338,N_13318);
nand U16653 (N_16653,N_12599,N_12842);
xor U16654 (N_16654,N_14505,N_12689);
or U16655 (N_16655,N_14720,N_13949);
or U16656 (N_16656,N_14019,N_14526);
and U16657 (N_16657,N_13076,N_13127);
nand U16658 (N_16658,N_12653,N_14957);
nor U16659 (N_16659,N_14250,N_12867);
xor U16660 (N_16660,N_13047,N_13271);
xor U16661 (N_16661,N_12669,N_14820);
nand U16662 (N_16662,N_13818,N_13613);
and U16663 (N_16663,N_12512,N_14433);
nand U16664 (N_16664,N_14146,N_13977);
and U16665 (N_16665,N_13053,N_13919);
nand U16666 (N_16666,N_14639,N_13586);
nor U16667 (N_16667,N_13284,N_14874);
or U16668 (N_16668,N_12951,N_13330);
nand U16669 (N_16669,N_12505,N_13064);
nand U16670 (N_16670,N_13060,N_13864);
xnor U16671 (N_16671,N_13926,N_14739);
and U16672 (N_16672,N_13650,N_13537);
nor U16673 (N_16673,N_13276,N_14816);
nor U16674 (N_16674,N_14069,N_14874);
or U16675 (N_16675,N_14718,N_12734);
and U16676 (N_16676,N_14352,N_12714);
nor U16677 (N_16677,N_12544,N_14781);
or U16678 (N_16678,N_14721,N_13067);
or U16679 (N_16679,N_14291,N_13421);
nor U16680 (N_16680,N_12986,N_13009);
or U16681 (N_16681,N_14284,N_12616);
nor U16682 (N_16682,N_14215,N_14137);
nand U16683 (N_16683,N_13906,N_13496);
and U16684 (N_16684,N_12622,N_13779);
and U16685 (N_16685,N_14290,N_14848);
nor U16686 (N_16686,N_14248,N_13693);
nor U16687 (N_16687,N_13567,N_13123);
nand U16688 (N_16688,N_12832,N_13135);
xnor U16689 (N_16689,N_14904,N_12868);
xnor U16690 (N_16690,N_13347,N_13431);
nand U16691 (N_16691,N_12967,N_13125);
or U16692 (N_16692,N_14147,N_14836);
and U16693 (N_16693,N_14510,N_12641);
and U16694 (N_16694,N_14796,N_14620);
or U16695 (N_16695,N_13565,N_14882);
and U16696 (N_16696,N_14355,N_12707);
nor U16697 (N_16697,N_13947,N_14633);
xnor U16698 (N_16698,N_12937,N_12555);
and U16699 (N_16699,N_13206,N_14460);
and U16700 (N_16700,N_14330,N_14157);
and U16701 (N_16701,N_14450,N_13000);
and U16702 (N_16702,N_13026,N_14895);
and U16703 (N_16703,N_13533,N_14759);
nand U16704 (N_16704,N_12661,N_12577);
xnor U16705 (N_16705,N_13711,N_12657);
nor U16706 (N_16706,N_14605,N_12982);
or U16707 (N_16707,N_13244,N_12506);
and U16708 (N_16708,N_13120,N_14210);
and U16709 (N_16709,N_12514,N_14228);
or U16710 (N_16710,N_14060,N_14858);
or U16711 (N_16711,N_13505,N_13756);
nor U16712 (N_16712,N_12880,N_12981);
or U16713 (N_16713,N_13956,N_14817);
and U16714 (N_16714,N_13987,N_13909);
xor U16715 (N_16715,N_13745,N_12559);
and U16716 (N_16716,N_14264,N_13081);
and U16717 (N_16717,N_14591,N_12663);
nor U16718 (N_16718,N_13703,N_13052);
nand U16719 (N_16719,N_14609,N_14913);
xor U16720 (N_16720,N_12994,N_12581);
or U16721 (N_16721,N_14170,N_14711);
and U16722 (N_16722,N_13415,N_13877);
xnor U16723 (N_16723,N_13014,N_13085);
and U16724 (N_16724,N_14649,N_12966);
xnor U16725 (N_16725,N_12826,N_12776);
and U16726 (N_16726,N_14297,N_14059);
nor U16727 (N_16727,N_14330,N_13341);
or U16728 (N_16728,N_14367,N_14821);
nor U16729 (N_16729,N_14822,N_13872);
xnor U16730 (N_16730,N_14840,N_14320);
nand U16731 (N_16731,N_14396,N_12602);
nand U16732 (N_16732,N_13240,N_13612);
or U16733 (N_16733,N_14630,N_14360);
or U16734 (N_16734,N_14477,N_12621);
nor U16735 (N_16735,N_13021,N_14441);
or U16736 (N_16736,N_13286,N_12626);
nand U16737 (N_16737,N_13912,N_12897);
and U16738 (N_16738,N_13106,N_14946);
or U16739 (N_16739,N_14474,N_12786);
and U16740 (N_16740,N_14015,N_13161);
nor U16741 (N_16741,N_13989,N_13889);
nand U16742 (N_16742,N_13593,N_13612);
nor U16743 (N_16743,N_14607,N_12536);
xnor U16744 (N_16744,N_14013,N_14858);
and U16745 (N_16745,N_12688,N_14259);
nand U16746 (N_16746,N_13691,N_13154);
xnor U16747 (N_16747,N_13990,N_13346);
nand U16748 (N_16748,N_13875,N_12905);
xor U16749 (N_16749,N_13680,N_13765);
xnor U16750 (N_16750,N_14291,N_13639);
nor U16751 (N_16751,N_13794,N_14627);
nor U16752 (N_16752,N_14942,N_13864);
xnor U16753 (N_16753,N_13176,N_14718);
and U16754 (N_16754,N_13880,N_14954);
or U16755 (N_16755,N_14295,N_14282);
or U16756 (N_16756,N_14997,N_14382);
and U16757 (N_16757,N_14823,N_14352);
xnor U16758 (N_16758,N_13741,N_12868);
xnor U16759 (N_16759,N_12539,N_13262);
nor U16760 (N_16760,N_14974,N_14186);
nand U16761 (N_16761,N_14534,N_14497);
nor U16762 (N_16762,N_14709,N_12645);
nand U16763 (N_16763,N_12907,N_13056);
nor U16764 (N_16764,N_13642,N_14392);
or U16765 (N_16765,N_13496,N_12580);
xor U16766 (N_16766,N_14966,N_12710);
xnor U16767 (N_16767,N_12845,N_14632);
xnor U16768 (N_16768,N_12923,N_14891);
and U16769 (N_16769,N_14491,N_14676);
xor U16770 (N_16770,N_13265,N_14527);
and U16771 (N_16771,N_14932,N_13793);
xnor U16772 (N_16772,N_12997,N_12643);
xnor U16773 (N_16773,N_14251,N_14377);
nand U16774 (N_16774,N_13852,N_13000);
and U16775 (N_16775,N_14566,N_12797);
and U16776 (N_16776,N_13993,N_14117);
nand U16777 (N_16777,N_13720,N_14937);
xor U16778 (N_16778,N_14445,N_14891);
nand U16779 (N_16779,N_14612,N_13472);
and U16780 (N_16780,N_14855,N_14282);
xnor U16781 (N_16781,N_14539,N_12785);
and U16782 (N_16782,N_14954,N_13288);
and U16783 (N_16783,N_14248,N_12909);
nand U16784 (N_16784,N_12934,N_14553);
and U16785 (N_16785,N_13146,N_12930);
or U16786 (N_16786,N_13231,N_13651);
and U16787 (N_16787,N_13763,N_14478);
or U16788 (N_16788,N_13076,N_14875);
and U16789 (N_16789,N_14406,N_12623);
xor U16790 (N_16790,N_12514,N_13579);
or U16791 (N_16791,N_13530,N_13185);
nand U16792 (N_16792,N_14974,N_12550);
nand U16793 (N_16793,N_14814,N_13551);
nor U16794 (N_16794,N_14176,N_13355);
nand U16795 (N_16795,N_14362,N_13211);
xnor U16796 (N_16796,N_13826,N_13284);
or U16797 (N_16797,N_12817,N_13732);
or U16798 (N_16798,N_14368,N_13868);
nand U16799 (N_16799,N_13435,N_13042);
nand U16800 (N_16800,N_13073,N_14300);
xor U16801 (N_16801,N_13066,N_14224);
nand U16802 (N_16802,N_12947,N_13684);
or U16803 (N_16803,N_14730,N_13767);
nand U16804 (N_16804,N_13587,N_14758);
or U16805 (N_16805,N_14239,N_13356);
and U16806 (N_16806,N_12852,N_13306);
nor U16807 (N_16807,N_13247,N_12922);
nand U16808 (N_16808,N_13341,N_14570);
nor U16809 (N_16809,N_13549,N_14980);
nand U16810 (N_16810,N_14398,N_13560);
and U16811 (N_16811,N_13532,N_13404);
xor U16812 (N_16812,N_14254,N_13357);
and U16813 (N_16813,N_14497,N_13994);
or U16814 (N_16814,N_13043,N_12959);
or U16815 (N_16815,N_13175,N_14355);
xor U16816 (N_16816,N_13697,N_12901);
xor U16817 (N_16817,N_14951,N_14841);
and U16818 (N_16818,N_13601,N_13101);
nor U16819 (N_16819,N_14567,N_14990);
or U16820 (N_16820,N_13117,N_13646);
or U16821 (N_16821,N_14597,N_13322);
or U16822 (N_16822,N_14499,N_12712);
nor U16823 (N_16823,N_14902,N_14528);
nand U16824 (N_16824,N_13707,N_12535);
and U16825 (N_16825,N_13569,N_12565);
or U16826 (N_16826,N_13256,N_14959);
and U16827 (N_16827,N_12808,N_12879);
or U16828 (N_16828,N_14902,N_13396);
nand U16829 (N_16829,N_13898,N_13359);
and U16830 (N_16830,N_12922,N_12815);
nand U16831 (N_16831,N_14497,N_14762);
or U16832 (N_16832,N_13114,N_13163);
nand U16833 (N_16833,N_13286,N_12864);
nor U16834 (N_16834,N_14969,N_12567);
nor U16835 (N_16835,N_14281,N_14303);
or U16836 (N_16836,N_12798,N_13027);
nand U16837 (N_16837,N_13800,N_12545);
or U16838 (N_16838,N_13875,N_13946);
and U16839 (N_16839,N_13358,N_13861);
xor U16840 (N_16840,N_14011,N_13751);
nand U16841 (N_16841,N_12845,N_14119);
nand U16842 (N_16842,N_12614,N_12703);
nand U16843 (N_16843,N_13736,N_12511);
or U16844 (N_16844,N_14136,N_14747);
or U16845 (N_16845,N_14222,N_14871);
xor U16846 (N_16846,N_14888,N_12585);
xnor U16847 (N_16847,N_12828,N_13602);
nor U16848 (N_16848,N_13059,N_12973);
xor U16849 (N_16849,N_14713,N_14579);
or U16850 (N_16850,N_13338,N_13911);
or U16851 (N_16851,N_12853,N_14840);
nor U16852 (N_16852,N_12939,N_14015);
xnor U16853 (N_16853,N_14706,N_12824);
nor U16854 (N_16854,N_14603,N_13030);
nand U16855 (N_16855,N_14277,N_13770);
and U16856 (N_16856,N_13448,N_13996);
and U16857 (N_16857,N_14136,N_13004);
nand U16858 (N_16858,N_14420,N_14964);
nor U16859 (N_16859,N_14088,N_14304);
xor U16860 (N_16860,N_14439,N_13173);
xor U16861 (N_16861,N_14596,N_13920);
or U16862 (N_16862,N_14469,N_14867);
or U16863 (N_16863,N_13428,N_13647);
or U16864 (N_16864,N_12705,N_14329);
and U16865 (N_16865,N_14864,N_14006);
and U16866 (N_16866,N_13497,N_14560);
or U16867 (N_16867,N_13254,N_12754);
or U16868 (N_16868,N_12881,N_13373);
nand U16869 (N_16869,N_12749,N_13350);
xnor U16870 (N_16870,N_13033,N_14700);
xnor U16871 (N_16871,N_12682,N_12750);
nor U16872 (N_16872,N_13083,N_12853);
nand U16873 (N_16873,N_12590,N_13587);
and U16874 (N_16874,N_12692,N_13652);
xor U16875 (N_16875,N_14396,N_12639);
nand U16876 (N_16876,N_13315,N_12884);
and U16877 (N_16877,N_13216,N_14112);
or U16878 (N_16878,N_14211,N_14131);
or U16879 (N_16879,N_12533,N_14326);
xor U16880 (N_16880,N_13853,N_13872);
and U16881 (N_16881,N_13682,N_14755);
and U16882 (N_16882,N_14121,N_14279);
nand U16883 (N_16883,N_14728,N_14188);
or U16884 (N_16884,N_14180,N_13145);
and U16885 (N_16885,N_14162,N_13759);
and U16886 (N_16886,N_13956,N_12685);
and U16887 (N_16887,N_14903,N_14449);
xnor U16888 (N_16888,N_13093,N_12954);
nand U16889 (N_16889,N_14595,N_12954);
nand U16890 (N_16890,N_13667,N_14612);
and U16891 (N_16891,N_13537,N_13126);
or U16892 (N_16892,N_13512,N_14187);
nor U16893 (N_16893,N_13853,N_13431);
and U16894 (N_16894,N_14548,N_13115);
nand U16895 (N_16895,N_14491,N_14477);
nor U16896 (N_16896,N_14742,N_13889);
or U16897 (N_16897,N_13939,N_13614);
or U16898 (N_16898,N_14382,N_14751);
or U16899 (N_16899,N_14506,N_13305);
nand U16900 (N_16900,N_13230,N_13757);
or U16901 (N_16901,N_13929,N_13924);
nor U16902 (N_16902,N_13347,N_14778);
and U16903 (N_16903,N_13410,N_13188);
nand U16904 (N_16904,N_14162,N_12964);
nand U16905 (N_16905,N_14343,N_12830);
nor U16906 (N_16906,N_14118,N_13533);
nor U16907 (N_16907,N_13151,N_13420);
nor U16908 (N_16908,N_14429,N_14802);
and U16909 (N_16909,N_14120,N_14128);
xor U16910 (N_16910,N_14262,N_13563);
and U16911 (N_16911,N_14000,N_14400);
nand U16912 (N_16912,N_13695,N_12848);
nor U16913 (N_16913,N_12884,N_14260);
xnor U16914 (N_16914,N_12825,N_13248);
nor U16915 (N_16915,N_12665,N_12778);
or U16916 (N_16916,N_14559,N_12701);
nand U16917 (N_16917,N_14661,N_12717);
and U16918 (N_16918,N_12742,N_12882);
xnor U16919 (N_16919,N_14176,N_14167);
xor U16920 (N_16920,N_12587,N_13780);
or U16921 (N_16921,N_14012,N_13213);
nand U16922 (N_16922,N_14388,N_12829);
nor U16923 (N_16923,N_13136,N_13015);
nand U16924 (N_16924,N_13013,N_13848);
and U16925 (N_16925,N_13664,N_12843);
nand U16926 (N_16926,N_12809,N_13725);
xnor U16927 (N_16927,N_13726,N_13337);
nor U16928 (N_16928,N_14093,N_14656);
xnor U16929 (N_16929,N_12789,N_13718);
and U16930 (N_16930,N_14277,N_14084);
xnor U16931 (N_16931,N_12633,N_13695);
nor U16932 (N_16932,N_13377,N_12926);
nand U16933 (N_16933,N_13193,N_12762);
xor U16934 (N_16934,N_14485,N_13052);
and U16935 (N_16935,N_13223,N_14406);
and U16936 (N_16936,N_13688,N_13974);
nand U16937 (N_16937,N_14098,N_14523);
or U16938 (N_16938,N_14963,N_12552);
nand U16939 (N_16939,N_14311,N_13053);
xor U16940 (N_16940,N_14294,N_14846);
nor U16941 (N_16941,N_12631,N_13318);
or U16942 (N_16942,N_12623,N_14721);
and U16943 (N_16943,N_14435,N_12995);
or U16944 (N_16944,N_13312,N_12589);
nor U16945 (N_16945,N_14222,N_13127);
nor U16946 (N_16946,N_14018,N_14364);
or U16947 (N_16947,N_12992,N_14605);
nand U16948 (N_16948,N_13771,N_13257);
nand U16949 (N_16949,N_14066,N_14430);
xnor U16950 (N_16950,N_14768,N_14294);
nand U16951 (N_16951,N_13026,N_14216);
xnor U16952 (N_16952,N_13515,N_14882);
xnor U16953 (N_16953,N_14796,N_14019);
xnor U16954 (N_16954,N_12981,N_12520);
or U16955 (N_16955,N_13305,N_14310);
and U16956 (N_16956,N_12811,N_14399);
nand U16957 (N_16957,N_14261,N_14542);
nor U16958 (N_16958,N_13279,N_13688);
nor U16959 (N_16959,N_13686,N_13284);
nand U16960 (N_16960,N_13812,N_14041);
nor U16961 (N_16961,N_14542,N_14376);
nand U16962 (N_16962,N_13506,N_13085);
nand U16963 (N_16963,N_14552,N_13259);
xor U16964 (N_16964,N_13670,N_12797);
and U16965 (N_16965,N_14052,N_13471);
nand U16966 (N_16966,N_14890,N_14526);
or U16967 (N_16967,N_14077,N_14130);
and U16968 (N_16968,N_13982,N_12624);
or U16969 (N_16969,N_13254,N_13379);
or U16970 (N_16970,N_14771,N_12694);
nor U16971 (N_16971,N_14121,N_14625);
xor U16972 (N_16972,N_13897,N_13501);
and U16973 (N_16973,N_14555,N_14653);
and U16974 (N_16974,N_14803,N_12726);
or U16975 (N_16975,N_13707,N_14509);
and U16976 (N_16976,N_13271,N_13821);
nand U16977 (N_16977,N_13355,N_12714);
or U16978 (N_16978,N_12614,N_14926);
xor U16979 (N_16979,N_13507,N_13082);
xor U16980 (N_16980,N_12985,N_13934);
nor U16981 (N_16981,N_13627,N_14042);
nand U16982 (N_16982,N_14983,N_14626);
or U16983 (N_16983,N_12975,N_13843);
and U16984 (N_16984,N_13631,N_14125);
nor U16985 (N_16985,N_13289,N_13968);
xor U16986 (N_16986,N_14756,N_12810);
nand U16987 (N_16987,N_13549,N_14368);
nor U16988 (N_16988,N_12796,N_13489);
nor U16989 (N_16989,N_14408,N_13319);
xor U16990 (N_16990,N_12968,N_13420);
or U16991 (N_16991,N_14351,N_14309);
nor U16992 (N_16992,N_13777,N_14912);
or U16993 (N_16993,N_12581,N_13651);
and U16994 (N_16994,N_13683,N_12898);
nor U16995 (N_16995,N_12876,N_13624);
nor U16996 (N_16996,N_13303,N_14642);
xnor U16997 (N_16997,N_13711,N_13135);
and U16998 (N_16998,N_14400,N_12648);
xor U16999 (N_16999,N_12654,N_14675);
nor U17000 (N_17000,N_13770,N_13236);
or U17001 (N_17001,N_13905,N_12689);
xor U17002 (N_17002,N_14276,N_13070);
xnor U17003 (N_17003,N_14478,N_12863);
and U17004 (N_17004,N_13429,N_14557);
or U17005 (N_17005,N_13252,N_14129);
xnor U17006 (N_17006,N_14909,N_13771);
xnor U17007 (N_17007,N_13083,N_14797);
nand U17008 (N_17008,N_12905,N_14261);
nand U17009 (N_17009,N_14037,N_14098);
and U17010 (N_17010,N_13379,N_12540);
and U17011 (N_17011,N_14687,N_12837);
and U17012 (N_17012,N_12745,N_14395);
nor U17013 (N_17013,N_13510,N_13353);
nand U17014 (N_17014,N_13097,N_12685);
xor U17015 (N_17015,N_13593,N_13307);
or U17016 (N_17016,N_14056,N_14630);
or U17017 (N_17017,N_13918,N_14660);
xor U17018 (N_17018,N_13126,N_14214);
nor U17019 (N_17019,N_13977,N_14037);
or U17020 (N_17020,N_12989,N_13018);
or U17021 (N_17021,N_12845,N_13643);
xnor U17022 (N_17022,N_13797,N_14500);
or U17023 (N_17023,N_12745,N_14322);
and U17024 (N_17024,N_13959,N_13615);
xor U17025 (N_17025,N_12926,N_14741);
xnor U17026 (N_17026,N_13979,N_12888);
and U17027 (N_17027,N_14449,N_13963);
and U17028 (N_17028,N_14286,N_14179);
xnor U17029 (N_17029,N_14476,N_13636);
and U17030 (N_17030,N_13363,N_14624);
nand U17031 (N_17031,N_12609,N_12804);
or U17032 (N_17032,N_12992,N_14898);
and U17033 (N_17033,N_14972,N_14412);
or U17034 (N_17034,N_14623,N_14532);
xor U17035 (N_17035,N_13137,N_12514);
xor U17036 (N_17036,N_12817,N_12873);
nand U17037 (N_17037,N_13886,N_13043);
xor U17038 (N_17038,N_14533,N_14303);
and U17039 (N_17039,N_12579,N_13218);
nor U17040 (N_17040,N_13156,N_13161);
xor U17041 (N_17041,N_12651,N_14179);
or U17042 (N_17042,N_14205,N_14829);
or U17043 (N_17043,N_12557,N_12937);
xor U17044 (N_17044,N_14288,N_14921);
and U17045 (N_17045,N_13626,N_12976);
xor U17046 (N_17046,N_13599,N_13794);
nor U17047 (N_17047,N_12747,N_14591);
and U17048 (N_17048,N_14222,N_13717);
nor U17049 (N_17049,N_14111,N_13543);
nor U17050 (N_17050,N_14252,N_12923);
and U17051 (N_17051,N_13030,N_12793);
xnor U17052 (N_17052,N_12888,N_14852);
nand U17053 (N_17053,N_14935,N_13977);
and U17054 (N_17054,N_14309,N_13777);
nor U17055 (N_17055,N_14681,N_12849);
and U17056 (N_17056,N_12512,N_13507);
nor U17057 (N_17057,N_12647,N_14908);
and U17058 (N_17058,N_14289,N_13573);
nor U17059 (N_17059,N_13681,N_14893);
and U17060 (N_17060,N_14886,N_14577);
nand U17061 (N_17061,N_14706,N_14004);
or U17062 (N_17062,N_13226,N_12916);
nand U17063 (N_17063,N_13287,N_12803);
nand U17064 (N_17064,N_12770,N_13142);
and U17065 (N_17065,N_14303,N_13236);
or U17066 (N_17066,N_14916,N_14350);
xor U17067 (N_17067,N_13357,N_12509);
or U17068 (N_17068,N_13831,N_14673);
or U17069 (N_17069,N_14518,N_13111);
and U17070 (N_17070,N_13982,N_14800);
nand U17071 (N_17071,N_13928,N_12578);
and U17072 (N_17072,N_13868,N_13933);
nor U17073 (N_17073,N_14120,N_14584);
and U17074 (N_17074,N_12612,N_14242);
xnor U17075 (N_17075,N_14256,N_13589);
and U17076 (N_17076,N_12966,N_13793);
or U17077 (N_17077,N_13152,N_12548);
or U17078 (N_17078,N_13435,N_12944);
nand U17079 (N_17079,N_13854,N_13436);
nor U17080 (N_17080,N_13572,N_14695);
xor U17081 (N_17081,N_14504,N_13065);
nor U17082 (N_17082,N_12523,N_13542);
and U17083 (N_17083,N_13631,N_14958);
xor U17084 (N_17084,N_13180,N_14824);
nor U17085 (N_17085,N_14805,N_14659);
or U17086 (N_17086,N_12742,N_12703);
nor U17087 (N_17087,N_13315,N_13867);
nor U17088 (N_17088,N_14482,N_14319);
nand U17089 (N_17089,N_12857,N_13978);
nor U17090 (N_17090,N_14340,N_13863);
nand U17091 (N_17091,N_14776,N_12558);
and U17092 (N_17092,N_12836,N_14782);
and U17093 (N_17093,N_13023,N_12687);
xnor U17094 (N_17094,N_13324,N_14472);
nand U17095 (N_17095,N_12798,N_13411);
xnor U17096 (N_17096,N_14161,N_14568);
or U17097 (N_17097,N_12990,N_14631);
xor U17098 (N_17098,N_13127,N_12747);
nor U17099 (N_17099,N_13734,N_14334);
nand U17100 (N_17100,N_13808,N_12556);
and U17101 (N_17101,N_13437,N_14588);
or U17102 (N_17102,N_13257,N_14109);
xor U17103 (N_17103,N_14419,N_13166);
xor U17104 (N_17104,N_14190,N_13916);
xor U17105 (N_17105,N_14914,N_13899);
nand U17106 (N_17106,N_14035,N_14994);
nand U17107 (N_17107,N_13035,N_13850);
nor U17108 (N_17108,N_13702,N_13874);
xor U17109 (N_17109,N_14894,N_13313);
nand U17110 (N_17110,N_13521,N_14123);
and U17111 (N_17111,N_13804,N_14851);
and U17112 (N_17112,N_14118,N_12997);
nor U17113 (N_17113,N_13642,N_12901);
nor U17114 (N_17114,N_13418,N_14725);
xnor U17115 (N_17115,N_12752,N_13013);
nor U17116 (N_17116,N_14287,N_13654);
or U17117 (N_17117,N_14381,N_13192);
or U17118 (N_17118,N_13025,N_12536);
nor U17119 (N_17119,N_14540,N_14831);
or U17120 (N_17120,N_14450,N_13193);
nor U17121 (N_17121,N_14009,N_13983);
and U17122 (N_17122,N_13678,N_14985);
and U17123 (N_17123,N_12701,N_13603);
and U17124 (N_17124,N_14491,N_14403);
xor U17125 (N_17125,N_12796,N_14844);
or U17126 (N_17126,N_13986,N_13144);
nor U17127 (N_17127,N_12745,N_13707);
nor U17128 (N_17128,N_14774,N_14325);
and U17129 (N_17129,N_14661,N_14952);
or U17130 (N_17130,N_13325,N_12562);
nor U17131 (N_17131,N_13043,N_13673);
and U17132 (N_17132,N_13059,N_14814);
nand U17133 (N_17133,N_12623,N_14746);
xnor U17134 (N_17134,N_12525,N_14806);
xnor U17135 (N_17135,N_13321,N_13560);
or U17136 (N_17136,N_14974,N_14834);
xnor U17137 (N_17137,N_14794,N_13121);
nor U17138 (N_17138,N_14465,N_13602);
or U17139 (N_17139,N_12788,N_13750);
nor U17140 (N_17140,N_14570,N_13032);
and U17141 (N_17141,N_13650,N_13509);
or U17142 (N_17142,N_12558,N_13547);
xor U17143 (N_17143,N_12958,N_13481);
xnor U17144 (N_17144,N_14848,N_14197);
or U17145 (N_17145,N_14271,N_12801);
and U17146 (N_17146,N_13462,N_14496);
xnor U17147 (N_17147,N_13026,N_12644);
xor U17148 (N_17148,N_14358,N_13403);
or U17149 (N_17149,N_13871,N_13895);
or U17150 (N_17150,N_13532,N_13053);
and U17151 (N_17151,N_14512,N_12962);
nor U17152 (N_17152,N_14402,N_14581);
and U17153 (N_17153,N_14013,N_13077);
nor U17154 (N_17154,N_13855,N_13500);
and U17155 (N_17155,N_14179,N_14851);
xnor U17156 (N_17156,N_14678,N_12805);
and U17157 (N_17157,N_14929,N_13219);
xor U17158 (N_17158,N_13526,N_13541);
nor U17159 (N_17159,N_13844,N_13581);
or U17160 (N_17160,N_14577,N_13882);
or U17161 (N_17161,N_14528,N_13217);
nor U17162 (N_17162,N_14466,N_13258);
nand U17163 (N_17163,N_13424,N_12700);
nand U17164 (N_17164,N_13558,N_13278);
or U17165 (N_17165,N_13727,N_14420);
and U17166 (N_17166,N_12596,N_14952);
nand U17167 (N_17167,N_13649,N_12574);
and U17168 (N_17168,N_14587,N_14284);
nor U17169 (N_17169,N_14779,N_12983);
nor U17170 (N_17170,N_13585,N_12955);
and U17171 (N_17171,N_13710,N_12928);
nor U17172 (N_17172,N_13946,N_14214);
and U17173 (N_17173,N_13547,N_14497);
xnor U17174 (N_17174,N_13238,N_13946);
or U17175 (N_17175,N_13277,N_14957);
or U17176 (N_17176,N_14161,N_12651);
and U17177 (N_17177,N_12517,N_14272);
and U17178 (N_17178,N_12519,N_14637);
xnor U17179 (N_17179,N_14866,N_14036);
nor U17180 (N_17180,N_14596,N_12831);
or U17181 (N_17181,N_13005,N_14643);
and U17182 (N_17182,N_14597,N_13815);
nand U17183 (N_17183,N_13352,N_13345);
and U17184 (N_17184,N_14857,N_12983);
and U17185 (N_17185,N_13614,N_13322);
and U17186 (N_17186,N_12740,N_14468);
xor U17187 (N_17187,N_12564,N_13809);
or U17188 (N_17188,N_13574,N_14344);
nand U17189 (N_17189,N_14171,N_13727);
xnor U17190 (N_17190,N_12904,N_13121);
nor U17191 (N_17191,N_13126,N_14728);
nor U17192 (N_17192,N_13582,N_12638);
and U17193 (N_17193,N_14875,N_14257);
or U17194 (N_17194,N_13898,N_13780);
nand U17195 (N_17195,N_12785,N_14518);
or U17196 (N_17196,N_14042,N_13483);
nor U17197 (N_17197,N_14237,N_14285);
nor U17198 (N_17198,N_12720,N_13154);
and U17199 (N_17199,N_12769,N_14518);
xnor U17200 (N_17200,N_14854,N_14435);
nand U17201 (N_17201,N_13914,N_12947);
or U17202 (N_17202,N_14902,N_13306);
nand U17203 (N_17203,N_14430,N_12763);
and U17204 (N_17204,N_14619,N_14716);
nor U17205 (N_17205,N_12862,N_12703);
nor U17206 (N_17206,N_14326,N_14661);
nor U17207 (N_17207,N_14467,N_12689);
xnor U17208 (N_17208,N_14858,N_13492);
and U17209 (N_17209,N_13337,N_14102);
or U17210 (N_17210,N_14365,N_14206);
xor U17211 (N_17211,N_13451,N_13177);
xor U17212 (N_17212,N_14287,N_13789);
or U17213 (N_17213,N_14922,N_14663);
nand U17214 (N_17214,N_14591,N_14095);
nand U17215 (N_17215,N_13488,N_14109);
and U17216 (N_17216,N_14557,N_13506);
nand U17217 (N_17217,N_14602,N_14432);
xor U17218 (N_17218,N_12874,N_14886);
nand U17219 (N_17219,N_12783,N_14348);
and U17220 (N_17220,N_14172,N_12773);
xor U17221 (N_17221,N_13996,N_14083);
nand U17222 (N_17222,N_13488,N_12509);
or U17223 (N_17223,N_14645,N_12534);
nor U17224 (N_17224,N_12640,N_13301);
nor U17225 (N_17225,N_14426,N_13747);
nor U17226 (N_17226,N_13290,N_12606);
and U17227 (N_17227,N_13876,N_14248);
nand U17228 (N_17228,N_14402,N_14962);
and U17229 (N_17229,N_14501,N_13817);
nor U17230 (N_17230,N_13793,N_14032);
nor U17231 (N_17231,N_13806,N_14815);
nand U17232 (N_17232,N_13360,N_14095);
nand U17233 (N_17233,N_14321,N_14819);
nand U17234 (N_17234,N_13105,N_12889);
and U17235 (N_17235,N_12580,N_14405);
and U17236 (N_17236,N_13170,N_12638);
or U17237 (N_17237,N_12866,N_13766);
and U17238 (N_17238,N_14722,N_14659);
or U17239 (N_17239,N_12823,N_12766);
and U17240 (N_17240,N_14914,N_14698);
xor U17241 (N_17241,N_12582,N_12562);
nand U17242 (N_17242,N_14277,N_14650);
xnor U17243 (N_17243,N_12875,N_14995);
or U17244 (N_17244,N_12873,N_14619);
nand U17245 (N_17245,N_13319,N_12657);
nand U17246 (N_17246,N_14040,N_13420);
nor U17247 (N_17247,N_12550,N_14391);
or U17248 (N_17248,N_14001,N_13631);
and U17249 (N_17249,N_13247,N_12631);
or U17250 (N_17250,N_13518,N_14119);
nand U17251 (N_17251,N_14187,N_12898);
nor U17252 (N_17252,N_13434,N_13983);
or U17253 (N_17253,N_14180,N_14225);
or U17254 (N_17254,N_13666,N_14880);
xnor U17255 (N_17255,N_13528,N_13366);
nor U17256 (N_17256,N_14430,N_13575);
and U17257 (N_17257,N_12768,N_13946);
or U17258 (N_17258,N_13651,N_13029);
xor U17259 (N_17259,N_12505,N_14462);
and U17260 (N_17260,N_13452,N_13557);
and U17261 (N_17261,N_14660,N_14419);
nand U17262 (N_17262,N_12501,N_14777);
or U17263 (N_17263,N_14068,N_14740);
or U17264 (N_17264,N_12979,N_13987);
and U17265 (N_17265,N_14680,N_13201);
nor U17266 (N_17266,N_12666,N_13564);
xor U17267 (N_17267,N_13278,N_12780);
or U17268 (N_17268,N_14873,N_12795);
or U17269 (N_17269,N_13973,N_14988);
and U17270 (N_17270,N_13649,N_14559);
nor U17271 (N_17271,N_13561,N_13894);
or U17272 (N_17272,N_14566,N_12691);
nor U17273 (N_17273,N_13694,N_14876);
or U17274 (N_17274,N_14515,N_12722);
or U17275 (N_17275,N_12579,N_13831);
or U17276 (N_17276,N_12784,N_12566);
nand U17277 (N_17277,N_13362,N_13211);
xor U17278 (N_17278,N_13445,N_14656);
nor U17279 (N_17279,N_14368,N_12811);
and U17280 (N_17280,N_12961,N_14973);
or U17281 (N_17281,N_14787,N_12914);
or U17282 (N_17282,N_14111,N_13931);
xor U17283 (N_17283,N_13779,N_12922);
and U17284 (N_17284,N_12986,N_12818);
nor U17285 (N_17285,N_14016,N_14832);
nor U17286 (N_17286,N_12659,N_14979);
xnor U17287 (N_17287,N_13700,N_14368);
and U17288 (N_17288,N_13684,N_13036);
or U17289 (N_17289,N_13480,N_14057);
and U17290 (N_17290,N_13883,N_12974);
nand U17291 (N_17291,N_14977,N_13672);
xnor U17292 (N_17292,N_13702,N_13535);
nor U17293 (N_17293,N_12599,N_13024);
nor U17294 (N_17294,N_13035,N_13083);
or U17295 (N_17295,N_13111,N_14039);
and U17296 (N_17296,N_13744,N_14166);
and U17297 (N_17297,N_13299,N_13382);
and U17298 (N_17298,N_14112,N_13597);
or U17299 (N_17299,N_13618,N_13328);
nand U17300 (N_17300,N_12618,N_13048);
xnor U17301 (N_17301,N_13644,N_13120);
and U17302 (N_17302,N_14974,N_13479);
xnor U17303 (N_17303,N_13290,N_13046);
nor U17304 (N_17304,N_13295,N_12628);
nand U17305 (N_17305,N_14751,N_12610);
nor U17306 (N_17306,N_13976,N_14596);
nand U17307 (N_17307,N_14874,N_14212);
and U17308 (N_17308,N_13558,N_13343);
and U17309 (N_17309,N_14387,N_13106);
nand U17310 (N_17310,N_13126,N_14882);
nor U17311 (N_17311,N_12569,N_13879);
nor U17312 (N_17312,N_14986,N_12564);
xor U17313 (N_17313,N_14775,N_12894);
and U17314 (N_17314,N_13709,N_12600);
and U17315 (N_17315,N_14411,N_14005);
xnor U17316 (N_17316,N_14740,N_13163);
and U17317 (N_17317,N_14898,N_14874);
xor U17318 (N_17318,N_14979,N_13931);
and U17319 (N_17319,N_14162,N_12963);
xor U17320 (N_17320,N_13151,N_14167);
nand U17321 (N_17321,N_12527,N_14060);
or U17322 (N_17322,N_14605,N_14204);
nor U17323 (N_17323,N_12548,N_13104);
and U17324 (N_17324,N_13621,N_12890);
nor U17325 (N_17325,N_14912,N_12712);
nor U17326 (N_17326,N_14530,N_12694);
nor U17327 (N_17327,N_13073,N_13037);
and U17328 (N_17328,N_14106,N_14965);
or U17329 (N_17329,N_13610,N_12699);
xnor U17330 (N_17330,N_14063,N_14770);
xor U17331 (N_17331,N_14050,N_14553);
nand U17332 (N_17332,N_13704,N_13967);
xnor U17333 (N_17333,N_13830,N_14945);
xnor U17334 (N_17334,N_14007,N_14541);
nor U17335 (N_17335,N_13679,N_13636);
and U17336 (N_17336,N_12928,N_12765);
xor U17337 (N_17337,N_13844,N_12562);
or U17338 (N_17338,N_13281,N_13176);
nand U17339 (N_17339,N_13020,N_13100);
nand U17340 (N_17340,N_12571,N_13022);
and U17341 (N_17341,N_13815,N_14925);
or U17342 (N_17342,N_14300,N_14952);
nand U17343 (N_17343,N_13239,N_13433);
nor U17344 (N_17344,N_13653,N_12663);
xor U17345 (N_17345,N_13405,N_14593);
or U17346 (N_17346,N_12579,N_14801);
nand U17347 (N_17347,N_13330,N_14354);
xnor U17348 (N_17348,N_14380,N_12737);
nor U17349 (N_17349,N_12949,N_13556);
or U17350 (N_17350,N_14867,N_14175);
nand U17351 (N_17351,N_13058,N_12851);
nand U17352 (N_17352,N_13785,N_14093);
nor U17353 (N_17353,N_13403,N_12750);
nor U17354 (N_17354,N_13014,N_13381);
or U17355 (N_17355,N_14733,N_12783);
nand U17356 (N_17356,N_14524,N_12526);
xnor U17357 (N_17357,N_13670,N_13284);
nor U17358 (N_17358,N_13979,N_14079);
xnor U17359 (N_17359,N_13833,N_13979);
and U17360 (N_17360,N_14616,N_13335);
or U17361 (N_17361,N_13223,N_12514);
nor U17362 (N_17362,N_14010,N_14839);
or U17363 (N_17363,N_13395,N_12814);
or U17364 (N_17364,N_14638,N_13164);
and U17365 (N_17365,N_13792,N_13830);
xor U17366 (N_17366,N_13084,N_13088);
and U17367 (N_17367,N_12843,N_13873);
xor U17368 (N_17368,N_14246,N_13663);
and U17369 (N_17369,N_13687,N_13645);
nand U17370 (N_17370,N_12930,N_13109);
nand U17371 (N_17371,N_14816,N_14347);
xnor U17372 (N_17372,N_13601,N_14593);
nor U17373 (N_17373,N_13328,N_13246);
or U17374 (N_17374,N_12724,N_12964);
nand U17375 (N_17375,N_14823,N_12981);
xnor U17376 (N_17376,N_13029,N_13972);
xor U17377 (N_17377,N_13993,N_12694);
nand U17378 (N_17378,N_14254,N_13798);
and U17379 (N_17379,N_14488,N_12810);
or U17380 (N_17380,N_14773,N_13440);
xor U17381 (N_17381,N_13353,N_13955);
xnor U17382 (N_17382,N_14597,N_13162);
or U17383 (N_17383,N_14820,N_12786);
nand U17384 (N_17384,N_14253,N_14589);
nand U17385 (N_17385,N_12876,N_12855);
nor U17386 (N_17386,N_12861,N_12770);
xor U17387 (N_17387,N_13612,N_14854);
nor U17388 (N_17388,N_13680,N_14847);
xnor U17389 (N_17389,N_14985,N_13459);
nand U17390 (N_17390,N_14713,N_13225);
nand U17391 (N_17391,N_13330,N_14865);
nor U17392 (N_17392,N_12539,N_13480);
nand U17393 (N_17393,N_14157,N_13219);
and U17394 (N_17394,N_12956,N_14119);
nand U17395 (N_17395,N_13315,N_14655);
or U17396 (N_17396,N_13420,N_13504);
nor U17397 (N_17397,N_14734,N_14668);
or U17398 (N_17398,N_14670,N_14684);
xnor U17399 (N_17399,N_14675,N_12771);
xnor U17400 (N_17400,N_13549,N_13539);
and U17401 (N_17401,N_12922,N_14391);
nand U17402 (N_17402,N_13896,N_14243);
nor U17403 (N_17403,N_13536,N_13187);
and U17404 (N_17404,N_12681,N_13735);
nor U17405 (N_17405,N_14303,N_12799);
xor U17406 (N_17406,N_13951,N_14703);
nand U17407 (N_17407,N_12676,N_13542);
or U17408 (N_17408,N_14620,N_13595);
xnor U17409 (N_17409,N_13977,N_14643);
xnor U17410 (N_17410,N_13998,N_13083);
and U17411 (N_17411,N_12678,N_13347);
or U17412 (N_17412,N_13339,N_14193);
nand U17413 (N_17413,N_14897,N_14177);
or U17414 (N_17414,N_13097,N_12923);
nand U17415 (N_17415,N_13026,N_14032);
xor U17416 (N_17416,N_12901,N_13409);
nand U17417 (N_17417,N_12976,N_13231);
xor U17418 (N_17418,N_14182,N_12557);
nand U17419 (N_17419,N_12622,N_13158);
or U17420 (N_17420,N_14649,N_14927);
or U17421 (N_17421,N_12917,N_13153);
or U17422 (N_17422,N_14638,N_13987);
and U17423 (N_17423,N_13190,N_14121);
xor U17424 (N_17424,N_13747,N_14994);
nand U17425 (N_17425,N_12650,N_13409);
nand U17426 (N_17426,N_14446,N_14322);
or U17427 (N_17427,N_13894,N_13806);
nand U17428 (N_17428,N_12507,N_13267);
nor U17429 (N_17429,N_14259,N_13984);
or U17430 (N_17430,N_14997,N_14861);
xnor U17431 (N_17431,N_14057,N_14453);
xnor U17432 (N_17432,N_13672,N_12579);
nand U17433 (N_17433,N_14319,N_13093);
and U17434 (N_17434,N_13581,N_12750);
nand U17435 (N_17435,N_13977,N_14668);
nor U17436 (N_17436,N_12959,N_13764);
xnor U17437 (N_17437,N_14077,N_14619);
nor U17438 (N_17438,N_14943,N_14083);
nor U17439 (N_17439,N_12694,N_13009);
xnor U17440 (N_17440,N_13116,N_12874);
nor U17441 (N_17441,N_12903,N_13635);
nand U17442 (N_17442,N_13536,N_12812);
nor U17443 (N_17443,N_13644,N_12635);
and U17444 (N_17444,N_14839,N_14896);
or U17445 (N_17445,N_14082,N_13438);
or U17446 (N_17446,N_14281,N_13510);
nor U17447 (N_17447,N_12812,N_14074);
and U17448 (N_17448,N_13931,N_14154);
nor U17449 (N_17449,N_14157,N_14668);
nand U17450 (N_17450,N_12707,N_13887);
nand U17451 (N_17451,N_14062,N_14852);
nand U17452 (N_17452,N_14773,N_13178);
xor U17453 (N_17453,N_13085,N_12900);
xor U17454 (N_17454,N_13544,N_14113);
nand U17455 (N_17455,N_14629,N_13875);
or U17456 (N_17456,N_14699,N_14520);
nor U17457 (N_17457,N_14302,N_14280);
or U17458 (N_17458,N_13522,N_13993);
and U17459 (N_17459,N_13997,N_13404);
or U17460 (N_17460,N_13080,N_13091);
and U17461 (N_17461,N_12685,N_13154);
and U17462 (N_17462,N_14977,N_13889);
nand U17463 (N_17463,N_13130,N_14673);
xor U17464 (N_17464,N_12938,N_13099);
or U17465 (N_17465,N_13027,N_13679);
nor U17466 (N_17466,N_12534,N_13703);
nand U17467 (N_17467,N_14241,N_12786);
or U17468 (N_17468,N_14886,N_13945);
nor U17469 (N_17469,N_12728,N_12710);
and U17470 (N_17470,N_14692,N_13775);
nand U17471 (N_17471,N_14805,N_13098);
or U17472 (N_17472,N_13854,N_14558);
or U17473 (N_17473,N_12914,N_13790);
xnor U17474 (N_17474,N_13547,N_14709);
nand U17475 (N_17475,N_14435,N_14525);
nor U17476 (N_17476,N_14116,N_14937);
nand U17477 (N_17477,N_12794,N_12666);
xnor U17478 (N_17478,N_12853,N_14026);
and U17479 (N_17479,N_14136,N_13889);
xor U17480 (N_17480,N_14419,N_12662);
nor U17481 (N_17481,N_13779,N_13576);
nand U17482 (N_17482,N_13621,N_12563);
nand U17483 (N_17483,N_12576,N_12716);
nor U17484 (N_17484,N_13063,N_14870);
nand U17485 (N_17485,N_14677,N_14115);
nand U17486 (N_17486,N_14147,N_14274);
xnor U17487 (N_17487,N_13114,N_13728);
nand U17488 (N_17488,N_13307,N_12925);
xnor U17489 (N_17489,N_12621,N_13822);
nor U17490 (N_17490,N_14735,N_14827);
nor U17491 (N_17491,N_13217,N_13573);
nand U17492 (N_17492,N_14977,N_12990);
xnor U17493 (N_17493,N_14090,N_14676);
nand U17494 (N_17494,N_13172,N_14289);
nand U17495 (N_17495,N_14929,N_13768);
xor U17496 (N_17496,N_13226,N_14323);
or U17497 (N_17497,N_12794,N_13265);
and U17498 (N_17498,N_14812,N_12999);
nor U17499 (N_17499,N_12654,N_14878);
or U17500 (N_17500,N_15965,N_15120);
nor U17501 (N_17501,N_16053,N_16860);
xor U17502 (N_17502,N_17357,N_16259);
or U17503 (N_17503,N_16244,N_16348);
xor U17504 (N_17504,N_15998,N_16703);
and U17505 (N_17505,N_16377,N_15489);
nand U17506 (N_17506,N_15181,N_15964);
nor U17507 (N_17507,N_15567,N_15338);
or U17508 (N_17508,N_17034,N_15179);
nor U17509 (N_17509,N_15246,N_16935);
xor U17510 (N_17510,N_15766,N_15696);
or U17511 (N_17511,N_17386,N_16832);
xnor U17512 (N_17512,N_16503,N_15382);
xor U17513 (N_17513,N_15924,N_16679);
or U17514 (N_17514,N_15054,N_16313);
nor U17515 (N_17515,N_16496,N_15042);
nand U17516 (N_17516,N_16559,N_16073);
nor U17517 (N_17517,N_16554,N_15647);
xor U17518 (N_17518,N_16278,N_15517);
nand U17519 (N_17519,N_15968,N_15421);
nor U17520 (N_17520,N_16697,N_16119);
xnor U17521 (N_17521,N_17311,N_17331);
and U17522 (N_17522,N_15084,N_15570);
and U17523 (N_17523,N_17318,N_17250);
or U17524 (N_17524,N_16965,N_16153);
or U17525 (N_17525,N_17160,N_16523);
nand U17526 (N_17526,N_16071,N_16729);
and U17527 (N_17527,N_16213,N_15746);
nand U17528 (N_17528,N_17452,N_15863);
nand U17529 (N_17529,N_15367,N_15869);
xor U17530 (N_17530,N_16366,N_15558);
or U17531 (N_17531,N_17280,N_16945);
and U17532 (N_17532,N_16401,N_16558);
or U17533 (N_17533,N_16604,N_15698);
or U17534 (N_17534,N_17399,N_16130);
xnor U17535 (N_17535,N_17110,N_16795);
nor U17536 (N_17536,N_17328,N_17231);
xnor U17537 (N_17537,N_17142,N_15827);
xor U17538 (N_17538,N_16685,N_16952);
or U17539 (N_17539,N_16910,N_16658);
nor U17540 (N_17540,N_15520,N_15473);
xnor U17541 (N_17541,N_15554,N_16369);
xor U17542 (N_17542,N_15920,N_17052);
xor U17543 (N_17543,N_17249,N_17405);
xnor U17544 (N_17544,N_16903,N_15887);
nor U17545 (N_17545,N_15342,N_15436);
nor U17546 (N_17546,N_15643,N_17068);
nand U17547 (N_17547,N_16004,N_16502);
xnor U17548 (N_17548,N_15224,N_16957);
and U17549 (N_17549,N_15127,N_15066);
and U17550 (N_17550,N_16694,N_15569);
and U17551 (N_17551,N_15144,N_15034);
and U17552 (N_17552,N_16270,N_16659);
or U17553 (N_17553,N_15991,N_17055);
and U17554 (N_17554,N_17212,N_15079);
nor U17555 (N_17555,N_15892,N_17494);
nor U17556 (N_17556,N_16819,N_17143);
nor U17557 (N_17557,N_15493,N_15539);
or U17558 (N_17558,N_15491,N_15404);
nor U17559 (N_17559,N_16243,N_16564);
or U17560 (N_17560,N_16762,N_17097);
and U17561 (N_17561,N_16676,N_16322);
nand U17562 (N_17562,N_15700,N_15780);
nor U17563 (N_17563,N_17333,N_16985);
nor U17564 (N_17564,N_15156,N_15061);
nor U17565 (N_17565,N_16672,N_16532);
nand U17566 (N_17566,N_15791,N_17077);
and U17567 (N_17567,N_16192,N_15363);
nor U17568 (N_17568,N_16804,N_15538);
nor U17569 (N_17569,N_15242,N_17471);
nor U17570 (N_17570,N_17429,N_16383);
and U17571 (N_17571,N_16831,N_15312);
and U17572 (N_17572,N_17257,N_17123);
nor U17573 (N_17573,N_15065,N_15919);
nor U17574 (N_17574,N_16520,N_15056);
and U17575 (N_17575,N_15727,N_17381);
xor U17576 (N_17576,N_16177,N_17245);
or U17577 (N_17577,N_16370,N_16929);
or U17578 (N_17578,N_16590,N_16197);
nand U17579 (N_17579,N_15632,N_16483);
nor U17580 (N_17580,N_15479,N_16481);
or U17581 (N_17581,N_16498,N_15143);
or U17582 (N_17582,N_15463,N_16253);
and U17583 (N_17583,N_17465,N_17206);
nand U17584 (N_17584,N_17324,N_15197);
nand U17585 (N_17585,N_16067,N_15110);
and U17586 (N_17586,N_15255,N_15376);
nor U17587 (N_17587,N_16393,N_17168);
or U17588 (N_17588,N_17009,N_15490);
and U17589 (N_17589,N_17427,N_16859);
and U17590 (N_17590,N_16199,N_17102);
or U17591 (N_17591,N_16912,N_17173);
nor U17592 (N_17592,N_17347,N_15831);
nor U17593 (N_17593,N_16678,N_17223);
nand U17594 (N_17594,N_16200,N_16951);
xnor U17595 (N_17595,N_15899,N_17027);
or U17596 (N_17596,N_17379,N_17462);
nor U17597 (N_17597,N_16711,N_15770);
and U17598 (N_17598,N_15228,N_16389);
and U17599 (N_17599,N_16332,N_16204);
nand U17600 (N_17600,N_15748,N_15315);
or U17601 (N_17601,N_16886,N_15214);
nand U17602 (N_17602,N_15756,N_17035);
xnor U17603 (N_17603,N_15853,N_16136);
nor U17604 (N_17604,N_15534,N_17273);
and U17605 (N_17605,N_15828,N_17109);
xnor U17606 (N_17606,N_16104,N_15243);
nor U17607 (N_17607,N_15150,N_15693);
xnor U17608 (N_17608,N_15523,N_15196);
nand U17609 (N_17609,N_15321,N_16514);
nor U17610 (N_17610,N_15716,N_16344);
nor U17611 (N_17611,N_16091,N_15714);
or U17612 (N_17612,N_15074,N_16290);
nand U17613 (N_17613,N_15631,N_16343);
nand U17614 (N_17614,N_17221,N_15271);
nor U17615 (N_17615,N_16317,N_16544);
xnor U17616 (N_17616,N_16636,N_15916);
nand U17617 (N_17617,N_17135,N_15102);
and U17618 (N_17618,N_16986,N_16328);
xor U17619 (N_17619,N_15680,N_15986);
xor U17620 (N_17620,N_15636,N_15131);
and U17621 (N_17621,N_16407,N_15139);
xnor U17622 (N_17622,N_16072,N_17489);
or U17623 (N_17623,N_15132,N_17202);
or U17624 (N_17624,N_16125,N_15007);
xnor U17625 (N_17625,N_17140,N_15417);
nor U17626 (N_17626,N_15880,N_16684);
or U17627 (N_17627,N_16633,N_15318);
nand U17628 (N_17628,N_17370,N_16115);
xor U17629 (N_17629,N_17404,N_17434);
or U17630 (N_17630,N_17411,N_16228);
and U17631 (N_17631,N_15768,N_15108);
nor U17632 (N_17632,N_17122,N_16997);
xnor U17633 (N_17633,N_16789,N_17059);
or U17634 (N_17634,N_16166,N_16572);
and U17635 (N_17635,N_17466,N_15835);
or U17636 (N_17636,N_15453,N_15137);
and U17637 (N_17637,N_17486,N_16648);
nor U17638 (N_17638,N_15803,N_15855);
and U17639 (N_17639,N_15667,N_17442);
xor U17640 (N_17640,N_16225,N_15050);
or U17641 (N_17641,N_15515,N_17332);
nor U17642 (N_17642,N_16400,N_16628);
and U17643 (N_17643,N_16509,N_15116);
xor U17644 (N_17644,N_15531,N_15337);
nor U17645 (N_17645,N_15655,N_15948);
or U17646 (N_17646,N_17073,N_16974);
nor U17647 (N_17647,N_15682,N_15291);
or U17648 (N_17648,N_16733,N_15934);
nand U17649 (N_17649,N_16363,N_15280);
nor U17650 (N_17650,N_15870,N_16327);
nor U17651 (N_17651,N_17416,N_17453);
nor U17652 (N_17652,N_16978,N_15737);
nand U17653 (N_17653,N_15470,N_16388);
xnor U17654 (N_17654,N_15406,N_17066);
xnor U17655 (N_17655,N_15250,N_15507);
nor U17656 (N_17656,N_16022,N_15929);
or U17657 (N_17657,N_15435,N_15414);
xor U17658 (N_17658,N_17430,N_15778);
nor U17659 (N_17659,N_15506,N_17174);
nand U17660 (N_17660,N_15049,N_15537);
or U17661 (N_17661,N_15789,N_16999);
nand U17662 (N_17662,N_17480,N_16482);
nor U17663 (N_17663,N_15583,N_17190);
nand U17664 (N_17664,N_16390,N_15782);
and U17665 (N_17665,N_15472,N_16391);
nand U17666 (N_17666,N_17485,N_16459);
or U17667 (N_17667,N_16149,N_17082);
nand U17668 (N_17668,N_16062,N_16698);
nand U17669 (N_17669,N_16640,N_16222);
nand U17670 (N_17670,N_15186,N_15254);
nand U17671 (N_17671,N_15184,N_17417);
or U17672 (N_17672,N_16656,N_15294);
and U17673 (N_17673,N_15595,N_16522);
and U17674 (N_17674,N_16955,N_16298);
and U17675 (N_17675,N_17036,N_15136);
xor U17676 (N_17676,N_15957,N_17474);
nor U17677 (N_17677,N_16537,N_15518);
or U17678 (N_17678,N_16591,N_15597);
nand U17679 (N_17679,N_17226,N_16092);
nor U17680 (N_17680,N_17219,N_15457);
and U17681 (N_17681,N_16937,N_15813);
and U17682 (N_17682,N_15476,N_15985);
and U17683 (N_17683,N_16135,N_16487);
nand U17684 (N_17684,N_15174,N_17230);
or U17685 (N_17685,N_15212,N_17440);
and U17686 (N_17686,N_17112,N_15456);
xnor U17687 (N_17687,N_16036,N_16970);
and U17688 (N_17688,N_16643,N_16977);
and U17689 (N_17689,N_17421,N_16950);
or U17690 (N_17690,N_15233,N_16586);
nor U17691 (N_17691,N_16013,N_16320);
nor U17692 (N_17692,N_17234,N_15949);
or U17693 (N_17693,N_15109,N_17222);
nand U17694 (N_17694,N_15252,N_17111);
nand U17695 (N_17695,N_17336,N_15839);
nor U17696 (N_17696,N_15001,N_15510);
and U17697 (N_17697,N_17133,N_17119);
xnor U17698 (N_17698,N_17287,N_16094);
and U17699 (N_17699,N_17118,N_15475);
nor U17700 (N_17700,N_15654,N_16452);
nor U17701 (N_17701,N_17029,N_16907);
nand U17702 (N_17702,N_17389,N_15175);
xnor U17703 (N_17703,N_16661,N_15584);
xor U17704 (N_17704,N_15917,N_16737);
and U17705 (N_17705,N_17444,N_17037);
and U17706 (N_17706,N_17194,N_16829);
or U17707 (N_17707,N_15033,N_16495);
or U17708 (N_17708,N_15171,N_16041);
xor U17709 (N_17709,N_17458,N_16264);
or U17710 (N_17710,N_17121,N_15162);
nand U17711 (N_17711,N_16272,N_16506);
nor U17712 (N_17712,N_16949,N_16934);
xor U17713 (N_17713,N_16142,N_15850);
nand U17714 (N_17714,N_16218,N_16157);
and U17715 (N_17715,N_16237,N_16240);
and U17716 (N_17716,N_15977,N_16624);
nand U17717 (N_17717,N_15410,N_16567);
nand U17718 (N_17718,N_17218,N_16880);
xor U17719 (N_17719,N_15481,N_16782);
xor U17720 (N_17720,N_15692,N_16242);
nand U17721 (N_17721,N_17013,N_16916);
nor U17722 (N_17722,N_16176,N_16444);
and U17723 (N_17723,N_16494,N_17482);
and U17724 (N_17724,N_15677,N_15976);
nand U17725 (N_17725,N_15052,N_16542);
xnor U17726 (N_17726,N_15449,N_15273);
nand U17727 (N_17727,N_15101,N_15730);
and U17728 (N_17728,N_16287,N_15117);
nor U17729 (N_17729,N_15094,N_16282);
nor U17730 (N_17730,N_16175,N_15847);
and U17731 (N_17731,N_17182,N_15541);
or U17732 (N_17732,N_16754,N_16990);
nand U17733 (N_17733,N_15710,N_15563);
or U17734 (N_17734,N_17369,N_15725);
nor U17735 (N_17735,N_15704,N_16260);
xnor U17736 (N_17736,N_16038,N_16879);
xor U17737 (N_17737,N_16068,N_15209);
and U17738 (N_17738,N_17334,N_17127);
nand U17739 (N_17739,N_16919,N_15885);
and U17740 (N_17740,N_16280,N_15702);
or U17741 (N_17741,N_16475,N_17115);
nor U17742 (N_17742,N_17390,N_16601);
xnor U17743 (N_17743,N_15540,N_16141);
or U17744 (N_17744,N_15051,N_15307);
and U17745 (N_17745,N_15332,N_15459);
and U17746 (N_17746,N_16896,N_15878);
or U17747 (N_17747,N_15502,N_15607);
nand U17748 (N_17748,N_16803,N_15237);
nand U17749 (N_17749,N_16666,N_15794);
xor U17750 (N_17750,N_16023,N_16269);
xor U17751 (N_17751,N_17468,N_15422);
nor U17752 (N_17752,N_17196,N_16011);
nor U17753 (N_17753,N_16635,N_15428);
xor U17754 (N_17754,N_15275,N_15093);
and U17755 (N_17755,N_15343,N_16156);
nand U17756 (N_17756,N_17436,N_16455);
xor U17757 (N_17757,N_15225,N_16589);
nor U17758 (N_17758,N_16593,N_16606);
or U17759 (N_17759,N_16336,N_15774);
nand U17760 (N_17760,N_15441,N_15360);
or U17761 (N_17761,N_16231,N_17031);
xor U17762 (N_17762,N_15621,N_15944);
and U17763 (N_17763,N_15402,N_15818);
and U17764 (N_17764,N_17152,N_15088);
nor U17765 (N_17765,N_16417,N_15912);
and U17766 (N_17766,N_17254,N_15443);
nor U17767 (N_17767,N_15433,N_15829);
xnor U17768 (N_17768,N_15474,N_15645);
nand U17769 (N_17769,N_16644,N_15005);
nand U17770 (N_17770,N_16619,N_16405);
nand U17771 (N_17771,N_17356,N_17158);
or U17772 (N_17772,N_16602,N_16026);
or U17773 (N_17773,N_15465,N_15285);
xor U17774 (N_17774,N_15528,N_15147);
xnor U17775 (N_17775,N_15656,N_15378);
nand U17776 (N_17776,N_16054,N_15573);
xor U17777 (N_17777,N_15905,N_15266);
nand U17778 (N_17778,N_15241,N_17397);
nor U17779 (N_17779,N_15014,N_16858);
xor U17780 (N_17780,N_15339,N_16816);
and U17781 (N_17781,N_16847,N_15571);
nand U17782 (N_17782,N_15660,N_16569);
nand U17783 (N_17783,N_16761,N_16372);
or U17784 (N_17784,N_16032,N_16866);
xor U17785 (N_17785,N_16184,N_15355);
xnor U17786 (N_17786,N_15028,N_16172);
nor U17787 (N_17787,N_16430,N_16581);
nand U17788 (N_17788,N_17063,N_17006);
or U17789 (N_17789,N_16394,N_15015);
xnor U17790 (N_17790,N_17238,N_15796);
nor U17791 (N_17791,N_15030,N_16682);
xor U17792 (N_17792,N_15723,N_16534);
or U17793 (N_17793,N_15519,N_16453);
nand U17794 (N_17794,N_17293,N_15875);
nand U17795 (N_17795,N_16028,N_15936);
nor U17796 (N_17796,N_16012,N_15691);
and U17797 (N_17797,N_15729,N_16627);
nor U17798 (N_17798,N_15046,N_16812);
or U17799 (N_17799,N_15055,N_16330);
or U17800 (N_17800,N_16731,N_15872);
or U17801 (N_17801,N_16758,N_15036);
nand U17802 (N_17802,N_17358,N_16059);
and U17803 (N_17803,N_17211,N_15299);
xnor U17804 (N_17804,N_16263,N_16850);
and U17805 (N_17805,N_15302,N_17054);
xor U17806 (N_17806,N_15641,N_16660);
and U17807 (N_17807,N_16843,N_16404);
or U17808 (N_17808,N_16357,N_16655);
nand U17809 (N_17809,N_17060,N_15384);
or U17810 (N_17810,N_16851,N_15959);
nand U17811 (N_17811,N_17005,N_15599);
xnor U17812 (N_17812,N_16379,N_16232);
and U17813 (N_17813,N_16374,N_15089);
or U17814 (N_17814,N_17274,N_17235);
nand U17815 (N_17815,N_15659,N_15933);
or U17816 (N_17816,N_16205,N_17275);
nand U17817 (N_17817,N_16465,N_17237);
nand U17818 (N_17818,N_16821,N_17107);
and U17819 (N_17819,N_16550,N_15990);
nor U17820 (N_17820,N_16811,N_15446);
and U17821 (N_17821,N_17481,N_16463);
nor U17822 (N_17822,N_17377,N_15927);
and U17823 (N_17823,N_17185,N_15635);
xor U17824 (N_17824,N_15247,N_16508);
nand U17825 (N_17825,N_16342,N_16667);
nand U17826 (N_17826,N_17343,N_15845);
or U17827 (N_17827,N_16331,N_17010);
or U17828 (N_17828,N_15270,N_15129);
xor U17829 (N_17829,N_17281,N_15579);
xor U17830 (N_17830,N_16958,N_15059);
nor U17831 (N_17831,N_15035,N_16566);
and U17832 (N_17832,N_17091,N_17294);
nor U17833 (N_17833,N_17016,N_17247);
xor U17834 (N_17834,N_15889,N_15206);
or U17835 (N_17835,N_16897,N_16245);
nand U17836 (N_17836,N_17265,N_15591);
nor U17837 (N_17837,N_17108,N_15146);
and U17838 (N_17838,N_15904,N_15154);
nor U17839 (N_17839,N_17312,N_16800);
xor U17840 (N_17840,N_15153,N_16750);
nor U17841 (N_17841,N_17251,N_16705);
nor U17842 (N_17842,N_15322,N_16971);
xor U17843 (N_17843,N_17259,N_15582);
nand U17844 (N_17844,N_15619,N_15073);
nand U17845 (N_17845,N_15201,N_16474);
or U17846 (N_17846,N_16780,N_16521);
or U17847 (N_17847,N_17162,N_15278);
nor U17848 (N_17848,N_15283,N_17072);
or U17849 (N_17849,N_15119,N_15100);
nor U17850 (N_17850,N_16936,N_15555);
nand U17851 (N_17851,N_15810,N_16626);
nor U17852 (N_17852,N_15039,N_15706);
nand U17853 (N_17853,N_16296,N_15395);
and U17854 (N_17854,N_16966,N_17098);
nor U17855 (N_17855,N_15353,N_16093);
and U17856 (N_17856,N_16973,N_17058);
and U17857 (N_17857,N_17184,N_15077);
xor U17858 (N_17858,N_16064,N_17306);
and U17859 (N_17859,N_15564,N_15464);
and U17860 (N_17860,N_16285,N_16629);
nand U17861 (N_17861,N_16609,N_16798);
and U17862 (N_17862,N_17288,N_16852);
nor U17863 (N_17863,N_17243,N_16020);
nand U17864 (N_17864,N_16546,N_17422);
xor U17865 (N_17865,N_15424,N_15744);
or U17866 (N_17866,N_17391,N_16471);
nor U17867 (N_17867,N_16749,N_16333);
nor U17868 (N_17868,N_16857,N_17497);
or U17869 (N_17869,N_16930,N_16620);
and U17870 (N_17870,N_15514,N_15076);
nand U17871 (N_17871,N_15207,N_16460);
nor U17872 (N_17872,N_16841,N_15600);
nor U17873 (N_17873,N_16894,N_15525);
or U17874 (N_17874,N_17065,N_15060);
xnor U17875 (N_17875,N_16665,N_15263);
or U17876 (N_17876,N_15387,N_17020);
and U17877 (N_17877,N_15745,N_16210);
and U17878 (N_17878,N_17487,N_15265);
and U17879 (N_17879,N_16061,N_15950);
or U17880 (N_17880,N_16646,N_16443);
xor U17881 (N_17881,N_16128,N_16801);
nand U17882 (N_17882,N_16185,N_15081);
nand U17883 (N_17883,N_17423,N_16844);
nand U17884 (N_17884,N_16238,N_16726);
and U17885 (N_17885,N_15155,N_16437);
and U17886 (N_17886,N_15792,N_16909);
nor U17887 (N_17887,N_17303,N_15664);
or U17888 (N_17888,N_16148,N_15793);
xor U17889 (N_17889,N_16526,N_15350);
nor U17890 (N_17890,N_17325,N_17420);
nor U17891 (N_17891,N_15151,N_15755);
xor U17892 (N_17892,N_17137,N_16713);
nand U17893 (N_17893,N_15408,N_17090);
xor U17894 (N_17894,N_17476,N_15420);
and U17895 (N_17895,N_15652,N_15572);
or U17896 (N_17896,N_17124,N_16637);
and U17897 (N_17897,N_15053,N_17043);
nor U17898 (N_17898,N_15145,N_16615);
nor U17899 (N_17899,N_15170,N_15032);
xnor U17900 (N_17900,N_15527,N_15533);
and U17901 (N_17901,N_15697,N_16574);
and U17902 (N_17902,N_15958,N_15165);
nand U17903 (N_17903,N_16375,N_15568);
and U17904 (N_17904,N_15972,N_17075);
or U17905 (N_17905,N_16917,N_17256);
nor U17906 (N_17906,N_16358,N_16355);
xor U17907 (N_17907,N_17407,N_15366);
and U17908 (N_17908,N_15666,N_15008);
and U17909 (N_17909,N_15921,N_16868);
nand U17910 (N_17910,N_15295,N_15169);
and U17911 (N_17911,N_16385,N_16265);
nor U17912 (N_17912,N_16944,N_16884);
nor U17913 (N_17913,N_15671,N_16900);
nand U17914 (N_17914,N_17375,N_16346);
and U17915 (N_17915,N_16785,N_16337);
or U17916 (N_17916,N_17344,N_15799);
and U17917 (N_17917,N_15269,N_16410);
nor U17918 (N_17918,N_16368,N_16557);
xor U17919 (N_17919,N_16928,N_16582);
or U17920 (N_17920,N_15164,N_17359);
and U17921 (N_17921,N_16063,N_16239);
xor U17922 (N_17922,N_16740,N_16403);
xnor U17923 (N_17923,N_17236,N_16031);
nor U17924 (N_17924,N_17093,N_15394);
or U17925 (N_17925,N_16089,N_16101);
xnor U17926 (N_17926,N_15057,N_16009);
and U17927 (N_17927,N_15876,N_17302);
nand U17928 (N_17928,N_16998,N_15542);
and U17929 (N_17929,N_15626,N_15719);
and U17930 (N_17930,N_15738,N_15646);
nand U17931 (N_17931,N_17353,N_16480);
nand U17932 (N_17932,N_15906,N_16600);
and U17933 (N_17933,N_17425,N_16766);
nand U17934 (N_17934,N_16543,N_16353);
nand U17935 (N_17935,N_16439,N_16100);
xor U17936 (N_17936,N_16926,N_16014);
or U17937 (N_17937,N_17099,N_15685);
xnor U17938 (N_17938,N_15112,N_16131);
xor U17939 (N_17939,N_16826,N_17248);
or U17940 (N_17940,N_17130,N_15442);
xnor U17941 (N_17941,N_15801,N_17492);
and U17942 (N_17942,N_16623,N_15448);
nand U17943 (N_17943,N_16295,N_16641);
xor U17944 (N_17944,N_16447,N_16892);
or U17945 (N_17945,N_15765,N_16442);
and U17946 (N_17946,N_16008,N_16702);
nor U17947 (N_17947,N_16889,N_16325);
and U17948 (N_17948,N_16381,N_15258);
nand U17949 (N_17949,N_16898,N_15226);
nor U17950 (N_17950,N_16329,N_16435);
xor U17951 (N_17951,N_15838,N_17301);
xnor U17952 (N_17952,N_15996,N_17136);
xnor U17953 (N_17953,N_15858,N_16796);
or U17954 (N_17954,N_15095,N_15082);
nand U17955 (N_17955,N_16943,N_16083);
and U17956 (N_17956,N_17305,N_16836);
nor U17957 (N_17957,N_16186,N_15090);
xor U17958 (N_17958,N_16107,N_15628);
nand U17959 (N_17959,N_16735,N_17401);
or U17960 (N_17960,N_15807,N_16468);
or U17961 (N_17961,N_17050,N_16426);
or U17962 (N_17962,N_17433,N_16772);
xnor U17963 (N_17963,N_17414,N_16721);
nor U17964 (N_17964,N_15808,N_16902);
nor U17965 (N_17965,N_16939,N_15282);
nor U17966 (N_17966,N_17167,N_15460);
nand U17967 (N_17967,N_15157,N_15788);
nand U17968 (N_17968,N_16042,N_15004);
nor U17969 (N_17969,N_16145,N_16436);
or U17970 (N_17970,N_16469,N_16314);
and U17971 (N_17971,N_16645,N_16548);
nand U17972 (N_17972,N_17269,N_16476);
and U17973 (N_17973,N_16788,N_15651);
xnor U17974 (N_17974,N_17120,N_16835);
nor U17975 (N_17975,N_15287,N_16639);
xnor U17976 (N_17976,N_15763,N_15140);
xor U17977 (N_17977,N_16276,N_15290);
or U17978 (N_17978,N_17496,N_15022);
and U17979 (N_17979,N_16085,N_15707);
xnor U17980 (N_17980,N_17284,N_16075);
nor U17981 (N_17981,N_16670,N_15231);
nor U17982 (N_17982,N_15205,N_16096);
and U17983 (N_17983,N_16561,N_16473);
xnor U17984 (N_17984,N_16991,N_16201);
and U17985 (N_17985,N_16555,N_17323);
and U17986 (N_17986,N_16082,N_15982);
or U17987 (N_17987,N_15286,N_16677);
or U17988 (N_17988,N_16838,N_15178);
or U17989 (N_17989,N_17443,N_17049);
xor U17990 (N_17990,N_16163,N_16883);
nor U17991 (N_17991,N_16140,N_15951);
xnor U17992 (N_17992,N_16875,N_15758);
nand U17993 (N_17993,N_16757,N_16708);
nor U17994 (N_17994,N_15388,N_15105);
or U17995 (N_17995,N_17106,N_15375);
and U17996 (N_17996,N_16428,N_16560);
or U17997 (N_17997,N_15743,N_16499);
and U17998 (N_17998,N_16043,N_17455);
nor U17999 (N_17999,N_17080,N_16122);
and U18000 (N_18000,N_15351,N_15306);
nor U18001 (N_18001,N_16517,N_15556);
nor U18002 (N_18002,N_15264,N_15023);
and U18003 (N_18003,N_15967,N_17081);
nor U18004 (N_18004,N_17132,N_16015);
xnor U18005 (N_18005,N_16577,N_17131);
nor U18006 (N_18006,N_17141,N_16552);
nand U18007 (N_18007,N_15911,N_16599);
and U18008 (N_18008,N_17395,N_16792);
nor U18009 (N_18009,N_15213,N_16529);
or U18010 (N_18010,N_15938,N_15909);
or U18011 (N_18011,N_15027,N_15204);
nor U18012 (N_18012,N_16221,N_15326);
nand U18013 (N_18013,N_16121,N_16212);
and U18014 (N_18014,N_17400,N_16219);
xnor U18015 (N_18015,N_17337,N_15864);
or U18016 (N_18016,N_16538,N_17026);
nand U18017 (N_18017,N_15461,N_15431);
nor U18018 (N_18018,N_17169,N_16432);
xor U18019 (N_18019,N_17070,N_15425);
nand U18020 (N_18020,N_16309,N_16824);
xor U18021 (N_18021,N_15547,N_16214);
or U18022 (N_18022,N_16587,N_15328);
nand U18023 (N_18023,N_16159,N_16361);
nand U18024 (N_18024,N_15293,N_16720);
nor U18025 (N_18025,N_15199,N_15804);
xor U18026 (N_18026,N_15331,N_16732);
xor U18027 (N_18027,N_17364,N_17410);
xnor U18028 (N_18028,N_15118,N_15288);
or U18029 (N_18029,N_16638,N_15202);
and U18030 (N_18030,N_16893,N_17125);
and U18031 (N_18031,N_16268,N_17408);
and U18032 (N_18032,N_15915,N_16771);
nand U18033 (N_18033,N_15096,N_15585);
or U18034 (N_18034,N_16778,N_16825);
xnor U18035 (N_18035,N_16165,N_15592);
nor U18036 (N_18036,N_16086,N_15511);
nand U18037 (N_18037,N_17187,N_15873);
nor U18038 (N_18038,N_16467,N_15627);
xnor U18039 (N_18039,N_16256,N_16863);
or U18040 (N_18040,N_16607,N_15327);
xor U18041 (N_18041,N_15999,N_16760);
and U18042 (N_18042,N_16380,N_17022);
nor U18043 (N_18043,N_17450,N_17228);
and U18044 (N_18044,N_16161,N_15953);
nor U18045 (N_18045,N_15854,N_15423);
and U18046 (N_18046,N_16226,N_15346);
nand U18047 (N_18047,N_17084,N_15639);
xor U18048 (N_18048,N_15062,N_15913);
xor U18049 (N_18049,N_16224,N_15675);
and U18050 (N_18050,N_15069,N_16683);
nand U18051 (N_18051,N_17001,N_15415);
or U18052 (N_18052,N_16802,N_16392);
or U18053 (N_18053,N_15189,N_16914);
and U18054 (N_18054,N_15236,N_17300);
or U18055 (N_18055,N_17239,N_16029);
nand U18056 (N_18056,N_15935,N_15760);
xor U18057 (N_18057,N_17224,N_17163);
or U18058 (N_18058,N_16084,N_17104);
nor U18059 (N_18059,N_17330,N_16273);
xor U18060 (N_18060,N_16450,N_15330);
nand U18061 (N_18061,N_15396,N_16194);
nor U18062 (N_18062,N_16598,N_15529);
xor U18063 (N_18063,N_15021,N_15058);
nand U18064 (N_18064,N_17146,N_15063);
nand U18065 (N_18065,N_16006,N_15732);
and U18066 (N_18066,N_17467,N_15440);
nand U18067 (N_18067,N_15043,N_15390);
nand U18068 (N_18068,N_17350,N_16479);
nor U18069 (N_18069,N_16223,N_16252);
nor U18070 (N_18070,N_16069,N_15133);
xor U18071 (N_18071,N_16776,N_17051);
or U18072 (N_18072,N_15114,N_17024);
and U18073 (N_18073,N_17308,N_15811);
and U18074 (N_18074,N_15485,N_17021);
xor U18075 (N_18075,N_17415,N_15411);
nor U18076 (N_18076,N_16765,N_17488);
xor U18077 (N_18077,N_15006,N_16960);
and U18078 (N_18078,N_15941,N_15699);
and U18079 (N_18079,N_16323,N_15586);
xnor U18080 (N_18080,N_16236,N_16286);
nand U18081 (N_18081,N_17479,N_15663);
xnor U18082 (N_18082,N_15578,N_17004);
nor U18083 (N_18083,N_16931,N_16123);
xnor U18084 (N_18084,N_16291,N_15230);
or U18085 (N_18085,N_15978,N_16664);
xnor U18086 (N_18086,N_17057,N_15092);
xor U18087 (N_18087,N_16592,N_16845);
nor U18088 (N_18088,N_15713,N_15893);
or U18089 (N_18089,N_16608,N_17339);
or U18090 (N_18090,N_16440,N_15594);
or U18091 (N_18091,N_16745,N_16017);
and U18092 (N_18092,N_15975,N_15166);
or U18093 (N_18093,N_15445,N_15530);
and U18094 (N_18094,N_15373,N_15602);
xnor U18095 (N_18095,N_15574,N_16039);
xor U18096 (N_18096,N_15840,N_15276);
and U18097 (N_18097,N_16005,N_17172);
nand U18098 (N_18098,N_16457,N_16173);
xnor U18099 (N_18099,N_16216,N_16129);
and U18100 (N_18100,N_16284,N_16266);
xnor U18101 (N_18101,N_16220,N_15994);
nor U18102 (N_18102,N_15817,N_17366);
and U18103 (N_18103,N_16103,N_16650);
xor U18104 (N_18104,N_17313,N_17056);
and U18105 (N_18105,N_16301,N_16267);
or U18106 (N_18106,N_17017,N_15310);
nand U18107 (N_18107,N_16080,N_15879);
xor U18108 (N_18108,N_15504,N_17432);
or U18109 (N_18109,N_16775,N_17361);
nor U18110 (N_18110,N_15989,N_15256);
xor U18111 (N_18111,N_15741,N_16580);
or U18112 (N_18112,N_16445,N_16076);
or U18113 (N_18113,N_15313,N_16817);
or U18114 (N_18114,N_15781,N_17138);
nand U18115 (N_18115,N_16050,N_16170);
nand U18116 (N_18116,N_16397,N_17352);
nand U18117 (N_18117,N_16334,N_15268);
nand U18118 (N_18118,N_15695,N_16562);
or U18119 (N_18119,N_17253,N_15172);
or U18120 (N_18120,N_16887,N_16155);
nand U18121 (N_18121,N_16431,N_16490);
xor U18122 (N_18122,N_15836,N_17008);
xor U18123 (N_18123,N_17210,N_16992);
nor U18124 (N_18124,N_17451,N_15981);
nor U18125 (N_18125,N_17113,N_15610);
or U18126 (N_18126,N_15939,N_15842);
and U18127 (N_18127,N_15673,N_16657);
or U18128 (N_18128,N_15980,N_17297);
nor U18129 (N_18129,N_16037,N_16341);
nor U18130 (N_18130,N_17322,N_16595);
nand U18131 (N_18131,N_15816,N_17208);
and U18132 (N_18132,N_16980,N_16653);
nor U18133 (N_18133,N_16675,N_15825);
or U18134 (N_18134,N_16491,N_17209);
nand U18135 (N_18135,N_16102,N_16497);
or U18136 (N_18136,N_16513,N_17477);
nor U18137 (N_18137,N_16492,N_17047);
nor U18138 (N_18138,N_16202,N_16486);
nand U18139 (N_18139,N_16302,N_17438);
and U18140 (N_18140,N_15468,N_16680);
nand U18141 (N_18141,N_16150,N_17155);
or U18142 (N_18142,N_15687,N_15790);
and U18143 (N_18143,N_16500,N_16967);
nand U18144 (N_18144,N_15890,N_17382);
or U18145 (N_18145,N_15857,N_17282);
xnor U18146 (N_18146,N_16258,N_16060);
and U18147 (N_18147,N_17101,N_17351);
and U18148 (N_18148,N_17042,N_16109);
xnor U18149 (N_18149,N_15598,N_15480);
nand U18150 (N_18150,N_15708,N_15123);
nand U18151 (N_18151,N_16250,N_16585);
or U18152 (N_18152,N_16818,N_15513);
or U18153 (N_18153,N_15185,N_15688);
xor U18154 (N_18154,N_16462,N_15419);
xnor U18155 (N_18155,N_15851,N_15413);
xor U18156 (N_18156,N_15200,N_15381);
or U18157 (N_18157,N_16687,N_17412);
and U18158 (N_18158,N_15031,N_16541);
or U18159 (N_18159,N_15800,N_16617);
nand U18160 (N_18160,N_17319,N_15823);
xnor U18161 (N_18161,N_15320,N_16891);
nand U18162 (N_18162,N_17266,N_15987);
nor U18163 (N_18163,N_17149,N_16748);
and U18164 (N_18164,N_17217,N_17449);
xnor U18165 (N_18165,N_16262,N_16078);
nor U18166 (N_18166,N_15325,N_15877);
or U18167 (N_18167,N_15192,N_15926);
xnor U18168 (N_18168,N_16211,N_16551);
xnor U18169 (N_18169,N_15244,N_15483);
nand U18170 (N_18170,N_17044,N_16964);
nor U18171 (N_18171,N_17246,N_15478);
xor U18172 (N_18172,N_15173,N_17053);
and U18173 (N_18173,N_15167,N_15862);
nand U18174 (N_18174,N_16853,N_16594);
nor U18175 (N_18175,N_15674,N_17252);
nand U18176 (N_18176,N_17216,N_17156);
and U18177 (N_18177,N_15952,N_16779);
or U18178 (N_18178,N_15300,N_16618);
and U18179 (N_18179,N_16865,N_16613);
or U18180 (N_18180,N_16077,N_16402);
nor U18181 (N_18181,N_16527,N_16255);
nand U18182 (N_18182,N_17299,N_15392);
nand U18183 (N_18183,N_16099,N_15319);
nand U18184 (N_18184,N_16822,N_16915);
or U18185 (N_18185,N_15971,N_15409);
or U18186 (N_18186,N_15251,N_15724);
or U18187 (N_18187,N_15349,N_15928);
xor U18188 (N_18188,N_16485,N_15612);
xnor U18189 (N_18189,N_16367,N_16616);
nor U18190 (N_18190,N_15227,N_16168);
xnor U18191 (N_18191,N_16147,N_16905);
and U18192 (N_18192,N_16727,N_17384);
or U18193 (N_18193,N_17227,N_15078);
xor U18194 (N_18194,N_17011,N_16303);
nand U18195 (N_18195,N_15786,N_16710);
nor U18196 (N_18196,N_16398,N_15374);
and U18197 (N_18197,N_15203,N_16854);
nor U18198 (N_18198,N_15805,N_16354);
nand U18199 (N_18199,N_15305,N_16755);
and U18200 (N_18200,N_15019,N_15248);
or U18201 (N_18201,N_16519,N_16279);
and U18202 (N_18202,N_16947,N_16137);
xnor U18203 (N_18203,N_15012,N_15565);
xor U18204 (N_18204,N_16840,N_16921);
nand U18205 (N_18205,N_16052,N_16016);
xnor U18206 (N_18206,N_15486,N_17341);
and U18207 (N_18207,N_15148,N_15277);
nor U18208 (N_18208,N_17260,N_16230);
or U18209 (N_18209,N_16524,N_16806);
nand U18210 (N_18210,N_16938,N_16813);
nand U18211 (N_18211,N_15168,N_16472);
nand U18212 (N_18212,N_16274,N_17199);
xnor U18213 (N_18213,N_15107,N_17233);
and U18214 (N_18214,N_15358,N_15126);
and U18215 (N_18215,N_17262,N_15672);
or U18216 (N_18216,N_17435,N_15067);
nand U18217 (N_18217,N_16696,N_15625);
xor U18218 (N_18218,N_16422,N_16106);
and U18219 (N_18219,N_16864,N_15559);
xor U18220 (N_18220,N_15072,N_16033);
xor U18221 (N_18221,N_16895,N_16873);
nand U18222 (N_18222,N_17371,N_16198);
or U18223 (N_18223,N_15365,N_15670);
xor U18224 (N_18224,N_15177,N_15819);
and U18225 (N_18225,N_15386,N_16151);
nor U18226 (N_18226,N_17126,N_16714);
or U18227 (N_18227,N_16164,N_16764);
xor U18228 (N_18228,N_17041,N_15217);
or U18229 (N_18229,N_16057,N_17380);
or U18230 (N_18230,N_15617,N_16416);
nor U18231 (N_18231,N_15615,N_16652);
nor U18232 (N_18232,N_15946,N_17290);
nand U18233 (N_18233,N_15546,N_16419);
or U18234 (N_18234,N_17470,N_16293);
nor U18235 (N_18235,N_15357,N_15560);
or U18236 (N_18236,N_17128,N_17413);
nor U18237 (N_18237,N_17483,N_17144);
and U18238 (N_18238,N_17147,N_15340);
nand U18239 (N_18239,N_16662,N_15979);
and U18240 (N_18240,N_15642,N_16849);
or U18241 (N_18241,N_17310,N_15925);
xnor U18242 (N_18242,N_15797,N_16501);
xor U18243 (N_18243,N_17177,N_17002);
or U18244 (N_18244,N_15455,N_16908);
nor U18245 (N_18245,N_17441,N_15134);
and U18246 (N_18246,N_17493,N_17116);
nor U18247 (N_18247,N_16719,N_16742);
and U18248 (N_18248,N_15684,N_15223);
nor U18249 (N_18249,N_15566,N_17376);
xor U18250 (N_18250,N_17426,N_17258);
or U18251 (N_18251,N_16399,N_16654);
and U18252 (N_18252,N_15180,N_16339);
and U18253 (N_18253,N_17165,N_15354);
nor U18254 (N_18254,N_16261,N_17406);
and U18255 (N_18255,N_16774,N_15992);
xnor U18256 (N_18256,N_15779,N_16699);
nand U18257 (N_18257,N_17076,N_16747);
or U18258 (N_18258,N_16563,N_16738);
and U18259 (N_18259,N_15712,N_15865);
xor U18260 (N_18260,N_16768,N_15711);
or U18261 (N_18261,N_16359,N_16556);
or U18262 (N_18262,N_16979,N_15689);
or U18263 (N_18263,N_16961,N_15222);
xnor U18264 (N_18264,N_16794,N_15405);
nand U18265 (N_18265,N_16611,N_17355);
or U18266 (N_18266,N_16767,N_15097);
and U18267 (N_18267,N_15138,N_17495);
xor U18268 (N_18268,N_15304,N_16972);
and U18269 (N_18269,N_15142,N_16786);
nor U18270 (N_18270,N_15901,N_15649);
nor U18271 (N_18271,N_16540,N_17475);
or U18272 (N_18272,N_17321,N_16575);
xor U18273 (N_18273,N_16995,N_16781);
and U18274 (N_18274,N_15104,N_17204);
or U18275 (N_18275,N_17261,N_15018);
nor U18276 (N_18276,N_17114,N_15303);
nor U18277 (N_18277,N_15802,N_17030);
and U18278 (N_18278,N_15427,N_15961);
and U18279 (N_18279,N_17213,N_16746);
or U18280 (N_18280,N_16378,N_15783);
and U18281 (N_18281,N_16597,N_15398);
nand U18282 (N_18282,N_15881,N_15606);
nor U18283 (N_18283,N_16154,N_17189);
and U18284 (N_18284,N_16318,N_15947);
or U18285 (N_18285,N_16605,N_15681);
or U18286 (N_18286,N_15372,N_16427);
nor U18287 (N_18287,N_16229,N_16215);
xor U18288 (N_18288,N_15640,N_17314);
or U18289 (N_18289,N_16871,N_15942);
or U18290 (N_18290,N_17267,N_16877);
nor U18291 (N_18291,N_15798,N_15176);
and U18292 (N_18292,N_16189,N_16449);
xor U18293 (N_18293,N_16959,N_15613);
xor U18294 (N_18294,N_17148,N_15220);
or U18295 (N_18295,N_15211,N_17061);
and U18296 (N_18296,N_15362,N_15883);
or U18297 (N_18297,N_16777,N_16438);
or U18298 (N_18298,N_17183,N_15025);
nor U18299 (N_18299,N_15931,N_16456);
or U18300 (N_18300,N_15551,N_17150);
nand U18301 (N_18301,N_16044,N_15369);
nand U18302 (N_18302,N_17484,N_17373);
nand U18303 (N_18303,N_17419,N_15234);
or U18304 (N_18304,N_16420,N_16195);
nor U18305 (N_18305,N_16673,N_15393);
nand U18306 (N_18306,N_15960,N_17192);
or U18307 (N_18307,N_15832,N_15962);
nand U18308 (N_18308,N_15345,N_15902);
nor U18309 (N_18309,N_17271,N_17240);
or U18310 (N_18310,N_15454,N_15281);
nand U18311 (N_18311,N_17463,N_17186);
nand U18312 (N_18312,N_15849,N_15048);
and U18313 (N_18313,N_16307,N_17279);
xnor U18314 (N_18314,N_15494,N_17205);
xor U18315 (N_18315,N_15683,N_15040);
nor U18316 (N_18316,N_16275,N_16466);
nand U18317 (N_18317,N_17176,N_16528);
nor U18318 (N_18318,N_16413,N_16797);
nor U18319 (N_18319,N_15334,N_16759);
and U18320 (N_18320,N_17129,N_16913);
xnor U18321 (N_18321,N_16408,N_15128);
nor U18322 (N_18322,N_15198,N_16870);
and U18323 (N_18323,N_15403,N_16862);
or U18324 (N_18324,N_15484,N_17354);
nand U18325 (N_18325,N_15013,N_16872);
and U18326 (N_18326,N_15000,N_17268);
or U18327 (N_18327,N_17145,N_15160);
xnor U18328 (N_18328,N_17151,N_17229);
and U18329 (N_18329,N_17456,N_15773);
or U18330 (N_18330,N_16881,N_15407);
nand U18331 (N_18331,N_16885,N_17447);
and U18332 (N_18332,N_15762,N_16045);
and U18333 (N_18333,N_16924,N_15648);
or U18334 (N_18334,N_15581,N_17014);
nor U18335 (N_18335,N_16000,N_15333);
or U18336 (N_18336,N_17048,N_17023);
nor U18337 (N_18337,N_15826,N_15221);
nor U18338 (N_18338,N_17464,N_16396);
or U18339 (N_18339,N_15437,N_15500);
nor U18340 (N_18340,N_15561,N_15412);
or U18341 (N_18341,N_16294,N_16035);
xor U18342 (N_18342,N_16425,N_15722);
nand U18343 (N_18343,N_15603,N_15846);
nor U18344 (N_18344,N_15701,N_16288);
and U18345 (N_18345,N_15106,N_16340);
or U18346 (N_18346,N_15444,N_15267);
nor U18347 (N_18347,N_15216,N_15866);
and U18348 (N_18348,N_16117,N_15888);
xnor U18349 (N_18349,N_15044,N_17291);
or U18350 (N_18350,N_15308,N_15447);
or U18351 (N_18351,N_15020,N_16306);
and U18352 (N_18352,N_15633,N_16174);
nand U18353 (N_18353,N_16002,N_16674);
and U18354 (N_18354,N_15757,N_16647);
xor U18355 (N_18355,N_15482,N_15279);
xnor U18356 (N_18356,N_16763,N_15451);
and U18357 (N_18357,N_16003,N_17457);
and U18358 (N_18358,N_15535,N_15370);
and U18359 (N_18359,N_15344,N_17409);
nor U18360 (N_18360,N_16206,N_15657);
or U18361 (N_18361,N_15371,N_17033);
nor U18362 (N_18362,N_15638,N_16406);
and U18363 (N_18363,N_17179,N_16752);
or U18364 (N_18364,N_16120,N_15253);
nor U18365 (N_18365,N_15814,N_16488);
nor U18366 (N_18366,N_17428,N_16805);
or U18367 (N_18367,N_15187,N_15532);
xor U18368 (N_18368,N_17461,N_16988);
and U18369 (N_18369,N_17203,N_15650);
xor U18370 (N_18370,N_16799,N_17304);
xor U18371 (N_18371,N_15973,N_17007);
or U18372 (N_18372,N_16047,N_15219);
nor U18373 (N_18373,N_17424,N_16188);
and U18374 (N_18374,N_16741,N_15553);
nand U18375 (N_18375,N_16603,N_16144);
and U18376 (N_18376,N_15611,N_15467);
and U18377 (N_18377,N_15589,N_15240);
or U18378 (N_18378,N_15292,N_17040);
nor U18379 (N_18379,N_17188,N_17028);
or U18380 (N_18380,N_16304,N_16669);
nand U18381 (N_18381,N_16193,N_16704);
or U18382 (N_18382,N_17316,N_16387);
and U18383 (N_18383,N_17385,N_15024);
nand U18384 (N_18384,N_15966,N_15161);
or U18385 (N_18385,N_16146,N_16025);
nand U18386 (N_18386,N_15945,N_16454);
or U18387 (N_18387,N_15587,N_17392);
or U18388 (N_18388,N_16190,N_15772);
nor U18389 (N_18389,N_15739,N_17087);
nor U18390 (N_18390,N_15974,N_16300);
or U18391 (N_18391,N_15970,N_16933);
nor U18392 (N_18392,N_16568,N_15498);
nor U18393 (N_18393,N_16116,N_16248);
nand U18394 (N_18394,N_16783,N_16596);
nand U18395 (N_18395,N_15439,N_16956);
xnor U18396 (N_18396,N_15314,N_16203);
or U18397 (N_18397,N_15616,N_15740);
nor U18398 (N_18398,N_17469,N_17154);
nor U18399 (N_18399,N_17241,N_16830);
nand U18400 (N_18400,N_15785,N_15499);
xor U18401 (N_18401,N_16019,N_15824);
or U18402 (N_18402,N_16055,N_16736);
nor U18403 (N_18403,N_15130,N_17278);
and U18404 (N_18404,N_17388,N_16570);
xor U18405 (N_18405,N_15609,N_17439);
nor U18406 (N_18406,N_16321,N_17272);
nand U18407 (N_18407,N_17383,N_17244);
nor U18408 (N_18408,N_15608,N_15891);
and U18409 (N_18409,N_15868,N_15141);
and U18410 (N_18410,N_16583,N_15544);
xor U18411 (N_18411,N_15550,N_16127);
nand U18412 (N_18412,N_16906,N_17473);
nand U18413 (N_18413,N_15083,N_16649);
or U18414 (N_18414,N_16904,N_16233);
xor U18415 (N_18415,N_15761,N_15232);
or U18416 (N_18416,N_16087,N_15605);
xnor U18417 (N_18417,N_16090,N_15503);
and U18418 (N_18418,N_16133,N_15593);
or U18419 (N_18419,N_16316,N_15261);
and U18420 (N_18420,N_16365,N_15111);
and U18421 (N_18421,N_15775,N_16612);
and U18422 (N_18422,N_17214,N_17491);
or U18423 (N_18423,N_15669,N_15715);
or U18424 (N_18424,N_17393,N_15298);
nor U18425 (N_18425,N_15210,N_17374);
and U18426 (N_18426,N_16809,N_16989);
or U18427 (N_18427,N_16734,N_15705);
nor U18428 (N_18428,N_17038,N_16362);
nand U18429 (N_18429,N_16547,N_16725);
or U18430 (N_18430,N_16588,N_16715);
or U18431 (N_18431,N_15158,N_15895);
nand U18432 (N_18432,N_17191,N_16962);
nand U18433 (N_18433,N_16890,N_17157);
xnor U18434 (N_18434,N_16968,N_17342);
xor U18435 (N_18435,N_15401,N_15848);
or U18436 (N_18436,N_15918,N_17074);
and U18437 (N_18437,N_15377,N_15526);
or U18438 (N_18438,N_15769,N_15149);
nor U18439 (N_18439,N_17372,N_17197);
nor U18440 (N_18440,N_15662,N_15301);
nor U18441 (N_18441,N_16505,N_16814);
nor U18442 (N_18442,N_17437,N_15215);
nand U18443 (N_18443,N_15003,N_16511);
nand U18444 (N_18444,N_15041,N_16925);
nand U18445 (N_18445,N_15752,N_16923);
and U18446 (N_18446,N_15717,N_17079);
or U18447 (N_18447,N_15163,N_15289);
nor U18448 (N_18448,N_16842,N_15955);
xnor U18449 (N_18449,N_17180,N_15159);
and U18450 (N_18450,N_17387,N_16808);
and U18451 (N_18451,N_15348,N_16716);
nand U18452 (N_18452,N_15993,N_16114);
nor U18453 (N_18453,N_16975,N_17096);
and U18454 (N_18454,N_15075,N_15487);
nor U18455 (N_18455,N_16784,N_16536);
nor U18456 (N_18456,N_16911,N_16791);
xnor U18457 (N_18457,N_17117,N_15822);
or U18458 (N_18458,N_15496,N_16191);
nand U18459 (N_18459,N_16178,N_16351);
nor U18460 (N_18460,N_15121,N_15011);
and U18461 (N_18461,N_16478,N_15017);
or U18462 (N_18462,N_16451,N_15379);
or U18463 (N_18463,N_16823,N_15389);
nand U18464 (N_18464,N_15709,N_16573);
xnor U18465 (N_18465,N_16706,N_16433);
nand U18466 (N_18466,N_17283,N_15548);
or U18467 (N_18467,N_15896,N_15997);
and U18468 (N_18468,N_15512,N_16692);
nor U18469 (N_18469,N_15562,N_17064);
nand U18470 (N_18470,N_15208,N_16349);
xnor U18471 (N_18471,N_16504,N_16074);
or U18472 (N_18472,N_17094,N_16423);
nand U18473 (N_18473,N_16634,N_15721);
and U18474 (N_18474,N_15665,N_16932);
nor U18475 (N_18475,N_16946,N_15309);
xor U18476 (N_18476,N_17018,N_15249);
xor U18477 (N_18477,N_16034,N_15620);
and U18478 (N_18478,N_15450,N_15391);
nor U18479 (N_18479,N_17320,N_16489);
or U18480 (N_18480,N_15898,N_16169);
or U18481 (N_18481,N_16695,N_15364);
nand U18482 (N_18482,N_16179,N_17345);
nand U18483 (N_18483,N_15400,N_15497);
nand U18484 (N_18484,N_16477,N_16927);
nand U18485 (N_18485,N_15726,N_16878);
or U18486 (N_18486,N_17348,N_16942);
and U18487 (N_18487,N_16724,N_15742);
and U18488 (N_18488,N_16126,N_15852);
nor U18489 (N_18489,N_15750,N_16241);
or U18490 (N_18490,N_15751,N_15521);
or U18491 (N_18491,N_16510,N_16535);
nand U18492 (N_18492,N_17490,N_15787);
xor U18493 (N_18493,N_16134,N_15262);
nand U18494 (N_18494,N_16545,N_15047);
and U18495 (N_18495,N_16371,N_16518);
nor U18496 (N_18496,N_16525,N_15956);
nand U18497 (N_18497,N_15429,N_16311);
xnor U18498 (N_18498,N_16118,N_15195);
xor U18499 (N_18499,N_16434,N_17363);
nand U18500 (N_18500,N_16139,N_16993);
xor U18501 (N_18501,N_15182,N_16030);
nand U18502 (N_18502,N_15575,N_16297);
and U18503 (N_18503,N_15576,N_16941);
and U18504 (N_18504,N_16553,N_16051);
and U18505 (N_18505,N_16418,N_15580);
and U18506 (N_18506,N_15747,N_17309);
nor U18507 (N_18507,N_16807,N_17295);
nand U18508 (N_18508,N_17181,N_15122);
nor U18509 (N_18509,N_16856,N_16111);
or U18510 (N_18510,N_15016,N_15784);
or U18511 (N_18511,N_16983,N_15522);
nand U18512 (N_18512,N_15995,N_15469);
xnor U18513 (N_18513,N_17276,N_15124);
xor U18514 (N_18514,N_16040,N_16152);
nand U18515 (N_18515,N_16046,N_15235);
xnor U18516 (N_18516,N_17499,N_15471);
or U18517 (N_18517,N_16010,N_16360);
nor U18518 (N_18518,N_16576,N_16049);
or U18519 (N_18519,N_15091,N_17166);
or U18520 (N_18520,N_15274,N_15399);
nor U18521 (N_18521,N_16882,N_15867);
nor U18522 (N_18522,N_16728,N_16867);
nand U18523 (N_18523,N_15894,N_15644);
nand U18524 (N_18524,N_16097,N_15545);
nand U18525 (N_18525,N_15859,N_15324);
nor U18526 (N_18526,N_16688,N_16827);
and U18527 (N_18527,N_15988,N_16982);
xor U18528 (N_18528,N_15577,N_16305);
nor U18529 (N_18529,N_15771,N_17329);
or U18530 (N_18530,N_16512,N_17069);
nor U18531 (N_18531,N_15009,N_15239);
nor U18532 (N_18532,N_15086,N_16079);
nand U18533 (N_18533,N_17032,N_17277);
xor U18534 (N_18534,N_15903,N_15341);
and U18535 (N_18535,N_16376,N_16386);
xnor U18536 (N_18536,N_17086,N_16112);
and U18537 (N_18537,N_15010,N_16217);
nand U18538 (N_18538,N_16066,N_16338);
nor U18539 (N_18539,N_15430,N_15937);
and U18540 (N_18540,N_15505,N_16271);
nand U18541 (N_18541,N_15488,N_17215);
xnor U18542 (N_18542,N_16515,N_16181);
nand U18543 (N_18543,N_17403,N_16373);
nand U18544 (N_18544,N_16981,N_17039);
xnor U18545 (N_18545,N_17263,N_15630);
nor U18546 (N_18546,N_16249,N_16976);
nor U18547 (N_18547,N_15658,N_15509);
or U18548 (N_18548,N_15963,N_17100);
and U18549 (N_18549,N_16837,N_17418);
xnor U18550 (N_18550,N_16356,N_16251);
nor U18551 (N_18551,N_16839,N_15113);
nand U18552 (N_18552,N_15549,N_15733);
nand U18553 (N_18553,N_15777,N_15190);
nor U18554 (N_18554,N_16421,N_15317);
or U18555 (N_18555,N_15516,N_15426);
and U18556 (N_18556,N_16254,N_17285);
and U18557 (N_18557,N_17338,N_15080);
and U18558 (N_18558,N_17078,N_15983);
or U18559 (N_18559,N_15590,N_15368);
or U18560 (N_18560,N_15064,N_16132);
and U18561 (N_18561,N_17170,N_16105);
and U18562 (N_18562,N_16124,N_16289);
or U18563 (N_18563,N_15329,N_16948);
xnor U18564 (N_18564,N_15604,N_16461);
nor U18565 (N_18565,N_16484,N_17232);
or U18566 (N_18566,N_15316,N_17460);
xor U18567 (N_18567,N_15418,N_15720);
xor U18568 (N_18568,N_16021,N_16565);
nor U18569 (N_18569,N_17346,N_15135);
and U18570 (N_18570,N_17071,N_15085);
nor U18571 (N_18571,N_15311,N_15679);
and U18572 (N_18572,N_17083,N_17446);
xor U18573 (N_18573,N_17315,N_17242);
or U18574 (N_18574,N_15452,N_16869);
nor U18575 (N_18575,N_17045,N_15833);
and U18576 (N_18576,N_15623,N_15238);
nor U18577 (N_18577,N_17398,N_16723);
nand U18578 (N_18578,N_16614,N_17161);
nand U18579 (N_18579,N_15272,N_16395);
nand U18580 (N_18580,N_17317,N_16987);
or U18581 (N_18581,N_16701,N_15543);
nand U18582 (N_18582,N_15458,N_16352);
nand U18583 (N_18583,N_16281,N_16578);
nor U18584 (N_18584,N_17164,N_17193);
or U18585 (N_18585,N_15969,N_16065);
nand U18586 (N_18586,N_15907,N_16953);
or U18587 (N_18587,N_16048,N_16171);
xnor U18588 (N_18588,N_16283,N_15922);
and U18589 (N_18589,N_16018,N_16081);
or U18590 (N_18590,N_16458,N_15749);
nor U18591 (N_18591,N_15634,N_16448);
xnor U18592 (N_18592,N_16227,N_16730);
nand U18593 (N_18593,N_15087,N_15764);
and U18594 (N_18594,N_15900,N_16888);
and U18595 (N_18595,N_17307,N_15614);
nand U18596 (N_18596,N_15841,N_16718);
or U18597 (N_18597,N_16070,N_16739);
or U18598 (N_18598,N_17171,N_15930);
nor U18599 (N_18599,N_15462,N_15736);
xor U18600 (N_18600,N_17472,N_16196);
or U18601 (N_18601,N_16663,N_17046);
or U18602 (N_18602,N_16770,N_16350);
nor U18603 (N_18603,N_16709,N_15629);
and U18604 (N_18604,N_15795,N_15860);
xnor U18605 (N_18605,N_16994,N_17153);
and U18606 (N_18606,N_16848,N_16409);
xnor U18607 (N_18607,N_15882,N_15820);
and U18608 (N_18608,N_16922,N_16549);
nand U18609 (N_18609,N_17015,N_16671);
and U18610 (N_18610,N_15731,N_16160);
and U18611 (N_18611,N_17003,N_15914);
and U18612 (N_18612,N_16493,N_16610);
nand U18613 (N_18613,N_15466,N_15637);
xnor U18614 (N_18614,N_16007,N_16470);
or U18615 (N_18615,N_16773,N_15661);
xor U18616 (N_18616,N_15815,N_15734);
or U18617 (N_18617,N_16632,N_15718);
or U18618 (N_18618,N_16312,N_16969);
xnor U18619 (N_18619,N_15694,N_15843);
nand U18620 (N_18620,N_15984,N_16531);
or U18621 (N_18621,N_16918,N_17178);
nand U18622 (N_18622,N_15183,N_15495);
xnor U18623 (N_18623,N_15125,N_16516);
nand U18624 (N_18624,N_17396,N_15383);
xnor U18625 (N_18625,N_15767,N_16996);
or U18626 (N_18626,N_17200,N_15690);
nor U18627 (N_18627,N_15856,N_15071);
nor U18628 (N_18628,N_16056,N_16292);
and U18629 (N_18629,N_17201,N_17105);
or U18630 (N_18630,N_16681,N_15552);
nor U18631 (N_18631,N_17402,N_16299);
nand U18632 (N_18632,N_17349,N_16963);
or U18633 (N_18633,N_17198,N_15703);
xnor U18634 (N_18634,N_16790,N_15029);
xnor U18635 (N_18635,N_16689,N_16001);
nand U18636 (N_18636,N_16920,N_16793);
xor U18637 (N_18637,N_17362,N_17368);
xnor U18638 (N_18638,N_16530,N_17431);
nor U18639 (N_18639,N_16984,N_16954);
nand U18640 (N_18640,N_16621,N_17139);
xor U18641 (N_18641,N_15759,N_17095);
xor U18642 (N_18642,N_17159,N_17019);
nand U18643 (N_18643,N_16717,N_16308);
nand U18644 (N_18644,N_16207,N_16384);
nor U18645 (N_18645,N_15753,N_16855);
nor U18646 (N_18646,N_15524,N_15910);
nand U18647 (N_18647,N_15229,N_16631);
nand U18648 (N_18648,N_15809,N_15194);
or U18649 (N_18649,N_16319,N_16584);
xor U18650 (N_18650,N_15830,N_16158);
or U18651 (N_18651,N_17360,N_17448);
nand U18652 (N_18652,N_15477,N_17327);
and U18653 (N_18653,N_17264,N_15844);
or U18654 (N_18654,N_15618,N_15323);
xnor U18655 (N_18655,N_16235,N_15601);
xnor U18656 (N_18656,N_16411,N_16424);
nor U18657 (N_18657,N_16901,N_15188);
and U18658 (N_18658,N_16415,N_15038);
nor U18659 (N_18659,N_16707,N_15821);
or U18660 (N_18660,N_16861,N_15380);
or U18661 (N_18661,N_15806,N_15296);
nor U18662 (N_18662,N_17326,N_17067);
nand U18663 (N_18663,N_15653,N_16108);
or U18664 (N_18664,N_16712,N_16246);
nand U18665 (N_18665,N_16686,N_16571);
or U18666 (N_18666,N_15297,N_16625);
or U18667 (N_18667,N_16234,N_15776);
and U18668 (N_18668,N_17000,N_16539);
and U18669 (N_18669,N_15492,N_16110);
nand U18670 (N_18670,N_15245,N_16167);
nor U18671 (N_18671,N_16668,N_16828);
and U18672 (N_18672,N_17454,N_15812);
and U18673 (N_18673,N_17286,N_16899);
nor U18674 (N_18674,N_16642,N_16722);
and U18675 (N_18675,N_16874,N_16027);
nand U18676 (N_18676,N_15886,N_16324);
and U18677 (N_18677,N_15352,N_15037);
nand U18678 (N_18678,N_16756,N_17365);
or U18679 (N_18679,N_15728,N_15068);
or U18680 (N_18680,N_16310,N_17367);
xnor U18681 (N_18681,N_15259,N_15908);
or U18682 (N_18682,N_16751,N_16744);
and U18683 (N_18683,N_15218,N_16183);
nand U18684 (N_18684,N_17340,N_16277);
nor U18685 (N_18685,N_15871,N_16743);
nand U18686 (N_18686,N_16412,N_16833);
nand U18687 (N_18687,N_15536,N_15284);
nand U18688 (N_18688,N_17478,N_16693);
or U18689 (N_18689,N_16345,N_15002);
nand U18690 (N_18690,N_15098,N_16247);
and U18691 (N_18691,N_16876,N_15754);
nand U18692 (N_18692,N_17378,N_15588);
nand U18693 (N_18693,N_16058,N_15099);
and U18694 (N_18694,N_15932,N_16315);
and U18695 (N_18695,N_15943,N_15356);
nor U18696 (N_18696,N_17134,N_15940);
nor U18697 (N_18697,N_15336,N_17445);
xor U18698 (N_18698,N_17089,N_15834);
nand U18699 (N_18699,N_15897,N_17255);
and U18700 (N_18700,N_16753,N_16810);
xnor U18701 (N_18701,N_15115,N_16769);
or U18702 (N_18702,N_16208,N_16846);
xnor U18703 (N_18703,N_15624,N_15501);
and U18704 (N_18704,N_16630,N_16622);
or U18705 (N_18705,N_16098,N_17085);
or U18706 (N_18706,N_16088,N_16382);
xnor U18707 (N_18707,N_15434,N_15678);
nor U18708 (N_18708,N_16364,N_15668);
or U18709 (N_18709,N_15193,N_15045);
or U18710 (N_18710,N_17207,N_16335);
nand U18711 (N_18711,N_15191,N_15070);
and U18712 (N_18712,N_16533,N_17025);
or U18713 (N_18713,N_17175,N_15884);
nand U18714 (N_18714,N_15622,N_16690);
or U18715 (N_18715,N_17225,N_16187);
nand U18716 (N_18716,N_15361,N_17062);
or U18717 (N_18717,N_16820,N_17459);
nor U18718 (N_18718,N_17012,N_17195);
xor U18719 (N_18719,N_17270,N_15347);
or U18720 (N_18720,N_15385,N_17335);
nand U18721 (N_18721,N_16414,N_15438);
xnor U18722 (N_18722,N_15335,N_17289);
xnor U18723 (N_18723,N_15103,N_16326);
xnor U18724 (N_18724,N_15676,N_15596);
nand U18725 (N_18725,N_15954,N_15152);
xor U18726 (N_18726,N_16180,N_16162);
nand U18727 (N_18727,N_15432,N_16347);
nand U18728 (N_18728,N_16940,N_16143);
or U18729 (N_18729,N_15874,N_16579);
xor U18730 (N_18730,N_16787,N_15416);
or U18731 (N_18731,N_15026,N_15257);
and U18732 (N_18732,N_16257,N_16209);
or U18733 (N_18733,N_16441,N_15508);
xor U18734 (N_18734,N_15735,N_15923);
or U18735 (N_18735,N_15260,N_16464);
nor U18736 (N_18736,N_17088,N_17298);
or U18737 (N_18737,N_17498,N_16446);
xnor U18738 (N_18738,N_17296,N_16507);
xor U18739 (N_18739,N_16024,N_17092);
nand U18740 (N_18740,N_17394,N_16834);
or U18741 (N_18741,N_17103,N_15557);
xor U18742 (N_18742,N_16182,N_15359);
and U18743 (N_18743,N_15686,N_16651);
and U18744 (N_18744,N_16815,N_16429);
nor U18745 (N_18745,N_16691,N_16095);
or U18746 (N_18746,N_17220,N_16138);
or U18747 (N_18747,N_15397,N_16113);
nor U18748 (N_18748,N_16700,N_17292);
xnor U18749 (N_18749,N_15837,N_15861);
nand U18750 (N_18750,N_16595,N_15403);
xor U18751 (N_18751,N_15784,N_15849);
xnor U18752 (N_18752,N_15601,N_16009);
nand U18753 (N_18753,N_16627,N_15302);
xnor U18754 (N_18754,N_16794,N_16608);
nand U18755 (N_18755,N_17180,N_15986);
xor U18756 (N_18756,N_16133,N_15719);
or U18757 (N_18757,N_15723,N_16321);
nand U18758 (N_18758,N_16673,N_16696);
or U18759 (N_18759,N_17299,N_17202);
or U18760 (N_18760,N_17020,N_16779);
nor U18761 (N_18761,N_15717,N_16014);
xnor U18762 (N_18762,N_17064,N_16158);
nand U18763 (N_18763,N_17307,N_15516);
nor U18764 (N_18764,N_16875,N_15321);
or U18765 (N_18765,N_15487,N_16398);
or U18766 (N_18766,N_16653,N_17334);
nor U18767 (N_18767,N_17148,N_15692);
nor U18768 (N_18768,N_17260,N_15272);
or U18769 (N_18769,N_17289,N_16725);
or U18770 (N_18770,N_16478,N_15530);
or U18771 (N_18771,N_15136,N_16369);
nor U18772 (N_18772,N_16021,N_15483);
and U18773 (N_18773,N_16708,N_15655);
and U18774 (N_18774,N_16415,N_17118);
nand U18775 (N_18775,N_16628,N_16573);
nor U18776 (N_18776,N_16421,N_16921);
nand U18777 (N_18777,N_16899,N_15007);
xnor U18778 (N_18778,N_15081,N_16169);
xor U18779 (N_18779,N_17466,N_15529);
and U18780 (N_18780,N_15387,N_17450);
nor U18781 (N_18781,N_15017,N_15277);
nor U18782 (N_18782,N_16800,N_17437);
nor U18783 (N_18783,N_15483,N_15348);
nand U18784 (N_18784,N_16703,N_17450);
nand U18785 (N_18785,N_15505,N_15799);
xnor U18786 (N_18786,N_16347,N_16221);
nor U18787 (N_18787,N_15600,N_16541);
or U18788 (N_18788,N_15354,N_17299);
nand U18789 (N_18789,N_17455,N_15915);
or U18790 (N_18790,N_15629,N_17026);
xnor U18791 (N_18791,N_16546,N_15534);
or U18792 (N_18792,N_16267,N_15459);
nor U18793 (N_18793,N_16299,N_16093);
nand U18794 (N_18794,N_16411,N_16703);
xnor U18795 (N_18795,N_16154,N_15243);
nand U18796 (N_18796,N_17484,N_16858);
and U18797 (N_18797,N_15301,N_15285);
xnor U18798 (N_18798,N_16864,N_15115);
xnor U18799 (N_18799,N_17158,N_17182);
and U18800 (N_18800,N_16683,N_17373);
xor U18801 (N_18801,N_16010,N_15540);
nor U18802 (N_18802,N_16672,N_16417);
or U18803 (N_18803,N_15449,N_17424);
and U18804 (N_18804,N_16297,N_16338);
xor U18805 (N_18805,N_15196,N_15022);
and U18806 (N_18806,N_16930,N_15943);
nand U18807 (N_18807,N_15912,N_15446);
xor U18808 (N_18808,N_16615,N_17340);
xor U18809 (N_18809,N_17245,N_17288);
or U18810 (N_18810,N_17389,N_16928);
xor U18811 (N_18811,N_15062,N_16671);
or U18812 (N_18812,N_16132,N_16974);
xnor U18813 (N_18813,N_15791,N_16962);
nor U18814 (N_18814,N_15434,N_15044);
nor U18815 (N_18815,N_16597,N_15798);
or U18816 (N_18816,N_16967,N_15256);
nand U18817 (N_18817,N_15080,N_16460);
xor U18818 (N_18818,N_16864,N_15312);
nand U18819 (N_18819,N_16946,N_16819);
or U18820 (N_18820,N_17142,N_16481);
nor U18821 (N_18821,N_17030,N_17175);
nor U18822 (N_18822,N_17017,N_15979);
xor U18823 (N_18823,N_17367,N_16184);
nand U18824 (N_18824,N_16152,N_15385);
and U18825 (N_18825,N_15857,N_16651);
nor U18826 (N_18826,N_15968,N_17241);
nor U18827 (N_18827,N_15111,N_15152);
or U18828 (N_18828,N_15932,N_15215);
nand U18829 (N_18829,N_16190,N_17289);
nand U18830 (N_18830,N_15009,N_16820);
or U18831 (N_18831,N_15280,N_16241);
and U18832 (N_18832,N_15782,N_15789);
nor U18833 (N_18833,N_15210,N_16620);
xor U18834 (N_18834,N_17026,N_17426);
and U18835 (N_18835,N_15402,N_15987);
and U18836 (N_18836,N_15913,N_17242);
nor U18837 (N_18837,N_16559,N_15928);
or U18838 (N_18838,N_16981,N_15122);
and U18839 (N_18839,N_17304,N_16650);
nor U18840 (N_18840,N_16861,N_16609);
xnor U18841 (N_18841,N_16714,N_16381);
and U18842 (N_18842,N_15466,N_15384);
xnor U18843 (N_18843,N_16004,N_15892);
nor U18844 (N_18844,N_16584,N_15143);
or U18845 (N_18845,N_15427,N_15715);
or U18846 (N_18846,N_15055,N_16634);
xor U18847 (N_18847,N_15772,N_16001);
nand U18848 (N_18848,N_16638,N_15184);
nor U18849 (N_18849,N_16157,N_16499);
xor U18850 (N_18850,N_17470,N_17395);
xnor U18851 (N_18851,N_15498,N_15272);
nor U18852 (N_18852,N_17442,N_16348);
and U18853 (N_18853,N_16212,N_16617);
nand U18854 (N_18854,N_15076,N_15116);
xor U18855 (N_18855,N_16073,N_17491);
xor U18856 (N_18856,N_17435,N_17037);
nand U18857 (N_18857,N_16409,N_15624);
or U18858 (N_18858,N_16867,N_16083);
xor U18859 (N_18859,N_15020,N_17196);
or U18860 (N_18860,N_15211,N_15540);
nor U18861 (N_18861,N_16658,N_15261);
xor U18862 (N_18862,N_16947,N_17383);
and U18863 (N_18863,N_16062,N_16643);
nor U18864 (N_18864,N_15824,N_16074);
nand U18865 (N_18865,N_16172,N_16549);
xor U18866 (N_18866,N_16102,N_15371);
xnor U18867 (N_18867,N_15120,N_16778);
or U18868 (N_18868,N_17220,N_16839);
nand U18869 (N_18869,N_17375,N_15372);
xnor U18870 (N_18870,N_15460,N_15739);
nand U18871 (N_18871,N_15696,N_16744);
xnor U18872 (N_18872,N_17307,N_17470);
nand U18873 (N_18873,N_16037,N_15120);
nand U18874 (N_18874,N_15155,N_15883);
nand U18875 (N_18875,N_16416,N_16822);
or U18876 (N_18876,N_16423,N_17448);
xor U18877 (N_18877,N_15184,N_16315);
or U18878 (N_18878,N_17015,N_17456);
nor U18879 (N_18879,N_16697,N_16542);
nor U18880 (N_18880,N_16863,N_16635);
and U18881 (N_18881,N_17473,N_16577);
xnor U18882 (N_18882,N_15247,N_16169);
nand U18883 (N_18883,N_16714,N_15643);
nor U18884 (N_18884,N_17487,N_16506);
nor U18885 (N_18885,N_16428,N_16593);
or U18886 (N_18886,N_17176,N_16759);
xor U18887 (N_18887,N_15979,N_16739);
or U18888 (N_18888,N_15553,N_15678);
nand U18889 (N_18889,N_15883,N_15149);
xnor U18890 (N_18890,N_16615,N_15069);
or U18891 (N_18891,N_16413,N_17172);
xnor U18892 (N_18892,N_16577,N_17143);
nand U18893 (N_18893,N_15634,N_15292);
xor U18894 (N_18894,N_15715,N_16253);
and U18895 (N_18895,N_16094,N_16217);
or U18896 (N_18896,N_17204,N_16883);
nor U18897 (N_18897,N_17332,N_15397);
or U18898 (N_18898,N_15231,N_16988);
and U18899 (N_18899,N_15942,N_16916);
nor U18900 (N_18900,N_16915,N_15423);
nor U18901 (N_18901,N_17140,N_15562);
and U18902 (N_18902,N_15275,N_15876);
nor U18903 (N_18903,N_15398,N_16112);
xor U18904 (N_18904,N_16295,N_16764);
nand U18905 (N_18905,N_17052,N_16039);
nand U18906 (N_18906,N_16559,N_15083);
or U18907 (N_18907,N_16027,N_15771);
nor U18908 (N_18908,N_15981,N_17449);
nand U18909 (N_18909,N_15338,N_16229);
nand U18910 (N_18910,N_15154,N_17179);
xnor U18911 (N_18911,N_17131,N_17054);
and U18912 (N_18912,N_16094,N_15553);
nand U18913 (N_18913,N_15566,N_17411);
xnor U18914 (N_18914,N_16746,N_17487);
xor U18915 (N_18915,N_15667,N_16205);
and U18916 (N_18916,N_15374,N_15595);
nor U18917 (N_18917,N_16471,N_15930);
and U18918 (N_18918,N_15977,N_15385);
nand U18919 (N_18919,N_15264,N_16501);
and U18920 (N_18920,N_16818,N_16497);
nand U18921 (N_18921,N_16685,N_16798);
and U18922 (N_18922,N_15763,N_16096);
nand U18923 (N_18923,N_16649,N_16394);
nor U18924 (N_18924,N_17248,N_15895);
xor U18925 (N_18925,N_15455,N_17043);
xor U18926 (N_18926,N_16407,N_16192);
xor U18927 (N_18927,N_16495,N_17071);
and U18928 (N_18928,N_15617,N_16138);
nor U18929 (N_18929,N_15530,N_16743);
xor U18930 (N_18930,N_15669,N_16039);
nand U18931 (N_18931,N_17044,N_16093);
nor U18932 (N_18932,N_17460,N_16883);
xor U18933 (N_18933,N_15119,N_15072);
or U18934 (N_18934,N_17333,N_17112);
and U18935 (N_18935,N_16739,N_17461);
xnor U18936 (N_18936,N_16145,N_16049);
nand U18937 (N_18937,N_15757,N_16177);
and U18938 (N_18938,N_16057,N_16276);
nand U18939 (N_18939,N_16949,N_16992);
or U18940 (N_18940,N_15372,N_15562);
or U18941 (N_18941,N_16093,N_15735);
and U18942 (N_18942,N_16022,N_16358);
or U18943 (N_18943,N_16324,N_17188);
xnor U18944 (N_18944,N_16319,N_15671);
or U18945 (N_18945,N_17428,N_17285);
xor U18946 (N_18946,N_15610,N_16537);
xor U18947 (N_18947,N_16321,N_16715);
xnor U18948 (N_18948,N_15435,N_15734);
nand U18949 (N_18949,N_17358,N_15078);
nand U18950 (N_18950,N_15227,N_15664);
nand U18951 (N_18951,N_16485,N_17049);
nor U18952 (N_18952,N_15817,N_16744);
and U18953 (N_18953,N_17274,N_16875);
or U18954 (N_18954,N_15796,N_16289);
xnor U18955 (N_18955,N_16404,N_16396);
nand U18956 (N_18956,N_17460,N_17047);
or U18957 (N_18957,N_15294,N_16800);
and U18958 (N_18958,N_17167,N_16838);
and U18959 (N_18959,N_15815,N_16788);
nand U18960 (N_18960,N_15010,N_16737);
nor U18961 (N_18961,N_16972,N_17373);
xor U18962 (N_18962,N_15703,N_15487);
and U18963 (N_18963,N_17100,N_15661);
xor U18964 (N_18964,N_15876,N_15197);
or U18965 (N_18965,N_17409,N_15637);
and U18966 (N_18966,N_15613,N_15076);
nor U18967 (N_18967,N_17409,N_16603);
xor U18968 (N_18968,N_16484,N_15001);
nand U18969 (N_18969,N_16372,N_16409);
nor U18970 (N_18970,N_16406,N_17001);
xnor U18971 (N_18971,N_17041,N_17339);
nand U18972 (N_18972,N_16344,N_16273);
nand U18973 (N_18973,N_15836,N_15659);
xor U18974 (N_18974,N_15372,N_15028);
and U18975 (N_18975,N_16849,N_17026);
or U18976 (N_18976,N_15307,N_16306);
nand U18977 (N_18977,N_15834,N_17424);
or U18978 (N_18978,N_15346,N_17317);
xor U18979 (N_18979,N_16774,N_16948);
and U18980 (N_18980,N_17348,N_15486);
and U18981 (N_18981,N_15877,N_16395);
or U18982 (N_18982,N_16503,N_16444);
nor U18983 (N_18983,N_16920,N_16657);
nand U18984 (N_18984,N_16675,N_16692);
nand U18985 (N_18985,N_16474,N_15461);
and U18986 (N_18986,N_17020,N_15241);
xnor U18987 (N_18987,N_15307,N_15914);
xor U18988 (N_18988,N_17344,N_16022);
and U18989 (N_18989,N_16430,N_15135);
xnor U18990 (N_18990,N_16824,N_15426);
or U18991 (N_18991,N_15019,N_16093);
xnor U18992 (N_18992,N_17088,N_16702);
nand U18993 (N_18993,N_17387,N_16051);
nor U18994 (N_18994,N_16810,N_16200);
xor U18995 (N_18995,N_17340,N_16883);
xnor U18996 (N_18996,N_16208,N_16070);
and U18997 (N_18997,N_15333,N_15219);
nor U18998 (N_18998,N_15905,N_15688);
xnor U18999 (N_18999,N_15024,N_16832);
or U19000 (N_19000,N_15211,N_16240);
or U19001 (N_19001,N_16689,N_17148);
or U19002 (N_19002,N_17171,N_16805);
and U19003 (N_19003,N_16387,N_15236);
nand U19004 (N_19004,N_16608,N_15263);
nor U19005 (N_19005,N_17361,N_16022);
and U19006 (N_19006,N_15691,N_16106);
xnor U19007 (N_19007,N_16804,N_16776);
or U19008 (N_19008,N_16189,N_15667);
nand U19009 (N_19009,N_16516,N_17300);
nand U19010 (N_19010,N_15370,N_15869);
and U19011 (N_19011,N_15555,N_15614);
nand U19012 (N_19012,N_17265,N_15168);
and U19013 (N_19013,N_15726,N_17357);
or U19014 (N_19014,N_16428,N_15206);
and U19015 (N_19015,N_17042,N_16087);
or U19016 (N_19016,N_15270,N_15383);
nand U19017 (N_19017,N_17492,N_15836);
nand U19018 (N_19018,N_16823,N_15862);
and U19019 (N_19019,N_16182,N_16806);
and U19020 (N_19020,N_16820,N_15741);
xor U19021 (N_19021,N_15124,N_16512);
xor U19022 (N_19022,N_16777,N_15777);
nor U19023 (N_19023,N_16127,N_16953);
and U19024 (N_19024,N_16991,N_16360);
or U19025 (N_19025,N_15780,N_16282);
and U19026 (N_19026,N_15207,N_16243);
and U19027 (N_19027,N_17003,N_16229);
and U19028 (N_19028,N_16159,N_16177);
xor U19029 (N_19029,N_16095,N_15629);
and U19030 (N_19030,N_15841,N_16550);
and U19031 (N_19031,N_17163,N_16166);
xor U19032 (N_19032,N_15459,N_17342);
and U19033 (N_19033,N_16949,N_15691);
xor U19034 (N_19034,N_15806,N_15664);
and U19035 (N_19035,N_16352,N_16652);
or U19036 (N_19036,N_15995,N_16444);
nor U19037 (N_19037,N_15229,N_15955);
nand U19038 (N_19038,N_15637,N_15288);
and U19039 (N_19039,N_15882,N_17302);
xor U19040 (N_19040,N_16900,N_17395);
and U19041 (N_19041,N_16658,N_17078);
and U19042 (N_19042,N_15117,N_15689);
xor U19043 (N_19043,N_17011,N_17434);
and U19044 (N_19044,N_15631,N_16838);
nor U19045 (N_19045,N_15437,N_16173);
nor U19046 (N_19046,N_15556,N_16756);
and U19047 (N_19047,N_15289,N_15778);
or U19048 (N_19048,N_17003,N_17141);
or U19049 (N_19049,N_16352,N_16460);
or U19050 (N_19050,N_15559,N_16053);
xnor U19051 (N_19051,N_16253,N_15678);
xor U19052 (N_19052,N_16756,N_16939);
nor U19053 (N_19053,N_16435,N_16069);
xor U19054 (N_19054,N_16389,N_16676);
xnor U19055 (N_19055,N_16319,N_17088);
or U19056 (N_19056,N_15091,N_16105);
nor U19057 (N_19057,N_16496,N_16910);
nand U19058 (N_19058,N_16231,N_16948);
xor U19059 (N_19059,N_15317,N_17187);
nand U19060 (N_19060,N_15706,N_16568);
nand U19061 (N_19061,N_16919,N_17131);
or U19062 (N_19062,N_16969,N_16663);
xor U19063 (N_19063,N_16756,N_17318);
or U19064 (N_19064,N_15861,N_16390);
and U19065 (N_19065,N_16921,N_17196);
xor U19066 (N_19066,N_15273,N_17231);
nand U19067 (N_19067,N_16170,N_16453);
and U19068 (N_19068,N_16332,N_15433);
and U19069 (N_19069,N_17296,N_15594);
nor U19070 (N_19070,N_15760,N_16792);
or U19071 (N_19071,N_15130,N_15569);
xnor U19072 (N_19072,N_15898,N_15756);
and U19073 (N_19073,N_17003,N_15357);
nand U19074 (N_19074,N_17357,N_15775);
nand U19075 (N_19075,N_15054,N_15914);
nor U19076 (N_19076,N_15906,N_17367);
and U19077 (N_19077,N_16051,N_15370);
nand U19078 (N_19078,N_15208,N_17256);
xnor U19079 (N_19079,N_15330,N_15871);
and U19080 (N_19080,N_16857,N_15235);
nor U19081 (N_19081,N_16989,N_16150);
nor U19082 (N_19082,N_15901,N_16971);
nor U19083 (N_19083,N_15710,N_17343);
xnor U19084 (N_19084,N_15235,N_16545);
nor U19085 (N_19085,N_15085,N_16579);
or U19086 (N_19086,N_15791,N_16844);
or U19087 (N_19087,N_17486,N_16393);
and U19088 (N_19088,N_15249,N_15709);
xor U19089 (N_19089,N_16971,N_15970);
nand U19090 (N_19090,N_16912,N_17101);
nor U19091 (N_19091,N_17129,N_15709);
xnor U19092 (N_19092,N_17451,N_16878);
nor U19093 (N_19093,N_15356,N_16528);
nor U19094 (N_19094,N_16190,N_15411);
or U19095 (N_19095,N_15275,N_17062);
xnor U19096 (N_19096,N_16622,N_17430);
nand U19097 (N_19097,N_16610,N_15332);
nor U19098 (N_19098,N_16354,N_17320);
or U19099 (N_19099,N_16115,N_15796);
or U19100 (N_19100,N_16615,N_15787);
nor U19101 (N_19101,N_15493,N_16682);
nor U19102 (N_19102,N_16054,N_16269);
xnor U19103 (N_19103,N_15008,N_15107);
nand U19104 (N_19104,N_15144,N_15121);
xor U19105 (N_19105,N_16757,N_15190);
xnor U19106 (N_19106,N_15264,N_15173);
nand U19107 (N_19107,N_17089,N_16628);
or U19108 (N_19108,N_17269,N_15989);
nand U19109 (N_19109,N_15157,N_17440);
xnor U19110 (N_19110,N_17382,N_15443);
nor U19111 (N_19111,N_16269,N_17072);
nor U19112 (N_19112,N_16441,N_17003);
or U19113 (N_19113,N_15424,N_17199);
and U19114 (N_19114,N_17206,N_17440);
and U19115 (N_19115,N_17073,N_15375);
nor U19116 (N_19116,N_16290,N_16398);
nor U19117 (N_19117,N_16774,N_15200);
xor U19118 (N_19118,N_16555,N_16158);
or U19119 (N_19119,N_15644,N_16325);
or U19120 (N_19120,N_15482,N_15006);
and U19121 (N_19121,N_17182,N_16390);
nand U19122 (N_19122,N_15958,N_15565);
xor U19123 (N_19123,N_15096,N_17470);
xnor U19124 (N_19124,N_16776,N_17351);
xnor U19125 (N_19125,N_16877,N_16695);
nor U19126 (N_19126,N_17240,N_17037);
nor U19127 (N_19127,N_15349,N_16983);
or U19128 (N_19128,N_16444,N_16311);
nor U19129 (N_19129,N_16059,N_16292);
nand U19130 (N_19130,N_15418,N_15339);
nor U19131 (N_19131,N_16466,N_16884);
xnor U19132 (N_19132,N_16654,N_16451);
nand U19133 (N_19133,N_15111,N_17298);
and U19134 (N_19134,N_15886,N_16576);
nand U19135 (N_19135,N_15148,N_15691);
nor U19136 (N_19136,N_16506,N_15563);
nor U19137 (N_19137,N_16418,N_16629);
and U19138 (N_19138,N_17120,N_15647);
nor U19139 (N_19139,N_16606,N_16897);
and U19140 (N_19140,N_16330,N_17303);
nor U19141 (N_19141,N_17095,N_15419);
or U19142 (N_19142,N_16429,N_15902);
nand U19143 (N_19143,N_16835,N_16868);
and U19144 (N_19144,N_17146,N_15218);
nor U19145 (N_19145,N_17387,N_17338);
nor U19146 (N_19146,N_15393,N_15431);
and U19147 (N_19147,N_17060,N_17231);
nor U19148 (N_19148,N_16180,N_15442);
nand U19149 (N_19149,N_17377,N_15258);
xor U19150 (N_19150,N_16396,N_15166);
or U19151 (N_19151,N_16034,N_15858);
and U19152 (N_19152,N_15362,N_16971);
nor U19153 (N_19153,N_16084,N_16799);
nor U19154 (N_19154,N_15728,N_15503);
nor U19155 (N_19155,N_16736,N_15485);
and U19156 (N_19156,N_16637,N_16333);
and U19157 (N_19157,N_16408,N_17243);
xnor U19158 (N_19158,N_16330,N_15019);
and U19159 (N_19159,N_16812,N_16987);
nand U19160 (N_19160,N_15227,N_16914);
nor U19161 (N_19161,N_15160,N_16980);
nor U19162 (N_19162,N_16081,N_17226);
nor U19163 (N_19163,N_15978,N_15950);
and U19164 (N_19164,N_17480,N_15020);
nor U19165 (N_19165,N_16826,N_17000);
nor U19166 (N_19166,N_15306,N_15301);
nor U19167 (N_19167,N_16914,N_15093);
nor U19168 (N_19168,N_15992,N_15599);
or U19169 (N_19169,N_15029,N_15637);
xor U19170 (N_19170,N_15825,N_15703);
nor U19171 (N_19171,N_15425,N_16055);
or U19172 (N_19172,N_16642,N_17049);
nand U19173 (N_19173,N_16320,N_16331);
nand U19174 (N_19174,N_15651,N_16774);
or U19175 (N_19175,N_16356,N_17352);
or U19176 (N_19176,N_15051,N_16817);
nand U19177 (N_19177,N_17470,N_15827);
xnor U19178 (N_19178,N_15367,N_16558);
and U19179 (N_19179,N_16444,N_16078);
and U19180 (N_19180,N_15917,N_16071);
xor U19181 (N_19181,N_17250,N_16878);
or U19182 (N_19182,N_16954,N_16932);
or U19183 (N_19183,N_16594,N_17477);
nand U19184 (N_19184,N_16098,N_15595);
or U19185 (N_19185,N_15234,N_15306);
nand U19186 (N_19186,N_17037,N_15968);
or U19187 (N_19187,N_17111,N_16493);
xnor U19188 (N_19188,N_16066,N_16128);
nor U19189 (N_19189,N_16626,N_17434);
nor U19190 (N_19190,N_16310,N_16756);
nor U19191 (N_19191,N_15153,N_16944);
nor U19192 (N_19192,N_16184,N_16868);
or U19193 (N_19193,N_17227,N_16659);
nand U19194 (N_19194,N_15515,N_16775);
nand U19195 (N_19195,N_17062,N_16718);
xor U19196 (N_19196,N_16639,N_15147);
xnor U19197 (N_19197,N_15271,N_16799);
xor U19198 (N_19198,N_17103,N_17137);
xor U19199 (N_19199,N_15307,N_16898);
or U19200 (N_19200,N_17104,N_15597);
nand U19201 (N_19201,N_15358,N_15060);
and U19202 (N_19202,N_16176,N_17092);
xnor U19203 (N_19203,N_17305,N_15627);
nand U19204 (N_19204,N_15587,N_15080);
or U19205 (N_19205,N_16455,N_17464);
or U19206 (N_19206,N_15002,N_15501);
or U19207 (N_19207,N_17236,N_16133);
nand U19208 (N_19208,N_15672,N_15355);
nand U19209 (N_19209,N_16240,N_15634);
xnor U19210 (N_19210,N_16030,N_17476);
nand U19211 (N_19211,N_16719,N_16105);
nor U19212 (N_19212,N_15033,N_15723);
or U19213 (N_19213,N_17459,N_15833);
xor U19214 (N_19214,N_16323,N_16664);
xnor U19215 (N_19215,N_16723,N_16107);
nor U19216 (N_19216,N_15094,N_17407);
nor U19217 (N_19217,N_15797,N_17162);
nand U19218 (N_19218,N_17471,N_16149);
nand U19219 (N_19219,N_15010,N_16444);
nand U19220 (N_19220,N_17404,N_15704);
and U19221 (N_19221,N_16485,N_17128);
and U19222 (N_19222,N_15178,N_15866);
or U19223 (N_19223,N_16891,N_15764);
xor U19224 (N_19224,N_15426,N_15023);
nand U19225 (N_19225,N_15688,N_16282);
nand U19226 (N_19226,N_16252,N_16249);
or U19227 (N_19227,N_15087,N_16967);
nand U19228 (N_19228,N_15960,N_15653);
xor U19229 (N_19229,N_15215,N_17177);
nand U19230 (N_19230,N_15284,N_15633);
and U19231 (N_19231,N_16998,N_17326);
and U19232 (N_19232,N_15243,N_17142);
or U19233 (N_19233,N_16921,N_17074);
or U19234 (N_19234,N_17069,N_15762);
xnor U19235 (N_19235,N_16674,N_16017);
nand U19236 (N_19236,N_16149,N_16580);
and U19237 (N_19237,N_16276,N_17324);
and U19238 (N_19238,N_15992,N_15290);
or U19239 (N_19239,N_15835,N_15935);
or U19240 (N_19240,N_16757,N_15295);
nand U19241 (N_19241,N_15314,N_15569);
nand U19242 (N_19242,N_16593,N_16444);
nor U19243 (N_19243,N_17241,N_15529);
and U19244 (N_19244,N_16395,N_16353);
and U19245 (N_19245,N_15248,N_15995);
nor U19246 (N_19246,N_16109,N_17045);
or U19247 (N_19247,N_15234,N_15578);
and U19248 (N_19248,N_16902,N_17303);
nor U19249 (N_19249,N_16495,N_16600);
or U19250 (N_19250,N_16430,N_17393);
and U19251 (N_19251,N_15708,N_16151);
and U19252 (N_19252,N_16546,N_15480);
and U19253 (N_19253,N_15207,N_16693);
xnor U19254 (N_19254,N_15518,N_16027);
xnor U19255 (N_19255,N_16168,N_15846);
or U19256 (N_19256,N_16479,N_16357);
or U19257 (N_19257,N_15158,N_15651);
xnor U19258 (N_19258,N_16256,N_16502);
or U19259 (N_19259,N_16407,N_16540);
or U19260 (N_19260,N_16730,N_16660);
nor U19261 (N_19261,N_15792,N_17425);
or U19262 (N_19262,N_16648,N_16653);
nor U19263 (N_19263,N_17150,N_15401);
nor U19264 (N_19264,N_16883,N_15784);
or U19265 (N_19265,N_17163,N_16941);
xnor U19266 (N_19266,N_15488,N_16583);
and U19267 (N_19267,N_16171,N_15929);
or U19268 (N_19268,N_16969,N_15623);
xnor U19269 (N_19269,N_15916,N_17321);
nor U19270 (N_19270,N_15468,N_16412);
nand U19271 (N_19271,N_16135,N_16654);
nand U19272 (N_19272,N_16470,N_16247);
or U19273 (N_19273,N_17262,N_16357);
nand U19274 (N_19274,N_16968,N_15413);
or U19275 (N_19275,N_17246,N_15401);
nor U19276 (N_19276,N_16687,N_15038);
nand U19277 (N_19277,N_16682,N_16444);
and U19278 (N_19278,N_17363,N_16016);
or U19279 (N_19279,N_15200,N_16819);
xnor U19280 (N_19280,N_15476,N_17442);
nand U19281 (N_19281,N_17064,N_17459);
xnor U19282 (N_19282,N_17282,N_16726);
or U19283 (N_19283,N_16555,N_15607);
nand U19284 (N_19284,N_15199,N_16163);
xnor U19285 (N_19285,N_15757,N_15972);
xor U19286 (N_19286,N_16649,N_17298);
xor U19287 (N_19287,N_16524,N_15409);
or U19288 (N_19288,N_16593,N_16185);
or U19289 (N_19289,N_16301,N_15079);
nor U19290 (N_19290,N_16315,N_15059);
nand U19291 (N_19291,N_16235,N_15128);
and U19292 (N_19292,N_17408,N_15272);
nand U19293 (N_19293,N_15312,N_16394);
and U19294 (N_19294,N_17344,N_15832);
nand U19295 (N_19295,N_15345,N_15774);
and U19296 (N_19296,N_15837,N_17043);
or U19297 (N_19297,N_16916,N_17409);
nand U19298 (N_19298,N_15373,N_15004);
nand U19299 (N_19299,N_15747,N_16666);
nor U19300 (N_19300,N_17271,N_16230);
nand U19301 (N_19301,N_15246,N_16657);
and U19302 (N_19302,N_16820,N_16951);
nand U19303 (N_19303,N_16772,N_15942);
nand U19304 (N_19304,N_17269,N_16168);
and U19305 (N_19305,N_17397,N_15144);
nor U19306 (N_19306,N_15089,N_15037);
or U19307 (N_19307,N_15908,N_15803);
and U19308 (N_19308,N_16533,N_16756);
nor U19309 (N_19309,N_15291,N_16788);
or U19310 (N_19310,N_15466,N_16360);
and U19311 (N_19311,N_15413,N_15162);
and U19312 (N_19312,N_16876,N_15977);
and U19313 (N_19313,N_15896,N_16330);
or U19314 (N_19314,N_16669,N_17421);
nor U19315 (N_19315,N_15339,N_17219);
nor U19316 (N_19316,N_17114,N_16827);
and U19317 (N_19317,N_15097,N_15686);
xor U19318 (N_19318,N_17200,N_16881);
or U19319 (N_19319,N_16921,N_15615);
nor U19320 (N_19320,N_17443,N_16646);
nand U19321 (N_19321,N_17048,N_16404);
and U19322 (N_19322,N_17396,N_16137);
and U19323 (N_19323,N_15275,N_17424);
xor U19324 (N_19324,N_16314,N_15145);
xor U19325 (N_19325,N_15600,N_17465);
or U19326 (N_19326,N_17284,N_16659);
xor U19327 (N_19327,N_17143,N_15331);
nand U19328 (N_19328,N_16693,N_17356);
xnor U19329 (N_19329,N_15708,N_17182);
and U19330 (N_19330,N_15456,N_15069);
nand U19331 (N_19331,N_15616,N_15784);
nor U19332 (N_19332,N_16337,N_16872);
xor U19333 (N_19333,N_16476,N_15878);
nor U19334 (N_19334,N_15471,N_17496);
xor U19335 (N_19335,N_15235,N_17052);
xor U19336 (N_19336,N_16363,N_16045);
or U19337 (N_19337,N_16788,N_15339);
and U19338 (N_19338,N_15534,N_17422);
xor U19339 (N_19339,N_15428,N_15339);
nor U19340 (N_19340,N_15446,N_15268);
xnor U19341 (N_19341,N_17079,N_15023);
or U19342 (N_19342,N_16259,N_16556);
nand U19343 (N_19343,N_15929,N_16968);
xor U19344 (N_19344,N_16480,N_15082);
xor U19345 (N_19345,N_15769,N_17330);
or U19346 (N_19346,N_16230,N_16122);
and U19347 (N_19347,N_15255,N_17197);
xnor U19348 (N_19348,N_16629,N_17002);
nor U19349 (N_19349,N_15028,N_15324);
nor U19350 (N_19350,N_15723,N_15310);
xor U19351 (N_19351,N_15372,N_15648);
xnor U19352 (N_19352,N_16115,N_16362);
and U19353 (N_19353,N_16075,N_15542);
xnor U19354 (N_19354,N_16102,N_16386);
xnor U19355 (N_19355,N_16624,N_15119);
and U19356 (N_19356,N_16565,N_17216);
or U19357 (N_19357,N_15089,N_16731);
or U19358 (N_19358,N_16503,N_17303);
xor U19359 (N_19359,N_17356,N_17102);
or U19360 (N_19360,N_16551,N_17451);
xnor U19361 (N_19361,N_16511,N_17315);
nand U19362 (N_19362,N_16987,N_16768);
and U19363 (N_19363,N_16590,N_17000);
or U19364 (N_19364,N_15600,N_16484);
xor U19365 (N_19365,N_16536,N_15395);
xnor U19366 (N_19366,N_16237,N_16845);
nand U19367 (N_19367,N_16240,N_16775);
or U19368 (N_19368,N_15897,N_15892);
xor U19369 (N_19369,N_15847,N_16376);
or U19370 (N_19370,N_16804,N_15856);
xor U19371 (N_19371,N_16320,N_15037);
nand U19372 (N_19372,N_16737,N_15011);
nand U19373 (N_19373,N_16240,N_16305);
nor U19374 (N_19374,N_16917,N_16554);
and U19375 (N_19375,N_17288,N_17326);
xnor U19376 (N_19376,N_15855,N_15611);
nor U19377 (N_19377,N_15601,N_16567);
nand U19378 (N_19378,N_15215,N_15422);
xor U19379 (N_19379,N_15246,N_16930);
nand U19380 (N_19380,N_17301,N_15180);
or U19381 (N_19381,N_16995,N_17296);
nand U19382 (N_19382,N_15832,N_16080);
nor U19383 (N_19383,N_15320,N_16945);
xnor U19384 (N_19384,N_15563,N_15480);
nor U19385 (N_19385,N_16097,N_16083);
or U19386 (N_19386,N_15667,N_15558);
xor U19387 (N_19387,N_16070,N_16777);
or U19388 (N_19388,N_15744,N_16634);
xor U19389 (N_19389,N_16014,N_17192);
or U19390 (N_19390,N_16749,N_15328);
nor U19391 (N_19391,N_15316,N_15022);
and U19392 (N_19392,N_15107,N_16579);
nand U19393 (N_19393,N_17359,N_16411);
nor U19394 (N_19394,N_15684,N_17302);
xor U19395 (N_19395,N_17265,N_15571);
and U19396 (N_19396,N_17031,N_17305);
and U19397 (N_19397,N_15798,N_16235);
or U19398 (N_19398,N_16563,N_16171);
xor U19399 (N_19399,N_16224,N_16202);
nor U19400 (N_19400,N_16171,N_17490);
and U19401 (N_19401,N_15119,N_16805);
xor U19402 (N_19402,N_16440,N_15462);
nand U19403 (N_19403,N_15826,N_15531);
nor U19404 (N_19404,N_16191,N_15115);
and U19405 (N_19405,N_16506,N_16993);
nand U19406 (N_19406,N_17077,N_15346);
nor U19407 (N_19407,N_16251,N_15120);
xnor U19408 (N_19408,N_16939,N_15799);
and U19409 (N_19409,N_17400,N_16936);
and U19410 (N_19410,N_17472,N_15285);
nor U19411 (N_19411,N_16589,N_16381);
nand U19412 (N_19412,N_15736,N_17384);
nor U19413 (N_19413,N_15274,N_17319);
nand U19414 (N_19414,N_15115,N_16423);
nand U19415 (N_19415,N_15628,N_15956);
xnor U19416 (N_19416,N_17272,N_15242);
xor U19417 (N_19417,N_15391,N_15143);
xor U19418 (N_19418,N_17387,N_15253);
nand U19419 (N_19419,N_16525,N_15336);
nor U19420 (N_19420,N_17037,N_15997);
and U19421 (N_19421,N_15148,N_16540);
and U19422 (N_19422,N_17246,N_15270);
nand U19423 (N_19423,N_15179,N_16845);
nor U19424 (N_19424,N_17241,N_15334);
or U19425 (N_19425,N_16981,N_16500);
nor U19426 (N_19426,N_15350,N_16795);
and U19427 (N_19427,N_16213,N_16459);
nor U19428 (N_19428,N_15574,N_16776);
nor U19429 (N_19429,N_15223,N_15786);
xnor U19430 (N_19430,N_16752,N_15403);
and U19431 (N_19431,N_16707,N_16750);
and U19432 (N_19432,N_16142,N_17455);
or U19433 (N_19433,N_15941,N_16209);
xor U19434 (N_19434,N_15793,N_16261);
and U19435 (N_19435,N_15622,N_16031);
xor U19436 (N_19436,N_16411,N_15333);
xor U19437 (N_19437,N_15794,N_16251);
xnor U19438 (N_19438,N_16191,N_15654);
or U19439 (N_19439,N_16348,N_16104);
and U19440 (N_19440,N_16596,N_15519);
and U19441 (N_19441,N_15977,N_17464);
nand U19442 (N_19442,N_16563,N_15756);
and U19443 (N_19443,N_16861,N_16305);
nand U19444 (N_19444,N_17112,N_15241);
or U19445 (N_19445,N_17463,N_17028);
nor U19446 (N_19446,N_17479,N_16102);
nor U19447 (N_19447,N_15805,N_16311);
nand U19448 (N_19448,N_15792,N_16017);
xor U19449 (N_19449,N_17253,N_16191);
nor U19450 (N_19450,N_16880,N_15759);
or U19451 (N_19451,N_17072,N_16530);
nor U19452 (N_19452,N_15123,N_15387);
and U19453 (N_19453,N_15698,N_16681);
or U19454 (N_19454,N_16456,N_15897);
or U19455 (N_19455,N_17002,N_15676);
nor U19456 (N_19456,N_17157,N_17161);
and U19457 (N_19457,N_16836,N_16920);
and U19458 (N_19458,N_16558,N_15257);
and U19459 (N_19459,N_16126,N_17098);
or U19460 (N_19460,N_15010,N_16928);
nand U19461 (N_19461,N_16711,N_16680);
nor U19462 (N_19462,N_15343,N_16632);
nor U19463 (N_19463,N_15868,N_15740);
or U19464 (N_19464,N_16799,N_15665);
nor U19465 (N_19465,N_15474,N_15354);
xor U19466 (N_19466,N_15327,N_15353);
or U19467 (N_19467,N_16633,N_17475);
nand U19468 (N_19468,N_16332,N_15118);
xor U19469 (N_19469,N_16833,N_15720);
xnor U19470 (N_19470,N_15466,N_15004);
nor U19471 (N_19471,N_17346,N_16253);
or U19472 (N_19472,N_16343,N_15005);
or U19473 (N_19473,N_16573,N_15983);
and U19474 (N_19474,N_16885,N_15380);
or U19475 (N_19475,N_16866,N_15349);
nor U19476 (N_19476,N_17386,N_17260);
nor U19477 (N_19477,N_15790,N_17201);
xor U19478 (N_19478,N_15778,N_16506);
and U19479 (N_19479,N_16833,N_16482);
or U19480 (N_19480,N_15247,N_15846);
xor U19481 (N_19481,N_15983,N_15965);
nor U19482 (N_19482,N_15927,N_17233);
nand U19483 (N_19483,N_16504,N_16709);
and U19484 (N_19484,N_15411,N_16876);
or U19485 (N_19485,N_17408,N_15165);
nor U19486 (N_19486,N_15014,N_17011);
xnor U19487 (N_19487,N_17228,N_15088);
nand U19488 (N_19488,N_15748,N_16002);
or U19489 (N_19489,N_15468,N_17100);
nand U19490 (N_19490,N_17394,N_16175);
and U19491 (N_19491,N_15653,N_15701);
nand U19492 (N_19492,N_17291,N_16611);
nand U19493 (N_19493,N_17467,N_16339);
nor U19494 (N_19494,N_17486,N_15329);
xnor U19495 (N_19495,N_15608,N_15867);
nand U19496 (N_19496,N_16291,N_16678);
xor U19497 (N_19497,N_15164,N_16661);
and U19498 (N_19498,N_15825,N_15206);
xnor U19499 (N_19499,N_15437,N_16598);
xnor U19500 (N_19500,N_15771,N_15514);
or U19501 (N_19501,N_15580,N_17158);
or U19502 (N_19502,N_17456,N_17210);
nand U19503 (N_19503,N_16187,N_15866);
nor U19504 (N_19504,N_17100,N_17311);
or U19505 (N_19505,N_15304,N_17292);
or U19506 (N_19506,N_16137,N_17161);
or U19507 (N_19507,N_17450,N_15262);
nand U19508 (N_19508,N_17222,N_17157);
nor U19509 (N_19509,N_15177,N_17412);
nor U19510 (N_19510,N_17186,N_15146);
xor U19511 (N_19511,N_15093,N_16030);
nor U19512 (N_19512,N_16349,N_16804);
xnor U19513 (N_19513,N_17064,N_17468);
nand U19514 (N_19514,N_16082,N_17066);
nor U19515 (N_19515,N_16010,N_15031);
nand U19516 (N_19516,N_17092,N_15081);
or U19517 (N_19517,N_16292,N_16614);
nand U19518 (N_19518,N_16272,N_17073);
nor U19519 (N_19519,N_15481,N_17395);
or U19520 (N_19520,N_16065,N_16549);
nor U19521 (N_19521,N_17441,N_15469);
nand U19522 (N_19522,N_16159,N_15886);
nor U19523 (N_19523,N_17448,N_16414);
or U19524 (N_19524,N_16468,N_16830);
xor U19525 (N_19525,N_16548,N_17256);
nor U19526 (N_19526,N_16612,N_17062);
xor U19527 (N_19527,N_15884,N_16956);
nand U19528 (N_19528,N_15710,N_16080);
and U19529 (N_19529,N_16689,N_17480);
and U19530 (N_19530,N_17273,N_16612);
xnor U19531 (N_19531,N_16635,N_15035);
or U19532 (N_19532,N_16496,N_16475);
or U19533 (N_19533,N_15102,N_15654);
xnor U19534 (N_19534,N_15846,N_17406);
nor U19535 (N_19535,N_17097,N_16593);
nor U19536 (N_19536,N_17187,N_16942);
and U19537 (N_19537,N_17470,N_16279);
or U19538 (N_19538,N_16325,N_15570);
nor U19539 (N_19539,N_15448,N_16581);
xor U19540 (N_19540,N_15872,N_15967);
and U19541 (N_19541,N_16589,N_15234);
nor U19542 (N_19542,N_15022,N_15770);
or U19543 (N_19543,N_16717,N_16499);
nand U19544 (N_19544,N_16568,N_17017);
nor U19545 (N_19545,N_15640,N_16614);
nor U19546 (N_19546,N_17024,N_16997);
nand U19547 (N_19547,N_16800,N_16580);
or U19548 (N_19548,N_16151,N_17014);
nor U19549 (N_19549,N_16994,N_17160);
nand U19550 (N_19550,N_15356,N_15327);
or U19551 (N_19551,N_16824,N_17471);
or U19552 (N_19552,N_17241,N_15473);
nor U19553 (N_19553,N_16484,N_17395);
nand U19554 (N_19554,N_16421,N_17357);
nand U19555 (N_19555,N_15254,N_16093);
nor U19556 (N_19556,N_15625,N_15609);
and U19557 (N_19557,N_17399,N_16462);
nor U19558 (N_19558,N_16821,N_16199);
nand U19559 (N_19559,N_17179,N_17416);
xor U19560 (N_19560,N_16303,N_15301);
or U19561 (N_19561,N_16086,N_15938);
or U19562 (N_19562,N_17151,N_15909);
nor U19563 (N_19563,N_17434,N_17151);
or U19564 (N_19564,N_17340,N_16199);
nand U19565 (N_19565,N_16048,N_15924);
nor U19566 (N_19566,N_15912,N_15247);
or U19567 (N_19567,N_16821,N_15076);
nand U19568 (N_19568,N_17222,N_15669);
xor U19569 (N_19569,N_16415,N_15768);
and U19570 (N_19570,N_16461,N_16602);
xnor U19571 (N_19571,N_16852,N_15969);
nor U19572 (N_19572,N_17337,N_17138);
and U19573 (N_19573,N_15115,N_15901);
nor U19574 (N_19574,N_16782,N_15960);
nor U19575 (N_19575,N_15559,N_15507);
nand U19576 (N_19576,N_17326,N_16932);
and U19577 (N_19577,N_17243,N_16173);
and U19578 (N_19578,N_17079,N_15823);
xnor U19579 (N_19579,N_17184,N_17225);
or U19580 (N_19580,N_15863,N_17470);
or U19581 (N_19581,N_16557,N_16643);
or U19582 (N_19582,N_17240,N_16164);
and U19583 (N_19583,N_15173,N_16404);
or U19584 (N_19584,N_16600,N_16238);
nor U19585 (N_19585,N_16997,N_15200);
xnor U19586 (N_19586,N_16253,N_15263);
nor U19587 (N_19587,N_17472,N_16667);
nand U19588 (N_19588,N_15231,N_16740);
xnor U19589 (N_19589,N_16834,N_15425);
xnor U19590 (N_19590,N_15983,N_16412);
xor U19591 (N_19591,N_16739,N_16194);
and U19592 (N_19592,N_16943,N_17162);
nand U19593 (N_19593,N_16307,N_15989);
and U19594 (N_19594,N_16909,N_15375);
or U19595 (N_19595,N_15707,N_17480);
or U19596 (N_19596,N_15682,N_17229);
xor U19597 (N_19597,N_15444,N_15889);
nand U19598 (N_19598,N_16292,N_16457);
xor U19599 (N_19599,N_15154,N_16021);
xnor U19600 (N_19600,N_17412,N_16226);
xor U19601 (N_19601,N_17254,N_17337);
and U19602 (N_19602,N_15210,N_15987);
nor U19603 (N_19603,N_16076,N_15782);
and U19604 (N_19604,N_15312,N_16421);
and U19605 (N_19605,N_16168,N_16083);
and U19606 (N_19606,N_16966,N_17438);
or U19607 (N_19607,N_17296,N_16292);
xor U19608 (N_19608,N_16140,N_17486);
or U19609 (N_19609,N_16045,N_17409);
nor U19610 (N_19610,N_17277,N_15951);
and U19611 (N_19611,N_17368,N_15486);
and U19612 (N_19612,N_16667,N_17278);
xor U19613 (N_19613,N_17484,N_16749);
nor U19614 (N_19614,N_15070,N_15000);
xor U19615 (N_19615,N_15617,N_15118);
xor U19616 (N_19616,N_16733,N_15568);
or U19617 (N_19617,N_15917,N_17305);
xor U19618 (N_19618,N_16983,N_17080);
xnor U19619 (N_19619,N_17462,N_15214);
or U19620 (N_19620,N_16875,N_17320);
nor U19621 (N_19621,N_16866,N_15059);
nor U19622 (N_19622,N_16254,N_15836);
nand U19623 (N_19623,N_17449,N_17090);
and U19624 (N_19624,N_15727,N_16113);
nand U19625 (N_19625,N_17215,N_16894);
and U19626 (N_19626,N_16145,N_15362);
nand U19627 (N_19627,N_15537,N_16495);
xnor U19628 (N_19628,N_17214,N_16764);
nand U19629 (N_19629,N_17243,N_17016);
nor U19630 (N_19630,N_15685,N_17159);
nand U19631 (N_19631,N_17402,N_17150);
and U19632 (N_19632,N_16230,N_15423);
and U19633 (N_19633,N_15553,N_15922);
nor U19634 (N_19634,N_15375,N_16896);
xor U19635 (N_19635,N_15276,N_17211);
nor U19636 (N_19636,N_16548,N_15290);
nor U19637 (N_19637,N_16798,N_16659);
or U19638 (N_19638,N_15964,N_15750);
xor U19639 (N_19639,N_15152,N_16323);
nand U19640 (N_19640,N_17192,N_16350);
or U19641 (N_19641,N_15465,N_16072);
or U19642 (N_19642,N_15054,N_15907);
and U19643 (N_19643,N_15880,N_16665);
and U19644 (N_19644,N_15487,N_16583);
or U19645 (N_19645,N_17212,N_16139);
nand U19646 (N_19646,N_16797,N_16247);
nand U19647 (N_19647,N_16816,N_17184);
and U19648 (N_19648,N_15145,N_17325);
xor U19649 (N_19649,N_15998,N_17328);
and U19650 (N_19650,N_17398,N_17326);
xnor U19651 (N_19651,N_15512,N_16031);
xor U19652 (N_19652,N_15105,N_17420);
nand U19653 (N_19653,N_15677,N_15128);
and U19654 (N_19654,N_15201,N_16248);
nand U19655 (N_19655,N_15135,N_15585);
nand U19656 (N_19656,N_17302,N_16916);
xor U19657 (N_19657,N_15123,N_15225);
xor U19658 (N_19658,N_16396,N_16034);
or U19659 (N_19659,N_17011,N_16120);
xnor U19660 (N_19660,N_17417,N_16995);
nand U19661 (N_19661,N_17121,N_15542);
nor U19662 (N_19662,N_15287,N_16110);
and U19663 (N_19663,N_16864,N_15153);
xnor U19664 (N_19664,N_16073,N_17494);
or U19665 (N_19665,N_15224,N_16231);
nand U19666 (N_19666,N_16074,N_16003);
or U19667 (N_19667,N_16979,N_15885);
and U19668 (N_19668,N_16200,N_15636);
nand U19669 (N_19669,N_15997,N_17474);
or U19670 (N_19670,N_16789,N_15698);
xor U19671 (N_19671,N_16328,N_17449);
xor U19672 (N_19672,N_17431,N_16780);
or U19673 (N_19673,N_15129,N_16890);
nor U19674 (N_19674,N_15319,N_16491);
or U19675 (N_19675,N_15706,N_15174);
and U19676 (N_19676,N_16876,N_15954);
or U19677 (N_19677,N_15748,N_17163);
nand U19678 (N_19678,N_16013,N_15649);
xnor U19679 (N_19679,N_15746,N_16679);
and U19680 (N_19680,N_15568,N_15552);
or U19681 (N_19681,N_17227,N_17021);
nor U19682 (N_19682,N_15593,N_15612);
xor U19683 (N_19683,N_15969,N_15268);
xnor U19684 (N_19684,N_15223,N_17448);
nand U19685 (N_19685,N_16434,N_15344);
nand U19686 (N_19686,N_15709,N_16561);
nor U19687 (N_19687,N_16993,N_16933);
nor U19688 (N_19688,N_16108,N_16196);
or U19689 (N_19689,N_16760,N_17167);
xor U19690 (N_19690,N_15463,N_17421);
xnor U19691 (N_19691,N_15906,N_15358);
nand U19692 (N_19692,N_16852,N_16465);
or U19693 (N_19693,N_15656,N_16455);
xor U19694 (N_19694,N_16987,N_16143);
nand U19695 (N_19695,N_17117,N_15658);
xnor U19696 (N_19696,N_15976,N_15466);
nor U19697 (N_19697,N_15093,N_15596);
xnor U19698 (N_19698,N_15904,N_17268);
nor U19699 (N_19699,N_15289,N_15113);
nand U19700 (N_19700,N_15825,N_16246);
nand U19701 (N_19701,N_16334,N_15498);
xnor U19702 (N_19702,N_15610,N_15663);
and U19703 (N_19703,N_15197,N_15003);
xnor U19704 (N_19704,N_15698,N_15211);
xnor U19705 (N_19705,N_15920,N_16811);
nand U19706 (N_19706,N_17243,N_15085);
nand U19707 (N_19707,N_15509,N_15413);
or U19708 (N_19708,N_15588,N_16506);
nand U19709 (N_19709,N_15819,N_16369);
nor U19710 (N_19710,N_16276,N_16174);
nand U19711 (N_19711,N_15220,N_17088);
and U19712 (N_19712,N_15356,N_17412);
xnor U19713 (N_19713,N_15157,N_15022);
and U19714 (N_19714,N_15084,N_16882);
nor U19715 (N_19715,N_15121,N_16323);
nand U19716 (N_19716,N_16788,N_17059);
or U19717 (N_19717,N_15284,N_17393);
or U19718 (N_19718,N_15301,N_16380);
or U19719 (N_19719,N_15589,N_17191);
nor U19720 (N_19720,N_15332,N_16959);
xnor U19721 (N_19721,N_15317,N_17387);
or U19722 (N_19722,N_16747,N_15708);
nand U19723 (N_19723,N_15357,N_17075);
and U19724 (N_19724,N_17118,N_15428);
nor U19725 (N_19725,N_15335,N_16142);
xor U19726 (N_19726,N_17266,N_17486);
or U19727 (N_19727,N_15334,N_15099);
or U19728 (N_19728,N_15555,N_17128);
nor U19729 (N_19729,N_16565,N_16175);
and U19730 (N_19730,N_16469,N_16678);
or U19731 (N_19731,N_15725,N_16446);
nor U19732 (N_19732,N_15012,N_15208);
xor U19733 (N_19733,N_15812,N_16008);
nand U19734 (N_19734,N_16869,N_16485);
and U19735 (N_19735,N_16559,N_16916);
nand U19736 (N_19736,N_16226,N_15405);
nand U19737 (N_19737,N_16593,N_15810);
nor U19738 (N_19738,N_16829,N_15137);
and U19739 (N_19739,N_15364,N_17184);
nor U19740 (N_19740,N_15269,N_16070);
nor U19741 (N_19741,N_17435,N_15658);
nor U19742 (N_19742,N_16466,N_16408);
or U19743 (N_19743,N_17115,N_16732);
or U19744 (N_19744,N_16621,N_16434);
xor U19745 (N_19745,N_15381,N_16351);
and U19746 (N_19746,N_16785,N_15904);
nand U19747 (N_19747,N_16679,N_16175);
and U19748 (N_19748,N_16632,N_17370);
xor U19749 (N_19749,N_15823,N_15909);
and U19750 (N_19750,N_17467,N_16940);
nand U19751 (N_19751,N_16418,N_15904);
xor U19752 (N_19752,N_17243,N_16751);
nand U19753 (N_19753,N_16975,N_15846);
and U19754 (N_19754,N_17371,N_17004);
nand U19755 (N_19755,N_16628,N_17002);
and U19756 (N_19756,N_16006,N_16855);
nand U19757 (N_19757,N_16291,N_15472);
or U19758 (N_19758,N_15179,N_15336);
xnor U19759 (N_19759,N_15114,N_16218);
and U19760 (N_19760,N_16197,N_17107);
xor U19761 (N_19761,N_16786,N_17381);
nor U19762 (N_19762,N_16414,N_15512);
nand U19763 (N_19763,N_16939,N_17355);
or U19764 (N_19764,N_16023,N_15077);
xnor U19765 (N_19765,N_16884,N_17140);
or U19766 (N_19766,N_15927,N_16187);
xor U19767 (N_19767,N_16977,N_16631);
nand U19768 (N_19768,N_15837,N_16920);
and U19769 (N_19769,N_15290,N_17464);
xnor U19770 (N_19770,N_15901,N_17415);
and U19771 (N_19771,N_15124,N_15336);
nand U19772 (N_19772,N_15483,N_15942);
and U19773 (N_19773,N_17001,N_17342);
nand U19774 (N_19774,N_15911,N_16078);
or U19775 (N_19775,N_16987,N_16471);
nand U19776 (N_19776,N_15964,N_16041);
nand U19777 (N_19777,N_16519,N_15200);
or U19778 (N_19778,N_15779,N_17478);
or U19779 (N_19779,N_15882,N_16651);
or U19780 (N_19780,N_16420,N_17415);
nor U19781 (N_19781,N_17280,N_15158);
and U19782 (N_19782,N_15427,N_15692);
nand U19783 (N_19783,N_16489,N_16273);
and U19784 (N_19784,N_16993,N_16629);
or U19785 (N_19785,N_16465,N_16866);
or U19786 (N_19786,N_16656,N_16659);
nand U19787 (N_19787,N_15941,N_16964);
nand U19788 (N_19788,N_16388,N_15972);
or U19789 (N_19789,N_16961,N_17374);
nand U19790 (N_19790,N_16698,N_15044);
and U19791 (N_19791,N_16647,N_15547);
nand U19792 (N_19792,N_16203,N_15716);
xnor U19793 (N_19793,N_16864,N_17421);
or U19794 (N_19794,N_16631,N_16865);
xor U19795 (N_19795,N_17482,N_15334);
and U19796 (N_19796,N_15835,N_17072);
xnor U19797 (N_19797,N_15283,N_15674);
and U19798 (N_19798,N_16085,N_15618);
nand U19799 (N_19799,N_15228,N_15575);
and U19800 (N_19800,N_16016,N_17012);
nand U19801 (N_19801,N_15870,N_17291);
or U19802 (N_19802,N_16305,N_17466);
nand U19803 (N_19803,N_16670,N_16920);
or U19804 (N_19804,N_17061,N_15763);
and U19805 (N_19805,N_16264,N_17067);
nand U19806 (N_19806,N_15549,N_16482);
xor U19807 (N_19807,N_15843,N_17383);
xnor U19808 (N_19808,N_17021,N_16415);
nor U19809 (N_19809,N_16306,N_16235);
nor U19810 (N_19810,N_16385,N_16943);
xor U19811 (N_19811,N_15562,N_15848);
nand U19812 (N_19812,N_16143,N_15908);
xnor U19813 (N_19813,N_16651,N_17300);
xnor U19814 (N_19814,N_17169,N_16436);
xnor U19815 (N_19815,N_15786,N_15178);
xor U19816 (N_19816,N_16953,N_16850);
nor U19817 (N_19817,N_16548,N_15324);
and U19818 (N_19818,N_17273,N_16265);
nand U19819 (N_19819,N_16034,N_15197);
or U19820 (N_19820,N_15717,N_15551);
and U19821 (N_19821,N_15071,N_15772);
nand U19822 (N_19822,N_15686,N_15603);
and U19823 (N_19823,N_16741,N_16899);
and U19824 (N_19824,N_17237,N_17157);
or U19825 (N_19825,N_16297,N_15349);
or U19826 (N_19826,N_16741,N_17286);
nor U19827 (N_19827,N_15213,N_16405);
and U19828 (N_19828,N_16926,N_15268);
xor U19829 (N_19829,N_16791,N_16982);
or U19830 (N_19830,N_15595,N_16587);
nor U19831 (N_19831,N_15756,N_17228);
nand U19832 (N_19832,N_16718,N_15244);
or U19833 (N_19833,N_15044,N_16592);
or U19834 (N_19834,N_16088,N_16796);
nor U19835 (N_19835,N_17395,N_16187);
and U19836 (N_19836,N_15429,N_17497);
nand U19837 (N_19837,N_15165,N_15555);
xnor U19838 (N_19838,N_17497,N_15057);
or U19839 (N_19839,N_17044,N_17066);
nor U19840 (N_19840,N_16902,N_15371);
nand U19841 (N_19841,N_16752,N_17274);
nand U19842 (N_19842,N_15230,N_16318);
or U19843 (N_19843,N_16180,N_16553);
and U19844 (N_19844,N_16662,N_16351);
or U19845 (N_19845,N_17277,N_17331);
nor U19846 (N_19846,N_17392,N_16471);
nand U19847 (N_19847,N_15592,N_17417);
and U19848 (N_19848,N_16449,N_16126);
xor U19849 (N_19849,N_16527,N_16902);
and U19850 (N_19850,N_16263,N_16951);
and U19851 (N_19851,N_15183,N_15917);
and U19852 (N_19852,N_17319,N_16141);
nand U19853 (N_19853,N_15696,N_16239);
and U19854 (N_19854,N_15064,N_17339);
or U19855 (N_19855,N_16410,N_16754);
nor U19856 (N_19856,N_17124,N_15404);
and U19857 (N_19857,N_17461,N_15462);
or U19858 (N_19858,N_15862,N_17347);
and U19859 (N_19859,N_15785,N_17138);
or U19860 (N_19860,N_15230,N_15719);
nand U19861 (N_19861,N_16255,N_16148);
nand U19862 (N_19862,N_17142,N_17077);
or U19863 (N_19863,N_15824,N_16972);
nor U19864 (N_19864,N_16975,N_16947);
nor U19865 (N_19865,N_16624,N_17409);
and U19866 (N_19866,N_15771,N_15579);
or U19867 (N_19867,N_15331,N_15285);
or U19868 (N_19868,N_17451,N_16540);
xnor U19869 (N_19869,N_16475,N_17438);
xor U19870 (N_19870,N_16087,N_17401);
nand U19871 (N_19871,N_16921,N_15930);
or U19872 (N_19872,N_15801,N_16214);
and U19873 (N_19873,N_16930,N_15463);
xnor U19874 (N_19874,N_16466,N_16727);
and U19875 (N_19875,N_16940,N_15247);
nand U19876 (N_19876,N_15114,N_15068);
or U19877 (N_19877,N_15519,N_15933);
or U19878 (N_19878,N_17112,N_15802);
nand U19879 (N_19879,N_16517,N_16071);
nand U19880 (N_19880,N_17309,N_15461);
and U19881 (N_19881,N_15986,N_16056);
and U19882 (N_19882,N_16542,N_17385);
or U19883 (N_19883,N_16324,N_17230);
or U19884 (N_19884,N_17039,N_15834);
nor U19885 (N_19885,N_15907,N_15871);
or U19886 (N_19886,N_17364,N_17116);
xor U19887 (N_19887,N_16714,N_16715);
xnor U19888 (N_19888,N_17292,N_15412);
or U19889 (N_19889,N_17073,N_15983);
and U19890 (N_19890,N_15422,N_17241);
nand U19891 (N_19891,N_16010,N_16343);
nand U19892 (N_19892,N_16962,N_17151);
nand U19893 (N_19893,N_16339,N_15288);
and U19894 (N_19894,N_17326,N_15874);
nand U19895 (N_19895,N_16709,N_15056);
or U19896 (N_19896,N_17491,N_15865);
or U19897 (N_19897,N_16296,N_15272);
nand U19898 (N_19898,N_15364,N_17224);
and U19899 (N_19899,N_17313,N_16186);
nor U19900 (N_19900,N_15387,N_15354);
and U19901 (N_19901,N_15982,N_16176);
nand U19902 (N_19902,N_15257,N_17000);
or U19903 (N_19903,N_15678,N_15127);
xor U19904 (N_19904,N_17097,N_16722);
nor U19905 (N_19905,N_15491,N_16195);
or U19906 (N_19906,N_15082,N_15472);
and U19907 (N_19907,N_17235,N_17285);
and U19908 (N_19908,N_15788,N_15283);
and U19909 (N_19909,N_15160,N_17088);
and U19910 (N_19910,N_15463,N_17479);
or U19911 (N_19911,N_16815,N_16887);
or U19912 (N_19912,N_16128,N_16458);
xnor U19913 (N_19913,N_15138,N_15685);
or U19914 (N_19914,N_15449,N_15396);
and U19915 (N_19915,N_16484,N_16407);
xor U19916 (N_19916,N_16948,N_16830);
xor U19917 (N_19917,N_15691,N_17095);
xor U19918 (N_19918,N_17280,N_16166);
xnor U19919 (N_19919,N_15334,N_16579);
and U19920 (N_19920,N_15219,N_16615);
nand U19921 (N_19921,N_15598,N_16798);
xnor U19922 (N_19922,N_17436,N_16496);
nand U19923 (N_19923,N_15717,N_16477);
nor U19924 (N_19924,N_15136,N_16492);
nand U19925 (N_19925,N_17403,N_16052);
nand U19926 (N_19926,N_16030,N_17146);
and U19927 (N_19927,N_15151,N_17419);
nor U19928 (N_19928,N_15896,N_15565);
nor U19929 (N_19929,N_16603,N_17488);
and U19930 (N_19930,N_16611,N_15731);
and U19931 (N_19931,N_15030,N_16832);
and U19932 (N_19932,N_17460,N_17224);
nor U19933 (N_19933,N_15156,N_15050);
xor U19934 (N_19934,N_16353,N_15378);
nand U19935 (N_19935,N_15670,N_15760);
nand U19936 (N_19936,N_15889,N_15970);
nor U19937 (N_19937,N_16232,N_17438);
nor U19938 (N_19938,N_15274,N_15397);
and U19939 (N_19939,N_16948,N_17484);
and U19940 (N_19940,N_15813,N_15499);
nand U19941 (N_19941,N_15039,N_17436);
xnor U19942 (N_19942,N_16762,N_16531);
nand U19943 (N_19943,N_17078,N_15447);
xnor U19944 (N_19944,N_15410,N_16529);
xnor U19945 (N_19945,N_16739,N_16742);
and U19946 (N_19946,N_17335,N_17316);
or U19947 (N_19947,N_15620,N_17072);
xor U19948 (N_19948,N_15942,N_15381);
xnor U19949 (N_19949,N_15753,N_16484);
nor U19950 (N_19950,N_15673,N_17454);
nand U19951 (N_19951,N_15285,N_16321);
nor U19952 (N_19952,N_16336,N_15724);
xnor U19953 (N_19953,N_16369,N_16940);
nor U19954 (N_19954,N_15702,N_16413);
nand U19955 (N_19955,N_16226,N_15610);
and U19956 (N_19956,N_17368,N_17144);
or U19957 (N_19957,N_15919,N_15753);
nor U19958 (N_19958,N_15187,N_15908);
nor U19959 (N_19959,N_16935,N_16536);
nor U19960 (N_19960,N_15846,N_17139);
and U19961 (N_19961,N_16116,N_16980);
or U19962 (N_19962,N_15246,N_15918);
or U19963 (N_19963,N_15020,N_15051);
and U19964 (N_19964,N_16767,N_16281);
and U19965 (N_19965,N_15038,N_15283);
or U19966 (N_19966,N_15542,N_16160);
and U19967 (N_19967,N_16462,N_16289);
nor U19968 (N_19968,N_17453,N_15174);
and U19969 (N_19969,N_15449,N_16594);
xor U19970 (N_19970,N_16283,N_15345);
nor U19971 (N_19971,N_16901,N_15693);
nor U19972 (N_19972,N_15023,N_16885);
and U19973 (N_19973,N_17317,N_16798);
nor U19974 (N_19974,N_16046,N_16473);
xnor U19975 (N_19975,N_16945,N_16498);
nor U19976 (N_19976,N_17093,N_15795);
or U19977 (N_19977,N_16517,N_16167);
xnor U19978 (N_19978,N_15003,N_16572);
and U19979 (N_19979,N_15427,N_15931);
nor U19980 (N_19980,N_16363,N_15795);
or U19981 (N_19981,N_15532,N_16389);
xnor U19982 (N_19982,N_16545,N_15433);
nand U19983 (N_19983,N_16125,N_15621);
nand U19984 (N_19984,N_16011,N_16286);
and U19985 (N_19985,N_16304,N_15287);
nand U19986 (N_19986,N_15913,N_16379);
nand U19987 (N_19987,N_16552,N_17379);
and U19988 (N_19988,N_16877,N_16850);
nand U19989 (N_19989,N_17298,N_15587);
nor U19990 (N_19990,N_15330,N_15815);
nand U19991 (N_19991,N_17361,N_15622);
and U19992 (N_19992,N_16658,N_17246);
xnor U19993 (N_19993,N_15047,N_15628);
nand U19994 (N_19994,N_15824,N_17380);
nand U19995 (N_19995,N_15712,N_15972);
nand U19996 (N_19996,N_16214,N_16712);
and U19997 (N_19997,N_16272,N_16087);
xnor U19998 (N_19998,N_15648,N_15868);
nand U19999 (N_19999,N_16965,N_16964);
and U20000 (N_20000,N_19542,N_18756);
nor U20001 (N_20001,N_18368,N_17550);
and U20002 (N_20002,N_19582,N_18636);
and U20003 (N_20003,N_19404,N_19368);
xnor U20004 (N_20004,N_17542,N_18408);
nand U20005 (N_20005,N_17750,N_19362);
and U20006 (N_20006,N_19793,N_19147);
nand U20007 (N_20007,N_18290,N_17844);
nor U20008 (N_20008,N_19451,N_19191);
nor U20009 (N_20009,N_19099,N_19736);
nor U20010 (N_20010,N_19781,N_19774);
or U20011 (N_20011,N_18224,N_19279);
or U20012 (N_20012,N_19919,N_18442);
nor U20013 (N_20013,N_19879,N_19361);
nor U20014 (N_20014,N_19274,N_19051);
and U20015 (N_20015,N_17704,N_19121);
xnor U20016 (N_20016,N_18245,N_18816);
and U20017 (N_20017,N_18903,N_17596);
xnor U20018 (N_20018,N_18863,N_18455);
xnor U20019 (N_20019,N_19253,N_18026);
xnor U20020 (N_20020,N_19620,N_18591);
or U20021 (N_20021,N_17610,N_18631);
nor U20022 (N_20022,N_17838,N_17567);
or U20023 (N_20023,N_19876,N_17973);
or U20024 (N_20024,N_19042,N_19011);
and U20025 (N_20025,N_18091,N_18694);
nor U20026 (N_20026,N_18189,N_19201);
and U20027 (N_20027,N_18963,N_18471);
or U20028 (N_20028,N_17728,N_17963);
nand U20029 (N_20029,N_18074,N_18649);
xnor U20030 (N_20030,N_19431,N_19033);
or U20031 (N_20031,N_19839,N_18492);
or U20032 (N_20032,N_18698,N_19588);
nand U20033 (N_20033,N_18771,N_18937);
and U20034 (N_20034,N_18036,N_19997);
or U20035 (N_20035,N_19733,N_17560);
nor U20036 (N_20036,N_17531,N_19570);
nand U20037 (N_20037,N_19089,N_19882);
xor U20038 (N_20038,N_18302,N_17732);
nand U20039 (N_20039,N_19034,N_18068);
xor U20040 (N_20040,N_19081,N_19382);
xor U20041 (N_20041,N_19547,N_17516);
or U20042 (N_20042,N_18174,N_18933);
nor U20043 (N_20043,N_18745,N_19463);
or U20044 (N_20044,N_19596,N_18237);
nor U20045 (N_20045,N_18219,N_17926);
nand U20046 (N_20046,N_18128,N_19068);
xnor U20047 (N_20047,N_19900,N_19385);
xnor U20048 (N_20048,N_19727,N_19327);
nand U20049 (N_20049,N_18549,N_17943);
or U20050 (N_20050,N_19895,N_19260);
or U20051 (N_20051,N_18513,N_18375);
nand U20052 (N_20052,N_18864,N_18055);
xor U20053 (N_20053,N_17678,N_18930);
nand U20054 (N_20054,N_18583,N_17912);
or U20055 (N_20055,N_18281,N_18612);
xnor U20056 (N_20056,N_18314,N_19521);
and U20057 (N_20057,N_19240,N_18126);
and U20058 (N_20058,N_17514,N_19067);
xor U20059 (N_20059,N_19710,N_17918);
nor U20060 (N_20060,N_18880,N_18618);
or U20061 (N_20061,N_17636,N_19120);
or U20062 (N_20062,N_18094,N_18845);
and U20063 (N_20063,N_19851,N_19869);
or U20064 (N_20064,N_18283,N_19835);
nor U20065 (N_20065,N_18517,N_19225);
nand U20066 (N_20066,N_17687,N_17934);
or U20067 (N_20067,N_19992,N_18855);
and U20068 (N_20068,N_17548,N_19052);
xor U20069 (N_20069,N_19455,N_18954);
or U20070 (N_20070,N_19910,N_19885);
nor U20071 (N_20071,N_19566,N_18508);
xor U20072 (N_20072,N_18156,N_18432);
and U20073 (N_20073,N_17651,N_17673);
nor U20074 (N_20074,N_18522,N_17999);
xnor U20075 (N_20075,N_18383,N_18087);
xor U20076 (N_20076,N_18897,N_19234);
nor U20077 (N_20077,N_19724,N_18066);
xor U20078 (N_20078,N_18892,N_18460);
xor U20079 (N_20079,N_17527,N_19574);
or U20080 (N_20080,N_19152,N_18944);
and U20081 (N_20081,N_17522,N_18685);
nand U20082 (N_20082,N_18960,N_17798);
nor U20083 (N_20083,N_19071,N_17683);
nand U20084 (N_20084,N_19397,N_18321);
and U20085 (N_20085,N_17925,N_18208);
nand U20086 (N_20086,N_18758,N_17776);
xor U20087 (N_20087,N_18425,N_19432);
and U20088 (N_20088,N_18740,N_18424);
xor U20089 (N_20089,N_17581,N_19217);
and U20090 (N_20090,N_19079,N_18790);
and U20091 (N_20091,N_19353,N_17536);
nor U20092 (N_20092,N_17994,N_19140);
and U20093 (N_20093,N_19658,N_19514);
or U20094 (N_20094,N_19183,N_19539);
and U20095 (N_20095,N_19677,N_17786);
nand U20096 (N_20096,N_19290,N_18085);
nor U20097 (N_20097,N_19129,N_17731);
xnor U20098 (N_20098,N_18057,N_17974);
or U20099 (N_20099,N_19532,N_18556);
nor U20100 (N_20100,N_19780,N_19429);
or U20101 (N_20101,N_19436,N_18239);
and U20102 (N_20102,N_19255,N_18762);
nor U20103 (N_20103,N_18768,N_19370);
and U20104 (N_20104,N_19728,N_19916);
xnor U20105 (N_20105,N_18078,N_17637);
nor U20106 (N_20106,N_19921,N_19784);
xor U20107 (N_20107,N_18754,N_19012);
or U20108 (N_20108,N_17722,N_18297);
nand U20109 (N_20109,N_18214,N_18354);
nand U20110 (N_20110,N_18121,N_19203);
xnor U20111 (N_20111,N_19095,N_18682);
or U20112 (N_20112,N_19014,N_17590);
nor U20113 (N_20113,N_18491,N_19466);
nand U20114 (N_20114,N_18988,N_18201);
and U20115 (N_20115,N_18351,N_17743);
or U20116 (N_20116,N_18435,N_18728);
or U20117 (N_20117,N_17952,N_19286);
and U20118 (N_20118,N_18238,N_19096);
or U20119 (N_20119,N_17717,N_17933);
nand U20120 (N_20120,N_18700,N_18851);
xor U20121 (N_20121,N_18914,N_19942);
nand U20122 (N_20122,N_19703,N_18114);
nor U20123 (N_20123,N_19263,N_19220);
or U20124 (N_20124,N_17625,N_19557);
xnor U20125 (N_20125,N_17710,N_18994);
xor U20126 (N_20126,N_18441,N_17945);
or U20127 (N_20127,N_19280,N_19980);
nand U20128 (N_20128,N_17808,N_18382);
nor U20129 (N_20129,N_17919,N_17521);
and U20130 (N_20130,N_19770,N_17816);
and U20131 (N_20131,N_19896,N_18941);
nor U20132 (N_20132,N_17902,N_18462);
and U20133 (N_20133,N_18360,N_18160);
nand U20134 (N_20134,N_19157,N_19573);
or U20135 (N_20135,N_17761,N_19714);
or U20136 (N_20136,N_18456,N_18499);
nand U20137 (N_20137,N_18961,N_19330);
nor U20138 (N_20138,N_19039,N_18002);
and U20139 (N_20139,N_17889,N_18269);
nand U20140 (N_20140,N_19639,N_18362);
nand U20141 (N_20141,N_19338,N_19863);
and U20142 (N_20142,N_18555,N_19927);
nand U20143 (N_20143,N_19510,N_18440);
and U20144 (N_20144,N_18964,N_19126);
nand U20145 (N_20145,N_18610,N_19438);
and U20146 (N_20146,N_18211,N_18379);
and U20147 (N_20147,N_18877,N_18343);
xor U20148 (N_20148,N_19968,N_18466);
nor U20149 (N_20149,N_19858,N_18277);
or U20150 (N_20150,N_18785,N_19301);
nand U20151 (N_20151,N_18086,N_19426);
nor U20152 (N_20152,N_17815,N_18388);
and U20153 (N_20153,N_17855,N_17615);
or U20154 (N_20154,N_18688,N_19139);
nor U20155 (N_20155,N_17895,N_19555);
nand U20156 (N_20156,N_18065,N_18274);
and U20157 (N_20157,N_18474,N_18100);
xor U20158 (N_20158,N_18609,N_19753);
or U20159 (N_20159,N_18199,N_19453);
nand U20160 (N_20160,N_17972,N_18198);
and U20161 (N_20161,N_19966,N_19090);
xor U20162 (N_20162,N_17837,N_19424);
and U20163 (N_20163,N_19956,N_18380);
nor U20164 (N_20164,N_18257,N_19124);
xor U20165 (N_20165,N_18828,N_19227);
or U20166 (N_20166,N_18447,N_19377);
and U20167 (N_20167,N_18686,N_17553);
nand U20168 (N_20168,N_17692,N_18893);
xnor U20169 (N_20169,N_17505,N_19141);
or U20170 (N_20170,N_18465,N_17783);
nor U20171 (N_20171,N_18955,N_17696);
and U20172 (N_20172,N_18966,N_19374);
and U20173 (N_20173,N_18817,N_19782);
xor U20174 (N_20174,N_19976,N_17916);
xnor U20175 (N_20175,N_19146,N_18521);
and U20176 (N_20176,N_19036,N_19343);
and U20177 (N_20177,N_18376,N_18545);
or U20178 (N_20178,N_18904,N_18401);
or U20179 (N_20179,N_19899,N_17624);
xnor U20180 (N_20180,N_18072,N_19023);
and U20181 (N_20181,N_19518,N_17813);
or U20182 (N_20182,N_18047,N_19949);
xor U20183 (N_20183,N_18727,N_18601);
nand U20184 (N_20184,N_17688,N_19421);
nor U20185 (N_20185,N_18755,N_19437);
nand U20186 (N_20186,N_19294,N_18405);
or U20187 (N_20187,N_18919,N_19776);
or U20188 (N_20188,N_17579,N_18217);
and U20189 (N_20189,N_18143,N_18037);
and U20190 (N_20190,N_19307,N_19541);
and U20191 (N_20191,N_17839,N_18912);
nand U20192 (N_20192,N_19066,N_19577);
nor U20193 (N_20193,N_18546,N_19722);
nor U20194 (N_20194,N_18421,N_19845);
nand U20195 (N_20195,N_19304,N_17773);
nor U20196 (N_20196,N_17795,N_18137);
or U20197 (N_20197,N_18623,N_18596);
nand U20198 (N_20198,N_18789,N_18588);
nand U20199 (N_20199,N_19475,N_18722);
xor U20200 (N_20200,N_19419,N_19638);
and U20201 (N_20201,N_19193,N_17616);
nand U20202 (N_20202,N_19901,N_19352);
nand U20203 (N_20203,N_19258,N_18574);
or U20204 (N_20204,N_17980,N_19777);
nand U20205 (N_20205,N_19551,N_19093);
nor U20206 (N_20206,N_18018,N_18357);
or U20207 (N_20207,N_18475,N_18769);
xnor U20208 (N_20208,N_17599,N_18080);
xor U20209 (N_20209,N_18626,N_18258);
and U20210 (N_20210,N_17532,N_17903);
nand U20211 (N_20211,N_19055,N_18822);
nor U20212 (N_20212,N_17981,N_19686);
nand U20213 (N_20213,N_18720,N_18561);
or U20214 (N_20214,N_18389,N_17823);
nand U20215 (N_20215,N_17629,N_18586);
and U20216 (N_20216,N_19932,N_17971);
and U20217 (N_20217,N_18320,N_18662);
and U20218 (N_20218,N_19190,N_19534);
nand U20219 (N_20219,N_18957,N_17924);
xnor U20220 (N_20220,N_19192,N_17819);
and U20221 (N_20221,N_18878,N_19392);
or U20222 (N_20222,N_19685,N_18641);
or U20223 (N_20223,N_19484,N_18613);
or U20224 (N_20224,N_19801,N_17881);
nor U20225 (N_20225,N_19000,N_18625);
nor U20226 (N_20226,N_18325,N_19237);
xor U20227 (N_20227,N_18597,N_19684);
nor U20228 (N_20228,N_19349,N_19855);
and U20229 (N_20229,N_18691,N_18542);
nand U20230 (N_20230,N_18312,N_19402);
nand U20231 (N_20231,N_19856,N_19344);
nor U20232 (N_20232,N_19533,N_19877);
and U20233 (N_20233,N_17698,N_19127);
xor U20234 (N_20234,N_17591,N_19786);
xnor U20235 (N_20235,N_17998,N_18176);
nor U20236 (N_20236,N_19970,N_18235);
nand U20237 (N_20237,N_19222,N_18882);
or U20238 (N_20238,N_19676,N_18655);
or U20239 (N_20239,N_18001,N_19365);
or U20240 (N_20240,N_19982,N_18182);
nand U20241 (N_20241,N_19729,N_18154);
nor U20242 (N_20242,N_18890,N_18835);
and U20243 (N_20243,N_18520,N_17621);
xnor U20244 (N_20244,N_18348,N_17622);
nor U20245 (N_20245,N_18825,N_19180);
nor U20246 (N_20246,N_18384,N_18180);
nand U20247 (N_20247,N_19358,N_18945);
and U20248 (N_20248,N_18997,N_19866);
and U20249 (N_20249,N_19825,N_18734);
or U20250 (N_20250,N_19669,N_18593);
or U20251 (N_20251,N_17569,N_18426);
nor U20252 (N_20252,N_19559,N_19242);
nand U20253 (N_20253,N_19312,N_19578);
or U20254 (N_20254,N_19946,N_19792);
and U20255 (N_20255,N_19202,N_18118);
nor U20256 (N_20256,N_19238,N_19423);
nor U20257 (N_20257,N_17932,N_19730);
nand U20258 (N_20258,N_18285,N_18342);
and U20259 (N_20259,N_19491,N_19446);
and U20260 (N_20260,N_18512,N_19527);
xor U20261 (N_20261,N_19704,N_18661);
xor U20262 (N_20262,N_18515,N_18854);
and U20263 (N_20263,N_17899,N_18744);
and U20264 (N_20264,N_17570,N_18876);
or U20265 (N_20265,N_18363,N_18053);
nand U20266 (N_20266,N_17949,N_19218);
xnor U20267 (N_20267,N_19687,N_18753);
and U20268 (N_20268,N_18995,N_18949);
nand U20269 (N_20269,N_18319,N_19028);
nand U20270 (N_20270,N_19944,N_19091);
and U20271 (N_20271,N_18735,N_18242);
nand U20272 (N_20272,N_18853,N_19644);
or U20273 (N_20273,N_18659,N_19673);
nor U20274 (N_20274,N_17675,N_18965);
xnor U20275 (N_20275,N_19892,N_17957);
or U20276 (N_20276,N_19176,N_19528);
and U20277 (N_20277,N_19371,N_17807);
or U20278 (N_20278,N_19049,N_19509);
nand U20279 (N_20279,N_18496,N_19967);
xnor U20280 (N_20280,N_18717,N_18538);
xor U20281 (N_20281,N_19571,N_18092);
xor U20282 (N_20282,N_19412,N_19341);
nand U20283 (N_20283,N_19390,N_18948);
or U20284 (N_20284,N_18399,N_19590);
nand U20285 (N_20285,N_18602,N_18070);
nor U20286 (N_20286,N_17526,N_18478);
and U20287 (N_20287,N_19077,N_19305);
nand U20288 (N_20288,N_18102,N_17879);
xor U20289 (N_20289,N_17524,N_18397);
and U20290 (N_20290,N_19300,N_18185);
nand U20291 (N_20291,N_19647,N_17628);
xnor U20292 (N_20292,N_18974,N_19803);
nor U20293 (N_20293,N_18450,N_18493);
xnor U20294 (N_20294,N_18887,N_17996);
and U20295 (N_20295,N_18811,N_18200);
xnor U20296 (N_20296,N_19470,N_19293);
xor U20297 (N_20297,N_18009,N_19958);
nor U20298 (N_20298,N_17512,N_17735);
nand U20299 (N_20299,N_19670,N_19756);
nand U20300 (N_20300,N_19779,N_18192);
or U20301 (N_20301,N_18259,N_19883);
xor U20302 (N_20302,N_18934,N_18850);
and U20303 (N_20303,N_19619,N_17936);
xor U20304 (N_20304,N_19132,N_18136);
and U20305 (N_20305,N_18742,N_18016);
and U20306 (N_20306,N_17541,N_19741);
nor U20307 (N_20307,N_18540,N_18888);
or U20308 (N_20308,N_19478,N_19372);
nor U20309 (N_20309,N_17875,N_18579);
xor U20310 (N_20310,N_17860,N_19654);
xnor U20311 (N_20311,N_19032,N_17680);
nand U20312 (N_20312,N_19134,N_19481);
or U20313 (N_20313,N_19544,N_17968);
xnor U20314 (N_20314,N_18548,N_18204);
and U20315 (N_20315,N_18746,N_19824);
or U20316 (N_20316,N_18067,N_19080);
nand U20317 (N_20317,N_19785,N_18227);
or U20318 (N_20318,N_18869,N_19233);
xor U20319 (N_20319,N_19600,N_19272);
xor U20320 (N_20320,N_19973,N_19752);
or U20321 (N_20321,N_19076,N_18606);
or U20322 (N_20322,N_19734,N_19289);
nor U20323 (N_20323,N_17915,N_19232);
or U20324 (N_20324,N_19430,N_19322);
nor U20325 (N_20325,N_18300,N_17812);
or U20326 (N_20326,N_19447,N_19065);
nand U20327 (N_20327,N_18260,N_18761);
xor U20328 (N_20328,N_17827,N_19007);
and U20329 (N_20329,N_18594,N_18633);
nand U20330 (N_20330,N_18537,N_19920);
and U20331 (N_20331,N_17755,N_19306);
nor U20332 (N_20332,N_19018,N_18923);
nor U20333 (N_20333,N_18256,N_18999);
or U20334 (N_20334,N_19831,N_18205);
or U20335 (N_20335,N_17766,N_19884);
nor U20336 (N_20336,N_19611,N_18833);
nor U20337 (N_20337,N_18031,N_19584);
and U20338 (N_20338,N_18138,N_18461);
or U20339 (N_20339,N_18063,N_19764);
or U20340 (N_20340,N_18837,N_19961);
xor U20341 (N_20341,N_17878,N_17749);
nand U20342 (N_20342,N_19410,N_18983);
nand U20343 (N_20343,N_18842,N_18341);
or U20344 (N_20344,N_19864,N_19084);
nand U20345 (N_20345,N_17894,N_18406);
nor U20346 (N_20346,N_18434,N_18041);
and U20347 (N_20347,N_17583,N_18826);
and U20348 (N_20348,N_17605,N_18946);
nand U20349 (N_20349,N_17632,N_18939);
nand U20350 (N_20350,N_19044,N_19550);
or U20351 (N_20351,N_18386,N_18696);
or U20352 (N_20352,N_18721,N_17898);
and U20353 (N_20353,N_17565,N_18551);
nor U20354 (N_20354,N_19746,N_19271);
nand U20355 (N_20355,N_19675,N_19612);
xor U20356 (N_20356,N_18781,N_17908);
nor U20357 (N_20357,N_18374,N_19716);
or U20358 (N_20358,N_17537,N_19262);
nand U20359 (N_20359,N_18364,N_18096);
or U20360 (N_20360,N_19137,N_17790);
or U20361 (N_20361,N_18190,N_18577);
nand U20362 (N_20362,N_19297,N_17600);
or U20363 (N_20363,N_17572,N_19409);
and U20364 (N_20364,N_18133,N_17658);
xor U20365 (N_20365,N_19405,N_19806);
and U20366 (N_20366,N_19199,N_19552);
nor U20367 (N_20367,N_17549,N_19482);
nor U20368 (N_20368,N_19615,N_17694);
nor U20369 (N_20369,N_19101,N_17715);
nor U20370 (N_20370,N_19239,N_18729);
and U20371 (N_20371,N_19838,N_19145);
and U20372 (N_20372,N_19467,N_18395);
nor U20373 (N_20373,N_17725,N_19172);
xor U20374 (N_20374,N_19104,N_19893);
nand U20375 (N_20375,N_19457,N_18316);
nand U20376 (N_20376,N_19422,N_17627);
nand U20377 (N_20377,N_19298,N_18763);
xor U20378 (N_20378,N_19915,N_17910);
and U20379 (N_20379,N_18747,N_18503);
nand U20380 (N_20380,N_19860,N_18233);
and U20381 (N_20381,N_17529,N_18901);
xor U20382 (N_20382,N_19395,N_17573);
nor U20383 (N_20383,N_19248,N_18514);
nand U20384 (N_20384,N_19701,N_19659);
or U20385 (N_20385,N_17892,N_18794);
nand U20386 (N_20386,N_19898,N_17700);
nand U20387 (N_20387,N_18519,N_19626);
and U20388 (N_20388,N_19621,N_17662);
xor U20389 (N_20389,N_18170,N_19460);
or U20390 (N_20390,N_19700,N_18095);
nand U20391 (N_20391,N_19594,N_17901);
or U20392 (N_20392,N_18369,N_18846);
or U20393 (N_20393,N_19788,N_19795);
nand U20394 (N_20394,N_19748,N_18952);
nand U20395 (N_20395,N_18932,N_19062);
xnor U20396 (N_20396,N_18048,N_19575);
nand U20397 (N_20397,N_19489,N_19401);
nand U20398 (N_20398,N_18079,N_19671);
nand U20399 (N_20399,N_18467,N_19094);
and U20400 (N_20400,N_18402,N_19585);
xor U20401 (N_20401,N_19513,N_18532);
xnor U20402 (N_20402,N_17585,N_18370);
nor U20403 (N_20403,N_18184,N_18145);
or U20404 (N_20404,N_19543,N_18982);
or U20405 (N_20405,N_18856,N_18801);
or U20406 (N_20406,N_18381,N_18687);
xnor U20407 (N_20407,N_18681,N_19149);
or U20408 (N_20408,N_17668,N_19914);
and U20409 (N_20409,N_17703,N_19411);
nor U20410 (N_20410,N_18500,N_19723);
or U20411 (N_20411,N_19807,N_19135);
nor U20412 (N_20412,N_17862,N_18069);
or U20413 (N_20413,N_18886,N_19252);
nor U20414 (N_20414,N_19270,N_18355);
and U20415 (N_20415,N_17863,N_18273);
nand U20416 (N_20416,N_18255,N_17641);
xor U20417 (N_20417,N_19143,N_18866);
nand U20418 (N_20418,N_17979,N_19398);
nor U20419 (N_20419,N_18081,N_18410);
nand U20420 (N_20420,N_19894,N_18459);
and U20421 (N_20421,N_19243,N_19680);
or U20422 (N_20422,N_18109,N_17752);
and U20423 (N_20423,N_18112,N_18884);
nand U20424 (N_20424,N_19763,N_19606);
nor U20425 (N_20425,N_19295,N_18101);
xnor U20426 (N_20426,N_18050,N_18264);
xnor U20427 (N_20427,N_19511,N_18920);
xor U20428 (N_20428,N_18090,N_18293);
xor U20429 (N_20429,N_17840,N_18163);
and U20430 (N_20430,N_19445,N_17754);
or U20431 (N_20431,N_18262,N_19889);
nor U20432 (N_20432,N_18029,N_17779);
and U20433 (N_20433,N_18151,N_19568);
xor U20434 (N_20434,N_19391,N_18975);
nor U20435 (N_20435,N_17826,N_17841);
nor U20436 (N_20436,N_19840,N_19384);
xnor U20437 (N_20437,N_19020,N_18584);
nor U20438 (N_20438,N_17519,N_18894);
or U20439 (N_20439,N_19661,N_17751);
or U20440 (N_20440,N_19309,N_19151);
xnor U20441 (N_20441,N_19009,N_17689);
or U20442 (N_20442,N_18153,N_18433);
nand U20443 (N_20443,N_19078,N_19999);
and U20444 (N_20444,N_18495,N_17762);
xnor U20445 (N_20445,N_19486,N_18665);
and U20446 (N_20446,N_19414,N_17931);
or U20447 (N_20447,N_18678,N_19406);
or U20448 (N_20448,N_17911,N_17978);
or U20449 (N_20449,N_19591,N_18523);
and U20450 (N_20450,N_17801,N_19592);
xor U20451 (N_20451,N_17562,N_19681);
nor U20452 (N_20452,N_17525,N_17880);
xor U20453 (N_20453,N_17989,N_19163);
nand U20454 (N_20454,N_19458,N_19649);
nand U20455 (N_20455,N_18818,N_19452);
and U20456 (N_20456,N_17849,N_18578);
or U20457 (N_20457,N_17928,N_19751);
and U20458 (N_20458,N_19875,N_17935);
nand U20459 (N_20459,N_17594,N_19155);
nor U20460 (N_20460,N_19991,N_18428);
nand U20461 (N_20461,N_18110,N_19500);
nor U20462 (N_20462,N_19563,N_18857);
nor U20463 (N_20463,N_17868,N_17929);
and U20464 (N_20464,N_18527,N_18075);
nand U20465 (N_20465,N_18215,N_18298);
nor U20466 (N_20466,N_19633,N_19026);
or U20467 (N_20467,N_17500,N_18306);
nand U20468 (N_20468,N_17986,N_18774);
nand U20469 (N_20469,N_18968,N_18310);
and U20470 (N_20470,N_19928,N_18147);
nor U20471 (N_20471,N_19400,N_18536);
nor U20472 (N_20472,N_19978,N_19537);
xor U20473 (N_20473,N_18385,N_18261);
nand U20474 (N_20474,N_18671,N_17720);
or U20475 (N_20475,N_18438,N_18352);
or U20476 (N_20476,N_17744,N_18144);
xnor U20477 (N_20477,N_18116,N_19862);
or U20478 (N_20478,N_19903,N_17985);
nand U20479 (N_20479,N_19945,N_19739);
or U20480 (N_20480,N_17920,N_17959);
or U20481 (N_20481,N_17997,N_17909);
nand U20482 (N_20482,N_19013,N_19200);
nor U20483 (N_20483,N_19988,N_19947);
xnor U20484 (N_20484,N_17665,N_18783);
nand U20485 (N_20485,N_19363,N_17726);
xnor U20486 (N_20486,N_18282,N_19586);
xnor U20487 (N_20487,N_17571,N_18852);
nand U20488 (N_20488,N_19229,N_18034);
xor U20489 (N_20489,N_19197,N_17699);
nor U20490 (N_20490,N_19497,N_18705);
nor U20491 (N_20491,N_18821,N_18797);
nand U20492 (N_20492,N_19214,N_18553);
nand U20493 (N_20493,N_19257,N_18568);
xnor U20494 (N_20494,N_19336,N_18323);
nor U20495 (N_20495,N_18980,N_18617);
xnor U20496 (N_20496,N_18335,N_17967);
and U20497 (N_20497,N_19103,N_17853);
nand U20498 (N_20498,N_18674,N_18531);
and U20499 (N_20499,N_18089,N_17612);
or U20500 (N_20500,N_18838,N_19783);
and U20501 (N_20501,N_19762,N_18431);
nor U20502 (N_20502,N_19941,N_19854);
and U20503 (N_20503,N_17538,N_19442);
and U20504 (N_20504,N_17589,N_18150);
and U20505 (N_20505,N_19417,N_17518);
nor U20506 (N_20506,N_19359,N_18718);
xor U20507 (N_20507,N_18638,N_19822);
nor U20508 (N_20508,N_18627,N_18097);
nor U20509 (N_20509,N_18978,N_17778);
or U20510 (N_20510,N_18844,N_18823);
or U20511 (N_20511,N_19464,N_18326);
or U20512 (N_20512,N_17982,N_18582);
nand U20513 (N_20513,N_19623,N_19108);
xnor U20514 (N_20514,N_18782,N_18498);
or U20515 (N_20515,N_19100,N_17810);
nand U20516 (N_20516,N_18525,N_18787);
nand U20517 (N_20517,N_18929,N_19056);
xor U20518 (N_20518,N_17509,N_17551);
nand U20519 (N_20519,N_18212,N_17962);
nand U20520 (N_20520,N_17858,N_18793);
and U20521 (N_20521,N_17721,N_18124);
and U20522 (N_20522,N_18171,N_17738);
nor U20523 (N_20523,N_19705,N_19035);
nor U20524 (N_20524,N_17682,N_18263);
or U20525 (N_20525,N_18719,N_19975);
and U20526 (N_20526,N_19861,N_17580);
or U20527 (N_20527,N_19003,N_18509);
xor U20528 (N_20528,N_17772,N_17767);
nand U20529 (N_20529,N_17913,N_18209);
nor U20530 (N_20530,N_18332,N_18027);
nand U20531 (N_20531,N_18266,N_19109);
or U20532 (N_20532,N_18279,N_17977);
or U20533 (N_20533,N_19599,N_19699);
or U20534 (N_20534,N_18411,N_17995);
xnor U20535 (N_20535,N_19275,N_18979);
nor U20536 (N_20536,N_18764,N_17657);
xor U20537 (N_20537,N_19749,N_17539);
xnor U20538 (N_20538,N_18731,N_18115);
and U20539 (N_20539,N_17739,N_18563);
and U20540 (N_20540,N_18628,N_17661);
nor U20541 (N_20541,N_19937,N_19226);
nand U20542 (N_20542,N_19105,N_19287);
xnor U20543 (N_20543,N_19278,N_19331);
nand U20544 (N_20544,N_18328,N_19379);
or U20545 (N_20545,N_18008,N_19549);
and U20546 (N_20546,N_18716,N_19198);
or U20547 (N_20547,N_19030,N_19936);
and U20548 (N_20548,N_19407,N_19002);
nor U20549 (N_20549,N_18146,N_17820);
nor U20550 (N_20550,N_19887,N_17702);
and U20551 (N_20551,N_18862,N_18403);
and U20552 (N_20552,N_18329,N_17652);
nor U20553 (N_20553,N_18570,N_19721);
nor U20554 (N_20554,N_18843,N_18879);
nor U20555 (N_20555,N_18598,N_17842);
nor U20556 (N_20556,N_19154,N_19765);
and U20557 (N_20557,N_19085,N_17506);
or U20558 (N_20558,N_17764,N_18162);
or U20559 (N_20559,N_19580,N_17686);
xnor U20560 (N_20560,N_19702,N_17719);
nand U20561 (N_20561,N_19834,N_18506);
nor U20562 (N_20562,N_19688,N_18581);
and U20563 (N_20563,N_17507,N_19061);
or U20564 (N_20564,N_19195,N_18158);
nand U20565 (N_20565,N_19112,N_18604);
xor U20566 (N_20566,N_18148,N_17796);
xnor U20567 (N_20567,N_19416,N_19694);
nand U20568 (N_20568,N_19043,N_18165);
nor U20569 (N_20569,N_18052,N_17983);
and U20570 (N_20570,N_18639,N_17905);
nand U20571 (N_20571,N_17793,N_19219);
nand U20572 (N_20572,N_18241,N_17961);
nand U20573 (N_20573,N_18590,N_18387);
or U20574 (N_20574,N_17684,N_18276);
and U20575 (N_20575,N_18019,N_18014);
nand U20576 (N_20576,N_18446,N_19827);
or U20577 (N_20577,N_19554,N_17753);
xnor U20578 (N_20578,N_19017,N_18738);
and U20579 (N_20579,N_17633,N_18003);
nor U20580 (N_20580,N_19816,N_18448);
xor U20581 (N_20581,N_18798,N_18668);
nor U20582 (N_20582,N_18804,N_18889);
or U20583 (N_20583,N_19823,N_19211);
nand U20584 (N_20584,N_18543,N_18615);
xor U20585 (N_20585,N_18301,N_19318);
nand U20586 (N_20586,N_17745,N_18922);
and U20587 (N_20587,N_17763,N_19299);
xor U20588 (N_20588,N_18780,N_19576);
nor U20589 (N_20589,N_19107,N_19373);
xor U20590 (N_20590,N_18680,N_18739);
or U20591 (N_20591,N_18679,N_17611);
nor U20592 (N_20592,N_17794,N_19029);
and U20593 (N_20593,N_18006,N_17800);
nor U20594 (N_20594,N_17642,N_19116);
or U20595 (N_20595,N_17948,N_18749);
or U20596 (N_20596,N_19567,N_18737);
or U20597 (N_20597,N_18605,N_17640);
nor U20598 (N_20598,N_17654,N_18760);
nand U20599 (N_20599,N_19603,N_19092);
xnor U20600 (N_20600,N_18667,N_19668);
nor U20601 (N_20601,N_17619,N_19118);
nor U20602 (N_20602,N_19939,N_19502);
xor U20603 (N_20603,N_18197,N_18558);
xor U20604 (N_20604,N_18516,N_18827);
nand U20605 (N_20605,N_19522,N_18875);
nand U20606 (N_20606,N_19325,N_19246);
and U20607 (N_20607,N_18142,N_18022);
xor U20608 (N_20608,N_19487,N_18710);
nand U20609 (N_20609,N_18723,N_19216);
nand U20610 (N_20610,N_19535,N_19444);
nor U20611 (N_20611,N_17586,N_18394);
and U20612 (N_20612,N_18533,N_18539);
nor U20613 (N_20613,N_18464,N_17846);
or U20614 (N_20614,N_19106,N_18925);
or U20615 (N_20615,N_17653,N_18534);
nor U20616 (N_20616,N_19698,N_18045);
nor U20617 (N_20617,N_18913,N_19130);
nand U20618 (N_20618,N_19040,N_19597);
and U20619 (N_20619,N_18881,N_19872);
xnor U20620 (N_20620,N_17647,N_18330);
and U20621 (N_20621,N_17757,N_19874);
or U20622 (N_20622,N_19726,N_17822);
nor U20623 (N_20623,N_18005,N_18805);
nand U20624 (N_20624,N_17896,N_18409);
xnor U20625 (N_20625,N_19133,N_18559);
nand U20626 (N_20626,N_19461,N_19624);
or U20627 (N_20627,N_17577,N_18304);
and U20628 (N_20628,N_18786,N_19387);
or U20629 (N_20629,N_18819,N_17543);
xor U20630 (N_20630,N_19473,N_17774);
or U20631 (N_20631,N_17791,N_19691);
nor U20632 (N_20632,N_18947,N_19328);
and U20633 (N_20633,N_19439,N_19672);
nand U20634 (N_20634,N_17555,N_17552);
nor U20635 (N_20635,N_17865,N_17866);
and U20636 (N_20636,N_17884,N_19221);
and U20637 (N_20637,N_19173,N_18129);
xnor U20638 (N_20638,N_18223,N_18453);
and U20639 (N_20639,N_19754,N_18327);
and U20640 (N_20640,N_18859,N_18704);
xnor U20641 (N_20641,N_18750,N_19162);
or U20642 (N_20642,N_18175,N_18073);
nor U20643 (N_20643,N_18663,N_18353);
or U20644 (N_20644,N_19912,N_18841);
or U20645 (N_20645,N_19609,N_18535);
or U20646 (N_20646,N_19523,N_19504);
xnor U20647 (N_20647,N_19998,N_17797);
nand U20648 (N_20648,N_18344,N_19761);
nand U20649 (N_20649,N_19053,N_19536);
and U20650 (N_20650,N_18571,N_19595);
xnor U20651 (N_20651,N_19206,N_17804);
xnor U20652 (N_20652,N_18572,N_19911);
nor U20653 (N_20653,N_19082,N_19375);
nand U20654 (N_20654,N_19849,N_19496);
nand U20655 (N_20655,N_19720,N_19250);
xor U20656 (N_20656,N_18885,N_18832);
and U20657 (N_20657,N_19503,N_18993);
nor U20658 (N_20658,N_19653,N_17511);
nor U20659 (N_20659,N_19622,N_18181);
nor U20660 (N_20660,N_18088,N_19168);
nor U20661 (N_20661,N_19164,N_19069);
xnor U20662 (N_20662,N_18573,N_19813);
nor U20663 (N_20663,N_18172,N_19985);
and U20664 (N_20664,N_18985,N_18367);
and U20665 (N_20665,N_19818,N_18646);
xor U20666 (N_20666,N_19641,N_19208);
and U20667 (N_20667,N_18830,N_18232);
or U20668 (N_20668,N_19908,N_17965);
nand U20669 (N_20669,N_19954,N_18105);
and U20670 (N_20670,N_18616,N_19581);
nor U20671 (N_20671,N_17883,N_19265);
and U20672 (N_20672,N_19230,N_18732);
or U20673 (N_20673,N_17714,N_18630);
nor U20674 (N_20674,N_18831,N_17648);
nor U20675 (N_20675,N_19737,N_18675);
xnor U20676 (N_20676,N_17693,N_18653);
and U20677 (N_20677,N_18924,N_19212);
nand U20678 (N_20678,N_18249,N_17843);
and U20679 (N_20679,N_17930,N_18918);
and U20680 (N_20680,N_18015,N_19476);
nand U20681 (N_20681,N_19972,N_19369);
or U20682 (N_20682,N_18647,N_18248);
xor U20683 (N_20683,N_18940,N_17620);
nor U20684 (N_20684,N_18366,N_19977);
xor U20685 (N_20685,N_18969,N_17861);
nand U20686 (N_20686,N_18733,N_18715);
nor U20687 (N_20687,N_19420,N_18033);
and U20688 (N_20688,N_19449,N_19448);
nand U20689 (N_20689,N_19682,N_19110);
or U20690 (N_20690,N_18324,N_19712);
or U20691 (N_20691,N_18222,N_18709);
or U20692 (N_20692,N_19613,N_17713);
nor U20693 (N_20693,N_18936,N_17771);
or U20694 (N_20694,N_19974,N_18451);
xor U20695 (N_20695,N_19354,N_17914);
xnor U20696 (N_20696,N_18359,N_18206);
or U20697 (N_20697,N_17876,N_18267);
nand U20698 (N_20698,N_18935,N_18664);
and U20699 (N_20699,N_18921,N_18895);
nor U20700 (N_20700,N_19938,N_18333);
nand U20701 (N_20701,N_19231,N_19990);
or U20702 (N_20702,N_19188,N_17781);
nor U20703 (N_20703,N_18104,N_18444);
nand U20704 (N_20704,N_19165,N_18926);
or U20705 (N_20705,N_18280,N_18713);
and U20706 (N_20706,N_19228,N_18318);
nand U20707 (N_20707,N_17533,N_17785);
nand U20708 (N_20708,N_17787,N_18480);
nor U20709 (N_20709,N_18400,N_19789);
xor U20710 (N_20710,N_19024,N_18836);
nor U20711 (N_20711,N_18566,N_18393);
nor U20712 (N_20712,N_17663,N_19993);
and U20713 (N_20713,N_19740,N_19019);
nand U20714 (N_20714,N_17821,N_19269);
nand U20715 (N_20715,N_17877,N_19553);
or U20716 (N_20716,N_18977,N_18228);
nand U20717 (N_20717,N_19223,N_17993);
or U20718 (N_20718,N_19935,N_19435);
nor U20719 (N_20719,N_17701,N_18896);
xnor U20720 (N_20720,N_18141,N_18501);
nand U20721 (N_20721,N_18250,N_19924);
nor U20722 (N_20722,N_17938,N_19904);
nand U20723 (N_20723,N_18247,N_17617);
nor U20724 (N_20724,N_18595,N_17664);
nand U20725 (N_20725,N_18690,N_19088);
nand U20726 (N_20726,N_19709,N_18291);
and U20727 (N_20727,N_17520,N_18123);
nand U20728 (N_20728,N_17953,N_19314);
nor U20729 (N_20729,N_18998,N_17964);
xor U20730 (N_20730,N_19706,N_18554);
nand U20731 (N_20731,N_19747,N_17954);
and U20732 (N_20732,N_18765,N_18012);
xnor U20733 (N_20733,N_17937,N_19471);
xor U20734 (N_20734,N_18454,N_18849);
xor U20735 (N_20735,N_19450,N_18071);
and U20736 (N_20736,N_19815,N_18898);
nor U20737 (N_20737,N_17643,N_18575);
nand U20738 (N_20738,N_18221,N_19266);
nor U20739 (N_20739,N_18803,N_18131);
xor U20740 (N_20740,N_19742,N_18305);
nor U20741 (N_20741,N_18207,N_18195);
nand U20742 (N_20742,N_18772,N_18130);
or U20743 (N_20743,N_17712,N_19870);
nor U20744 (N_20744,N_19663,N_19083);
and U20745 (N_20745,N_19153,N_19001);
xor U20746 (N_20746,N_19408,N_19897);
nand U20747 (N_20747,N_19656,N_18970);
nand U20748 (N_20748,N_18654,N_17770);
xnor U20749 (N_20749,N_19925,N_18309);
or U20750 (N_20750,N_19477,N_17941);
xnor U20751 (N_20751,N_18317,N_19800);
and U20752 (N_20752,N_18152,N_17607);
or U20753 (N_20753,N_18911,N_18962);
nor U20754 (N_20754,N_19693,N_18186);
xnor U20755 (N_20755,N_19131,N_19890);
and U20756 (N_20756,N_18910,N_18791);
xnor U20757 (N_20757,N_19651,N_19725);
and U20758 (N_20758,N_19768,N_18867);
nand U20759 (N_20759,N_17603,N_19334);
xnor U20760 (N_20760,N_19923,N_18417);
nand U20761 (N_20761,N_18824,N_18251);
nor U20762 (N_20762,N_17558,N_18576);
nor U20763 (N_20763,N_17530,N_17606);
xnor U20764 (N_20764,N_19282,N_18337);
nor U20765 (N_20765,N_18708,N_17832);
or U20766 (N_20766,N_18839,N_18528);
nor U20767 (N_20767,N_18773,N_19650);
xor U20768 (N_20768,N_19689,N_17723);
or U20769 (N_20769,N_19888,N_19617);
nor U20770 (N_20770,N_18858,N_17802);
or U20771 (N_20771,N_18308,N_19213);
xor U20772 (N_20772,N_19646,N_18642);
and U20773 (N_20773,N_17864,N_17513);
and U20774 (N_20774,N_17970,N_18637);
nor U20775 (N_20775,N_19632,N_19004);
nor U20776 (N_20776,N_19909,N_18644);
and U20777 (N_20777,N_19204,N_19215);
and U20778 (N_20778,N_17882,N_17685);
nor U20779 (N_20779,N_19356,N_19086);
xor U20780 (N_20780,N_17927,N_18203);
xnor U20781 (N_20781,N_18524,N_19321);
and U20782 (N_20782,N_18463,N_19812);
nor U20783 (N_20783,N_18371,N_17670);
nor U20784 (N_20784,N_17939,N_19926);
nor U20785 (N_20785,N_19602,N_19483);
and U20786 (N_20786,N_18025,N_18777);
nand U20787 (N_20787,N_18484,N_18802);
or U20788 (N_20788,N_18108,N_19236);
nand U20789 (N_20789,N_19828,N_19814);
xor U20790 (N_20790,N_19465,N_18829);
nor U20791 (N_20791,N_19907,N_17674);
nand U20792 (N_20792,N_19235,N_18191);
xnor U20793 (N_20793,N_18976,N_18244);
nor U20794 (N_20794,N_19605,N_18906);
and U20795 (N_20795,N_19719,N_19931);
and U20796 (N_20796,N_18107,N_19760);
nor U20797 (N_20797,N_19184,N_18082);
xnor U20798 (N_20798,N_17681,N_19505);
nand U20799 (N_20799,N_19796,N_19713);
nor U20800 (N_20800,N_18959,N_17769);
xnor U20801 (N_20801,N_18187,N_19902);
xnor U20802 (N_20802,N_18603,N_18767);
nor U20803 (N_20803,N_19964,N_17955);
nand U20804 (N_20804,N_19579,N_17777);
and U20805 (N_20805,N_18004,N_18950);
and U20806 (N_20806,N_19871,N_19311);
or U20807 (N_20807,N_18490,N_19962);
xnor U20808 (N_20808,N_17756,N_19531);
or U20809 (N_20809,N_19731,N_19791);
and U20810 (N_20810,N_17564,N_19025);
xor U20811 (N_20811,N_19771,N_18021);
nand U20812 (N_20812,N_19156,N_18111);
nand U20813 (N_20813,N_17582,N_19224);
nor U20814 (N_20814,N_19821,N_19868);
nor U20815 (N_20815,N_18795,N_19799);
nand U20816 (N_20816,N_19474,N_19628);
xnor U20817 (N_20817,N_19378,N_19940);
xnor U20818 (N_20818,N_19498,N_18987);
nand U20819 (N_20819,N_19811,N_19054);
xor U20820 (N_20820,N_18288,N_17923);
or U20821 (N_20821,N_19469,N_18167);
and U20822 (N_20822,N_19494,N_19185);
nor U20823 (N_20823,N_17799,N_18776);
nand U20824 (N_20824,N_19073,N_19959);
xor U20825 (N_20825,N_19468,N_18420);
and U20826 (N_20826,N_17854,N_19046);
nand U20827 (N_20827,N_19957,N_19520);
nor U20828 (N_20828,N_18289,N_17695);
nand U20829 (N_20829,N_18766,N_19548);
nor U20830 (N_20830,N_17856,N_18743);
nand U20831 (N_20831,N_17574,N_18927);
xnor U20832 (N_20832,N_19804,N_18775);
nand U20833 (N_20833,N_18039,N_19995);
xnor U20834 (N_20834,N_17706,N_17515);
nor U20835 (N_20835,N_18230,N_18166);
xnor U20836 (N_20836,N_18054,N_17690);
xor U20837 (N_20837,N_18990,N_18336);
xnor U20838 (N_20838,N_18038,N_19717);
and U20839 (N_20839,N_19125,N_19332);
xnor U20840 (N_20840,N_18157,N_18651);
xnor U20841 (N_20841,N_19766,N_19087);
nand U20842 (N_20842,N_18210,N_18689);
and U20843 (N_20843,N_17831,N_17784);
xnor U20844 (N_20844,N_19755,N_19366);
and U20845 (N_20845,N_18265,N_19119);
xor U20846 (N_20846,N_17502,N_17987);
or U20847 (N_20847,N_17847,N_19750);
or U20848 (N_20848,N_19285,N_19171);
and U20849 (N_20849,N_19683,N_19283);
xor U20850 (N_20850,N_19930,N_18942);
or U20851 (N_20851,N_18056,N_19148);
nand U20852 (N_20852,N_18084,N_18064);
nand U20853 (N_20853,N_19456,N_18648);
nand U20854 (N_20854,N_17737,N_18468);
xor U20855 (N_20855,N_18547,N_17718);
or U20856 (N_20856,N_17897,N_19027);
or U20857 (N_20857,N_17644,N_17677);
nor U20858 (N_20858,N_18815,N_18872);
nand U20859 (N_20859,N_19381,N_19355);
xor U20860 (N_20860,N_19308,N_18494);
or U20861 (N_20861,N_19284,N_19256);
nor U20862 (N_20862,N_17716,N_18693);
xnor U20863 (N_20863,N_17833,N_18621);
xnor U20864 (N_20864,N_17707,N_17733);
and U20865 (N_20865,N_18656,N_18725);
and U20866 (N_20866,N_18847,N_19565);
nor U20867 (N_20867,N_19488,N_17988);
nor U20868 (N_20868,N_19485,N_17742);
nand U20869 (N_20869,N_18430,N_18365);
or U20870 (N_20870,N_17724,N_17535);
and U20871 (N_20871,N_19389,N_17765);
xnor U20872 (N_20872,N_19630,N_18155);
xor U20873 (N_20873,N_19524,N_17729);
nand U20874 (N_20874,N_19859,N_19735);
nor U20875 (N_20875,N_17960,N_19276);
and U20876 (N_20876,N_18608,N_19501);
nand U20877 (N_20877,N_19950,N_18188);
xnor U20878 (N_20878,N_18345,N_17828);
xnor U20879 (N_20879,N_17730,N_19045);
nand U20880 (N_20880,N_18748,N_18196);
and U20881 (N_20881,N_19320,N_19562);
nor U20882 (N_20882,N_19058,N_17646);
nor U20883 (N_20883,N_19346,N_17660);
and U20884 (N_20884,N_19115,N_18848);
or U20885 (N_20885,N_19951,N_18356);
nand U20886 (N_20886,N_19852,N_19540);
nand U20887 (N_20887,N_18868,N_17873);
xnor U20888 (N_20888,N_18252,N_19512);
xnor U20889 (N_20889,N_18099,N_19006);
xnor U20890 (N_20890,N_19113,N_18024);
and U20891 (N_20891,N_18600,N_19778);
or U20892 (N_20892,N_19418,N_18149);
nor U20893 (N_20893,N_18350,N_19177);
or U20894 (N_20894,N_18042,N_17587);
and U20895 (N_20895,N_18799,N_18569);
and U20896 (N_20896,N_18007,N_18778);
nand U20897 (N_20897,N_18392,N_19021);
nand U20898 (N_20898,N_19986,N_19329);
xor U20899 (N_20899,N_18635,N_19005);
nand U20900 (N_20900,N_18915,N_19994);
xnor U20901 (N_20901,N_18820,N_19773);
and U20902 (N_20902,N_17634,N_18684);
xor U20903 (N_20903,N_17736,N_19843);
or U20904 (N_20904,N_19969,N_19310);
nor U20905 (N_20905,N_18951,N_19886);
or U20906 (N_20906,N_19538,N_19853);
and U20907 (N_20907,N_19880,N_19057);
or U20908 (N_20908,N_17829,N_18373);
nand U20909 (N_20909,N_17803,N_19787);
and U20910 (N_20910,N_18530,N_18414);
and U20911 (N_20911,N_17709,N_19317);
xnor U20912 (N_20912,N_18812,N_19393);
and U20913 (N_20913,N_18991,N_18808);
and U20914 (N_20914,N_17817,N_18194);
xnor U20915 (N_20915,N_18672,N_18483);
xnor U20916 (N_20916,N_19288,N_17554);
xnor U20917 (N_20917,N_19556,N_19249);
or U20918 (N_20918,N_18139,N_17890);
nor U20919 (N_20919,N_18046,N_19829);
nor U20920 (N_20920,N_18810,N_18470);
or U20921 (N_20921,N_19943,N_17852);
nor U20922 (N_20922,N_19326,N_18458);
nor U20923 (N_20923,N_18299,N_18135);
nor U20924 (N_20924,N_17547,N_19247);
or U20925 (N_20925,N_19922,N_17944);
nand U20926 (N_20926,N_19983,N_18726);
nand U20927 (N_20927,N_17921,N_19696);
and U20928 (N_20928,N_18683,N_18286);
nand U20929 (N_20929,N_18599,N_19367);
or U20930 (N_20930,N_18692,N_17818);
nor U20931 (N_20931,N_17559,N_17874);
xor U20932 (N_20932,N_18580,N_18557);
nor U20933 (N_20933,N_18361,N_19291);
nand U20934 (N_20934,N_17649,N_17656);
nor U20935 (N_20935,N_17544,N_17563);
or U20936 (N_20936,N_19820,N_18473);
nor U20937 (N_20937,N_19906,N_18552);
or U20938 (N_20938,N_18564,N_18051);
or U20939 (N_20939,N_18413,N_19167);
xnor U20940 (N_20940,N_18860,N_18701);
and U20941 (N_20941,N_18338,N_19841);
nor U20942 (N_20942,N_18346,N_19427);
nor U20943 (N_20943,N_18931,N_17768);
nand U20944 (N_20944,N_19826,N_19598);
and U20945 (N_20945,N_18806,N_17578);
xnor U20946 (N_20946,N_19059,N_19138);
nor U20947 (N_20947,N_19643,N_19194);
xor U20948 (N_20948,N_19454,N_19472);
or U20949 (N_20949,N_19744,N_19399);
or U20950 (N_20950,N_18908,N_19315);
nand U20951 (N_20951,N_17602,N_17830);
nand U20952 (N_20952,N_17814,N_17645);
nand U20953 (N_20953,N_18311,N_17691);
and U20954 (N_20954,N_18193,N_18032);
nand U20955 (N_20955,N_17676,N_18429);
or U20956 (N_20956,N_18620,N_18902);
nand U20957 (N_20957,N_19881,N_17540);
nor U20958 (N_20958,N_17545,N_17501);
nor U20959 (N_20959,N_17508,N_18423);
nor U20960 (N_20960,N_18427,N_19865);
nand U20961 (N_20961,N_18650,N_17592);
nand U20962 (N_20962,N_19244,N_17922);
and U20963 (N_20963,N_18436,N_19732);
nand U20964 (N_20964,N_19267,N_18076);
nand U20965 (N_20965,N_18472,N_18407);
xor U20966 (N_20966,N_19264,N_19403);
nand U20967 (N_20967,N_18294,N_18202);
or U20968 (N_20968,N_18611,N_19979);
or U20969 (N_20969,N_18093,N_19186);
and U20970 (N_20970,N_18550,N_19560);
or U20971 (N_20971,N_17836,N_18752);
nor U20972 (N_20972,N_17904,N_19507);
nand U20973 (N_20973,N_18814,N_18634);
or U20974 (N_20974,N_18404,N_18809);
xnor U20975 (N_20975,N_17523,N_17811);
or U20976 (N_20976,N_17947,N_18140);
or U20977 (N_20977,N_19665,N_18278);
xnor U20978 (N_20978,N_18938,N_18796);
or U20979 (N_20979,N_19847,N_19601);
nor U20980 (N_20980,N_18437,N_17639);
or U20981 (N_20981,N_18800,N_18119);
xor U20982 (N_20982,N_18861,N_18488);
and U20983 (N_20983,N_19376,N_19339);
nand U20984 (N_20984,N_17630,N_18416);
nor U20985 (N_20985,N_17886,N_19205);
and U20986 (N_20986,N_18169,N_19692);
or U20987 (N_20987,N_19657,N_18917);
and U20988 (N_20988,N_18624,N_18220);
or U20989 (N_20989,N_18712,N_19798);
xnor U20990 (N_20990,N_17597,N_19809);
xnor U20991 (N_20991,N_18443,N_18313);
or U20992 (N_20992,N_18347,N_18907);
or U20993 (N_20993,N_18231,N_19144);
xor U20994 (N_20994,N_18043,N_19960);
nor U20995 (N_20995,N_18660,N_19627);
nor U20996 (N_20996,N_17517,N_19837);
or U20997 (N_20997,N_18703,N_18632);
or U20998 (N_20998,N_17747,N_19634);
nand U20999 (N_20999,N_17598,N_19636);
xnor U21000 (N_21000,N_19182,N_19038);
nand U21001 (N_21001,N_19836,N_19517);
nand U21002 (N_21002,N_19674,N_18658);
xor U21003 (N_21003,N_18061,N_19873);
nand U21004 (N_21004,N_19340,N_19530);
nand U21005 (N_21005,N_19016,N_18013);
nor U21006 (N_21006,N_19342,N_19981);
or U21007 (N_21007,N_18295,N_18770);
nand U21008 (N_21008,N_18023,N_18030);
nor U21009 (N_21009,N_18315,N_17705);
and U21010 (N_21010,N_19878,N_17618);
nor U21011 (N_21011,N_19345,N_17942);
xor U21012 (N_21012,N_17885,N_19161);
nor U21013 (N_21013,N_19987,N_18482);
xnor U21014 (N_21014,N_19697,N_18619);
nand U21015 (N_21015,N_17848,N_18011);
nor U21016 (N_21016,N_18243,N_17614);
xor U21017 (N_21017,N_19631,N_19348);
nand U21018 (N_21018,N_17990,N_18117);
nor U21019 (N_21019,N_18270,N_19508);
nor U21020 (N_21020,N_17788,N_18476);
nor U21021 (N_21021,N_17601,N_19905);
nor U21022 (N_21022,N_19316,N_18253);
nand U21023 (N_21023,N_18229,N_19493);
or U21024 (N_21024,N_17871,N_19187);
xor U21025 (N_21025,N_18173,N_17789);
and U21026 (N_21026,N_18017,N_18751);
xnor U21027 (N_21027,N_18873,N_18981);
xnor U21028 (N_21028,N_19207,N_19490);
or U21029 (N_21029,N_19690,N_18587);
nand U21030 (N_21030,N_19102,N_18303);
nor U21031 (N_21031,N_19123,N_18419);
nor U21032 (N_21032,N_19189,N_19625);
and U21033 (N_21033,N_19971,N_19569);
or U21034 (N_21034,N_18562,N_18614);
nor U21035 (N_21035,N_18657,N_19324);
and U21036 (N_21036,N_19984,N_19050);
nand U21037 (N_21037,N_19519,N_19313);
nand U21038 (N_21038,N_17510,N_17870);
nor U21039 (N_21039,N_18697,N_19254);
nor U21040 (N_21040,N_17859,N_19948);
nor U21041 (N_21041,N_18183,N_19428);
nand U21042 (N_21042,N_17734,N_18741);
or U21043 (N_21043,N_18125,N_19388);
nand U21044 (N_21044,N_19170,N_19516);
or U21045 (N_21045,N_18083,N_19772);
xnor U21046 (N_21046,N_18396,N_19867);
or U21047 (N_21047,N_17659,N_17557);
nor U21048 (N_21048,N_17867,N_18736);
nand U21049 (N_21049,N_19589,N_17669);
or U21050 (N_21050,N_19715,N_18479);
or U21051 (N_21051,N_17576,N_17891);
or U21052 (N_21052,N_17697,N_17556);
or U21053 (N_21053,N_18916,N_17504);
nand U21054 (N_21054,N_17609,N_17667);
or U21055 (N_21055,N_18629,N_18469);
nand U21056 (N_21056,N_19070,N_17759);
or U21057 (N_21057,N_19743,N_19955);
or U21058 (N_21058,N_17887,N_19031);
or U21059 (N_21059,N_17711,N_19241);
or U21060 (N_21060,N_19433,N_18497);
nor U21061 (N_21061,N_19122,N_19150);
nor U21062 (N_21062,N_18953,N_19041);
or U21063 (N_21063,N_18254,N_19572);
or U21064 (N_21064,N_19347,N_18505);
nor U21065 (N_21065,N_19178,N_18457);
xnor U21066 (N_21066,N_18840,N_19022);
xor U21067 (N_21067,N_17940,N_18670);
and U21068 (N_21068,N_19209,N_18788);
xnor U21069 (N_21069,N_18339,N_17613);
or U21070 (N_21070,N_19075,N_17775);
xnor U21071 (N_21071,N_18507,N_19303);
or U21072 (N_21072,N_19459,N_19196);
and U21073 (N_21073,N_18284,N_19810);
nor U21074 (N_21074,N_19616,N_18585);
nor U21075 (N_21075,N_18035,N_19667);
xnor U21076 (N_21076,N_18077,N_19210);
xnor U21077 (N_21077,N_19281,N_19660);
nor U21078 (N_21078,N_17635,N_19529);
and U21079 (N_21079,N_19652,N_17950);
nor U21080 (N_21080,N_19525,N_17528);
nand U21081 (N_21081,N_19738,N_17780);
nand U21082 (N_21082,N_18164,N_19918);
and U21083 (N_21083,N_17623,N_18322);
or U21084 (N_21084,N_19608,N_18502);
xnor U21085 (N_21085,N_19629,N_17593);
nand U21086 (N_21086,N_19166,N_19350);
and U21087 (N_21087,N_18958,N_17758);
xnor U21088 (N_21088,N_18178,N_19610);
nand U21089 (N_21089,N_19679,N_18044);
and U21090 (N_21090,N_17672,N_18246);
nand U21091 (N_21091,N_17575,N_19618);
nor U21092 (N_21092,N_19758,N_17546);
and U21093 (N_21093,N_19965,N_19174);
nor U21094 (N_21094,N_18272,N_18643);
xor U21095 (N_21095,N_17869,N_19337);
nor U21096 (N_21096,N_18372,N_19492);
xnor U21097 (N_21097,N_19558,N_17992);
nor U21098 (N_21098,N_18560,N_18489);
and U21099 (N_21099,N_18989,N_19386);
or U21100 (N_21100,N_18652,N_19891);
xnor U21101 (N_21101,N_19526,N_17741);
nand U21102 (N_21102,N_18622,N_17857);
and U21103 (N_21103,N_18510,N_18159);
and U21104 (N_21104,N_18179,N_18529);
nand U21105 (N_21105,N_18268,N_18486);
nor U21106 (N_21106,N_17671,N_19008);
nand U21107 (N_21107,N_19775,N_19158);
and U21108 (N_21108,N_18730,N_19047);
xor U21109 (N_21109,N_17631,N_17806);
nor U21110 (N_21110,N_18996,N_18899);
nand U21111 (N_21111,N_17746,N_17893);
and U21112 (N_21112,N_19268,N_18412);
xnor U21113 (N_21113,N_19515,N_18640);
nand U21114 (N_21114,N_18865,N_18702);
nand U21115 (N_21115,N_18340,N_18714);
xnor U21116 (N_21116,N_19425,N_18900);
and U21117 (N_21117,N_18943,N_18132);
and U21118 (N_21118,N_19351,N_19074);
and U21119 (N_21119,N_17760,N_17917);
nand U21120 (N_21120,N_19607,N_19333);
or U21121 (N_21121,N_18234,N_19917);
nand U21122 (N_21122,N_19479,N_19604);
or U21123 (N_21123,N_17626,N_19846);
xnor U21124 (N_21124,N_18213,N_19745);
nand U21125 (N_21125,N_18677,N_19296);
or U21126 (N_21126,N_18699,N_18589);
nand U21127 (N_21127,N_19060,N_19010);
xor U21128 (N_21128,N_19805,N_18120);
nand U21129 (N_21129,N_19614,N_19587);
and U21130 (N_21130,N_17888,N_19097);
and U21131 (N_21131,N_17566,N_18707);
nand U21132 (N_21132,N_17975,N_18000);
nor U21133 (N_21133,N_17584,N_18334);
xor U21134 (N_21134,N_19114,N_18236);
nand U21135 (N_21135,N_18390,N_18226);
and U21136 (N_21136,N_19564,N_19953);
and U21137 (N_21137,N_18759,N_17595);
nor U21138 (N_21138,N_18807,N_17991);
and U21139 (N_21139,N_18792,N_19499);
and U21140 (N_21140,N_19830,N_18127);
nor U21141 (N_21141,N_18422,N_19802);
xor U21142 (N_21142,N_19933,N_18971);
and U21143 (N_21143,N_19142,N_18060);
nand U21144 (N_21144,N_18986,N_19794);
nor U21145 (N_21145,N_19277,N_17638);
nand U21146 (N_21146,N_17503,N_18874);
or U21147 (N_21147,N_18504,N_18445);
nand U21148 (N_21148,N_18225,N_17534);
and U21149 (N_21149,N_19952,N_18020);
nor U21150 (N_21150,N_18526,N_17568);
nand U21151 (N_21151,N_17825,N_17984);
and U21152 (N_21152,N_18669,N_18724);
xor U21153 (N_21153,N_17809,N_19259);
and U21154 (N_21154,N_18905,N_19913);
xor U21155 (N_21155,N_18358,N_19707);
nand U21156 (N_21156,N_18487,N_18287);
xnor U21157 (N_21157,N_17792,N_19117);
and U21158 (N_21158,N_18666,N_17708);
xnor U21159 (N_21159,N_18757,N_18870);
and U21160 (N_21160,N_19261,N_17740);
xor U21161 (N_21161,N_19015,N_19440);
xor U21162 (N_21162,N_19655,N_18973);
xor U21163 (N_21163,N_18695,N_17900);
nand U21164 (N_21164,N_19678,N_18485);
nand U21165 (N_21165,N_18106,N_19443);
nand U21166 (N_21166,N_19635,N_18967);
xnor U21167 (N_21167,N_18452,N_19844);
or U21168 (N_21168,N_18481,N_18377);
and U21169 (N_21169,N_19413,N_17824);
xnor U21170 (N_21170,N_18676,N_18161);
nor U21171 (N_21171,N_19642,N_19545);
or U21172 (N_21172,N_18296,N_19850);
nand U21173 (N_21173,N_18992,N_19546);
and U21174 (N_21174,N_19434,N_18645);
xnor U21175 (N_21175,N_19857,N_19808);
xnor U21176 (N_21176,N_18439,N_17748);
xnor U21177 (N_21177,N_19662,N_19711);
and U21178 (N_21178,N_17958,N_17782);
nor U21179 (N_21179,N_18711,N_19335);
or U21180 (N_21180,N_19245,N_18592);
nor U21181 (N_21181,N_19251,N_19160);
and U21182 (N_21182,N_18706,N_19169);
nand U21183 (N_21183,N_19323,N_18307);
or U21184 (N_21184,N_18477,N_19934);
xor U21185 (N_21185,N_18813,N_19929);
xnor U21186 (N_21186,N_17845,N_18511);
xnor U21187 (N_21187,N_19360,N_17850);
xor U21188 (N_21188,N_19302,N_18028);
or U21189 (N_21189,N_19383,N_18891);
nand U21190 (N_21190,N_19645,N_18544);
xor U21191 (N_21191,N_18177,N_18883);
xnor U21192 (N_21192,N_17956,N_18271);
or U21193 (N_21193,N_18956,N_17907);
and U21194 (N_21194,N_18275,N_19996);
and U21195 (N_21195,N_18240,N_19415);
or U21196 (N_21196,N_17872,N_19396);
and U21197 (N_21197,N_19648,N_17851);
nor U21198 (N_21198,N_19292,N_18103);
xnor U21199 (N_21199,N_19695,N_17561);
nor U21200 (N_21200,N_19394,N_19989);
nand U21201 (N_21201,N_19506,N_17976);
and U21202 (N_21202,N_19098,N_17946);
or U21203 (N_21203,N_19441,N_19640);
nor U21204 (N_21204,N_18784,N_19179);
nand U21205 (N_21205,N_18415,N_19759);
and U21206 (N_21206,N_18058,N_18607);
nor U21207 (N_21207,N_18871,N_18518);
and U21208 (N_21208,N_18010,N_18349);
nor U21209 (N_21209,N_19380,N_18391);
nor U21210 (N_21210,N_18928,N_19064);
xnor U21211 (N_21211,N_19767,N_18909);
xor U21212 (N_21212,N_17805,N_19037);
nor U21213 (N_21213,N_19583,N_19666);
xor U21214 (N_21214,N_19111,N_19273);
nor U21215 (N_21215,N_17727,N_19480);
xnor U21216 (N_21216,N_18779,N_18040);
xor U21217 (N_21217,N_18449,N_18565);
xnor U21218 (N_21218,N_19757,N_19832);
nand U21219 (N_21219,N_17966,N_18122);
xnor U21220 (N_21220,N_19128,N_18567);
or U21221 (N_21221,N_19769,N_17666);
nand U21222 (N_21222,N_19181,N_18673);
nand U21223 (N_21223,N_19842,N_19664);
and U21224 (N_21224,N_19790,N_18541);
and U21225 (N_21225,N_18972,N_18398);
xnor U21226 (N_21226,N_19048,N_18216);
nand U21227 (N_21227,N_18098,N_19072);
and U21228 (N_21228,N_19495,N_19637);
nand U21229 (N_21229,N_19848,N_17604);
xnor U21230 (N_21230,N_18331,N_19319);
nand U21231 (N_21231,N_19364,N_18292);
and U21232 (N_21232,N_19462,N_17650);
nand U21233 (N_21233,N_17834,N_18062);
nand U21234 (N_21234,N_18218,N_19136);
nor U21235 (N_21235,N_19718,N_17951);
nand U21236 (N_21236,N_17608,N_17679);
nor U21237 (N_21237,N_19175,N_19819);
and U21238 (N_21238,N_18984,N_19357);
and U21239 (N_21239,N_19159,N_17655);
and U21240 (N_21240,N_18834,N_19063);
nand U21241 (N_21241,N_19817,N_18168);
or U21242 (N_21242,N_18049,N_17906);
nor U21243 (N_21243,N_19708,N_19833);
or U21244 (N_21244,N_19593,N_17969);
and U21245 (N_21245,N_19797,N_19963);
nor U21246 (N_21246,N_18378,N_18418);
or U21247 (N_21247,N_19561,N_18134);
nand U21248 (N_21248,N_18113,N_17835);
nand U21249 (N_21249,N_18059,N_17588);
nand U21250 (N_21250,N_18319,N_19444);
xnor U21251 (N_21251,N_19555,N_18144);
or U21252 (N_21252,N_18198,N_19400);
nand U21253 (N_21253,N_17692,N_19912);
and U21254 (N_21254,N_19745,N_19525);
nand U21255 (N_21255,N_17760,N_18732);
xnor U21256 (N_21256,N_19003,N_19608);
nand U21257 (N_21257,N_19294,N_18605);
xnor U21258 (N_21258,N_19196,N_18626);
and U21259 (N_21259,N_19010,N_17607);
xor U21260 (N_21260,N_18804,N_19678);
xor U21261 (N_21261,N_19112,N_17638);
and U21262 (N_21262,N_19171,N_18894);
or U21263 (N_21263,N_19050,N_19906);
nand U21264 (N_21264,N_18109,N_19409);
xnor U21265 (N_21265,N_18566,N_18165);
or U21266 (N_21266,N_19705,N_18583);
and U21267 (N_21267,N_18544,N_18791);
and U21268 (N_21268,N_18512,N_17916);
xnor U21269 (N_21269,N_18102,N_19235);
xor U21270 (N_21270,N_18628,N_19569);
xor U21271 (N_21271,N_18214,N_19944);
xor U21272 (N_21272,N_19299,N_19064);
nor U21273 (N_21273,N_17884,N_18638);
nor U21274 (N_21274,N_19356,N_19476);
and U21275 (N_21275,N_19061,N_17882);
nor U21276 (N_21276,N_18299,N_18790);
xor U21277 (N_21277,N_19141,N_18757);
nor U21278 (N_21278,N_19771,N_18099);
or U21279 (N_21279,N_17974,N_18416);
and U21280 (N_21280,N_17989,N_18486);
or U21281 (N_21281,N_18183,N_18366);
nand U21282 (N_21282,N_19469,N_18496);
nand U21283 (N_21283,N_19591,N_18540);
xnor U21284 (N_21284,N_18144,N_17988);
or U21285 (N_21285,N_17919,N_17868);
nand U21286 (N_21286,N_17728,N_17788);
nor U21287 (N_21287,N_19760,N_19315);
nor U21288 (N_21288,N_19458,N_17597);
or U21289 (N_21289,N_19751,N_17674);
or U21290 (N_21290,N_19254,N_18778);
and U21291 (N_21291,N_18275,N_18740);
xnor U21292 (N_21292,N_18949,N_17648);
and U21293 (N_21293,N_18007,N_19006);
nand U21294 (N_21294,N_17663,N_19975);
and U21295 (N_21295,N_18236,N_18267);
or U21296 (N_21296,N_18001,N_19614);
xor U21297 (N_21297,N_19769,N_19197);
xnor U21298 (N_21298,N_19210,N_19459);
or U21299 (N_21299,N_19487,N_19123);
and U21300 (N_21300,N_18942,N_18100);
or U21301 (N_21301,N_18843,N_19015);
or U21302 (N_21302,N_17535,N_18728);
nand U21303 (N_21303,N_18942,N_17816);
or U21304 (N_21304,N_19021,N_18464);
nor U21305 (N_21305,N_19960,N_18188);
or U21306 (N_21306,N_18668,N_19414);
nand U21307 (N_21307,N_18080,N_19863);
or U21308 (N_21308,N_18432,N_19678);
xor U21309 (N_21309,N_18728,N_17961);
nand U21310 (N_21310,N_18242,N_19916);
or U21311 (N_21311,N_18031,N_18235);
and U21312 (N_21312,N_18744,N_18486);
and U21313 (N_21313,N_18986,N_17730);
and U21314 (N_21314,N_18520,N_18178);
xnor U21315 (N_21315,N_18108,N_18121);
nor U21316 (N_21316,N_19248,N_17562);
nand U21317 (N_21317,N_19740,N_17938);
nand U21318 (N_21318,N_17614,N_18352);
and U21319 (N_21319,N_18550,N_18008);
xnor U21320 (N_21320,N_18897,N_17597);
or U21321 (N_21321,N_19105,N_19213);
nand U21322 (N_21322,N_18649,N_18186);
and U21323 (N_21323,N_18903,N_18598);
nand U21324 (N_21324,N_19116,N_19576);
nor U21325 (N_21325,N_19391,N_17736);
nor U21326 (N_21326,N_18526,N_18140);
and U21327 (N_21327,N_19547,N_18347);
nand U21328 (N_21328,N_17921,N_19292);
nor U21329 (N_21329,N_19460,N_18951);
and U21330 (N_21330,N_19275,N_17605);
xnor U21331 (N_21331,N_18816,N_18041);
nor U21332 (N_21332,N_18124,N_18755);
xor U21333 (N_21333,N_18201,N_19147);
nand U21334 (N_21334,N_17942,N_18145);
or U21335 (N_21335,N_18513,N_18589);
or U21336 (N_21336,N_18292,N_19592);
or U21337 (N_21337,N_18466,N_18399);
xnor U21338 (N_21338,N_17882,N_19889);
and U21339 (N_21339,N_19768,N_17863);
nor U21340 (N_21340,N_18004,N_18937);
xnor U21341 (N_21341,N_19001,N_18886);
and U21342 (N_21342,N_19555,N_18161);
xor U21343 (N_21343,N_19345,N_19145);
and U21344 (N_21344,N_19476,N_18960);
or U21345 (N_21345,N_18608,N_19105);
xnor U21346 (N_21346,N_19257,N_19640);
and U21347 (N_21347,N_17639,N_19566);
and U21348 (N_21348,N_19895,N_17794);
xor U21349 (N_21349,N_18650,N_17585);
nand U21350 (N_21350,N_17519,N_19184);
nor U21351 (N_21351,N_18958,N_17524);
and U21352 (N_21352,N_18937,N_19727);
and U21353 (N_21353,N_18768,N_18181);
and U21354 (N_21354,N_18405,N_18998);
xor U21355 (N_21355,N_18497,N_17890);
xnor U21356 (N_21356,N_18763,N_18495);
nor U21357 (N_21357,N_18630,N_19869);
nor U21358 (N_21358,N_19156,N_19990);
or U21359 (N_21359,N_18017,N_18992);
nand U21360 (N_21360,N_17634,N_17728);
and U21361 (N_21361,N_19307,N_19816);
and U21362 (N_21362,N_18176,N_18480);
and U21363 (N_21363,N_18918,N_18588);
nand U21364 (N_21364,N_19564,N_18634);
nand U21365 (N_21365,N_17649,N_19784);
nand U21366 (N_21366,N_18261,N_19546);
and U21367 (N_21367,N_19690,N_17776);
or U21368 (N_21368,N_19289,N_18291);
nor U21369 (N_21369,N_18210,N_19378);
or U21370 (N_21370,N_19989,N_18621);
nor U21371 (N_21371,N_17577,N_19329);
and U21372 (N_21372,N_18497,N_18525);
nor U21373 (N_21373,N_19618,N_17840);
and U21374 (N_21374,N_18976,N_18557);
xnor U21375 (N_21375,N_19400,N_17552);
and U21376 (N_21376,N_19900,N_17722);
or U21377 (N_21377,N_17954,N_19643);
nand U21378 (N_21378,N_19727,N_19513);
nand U21379 (N_21379,N_17981,N_19572);
or U21380 (N_21380,N_17624,N_19177);
nand U21381 (N_21381,N_17952,N_18543);
and U21382 (N_21382,N_19196,N_17933);
nand U21383 (N_21383,N_19328,N_18292);
xor U21384 (N_21384,N_18910,N_19191);
nand U21385 (N_21385,N_18819,N_19733);
xnor U21386 (N_21386,N_18033,N_18289);
nand U21387 (N_21387,N_18310,N_18089);
nor U21388 (N_21388,N_18565,N_18377);
nor U21389 (N_21389,N_19385,N_19202);
or U21390 (N_21390,N_18460,N_17823);
or U21391 (N_21391,N_17692,N_18607);
and U21392 (N_21392,N_18657,N_18164);
or U21393 (N_21393,N_18122,N_17771);
or U21394 (N_21394,N_19866,N_18450);
nor U21395 (N_21395,N_18263,N_19700);
nand U21396 (N_21396,N_18144,N_18762);
nand U21397 (N_21397,N_18949,N_18148);
nor U21398 (N_21398,N_19651,N_17646);
and U21399 (N_21399,N_19329,N_18341);
nand U21400 (N_21400,N_18558,N_17633);
or U21401 (N_21401,N_19456,N_17899);
or U21402 (N_21402,N_19953,N_19095);
xor U21403 (N_21403,N_19364,N_19818);
nor U21404 (N_21404,N_17757,N_19088);
and U21405 (N_21405,N_17533,N_18107);
xnor U21406 (N_21406,N_19878,N_19117);
and U21407 (N_21407,N_19859,N_18329);
nand U21408 (N_21408,N_18394,N_18907);
xor U21409 (N_21409,N_17995,N_18056);
nor U21410 (N_21410,N_19013,N_18067);
and U21411 (N_21411,N_18224,N_18772);
nand U21412 (N_21412,N_18519,N_19150);
nor U21413 (N_21413,N_17902,N_19210);
nor U21414 (N_21414,N_17530,N_18777);
or U21415 (N_21415,N_17942,N_19448);
xnor U21416 (N_21416,N_18371,N_17771);
and U21417 (N_21417,N_19871,N_19947);
xor U21418 (N_21418,N_18574,N_17619);
and U21419 (N_21419,N_18474,N_19173);
and U21420 (N_21420,N_17579,N_17930);
nand U21421 (N_21421,N_18159,N_18521);
nor U21422 (N_21422,N_17675,N_19190);
nand U21423 (N_21423,N_19935,N_19454);
nand U21424 (N_21424,N_18009,N_18975);
nand U21425 (N_21425,N_18898,N_18483);
xnor U21426 (N_21426,N_17821,N_17501);
nand U21427 (N_21427,N_18777,N_17872);
and U21428 (N_21428,N_18271,N_18886);
and U21429 (N_21429,N_18303,N_17928);
or U21430 (N_21430,N_19513,N_18292);
xnor U21431 (N_21431,N_18577,N_19272);
nor U21432 (N_21432,N_17882,N_18797);
xor U21433 (N_21433,N_19516,N_19308);
or U21434 (N_21434,N_17672,N_19274);
and U21435 (N_21435,N_17671,N_19012);
or U21436 (N_21436,N_17734,N_19101);
nor U21437 (N_21437,N_17645,N_18005);
nand U21438 (N_21438,N_17664,N_19926);
nor U21439 (N_21439,N_18862,N_18331);
nor U21440 (N_21440,N_17724,N_18829);
or U21441 (N_21441,N_18917,N_18514);
nor U21442 (N_21442,N_18486,N_18464);
xor U21443 (N_21443,N_19451,N_19670);
and U21444 (N_21444,N_18114,N_19157);
or U21445 (N_21445,N_18008,N_18049);
nor U21446 (N_21446,N_19373,N_18589);
nor U21447 (N_21447,N_18860,N_19400);
nand U21448 (N_21448,N_19360,N_19374);
nand U21449 (N_21449,N_19435,N_19021);
nand U21450 (N_21450,N_17755,N_18966);
and U21451 (N_21451,N_19937,N_19264);
and U21452 (N_21452,N_19756,N_18026);
nor U21453 (N_21453,N_18424,N_18346);
and U21454 (N_21454,N_19785,N_19544);
or U21455 (N_21455,N_18613,N_18475);
xor U21456 (N_21456,N_19970,N_19333);
xor U21457 (N_21457,N_18995,N_19143);
and U21458 (N_21458,N_19868,N_18092);
or U21459 (N_21459,N_18373,N_19873);
nor U21460 (N_21460,N_19204,N_19092);
or U21461 (N_21461,N_19523,N_19509);
nand U21462 (N_21462,N_18661,N_19398);
nor U21463 (N_21463,N_18769,N_19107);
xnor U21464 (N_21464,N_18818,N_18082);
and U21465 (N_21465,N_19827,N_18955);
or U21466 (N_21466,N_18223,N_18177);
or U21467 (N_21467,N_18718,N_19600);
nand U21468 (N_21468,N_17657,N_18433);
nor U21469 (N_21469,N_19297,N_17749);
and U21470 (N_21470,N_18334,N_18868);
and U21471 (N_21471,N_19710,N_18027);
or U21472 (N_21472,N_18226,N_19974);
nand U21473 (N_21473,N_19250,N_19249);
or U21474 (N_21474,N_17691,N_17719);
xor U21475 (N_21475,N_19011,N_18113);
xor U21476 (N_21476,N_19113,N_18757);
nor U21477 (N_21477,N_19060,N_19103);
and U21478 (N_21478,N_17611,N_17758);
nor U21479 (N_21479,N_19772,N_17910);
xor U21480 (N_21480,N_17768,N_19237);
nor U21481 (N_21481,N_17796,N_17589);
nand U21482 (N_21482,N_17563,N_19744);
nor U21483 (N_21483,N_18424,N_18186);
nor U21484 (N_21484,N_17934,N_18677);
and U21485 (N_21485,N_19171,N_18150);
xnor U21486 (N_21486,N_18424,N_19849);
nand U21487 (N_21487,N_19460,N_18412);
and U21488 (N_21488,N_18002,N_19495);
nor U21489 (N_21489,N_17531,N_17631);
nand U21490 (N_21490,N_18871,N_19497);
or U21491 (N_21491,N_19343,N_19351);
and U21492 (N_21492,N_17735,N_19535);
nand U21493 (N_21493,N_19710,N_17715);
nand U21494 (N_21494,N_18086,N_18541);
or U21495 (N_21495,N_18456,N_17828);
and U21496 (N_21496,N_18991,N_18709);
and U21497 (N_21497,N_17958,N_19521);
nand U21498 (N_21498,N_18988,N_18425);
xnor U21499 (N_21499,N_19650,N_17570);
nand U21500 (N_21500,N_17507,N_17827);
or U21501 (N_21501,N_18797,N_17794);
and U21502 (N_21502,N_17914,N_19483);
xor U21503 (N_21503,N_18938,N_17658);
and U21504 (N_21504,N_17624,N_18517);
xnor U21505 (N_21505,N_18553,N_18724);
nor U21506 (N_21506,N_19730,N_17628);
xnor U21507 (N_21507,N_19395,N_19250);
or U21508 (N_21508,N_18915,N_17537);
and U21509 (N_21509,N_18167,N_17564);
nor U21510 (N_21510,N_19361,N_17818);
xor U21511 (N_21511,N_17566,N_18674);
nand U21512 (N_21512,N_19316,N_19289);
and U21513 (N_21513,N_19740,N_18329);
or U21514 (N_21514,N_18950,N_18159);
or U21515 (N_21515,N_18733,N_18003);
and U21516 (N_21516,N_19627,N_17796);
and U21517 (N_21517,N_19495,N_19675);
nor U21518 (N_21518,N_18990,N_19321);
nand U21519 (N_21519,N_19192,N_18206);
xor U21520 (N_21520,N_17913,N_18223);
or U21521 (N_21521,N_17874,N_17698);
nor U21522 (N_21522,N_19526,N_19048);
xnor U21523 (N_21523,N_17928,N_18051);
and U21524 (N_21524,N_18625,N_19784);
xnor U21525 (N_21525,N_17723,N_19848);
or U21526 (N_21526,N_19209,N_18118);
nand U21527 (N_21527,N_19197,N_18875);
xnor U21528 (N_21528,N_19038,N_18867);
nand U21529 (N_21529,N_19435,N_18359);
nor U21530 (N_21530,N_18555,N_19475);
or U21531 (N_21531,N_17767,N_18561);
and U21532 (N_21532,N_19726,N_17876);
nor U21533 (N_21533,N_17915,N_18827);
nand U21534 (N_21534,N_17594,N_17998);
and U21535 (N_21535,N_19839,N_19612);
xor U21536 (N_21536,N_19677,N_18583);
and U21537 (N_21537,N_17523,N_19887);
or U21538 (N_21538,N_19491,N_18125);
or U21539 (N_21539,N_18602,N_18094);
or U21540 (N_21540,N_17523,N_19035);
and U21541 (N_21541,N_19139,N_19376);
and U21542 (N_21542,N_18601,N_19407);
and U21543 (N_21543,N_18357,N_18686);
nand U21544 (N_21544,N_18161,N_18699);
or U21545 (N_21545,N_19545,N_19895);
and U21546 (N_21546,N_19283,N_18610);
or U21547 (N_21547,N_19557,N_17874);
nand U21548 (N_21548,N_19903,N_17976);
and U21549 (N_21549,N_19384,N_19998);
and U21550 (N_21550,N_18357,N_19791);
xor U21551 (N_21551,N_19288,N_18081);
or U21552 (N_21552,N_18860,N_18905);
or U21553 (N_21553,N_18523,N_17937);
xnor U21554 (N_21554,N_19090,N_18536);
and U21555 (N_21555,N_18950,N_18124);
nand U21556 (N_21556,N_18535,N_18972);
or U21557 (N_21557,N_17668,N_18430);
xor U21558 (N_21558,N_19984,N_18107);
nor U21559 (N_21559,N_17778,N_18239);
xnor U21560 (N_21560,N_19826,N_19265);
or U21561 (N_21561,N_19926,N_19563);
and U21562 (N_21562,N_18351,N_19408);
and U21563 (N_21563,N_18702,N_17820);
nor U21564 (N_21564,N_19340,N_19958);
nand U21565 (N_21565,N_17866,N_18126);
nand U21566 (N_21566,N_17677,N_19431);
and U21567 (N_21567,N_19521,N_18178);
and U21568 (N_21568,N_18668,N_19633);
and U21569 (N_21569,N_17743,N_18965);
xnor U21570 (N_21570,N_17625,N_19286);
xnor U21571 (N_21571,N_18245,N_19439);
or U21572 (N_21572,N_19916,N_18810);
nand U21573 (N_21573,N_19436,N_18501);
nand U21574 (N_21574,N_19970,N_19703);
and U21575 (N_21575,N_19838,N_17700);
nor U21576 (N_21576,N_18716,N_19093);
and U21577 (N_21577,N_17546,N_19619);
or U21578 (N_21578,N_19801,N_19314);
or U21579 (N_21579,N_19589,N_18865);
and U21580 (N_21580,N_18795,N_19144);
and U21581 (N_21581,N_19748,N_18612);
nor U21582 (N_21582,N_19605,N_18582);
or U21583 (N_21583,N_19041,N_19099);
nand U21584 (N_21584,N_18937,N_18554);
nand U21585 (N_21585,N_19434,N_18172);
nor U21586 (N_21586,N_18563,N_18780);
nor U21587 (N_21587,N_19454,N_19535);
nand U21588 (N_21588,N_18424,N_18889);
and U21589 (N_21589,N_19237,N_19525);
or U21590 (N_21590,N_17978,N_19719);
and U21591 (N_21591,N_19319,N_18930);
xnor U21592 (N_21592,N_18706,N_18002);
xor U21593 (N_21593,N_18920,N_17635);
and U21594 (N_21594,N_18776,N_19901);
nor U21595 (N_21595,N_19849,N_18889);
and U21596 (N_21596,N_18777,N_18374);
xnor U21597 (N_21597,N_19246,N_19490);
nor U21598 (N_21598,N_18847,N_18238);
xor U21599 (N_21599,N_17722,N_19985);
nand U21600 (N_21600,N_18499,N_19570);
nor U21601 (N_21601,N_17597,N_17933);
and U21602 (N_21602,N_19977,N_19698);
nor U21603 (N_21603,N_18298,N_17959);
xor U21604 (N_21604,N_17501,N_19594);
nand U21605 (N_21605,N_17588,N_18597);
and U21606 (N_21606,N_18574,N_18382);
xor U21607 (N_21607,N_18668,N_19489);
or U21608 (N_21608,N_18595,N_18429);
or U21609 (N_21609,N_19830,N_19278);
nor U21610 (N_21610,N_19543,N_19800);
or U21611 (N_21611,N_19608,N_19441);
or U21612 (N_21612,N_18274,N_17717);
and U21613 (N_21613,N_17847,N_18628);
nand U21614 (N_21614,N_18452,N_18550);
and U21615 (N_21615,N_19396,N_19684);
or U21616 (N_21616,N_19137,N_17796);
and U21617 (N_21617,N_19812,N_19329);
nand U21618 (N_21618,N_17954,N_18185);
nor U21619 (N_21619,N_18482,N_18505);
and U21620 (N_21620,N_18397,N_19140);
nand U21621 (N_21621,N_18523,N_19975);
nor U21622 (N_21622,N_17521,N_19234);
nor U21623 (N_21623,N_18868,N_19858);
nor U21624 (N_21624,N_17522,N_19671);
xnor U21625 (N_21625,N_18206,N_19850);
xnor U21626 (N_21626,N_19379,N_19467);
and U21627 (N_21627,N_17852,N_19590);
xnor U21628 (N_21628,N_19416,N_18969);
xnor U21629 (N_21629,N_18172,N_17747);
and U21630 (N_21630,N_18019,N_18235);
and U21631 (N_21631,N_19409,N_18269);
nor U21632 (N_21632,N_18364,N_19092);
nand U21633 (N_21633,N_17701,N_17774);
nor U21634 (N_21634,N_19642,N_18653);
xnor U21635 (N_21635,N_19247,N_19372);
nand U21636 (N_21636,N_18515,N_19112);
or U21637 (N_21637,N_18259,N_18845);
nor U21638 (N_21638,N_18027,N_18187);
nor U21639 (N_21639,N_19698,N_17946);
and U21640 (N_21640,N_18657,N_17776);
nand U21641 (N_21641,N_18483,N_17725);
and U21642 (N_21642,N_19916,N_18478);
nor U21643 (N_21643,N_18063,N_18094);
and U21644 (N_21644,N_18331,N_17937);
nand U21645 (N_21645,N_19740,N_18216);
or U21646 (N_21646,N_17582,N_18638);
and U21647 (N_21647,N_17733,N_18193);
xnor U21648 (N_21648,N_17916,N_18377);
nand U21649 (N_21649,N_18085,N_18325);
xnor U21650 (N_21650,N_18963,N_18218);
or U21651 (N_21651,N_18657,N_18303);
nand U21652 (N_21652,N_17882,N_17726);
nor U21653 (N_21653,N_18591,N_19695);
nor U21654 (N_21654,N_18534,N_18730);
nor U21655 (N_21655,N_19588,N_19726);
xor U21656 (N_21656,N_19637,N_18314);
nand U21657 (N_21657,N_17984,N_18776);
xor U21658 (N_21658,N_17501,N_17725);
and U21659 (N_21659,N_18332,N_19742);
nor U21660 (N_21660,N_18034,N_19870);
nand U21661 (N_21661,N_18498,N_18578);
nor U21662 (N_21662,N_18183,N_18764);
or U21663 (N_21663,N_18367,N_18585);
and U21664 (N_21664,N_19796,N_18437);
xnor U21665 (N_21665,N_18782,N_19078);
or U21666 (N_21666,N_19628,N_17845);
xnor U21667 (N_21667,N_19021,N_19581);
or U21668 (N_21668,N_17658,N_18167);
and U21669 (N_21669,N_17729,N_18015);
or U21670 (N_21670,N_18296,N_19269);
or U21671 (N_21671,N_19991,N_19381);
nand U21672 (N_21672,N_17561,N_18315);
and U21673 (N_21673,N_18442,N_18725);
nand U21674 (N_21674,N_19598,N_18709);
nand U21675 (N_21675,N_18979,N_17628);
xor U21676 (N_21676,N_18192,N_18161);
or U21677 (N_21677,N_19572,N_18231);
or U21678 (N_21678,N_19853,N_18690);
nor U21679 (N_21679,N_18356,N_18282);
xnor U21680 (N_21680,N_17763,N_18458);
xnor U21681 (N_21681,N_17915,N_18346);
nor U21682 (N_21682,N_18995,N_19636);
and U21683 (N_21683,N_19903,N_17947);
nand U21684 (N_21684,N_18383,N_17848);
or U21685 (N_21685,N_17849,N_18560);
nor U21686 (N_21686,N_17932,N_17506);
xor U21687 (N_21687,N_18985,N_17899);
nor U21688 (N_21688,N_18989,N_18298);
nand U21689 (N_21689,N_18710,N_18744);
xnor U21690 (N_21690,N_19397,N_19716);
or U21691 (N_21691,N_18715,N_18209);
nand U21692 (N_21692,N_17539,N_17933);
or U21693 (N_21693,N_18150,N_18258);
nor U21694 (N_21694,N_17574,N_19083);
or U21695 (N_21695,N_18834,N_19141);
or U21696 (N_21696,N_19425,N_18656);
or U21697 (N_21697,N_18550,N_19572);
and U21698 (N_21698,N_17725,N_19404);
nor U21699 (N_21699,N_18929,N_17871);
nand U21700 (N_21700,N_19741,N_18753);
nor U21701 (N_21701,N_17707,N_19024);
and U21702 (N_21702,N_19416,N_17545);
nand U21703 (N_21703,N_18533,N_18593);
and U21704 (N_21704,N_17712,N_18663);
nor U21705 (N_21705,N_18153,N_19420);
nor U21706 (N_21706,N_18512,N_19641);
xor U21707 (N_21707,N_18281,N_19841);
and U21708 (N_21708,N_18331,N_18644);
or U21709 (N_21709,N_19517,N_18187);
or U21710 (N_21710,N_18417,N_18753);
xor U21711 (N_21711,N_17716,N_19433);
xor U21712 (N_21712,N_19011,N_19446);
nor U21713 (N_21713,N_19126,N_17613);
xnor U21714 (N_21714,N_19960,N_18635);
nand U21715 (N_21715,N_17860,N_18985);
or U21716 (N_21716,N_19674,N_19921);
nand U21717 (N_21717,N_18330,N_18280);
nand U21718 (N_21718,N_18129,N_19663);
xnor U21719 (N_21719,N_18839,N_19994);
nand U21720 (N_21720,N_17878,N_19743);
nand U21721 (N_21721,N_17559,N_19616);
and U21722 (N_21722,N_19480,N_19699);
or U21723 (N_21723,N_18353,N_18263);
and U21724 (N_21724,N_18156,N_19972);
and U21725 (N_21725,N_17787,N_19330);
nand U21726 (N_21726,N_18351,N_18636);
and U21727 (N_21727,N_19735,N_18398);
nand U21728 (N_21728,N_19544,N_17909);
nor U21729 (N_21729,N_17903,N_18007);
and U21730 (N_21730,N_17955,N_18310);
nor U21731 (N_21731,N_19184,N_17636);
or U21732 (N_21732,N_18473,N_19933);
nand U21733 (N_21733,N_19975,N_18540);
or U21734 (N_21734,N_19355,N_17987);
xor U21735 (N_21735,N_17902,N_18666);
nor U21736 (N_21736,N_18105,N_19957);
nand U21737 (N_21737,N_18037,N_18927);
nor U21738 (N_21738,N_19839,N_17561);
nor U21739 (N_21739,N_19817,N_18054);
nand U21740 (N_21740,N_18748,N_17567);
nand U21741 (N_21741,N_18031,N_18180);
xnor U21742 (N_21742,N_18866,N_18830);
xor U21743 (N_21743,N_19454,N_19889);
and U21744 (N_21744,N_19682,N_18551);
xnor U21745 (N_21745,N_18915,N_19036);
and U21746 (N_21746,N_18581,N_18869);
nor U21747 (N_21747,N_18259,N_18994);
and U21748 (N_21748,N_17708,N_18525);
or U21749 (N_21749,N_17669,N_19417);
nor U21750 (N_21750,N_19419,N_19119);
xor U21751 (N_21751,N_17605,N_17896);
or U21752 (N_21752,N_18626,N_18115);
and U21753 (N_21753,N_17887,N_17907);
nand U21754 (N_21754,N_18036,N_18067);
and U21755 (N_21755,N_18882,N_18282);
xnor U21756 (N_21756,N_19349,N_19825);
and U21757 (N_21757,N_18496,N_18264);
and U21758 (N_21758,N_19323,N_19813);
and U21759 (N_21759,N_19923,N_17934);
and U21760 (N_21760,N_17535,N_18993);
nor U21761 (N_21761,N_19173,N_18924);
xor U21762 (N_21762,N_19846,N_18293);
or U21763 (N_21763,N_19875,N_19928);
nand U21764 (N_21764,N_18102,N_17799);
or U21765 (N_21765,N_19778,N_17743);
or U21766 (N_21766,N_17598,N_18700);
nor U21767 (N_21767,N_17766,N_18023);
or U21768 (N_21768,N_18611,N_19247);
or U21769 (N_21769,N_18354,N_18993);
or U21770 (N_21770,N_18204,N_18716);
nand U21771 (N_21771,N_19601,N_18557);
or U21772 (N_21772,N_19506,N_17749);
nand U21773 (N_21773,N_19302,N_17636);
nor U21774 (N_21774,N_17553,N_17688);
and U21775 (N_21775,N_18048,N_18627);
nor U21776 (N_21776,N_19202,N_19618);
nor U21777 (N_21777,N_18105,N_19841);
and U21778 (N_21778,N_18385,N_18742);
nor U21779 (N_21779,N_19963,N_17957);
nor U21780 (N_21780,N_19734,N_18229);
or U21781 (N_21781,N_17787,N_18908);
and U21782 (N_21782,N_18138,N_18177);
nand U21783 (N_21783,N_17893,N_17933);
xor U21784 (N_21784,N_18926,N_17837);
nand U21785 (N_21785,N_19511,N_18403);
nor U21786 (N_21786,N_18198,N_17720);
and U21787 (N_21787,N_18770,N_18497);
or U21788 (N_21788,N_19757,N_18178);
nand U21789 (N_21789,N_19427,N_18010);
xnor U21790 (N_21790,N_19505,N_18490);
nor U21791 (N_21791,N_18526,N_19786);
nor U21792 (N_21792,N_19536,N_19697);
nand U21793 (N_21793,N_17566,N_17581);
nor U21794 (N_21794,N_17623,N_18925);
nand U21795 (N_21795,N_19150,N_18328);
nor U21796 (N_21796,N_19021,N_17828);
and U21797 (N_21797,N_19544,N_18114);
and U21798 (N_21798,N_19158,N_18002);
or U21799 (N_21799,N_18226,N_17648);
and U21800 (N_21800,N_19103,N_19495);
xor U21801 (N_21801,N_19166,N_18350);
and U21802 (N_21802,N_18990,N_19530);
nor U21803 (N_21803,N_18758,N_17762);
nand U21804 (N_21804,N_19801,N_19557);
xor U21805 (N_21805,N_19548,N_18100);
nor U21806 (N_21806,N_19073,N_19549);
nand U21807 (N_21807,N_17586,N_18086);
nand U21808 (N_21808,N_19054,N_19189);
and U21809 (N_21809,N_19030,N_18355);
nor U21810 (N_21810,N_18672,N_19663);
xor U21811 (N_21811,N_19534,N_17832);
xnor U21812 (N_21812,N_19532,N_18758);
or U21813 (N_21813,N_19170,N_19872);
and U21814 (N_21814,N_17827,N_17522);
nand U21815 (N_21815,N_19504,N_19205);
or U21816 (N_21816,N_19817,N_18731);
xor U21817 (N_21817,N_18263,N_17731);
nor U21818 (N_21818,N_18706,N_17759);
xor U21819 (N_21819,N_19295,N_18543);
nor U21820 (N_21820,N_17649,N_19655);
xor U21821 (N_21821,N_17548,N_17926);
xor U21822 (N_21822,N_18065,N_18663);
and U21823 (N_21823,N_18615,N_18462);
and U21824 (N_21824,N_18649,N_19655);
and U21825 (N_21825,N_18362,N_19605);
nor U21826 (N_21826,N_19354,N_17856);
nand U21827 (N_21827,N_17778,N_19666);
or U21828 (N_21828,N_17566,N_18391);
nand U21829 (N_21829,N_18389,N_19629);
nand U21830 (N_21830,N_19690,N_19013);
or U21831 (N_21831,N_18955,N_17897);
nand U21832 (N_21832,N_17971,N_18876);
xor U21833 (N_21833,N_18403,N_17943);
xnor U21834 (N_21834,N_19662,N_18307);
nor U21835 (N_21835,N_19152,N_18924);
xnor U21836 (N_21836,N_19466,N_19025);
xnor U21837 (N_21837,N_17962,N_18041);
nand U21838 (N_21838,N_19952,N_19775);
nor U21839 (N_21839,N_19647,N_18832);
nor U21840 (N_21840,N_18998,N_17943);
or U21841 (N_21841,N_18828,N_18168);
nand U21842 (N_21842,N_19541,N_17741);
and U21843 (N_21843,N_19922,N_17747);
nand U21844 (N_21844,N_18829,N_19907);
and U21845 (N_21845,N_19269,N_19230);
nor U21846 (N_21846,N_19544,N_19461);
or U21847 (N_21847,N_17655,N_18499);
nor U21848 (N_21848,N_17971,N_18724);
or U21849 (N_21849,N_19726,N_17857);
and U21850 (N_21850,N_19665,N_18868);
and U21851 (N_21851,N_19469,N_17510);
or U21852 (N_21852,N_18035,N_18242);
and U21853 (N_21853,N_17855,N_19585);
or U21854 (N_21854,N_19393,N_17505);
nand U21855 (N_21855,N_17969,N_18251);
nor U21856 (N_21856,N_19817,N_19139);
xor U21857 (N_21857,N_17874,N_18514);
nand U21858 (N_21858,N_19008,N_19389);
nor U21859 (N_21859,N_18292,N_19647);
and U21860 (N_21860,N_19229,N_19505);
and U21861 (N_21861,N_19738,N_19516);
and U21862 (N_21862,N_18422,N_19665);
or U21863 (N_21863,N_17971,N_18971);
xnor U21864 (N_21864,N_19623,N_19138);
xnor U21865 (N_21865,N_18383,N_18983);
nor U21866 (N_21866,N_18202,N_18130);
and U21867 (N_21867,N_19561,N_19239);
nand U21868 (N_21868,N_17830,N_18956);
and U21869 (N_21869,N_19063,N_19449);
or U21870 (N_21870,N_18898,N_17961);
nand U21871 (N_21871,N_17790,N_18743);
nor U21872 (N_21872,N_17682,N_19587);
nor U21873 (N_21873,N_18781,N_18406);
and U21874 (N_21874,N_19315,N_17624);
and U21875 (N_21875,N_18390,N_19367);
or U21876 (N_21876,N_19380,N_18210);
or U21877 (N_21877,N_18064,N_19663);
nor U21878 (N_21878,N_17777,N_18538);
xor U21879 (N_21879,N_19766,N_19034);
or U21880 (N_21880,N_19194,N_19604);
or U21881 (N_21881,N_18415,N_19908);
and U21882 (N_21882,N_18921,N_17619);
xnor U21883 (N_21883,N_18356,N_17515);
xnor U21884 (N_21884,N_18380,N_18234);
or U21885 (N_21885,N_17650,N_19501);
xnor U21886 (N_21886,N_18753,N_19978);
or U21887 (N_21887,N_19951,N_18977);
nand U21888 (N_21888,N_19594,N_18098);
nor U21889 (N_21889,N_19782,N_18573);
xnor U21890 (N_21890,N_19989,N_19748);
nor U21891 (N_21891,N_19727,N_19587);
nor U21892 (N_21892,N_18460,N_18583);
xor U21893 (N_21893,N_18043,N_18864);
and U21894 (N_21894,N_17777,N_17811);
nor U21895 (N_21895,N_17620,N_17672);
and U21896 (N_21896,N_18554,N_18814);
and U21897 (N_21897,N_17838,N_18100);
nor U21898 (N_21898,N_18439,N_17590);
xor U21899 (N_21899,N_18414,N_18447);
nand U21900 (N_21900,N_19292,N_18031);
xor U21901 (N_21901,N_19945,N_19039);
xnor U21902 (N_21902,N_18688,N_18895);
nand U21903 (N_21903,N_17712,N_17919);
nand U21904 (N_21904,N_17504,N_17684);
nor U21905 (N_21905,N_18942,N_19426);
nor U21906 (N_21906,N_18428,N_18107);
nor U21907 (N_21907,N_19711,N_18447);
or U21908 (N_21908,N_18865,N_18652);
and U21909 (N_21909,N_18186,N_18326);
nor U21910 (N_21910,N_18638,N_18280);
nand U21911 (N_21911,N_18926,N_19636);
xor U21912 (N_21912,N_18246,N_19638);
xor U21913 (N_21913,N_17982,N_17875);
nand U21914 (N_21914,N_18708,N_19716);
xnor U21915 (N_21915,N_18636,N_18277);
or U21916 (N_21916,N_19661,N_19377);
xor U21917 (N_21917,N_18740,N_19360);
nor U21918 (N_21918,N_19162,N_18307);
or U21919 (N_21919,N_19410,N_18304);
xnor U21920 (N_21920,N_18643,N_19068);
or U21921 (N_21921,N_17531,N_18156);
nor U21922 (N_21922,N_19401,N_17531);
and U21923 (N_21923,N_17652,N_19245);
and U21924 (N_21924,N_18333,N_19423);
or U21925 (N_21925,N_18722,N_17802);
nor U21926 (N_21926,N_19485,N_17773);
nor U21927 (N_21927,N_18025,N_18309);
xnor U21928 (N_21928,N_17714,N_18291);
nor U21929 (N_21929,N_17572,N_18401);
or U21930 (N_21930,N_18707,N_17625);
and U21931 (N_21931,N_18591,N_19095);
nor U21932 (N_21932,N_18665,N_19007);
and U21933 (N_21933,N_19312,N_18487);
or U21934 (N_21934,N_18909,N_17657);
nand U21935 (N_21935,N_19031,N_19289);
nor U21936 (N_21936,N_19546,N_19024);
xor U21937 (N_21937,N_18396,N_18478);
or U21938 (N_21938,N_17708,N_17876);
xor U21939 (N_21939,N_19811,N_17692);
xnor U21940 (N_21940,N_19397,N_17511);
nand U21941 (N_21941,N_19334,N_19239);
and U21942 (N_21942,N_18819,N_17873);
and U21943 (N_21943,N_19973,N_18669);
xor U21944 (N_21944,N_19379,N_17867);
nor U21945 (N_21945,N_19265,N_18108);
nor U21946 (N_21946,N_19224,N_17776);
nor U21947 (N_21947,N_18552,N_19783);
and U21948 (N_21948,N_18831,N_18918);
nand U21949 (N_21949,N_18530,N_19225);
nor U21950 (N_21950,N_19963,N_19878);
xnor U21951 (N_21951,N_18901,N_17783);
xor U21952 (N_21952,N_19328,N_17708);
and U21953 (N_21953,N_18717,N_19207);
and U21954 (N_21954,N_19079,N_19050);
xnor U21955 (N_21955,N_18170,N_19810);
xor U21956 (N_21956,N_19282,N_19821);
nand U21957 (N_21957,N_19401,N_18126);
nor U21958 (N_21958,N_18750,N_18824);
nor U21959 (N_21959,N_18871,N_17750);
nor U21960 (N_21960,N_17605,N_19073);
or U21961 (N_21961,N_18659,N_19255);
xnor U21962 (N_21962,N_18356,N_19107);
nor U21963 (N_21963,N_18144,N_18855);
nand U21964 (N_21964,N_18673,N_17922);
or U21965 (N_21965,N_18936,N_19563);
xor U21966 (N_21966,N_18939,N_18179);
nand U21967 (N_21967,N_19088,N_19793);
nor U21968 (N_21968,N_18648,N_18965);
nor U21969 (N_21969,N_19967,N_19661);
nand U21970 (N_21970,N_18021,N_19508);
nor U21971 (N_21971,N_18678,N_19047);
xor U21972 (N_21972,N_17524,N_19527);
or U21973 (N_21973,N_17811,N_19729);
or U21974 (N_21974,N_18698,N_19757);
nand U21975 (N_21975,N_17568,N_19202);
and U21976 (N_21976,N_19256,N_18087);
xnor U21977 (N_21977,N_17914,N_19371);
xnor U21978 (N_21978,N_19167,N_18201);
and U21979 (N_21979,N_18019,N_17526);
or U21980 (N_21980,N_18363,N_18418);
nor U21981 (N_21981,N_18044,N_18133);
nand U21982 (N_21982,N_18976,N_19548);
or U21983 (N_21983,N_18230,N_19367);
nand U21984 (N_21984,N_18434,N_18985);
or U21985 (N_21985,N_18730,N_18355);
nand U21986 (N_21986,N_18260,N_18352);
xor U21987 (N_21987,N_18095,N_18519);
nand U21988 (N_21988,N_17944,N_19068);
or U21989 (N_21989,N_18935,N_17920);
xnor U21990 (N_21990,N_19367,N_17532);
nor U21991 (N_21991,N_18153,N_19640);
xor U21992 (N_21992,N_17778,N_17841);
nor U21993 (N_21993,N_19812,N_17666);
nand U21994 (N_21994,N_19014,N_19198);
nand U21995 (N_21995,N_17851,N_18435);
nand U21996 (N_21996,N_19790,N_17706);
nand U21997 (N_21997,N_17654,N_18469);
nor U21998 (N_21998,N_18582,N_19443);
nand U21999 (N_21999,N_18573,N_19504);
nand U22000 (N_22000,N_19788,N_19946);
xor U22001 (N_22001,N_18601,N_18726);
nand U22002 (N_22002,N_17551,N_18915);
or U22003 (N_22003,N_19570,N_18144);
nor U22004 (N_22004,N_19451,N_18127);
or U22005 (N_22005,N_18576,N_17700);
or U22006 (N_22006,N_19916,N_18886);
or U22007 (N_22007,N_19882,N_18846);
nand U22008 (N_22008,N_18660,N_19688);
and U22009 (N_22009,N_18871,N_17586);
or U22010 (N_22010,N_19943,N_18399);
and U22011 (N_22011,N_18135,N_19446);
or U22012 (N_22012,N_17542,N_17779);
or U22013 (N_22013,N_17639,N_17903);
and U22014 (N_22014,N_18854,N_19714);
nand U22015 (N_22015,N_19338,N_17725);
xor U22016 (N_22016,N_19104,N_18088);
nand U22017 (N_22017,N_17688,N_17811);
and U22018 (N_22018,N_19774,N_17771);
nor U22019 (N_22019,N_18142,N_18029);
or U22020 (N_22020,N_18468,N_19913);
nand U22021 (N_22021,N_19306,N_18466);
or U22022 (N_22022,N_18572,N_18723);
nor U22023 (N_22023,N_17792,N_19475);
nor U22024 (N_22024,N_19645,N_18985);
xor U22025 (N_22025,N_17990,N_17756);
and U22026 (N_22026,N_18710,N_18768);
nor U22027 (N_22027,N_19055,N_18760);
nand U22028 (N_22028,N_18377,N_18344);
xnor U22029 (N_22029,N_19255,N_19972);
nor U22030 (N_22030,N_19033,N_17614);
nor U22031 (N_22031,N_17763,N_18474);
nand U22032 (N_22032,N_17878,N_18558);
nor U22033 (N_22033,N_18270,N_18141);
and U22034 (N_22034,N_18532,N_19692);
or U22035 (N_22035,N_19942,N_18672);
xnor U22036 (N_22036,N_19613,N_19753);
nand U22037 (N_22037,N_19661,N_17721);
or U22038 (N_22038,N_18991,N_19026);
xnor U22039 (N_22039,N_18483,N_18514);
nand U22040 (N_22040,N_17624,N_19892);
nor U22041 (N_22041,N_19570,N_19408);
or U22042 (N_22042,N_19075,N_18844);
nor U22043 (N_22043,N_19508,N_19355);
and U22044 (N_22044,N_19299,N_18004);
nor U22045 (N_22045,N_19969,N_18878);
and U22046 (N_22046,N_18216,N_18192);
or U22047 (N_22047,N_19868,N_17508);
nor U22048 (N_22048,N_19346,N_18149);
nand U22049 (N_22049,N_19566,N_18484);
xor U22050 (N_22050,N_19639,N_17709);
or U22051 (N_22051,N_18054,N_18723);
nor U22052 (N_22052,N_19329,N_18926);
or U22053 (N_22053,N_18480,N_17840);
nand U22054 (N_22054,N_18650,N_18580);
and U22055 (N_22055,N_19306,N_19707);
or U22056 (N_22056,N_19440,N_18494);
and U22057 (N_22057,N_18279,N_18719);
nor U22058 (N_22058,N_18825,N_18790);
nor U22059 (N_22059,N_18229,N_17677);
or U22060 (N_22060,N_17778,N_19189);
xnor U22061 (N_22061,N_18189,N_19057);
xor U22062 (N_22062,N_18689,N_19239);
nor U22063 (N_22063,N_17702,N_19087);
nor U22064 (N_22064,N_19309,N_19883);
xor U22065 (N_22065,N_18753,N_19915);
nor U22066 (N_22066,N_19779,N_19267);
nand U22067 (N_22067,N_18975,N_17648);
and U22068 (N_22068,N_19599,N_18411);
xnor U22069 (N_22069,N_18121,N_19454);
and U22070 (N_22070,N_17925,N_18327);
nor U22071 (N_22071,N_17588,N_17533);
nor U22072 (N_22072,N_19087,N_19147);
nand U22073 (N_22073,N_18184,N_19287);
nand U22074 (N_22074,N_17923,N_18125);
nand U22075 (N_22075,N_17570,N_19353);
and U22076 (N_22076,N_17694,N_18790);
or U22077 (N_22077,N_18759,N_17962);
nand U22078 (N_22078,N_19313,N_17618);
and U22079 (N_22079,N_19460,N_17620);
nor U22080 (N_22080,N_18348,N_19990);
nor U22081 (N_22081,N_19664,N_17710);
xnor U22082 (N_22082,N_18142,N_18471);
xor U22083 (N_22083,N_18918,N_17782);
nor U22084 (N_22084,N_18547,N_18181);
nor U22085 (N_22085,N_18323,N_19928);
xnor U22086 (N_22086,N_19181,N_18569);
or U22087 (N_22087,N_19253,N_17863);
xor U22088 (N_22088,N_17948,N_18492);
nand U22089 (N_22089,N_18742,N_18596);
nand U22090 (N_22090,N_19529,N_18396);
and U22091 (N_22091,N_18424,N_19697);
nor U22092 (N_22092,N_18800,N_17923);
nand U22093 (N_22093,N_18450,N_19574);
xnor U22094 (N_22094,N_18525,N_18874);
nor U22095 (N_22095,N_18109,N_19784);
xnor U22096 (N_22096,N_19088,N_19624);
or U22097 (N_22097,N_19002,N_17799);
nor U22098 (N_22098,N_18972,N_17596);
nor U22099 (N_22099,N_19715,N_19714);
nor U22100 (N_22100,N_18762,N_18558);
xnor U22101 (N_22101,N_19023,N_18426);
nor U22102 (N_22102,N_18145,N_19105);
or U22103 (N_22103,N_18998,N_19022);
xor U22104 (N_22104,N_17867,N_18892);
or U22105 (N_22105,N_17612,N_19339);
xnor U22106 (N_22106,N_19315,N_17903);
and U22107 (N_22107,N_19334,N_18197);
nor U22108 (N_22108,N_19108,N_18507);
or U22109 (N_22109,N_19871,N_19886);
nand U22110 (N_22110,N_18217,N_19149);
or U22111 (N_22111,N_18170,N_19613);
xnor U22112 (N_22112,N_17692,N_19874);
xor U22113 (N_22113,N_18775,N_19211);
nand U22114 (N_22114,N_19044,N_19364);
xor U22115 (N_22115,N_18884,N_19504);
and U22116 (N_22116,N_17594,N_19924);
or U22117 (N_22117,N_18053,N_19029);
nor U22118 (N_22118,N_19298,N_19416);
nand U22119 (N_22119,N_19553,N_17764);
nand U22120 (N_22120,N_17880,N_17986);
or U22121 (N_22121,N_18022,N_18700);
and U22122 (N_22122,N_18142,N_19690);
or U22123 (N_22123,N_18921,N_17857);
or U22124 (N_22124,N_19169,N_19529);
nor U22125 (N_22125,N_19724,N_19683);
nand U22126 (N_22126,N_19930,N_17976);
xnor U22127 (N_22127,N_19126,N_18932);
or U22128 (N_22128,N_19613,N_18835);
nor U22129 (N_22129,N_18059,N_19817);
xnor U22130 (N_22130,N_19313,N_19949);
nand U22131 (N_22131,N_17631,N_19527);
nand U22132 (N_22132,N_19912,N_19673);
nor U22133 (N_22133,N_18174,N_18039);
or U22134 (N_22134,N_18875,N_19004);
nand U22135 (N_22135,N_19248,N_19711);
or U22136 (N_22136,N_18406,N_17602);
nand U22137 (N_22137,N_18024,N_19004);
nor U22138 (N_22138,N_17629,N_17944);
or U22139 (N_22139,N_19669,N_18345);
xor U22140 (N_22140,N_19173,N_18222);
nor U22141 (N_22141,N_17806,N_18314);
xor U22142 (N_22142,N_19383,N_19831);
xnor U22143 (N_22143,N_19861,N_18851);
nand U22144 (N_22144,N_18156,N_17509);
nand U22145 (N_22145,N_17801,N_19237);
and U22146 (N_22146,N_19600,N_19703);
nor U22147 (N_22147,N_18118,N_17914);
and U22148 (N_22148,N_18934,N_18402);
nor U22149 (N_22149,N_18881,N_17613);
xor U22150 (N_22150,N_18442,N_18699);
xor U22151 (N_22151,N_19363,N_19868);
xor U22152 (N_22152,N_19049,N_19038);
nor U22153 (N_22153,N_17622,N_17600);
nor U22154 (N_22154,N_19742,N_19004);
and U22155 (N_22155,N_19548,N_17519);
nor U22156 (N_22156,N_17944,N_19546);
and U22157 (N_22157,N_18828,N_17972);
nor U22158 (N_22158,N_19385,N_18032);
and U22159 (N_22159,N_18769,N_19049);
or U22160 (N_22160,N_19243,N_19682);
or U22161 (N_22161,N_19182,N_19601);
nand U22162 (N_22162,N_18993,N_17870);
or U22163 (N_22163,N_19497,N_18140);
nor U22164 (N_22164,N_19762,N_18223);
and U22165 (N_22165,N_18388,N_18925);
or U22166 (N_22166,N_18160,N_19170);
xor U22167 (N_22167,N_19170,N_19001);
nand U22168 (N_22168,N_18102,N_19976);
xor U22169 (N_22169,N_19573,N_17930);
xor U22170 (N_22170,N_19229,N_17660);
nand U22171 (N_22171,N_19463,N_18547);
nor U22172 (N_22172,N_19618,N_19133);
and U22173 (N_22173,N_19425,N_19027);
nor U22174 (N_22174,N_17649,N_18522);
nand U22175 (N_22175,N_18174,N_17968);
or U22176 (N_22176,N_17733,N_19583);
xor U22177 (N_22177,N_19475,N_18373);
nor U22178 (N_22178,N_19929,N_19324);
and U22179 (N_22179,N_18177,N_18272);
nor U22180 (N_22180,N_17913,N_19695);
or U22181 (N_22181,N_19610,N_18776);
nand U22182 (N_22182,N_17760,N_19551);
and U22183 (N_22183,N_19028,N_19470);
and U22184 (N_22184,N_18513,N_18501);
xnor U22185 (N_22185,N_19054,N_18361);
xor U22186 (N_22186,N_19604,N_19910);
and U22187 (N_22187,N_17938,N_19664);
nor U22188 (N_22188,N_19790,N_19017);
nor U22189 (N_22189,N_18810,N_18505);
nand U22190 (N_22190,N_19973,N_17512);
nor U22191 (N_22191,N_19294,N_18865);
nand U22192 (N_22192,N_18100,N_18776);
nand U22193 (N_22193,N_19117,N_19721);
or U22194 (N_22194,N_19506,N_18351);
xor U22195 (N_22195,N_18224,N_17696);
nand U22196 (N_22196,N_18734,N_18693);
or U22197 (N_22197,N_19617,N_19680);
or U22198 (N_22198,N_18835,N_18709);
nand U22199 (N_22199,N_17657,N_18691);
and U22200 (N_22200,N_19922,N_17976);
or U22201 (N_22201,N_19265,N_19502);
and U22202 (N_22202,N_18570,N_19243);
or U22203 (N_22203,N_19165,N_17676);
nor U22204 (N_22204,N_19958,N_19780);
nor U22205 (N_22205,N_19658,N_18597);
xor U22206 (N_22206,N_18604,N_18335);
xnor U22207 (N_22207,N_18602,N_18560);
and U22208 (N_22208,N_18917,N_18014);
nor U22209 (N_22209,N_19829,N_19410);
and U22210 (N_22210,N_18432,N_19821);
or U22211 (N_22211,N_18337,N_18750);
and U22212 (N_22212,N_18093,N_19535);
nand U22213 (N_22213,N_18798,N_19497);
and U22214 (N_22214,N_18462,N_17862);
nand U22215 (N_22215,N_17932,N_18721);
nor U22216 (N_22216,N_19766,N_19558);
nor U22217 (N_22217,N_19580,N_18382);
or U22218 (N_22218,N_18812,N_18275);
and U22219 (N_22219,N_19573,N_17680);
or U22220 (N_22220,N_18641,N_19506);
xor U22221 (N_22221,N_19335,N_17758);
or U22222 (N_22222,N_18221,N_19832);
or U22223 (N_22223,N_19880,N_18959);
or U22224 (N_22224,N_18775,N_18521);
or U22225 (N_22225,N_18270,N_18487);
nand U22226 (N_22226,N_19734,N_18445);
and U22227 (N_22227,N_17943,N_19903);
nor U22228 (N_22228,N_18010,N_19981);
and U22229 (N_22229,N_19411,N_18929);
or U22230 (N_22230,N_17545,N_19549);
and U22231 (N_22231,N_19010,N_17514);
nand U22232 (N_22232,N_19056,N_19951);
nand U22233 (N_22233,N_19185,N_18313);
nand U22234 (N_22234,N_18400,N_17506);
or U22235 (N_22235,N_18442,N_17551);
and U22236 (N_22236,N_18861,N_19280);
nand U22237 (N_22237,N_19710,N_19996);
or U22238 (N_22238,N_17764,N_19815);
xnor U22239 (N_22239,N_18361,N_18425);
or U22240 (N_22240,N_19433,N_19945);
xnor U22241 (N_22241,N_19570,N_19306);
or U22242 (N_22242,N_19565,N_17800);
nand U22243 (N_22243,N_19948,N_18292);
xnor U22244 (N_22244,N_19948,N_18420);
nand U22245 (N_22245,N_17740,N_19908);
xnor U22246 (N_22246,N_19453,N_18274);
nand U22247 (N_22247,N_18971,N_18657);
and U22248 (N_22248,N_18163,N_19414);
nand U22249 (N_22249,N_17729,N_18670);
and U22250 (N_22250,N_19382,N_18103);
nor U22251 (N_22251,N_19172,N_19971);
xor U22252 (N_22252,N_17888,N_17600);
xnor U22253 (N_22253,N_19373,N_17997);
nor U22254 (N_22254,N_19681,N_18998);
nand U22255 (N_22255,N_19884,N_19013);
nor U22256 (N_22256,N_19637,N_19348);
or U22257 (N_22257,N_19536,N_18877);
nand U22258 (N_22258,N_18051,N_19089);
and U22259 (N_22259,N_17633,N_18421);
xor U22260 (N_22260,N_18986,N_18203);
xor U22261 (N_22261,N_18115,N_18052);
nand U22262 (N_22262,N_17632,N_18517);
or U22263 (N_22263,N_19710,N_19890);
and U22264 (N_22264,N_19964,N_18182);
nand U22265 (N_22265,N_19563,N_19291);
nand U22266 (N_22266,N_18479,N_19048);
nand U22267 (N_22267,N_18760,N_18231);
nor U22268 (N_22268,N_17576,N_18995);
or U22269 (N_22269,N_19621,N_19041);
xor U22270 (N_22270,N_19618,N_19873);
and U22271 (N_22271,N_19624,N_19143);
and U22272 (N_22272,N_18782,N_18236);
nand U22273 (N_22273,N_19199,N_19783);
nand U22274 (N_22274,N_18095,N_18916);
or U22275 (N_22275,N_19014,N_17507);
xnor U22276 (N_22276,N_17764,N_18501);
or U22277 (N_22277,N_17633,N_18520);
nor U22278 (N_22278,N_19881,N_18033);
and U22279 (N_22279,N_18063,N_18726);
nand U22280 (N_22280,N_19146,N_19379);
or U22281 (N_22281,N_18563,N_19637);
nand U22282 (N_22282,N_18066,N_17545);
or U22283 (N_22283,N_19758,N_19689);
nor U22284 (N_22284,N_18805,N_17662);
and U22285 (N_22285,N_18908,N_19469);
and U22286 (N_22286,N_19125,N_18355);
or U22287 (N_22287,N_19148,N_18542);
or U22288 (N_22288,N_19019,N_18840);
or U22289 (N_22289,N_19760,N_18560);
nor U22290 (N_22290,N_17784,N_18530);
or U22291 (N_22291,N_19869,N_18192);
or U22292 (N_22292,N_17788,N_17725);
and U22293 (N_22293,N_17712,N_17714);
nand U22294 (N_22294,N_19459,N_18981);
nor U22295 (N_22295,N_18378,N_19318);
or U22296 (N_22296,N_18049,N_17793);
nand U22297 (N_22297,N_18482,N_18373);
nand U22298 (N_22298,N_19780,N_17608);
xnor U22299 (N_22299,N_18331,N_18099);
and U22300 (N_22300,N_17703,N_19160);
xor U22301 (N_22301,N_19696,N_19341);
nand U22302 (N_22302,N_18337,N_19602);
nor U22303 (N_22303,N_19883,N_17657);
and U22304 (N_22304,N_18356,N_18445);
nor U22305 (N_22305,N_17715,N_19269);
xor U22306 (N_22306,N_19579,N_19666);
xnor U22307 (N_22307,N_19606,N_17583);
and U22308 (N_22308,N_18653,N_18905);
nor U22309 (N_22309,N_19898,N_18149);
xor U22310 (N_22310,N_19525,N_18877);
and U22311 (N_22311,N_17672,N_18405);
nor U22312 (N_22312,N_18120,N_19737);
nand U22313 (N_22313,N_19897,N_17937);
nand U22314 (N_22314,N_18473,N_18670);
nor U22315 (N_22315,N_18584,N_19997);
nand U22316 (N_22316,N_17543,N_19501);
nor U22317 (N_22317,N_17906,N_19947);
nor U22318 (N_22318,N_18852,N_18902);
xnor U22319 (N_22319,N_19450,N_17607);
or U22320 (N_22320,N_19952,N_17813);
nor U22321 (N_22321,N_18348,N_19931);
nor U22322 (N_22322,N_19067,N_17593);
nand U22323 (N_22323,N_19307,N_18650);
nor U22324 (N_22324,N_18230,N_19277);
xor U22325 (N_22325,N_19263,N_19841);
xor U22326 (N_22326,N_19606,N_18822);
or U22327 (N_22327,N_17934,N_18299);
xnor U22328 (N_22328,N_18300,N_19091);
xnor U22329 (N_22329,N_19459,N_17912);
xnor U22330 (N_22330,N_19643,N_19297);
and U22331 (N_22331,N_18036,N_17882);
or U22332 (N_22332,N_18920,N_18362);
xor U22333 (N_22333,N_19377,N_18465);
nand U22334 (N_22334,N_18324,N_19677);
nor U22335 (N_22335,N_18428,N_19884);
nor U22336 (N_22336,N_18273,N_18048);
nor U22337 (N_22337,N_19087,N_19821);
nand U22338 (N_22338,N_19677,N_17602);
and U22339 (N_22339,N_19788,N_18922);
nand U22340 (N_22340,N_19011,N_19542);
nand U22341 (N_22341,N_19028,N_19377);
xnor U22342 (N_22342,N_18685,N_19853);
or U22343 (N_22343,N_18671,N_18912);
and U22344 (N_22344,N_19307,N_18896);
nor U22345 (N_22345,N_19870,N_19948);
xnor U22346 (N_22346,N_19748,N_18014);
nor U22347 (N_22347,N_19056,N_19522);
or U22348 (N_22348,N_19264,N_18513);
and U22349 (N_22349,N_17995,N_18585);
xnor U22350 (N_22350,N_18329,N_17937);
and U22351 (N_22351,N_19437,N_19686);
xor U22352 (N_22352,N_19525,N_19751);
nand U22353 (N_22353,N_18233,N_19641);
xor U22354 (N_22354,N_18334,N_18221);
and U22355 (N_22355,N_18627,N_19603);
or U22356 (N_22356,N_18944,N_18961);
nor U22357 (N_22357,N_17790,N_17703);
nor U22358 (N_22358,N_17606,N_18174);
and U22359 (N_22359,N_19490,N_19137);
nor U22360 (N_22360,N_18551,N_17797);
nor U22361 (N_22361,N_18604,N_17861);
nand U22362 (N_22362,N_18835,N_18010);
or U22363 (N_22363,N_19260,N_19072);
xnor U22364 (N_22364,N_18327,N_18308);
or U22365 (N_22365,N_17536,N_17906);
nand U22366 (N_22366,N_17642,N_18964);
and U22367 (N_22367,N_19929,N_19869);
xnor U22368 (N_22368,N_19038,N_17626);
or U22369 (N_22369,N_19187,N_18005);
xor U22370 (N_22370,N_17615,N_17506);
nor U22371 (N_22371,N_19171,N_17814);
nor U22372 (N_22372,N_19145,N_18942);
or U22373 (N_22373,N_19015,N_18504);
xor U22374 (N_22374,N_18266,N_18382);
and U22375 (N_22375,N_19307,N_19176);
and U22376 (N_22376,N_17855,N_18024);
nand U22377 (N_22377,N_18582,N_19691);
or U22378 (N_22378,N_17716,N_17841);
xor U22379 (N_22379,N_19106,N_19603);
nand U22380 (N_22380,N_18425,N_19916);
nor U22381 (N_22381,N_17711,N_17782);
nor U22382 (N_22382,N_19476,N_17764);
xnor U22383 (N_22383,N_19870,N_17773);
nor U22384 (N_22384,N_19656,N_18678);
nor U22385 (N_22385,N_19658,N_19091);
nand U22386 (N_22386,N_17967,N_18565);
or U22387 (N_22387,N_19567,N_19851);
nand U22388 (N_22388,N_18434,N_18444);
xnor U22389 (N_22389,N_19663,N_17694);
xor U22390 (N_22390,N_19199,N_19343);
or U22391 (N_22391,N_17983,N_19062);
or U22392 (N_22392,N_17795,N_18251);
xnor U22393 (N_22393,N_17896,N_19089);
nor U22394 (N_22394,N_17902,N_18833);
nand U22395 (N_22395,N_18011,N_19667);
xor U22396 (N_22396,N_18494,N_19258);
nor U22397 (N_22397,N_18209,N_19283);
and U22398 (N_22398,N_18583,N_18796);
or U22399 (N_22399,N_18180,N_17816);
and U22400 (N_22400,N_18498,N_17827);
nand U22401 (N_22401,N_17781,N_18622);
or U22402 (N_22402,N_19622,N_19693);
or U22403 (N_22403,N_17899,N_18317);
xor U22404 (N_22404,N_19398,N_19485);
nor U22405 (N_22405,N_19689,N_19701);
nand U22406 (N_22406,N_17984,N_19643);
nand U22407 (N_22407,N_19201,N_17556);
nor U22408 (N_22408,N_18684,N_17754);
nand U22409 (N_22409,N_19506,N_17997);
nor U22410 (N_22410,N_19932,N_19618);
nor U22411 (N_22411,N_18525,N_18807);
xor U22412 (N_22412,N_17530,N_18633);
and U22413 (N_22413,N_18347,N_18754);
nand U22414 (N_22414,N_18981,N_18451);
or U22415 (N_22415,N_18170,N_18604);
nor U22416 (N_22416,N_18499,N_19056);
nor U22417 (N_22417,N_18441,N_18905);
and U22418 (N_22418,N_18841,N_17648);
and U22419 (N_22419,N_19197,N_17730);
xnor U22420 (N_22420,N_18958,N_19073);
and U22421 (N_22421,N_18726,N_19202);
nor U22422 (N_22422,N_17904,N_18563);
and U22423 (N_22423,N_19883,N_18210);
nand U22424 (N_22424,N_18002,N_19312);
or U22425 (N_22425,N_19448,N_19371);
and U22426 (N_22426,N_19089,N_19583);
nand U22427 (N_22427,N_19969,N_19513);
or U22428 (N_22428,N_19917,N_18719);
nand U22429 (N_22429,N_17932,N_18963);
nand U22430 (N_22430,N_19853,N_17763);
or U22431 (N_22431,N_18827,N_19492);
or U22432 (N_22432,N_18816,N_19130);
nor U22433 (N_22433,N_17558,N_18872);
and U22434 (N_22434,N_19989,N_17993);
or U22435 (N_22435,N_19481,N_19914);
nor U22436 (N_22436,N_18808,N_18353);
nand U22437 (N_22437,N_19313,N_18765);
or U22438 (N_22438,N_19676,N_18317);
and U22439 (N_22439,N_18569,N_17637);
or U22440 (N_22440,N_19794,N_18228);
nand U22441 (N_22441,N_19953,N_18366);
and U22442 (N_22442,N_19709,N_18076);
or U22443 (N_22443,N_18917,N_19668);
nor U22444 (N_22444,N_19397,N_19923);
xor U22445 (N_22445,N_18261,N_19403);
xnor U22446 (N_22446,N_18771,N_19261);
nor U22447 (N_22447,N_17784,N_17869);
nand U22448 (N_22448,N_18212,N_17617);
and U22449 (N_22449,N_17938,N_18193);
nor U22450 (N_22450,N_17745,N_18968);
xor U22451 (N_22451,N_18516,N_17717);
or U22452 (N_22452,N_18384,N_18880);
nand U22453 (N_22453,N_17943,N_18750);
nor U22454 (N_22454,N_19056,N_18875);
xor U22455 (N_22455,N_19417,N_17586);
or U22456 (N_22456,N_19326,N_19284);
or U22457 (N_22457,N_19380,N_18020);
xor U22458 (N_22458,N_19000,N_18269);
nand U22459 (N_22459,N_19777,N_19997);
or U22460 (N_22460,N_19508,N_19647);
and U22461 (N_22461,N_18047,N_18678);
and U22462 (N_22462,N_18317,N_19036);
nor U22463 (N_22463,N_19941,N_19482);
and U22464 (N_22464,N_17569,N_19102);
xor U22465 (N_22465,N_18609,N_18881);
or U22466 (N_22466,N_19822,N_18037);
and U22467 (N_22467,N_17738,N_19774);
and U22468 (N_22468,N_19722,N_19157);
nor U22469 (N_22469,N_18940,N_18288);
or U22470 (N_22470,N_18396,N_19678);
xor U22471 (N_22471,N_17818,N_19278);
nand U22472 (N_22472,N_18052,N_18699);
and U22473 (N_22473,N_18473,N_18825);
nor U22474 (N_22474,N_19242,N_19030);
nor U22475 (N_22475,N_19909,N_17817);
nor U22476 (N_22476,N_18776,N_19788);
or U22477 (N_22477,N_18904,N_17620);
nor U22478 (N_22478,N_18143,N_18606);
or U22479 (N_22479,N_19296,N_17811);
nor U22480 (N_22480,N_17782,N_18239);
nand U22481 (N_22481,N_18598,N_18573);
xor U22482 (N_22482,N_18132,N_18364);
nand U22483 (N_22483,N_19934,N_19936);
xnor U22484 (N_22484,N_17851,N_18554);
or U22485 (N_22485,N_17971,N_19078);
or U22486 (N_22486,N_19091,N_17877);
and U22487 (N_22487,N_18792,N_19266);
or U22488 (N_22488,N_18807,N_19702);
and U22489 (N_22489,N_18015,N_18252);
or U22490 (N_22490,N_19942,N_18003);
and U22491 (N_22491,N_19855,N_19113);
and U22492 (N_22492,N_19325,N_18444);
nor U22493 (N_22493,N_18016,N_19892);
xor U22494 (N_22494,N_19902,N_17917);
and U22495 (N_22495,N_18790,N_19239);
or U22496 (N_22496,N_19303,N_19428);
or U22497 (N_22497,N_19142,N_19817);
and U22498 (N_22498,N_19131,N_19136);
or U22499 (N_22499,N_17984,N_18074);
nor U22500 (N_22500,N_20512,N_21183);
xnor U22501 (N_22501,N_21044,N_20671);
nand U22502 (N_22502,N_20128,N_21473);
xor U22503 (N_22503,N_21456,N_20100);
nor U22504 (N_22504,N_21233,N_20305);
or U22505 (N_22505,N_21595,N_20028);
nand U22506 (N_22506,N_22110,N_20034);
xor U22507 (N_22507,N_21737,N_20089);
nand U22508 (N_22508,N_21440,N_22035);
xnor U22509 (N_22509,N_20604,N_20590);
and U22510 (N_22510,N_21447,N_20229);
xnor U22511 (N_22511,N_20996,N_21139);
and U22512 (N_22512,N_21492,N_22150);
nand U22513 (N_22513,N_22442,N_21313);
or U22514 (N_22514,N_20791,N_21508);
nor U22515 (N_22515,N_20934,N_20209);
nand U22516 (N_22516,N_20396,N_21765);
or U22517 (N_22517,N_20851,N_21825);
nor U22518 (N_22518,N_21325,N_20634);
nor U22519 (N_22519,N_21503,N_20239);
nand U22520 (N_22520,N_22137,N_22472);
and U22521 (N_22521,N_22173,N_21471);
or U22522 (N_22522,N_20780,N_21498);
and U22523 (N_22523,N_21845,N_20811);
and U22524 (N_22524,N_20383,N_21510);
or U22525 (N_22525,N_20889,N_22389);
and U22526 (N_22526,N_20390,N_21267);
or U22527 (N_22527,N_21202,N_20092);
and U22528 (N_22528,N_21504,N_20877);
xor U22529 (N_22529,N_22046,N_20107);
nand U22530 (N_22530,N_20714,N_21703);
and U22531 (N_22531,N_22334,N_20806);
or U22532 (N_22532,N_21483,N_20730);
and U22533 (N_22533,N_20910,N_21063);
nand U22534 (N_22534,N_20621,N_20440);
xor U22535 (N_22535,N_20136,N_21236);
nand U22536 (N_22536,N_22380,N_21897);
xor U22537 (N_22537,N_21385,N_22415);
nand U22538 (N_22538,N_20000,N_21235);
or U22539 (N_22539,N_20443,N_22418);
or U22540 (N_22540,N_20564,N_20673);
xnor U22541 (N_22541,N_21232,N_22480);
or U22542 (N_22542,N_21931,N_22457);
nand U22543 (N_22543,N_21231,N_21149);
xnor U22544 (N_22544,N_21708,N_21197);
nand U22545 (N_22545,N_21328,N_21953);
nor U22546 (N_22546,N_22074,N_22305);
or U22547 (N_22547,N_21402,N_21570);
or U22548 (N_22548,N_20756,N_21962);
xor U22549 (N_22549,N_22090,N_21262);
nand U22550 (N_22550,N_21744,N_21212);
xor U22551 (N_22551,N_21283,N_20783);
nor U22552 (N_22552,N_21389,N_22177);
xnor U22553 (N_22553,N_20740,N_21830);
nand U22554 (N_22554,N_21653,N_20807);
nor U22555 (N_22555,N_20233,N_22080);
nor U22556 (N_22556,N_20678,N_20670);
xor U22557 (N_22557,N_22432,N_20257);
nand U22558 (N_22558,N_21330,N_20949);
nor U22559 (N_22559,N_21958,N_20118);
nand U22560 (N_22560,N_20700,N_22062);
and U22561 (N_22561,N_21700,N_20977);
or U22562 (N_22562,N_21843,N_20464);
nand U22563 (N_22563,N_20403,N_20758);
and U22564 (N_22564,N_20504,N_20148);
nand U22565 (N_22565,N_20494,N_21857);
nor U22566 (N_22566,N_21257,N_21869);
nor U22567 (N_22567,N_20063,N_21490);
nand U22568 (N_22568,N_21411,N_21917);
or U22569 (N_22569,N_21240,N_20820);
or U22570 (N_22570,N_20954,N_21655);
or U22571 (N_22571,N_20200,N_20695);
and U22572 (N_22572,N_20777,N_22373);
nor U22573 (N_22573,N_22321,N_20413);
xnor U22574 (N_22574,N_21156,N_20347);
nor U22575 (N_22575,N_22170,N_20058);
or U22576 (N_22576,N_20528,N_20854);
xnor U22577 (N_22577,N_20421,N_20732);
nand U22578 (N_22578,N_22214,N_21693);
and U22579 (N_22579,N_20081,N_20162);
nor U22580 (N_22580,N_22026,N_21896);
nor U22581 (N_22581,N_22422,N_20416);
nand U22582 (N_22582,N_20773,N_20880);
or U22583 (N_22583,N_20814,N_20753);
or U22584 (N_22584,N_20623,N_22447);
nor U22585 (N_22585,N_20252,N_22347);
or U22586 (N_22586,N_20916,N_21134);
xnor U22587 (N_22587,N_22015,N_21876);
nor U22588 (N_22588,N_21260,N_22149);
nor U22589 (N_22589,N_20800,N_20506);
nand U22590 (N_22590,N_21375,N_22124);
and U22591 (N_22591,N_20101,N_20462);
or U22592 (N_22592,N_20605,N_20618);
nor U22593 (N_22593,N_21996,N_20606);
or U22594 (N_22594,N_21726,N_20053);
and U22595 (N_22595,N_21000,N_22294);
nor U22596 (N_22596,N_21237,N_21647);
and U22597 (N_22597,N_21695,N_20307);
nor U22598 (N_22598,N_22135,N_20917);
and U22599 (N_22599,N_22461,N_21029);
or U22600 (N_22600,N_20398,N_21561);
or U22601 (N_22601,N_20550,N_20358);
and U22602 (N_22602,N_22220,N_22427);
nor U22603 (N_22603,N_21282,N_22444);
nand U22604 (N_22604,N_20833,N_20131);
xnor U22605 (N_22605,N_21716,N_20496);
and U22606 (N_22606,N_21436,N_20776);
nor U22607 (N_22607,N_20908,N_22290);
and U22608 (N_22608,N_21633,N_22104);
nor U22609 (N_22609,N_20223,N_20567);
nor U22610 (N_22610,N_21219,N_22082);
and U22611 (N_22611,N_21119,N_21192);
and U22612 (N_22612,N_21289,N_21999);
nand U22613 (N_22613,N_22333,N_20686);
nand U22614 (N_22614,N_21494,N_20304);
and U22615 (N_22615,N_20906,N_20692);
nor U22616 (N_22616,N_20277,N_20141);
or U22617 (N_22617,N_22190,N_21184);
nor U22618 (N_22618,N_22063,N_21667);
nand U22619 (N_22619,N_21345,N_21066);
and U22620 (N_22620,N_21381,N_21864);
and U22621 (N_22621,N_21438,N_20222);
xnor U22622 (N_22622,N_20580,N_20232);
or U22623 (N_22623,N_21548,N_20400);
or U22624 (N_22624,N_22358,N_22329);
or U22625 (N_22625,N_22235,N_21120);
nand U22626 (N_22626,N_22198,N_20386);
xnor U22627 (N_22627,N_20707,N_21244);
nand U22628 (N_22628,N_21264,N_22134);
or U22629 (N_22629,N_21762,N_20641);
or U22630 (N_22630,N_22208,N_21663);
nand U22631 (N_22631,N_21041,N_22429);
nor U22632 (N_22632,N_20351,N_21640);
nor U22633 (N_22633,N_21627,N_20153);
xor U22634 (N_22634,N_20765,N_22188);
xor U22635 (N_22635,N_22456,N_20620);
nand U22636 (N_22636,N_20006,N_21520);
xor U22637 (N_22637,N_21431,N_20407);
and U22638 (N_22638,N_21611,N_21446);
nand U22639 (N_22639,N_20940,N_20242);
and U22640 (N_22640,N_22205,N_20926);
xnor U22641 (N_22641,N_20346,N_22037);
and U22642 (N_22642,N_20023,N_21405);
nand U22643 (N_22643,N_21126,N_21565);
xnor U22644 (N_22644,N_20845,N_20380);
and U22645 (N_22645,N_21900,N_20899);
and U22646 (N_22646,N_21211,N_22322);
xnor U22647 (N_22647,N_20959,N_20744);
nand U22648 (N_22648,N_22230,N_22171);
xnor U22649 (N_22649,N_21851,N_21842);
nor U22650 (N_22650,N_20137,N_20286);
or U22651 (N_22651,N_20558,N_20873);
and U22652 (N_22652,N_21486,N_22040);
and U22653 (N_22653,N_21649,N_21168);
xor U22654 (N_22654,N_22196,N_21003);
and U22655 (N_22655,N_21977,N_20521);
or U22656 (N_22656,N_21318,N_21934);
or U22657 (N_22657,N_20344,N_20371);
or U22658 (N_22658,N_20608,N_22068);
nor U22659 (N_22659,N_22277,N_20037);
xor U22660 (N_22660,N_22255,N_21939);
or U22661 (N_22661,N_22440,N_20099);
nand U22662 (N_22662,N_20839,N_20560);
or U22663 (N_22663,N_21190,N_20062);
or U22664 (N_22664,N_20818,N_22095);
or U22665 (N_22665,N_20352,N_20936);
or U22666 (N_22666,N_20155,N_20706);
xor U22667 (N_22667,N_21948,N_21259);
nor U22668 (N_22668,N_22180,N_21828);
or U22669 (N_22669,N_22003,N_21204);
xnor U22670 (N_22670,N_21868,N_21092);
and U22671 (N_22671,N_22145,N_22218);
nand U22672 (N_22672,N_20029,N_21439);
nand U22673 (N_22673,N_21945,N_20696);
nor U22674 (N_22674,N_21174,N_22083);
or U22675 (N_22675,N_22278,N_21728);
or U22676 (N_22676,N_20507,N_20202);
and U22677 (N_22677,N_22211,N_21763);
and U22678 (N_22678,N_21861,N_21143);
nor U22679 (N_22679,N_20626,N_22477);
nor U22680 (N_22680,N_21847,N_21216);
xnor U22681 (N_22681,N_20527,N_20489);
nand U22682 (N_22682,N_21434,N_22401);
nand U22683 (N_22683,N_21449,N_20391);
nor U22684 (N_22684,N_22365,N_20828);
nor U22685 (N_22685,N_20600,N_21229);
or U22686 (N_22686,N_21954,N_22327);
nand U22687 (N_22687,N_21138,N_20822);
nand U22688 (N_22688,N_21821,N_21587);
or U22689 (N_22689,N_20685,N_22093);
xor U22690 (N_22690,N_20572,N_22437);
and U22691 (N_22691,N_21218,N_21902);
xnor U22692 (N_22692,N_21575,N_20184);
xor U22693 (N_22693,N_22379,N_22406);
xnor U22694 (N_22694,N_20984,N_22078);
and U22695 (N_22695,N_21337,N_20725);
and U22696 (N_22696,N_20636,N_21336);
and U22697 (N_22697,N_22405,N_22433);
xnor U22698 (N_22698,N_22317,N_20435);
nand U22699 (N_22699,N_21820,N_20312);
nor U22700 (N_22700,N_20441,N_21609);
nand U22701 (N_22701,N_21805,N_20804);
xnor U22702 (N_22702,N_22359,N_21136);
or U22703 (N_22703,N_20825,N_21493);
nor U22704 (N_22704,N_22451,N_21680);
nor U22705 (N_22705,N_20235,N_20942);
or U22706 (N_22706,N_22245,N_20759);
nor U22707 (N_22707,N_21038,N_20895);
xor U22708 (N_22708,N_20931,N_21031);
xor U22709 (N_22709,N_22029,N_21151);
or U22710 (N_22710,N_21108,N_22311);
and U22711 (N_22711,N_20970,N_20360);
xnor U22712 (N_22712,N_20088,N_21348);
xnor U22713 (N_22713,N_21109,N_22291);
or U22714 (N_22714,N_22320,N_21435);
nor U22715 (N_22715,N_21122,N_21578);
nor U22716 (N_22716,N_21555,N_20482);
nor U22717 (N_22717,N_21025,N_20071);
nand U22718 (N_22718,N_20104,N_22142);
nor U22719 (N_22719,N_21720,N_21601);
or U22720 (N_22720,N_21458,N_21266);
xnor U22721 (N_22721,N_20221,N_21974);
nand U22722 (N_22722,N_21055,N_20872);
nand U22723 (N_22723,N_21339,N_21919);
nand U22724 (N_22724,N_22497,N_21796);
xor U22725 (N_22725,N_20547,N_20569);
nor U22726 (N_22726,N_20473,N_22232);
nand U22727 (N_22727,N_21636,N_21321);
or U22728 (N_22728,N_21739,N_20332);
nor U22729 (N_22729,N_20296,N_22168);
and U22730 (N_22730,N_21497,N_20384);
nor U22731 (N_22731,N_22489,N_20268);
xnor U22732 (N_22732,N_21155,N_20893);
xor U22733 (N_22733,N_22324,N_21263);
nand U22734 (N_22734,N_21975,N_20587);
xnor U22735 (N_22735,N_21489,N_20331);
xor U22736 (N_22736,N_21074,N_22286);
xnor U22737 (N_22737,N_22425,N_20168);
nor U22738 (N_22738,N_21580,N_20329);
xor U22739 (N_22739,N_21514,N_20385);
xor U22740 (N_22740,N_22485,N_20042);
xnor U22741 (N_22741,N_22234,N_22079);
and U22742 (N_22742,N_21111,N_21172);
nand U22743 (N_22743,N_22166,N_21807);
or U22744 (N_22744,N_21697,N_22244);
and U22745 (N_22745,N_21512,N_21227);
nor U22746 (N_22746,N_20659,N_21735);
nor U22747 (N_22747,N_21024,N_20091);
nand U22748 (N_22748,N_20712,N_20579);
or U22749 (N_22749,N_22109,N_22355);
or U22750 (N_22750,N_21516,N_20105);
and U22751 (N_22751,N_20918,N_22096);
nor U22752 (N_22752,N_22413,N_21819);
or U22753 (N_22753,N_20985,N_21967);
or U22754 (N_22754,N_20291,N_21925);
and U22755 (N_22755,N_20717,N_20570);
nor U22756 (N_22756,N_21100,N_21065);
nand U22757 (N_22757,N_20836,N_20207);
or U22758 (N_22758,N_22225,N_20300);
nand U22759 (N_22759,N_22330,N_20502);
xor U22760 (N_22760,N_22416,N_21878);
nand U22761 (N_22761,N_22285,N_21463);
or U22762 (N_22762,N_21320,N_20317);
xor U22763 (N_22763,N_21563,N_22296);
or U22764 (N_22764,N_20561,N_20336);
and U22765 (N_22765,N_20874,N_20597);
xor U22766 (N_22766,N_20699,N_20905);
nor U22767 (N_22767,N_22383,N_20236);
xnor U22768 (N_22768,N_22038,N_22458);
or U22769 (N_22769,N_21681,N_21892);
or U22770 (N_22770,N_20026,N_21905);
nand U22771 (N_22771,N_20338,N_22275);
nor U22772 (N_22772,N_20613,N_22431);
and U22773 (N_22773,N_22131,N_20745);
nor U22774 (N_22774,N_22494,N_20907);
and U22775 (N_22775,N_21524,N_20897);
and U22776 (N_22776,N_20330,N_21152);
or U22777 (N_22777,N_20372,N_22010);
xor U22778 (N_22778,N_22346,N_21964);
and U22779 (N_22779,N_21009,N_21098);
or U22780 (N_22780,N_21288,N_20739);
nand U22781 (N_22781,N_20375,N_20333);
xnor U22782 (N_22782,N_20093,N_20077);
and U22783 (N_22783,N_20549,N_22197);
nor U22784 (N_22784,N_22319,N_21308);
nand U22785 (N_22785,N_20894,N_20963);
nor U22786 (N_22786,N_22008,N_21875);
nand U22787 (N_22787,N_20962,N_21077);
xor U22788 (N_22788,N_21064,N_21093);
and U22789 (N_22789,N_21421,N_21284);
xor U22790 (N_22790,N_20599,N_20399);
nand U22791 (N_22791,N_20174,N_21573);
nor U22792 (N_22792,N_21730,N_20001);
and U22793 (N_22793,N_20272,N_20869);
or U22794 (N_22794,N_21323,N_22222);
nand U22795 (N_22795,N_22268,N_21403);
and U22796 (N_22796,N_21200,N_21881);
nor U22797 (N_22797,N_20901,N_20812);
xnor U22798 (N_22798,N_20582,N_21075);
xor U22799 (N_22799,N_20120,N_21013);
nand U22800 (N_22800,N_21069,N_21599);
nor U22801 (N_22801,N_21956,N_21058);
nor U22802 (N_22802,N_21629,N_20929);
nor U22803 (N_22803,N_21993,N_21297);
xor U22804 (N_22804,N_21145,N_21027);
or U22805 (N_22805,N_21916,N_20716);
nor U22806 (N_22806,N_21099,N_20614);
xnor U22807 (N_22807,N_21544,N_21702);
nor U22808 (N_22808,N_22179,N_21793);
and U22809 (N_22809,N_20862,N_21005);
xnor U22810 (N_22810,N_22028,N_20679);
and U22811 (N_22811,N_22340,N_20896);
nor U22812 (N_22812,N_22479,N_21661);
and U22813 (N_22813,N_22376,N_20186);
nand U22814 (N_22814,N_20708,N_21026);
nor U22815 (N_22815,N_22438,N_21729);
xnor U22816 (N_22816,N_20958,N_21777);
nand U22817 (N_22817,N_21951,N_21180);
or U22818 (N_22818,N_20762,N_20838);
or U22819 (N_22819,N_20501,N_20941);
nand U22820 (N_22820,N_20288,N_20667);
nand U22821 (N_22821,N_21920,N_20420);
or U22822 (N_22822,N_21590,N_20302);
nor U22823 (N_22823,N_21388,N_21534);
nand U22824 (N_22824,N_21393,N_20159);
and U22825 (N_22825,N_20583,N_21105);
nand U22826 (N_22826,N_21969,N_21306);
nor U22827 (N_22827,N_22377,N_22146);
nor U22828 (N_22828,N_20735,N_21034);
or U22829 (N_22829,N_22192,N_22193);
nand U22830 (N_22830,N_20188,N_20713);
and U22831 (N_22831,N_22369,N_20316);
or U22832 (N_22832,N_21214,N_20556);
or U22833 (N_22833,N_20588,N_21015);
nor U22834 (N_22834,N_21983,N_22259);
nor U22835 (N_22835,N_21147,N_21530);
nor U22836 (N_22836,N_20596,N_22363);
nor U22837 (N_22837,N_20036,N_20244);
nand U22838 (N_22838,N_20051,N_21128);
nor U22839 (N_22839,N_21767,N_21946);
xnor U22840 (N_22840,N_20214,N_21314);
nor U22841 (N_22841,N_20925,N_21829);
and U22842 (N_22842,N_21252,N_20475);
nor U22843 (N_22843,N_22301,N_20827);
and U22844 (N_22844,N_20976,N_22167);
or U22845 (N_22845,N_20779,N_20943);
xor U22846 (N_22846,N_21274,N_22202);
and U22847 (N_22847,N_21322,N_22337);
or U22848 (N_22848,N_20546,N_21272);
nor U22849 (N_22849,N_21281,N_22044);
or U22850 (N_22850,N_20266,N_20370);
nand U22851 (N_22851,N_20010,N_22210);
xnor U22852 (N_22852,N_20313,N_20541);
and U22853 (N_22853,N_20289,N_20488);
nand U22854 (N_22854,N_20348,N_21541);
and U22855 (N_22855,N_22241,N_21791);
xor U22856 (N_22856,N_20427,N_22024);
xnor U22857 (N_22857,N_22120,N_21540);
nand U22858 (N_22858,N_20283,N_20944);
nand U22859 (N_22859,N_20160,N_21921);
and U22860 (N_22860,N_22470,N_20294);
nand U22861 (N_22861,N_21812,N_20350);
and U22862 (N_22862,N_21622,N_20785);
nor U22863 (N_22863,N_20412,N_21360);
xor U22864 (N_22864,N_22297,N_22140);
and U22865 (N_22865,N_20438,N_20871);
nand U22866 (N_22866,N_20228,N_21672);
and U22867 (N_22867,N_21273,N_22270);
xor U22868 (N_22868,N_20594,N_21602);
or U22869 (N_22869,N_22014,N_20457);
nor U22870 (N_22870,N_21460,N_22103);
or U22871 (N_22871,N_21850,N_22434);
nor U22872 (N_22872,N_20784,N_21338);
nor U22873 (N_22873,N_22036,N_22200);
xnor U22874 (N_22874,N_20491,N_20423);
and U22875 (N_22875,N_21344,N_21357);
xnor U22876 (N_22876,N_21811,N_22280);
or U22877 (N_22877,N_21226,N_20483);
or U22878 (N_22878,N_21674,N_22081);
or U22879 (N_22879,N_20477,N_21084);
or U22880 (N_22880,N_21641,N_20059);
nand U22881 (N_22881,N_20401,N_21893);
and U22882 (N_22882,N_21513,N_20829);
and U22883 (N_22883,N_20129,N_20852);
nor U22884 (N_22884,N_21201,N_21028);
and U22885 (N_22885,N_21890,N_21764);
or U22886 (N_22886,N_21331,N_20920);
nand U22887 (N_22887,N_22009,N_21732);
and U22888 (N_22888,N_21090,N_21943);
nand U22889 (N_22889,N_20287,N_21412);
nand U22890 (N_22890,N_22018,N_21371);
nand U22891 (N_22891,N_20526,N_20883);
nand U22892 (N_22892,N_20727,N_20094);
nor U22893 (N_22893,N_21186,N_22236);
or U22894 (N_22894,N_21255,N_21755);
xor U22895 (N_22895,N_22483,N_21210);
or U22896 (N_22896,N_21671,N_20284);
or U22897 (N_22897,N_21987,N_20853);
xor U22898 (N_22898,N_20267,N_21935);
or U22899 (N_22899,N_20308,N_21032);
nand U22900 (N_22900,N_21135,N_21746);
nor U22901 (N_22901,N_21205,N_20484);
nand U22902 (N_22902,N_20085,N_21007);
and U22903 (N_22903,N_21506,N_20250);
xor U22904 (N_22904,N_21877,N_22266);
xnor U22905 (N_22905,N_20553,N_20343);
or U22906 (N_22906,N_20449,N_21848);
nor U22907 (N_22907,N_21395,N_22315);
nand U22908 (N_22908,N_22257,N_21833);
or U22909 (N_22909,N_20922,N_20466);
nand U22910 (N_22910,N_21852,N_21740);
xor U22911 (N_22911,N_22227,N_21712);
or U22912 (N_22912,N_22426,N_22417);
and U22913 (N_22913,N_21675,N_21738);
xnor U22914 (N_22914,N_20103,N_20554);
nand U22915 (N_22915,N_20543,N_21023);
nand U22916 (N_22916,N_20075,N_21886);
nor U22917 (N_22917,N_21398,N_21078);
xnor U22918 (N_22918,N_21334,N_20049);
nand U22919 (N_22919,N_21907,N_21324);
or U22920 (N_22920,N_22341,N_21526);
xor U22921 (N_22921,N_20083,N_20589);
or U22922 (N_22922,N_20082,N_20365);
nand U22923 (N_22923,N_20956,N_20500);
or U22924 (N_22924,N_20536,N_21462);
or U22925 (N_22925,N_21269,N_20057);
xnor U22926 (N_22926,N_20480,N_20327);
xor U22927 (N_22927,N_21067,N_21639);
xor U22928 (N_22928,N_20662,N_20198);
nor U22929 (N_22929,N_21335,N_20715);
nor U22930 (N_22930,N_21124,N_20754);
xnor U22931 (N_22931,N_20231,N_20072);
nor U22932 (N_22932,N_21895,N_21731);
or U22933 (N_22933,N_22459,N_20404);
nand U22934 (N_22934,N_21170,N_21968);
or U22935 (N_22935,N_22246,N_20568);
nand U22936 (N_22936,N_20166,N_20486);
xnor U22937 (N_22937,N_20183,N_20324);
nand U22938 (N_22938,N_20180,N_20966);
and U22939 (N_22939,N_21553,N_20295);
xor U22940 (N_22940,N_21051,N_20681);
and U22941 (N_22941,N_21976,N_21824);
xor U22942 (N_22942,N_20345,N_20426);
nand U22943 (N_22943,N_20388,N_20455);
and U22944 (N_22944,N_20090,N_20980);
nor U22945 (N_22945,N_22248,N_20285);
nor U22946 (N_22946,N_20690,N_21300);
and U22947 (N_22947,N_21748,N_20009);
or U22948 (N_22948,N_22350,N_20971);
and U22949 (N_22949,N_21901,N_20591);
and U22950 (N_22950,N_21470,N_22007);
and U22951 (N_22951,N_20015,N_20911);
nor U22952 (N_22952,N_22141,N_20334);
xor U22953 (N_22953,N_20243,N_21814);
nand U22954 (N_22954,N_21118,N_20014);
nor U22955 (N_22955,N_21116,N_22474);
xor U22956 (N_22956,N_20193,N_21160);
and U22957 (N_22957,N_21474,N_20808);
nor U22958 (N_22958,N_20646,N_20326);
or U22959 (N_22959,N_21687,N_21991);
xor U22960 (N_22960,N_22371,N_20133);
or U22961 (N_22961,N_20353,N_21319);
or U22962 (N_22962,N_21496,N_22256);
and U22963 (N_22963,N_21176,N_21998);
and U22964 (N_22964,N_21428,N_20465);
and U22965 (N_22965,N_21188,N_20212);
and U22966 (N_22966,N_22282,N_20988);
xnor U22967 (N_22967,N_21567,N_22450);
and U22968 (N_22968,N_22191,N_21106);
xnor U22969 (N_22969,N_20781,N_21103);
xor U22970 (N_22970,N_22284,N_20790);
and U22971 (N_22971,N_21556,N_21607);
xor U22972 (N_22972,N_21046,N_21495);
nor U22973 (N_22973,N_21035,N_21608);
xnor U22974 (N_22974,N_20408,N_20511);
or U22975 (N_22975,N_21060,N_20628);
xnor U22976 (N_22976,N_21546,N_20045);
and U22977 (N_22977,N_22258,N_20601);
and U22978 (N_22978,N_21670,N_20602);
nor U22979 (N_22979,N_20282,N_21310);
and U22980 (N_22980,N_21642,N_20586);
nand U22981 (N_22981,N_22053,N_20691);
nor U22982 (N_22982,N_22430,N_21648);
nand U22983 (N_22983,N_20321,N_20824);
nor U22984 (N_22984,N_22332,N_22372);
nand U22985 (N_22985,N_20258,N_20146);
nor U22986 (N_22986,N_21760,N_21918);
xnor U22987 (N_22987,N_21299,N_20863);
nand U22988 (N_22988,N_21757,N_20719);
nor U22989 (N_22989,N_20428,N_20359);
nor U22990 (N_22990,N_20878,N_21140);
nor U22991 (N_22991,N_22254,N_20309);
or U22992 (N_22992,N_21794,N_21056);
nand U22993 (N_22993,N_22059,N_21042);
xor U22994 (N_22994,N_22027,N_22446);
xor U22995 (N_22995,N_22160,N_21963);
and U22996 (N_22996,N_21416,N_21157);
nand U22997 (N_22997,N_21261,N_20249);
nor U22998 (N_22998,N_21588,N_21409);
nand U22999 (N_22999,N_21685,N_20542);
nor U23000 (N_23000,N_20039,N_20796);
xnor U23001 (N_23001,N_22085,N_22264);
xnor U23002 (N_23002,N_21994,N_21898);
and U23003 (N_23003,N_22032,N_21761);
xor U23004 (N_23004,N_22408,N_20419);
or U23005 (N_23005,N_22001,N_21625);
nor U23006 (N_23006,N_21112,N_20616);
and U23007 (N_23007,N_21101,N_20932);
nor U23008 (N_23008,N_20322,N_21179);
xor U23009 (N_23009,N_21342,N_22482);
nand U23010 (N_23010,N_20415,N_20772);
nor U23011 (N_23011,N_21010,N_20454);
or U23012 (N_23012,N_21581,N_22449);
xnor U23013 (N_23013,N_22287,N_20179);
and U23014 (N_23014,N_21248,N_22123);
xor U23015 (N_23015,N_21756,N_20945);
nor U23016 (N_23016,N_21997,N_21882);
nand U23017 (N_23017,N_20782,N_20672);
and U23018 (N_23018,N_20111,N_20881);
xnor U23019 (N_23019,N_21694,N_20885);
and U23020 (N_23020,N_22387,N_21169);
and U23021 (N_23021,N_21538,N_21660);
and U23022 (N_23022,N_21624,N_20032);
and U23023 (N_23023,N_21924,N_20076);
xor U23024 (N_23024,N_21383,N_21933);
and U23025 (N_23025,N_22309,N_21096);
nor U23026 (N_23026,N_22157,N_21711);
and U23027 (N_23027,N_20933,N_22465);
and U23028 (N_23028,N_22049,N_20734);
nand U23029 (N_23029,N_22263,N_21018);
nand U23030 (N_23030,N_20342,N_20276);
nor U23031 (N_23031,N_21973,N_20904);
xnor U23032 (N_23032,N_20190,N_20434);
nor U23033 (N_23033,N_22323,N_20531);
or U23034 (N_23034,N_22165,N_21623);
xor U23035 (N_23035,N_21889,N_22384);
and U23036 (N_23036,N_21085,N_22155);
nor U23037 (N_23037,N_22331,N_21656);
nand U23038 (N_23038,N_21690,N_20020);
or U23039 (N_23039,N_20140,N_21144);
nor U23040 (N_23040,N_22033,N_20164);
or U23041 (N_23041,N_22325,N_22469);
or U23042 (N_23042,N_21254,N_21276);
xor U23043 (N_23043,N_20264,N_21666);
nand U23044 (N_23044,N_21426,N_22249);
xor U23045 (N_23045,N_20323,N_20581);
nand U23046 (N_23046,N_22342,N_21293);
nand U23047 (N_23047,N_21113,N_21367);
xnor U23048 (N_23048,N_22409,N_22176);
or U23049 (N_23049,N_22065,N_22119);
and U23050 (N_23050,N_20149,N_20157);
nor U23051 (N_23051,N_22388,N_20924);
or U23052 (N_23052,N_20930,N_20031);
or U23053 (N_23053,N_20640,N_20461);
xnor U23054 (N_23054,N_20135,N_20809);
and U23055 (N_23055,N_20612,N_21584);
nor U23056 (N_23056,N_20356,N_21246);
and U23057 (N_23057,N_21418,N_20968);
nand U23058 (N_23058,N_21453,N_21150);
and U23059 (N_23059,N_20281,N_21392);
xor U23060 (N_23060,N_21472,N_21121);
nor U23061 (N_23061,N_21558,N_20639);
and U23062 (N_23062,N_20802,N_20124);
nand U23063 (N_23063,N_20078,N_20156);
xnor U23064 (N_23064,N_22381,N_20701);
xor U23065 (N_23065,N_20532,N_22223);
xor U23066 (N_23066,N_22161,N_20098);
or U23067 (N_23067,N_22187,N_22186);
or U23068 (N_23068,N_20357,N_22126);
or U23069 (N_23069,N_20741,N_21709);
nand U23070 (N_23070,N_20151,N_21450);
and U23071 (N_23071,N_21592,N_21222);
nand U23072 (N_23072,N_21346,N_20913);
and U23073 (N_23073,N_21835,N_21941);
xor U23074 (N_23074,N_20525,N_20733);
nand U23075 (N_23075,N_20192,N_21662);
xor U23076 (N_23076,N_21872,N_20456);
or U23077 (N_23077,N_21505,N_20961);
and U23078 (N_23078,N_21195,N_21311);
nand U23079 (N_23079,N_20362,N_21130);
or U23080 (N_23080,N_20479,N_22060);
xor U23081 (N_23081,N_20064,N_20879);
or U23082 (N_23082,N_22056,N_20760);
nor U23083 (N_23083,N_21873,N_21658);
xnor U23084 (N_23084,N_20842,N_21596);
xor U23085 (N_23085,N_21836,N_20301);
nor U23086 (N_23086,N_21533,N_21487);
or U23087 (N_23087,N_22455,N_20247);
nand U23088 (N_23088,N_20948,N_20439);
xor U23089 (N_23089,N_21635,N_22127);
nor U23090 (N_23090,N_22138,N_20898);
or U23091 (N_23091,N_21822,N_21175);
xnor U23092 (N_23092,N_21786,N_21859);
nand U23093 (N_23093,N_20451,N_21250);
xor U23094 (N_23094,N_20215,N_21715);
and U23095 (N_23095,N_21097,N_21557);
nand U23096 (N_23096,N_20114,N_22339);
nor U23097 (N_23097,N_21380,N_21401);
and U23098 (N_23098,N_20577,N_20070);
nand U23099 (N_23099,N_22251,N_20850);
nor U23100 (N_23100,N_21193,N_22022);
xor U23101 (N_23101,N_21482,N_22113);
nor U23102 (N_23102,N_20723,N_21589);
xnor U23103 (N_23103,N_22058,N_22453);
nand U23104 (N_23104,N_21050,N_20251);
nand U23105 (N_23105,N_20424,N_20487);
xnor U23106 (N_23106,N_21048,N_21706);
nand U23107 (N_23107,N_20498,N_20805);
nor U23108 (N_23108,N_20847,N_21199);
or U23109 (N_23109,N_21718,N_22481);
or U23110 (N_23110,N_20478,N_21086);
or U23111 (N_23111,N_20722,N_21208);
and U23112 (N_23112,N_22094,N_20648);
or U23113 (N_23113,N_21692,N_21930);
xor U23114 (N_23114,N_20446,N_22398);
nor U23115 (N_23115,N_20130,N_21678);
xnor U23116 (N_23116,N_20445,N_20147);
or U23117 (N_23117,N_21950,N_22132);
nor U23118 (N_23118,N_22253,N_20866);
nor U23119 (N_23119,N_21354,N_21903);
or U23120 (N_23120,N_21659,N_21148);
nand U23121 (N_23121,N_21990,N_20655);
nor U23122 (N_23122,N_20684,N_20514);
nand U23123 (N_23123,N_21634,N_20306);
and U23124 (N_23124,N_22274,N_21185);
or U23125 (N_23125,N_20425,N_22492);
or U23126 (N_23126,N_22394,N_20084);
or U23127 (N_23127,N_20515,N_20658);
nor U23128 (N_23128,N_22215,N_20335);
and U23129 (N_23129,N_22112,N_20025);
xnor U23130 (N_23130,N_20683,N_20689);
nand U23131 (N_23131,N_22006,N_22072);
or U23132 (N_23132,N_21965,N_21107);
nand U23133 (N_23133,N_22017,N_20576);
nor U23134 (N_23134,N_20643,N_21970);
xor U23135 (N_23135,N_20065,N_20261);
nor U23136 (N_23136,N_21631,N_21879);
xor U23137 (N_23137,N_21089,N_21275);
nor U23138 (N_23138,N_20368,N_20429);
or U23139 (N_23139,N_21749,N_21909);
or U23140 (N_23140,N_21271,N_20038);
nor U23141 (N_23141,N_20736,N_21207);
or U23142 (N_23142,N_21509,N_20373);
and U23143 (N_23143,N_20680,N_20191);
nand U23144 (N_23144,N_21818,N_22139);
nand U23145 (N_23145,N_22463,N_22020);
xnor U23146 (N_23146,N_21955,N_21747);
and U23147 (N_23147,N_22421,N_20165);
or U23148 (N_23148,N_20593,N_20563);
and U23149 (N_23149,N_20876,N_20674);
or U23150 (N_23150,N_22092,N_21457);
nand U23151 (N_23151,N_21419,N_21384);
or U23152 (N_23152,N_20799,N_21464);
nor U23153 (N_23153,N_22393,N_21804);
nor U23154 (N_23154,N_21477,N_22283);
or U23155 (N_23155,N_20995,N_22075);
or U23156 (N_23156,N_21725,N_21479);
nor U23157 (N_23157,N_21080,N_22374);
nand U23158 (N_23158,N_21374,N_20774);
xor U23159 (N_23159,N_21583,N_21605);
xnor U23160 (N_23160,N_21979,N_21532);
or U23161 (N_23161,N_21936,N_21724);
xnor U23162 (N_23162,N_22195,N_22100);
or U23163 (N_23163,N_21571,N_20069);
nor U23164 (N_23164,N_20865,N_21645);
nand U23165 (N_23165,N_22021,N_20374);
nand U23166 (N_23166,N_21292,N_22288);
nor U23167 (N_23167,N_20769,N_22367);
or U23168 (N_23168,N_21673,N_21683);
and U23169 (N_23169,N_21177,N_20764);
or U23170 (N_23170,N_20697,N_21020);
and U23171 (N_23171,N_21350,N_20253);
xnor U23172 (N_23172,N_20468,N_22064);
nor U23173 (N_23173,N_22395,N_22084);
or U23174 (N_23174,N_22087,N_22302);
and U23175 (N_23175,N_22041,N_22343);
or U23176 (N_23176,N_20102,N_21410);
xor U23177 (N_23177,N_20019,N_20437);
nand U23178 (N_23178,N_21874,N_21072);
and U23179 (N_23179,N_20002,N_20219);
nand U23180 (N_23180,N_22069,N_21911);
and U23181 (N_23181,N_20048,N_21234);
and U23182 (N_23182,N_21727,N_22423);
nor U23183 (N_23183,N_22219,N_21628);
xnor U23184 (N_23184,N_20194,N_20068);
and U23185 (N_23185,N_21417,N_20378);
nor U23186 (N_23186,N_21572,N_21995);
nand U23187 (N_23187,N_22493,N_21733);
nand U23188 (N_23188,N_22011,N_21088);
nor U23189 (N_23189,N_20044,N_22169);
nor U23190 (N_23190,N_20185,N_21539);
or U23191 (N_23191,N_21430,N_21928);
and U23192 (N_23192,N_20397,N_20537);
xnor U23193 (N_23193,N_20566,N_22368);
nand U23194 (N_23194,N_20255,N_21826);
nor U23195 (N_23195,N_21569,N_21278);
and U23196 (N_23196,N_21316,N_22496);
or U23197 (N_23197,N_21853,N_21688);
or U23198 (N_23198,N_20645,N_20973);
and U23199 (N_23199,N_22025,N_21363);
nor U23200 (N_23200,N_20798,N_21249);
and U23201 (N_23201,N_22498,N_21043);
nor U23202 (N_23202,N_21413,N_21209);
or U23203 (N_23203,N_21832,N_21163);
xnor U23204 (N_23204,N_20414,N_20990);
or U23205 (N_23205,N_21855,N_22484);
nor U23206 (N_23206,N_22050,N_22047);
nand U23207 (N_23207,N_21871,N_21082);
nand U23208 (N_23208,N_20485,N_20615);
nand U23209 (N_23209,N_21582,N_20801);
and U23210 (N_23210,N_21059,N_20652);
or U23211 (N_23211,N_21591,N_21433);
nor U23212 (N_23212,N_21593,N_20238);
or U23213 (N_23213,N_21543,N_21361);
and U23214 (N_23214,N_20819,N_21932);
nand U23215 (N_23215,N_20139,N_22111);
or U23216 (N_23216,N_21554,N_22156);
nand U23217 (N_23217,N_20173,N_22107);
xor U23218 (N_23218,N_21391,N_21296);
nor U23219 (N_23219,N_21597,N_21287);
nor U23220 (N_23220,N_21870,N_22115);
and U23221 (N_23221,N_22091,N_22242);
nor U23222 (N_23222,N_21362,N_20275);
xnor U23223 (N_23223,N_21988,N_21722);
xor U23224 (N_23224,N_22108,N_20227);
nand U23225 (N_23225,N_21723,N_20022);
xnor U23226 (N_23226,N_20530,N_20571);
nand U23227 (N_23227,N_22229,N_21441);
or U23228 (N_23228,N_20050,N_20016);
or U23229 (N_23229,N_20047,N_22262);
nand U23230 (N_23230,N_20458,N_22077);
nand U23231 (N_23231,N_20831,N_20928);
or U23232 (N_23232,N_21341,N_21689);
nand U23233 (N_23233,N_22159,N_21914);
and U23234 (N_23234,N_22269,N_21049);
and U23235 (N_23235,N_22039,N_20143);
nor U23236 (N_23236,N_22441,N_20467);
and U23237 (N_23237,N_20260,N_20240);
xor U23238 (N_23238,N_20533,N_20548);
xor U23239 (N_23239,N_20816,N_20340);
and U23240 (N_23240,N_22265,N_20742);
xor U23241 (N_23241,N_20849,N_21182);
nand U23242 (N_23242,N_20813,N_20534);
or U23243 (N_23243,N_21251,N_22105);
nand U23244 (N_23244,N_21676,N_21942);
nand U23245 (N_23245,N_21125,N_20389);
and U23246 (N_23246,N_21952,N_21579);
or U23247 (N_23247,N_20121,N_21837);
and U23248 (N_23248,N_20199,N_20109);
nor U23249 (N_23249,N_22443,N_21795);
nor U23250 (N_23250,N_21775,N_20859);
xor U23251 (N_23251,N_20460,N_20205);
xor U23252 (N_23252,N_20524,N_22310);
and U23253 (N_23253,N_21815,N_21522);
nand U23254 (N_23254,N_21620,N_20704);
nand U23255 (N_23255,N_20017,N_22098);
xor U23256 (N_23256,N_20676,N_21650);
xor U23257 (N_23257,N_21785,N_22175);
nand U23258 (N_23258,N_22335,N_21253);
xnor U23259 (N_23259,N_22048,N_21131);
and U23260 (N_23260,N_20766,N_20220);
and U23261 (N_23261,N_20108,N_21265);
nand U23262 (N_23262,N_22164,N_22000);
nand U23263 (N_23263,N_22231,N_20861);
xnor U23264 (N_23264,N_20430,N_22306);
or U23265 (N_23265,N_20259,N_21223);
xnor U23266 (N_23266,N_21912,N_22207);
or U23267 (N_23267,N_22128,N_22271);
xnor U23268 (N_23268,N_22239,N_20463);
xnor U23269 (N_23269,N_20792,N_21637);
xor U23270 (N_23270,N_21586,N_22392);
xnor U23271 (N_23271,N_20448,N_21258);
nor U23272 (N_23272,N_20060,N_20731);
or U23273 (N_23273,N_22414,N_20024);
or U23274 (N_23274,N_21566,N_20562);
and U23275 (N_23275,N_21420,N_22261);
nor U23276 (N_23276,N_21545,N_21682);
or U23277 (N_23277,N_20142,N_21887);
xor U23278 (N_23278,N_21386,N_20953);
or U23279 (N_23279,N_21036,N_20919);
nor U23280 (N_23280,N_20355,N_22314);
nor U23281 (N_23281,N_22439,N_20939);
or U23282 (N_23282,N_21159,N_21929);
nor U23283 (N_23283,N_21792,N_20538);
or U23284 (N_23284,N_20273,N_21856);
nor U23285 (N_23285,N_20902,N_20575);
nor U23286 (N_23286,N_21745,N_20982);
and U23287 (N_23287,N_20718,N_21070);
xor U23288 (N_23288,N_20339,N_20172);
nand U23289 (N_23289,N_22348,N_20422);
or U23290 (N_23290,N_20767,N_22300);
and U23291 (N_23291,N_21782,N_21831);
xnor U23292 (N_23292,N_21443,N_21884);
xnor U23293 (N_23293,N_21705,N_22133);
xnor U23294 (N_23294,N_20490,N_22016);
xor U23295 (N_23295,N_20771,N_21630);
xnor U23296 (N_23296,N_22247,N_21638);
nor U23297 (N_23297,N_20974,N_22410);
nor U23298 (N_23298,N_22102,N_22201);
and U23299 (N_23299,N_21221,N_21617);
or U23300 (N_23300,N_21699,N_22448);
nand U23301 (N_23301,N_22354,N_20787);
and U23302 (N_23302,N_20433,N_20382);
nor U23303 (N_23303,N_21802,N_20544);
nor U23304 (N_23304,N_20794,N_21858);
and U23305 (N_23305,N_21158,N_20208);
or U23306 (N_23306,N_20752,N_21511);
xor U23307 (N_23307,N_22125,N_20709);
or U23308 (N_23308,N_21146,N_20960);
or U23309 (N_23309,N_20848,N_21390);
nor U23310 (N_23310,N_22385,N_21030);
nand U23311 (N_23311,N_21270,N_22152);
nor U23312 (N_23312,N_20256,N_21247);
nand U23313 (N_23313,N_20888,N_20748);
and U23314 (N_23314,N_21091,N_22204);
and U23315 (N_23315,N_22353,N_20837);
nand U23316 (N_23316,N_20644,N_20592);
nand U23317 (N_23317,N_21986,N_20314);
nor U23318 (N_23318,N_22391,N_20868);
nor U23319 (N_23319,N_21603,N_22351);
xor U23320 (N_23320,N_20021,N_21004);
or U23321 (N_23321,N_22464,N_20218);
and U23322 (N_23322,N_20432,N_21332);
nand U23323 (N_23323,N_21710,N_20993);
or U23324 (N_23324,N_21359,N_20923);
nor U23325 (N_23325,N_20262,N_21781);
nor U23326 (N_23326,N_21652,N_20650);
nor U23327 (N_23327,N_21776,N_21376);
nand U23328 (N_23328,N_22276,N_20112);
and U23329 (N_23329,N_21340,N_20005);
or U23330 (N_23330,N_20720,N_20823);
nor U23331 (N_23331,N_20617,N_20061);
nor U23332 (N_23332,N_21600,N_21957);
or U23333 (N_23333,N_20710,N_20751);
nand U23334 (N_23334,N_22424,N_22370);
nor U23335 (N_23335,N_21153,N_21329);
or U23336 (N_23336,N_20786,N_20635);
and U23337 (N_23337,N_21537,N_20937);
nor U23338 (N_23338,N_20043,N_20138);
or U23339 (N_23339,N_21165,N_20217);
nor U23340 (N_23340,N_21432,N_21860);
and U23341 (N_23341,N_20517,N_22435);
and U23342 (N_23342,N_21230,N_20263);
and U23343 (N_23343,N_21774,N_21424);
nand U23344 (N_23344,N_20211,N_21651);
or U23345 (N_23345,N_20497,N_21527);
xnor U23346 (N_23346,N_22316,N_21669);
nand U23347 (N_23347,N_22194,N_20054);
nor U23348 (N_23348,N_21286,N_20290);
nor U23349 (N_23349,N_20903,N_20299);
nor U23350 (N_23350,N_21326,N_21817);
nor U23351 (N_23351,N_21437,N_20349);
or U23352 (N_23352,N_22466,N_22181);
nand U23353 (N_23353,N_22228,N_20499);
nor U23354 (N_23354,N_21206,N_20665);
nor U23355 (N_23355,N_20201,N_20459);
or U23356 (N_23356,N_20341,N_21913);
or U23357 (N_23357,N_21215,N_22212);
xnor U23358 (N_23358,N_21379,N_21277);
or U23359 (N_23359,N_20206,N_21961);
nor U23360 (N_23360,N_20999,N_21422);
or U23361 (N_23361,N_20167,N_22488);
nor U23362 (N_23362,N_22289,N_21488);
nand U23363 (N_23363,N_20858,N_20318);
nand U23364 (N_23364,N_21110,N_21132);
nand U23365 (N_23365,N_21002,N_22312);
nor U23366 (N_23366,N_20637,N_20171);
or U23367 (N_23367,N_20551,N_22144);
and U23368 (N_23368,N_21501,N_20698);
and U23369 (N_23369,N_21577,N_20666);
nor U23370 (N_23370,N_20325,N_21621);
nor U23371 (N_23371,N_22397,N_21525);
or U23372 (N_23372,N_20216,N_21810);
or U23373 (N_23373,N_20163,N_22486);
nor U23374 (N_23374,N_20856,N_21838);
xnor U23375 (N_23375,N_21467,N_22318);
xor U23376 (N_23376,N_21940,N_20609);
or U23377 (N_23377,N_20187,N_21846);
nor U23378 (N_23378,N_21937,N_21461);
xnor U23379 (N_23379,N_20320,N_21542);
nand U23380 (N_23380,N_20481,N_20870);
nand U23381 (N_23381,N_22386,N_21515);
and U23382 (N_23382,N_20074,N_21366);
nand U23383 (N_23383,N_20030,N_20292);
or U23384 (N_23384,N_20447,N_22076);
and U23385 (N_23385,N_21268,N_21327);
nor U23386 (N_23386,N_21840,N_22034);
and U23387 (N_23387,N_21806,N_21549);
nand U23388 (N_23388,N_21312,N_21445);
nor U23389 (N_23389,N_21079,N_21618);
or U23390 (N_23390,N_22468,N_21162);
xor U23391 (N_23391,N_21228,N_20195);
xnor U23392 (N_23392,N_20529,N_21011);
xor U23393 (N_23393,N_22005,N_21619);
xnor U23394 (N_23394,N_21614,N_21938);
or U23395 (N_23395,N_20702,N_20226);
or U23396 (N_23396,N_21750,N_21280);
or U23397 (N_23397,N_22293,N_21904);
xnor U23398 (N_23398,N_21307,N_20585);
and U23399 (N_23399,N_20270,N_20040);
nand U23400 (N_23400,N_20337,N_20927);
xnor U23401 (N_23401,N_21016,N_21704);
nor U23402 (N_23402,N_21915,N_20152);
and U23403 (N_23403,N_22303,N_21425);
or U23404 (N_23404,N_21455,N_21369);
or U23405 (N_23405,N_21164,N_21094);
xnor U23406 (N_23406,N_20315,N_22336);
xnor U23407 (N_23407,N_21001,N_20117);
xnor U23408 (N_23408,N_20890,N_21076);
and U23409 (N_23409,N_20046,N_20864);
nor U23410 (N_23410,N_21243,N_20834);
and U23411 (N_23411,N_22174,N_21372);
nand U23412 (N_23412,N_22013,N_20768);
and U23413 (N_23413,N_21017,N_20688);
or U23414 (N_23414,N_20633,N_21423);
nand U23415 (N_23415,N_20097,N_21459);
nand U23416 (N_23416,N_20393,N_20778);
and U23417 (N_23417,N_21397,N_21037);
and U23418 (N_23418,N_21751,N_21491);
nand U23419 (N_23419,N_22121,N_20469);
nor U23420 (N_23420,N_21071,N_20274);
nor U23421 (N_23421,N_21813,N_21137);
nand U23422 (N_23422,N_22252,N_21220);
and U23423 (N_23423,N_21191,N_20381);
xnor U23424 (N_23424,N_21414,N_22185);
xnor U23425 (N_23425,N_21519,N_20743);
xnor U23426 (N_23426,N_21377,N_21081);
or U23427 (N_23427,N_21536,N_21910);
and U23428 (N_23428,N_21568,N_21294);
nand U23429 (N_23429,N_22452,N_21839);
or U23430 (N_23430,N_22445,N_20642);
xor U23431 (N_23431,N_20509,N_20442);
and U23432 (N_23432,N_20915,N_22403);
and U23433 (N_23433,N_21368,N_20630);
or U23434 (N_23434,N_20610,N_20994);
nor U23435 (N_23435,N_21052,N_21415);
nand U23436 (N_23436,N_22238,N_20354);
nor U23437 (N_23437,N_21550,N_20660);
or U23438 (N_23438,N_21798,N_20935);
or U23439 (N_23439,N_20826,N_22475);
and U23440 (N_23440,N_21985,N_22066);
and U23441 (N_23441,N_21452,N_21500);
and U23442 (N_23442,N_21396,N_21626);
nand U23443 (N_23443,N_20510,N_21816);
nand U23444 (N_23444,N_20964,N_20657);
xor U23445 (N_23445,N_21285,N_20298);
xor U23446 (N_23446,N_20409,N_20711);
xnor U23447 (N_23447,N_21758,N_21133);
xnor U23448 (N_23448,N_22183,N_21507);
or U23449 (N_23449,N_20573,N_20520);
xnor U23450 (N_23450,N_21803,N_21574);
and U23451 (N_23451,N_20557,N_21644);
nor U23452 (N_23452,N_21742,N_22476);
nor U23453 (N_23453,N_22061,N_20677);
xor U23454 (N_23454,N_22399,N_22428);
nor U23455 (N_23455,N_21612,N_20611);
nor U23456 (N_23456,N_21894,N_20492);
or U23457 (N_23457,N_21632,N_20377);
nand U23458 (N_23458,N_20418,N_21104);
or U23459 (N_23459,N_20417,N_22390);
xnor U23460 (N_23460,N_20649,N_20867);
nor U23461 (N_23461,N_21714,N_21187);
nor U23462 (N_23462,N_20729,N_22055);
nor U23463 (N_23463,N_20841,N_21333);
xor U23464 (N_23464,N_20855,N_21006);
xnor U23465 (N_23465,N_20675,N_21189);
nor U23466 (N_23466,N_20246,N_20625);
or U23467 (N_23467,N_20559,N_20979);
or U23468 (N_23468,N_21779,N_20952);
nor U23469 (N_23469,N_21387,N_20875);
or U23470 (N_23470,N_20476,N_20726);
or U23471 (N_23471,N_20033,N_21604);
and U23472 (N_23472,N_21980,N_20366);
and U23473 (N_23473,N_20411,N_20607);
xor U23474 (N_23474,N_20682,N_21073);
xnor U23475 (N_23475,N_20815,N_21684);
nor U23476 (N_23476,N_21053,N_20987);
or U23477 (N_23477,N_20651,N_20474);
or U23478 (N_23478,N_20254,N_20471);
nand U23479 (N_23479,N_20087,N_20603);
or U23480 (N_23480,N_20176,N_21834);
nand U23481 (N_23481,N_21485,N_22499);
nand U23482 (N_23482,N_21305,N_21129);
xnor U23483 (N_23483,N_20394,N_20303);
xnor U23484 (N_23484,N_21279,N_20797);
and U23485 (N_23485,N_20297,N_20882);
nand U23486 (N_23486,N_20189,N_20125);
xor U23487 (N_23487,N_21734,N_22362);
or U23488 (N_23488,N_21780,N_22364);
or U23489 (N_23489,N_20452,N_21679);
xor U23490 (N_23490,N_22136,N_21476);
nor U23491 (N_23491,N_20008,N_20664);
nor U23492 (N_23492,N_20169,N_20055);
and U23493 (N_23493,N_20132,N_21789);
or U23494 (N_23494,N_20013,N_22298);
nand U23495 (N_23495,N_21743,N_21173);
nand U23496 (N_23496,N_20997,N_21719);
nand U23497 (N_23497,N_21499,N_20840);
nor U23498 (N_23498,N_21347,N_22178);
xnor U23499 (N_23499,N_21444,N_21349);
and U23500 (N_23500,N_22147,N_21518);
or U23501 (N_23501,N_20110,N_20271);
and U23502 (N_23502,N_20379,N_20011);
nor U23503 (N_23503,N_20978,N_20361);
or U23504 (N_23504,N_20018,N_21899);
nand U23505 (N_23505,N_20598,N_21213);
nor U23506 (N_23506,N_21922,N_21484);
xor U23507 (N_23507,N_21057,N_21068);
nand U23508 (N_23508,N_21429,N_20788);
nor U23509 (N_23509,N_22478,N_21800);
nand U23510 (N_23510,N_21783,N_20123);
or U23511 (N_23511,N_21400,N_21972);
and U23512 (N_23512,N_20950,N_22184);
or U23513 (N_23513,N_21142,N_22143);
and U23514 (N_23514,N_20810,N_20967);
nand U23515 (N_23515,N_20749,N_21238);
nor U23516 (N_23516,N_22490,N_20981);
nor U23517 (N_23517,N_21117,N_20761);
xnor U23518 (N_23518,N_21242,N_20280);
nor U23519 (N_23519,N_22419,N_21290);
and U23520 (N_23520,N_22151,N_21022);
nand U23521 (N_23521,N_22400,N_21468);
nor U23522 (N_23522,N_21862,N_21301);
nor U23523 (N_23523,N_20086,N_21454);
xnor U23524 (N_23524,N_20969,N_21245);
xnor U23525 (N_23525,N_20402,N_22117);
nand U23526 (N_23526,N_20724,N_20545);
or U23527 (N_23527,N_22471,N_20746);
and U23528 (N_23528,N_22012,N_20663);
nor U23529 (N_23529,N_22213,N_21885);
nor U23530 (N_23530,N_22054,N_22382);
and U23531 (N_23531,N_20584,N_20067);
or U23532 (N_23532,N_20909,N_22002);
nand U23533 (N_23533,N_21665,N_21521);
nand U23534 (N_23534,N_20886,N_20096);
or U23535 (N_23535,N_21033,N_21809);
or U23536 (N_23536,N_21298,N_20027);
nand U23537 (N_23537,N_20269,N_21469);
or U23538 (N_23538,N_20134,N_20972);
nand U23539 (N_23539,N_20738,N_21014);
xnor U23540 (N_23540,N_22101,N_21295);
or U23541 (N_23541,N_21373,N_21535);
or U23542 (N_23542,N_21529,N_22043);
nor U23543 (N_23543,N_21949,N_21768);
or U23544 (N_23544,N_21823,N_21309);
nor U23545 (N_23545,N_21351,N_21047);
xor U23546 (N_23546,N_21196,N_20319);
and U23547 (N_23547,N_20860,N_21167);
xor U23548 (N_23548,N_20364,N_22057);
xnor U23549 (N_23549,N_21923,N_21291);
or U23550 (N_23550,N_22114,N_20647);
xor U23551 (N_23551,N_20376,N_21466);
and U23552 (N_23552,N_21598,N_22158);
or U23553 (N_23553,N_22243,N_21528);
nor U23554 (N_23554,N_22129,N_21203);
xnor U23555 (N_23555,N_20835,N_21754);
nor U23556 (N_23556,N_22404,N_20056);
xor U23557 (N_23557,N_22071,N_20007);
xor U23558 (N_23558,N_21039,N_22130);
nor U23559 (N_23559,N_21766,N_22070);
nand U23560 (N_23560,N_21613,N_21008);
or U23561 (N_23561,N_20750,N_21303);
or U23562 (N_23562,N_20203,N_20832);
or U23563 (N_23563,N_22118,N_22420);
nand U23564 (N_23564,N_20161,N_21606);
nor U23565 (N_23565,N_22240,N_22199);
xor U23566 (N_23566,N_20122,N_21404);
xnor U23567 (N_23567,N_20126,N_21194);
or U23568 (N_23568,N_20310,N_20113);
and U23569 (N_23569,N_20230,N_20369);
xnor U23570 (N_23570,N_20622,N_20817);
nand U23571 (N_23571,N_21906,N_21698);
xnor U23572 (N_23572,N_20627,N_21061);
and U23573 (N_23573,N_21616,N_21981);
nor U23574 (N_23574,N_22154,N_22436);
or U23575 (N_23575,N_20279,N_21547);
nor U23576 (N_23576,N_21442,N_21615);
and U23577 (N_23577,N_21773,N_21713);
or U23578 (N_23578,N_21161,N_20450);
or U23579 (N_23579,N_22073,N_22281);
xnor U23580 (N_23580,N_21888,N_21304);
or U23581 (N_23581,N_21095,N_21115);
and U23582 (N_23582,N_22412,N_20182);
nor U23583 (N_23583,N_20755,N_21102);
nand U23584 (N_23584,N_20793,N_21531);
and U23585 (N_23585,N_20119,N_21256);
or U23586 (N_23586,N_20947,N_22148);
or U23587 (N_23587,N_22473,N_20410);
and U23588 (N_23588,N_22106,N_21378);
xnor U23589 (N_23589,N_21891,N_20565);
xnor U23590 (N_23590,N_22217,N_21171);
and U23591 (N_23591,N_20012,N_20505);
and U23592 (N_23592,N_21480,N_21664);
or U23593 (N_23593,N_22051,N_20693);
nand U23594 (N_23594,N_21562,N_22260);
nand U23595 (N_23595,N_21394,N_21551);
and U23596 (N_23596,N_22162,N_20946);
and U23597 (N_23597,N_20293,N_20004);
xnor U23598 (N_23598,N_21564,N_20387);
nand U23599 (N_23599,N_22338,N_20516);
and U23600 (N_23600,N_21696,N_21944);
and U23601 (N_23601,N_20552,N_21370);
and U23602 (N_23602,N_20975,N_20770);
xor U23603 (N_23603,N_21677,N_20080);
nand U23604 (N_23604,N_20631,N_20619);
and U23605 (N_23605,N_22182,N_22487);
or U23606 (N_23606,N_22307,N_20694);
nand U23607 (N_23607,N_20405,N_20181);
and U23608 (N_23608,N_21040,N_20983);
xor U23609 (N_23609,N_20115,N_20127);
nand U23610 (N_23610,N_20957,N_22295);
and U23611 (N_23611,N_20955,N_20278);
or U23612 (N_23612,N_20436,N_20629);
and U23613 (N_23613,N_21769,N_22226);
or U23614 (N_23614,N_21239,N_21866);
nand U23615 (N_23615,N_20470,N_21523);
and U23616 (N_23616,N_20921,N_21478);
or U23617 (N_23617,N_20406,N_20066);
and U23618 (N_23618,N_22216,N_22031);
or U23619 (N_23619,N_22352,N_20992);
nor U23620 (N_23620,N_22460,N_21114);
or U23621 (N_23621,N_20495,N_21691);
xnor U23622 (N_23622,N_21741,N_21087);
nor U23623 (N_23623,N_21865,N_22375);
nand U23624 (N_23624,N_21517,N_22088);
and U23625 (N_23625,N_22221,N_20654);
xnor U23626 (N_23626,N_21083,N_22019);
xor U23627 (N_23627,N_20311,N_21654);
and U23628 (N_23628,N_20803,N_22237);
nor U23629 (N_23629,N_20965,N_21984);
nand U23630 (N_23630,N_20653,N_20241);
xor U23631 (N_23631,N_20444,N_20518);
or U23632 (N_23632,N_22023,N_20196);
and U23633 (N_23633,N_22099,N_20737);
and U23634 (N_23634,N_21302,N_22267);
nand U23635 (N_23635,N_21123,N_22360);
nor U23636 (N_23636,N_20523,N_22042);
nand U23637 (N_23637,N_21908,N_20900);
nor U23638 (N_23638,N_21982,N_21753);
and U23639 (N_23639,N_20846,N_20225);
and U23640 (N_23640,N_20843,N_20912);
nand U23641 (N_23641,N_20892,N_20248);
or U23642 (N_23642,N_20991,N_20453);
nand U23643 (N_23643,N_21686,N_21045);
or U23644 (N_23644,N_20224,N_21867);
and U23645 (N_23645,N_21224,N_21926);
xnor U23646 (N_23646,N_21560,N_22328);
xor U23647 (N_23647,N_21166,N_22272);
nand U23648 (N_23648,N_20757,N_20245);
xnor U23649 (N_23649,N_21849,N_21315);
nand U23650 (N_23650,N_20150,N_22304);
and U23651 (N_23651,N_21827,N_21759);
nand U23652 (N_23652,N_21552,N_20669);
nor U23653 (N_23653,N_21054,N_22313);
nor U23654 (N_23654,N_20503,N_21610);
xor U23655 (N_23655,N_20116,N_20951);
nor U23656 (N_23656,N_22052,N_20938);
nor U23657 (N_23657,N_21844,N_21966);
xnor U23658 (N_23658,N_20632,N_22411);
or U23659 (N_23659,N_22273,N_21971);
xor U23660 (N_23660,N_21481,N_22224);
and U23661 (N_23661,N_21019,N_21225);
nand U23662 (N_23662,N_21356,N_20392);
and U23663 (N_23663,N_20237,N_21752);
nand U23664 (N_23664,N_20687,N_20431);
xnor U23665 (N_23665,N_21797,N_21127);
or U23666 (N_23666,N_20539,N_22086);
and U23667 (N_23667,N_22378,N_21355);
nor U23668 (N_23668,N_22163,N_21643);
and U23669 (N_23669,N_21198,N_20795);
nor U23670 (N_23670,N_20705,N_21778);
and U23671 (N_23671,N_22067,N_20035);
or U23672 (N_23672,N_21668,N_22407);
nor U23673 (N_23673,N_21451,N_20210);
and U23674 (N_23674,N_21841,N_22344);
and U23675 (N_23675,N_20775,N_21448);
nor U23676 (N_23676,N_21790,N_21989);
nor U23677 (N_23677,N_21784,N_20519);
or U23678 (N_23678,N_22030,N_20891);
xor U23679 (N_23679,N_21576,N_21358);
nand U23680 (N_23680,N_22396,N_21365);
nand U23681 (N_23681,N_20213,N_22172);
nand U23682 (N_23682,N_20106,N_20508);
nand U23683 (N_23683,N_22345,N_21883);
xor U23684 (N_23684,N_20513,N_22250);
and U23685 (N_23685,N_22454,N_20721);
or U23686 (N_23686,N_21012,N_22122);
nand U23687 (N_23687,N_20763,N_20363);
nor U23688 (N_23688,N_20747,N_21717);
xnor U23689 (N_23689,N_22004,N_20493);
nand U23690 (N_23690,N_21657,N_20095);
nor U23691 (N_23691,N_22366,N_22089);
xor U23692 (N_23692,N_20998,N_21408);
nor U23693 (N_23693,N_20703,N_21154);
nand U23694 (N_23694,N_22357,N_22361);
nand U23695 (N_23695,N_20328,N_21788);
or U23696 (N_23696,N_20158,N_22402);
and U23697 (N_23697,N_21808,N_20522);
nand U23698 (N_23698,N_21217,N_22116);
or U23699 (N_23699,N_20830,N_21927);
nand U23700 (N_23700,N_20887,N_21407);
nor U23701 (N_23701,N_21863,N_20170);
or U23702 (N_23702,N_20540,N_21947);
or U23703 (N_23703,N_21594,N_20472);
nand U23704 (N_23704,N_21364,N_20789);
xnor U23705 (N_23705,N_20052,N_21343);
or U23706 (N_23706,N_21646,N_20177);
or U23707 (N_23707,N_21701,N_22233);
and U23708 (N_23708,N_20989,N_22356);
and U23709 (N_23709,N_20367,N_20395);
nor U23710 (N_23710,N_20914,N_20857);
nand U23711 (N_23711,N_22203,N_21399);
xor U23712 (N_23712,N_21317,N_20574);
and U23713 (N_23713,N_21141,N_21992);
and U23714 (N_23714,N_21502,N_21880);
or U23715 (N_23715,N_22153,N_22308);
and U23716 (N_23716,N_21770,N_20656);
xnor U23717 (N_23717,N_20986,N_20555);
nor U23718 (N_23718,N_21801,N_22279);
and U23719 (N_23719,N_20041,N_22495);
nor U23720 (N_23720,N_20884,N_21787);
or U23721 (N_23721,N_21559,N_21736);
nor U23722 (N_23722,N_20821,N_21585);
or U23723 (N_23723,N_21707,N_20844);
nor U23724 (N_23724,N_20265,N_20145);
nand U23725 (N_23725,N_20144,N_20624);
nor U23726 (N_23726,N_20154,N_21959);
nor U23727 (N_23727,N_22292,N_22299);
nand U23728 (N_23728,N_21854,N_21062);
xor U23729 (N_23729,N_21021,N_21475);
xor U23730 (N_23730,N_20175,N_22206);
nor U23731 (N_23731,N_21427,N_20535);
nor U23732 (N_23732,N_20668,N_21799);
or U23733 (N_23733,N_20204,N_21353);
and U23734 (N_23734,N_22045,N_20178);
or U23735 (N_23735,N_20197,N_22097);
nand U23736 (N_23736,N_20003,N_21178);
or U23737 (N_23737,N_20661,N_22326);
and U23738 (N_23738,N_21181,N_22209);
nand U23739 (N_23739,N_21465,N_21771);
nand U23740 (N_23740,N_20728,N_22189);
nand U23741 (N_23741,N_20638,N_20073);
or U23742 (N_23742,N_22462,N_20234);
or U23743 (N_23743,N_21721,N_21978);
xnor U23744 (N_23744,N_21382,N_20578);
nor U23745 (N_23745,N_21352,N_21241);
nand U23746 (N_23746,N_22467,N_21960);
and U23747 (N_23747,N_21772,N_22491);
nor U23748 (N_23748,N_21406,N_20079);
or U23749 (N_23749,N_20595,N_22349);
and U23750 (N_23750,N_21937,N_21017);
and U23751 (N_23751,N_20677,N_20909);
and U23752 (N_23752,N_21921,N_20261);
or U23753 (N_23753,N_21411,N_20176);
xnor U23754 (N_23754,N_22057,N_21384);
or U23755 (N_23755,N_21470,N_21794);
or U23756 (N_23756,N_20544,N_20302);
nand U23757 (N_23757,N_22068,N_22315);
nor U23758 (N_23758,N_20867,N_21010);
nor U23759 (N_23759,N_20870,N_20492);
xnor U23760 (N_23760,N_21426,N_22396);
xnor U23761 (N_23761,N_21167,N_21174);
or U23762 (N_23762,N_20024,N_20984);
or U23763 (N_23763,N_21665,N_20147);
nor U23764 (N_23764,N_20825,N_20380);
nor U23765 (N_23765,N_21878,N_20791);
nand U23766 (N_23766,N_22163,N_21856);
nor U23767 (N_23767,N_21911,N_20329);
xor U23768 (N_23768,N_20313,N_20998);
or U23769 (N_23769,N_20660,N_20060);
nor U23770 (N_23770,N_20337,N_22065);
xor U23771 (N_23771,N_22376,N_21325);
nor U23772 (N_23772,N_20940,N_21806);
xor U23773 (N_23773,N_20522,N_20331);
nor U23774 (N_23774,N_20417,N_21065);
xor U23775 (N_23775,N_21077,N_21428);
nor U23776 (N_23776,N_21945,N_20979);
nand U23777 (N_23777,N_21534,N_20122);
xor U23778 (N_23778,N_21962,N_21036);
nor U23779 (N_23779,N_20959,N_20589);
nand U23780 (N_23780,N_21903,N_22010);
or U23781 (N_23781,N_20232,N_22137);
xor U23782 (N_23782,N_20732,N_21641);
xor U23783 (N_23783,N_20582,N_21648);
xnor U23784 (N_23784,N_20093,N_21092);
nand U23785 (N_23785,N_21293,N_21198);
nand U23786 (N_23786,N_21239,N_20548);
and U23787 (N_23787,N_22282,N_20035);
nand U23788 (N_23788,N_20896,N_22235);
and U23789 (N_23789,N_20028,N_21074);
nand U23790 (N_23790,N_22475,N_22102);
nand U23791 (N_23791,N_21451,N_20278);
or U23792 (N_23792,N_21192,N_20724);
xor U23793 (N_23793,N_21590,N_22467);
xnor U23794 (N_23794,N_21031,N_20580);
and U23795 (N_23795,N_21747,N_21443);
nor U23796 (N_23796,N_20849,N_21017);
and U23797 (N_23797,N_20821,N_21469);
or U23798 (N_23798,N_20312,N_21525);
and U23799 (N_23799,N_22340,N_20976);
and U23800 (N_23800,N_21159,N_21267);
or U23801 (N_23801,N_22353,N_20515);
and U23802 (N_23802,N_20918,N_22346);
or U23803 (N_23803,N_20947,N_21567);
xor U23804 (N_23804,N_20778,N_21323);
nand U23805 (N_23805,N_20161,N_20143);
nor U23806 (N_23806,N_20636,N_20012);
or U23807 (N_23807,N_21005,N_20453);
or U23808 (N_23808,N_22242,N_21393);
or U23809 (N_23809,N_22455,N_21074);
and U23810 (N_23810,N_21257,N_22383);
and U23811 (N_23811,N_22134,N_22005);
and U23812 (N_23812,N_20478,N_20114);
and U23813 (N_23813,N_20487,N_20429);
and U23814 (N_23814,N_21698,N_20381);
or U23815 (N_23815,N_21752,N_21468);
nor U23816 (N_23816,N_22063,N_20460);
and U23817 (N_23817,N_21825,N_20950);
or U23818 (N_23818,N_22384,N_22033);
and U23819 (N_23819,N_22033,N_21733);
and U23820 (N_23820,N_20732,N_20306);
and U23821 (N_23821,N_21086,N_22058);
and U23822 (N_23822,N_21380,N_21892);
and U23823 (N_23823,N_20618,N_21566);
and U23824 (N_23824,N_22088,N_20547);
nor U23825 (N_23825,N_20579,N_22481);
and U23826 (N_23826,N_20195,N_22339);
nor U23827 (N_23827,N_21836,N_20207);
nor U23828 (N_23828,N_22040,N_21209);
nand U23829 (N_23829,N_22105,N_21911);
xor U23830 (N_23830,N_21017,N_20963);
nand U23831 (N_23831,N_20265,N_21680);
or U23832 (N_23832,N_22358,N_22495);
and U23833 (N_23833,N_22415,N_21509);
xnor U23834 (N_23834,N_21617,N_20967);
xnor U23835 (N_23835,N_22446,N_21832);
nand U23836 (N_23836,N_20889,N_20302);
nor U23837 (N_23837,N_20214,N_21855);
nand U23838 (N_23838,N_21506,N_21615);
nand U23839 (N_23839,N_22483,N_21933);
nand U23840 (N_23840,N_21804,N_22462);
nor U23841 (N_23841,N_21467,N_21644);
xor U23842 (N_23842,N_20392,N_21253);
or U23843 (N_23843,N_22440,N_20242);
nand U23844 (N_23844,N_20409,N_20659);
nand U23845 (N_23845,N_20108,N_20104);
xnor U23846 (N_23846,N_21574,N_20512);
nand U23847 (N_23847,N_21925,N_21932);
nor U23848 (N_23848,N_22312,N_20180);
or U23849 (N_23849,N_20489,N_21584);
or U23850 (N_23850,N_21073,N_22291);
xor U23851 (N_23851,N_20687,N_21218);
and U23852 (N_23852,N_22264,N_22004);
nand U23853 (N_23853,N_21290,N_21306);
xor U23854 (N_23854,N_20190,N_21610);
or U23855 (N_23855,N_22016,N_20697);
xnor U23856 (N_23856,N_21727,N_21154);
nand U23857 (N_23857,N_20652,N_21204);
xor U23858 (N_23858,N_20713,N_20042);
xnor U23859 (N_23859,N_20011,N_21465);
nor U23860 (N_23860,N_21694,N_20261);
or U23861 (N_23861,N_20326,N_21515);
xnor U23862 (N_23862,N_20464,N_21686);
nand U23863 (N_23863,N_21366,N_21442);
nand U23864 (N_23864,N_20736,N_21718);
and U23865 (N_23865,N_21295,N_20355);
xor U23866 (N_23866,N_20159,N_22021);
nand U23867 (N_23867,N_21449,N_21813);
nand U23868 (N_23868,N_20108,N_20578);
and U23869 (N_23869,N_22447,N_20744);
and U23870 (N_23870,N_20810,N_20071);
nand U23871 (N_23871,N_22196,N_21671);
or U23872 (N_23872,N_20915,N_20996);
nor U23873 (N_23873,N_21296,N_21068);
nor U23874 (N_23874,N_20364,N_21923);
nand U23875 (N_23875,N_20705,N_20320);
xnor U23876 (N_23876,N_21544,N_21721);
xnor U23877 (N_23877,N_20273,N_20637);
nand U23878 (N_23878,N_22468,N_20238);
and U23879 (N_23879,N_20329,N_20295);
and U23880 (N_23880,N_20195,N_21409);
xor U23881 (N_23881,N_22414,N_20547);
nand U23882 (N_23882,N_20246,N_21202);
and U23883 (N_23883,N_21107,N_22416);
and U23884 (N_23884,N_21836,N_20947);
xor U23885 (N_23885,N_21177,N_22203);
xor U23886 (N_23886,N_21516,N_20077);
or U23887 (N_23887,N_21591,N_20064);
or U23888 (N_23888,N_20990,N_21633);
and U23889 (N_23889,N_21712,N_20024);
xor U23890 (N_23890,N_20589,N_20310);
or U23891 (N_23891,N_21186,N_20400);
nor U23892 (N_23892,N_21017,N_20948);
nor U23893 (N_23893,N_21190,N_21955);
nand U23894 (N_23894,N_22057,N_20440);
nand U23895 (N_23895,N_20178,N_20433);
nand U23896 (N_23896,N_20589,N_21247);
or U23897 (N_23897,N_20964,N_21112);
xor U23898 (N_23898,N_21547,N_20599);
or U23899 (N_23899,N_20518,N_21764);
or U23900 (N_23900,N_20318,N_20989);
and U23901 (N_23901,N_21669,N_20268);
or U23902 (N_23902,N_21549,N_22157);
or U23903 (N_23903,N_21548,N_22000);
xnor U23904 (N_23904,N_21958,N_21986);
nand U23905 (N_23905,N_21210,N_21521);
xnor U23906 (N_23906,N_20192,N_20630);
xor U23907 (N_23907,N_20923,N_22388);
nand U23908 (N_23908,N_22362,N_21349);
xnor U23909 (N_23909,N_20649,N_21299);
nor U23910 (N_23910,N_21076,N_20617);
xor U23911 (N_23911,N_22187,N_21722);
or U23912 (N_23912,N_20138,N_20933);
and U23913 (N_23913,N_21354,N_21266);
and U23914 (N_23914,N_20818,N_21770);
xnor U23915 (N_23915,N_20566,N_21596);
nor U23916 (N_23916,N_22388,N_20002);
and U23917 (N_23917,N_20010,N_22055);
xor U23918 (N_23918,N_20833,N_22486);
nor U23919 (N_23919,N_20738,N_21901);
or U23920 (N_23920,N_22038,N_21029);
or U23921 (N_23921,N_21755,N_20698);
xnor U23922 (N_23922,N_20960,N_21349);
xnor U23923 (N_23923,N_21587,N_20167);
nand U23924 (N_23924,N_21255,N_20519);
xnor U23925 (N_23925,N_21727,N_22349);
nor U23926 (N_23926,N_22412,N_21730);
xnor U23927 (N_23927,N_22348,N_20044);
or U23928 (N_23928,N_22274,N_21096);
and U23929 (N_23929,N_20624,N_20965);
or U23930 (N_23930,N_20615,N_20402);
and U23931 (N_23931,N_21264,N_21268);
nor U23932 (N_23932,N_22458,N_21094);
and U23933 (N_23933,N_21251,N_22184);
xnor U23934 (N_23934,N_20768,N_21335);
or U23935 (N_23935,N_20085,N_20683);
nor U23936 (N_23936,N_22242,N_20502);
nor U23937 (N_23937,N_22002,N_22129);
or U23938 (N_23938,N_20672,N_22337);
and U23939 (N_23939,N_21652,N_21107);
xor U23940 (N_23940,N_20361,N_22136);
or U23941 (N_23941,N_22248,N_20397);
nor U23942 (N_23942,N_22185,N_20319);
and U23943 (N_23943,N_21170,N_21166);
and U23944 (N_23944,N_20738,N_21784);
and U23945 (N_23945,N_21883,N_21279);
nor U23946 (N_23946,N_20827,N_21640);
xnor U23947 (N_23947,N_20470,N_22097);
xnor U23948 (N_23948,N_21460,N_21354);
or U23949 (N_23949,N_22226,N_21571);
nor U23950 (N_23950,N_20793,N_20920);
nor U23951 (N_23951,N_20354,N_22251);
and U23952 (N_23952,N_20022,N_22218);
nand U23953 (N_23953,N_22414,N_21832);
or U23954 (N_23954,N_20105,N_21347);
nor U23955 (N_23955,N_21043,N_20338);
nand U23956 (N_23956,N_20285,N_20186);
xor U23957 (N_23957,N_22235,N_21078);
and U23958 (N_23958,N_22212,N_21220);
nand U23959 (N_23959,N_22017,N_21927);
xnor U23960 (N_23960,N_20511,N_21780);
nand U23961 (N_23961,N_21700,N_21755);
nor U23962 (N_23962,N_21928,N_20246);
or U23963 (N_23963,N_20740,N_20594);
xor U23964 (N_23964,N_21866,N_20239);
nand U23965 (N_23965,N_21629,N_22064);
xor U23966 (N_23966,N_20934,N_20240);
and U23967 (N_23967,N_21420,N_20361);
nor U23968 (N_23968,N_21535,N_20908);
and U23969 (N_23969,N_20287,N_20358);
nand U23970 (N_23970,N_22070,N_21952);
or U23971 (N_23971,N_20550,N_20737);
and U23972 (N_23972,N_20294,N_20098);
or U23973 (N_23973,N_22160,N_20345);
and U23974 (N_23974,N_21294,N_21454);
xor U23975 (N_23975,N_21934,N_21811);
and U23976 (N_23976,N_21529,N_20839);
xnor U23977 (N_23977,N_21375,N_20434);
and U23978 (N_23978,N_20044,N_21255);
nand U23979 (N_23979,N_20557,N_21053);
and U23980 (N_23980,N_21024,N_21133);
or U23981 (N_23981,N_21542,N_21085);
or U23982 (N_23982,N_21696,N_21058);
or U23983 (N_23983,N_20486,N_21305);
nand U23984 (N_23984,N_22149,N_20802);
xor U23985 (N_23985,N_21113,N_21543);
or U23986 (N_23986,N_20548,N_20131);
xor U23987 (N_23987,N_20922,N_21192);
nor U23988 (N_23988,N_21972,N_21601);
and U23989 (N_23989,N_20943,N_21103);
xnor U23990 (N_23990,N_21980,N_22377);
nand U23991 (N_23991,N_22072,N_20139);
or U23992 (N_23992,N_21094,N_20863);
and U23993 (N_23993,N_20391,N_20154);
nor U23994 (N_23994,N_20715,N_20891);
or U23995 (N_23995,N_21637,N_20234);
or U23996 (N_23996,N_21083,N_20765);
xor U23997 (N_23997,N_22260,N_21418);
xnor U23998 (N_23998,N_20305,N_21131);
or U23999 (N_23999,N_22249,N_22230);
nand U24000 (N_24000,N_22396,N_20934);
or U24001 (N_24001,N_21587,N_22065);
nand U24002 (N_24002,N_21913,N_22405);
xor U24003 (N_24003,N_21057,N_20137);
nor U24004 (N_24004,N_20605,N_20537);
xor U24005 (N_24005,N_21225,N_21436);
xor U24006 (N_24006,N_20395,N_21102);
and U24007 (N_24007,N_22368,N_20971);
or U24008 (N_24008,N_21241,N_21648);
and U24009 (N_24009,N_20589,N_20588);
or U24010 (N_24010,N_20243,N_22469);
nand U24011 (N_24011,N_20211,N_21859);
xnor U24012 (N_24012,N_21981,N_22255);
or U24013 (N_24013,N_20282,N_20320);
nand U24014 (N_24014,N_20171,N_21462);
xor U24015 (N_24015,N_21606,N_21865);
nand U24016 (N_24016,N_20246,N_21018);
nand U24017 (N_24017,N_20987,N_22191);
nor U24018 (N_24018,N_21673,N_20516);
xor U24019 (N_24019,N_20199,N_21120);
nand U24020 (N_24020,N_20376,N_21098);
nor U24021 (N_24021,N_22087,N_22426);
nand U24022 (N_24022,N_20827,N_20731);
and U24023 (N_24023,N_21711,N_20687);
nor U24024 (N_24024,N_21913,N_22021);
nor U24025 (N_24025,N_21881,N_20829);
xnor U24026 (N_24026,N_21658,N_20009);
or U24027 (N_24027,N_20486,N_20676);
xnor U24028 (N_24028,N_21513,N_21674);
nand U24029 (N_24029,N_21105,N_21922);
nand U24030 (N_24030,N_20572,N_22472);
nand U24031 (N_24031,N_22379,N_20729);
nand U24032 (N_24032,N_21664,N_21793);
nor U24033 (N_24033,N_22187,N_22345);
nor U24034 (N_24034,N_20454,N_20036);
and U24035 (N_24035,N_21088,N_21312);
nand U24036 (N_24036,N_21904,N_21340);
and U24037 (N_24037,N_20909,N_20810);
nor U24038 (N_24038,N_20716,N_22278);
or U24039 (N_24039,N_21328,N_22047);
xnor U24040 (N_24040,N_20254,N_22044);
nand U24041 (N_24041,N_20036,N_21098);
and U24042 (N_24042,N_20265,N_20688);
xnor U24043 (N_24043,N_20015,N_20768);
or U24044 (N_24044,N_20494,N_22308);
xnor U24045 (N_24045,N_20666,N_20037);
nor U24046 (N_24046,N_20816,N_21934);
xor U24047 (N_24047,N_20657,N_20756);
and U24048 (N_24048,N_20470,N_21373);
nor U24049 (N_24049,N_21013,N_21956);
nor U24050 (N_24050,N_20163,N_20450);
xor U24051 (N_24051,N_20409,N_22069);
nor U24052 (N_24052,N_20300,N_21290);
or U24053 (N_24053,N_20607,N_22256);
and U24054 (N_24054,N_22346,N_20670);
nor U24055 (N_24055,N_20212,N_22209);
nor U24056 (N_24056,N_20907,N_22314);
nor U24057 (N_24057,N_20883,N_22237);
nor U24058 (N_24058,N_22279,N_21373);
or U24059 (N_24059,N_20619,N_21828);
or U24060 (N_24060,N_20802,N_20334);
nor U24061 (N_24061,N_20648,N_22464);
nor U24062 (N_24062,N_21250,N_20785);
and U24063 (N_24063,N_20455,N_20127);
nand U24064 (N_24064,N_20699,N_21385);
xnor U24065 (N_24065,N_20743,N_20574);
or U24066 (N_24066,N_20103,N_21990);
nor U24067 (N_24067,N_21052,N_22238);
xnor U24068 (N_24068,N_21373,N_20499);
nand U24069 (N_24069,N_21577,N_21532);
nor U24070 (N_24070,N_20801,N_20516);
and U24071 (N_24071,N_21508,N_22135);
and U24072 (N_24072,N_21079,N_20717);
or U24073 (N_24073,N_20353,N_21673);
and U24074 (N_24074,N_20517,N_20884);
xnor U24075 (N_24075,N_21135,N_22011);
and U24076 (N_24076,N_22219,N_20978);
xnor U24077 (N_24077,N_22477,N_21377);
and U24078 (N_24078,N_21911,N_21444);
nand U24079 (N_24079,N_20318,N_21492);
xor U24080 (N_24080,N_22279,N_21032);
and U24081 (N_24081,N_22186,N_21149);
xor U24082 (N_24082,N_20226,N_20252);
nand U24083 (N_24083,N_21612,N_21519);
and U24084 (N_24084,N_20165,N_21550);
nor U24085 (N_24085,N_20817,N_20938);
xnor U24086 (N_24086,N_22061,N_20450);
and U24087 (N_24087,N_22348,N_20360);
and U24088 (N_24088,N_21753,N_20516);
xor U24089 (N_24089,N_20740,N_21943);
or U24090 (N_24090,N_20022,N_22048);
xor U24091 (N_24091,N_20911,N_20834);
or U24092 (N_24092,N_20949,N_20559);
nor U24093 (N_24093,N_20189,N_20354);
xnor U24094 (N_24094,N_20322,N_21608);
or U24095 (N_24095,N_22128,N_21020);
nand U24096 (N_24096,N_20820,N_21726);
xnor U24097 (N_24097,N_20856,N_22026);
and U24098 (N_24098,N_22034,N_21691);
or U24099 (N_24099,N_21586,N_21061);
xnor U24100 (N_24100,N_22443,N_20478);
xnor U24101 (N_24101,N_21690,N_21426);
and U24102 (N_24102,N_22028,N_20539);
or U24103 (N_24103,N_20000,N_22088);
or U24104 (N_24104,N_21226,N_20225);
or U24105 (N_24105,N_22432,N_22079);
nor U24106 (N_24106,N_21759,N_20725);
nand U24107 (N_24107,N_21464,N_21210);
nand U24108 (N_24108,N_21936,N_20781);
and U24109 (N_24109,N_20629,N_21765);
and U24110 (N_24110,N_22030,N_21083);
xor U24111 (N_24111,N_20814,N_20811);
nor U24112 (N_24112,N_22273,N_21609);
or U24113 (N_24113,N_21191,N_20161);
or U24114 (N_24114,N_20084,N_21067);
or U24115 (N_24115,N_21688,N_20471);
nor U24116 (N_24116,N_20605,N_22434);
or U24117 (N_24117,N_21096,N_21219);
or U24118 (N_24118,N_22306,N_21307);
xor U24119 (N_24119,N_21322,N_21390);
nand U24120 (N_24120,N_20995,N_20777);
and U24121 (N_24121,N_20524,N_21307);
nand U24122 (N_24122,N_21028,N_21986);
or U24123 (N_24123,N_20179,N_21011);
and U24124 (N_24124,N_22327,N_21295);
or U24125 (N_24125,N_21843,N_21589);
or U24126 (N_24126,N_20473,N_20820);
nand U24127 (N_24127,N_22452,N_21881);
xor U24128 (N_24128,N_21509,N_21461);
and U24129 (N_24129,N_21876,N_21961);
nand U24130 (N_24130,N_22443,N_21410);
and U24131 (N_24131,N_21658,N_21684);
nand U24132 (N_24132,N_22461,N_20270);
and U24133 (N_24133,N_20536,N_22037);
and U24134 (N_24134,N_20994,N_20595);
or U24135 (N_24135,N_21028,N_21692);
xnor U24136 (N_24136,N_22298,N_20026);
xor U24137 (N_24137,N_22215,N_21569);
and U24138 (N_24138,N_20873,N_22324);
and U24139 (N_24139,N_22230,N_22391);
nor U24140 (N_24140,N_20922,N_21066);
nand U24141 (N_24141,N_22448,N_20030);
or U24142 (N_24142,N_21663,N_20319);
nand U24143 (N_24143,N_21602,N_21207);
nor U24144 (N_24144,N_20568,N_21947);
nor U24145 (N_24145,N_20161,N_21013);
and U24146 (N_24146,N_20598,N_21572);
and U24147 (N_24147,N_21286,N_20212);
nor U24148 (N_24148,N_20260,N_20674);
nand U24149 (N_24149,N_20363,N_21373);
nor U24150 (N_24150,N_21744,N_20780);
or U24151 (N_24151,N_20497,N_21532);
or U24152 (N_24152,N_20580,N_21099);
and U24153 (N_24153,N_20852,N_21996);
xor U24154 (N_24154,N_21042,N_21735);
nor U24155 (N_24155,N_21474,N_21107);
and U24156 (N_24156,N_20832,N_20151);
xor U24157 (N_24157,N_20447,N_21559);
xor U24158 (N_24158,N_21011,N_20565);
xor U24159 (N_24159,N_21983,N_21848);
and U24160 (N_24160,N_20333,N_21115);
nor U24161 (N_24161,N_21508,N_21173);
xnor U24162 (N_24162,N_20488,N_20708);
or U24163 (N_24163,N_21156,N_21251);
nor U24164 (N_24164,N_20038,N_21195);
and U24165 (N_24165,N_22392,N_22025);
or U24166 (N_24166,N_20893,N_22375);
nor U24167 (N_24167,N_20142,N_20619);
or U24168 (N_24168,N_21177,N_21491);
nor U24169 (N_24169,N_22208,N_22005);
nand U24170 (N_24170,N_20298,N_22332);
nor U24171 (N_24171,N_20715,N_20342);
and U24172 (N_24172,N_20605,N_20016);
xor U24173 (N_24173,N_22003,N_21187);
nor U24174 (N_24174,N_20567,N_20440);
xnor U24175 (N_24175,N_21298,N_20155);
nand U24176 (N_24176,N_20912,N_21363);
xnor U24177 (N_24177,N_20343,N_22133);
or U24178 (N_24178,N_20396,N_22230);
nor U24179 (N_24179,N_22151,N_21780);
nand U24180 (N_24180,N_21292,N_22396);
nand U24181 (N_24181,N_20981,N_20230);
xnor U24182 (N_24182,N_20822,N_20689);
nor U24183 (N_24183,N_20972,N_22202);
xor U24184 (N_24184,N_21699,N_20250);
nor U24185 (N_24185,N_22463,N_20100);
xnor U24186 (N_24186,N_21729,N_20386);
nand U24187 (N_24187,N_21325,N_21431);
and U24188 (N_24188,N_22253,N_21880);
and U24189 (N_24189,N_21213,N_21741);
or U24190 (N_24190,N_20414,N_21325);
xor U24191 (N_24191,N_21236,N_21239);
xor U24192 (N_24192,N_21242,N_22144);
xor U24193 (N_24193,N_22023,N_21159);
nand U24194 (N_24194,N_21559,N_22356);
and U24195 (N_24195,N_20438,N_20471);
nand U24196 (N_24196,N_21860,N_20905);
nand U24197 (N_24197,N_21542,N_20006);
nand U24198 (N_24198,N_20167,N_21672);
or U24199 (N_24199,N_21636,N_22287);
nor U24200 (N_24200,N_20048,N_20741);
or U24201 (N_24201,N_22438,N_21942);
or U24202 (N_24202,N_22282,N_20808);
nand U24203 (N_24203,N_20454,N_20619);
xor U24204 (N_24204,N_20205,N_20642);
nor U24205 (N_24205,N_20728,N_20625);
nor U24206 (N_24206,N_21807,N_21988);
nand U24207 (N_24207,N_22373,N_22070);
or U24208 (N_24208,N_20208,N_20129);
xor U24209 (N_24209,N_21058,N_22366);
nor U24210 (N_24210,N_20983,N_20977);
and U24211 (N_24211,N_20609,N_21833);
nand U24212 (N_24212,N_20448,N_21861);
nor U24213 (N_24213,N_22082,N_22210);
xnor U24214 (N_24214,N_20525,N_22007);
nand U24215 (N_24215,N_22096,N_22031);
and U24216 (N_24216,N_21040,N_22420);
nor U24217 (N_24217,N_20419,N_22212);
and U24218 (N_24218,N_21011,N_20666);
nor U24219 (N_24219,N_22240,N_20066);
xor U24220 (N_24220,N_21308,N_20233);
nand U24221 (N_24221,N_21093,N_21018);
xor U24222 (N_24222,N_21512,N_20489);
nor U24223 (N_24223,N_21216,N_21586);
and U24224 (N_24224,N_20947,N_21868);
and U24225 (N_24225,N_21093,N_20031);
or U24226 (N_24226,N_21652,N_22209);
and U24227 (N_24227,N_22028,N_20327);
xnor U24228 (N_24228,N_20475,N_20712);
and U24229 (N_24229,N_21410,N_20085);
nor U24230 (N_24230,N_20511,N_20074);
nor U24231 (N_24231,N_22244,N_21013);
nor U24232 (N_24232,N_20103,N_21958);
and U24233 (N_24233,N_20041,N_21094);
xnor U24234 (N_24234,N_20788,N_20599);
nand U24235 (N_24235,N_20677,N_21096);
or U24236 (N_24236,N_20425,N_21219);
or U24237 (N_24237,N_20508,N_20721);
nor U24238 (N_24238,N_21742,N_20846);
nand U24239 (N_24239,N_20294,N_21594);
and U24240 (N_24240,N_21207,N_21693);
xor U24241 (N_24241,N_22475,N_20839);
nand U24242 (N_24242,N_21342,N_21878);
nor U24243 (N_24243,N_20875,N_21943);
nand U24244 (N_24244,N_21734,N_20223);
nor U24245 (N_24245,N_21929,N_20732);
and U24246 (N_24246,N_22032,N_20221);
nand U24247 (N_24247,N_22066,N_21815);
nand U24248 (N_24248,N_21876,N_20204);
and U24249 (N_24249,N_20971,N_20217);
xnor U24250 (N_24250,N_20126,N_20812);
and U24251 (N_24251,N_21357,N_21925);
xor U24252 (N_24252,N_22233,N_22294);
or U24253 (N_24253,N_21282,N_20775);
and U24254 (N_24254,N_20157,N_21121);
or U24255 (N_24255,N_22170,N_21833);
nand U24256 (N_24256,N_21092,N_21756);
nor U24257 (N_24257,N_21786,N_20083);
xor U24258 (N_24258,N_20640,N_22073);
and U24259 (N_24259,N_21882,N_20943);
nand U24260 (N_24260,N_21851,N_20869);
nand U24261 (N_24261,N_22248,N_20882);
and U24262 (N_24262,N_21305,N_22225);
xor U24263 (N_24263,N_20680,N_21899);
nor U24264 (N_24264,N_22171,N_22046);
xnor U24265 (N_24265,N_21867,N_22159);
or U24266 (N_24266,N_20400,N_21693);
xor U24267 (N_24267,N_20791,N_21783);
nand U24268 (N_24268,N_21047,N_22415);
and U24269 (N_24269,N_21794,N_20134);
nand U24270 (N_24270,N_21162,N_21110);
xor U24271 (N_24271,N_20097,N_22061);
xnor U24272 (N_24272,N_20904,N_21674);
xnor U24273 (N_24273,N_21746,N_22304);
and U24274 (N_24274,N_21464,N_22437);
and U24275 (N_24275,N_20599,N_20372);
nand U24276 (N_24276,N_20093,N_22419);
nand U24277 (N_24277,N_20149,N_21667);
or U24278 (N_24278,N_20086,N_21644);
xor U24279 (N_24279,N_21951,N_22065);
nand U24280 (N_24280,N_21494,N_20522);
or U24281 (N_24281,N_21196,N_21979);
or U24282 (N_24282,N_21678,N_20827);
xor U24283 (N_24283,N_22027,N_20687);
xor U24284 (N_24284,N_21103,N_21068);
and U24285 (N_24285,N_22381,N_20336);
or U24286 (N_24286,N_20267,N_21285);
nor U24287 (N_24287,N_20632,N_21971);
and U24288 (N_24288,N_20866,N_20187);
nor U24289 (N_24289,N_20883,N_22012);
or U24290 (N_24290,N_22018,N_21011);
xnor U24291 (N_24291,N_21728,N_20661);
and U24292 (N_24292,N_20597,N_20059);
nor U24293 (N_24293,N_21586,N_21060);
nand U24294 (N_24294,N_21157,N_20354);
nand U24295 (N_24295,N_21679,N_22351);
nor U24296 (N_24296,N_20186,N_21100);
nor U24297 (N_24297,N_21516,N_21111);
and U24298 (N_24298,N_21112,N_22259);
nand U24299 (N_24299,N_21948,N_20061);
or U24300 (N_24300,N_22373,N_21106);
nor U24301 (N_24301,N_21297,N_21050);
nor U24302 (N_24302,N_20907,N_21857);
nor U24303 (N_24303,N_21527,N_20302);
xor U24304 (N_24304,N_21107,N_20405);
nand U24305 (N_24305,N_20732,N_21632);
nor U24306 (N_24306,N_20955,N_21756);
xor U24307 (N_24307,N_20464,N_20515);
nor U24308 (N_24308,N_22173,N_22114);
or U24309 (N_24309,N_22487,N_22417);
and U24310 (N_24310,N_21985,N_22063);
or U24311 (N_24311,N_20223,N_20983);
nor U24312 (N_24312,N_20951,N_21831);
xnor U24313 (N_24313,N_21770,N_21692);
xor U24314 (N_24314,N_22407,N_21306);
and U24315 (N_24315,N_20662,N_22473);
or U24316 (N_24316,N_20402,N_21309);
xnor U24317 (N_24317,N_21586,N_21280);
or U24318 (N_24318,N_21612,N_21981);
or U24319 (N_24319,N_21737,N_20094);
nor U24320 (N_24320,N_22219,N_22235);
xnor U24321 (N_24321,N_20234,N_20238);
nand U24322 (N_24322,N_22113,N_21978);
or U24323 (N_24323,N_21939,N_20636);
nor U24324 (N_24324,N_22470,N_21605);
and U24325 (N_24325,N_20132,N_21863);
xnor U24326 (N_24326,N_21369,N_21080);
or U24327 (N_24327,N_20133,N_21255);
nand U24328 (N_24328,N_21336,N_20047);
and U24329 (N_24329,N_21329,N_22121);
nand U24330 (N_24330,N_20206,N_22425);
nand U24331 (N_24331,N_20724,N_20940);
xor U24332 (N_24332,N_21526,N_21325);
nand U24333 (N_24333,N_20883,N_21302);
nor U24334 (N_24334,N_22354,N_21071);
nor U24335 (N_24335,N_20570,N_21804);
nor U24336 (N_24336,N_20939,N_22394);
nand U24337 (N_24337,N_20518,N_22418);
and U24338 (N_24338,N_22123,N_20831);
or U24339 (N_24339,N_22122,N_22220);
nand U24340 (N_24340,N_22146,N_22481);
nor U24341 (N_24341,N_20477,N_20688);
and U24342 (N_24342,N_20030,N_20515);
and U24343 (N_24343,N_21700,N_20946);
xnor U24344 (N_24344,N_20051,N_20551);
or U24345 (N_24345,N_21080,N_20557);
or U24346 (N_24346,N_21425,N_20708);
or U24347 (N_24347,N_21300,N_21536);
xor U24348 (N_24348,N_20708,N_21888);
xor U24349 (N_24349,N_21305,N_22404);
nor U24350 (N_24350,N_20043,N_20037);
xor U24351 (N_24351,N_20267,N_20880);
or U24352 (N_24352,N_20042,N_21302);
nand U24353 (N_24353,N_21966,N_20809);
or U24354 (N_24354,N_21759,N_21720);
or U24355 (N_24355,N_21489,N_21792);
xnor U24356 (N_24356,N_21265,N_21356);
xor U24357 (N_24357,N_21329,N_21429);
xor U24358 (N_24358,N_22321,N_20888);
or U24359 (N_24359,N_20832,N_21606);
and U24360 (N_24360,N_20802,N_21396);
nand U24361 (N_24361,N_21191,N_21617);
and U24362 (N_24362,N_21874,N_21408);
xor U24363 (N_24363,N_22496,N_22370);
or U24364 (N_24364,N_21816,N_20107);
xnor U24365 (N_24365,N_20637,N_21133);
nor U24366 (N_24366,N_22457,N_20269);
or U24367 (N_24367,N_21792,N_21376);
nand U24368 (N_24368,N_21356,N_20539);
nor U24369 (N_24369,N_21356,N_22091);
xor U24370 (N_24370,N_21881,N_21286);
and U24371 (N_24371,N_21664,N_21536);
xor U24372 (N_24372,N_21260,N_21304);
or U24373 (N_24373,N_21110,N_21641);
or U24374 (N_24374,N_22083,N_21125);
xnor U24375 (N_24375,N_22359,N_22406);
xnor U24376 (N_24376,N_22221,N_20958);
xor U24377 (N_24377,N_20357,N_20120);
or U24378 (N_24378,N_20301,N_20590);
xnor U24379 (N_24379,N_20115,N_20747);
xor U24380 (N_24380,N_21161,N_20705);
xnor U24381 (N_24381,N_21159,N_22085);
or U24382 (N_24382,N_21674,N_21924);
nand U24383 (N_24383,N_21613,N_20527);
or U24384 (N_24384,N_20678,N_20988);
nor U24385 (N_24385,N_21424,N_20950);
xor U24386 (N_24386,N_21024,N_21890);
and U24387 (N_24387,N_20855,N_20465);
or U24388 (N_24388,N_22334,N_21780);
xnor U24389 (N_24389,N_20485,N_20647);
or U24390 (N_24390,N_21963,N_20575);
xor U24391 (N_24391,N_22019,N_20052);
xnor U24392 (N_24392,N_20457,N_20636);
nor U24393 (N_24393,N_21475,N_20127);
nor U24394 (N_24394,N_20444,N_22063);
or U24395 (N_24395,N_21111,N_20143);
xnor U24396 (N_24396,N_22226,N_21348);
xor U24397 (N_24397,N_20163,N_20027);
nor U24398 (N_24398,N_21414,N_21715);
nand U24399 (N_24399,N_21690,N_21661);
nand U24400 (N_24400,N_20484,N_21288);
xor U24401 (N_24401,N_20264,N_20668);
or U24402 (N_24402,N_21581,N_22124);
nand U24403 (N_24403,N_20634,N_21386);
nor U24404 (N_24404,N_20629,N_21435);
and U24405 (N_24405,N_20309,N_20971);
xor U24406 (N_24406,N_20446,N_20969);
nand U24407 (N_24407,N_21568,N_22055);
xor U24408 (N_24408,N_21661,N_20043);
or U24409 (N_24409,N_21760,N_21657);
or U24410 (N_24410,N_21061,N_21312);
nand U24411 (N_24411,N_20528,N_20086);
or U24412 (N_24412,N_20355,N_20122);
or U24413 (N_24413,N_22382,N_20484);
or U24414 (N_24414,N_20224,N_20904);
nand U24415 (N_24415,N_20274,N_20315);
nand U24416 (N_24416,N_21408,N_22287);
xor U24417 (N_24417,N_21891,N_21309);
or U24418 (N_24418,N_22216,N_21689);
and U24419 (N_24419,N_20314,N_21542);
xnor U24420 (N_24420,N_20007,N_20352);
and U24421 (N_24421,N_21401,N_21531);
nor U24422 (N_24422,N_20054,N_22359);
xnor U24423 (N_24423,N_21207,N_21491);
or U24424 (N_24424,N_21716,N_20964);
nor U24425 (N_24425,N_20440,N_21184);
or U24426 (N_24426,N_21664,N_20692);
or U24427 (N_24427,N_21220,N_21369);
nor U24428 (N_24428,N_21082,N_22082);
nand U24429 (N_24429,N_20706,N_21821);
nand U24430 (N_24430,N_21911,N_21739);
nor U24431 (N_24431,N_21791,N_21042);
nand U24432 (N_24432,N_20998,N_20948);
or U24433 (N_24433,N_20428,N_20462);
xnor U24434 (N_24434,N_21989,N_22047);
nor U24435 (N_24435,N_20279,N_22026);
nor U24436 (N_24436,N_20843,N_21729);
nor U24437 (N_24437,N_21369,N_21754);
nor U24438 (N_24438,N_20408,N_22110);
xor U24439 (N_24439,N_20388,N_21886);
or U24440 (N_24440,N_21246,N_21149);
or U24441 (N_24441,N_21096,N_22417);
nand U24442 (N_24442,N_20210,N_20945);
xnor U24443 (N_24443,N_22448,N_21338);
nand U24444 (N_24444,N_20315,N_20922);
and U24445 (N_24445,N_22270,N_21797);
or U24446 (N_24446,N_22129,N_20655);
nand U24447 (N_24447,N_22425,N_22382);
or U24448 (N_24448,N_21892,N_20213);
nand U24449 (N_24449,N_21785,N_20598);
xnor U24450 (N_24450,N_21080,N_22420);
and U24451 (N_24451,N_20272,N_20723);
and U24452 (N_24452,N_20661,N_21783);
and U24453 (N_24453,N_21704,N_22492);
nor U24454 (N_24454,N_21977,N_21539);
nand U24455 (N_24455,N_21003,N_22485);
xnor U24456 (N_24456,N_21930,N_22316);
nor U24457 (N_24457,N_21373,N_21912);
nor U24458 (N_24458,N_22425,N_21237);
xnor U24459 (N_24459,N_22337,N_20982);
nand U24460 (N_24460,N_21094,N_21700);
xnor U24461 (N_24461,N_21579,N_21169);
nor U24462 (N_24462,N_21809,N_20370);
and U24463 (N_24463,N_20824,N_21826);
nor U24464 (N_24464,N_22490,N_21221);
nor U24465 (N_24465,N_21034,N_21680);
nand U24466 (N_24466,N_22307,N_21677);
nand U24467 (N_24467,N_21903,N_20098);
and U24468 (N_24468,N_20734,N_22160);
or U24469 (N_24469,N_21434,N_20772);
nor U24470 (N_24470,N_22386,N_20073);
nand U24471 (N_24471,N_21105,N_20608);
nand U24472 (N_24472,N_20726,N_20481);
nor U24473 (N_24473,N_20660,N_22267);
nand U24474 (N_24474,N_20780,N_22093);
xor U24475 (N_24475,N_20352,N_21149);
nand U24476 (N_24476,N_20345,N_21795);
nand U24477 (N_24477,N_21199,N_21326);
and U24478 (N_24478,N_21486,N_21534);
or U24479 (N_24479,N_21067,N_20059);
xor U24480 (N_24480,N_22263,N_20634);
nor U24481 (N_24481,N_20604,N_20028);
xor U24482 (N_24482,N_21861,N_21379);
nor U24483 (N_24483,N_21115,N_21673);
xor U24484 (N_24484,N_20241,N_22430);
or U24485 (N_24485,N_22297,N_21833);
or U24486 (N_24486,N_21958,N_20714);
and U24487 (N_24487,N_20123,N_20945);
nand U24488 (N_24488,N_20443,N_22005);
nor U24489 (N_24489,N_22460,N_22499);
or U24490 (N_24490,N_22177,N_21574);
nand U24491 (N_24491,N_20597,N_20105);
nand U24492 (N_24492,N_21207,N_20482);
nor U24493 (N_24493,N_21402,N_20751);
nand U24494 (N_24494,N_22407,N_21419);
or U24495 (N_24495,N_21833,N_21102);
and U24496 (N_24496,N_20864,N_20943);
nor U24497 (N_24497,N_22189,N_21924);
xor U24498 (N_24498,N_22386,N_20079);
nor U24499 (N_24499,N_20660,N_20636);
xor U24500 (N_24500,N_21630,N_20403);
nand U24501 (N_24501,N_20294,N_21393);
or U24502 (N_24502,N_20183,N_22299);
and U24503 (N_24503,N_22058,N_20292);
and U24504 (N_24504,N_20659,N_21551);
and U24505 (N_24505,N_21360,N_22002);
nor U24506 (N_24506,N_22329,N_21359);
xor U24507 (N_24507,N_20010,N_21027);
and U24508 (N_24508,N_21267,N_20363);
xnor U24509 (N_24509,N_20737,N_20870);
and U24510 (N_24510,N_20486,N_20012);
nor U24511 (N_24511,N_21408,N_20124);
nor U24512 (N_24512,N_21506,N_20751);
nor U24513 (N_24513,N_21174,N_22133);
or U24514 (N_24514,N_21999,N_21409);
nor U24515 (N_24515,N_20215,N_22318);
xnor U24516 (N_24516,N_21433,N_21959);
or U24517 (N_24517,N_20016,N_20418);
xnor U24518 (N_24518,N_21770,N_20021);
xor U24519 (N_24519,N_22306,N_20199);
nor U24520 (N_24520,N_21011,N_22437);
and U24521 (N_24521,N_20200,N_21188);
nor U24522 (N_24522,N_21880,N_21735);
xor U24523 (N_24523,N_21959,N_20478);
nand U24524 (N_24524,N_22086,N_22068);
xor U24525 (N_24525,N_22481,N_22093);
and U24526 (N_24526,N_21990,N_21096);
or U24527 (N_24527,N_20734,N_22494);
nand U24528 (N_24528,N_20506,N_20163);
nor U24529 (N_24529,N_21715,N_21981);
and U24530 (N_24530,N_20760,N_20018);
xor U24531 (N_24531,N_21880,N_20071);
and U24532 (N_24532,N_20598,N_20050);
or U24533 (N_24533,N_22492,N_21287);
nor U24534 (N_24534,N_20454,N_20087);
or U24535 (N_24535,N_21665,N_21522);
nand U24536 (N_24536,N_20364,N_20927);
nand U24537 (N_24537,N_20236,N_22332);
xnor U24538 (N_24538,N_20182,N_20626);
xnor U24539 (N_24539,N_21124,N_20147);
and U24540 (N_24540,N_21878,N_21297);
nand U24541 (N_24541,N_21574,N_22041);
nand U24542 (N_24542,N_22013,N_21016);
nand U24543 (N_24543,N_22434,N_21575);
xor U24544 (N_24544,N_21203,N_21701);
nand U24545 (N_24545,N_20537,N_21770);
nand U24546 (N_24546,N_20112,N_22457);
xor U24547 (N_24547,N_21164,N_20746);
and U24548 (N_24548,N_20904,N_20827);
xnor U24549 (N_24549,N_20836,N_21637);
nor U24550 (N_24550,N_20124,N_20131);
and U24551 (N_24551,N_20667,N_21859);
xor U24552 (N_24552,N_22274,N_22445);
xnor U24553 (N_24553,N_21533,N_20334);
xnor U24554 (N_24554,N_20627,N_20427);
xor U24555 (N_24555,N_21492,N_21419);
xnor U24556 (N_24556,N_21984,N_21463);
nand U24557 (N_24557,N_20709,N_20547);
nor U24558 (N_24558,N_22336,N_22008);
nand U24559 (N_24559,N_21054,N_20827);
nand U24560 (N_24560,N_20482,N_21569);
xor U24561 (N_24561,N_21030,N_20668);
xor U24562 (N_24562,N_20443,N_21564);
and U24563 (N_24563,N_22307,N_21351);
xnor U24564 (N_24564,N_22176,N_20802);
nand U24565 (N_24565,N_22363,N_21348);
nor U24566 (N_24566,N_20420,N_20418);
nor U24567 (N_24567,N_21528,N_20301);
nor U24568 (N_24568,N_22312,N_21681);
nor U24569 (N_24569,N_21330,N_22324);
and U24570 (N_24570,N_20512,N_21098);
or U24571 (N_24571,N_21579,N_21087);
xnor U24572 (N_24572,N_21207,N_20672);
nor U24573 (N_24573,N_20072,N_21952);
nand U24574 (N_24574,N_20870,N_20780);
nor U24575 (N_24575,N_21559,N_22247);
nand U24576 (N_24576,N_20446,N_20063);
and U24577 (N_24577,N_20541,N_20269);
nor U24578 (N_24578,N_21758,N_21693);
nor U24579 (N_24579,N_22042,N_20425);
and U24580 (N_24580,N_22465,N_20280);
or U24581 (N_24581,N_21001,N_20578);
or U24582 (N_24582,N_20181,N_21113);
nand U24583 (N_24583,N_20715,N_21766);
and U24584 (N_24584,N_20591,N_20714);
xnor U24585 (N_24585,N_22470,N_22061);
xnor U24586 (N_24586,N_20558,N_21064);
nor U24587 (N_24587,N_22322,N_20220);
or U24588 (N_24588,N_22475,N_20030);
nand U24589 (N_24589,N_22277,N_21521);
nor U24590 (N_24590,N_21726,N_21703);
or U24591 (N_24591,N_20418,N_20298);
or U24592 (N_24592,N_20685,N_22129);
nor U24593 (N_24593,N_20711,N_21632);
nor U24594 (N_24594,N_22232,N_20129);
or U24595 (N_24595,N_21982,N_21439);
nor U24596 (N_24596,N_20877,N_22446);
and U24597 (N_24597,N_22367,N_21529);
nand U24598 (N_24598,N_22051,N_21363);
nand U24599 (N_24599,N_22411,N_20058);
xor U24600 (N_24600,N_20775,N_20680);
nand U24601 (N_24601,N_22245,N_22428);
xnor U24602 (N_24602,N_22056,N_22255);
nand U24603 (N_24603,N_21327,N_20987);
xnor U24604 (N_24604,N_21821,N_20156);
nand U24605 (N_24605,N_22153,N_22067);
xnor U24606 (N_24606,N_20349,N_22182);
nor U24607 (N_24607,N_20162,N_21044);
xor U24608 (N_24608,N_21742,N_21567);
or U24609 (N_24609,N_21501,N_20718);
xnor U24610 (N_24610,N_22328,N_20934);
and U24611 (N_24611,N_21865,N_22004);
nand U24612 (N_24612,N_21872,N_20058);
xnor U24613 (N_24613,N_22388,N_20694);
nand U24614 (N_24614,N_20552,N_22328);
nand U24615 (N_24615,N_20576,N_21279);
xor U24616 (N_24616,N_22328,N_21500);
nor U24617 (N_24617,N_22051,N_22046);
nand U24618 (N_24618,N_21405,N_20756);
or U24619 (N_24619,N_21776,N_20129);
xor U24620 (N_24620,N_22292,N_21330);
and U24621 (N_24621,N_20212,N_20715);
or U24622 (N_24622,N_20414,N_21399);
nor U24623 (N_24623,N_21659,N_22465);
nand U24624 (N_24624,N_22000,N_21307);
or U24625 (N_24625,N_20712,N_20072);
or U24626 (N_24626,N_21076,N_21719);
nand U24627 (N_24627,N_20473,N_20247);
or U24628 (N_24628,N_22212,N_21866);
and U24629 (N_24629,N_20441,N_22013);
nand U24630 (N_24630,N_20657,N_20024);
and U24631 (N_24631,N_21013,N_20868);
or U24632 (N_24632,N_20115,N_22312);
nand U24633 (N_24633,N_21416,N_21911);
or U24634 (N_24634,N_20851,N_21574);
or U24635 (N_24635,N_21763,N_21257);
or U24636 (N_24636,N_20021,N_20893);
nand U24637 (N_24637,N_20002,N_21567);
nand U24638 (N_24638,N_21467,N_22263);
and U24639 (N_24639,N_21887,N_21945);
and U24640 (N_24640,N_20922,N_21548);
nor U24641 (N_24641,N_22341,N_20213);
or U24642 (N_24642,N_21754,N_22068);
nand U24643 (N_24643,N_21887,N_21653);
nand U24644 (N_24644,N_20932,N_22261);
or U24645 (N_24645,N_21559,N_21488);
nor U24646 (N_24646,N_20077,N_22206);
nor U24647 (N_24647,N_20139,N_22038);
xnor U24648 (N_24648,N_21358,N_22136);
and U24649 (N_24649,N_22468,N_21707);
or U24650 (N_24650,N_21537,N_22154);
xor U24651 (N_24651,N_21510,N_20213);
or U24652 (N_24652,N_22231,N_21933);
xnor U24653 (N_24653,N_20291,N_20888);
nor U24654 (N_24654,N_20462,N_20393);
nand U24655 (N_24655,N_22105,N_22394);
and U24656 (N_24656,N_21476,N_21196);
and U24657 (N_24657,N_20456,N_22315);
and U24658 (N_24658,N_21474,N_21360);
xor U24659 (N_24659,N_21450,N_21315);
or U24660 (N_24660,N_20839,N_21802);
xnor U24661 (N_24661,N_21809,N_22023);
or U24662 (N_24662,N_22310,N_20088);
nor U24663 (N_24663,N_20520,N_22382);
and U24664 (N_24664,N_22024,N_21600);
nand U24665 (N_24665,N_21464,N_22441);
or U24666 (N_24666,N_21809,N_20312);
and U24667 (N_24667,N_21246,N_20059);
or U24668 (N_24668,N_20481,N_21256);
nand U24669 (N_24669,N_20684,N_21102);
nor U24670 (N_24670,N_20863,N_22289);
xnor U24671 (N_24671,N_21552,N_22028);
xnor U24672 (N_24672,N_21695,N_20727);
nor U24673 (N_24673,N_21880,N_20756);
xnor U24674 (N_24674,N_21223,N_21566);
and U24675 (N_24675,N_21239,N_21197);
nand U24676 (N_24676,N_21420,N_21959);
and U24677 (N_24677,N_21951,N_21753);
or U24678 (N_24678,N_20524,N_20839);
xor U24679 (N_24679,N_21495,N_20429);
nor U24680 (N_24680,N_21439,N_21415);
nor U24681 (N_24681,N_20331,N_20912);
nor U24682 (N_24682,N_20022,N_20582);
xor U24683 (N_24683,N_20596,N_20759);
nand U24684 (N_24684,N_20948,N_21123);
xnor U24685 (N_24685,N_21845,N_21249);
and U24686 (N_24686,N_20320,N_20266);
and U24687 (N_24687,N_20532,N_21552);
nand U24688 (N_24688,N_21188,N_21556);
xor U24689 (N_24689,N_21018,N_22128);
nand U24690 (N_24690,N_20567,N_21609);
or U24691 (N_24691,N_22045,N_21849);
or U24692 (N_24692,N_22377,N_20169);
nand U24693 (N_24693,N_21757,N_21100);
or U24694 (N_24694,N_21703,N_22357);
nor U24695 (N_24695,N_20074,N_20725);
nand U24696 (N_24696,N_22125,N_22384);
and U24697 (N_24697,N_20248,N_21043);
nand U24698 (N_24698,N_21476,N_21887);
and U24699 (N_24699,N_21822,N_20086);
or U24700 (N_24700,N_21683,N_22060);
or U24701 (N_24701,N_20150,N_21468);
nand U24702 (N_24702,N_21124,N_20361);
and U24703 (N_24703,N_20763,N_20310);
xor U24704 (N_24704,N_22116,N_20861);
or U24705 (N_24705,N_20559,N_20778);
xor U24706 (N_24706,N_20744,N_20945);
nand U24707 (N_24707,N_20796,N_21672);
nand U24708 (N_24708,N_22472,N_21095);
nand U24709 (N_24709,N_21541,N_22033);
nand U24710 (N_24710,N_20803,N_20692);
nor U24711 (N_24711,N_22019,N_21148);
nor U24712 (N_24712,N_22399,N_20612);
or U24713 (N_24713,N_21982,N_20693);
or U24714 (N_24714,N_20815,N_20161);
nor U24715 (N_24715,N_20159,N_20691);
nand U24716 (N_24716,N_22148,N_20783);
or U24717 (N_24717,N_21712,N_20695);
nor U24718 (N_24718,N_22308,N_22453);
nand U24719 (N_24719,N_20851,N_20013);
and U24720 (N_24720,N_21331,N_22063);
nand U24721 (N_24721,N_20774,N_21163);
and U24722 (N_24722,N_21976,N_20948);
xnor U24723 (N_24723,N_20070,N_21307);
xor U24724 (N_24724,N_21646,N_22016);
nand U24725 (N_24725,N_22430,N_21445);
nor U24726 (N_24726,N_22106,N_22477);
xor U24727 (N_24727,N_21950,N_21853);
and U24728 (N_24728,N_21837,N_22265);
nor U24729 (N_24729,N_21652,N_20930);
nand U24730 (N_24730,N_20685,N_22237);
nand U24731 (N_24731,N_21850,N_21833);
and U24732 (N_24732,N_22200,N_21968);
and U24733 (N_24733,N_21443,N_20181);
nor U24734 (N_24734,N_21614,N_21719);
xnor U24735 (N_24735,N_20237,N_21588);
and U24736 (N_24736,N_20092,N_21946);
and U24737 (N_24737,N_21292,N_20921);
nand U24738 (N_24738,N_21578,N_20507);
or U24739 (N_24739,N_20275,N_20935);
or U24740 (N_24740,N_22168,N_21992);
nor U24741 (N_24741,N_21146,N_22481);
nand U24742 (N_24742,N_22304,N_21297);
or U24743 (N_24743,N_21342,N_20590);
nand U24744 (N_24744,N_20917,N_20325);
xor U24745 (N_24745,N_22176,N_22142);
and U24746 (N_24746,N_21015,N_21124);
and U24747 (N_24747,N_22157,N_20752);
nor U24748 (N_24748,N_21017,N_20292);
and U24749 (N_24749,N_20356,N_22433);
nand U24750 (N_24750,N_21419,N_21136);
nand U24751 (N_24751,N_21021,N_21484);
nor U24752 (N_24752,N_22022,N_22294);
or U24753 (N_24753,N_21969,N_22426);
xnor U24754 (N_24754,N_20382,N_20185);
or U24755 (N_24755,N_20174,N_20445);
nand U24756 (N_24756,N_21093,N_22419);
xor U24757 (N_24757,N_21193,N_20206);
or U24758 (N_24758,N_22448,N_22218);
and U24759 (N_24759,N_20237,N_21263);
and U24760 (N_24760,N_21959,N_20058);
nand U24761 (N_24761,N_21201,N_22249);
nand U24762 (N_24762,N_20407,N_21139);
or U24763 (N_24763,N_21961,N_20535);
and U24764 (N_24764,N_22402,N_22260);
xor U24765 (N_24765,N_20682,N_21228);
and U24766 (N_24766,N_22048,N_22376);
nor U24767 (N_24767,N_20240,N_20282);
nand U24768 (N_24768,N_20220,N_20202);
or U24769 (N_24769,N_22128,N_21684);
xor U24770 (N_24770,N_20787,N_20862);
xnor U24771 (N_24771,N_20888,N_20296);
or U24772 (N_24772,N_21283,N_21148);
nor U24773 (N_24773,N_21901,N_21684);
xor U24774 (N_24774,N_20498,N_21790);
nor U24775 (N_24775,N_20951,N_22306);
nor U24776 (N_24776,N_21066,N_21321);
nand U24777 (N_24777,N_21531,N_22469);
or U24778 (N_24778,N_20192,N_20108);
nor U24779 (N_24779,N_20517,N_21993);
nor U24780 (N_24780,N_21586,N_21639);
xor U24781 (N_24781,N_20891,N_20038);
nor U24782 (N_24782,N_20923,N_21899);
nor U24783 (N_24783,N_20047,N_20918);
nor U24784 (N_24784,N_20967,N_20362);
and U24785 (N_24785,N_22053,N_21541);
and U24786 (N_24786,N_21059,N_21211);
nor U24787 (N_24787,N_21958,N_21966);
or U24788 (N_24788,N_21912,N_21958);
nand U24789 (N_24789,N_21144,N_22341);
nand U24790 (N_24790,N_22175,N_21941);
nor U24791 (N_24791,N_22032,N_21178);
nor U24792 (N_24792,N_20426,N_20096);
xnor U24793 (N_24793,N_21090,N_22498);
xor U24794 (N_24794,N_20666,N_21784);
and U24795 (N_24795,N_20891,N_22471);
nor U24796 (N_24796,N_22453,N_20887);
xnor U24797 (N_24797,N_22051,N_20627);
nand U24798 (N_24798,N_22464,N_22322);
xor U24799 (N_24799,N_20188,N_22147);
and U24800 (N_24800,N_20571,N_21184);
xnor U24801 (N_24801,N_22313,N_20432);
or U24802 (N_24802,N_20540,N_21195);
xor U24803 (N_24803,N_20175,N_22445);
and U24804 (N_24804,N_21842,N_22364);
nand U24805 (N_24805,N_21499,N_21352);
or U24806 (N_24806,N_20972,N_21624);
or U24807 (N_24807,N_22128,N_21447);
and U24808 (N_24808,N_21526,N_20631);
nor U24809 (N_24809,N_20604,N_20860);
xor U24810 (N_24810,N_21436,N_21070);
nand U24811 (N_24811,N_20200,N_21189);
and U24812 (N_24812,N_20927,N_20014);
xor U24813 (N_24813,N_20924,N_20919);
or U24814 (N_24814,N_20288,N_22319);
or U24815 (N_24815,N_21447,N_20680);
and U24816 (N_24816,N_21949,N_21845);
or U24817 (N_24817,N_22113,N_21889);
nand U24818 (N_24818,N_20406,N_21865);
xnor U24819 (N_24819,N_20981,N_20400);
nand U24820 (N_24820,N_20848,N_20581);
or U24821 (N_24821,N_20747,N_21811);
and U24822 (N_24822,N_20525,N_21034);
and U24823 (N_24823,N_20181,N_21817);
nand U24824 (N_24824,N_20785,N_20541);
nand U24825 (N_24825,N_20979,N_22003);
xnor U24826 (N_24826,N_22446,N_22315);
nor U24827 (N_24827,N_20330,N_20380);
or U24828 (N_24828,N_20087,N_21124);
nor U24829 (N_24829,N_20940,N_21967);
and U24830 (N_24830,N_21953,N_20601);
xnor U24831 (N_24831,N_21536,N_20603);
and U24832 (N_24832,N_21381,N_21599);
or U24833 (N_24833,N_22248,N_21382);
or U24834 (N_24834,N_20761,N_21257);
or U24835 (N_24835,N_22425,N_20148);
and U24836 (N_24836,N_22197,N_21394);
or U24837 (N_24837,N_20941,N_22372);
or U24838 (N_24838,N_21680,N_21096);
xor U24839 (N_24839,N_20691,N_20960);
and U24840 (N_24840,N_21445,N_22027);
xnor U24841 (N_24841,N_20802,N_20310);
and U24842 (N_24842,N_20987,N_20741);
and U24843 (N_24843,N_21707,N_20310);
nand U24844 (N_24844,N_20892,N_22215);
and U24845 (N_24845,N_20605,N_21382);
or U24846 (N_24846,N_22499,N_21570);
or U24847 (N_24847,N_22156,N_20149);
and U24848 (N_24848,N_22363,N_20593);
nand U24849 (N_24849,N_21362,N_22189);
and U24850 (N_24850,N_22372,N_20568);
nor U24851 (N_24851,N_20842,N_21480);
nor U24852 (N_24852,N_21645,N_22411);
and U24853 (N_24853,N_20566,N_21213);
xnor U24854 (N_24854,N_21253,N_21679);
xnor U24855 (N_24855,N_20194,N_22261);
xor U24856 (N_24856,N_20895,N_22106);
xnor U24857 (N_24857,N_20832,N_21682);
nor U24858 (N_24858,N_21650,N_20613);
or U24859 (N_24859,N_20337,N_21334);
or U24860 (N_24860,N_22100,N_22340);
or U24861 (N_24861,N_22032,N_21317);
xor U24862 (N_24862,N_20497,N_20185);
xnor U24863 (N_24863,N_22443,N_21864);
nor U24864 (N_24864,N_20471,N_20098);
nand U24865 (N_24865,N_20785,N_21165);
and U24866 (N_24866,N_20417,N_20682);
and U24867 (N_24867,N_21278,N_22330);
nor U24868 (N_24868,N_20908,N_21507);
xor U24869 (N_24869,N_22000,N_22134);
or U24870 (N_24870,N_20533,N_20977);
nor U24871 (N_24871,N_20193,N_22319);
or U24872 (N_24872,N_20629,N_22058);
and U24873 (N_24873,N_22136,N_21487);
nand U24874 (N_24874,N_21750,N_21851);
xor U24875 (N_24875,N_21752,N_21718);
xnor U24876 (N_24876,N_20259,N_20217);
nand U24877 (N_24877,N_21081,N_22420);
nor U24878 (N_24878,N_21387,N_20743);
and U24879 (N_24879,N_20277,N_21396);
nor U24880 (N_24880,N_21320,N_20257);
xnor U24881 (N_24881,N_21557,N_20527);
nor U24882 (N_24882,N_21754,N_22320);
nor U24883 (N_24883,N_20833,N_21149);
nor U24884 (N_24884,N_21618,N_20451);
nor U24885 (N_24885,N_21941,N_21640);
xor U24886 (N_24886,N_20736,N_21723);
nand U24887 (N_24887,N_22476,N_20021);
nor U24888 (N_24888,N_22419,N_20244);
and U24889 (N_24889,N_21719,N_21770);
and U24890 (N_24890,N_21854,N_21568);
xor U24891 (N_24891,N_22335,N_20001);
nor U24892 (N_24892,N_21071,N_21995);
or U24893 (N_24893,N_21024,N_22048);
xnor U24894 (N_24894,N_20470,N_21900);
or U24895 (N_24895,N_21884,N_21662);
and U24896 (N_24896,N_21432,N_22204);
or U24897 (N_24897,N_22437,N_21895);
nand U24898 (N_24898,N_22314,N_21097);
xnor U24899 (N_24899,N_21157,N_20591);
nand U24900 (N_24900,N_21114,N_21951);
nor U24901 (N_24901,N_20603,N_21951);
or U24902 (N_24902,N_20433,N_20057);
and U24903 (N_24903,N_22140,N_22295);
and U24904 (N_24904,N_20100,N_20055);
nand U24905 (N_24905,N_21913,N_21201);
xnor U24906 (N_24906,N_21666,N_20817);
nor U24907 (N_24907,N_21052,N_21832);
xnor U24908 (N_24908,N_20019,N_20477);
xor U24909 (N_24909,N_21327,N_21162);
nand U24910 (N_24910,N_21653,N_20490);
and U24911 (N_24911,N_21744,N_22071);
and U24912 (N_24912,N_22255,N_22274);
and U24913 (N_24913,N_20904,N_21710);
or U24914 (N_24914,N_21297,N_21667);
xor U24915 (N_24915,N_20323,N_20519);
nand U24916 (N_24916,N_21838,N_20532);
xor U24917 (N_24917,N_22449,N_20086);
or U24918 (N_24918,N_21030,N_22291);
xnor U24919 (N_24919,N_20199,N_22359);
nor U24920 (N_24920,N_20832,N_20257);
nand U24921 (N_24921,N_21989,N_22362);
nor U24922 (N_24922,N_21888,N_22193);
or U24923 (N_24923,N_20359,N_20455);
or U24924 (N_24924,N_22230,N_21896);
xor U24925 (N_24925,N_21914,N_21242);
nand U24926 (N_24926,N_20371,N_20544);
and U24927 (N_24927,N_21979,N_21453);
nand U24928 (N_24928,N_22426,N_20019);
nand U24929 (N_24929,N_22228,N_21961);
nor U24930 (N_24930,N_21844,N_20833);
xor U24931 (N_24931,N_20790,N_21710);
and U24932 (N_24932,N_20963,N_21340);
xor U24933 (N_24933,N_20640,N_20878);
and U24934 (N_24934,N_20595,N_21509);
xnor U24935 (N_24935,N_21394,N_22199);
or U24936 (N_24936,N_20429,N_22035);
or U24937 (N_24937,N_21447,N_20041);
nor U24938 (N_24938,N_21215,N_22440);
nand U24939 (N_24939,N_22404,N_21428);
or U24940 (N_24940,N_20852,N_20030);
or U24941 (N_24941,N_20607,N_22272);
and U24942 (N_24942,N_21529,N_21173);
nor U24943 (N_24943,N_20953,N_20474);
nor U24944 (N_24944,N_20306,N_22284);
nor U24945 (N_24945,N_20019,N_20104);
xor U24946 (N_24946,N_21106,N_21385);
and U24947 (N_24947,N_21830,N_21551);
xnor U24948 (N_24948,N_20331,N_20671);
or U24949 (N_24949,N_20487,N_21813);
and U24950 (N_24950,N_20575,N_22285);
or U24951 (N_24951,N_21898,N_21229);
nand U24952 (N_24952,N_21780,N_20210);
nor U24953 (N_24953,N_21448,N_20117);
xor U24954 (N_24954,N_21717,N_22280);
or U24955 (N_24955,N_20082,N_20999);
or U24956 (N_24956,N_20307,N_21723);
nor U24957 (N_24957,N_21494,N_21964);
and U24958 (N_24958,N_21498,N_20175);
nor U24959 (N_24959,N_20051,N_20908);
xnor U24960 (N_24960,N_20352,N_21760);
nor U24961 (N_24961,N_20347,N_20717);
nor U24962 (N_24962,N_21441,N_20710);
xnor U24963 (N_24963,N_21007,N_20475);
nor U24964 (N_24964,N_20715,N_20666);
nand U24965 (N_24965,N_22080,N_21791);
xor U24966 (N_24966,N_20558,N_20568);
and U24967 (N_24967,N_22083,N_20606);
xor U24968 (N_24968,N_20380,N_20483);
and U24969 (N_24969,N_20244,N_20074);
and U24970 (N_24970,N_22114,N_21033);
nand U24971 (N_24971,N_22276,N_21597);
or U24972 (N_24972,N_20373,N_21930);
nor U24973 (N_24973,N_21269,N_21604);
nand U24974 (N_24974,N_21448,N_20676);
nand U24975 (N_24975,N_20867,N_20361);
or U24976 (N_24976,N_21275,N_20517);
or U24977 (N_24977,N_21569,N_20959);
nand U24978 (N_24978,N_22274,N_20977);
and U24979 (N_24979,N_20267,N_21332);
or U24980 (N_24980,N_22091,N_22318);
and U24981 (N_24981,N_21498,N_22348);
xnor U24982 (N_24982,N_21144,N_21733);
and U24983 (N_24983,N_21233,N_20250);
or U24984 (N_24984,N_20077,N_21427);
nand U24985 (N_24985,N_22019,N_21538);
or U24986 (N_24986,N_21117,N_21887);
or U24987 (N_24987,N_20834,N_20461);
xor U24988 (N_24988,N_21894,N_20420);
and U24989 (N_24989,N_21690,N_20392);
xnor U24990 (N_24990,N_21031,N_20833);
nor U24991 (N_24991,N_20443,N_20727);
nor U24992 (N_24992,N_21003,N_20934);
nor U24993 (N_24993,N_20777,N_20568);
nor U24994 (N_24994,N_20557,N_21353);
and U24995 (N_24995,N_21899,N_20124);
or U24996 (N_24996,N_20614,N_21702);
or U24997 (N_24997,N_22171,N_20143);
or U24998 (N_24998,N_21016,N_21707);
nor U24999 (N_24999,N_21376,N_22163);
or UO_0 (O_0,N_24980,N_23579);
nand UO_1 (O_1,N_24152,N_23760);
xor UO_2 (O_2,N_23067,N_23309);
or UO_3 (O_3,N_22952,N_23127);
or UO_4 (O_4,N_24296,N_24375);
nor UO_5 (O_5,N_23892,N_24680);
nand UO_6 (O_6,N_24094,N_24808);
nor UO_7 (O_7,N_24549,N_22532);
nand UO_8 (O_8,N_23815,N_24718);
and UO_9 (O_9,N_22713,N_23420);
and UO_10 (O_10,N_23981,N_23820);
xnor UO_11 (O_11,N_23507,N_24875);
or UO_12 (O_12,N_22630,N_22628);
xnor UO_13 (O_13,N_22923,N_23167);
and UO_14 (O_14,N_22771,N_23359);
nor UO_15 (O_15,N_24521,N_24091);
nand UO_16 (O_16,N_24456,N_22649);
nand UO_17 (O_17,N_23193,N_23519);
and UO_18 (O_18,N_22530,N_23584);
nor UO_19 (O_19,N_24298,N_24915);
xor UO_20 (O_20,N_22586,N_24999);
and UO_21 (O_21,N_23395,N_23231);
and UO_22 (O_22,N_23611,N_23479);
nand UO_23 (O_23,N_23692,N_23762);
xnor UO_24 (O_24,N_23389,N_24837);
nor UO_25 (O_25,N_23713,N_23152);
xnor UO_26 (O_26,N_24936,N_24839);
xnor UO_27 (O_27,N_22857,N_23633);
nand UO_28 (O_28,N_24367,N_23012);
and UO_29 (O_29,N_23696,N_23266);
nand UO_30 (O_30,N_23553,N_24608);
or UO_31 (O_31,N_23404,N_24586);
xor UO_32 (O_32,N_24410,N_22892);
nand UO_33 (O_33,N_24990,N_24024);
or UO_34 (O_34,N_22871,N_24672);
and UO_35 (O_35,N_24222,N_23483);
nor UO_36 (O_36,N_24426,N_24106);
and UO_37 (O_37,N_23041,N_23379);
xor UO_38 (O_38,N_22656,N_24598);
nand UO_39 (O_39,N_24989,N_24658);
nand UO_40 (O_40,N_22813,N_23213);
or UO_41 (O_41,N_23077,N_23333);
or UO_42 (O_42,N_23651,N_24919);
or UO_43 (O_43,N_24757,N_23863);
nand UO_44 (O_44,N_22880,N_24218);
or UO_45 (O_45,N_24967,N_24749);
or UO_46 (O_46,N_22693,N_22531);
nor UO_47 (O_47,N_23295,N_24340);
and UO_48 (O_48,N_22641,N_22977);
and UO_49 (O_49,N_22972,N_23272);
xor UO_50 (O_50,N_23367,N_23150);
nor UO_51 (O_51,N_23253,N_24402);
or UO_52 (O_52,N_24711,N_23572);
and UO_53 (O_53,N_23598,N_23925);
and UO_54 (O_54,N_23825,N_24626);
or UO_55 (O_55,N_23997,N_24813);
nand UO_56 (O_56,N_22775,N_23455);
xnor UO_57 (O_57,N_23637,N_24307);
nand UO_58 (O_58,N_23618,N_23619);
xor UO_59 (O_59,N_24113,N_22637);
and UO_60 (O_60,N_22593,N_23254);
xnor UO_61 (O_61,N_24362,N_24075);
nor UO_62 (O_62,N_24349,N_22999);
xor UO_63 (O_63,N_23813,N_22779);
or UO_64 (O_64,N_24134,N_24700);
nor UO_65 (O_65,N_24171,N_23774);
nand UO_66 (O_66,N_24125,N_24484);
nand UO_67 (O_67,N_24578,N_23234);
nand UO_68 (O_68,N_22796,N_23019);
xnor UO_69 (O_69,N_23612,N_22602);
or UO_70 (O_70,N_24565,N_24946);
or UO_71 (O_71,N_22956,N_22581);
nor UO_72 (O_72,N_23228,N_23614);
and UO_73 (O_73,N_24668,N_24940);
or UO_74 (O_74,N_24846,N_24883);
and UO_75 (O_75,N_24379,N_23917);
nand UO_76 (O_76,N_22823,N_23967);
xnor UO_77 (O_77,N_24916,N_24845);
nor UO_78 (O_78,N_24269,N_23375);
nor UO_79 (O_79,N_24929,N_22691);
and UO_80 (O_80,N_23861,N_23057);
xor UO_81 (O_81,N_23730,N_22543);
nand UO_82 (O_82,N_23529,N_22720);
nand UO_83 (O_83,N_23064,N_22618);
nor UO_84 (O_84,N_22583,N_22712);
nand UO_85 (O_85,N_24086,N_23165);
nor UO_86 (O_86,N_24646,N_23946);
xor UO_87 (O_87,N_24329,N_24247);
nand UO_88 (O_88,N_24754,N_24544);
nand UO_89 (O_89,N_24099,N_23973);
and UO_90 (O_90,N_24158,N_23889);
and UO_91 (O_91,N_22559,N_22978);
nand UO_92 (O_92,N_23293,N_23400);
nor UO_93 (O_93,N_24976,N_24770);
nand UO_94 (O_94,N_24717,N_24424);
nand UO_95 (O_95,N_23025,N_22590);
nor UO_96 (O_96,N_24029,N_24290);
nand UO_97 (O_97,N_23303,N_23235);
or UO_98 (O_98,N_22874,N_23444);
xor UO_99 (O_99,N_24007,N_23194);
nand UO_100 (O_100,N_22560,N_22708);
nand UO_101 (O_101,N_24870,N_24283);
and UO_102 (O_102,N_24681,N_23219);
nand UO_103 (O_103,N_24862,N_23036);
nor UO_104 (O_104,N_23366,N_22899);
or UO_105 (O_105,N_22534,N_24743);
xnor UO_106 (O_106,N_24631,N_23856);
or UO_107 (O_107,N_24535,N_23123);
nand UO_108 (O_108,N_24339,N_24965);
or UO_109 (O_109,N_23211,N_24263);
and UO_110 (O_110,N_24249,N_23725);
nand UO_111 (O_111,N_23847,N_24709);
nand UO_112 (O_112,N_24244,N_23242);
and UO_113 (O_113,N_23520,N_23987);
nor UO_114 (O_114,N_23573,N_24702);
nand UO_115 (O_115,N_23363,N_24713);
or UO_116 (O_116,N_24648,N_23260);
and UO_117 (O_117,N_23864,N_24895);
nor UO_118 (O_118,N_22808,N_22938);
and UO_119 (O_119,N_24274,N_24464);
xor UO_120 (O_120,N_23467,N_23884);
nor UO_121 (O_121,N_22647,N_22685);
and UO_122 (O_122,N_22679,N_23620);
xor UO_123 (O_123,N_22844,N_23907);
and UO_124 (O_124,N_23498,N_23080);
and UO_125 (O_125,N_23735,N_24245);
or UO_126 (O_126,N_24460,N_24416);
nor UO_127 (O_127,N_22518,N_24315);
nand UO_128 (O_128,N_22984,N_23328);
nand UO_129 (O_129,N_23597,N_23671);
or UO_130 (O_130,N_24667,N_22895);
nor UO_131 (O_131,N_24949,N_23823);
xnor UO_132 (O_132,N_23758,N_24401);
nand UO_133 (O_133,N_24440,N_23493);
nand UO_134 (O_134,N_23175,N_24594);
xnor UO_135 (O_135,N_23416,N_23294);
xnor UO_136 (O_136,N_24259,N_24868);
or UO_137 (O_137,N_23163,N_22655);
nor UO_138 (O_138,N_24975,N_24825);
xor UO_139 (O_139,N_22785,N_23218);
and UO_140 (O_140,N_24695,N_24467);
or UO_141 (O_141,N_23459,N_22665);
nor UO_142 (O_142,N_24475,N_24746);
nor UO_143 (O_143,N_22615,N_22961);
or UO_144 (O_144,N_24877,N_24356);
or UO_145 (O_145,N_24554,N_24986);
nor UO_146 (O_146,N_23670,N_23866);
nand UO_147 (O_147,N_23723,N_23587);
nor UO_148 (O_148,N_24129,N_22503);
xnor UO_149 (O_149,N_24924,N_23939);
nand UO_150 (O_150,N_22768,N_24120);
xor UO_151 (O_151,N_23608,N_24122);
xnor UO_152 (O_152,N_22730,N_23792);
nand UO_153 (O_153,N_24844,N_24449);
and UO_154 (O_154,N_24812,N_22616);
or UO_155 (O_155,N_24637,N_24536);
nand UO_156 (O_156,N_24719,N_24133);
nand UO_157 (O_157,N_23296,N_22709);
or UO_158 (O_158,N_24557,N_23126);
nand UO_159 (O_159,N_24450,N_24607);
and UO_160 (O_160,N_24179,N_22798);
or UO_161 (O_161,N_22927,N_23945);
nor UO_162 (O_162,N_22722,N_23320);
and UO_163 (O_163,N_22941,N_22642);
or UO_164 (O_164,N_22930,N_24865);
xnor UO_165 (O_165,N_24435,N_22933);
xnor UO_166 (O_166,N_22605,N_24144);
xnor UO_167 (O_167,N_22867,N_23311);
nor UO_168 (O_168,N_22887,N_23094);
xnor UO_169 (O_169,N_24497,N_24828);
or UO_170 (O_170,N_23341,N_24323);
xor UO_171 (O_171,N_24013,N_23256);
and UO_172 (O_172,N_23771,N_24156);
and UO_173 (O_173,N_23969,N_23702);
nand UO_174 (O_174,N_23712,N_22985);
or UO_175 (O_175,N_23852,N_24590);
and UO_176 (O_176,N_24137,N_24320);
and UO_177 (O_177,N_24398,N_24944);
and UO_178 (O_178,N_22793,N_22717);
nand UO_179 (O_179,N_23594,N_24414);
and UO_180 (O_180,N_22815,N_23837);
and UO_181 (O_181,N_24425,N_22663);
nand UO_182 (O_182,N_23984,N_23943);
or UO_183 (O_183,N_22633,N_23634);
or UO_184 (O_184,N_23737,N_23107);
xor UO_185 (O_185,N_23525,N_22811);
or UO_186 (O_186,N_23665,N_22851);
or UO_187 (O_187,N_23136,N_24933);
nand UO_188 (O_188,N_22750,N_23415);
and UO_189 (O_189,N_23728,N_23096);
nor UO_190 (O_190,N_24026,N_24161);
and UO_191 (O_191,N_23583,N_24921);
and UO_192 (O_192,N_22542,N_24686);
and UO_193 (O_193,N_23916,N_24817);
and UO_194 (O_194,N_23487,N_23803);
or UO_195 (O_195,N_23691,N_23489);
nand UO_196 (O_196,N_24885,N_24553);
and UO_197 (O_197,N_23909,N_24318);
and UO_198 (O_198,N_23548,N_23840);
xor UO_199 (O_199,N_23870,N_24337);
nor UO_200 (O_200,N_23334,N_24308);
or UO_201 (O_201,N_22558,N_24173);
nand UO_202 (O_202,N_23893,N_22746);
nor UO_203 (O_203,N_23139,N_23667);
nand UO_204 (O_204,N_24305,N_23143);
xnor UO_205 (O_205,N_24714,N_24601);
and UO_206 (O_206,N_24853,N_24392);
xnor UO_207 (O_207,N_23247,N_22963);
nand UO_208 (O_208,N_24254,N_23227);
nand UO_209 (O_209,N_22986,N_24493);
or UO_210 (O_210,N_23120,N_22613);
or UO_211 (O_211,N_24645,N_24124);
nor UO_212 (O_212,N_23441,N_22789);
nor UO_213 (O_213,N_24240,N_24139);
or UO_214 (O_214,N_24831,N_22580);
or UO_215 (O_215,N_24256,N_24927);
or UO_216 (O_216,N_23274,N_23091);
nor UO_217 (O_217,N_22838,N_24063);
nor UO_218 (O_218,N_24533,N_24708);
nand UO_219 (O_219,N_24468,N_23115);
and UO_220 (O_220,N_23768,N_23576);
and UO_221 (O_221,N_24203,N_24176);
xnor UO_222 (O_222,N_24515,N_22918);
and UO_223 (O_223,N_24353,N_23027);
nand UO_224 (O_224,N_22758,N_23271);
nand UO_225 (O_225,N_23468,N_23518);
and UO_226 (O_226,N_22620,N_23054);
nor UO_227 (O_227,N_24181,N_23899);
xor UO_228 (O_228,N_24232,N_22890);
nand UO_229 (O_229,N_23411,N_23330);
nand UO_230 (O_230,N_23878,N_22736);
or UO_231 (O_231,N_23921,N_23699);
and UO_232 (O_232,N_23196,N_23674);
nor UO_233 (O_233,N_24923,N_24728);
xnor UO_234 (O_234,N_23440,N_23908);
nand UO_235 (O_235,N_24209,N_23537);
xnor UO_236 (O_236,N_23650,N_24178);
nand UO_237 (O_237,N_24331,N_23490);
and UO_238 (O_238,N_24282,N_24640);
xnor UO_239 (O_239,N_23010,N_23135);
nand UO_240 (O_240,N_24603,N_24233);
xnor UO_241 (O_241,N_23076,N_22925);
xor UO_242 (O_242,N_22849,N_24386);
or UO_243 (O_243,N_23159,N_23541);
nand UO_244 (O_244,N_24409,N_23239);
and UO_245 (O_245,N_23391,N_23024);
xnor UO_246 (O_246,N_24740,N_24248);
and UO_247 (O_247,N_22847,N_23613);
or UO_248 (O_248,N_24587,N_23668);
xnor UO_249 (O_249,N_24294,N_24145);
or UO_250 (O_250,N_23811,N_24052);
and UO_251 (O_251,N_24316,N_23049);
nand UO_252 (O_252,N_22910,N_24077);
nand UO_253 (O_253,N_23185,N_23170);
nor UO_254 (O_254,N_23063,N_22919);
nand UO_255 (O_255,N_22760,N_22929);
and UO_256 (O_256,N_22776,N_22512);
xnor UO_257 (O_257,N_23406,N_24734);
or UO_258 (O_258,N_23432,N_23681);
nor UO_259 (O_259,N_24751,N_24599);
nor UO_260 (O_260,N_23134,N_24031);
or UO_261 (O_261,N_24665,N_22585);
or UO_262 (O_262,N_23661,N_24074);
xor UO_263 (O_263,N_24583,N_22826);
and UO_264 (O_264,N_24429,N_24733);
nor UO_265 (O_265,N_24773,N_23308);
and UO_266 (O_266,N_24832,N_24012);
or UO_267 (O_267,N_24228,N_22519);
nor UO_268 (O_268,N_24299,N_22644);
nand UO_269 (O_269,N_22799,N_24487);
xnor UO_270 (O_270,N_24168,N_23220);
and UO_271 (O_271,N_23933,N_23377);
xnor UO_272 (O_272,N_23316,N_23471);
or UO_273 (O_273,N_23184,N_24874);
and UO_274 (O_274,N_24059,N_22646);
nand UO_275 (O_275,N_23644,N_23515);
nand UO_276 (O_276,N_22676,N_22928);
nand UO_277 (O_277,N_23051,N_24350);
xor UO_278 (O_278,N_22787,N_23215);
or UO_279 (O_279,N_24403,N_23779);
nor UO_280 (O_280,N_24042,N_24199);
nand UO_281 (O_281,N_24676,N_24462);
xnor UO_282 (O_282,N_22660,N_23977);
xor UO_283 (O_283,N_22595,N_23302);
nor UO_284 (O_284,N_23474,N_22802);
nor UO_285 (O_285,N_23996,N_24572);
and UO_286 (O_286,N_24663,N_23844);
xnor UO_287 (O_287,N_23182,N_22594);
nor UO_288 (O_288,N_23424,N_22979);
or UO_289 (O_289,N_23731,N_23224);
or UO_290 (O_290,N_22636,N_23764);
nor UO_291 (O_291,N_22924,N_22848);
and UO_292 (O_292,N_22725,N_22862);
nor UO_293 (O_293,N_23003,N_24242);
or UO_294 (O_294,N_24898,N_23890);
xor UO_295 (O_295,N_24098,N_23105);
and UO_296 (O_296,N_24067,N_23876);
and UO_297 (O_297,N_23141,N_24302);
or UO_298 (O_298,N_23947,N_22764);
or UO_299 (O_299,N_22962,N_23935);
and UO_300 (O_300,N_23007,N_22909);
xor UO_301 (O_301,N_23156,N_22711);
nand UO_302 (O_302,N_23606,N_24060);
nand UO_303 (O_303,N_24706,N_24418);
and UO_304 (O_304,N_22990,N_23694);
nand UO_305 (O_305,N_24739,N_23664);
nor UO_306 (O_306,N_22772,N_23124);
or UO_307 (O_307,N_23875,N_24900);
and UO_308 (O_308,N_24902,N_22666);
nor UO_309 (O_309,N_24476,N_24478);
or UO_310 (O_310,N_22680,N_23564);
or UO_311 (O_311,N_22840,N_24100);
nand UO_312 (O_312,N_23649,N_23682);
xnor UO_313 (O_313,N_23394,N_23970);
or UO_314 (O_314,N_24201,N_23172);
nor UO_315 (O_315,N_23477,N_24495);
nand UO_316 (O_316,N_23070,N_24576);
nor UO_317 (O_317,N_23798,N_23258);
nand UO_318 (O_318,N_24503,N_22675);
nor UO_319 (O_319,N_23140,N_23817);
nand UO_320 (O_320,N_23031,N_22548);
nand UO_321 (O_321,N_24281,N_24771);
nor UO_322 (O_322,N_24744,N_23784);
and UO_323 (O_323,N_24239,N_24022);
and UO_324 (O_324,N_24028,N_24219);
and UO_325 (O_325,N_23555,N_24348);
nor UO_326 (O_326,N_24689,N_23512);
and UO_327 (O_327,N_24035,N_23425);
nor UO_328 (O_328,N_22882,N_23419);
nand UO_329 (O_329,N_24579,N_23918);
and UO_330 (O_330,N_23563,N_23666);
and UO_331 (O_331,N_23009,N_23625);
or UO_332 (O_332,N_22582,N_22915);
nor UO_333 (O_333,N_24712,N_22721);
nor UO_334 (O_334,N_24947,N_22546);
nand UO_335 (O_335,N_24692,N_24146);
nand UO_336 (O_336,N_23885,N_22975);
or UO_337 (O_337,N_24559,N_24840);
or UO_338 (O_338,N_22669,N_23733);
and UO_339 (O_339,N_23785,N_23950);
xnor UO_340 (O_340,N_24538,N_23125);
nor UO_341 (O_341,N_22726,N_23292);
nand UO_342 (O_342,N_23362,N_24529);
or UO_343 (O_343,N_24661,N_23151);
nor UO_344 (O_344,N_23755,N_23998);
or UO_345 (O_345,N_23090,N_23089);
nand UO_346 (O_346,N_24395,N_23033);
nor UO_347 (O_347,N_24796,N_23566);
or UO_348 (O_348,N_24987,N_23062);
and UO_349 (O_349,N_24612,N_23045);
nor UO_350 (O_350,N_23804,N_24969);
nor UO_351 (O_351,N_22770,N_24730);
and UO_352 (O_352,N_24102,N_24285);
xor UO_353 (O_353,N_23248,N_24729);
xnor UO_354 (O_354,N_23800,N_24230);
nand UO_355 (O_355,N_23475,N_23093);
nand UO_356 (O_356,N_23204,N_23208);
or UO_357 (O_357,N_23679,N_24268);
nor UO_358 (O_358,N_23903,N_23137);
nor UO_359 (O_359,N_23491,N_24422);
nor UO_360 (O_360,N_22723,N_24621);
and UO_361 (O_361,N_22836,N_24473);
and UO_362 (O_362,N_22830,N_22877);
xnor UO_363 (O_363,N_23868,N_23663);
nand UO_364 (O_364,N_24342,N_24800);
nand UO_365 (O_365,N_23562,N_24160);
and UO_366 (O_366,N_22705,N_22997);
nor UO_367 (O_367,N_24913,N_23605);
and UO_368 (O_368,N_24271,N_24326);
xnor UO_369 (O_369,N_22936,N_23853);
nand UO_370 (O_370,N_23567,N_24439);
or UO_371 (O_371,N_22506,N_23516);
or UO_372 (O_372,N_24463,N_24447);
xnor UO_373 (O_373,N_22964,N_22747);
or UO_374 (O_374,N_23534,N_24205);
and UO_375 (O_375,N_24408,N_24480);
xnor UO_376 (O_376,N_23205,N_23277);
nor UO_377 (O_377,N_24566,N_24723);
nand UO_378 (O_378,N_23078,N_22607);
nor UO_379 (O_379,N_23810,N_22629);
nor UO_380 (O_380,N_22881,N_23177);
nand UO_381 (O_381,N_23287,N_23032);
and UO_382 (O_382,N_24202,N_23412);
nor UO_383 (O_383,N_22588,N_24011);
nor UO_384 (O_384,N_23683,N_23148);
nand UO_385 (O_385,N_22780,N_24289);
xor UO_386 (O_386,N_23550,N_23020);
or UO_387 (O_387,N_23857,N_23504);
or UO_388 (O_388,N_23403,N_23826);
and UO_389 (O_389,N_23638,N_23753);
and UO_390 (O_390,N_24284,N_24998);
nor UO_391 (O_391,N_24888,N_24679);
nand UO_392 (O_392,N_24255,N_24455);
xnor UO_393 (O_393,N_23531,N_22944);
nor UO_394 (O_394,N_24136,N_23206);
and UO_395 (O_395,N_23259,N_23799);
nor UO_396 (O_396,N_23326,N_24630);
nand UO_397 (O_397,N_22606,N_23600);
or UO_398 (O_398,N_24266,N_24351);
nor UO_399 (O_399,N_24185,N_24606);
nand UO_400 (O_400,N_24864,N_23348);
xor UO_401 (O_401,N_24653,N_23279);
or UO_402 (O_402,N_22983,N_24685);
nand UO_403 (O_403,N_23680,N_23354);
and UO_404 (O_404,N_24014,N_23435);
or UO_405 (O_405,N_24928,N_23250);
or UO_406 (O_406,N_23190,N_23662);
xor UO_407 (O_407,N_22673,N_22571);
xnor UO_408 (O_408,N_22741,N_24246);
and UO_409 (O_409,N_24991,N_22732);
nor UO_410 (O_410,N_23321,N_23743);
xnor UO_411 (O_411,N_23687,N_23936);
and UO_412 (O_412,N_23542,N_24520);
and UO_413 (O_413,N_24212,N_24815);
and UO_414 (O_414,N_24526,N_24677);
or UO_415 (O_415,N_24643,N_23988);
xnor UO_416 (O_416,N_24126,N_23299);
xor UO_417 (O_417,N_23690,N_22550);
and UO_418 (O_418,N_22539,N_22869);
or UO_419 (O_419,N_24541,N_24779);
or UO_420 (O_420,N_22812,N_23898);
or UO_421 (O_421,N_24964,N_24261);
nor UO_422 (O_422,N_24169,N_23047);
xnor UO_423 (O_423,N_24293,N_22687);
and UO_424 (O_424,N_24797,N_24225);
and UO_425 (O_425,N_22591,N_23241);
or UO_426 (O_426,N_24527,N_23154);
and UO_427 (O_427,N_23888,N_24431);
or UO_428 (O_428,N_23437,N_22966);
or UO_429 (O_429,N_24448,N_24978);
xor UO_430 (O_430,N_23016,N_22727);
nor UO_431 (O_431,N_23747,N_23886);
xor UO_432 (O_432,N_24427,N_24823);
nand UO_433 (O_433,N_23609,N_22957);
nand UO_434 (O_434,N_23181,N_23413);
and UO_435 (O_435,N_24119,N_23160);
nand UO_436 (O_436,N_23631,N_24413);
xnor UO_437 (O_437,N_23581,N_24019);
and UO_438 (O_438,N_23543,N_22751);
or UO_439 (O_439,N_24260,N_24968);
and UO_440 (O_440,N_24433,N_24363);
nor UO_441 (O_441,N_23353,N_22597);
nand UO_442 (O_442,N_24937,N_23186);
and UO_443 (O_443,N_22937,N_23993);
xnor UO_444 (O_444,N_24701,N_24932);
nor UO_445 (O_445,N_24802,N_22959);
nand UO_446 (O_446,N_23439,N_24569);
and UO_447 (O_447,N_23372,N_24693);
or UO_448 (O_448,N_23369,N_22541);
xnor UO_449 (O_449,N_23161,N_24444);
or UO_450 (O_450,N_23867,N_22853);
nor UO_451 (O_451,N_24666,N_23715);
xor UO_452 (O_452,N_23615,N_22843);
nand UO_453 (O_453,N_24217,N_24341);
or UO_454 (O_454,N_23118,N_24385);
nand UO_455 (O_455,N_24047,N_23307);
and UO_456 (O_456,N_23523,N_23698);
nand UO_457 (O_457,N_24258,N_23937);
xnor UO_458 (O_458,N_24938,N_24381);
nand UO_459 (O_459,N_24162,N_22540);
and UO_460 (O_460,N_23653,N_24200);
xnor UO_461 (O_461,N_24180,N_22701);
and UO_462 (O_462,N_24798,N_23245);
xor UO_463 (O_463,N_23270,N_23111);
nand UO_464 (O_464,N_23133,N_23360);
or UO_465 (O_465,N_24903,N_22600);
and UO_466 (O_466,N_22931,N_23102);
and UO_467 (O_467,N_24909,N_24871);
and UO_468 (O_468,N_23109,N_24390);
xor UO_469 (O_469,N_23500,N_22729);
xnor UO_470 (O_470,N_24304,N_23342);
and UO_471 (O_471,N_24384,N_24826);
xnor UO_472 (O_472,N_24278,N_24352);
or UO_473 (O_473,N_23176,N_24436);
nor UO_474 (O_474,N_24703,N_24918);
xor UO_475 (O_475,N_24108,N_23724);
nor UO_476 (O_476,N_22551,N_24881);
or UO_477 (O_477,N_24010,N_24112);
or UO_478 (O_478,N_22835,N_23450);
xnor UO_479 (O_479,N_23763,N_23282);
or UO_480 (O_480,N_22992,N_23081);
and UO_481 (O_481,N_24234,N_23897);
xor UO_482 (O_482,N_24405,N_24369);
or UO_483 (O_483,N_22858,N_23630);
nand UO_484 (O_484,N_24490,N_24966);
and UO_485 (O_485,N_23805,N_24333);
and UO_486 (O_486,N_24303,N_23560);
xnor UO_487 (O_487,N_22870,N_23381);
xnor UO_488 (O_488,N_24581,N_22831);
and UO_489 (O_489,N_24330,N_23203);
xnor UO_490 (O_490,N_24452,N_22536);
and UO_491 (O_491,N_22570,N_24505);
xnor UO_492 (O_492,N_23405,N_24006);
nand UO_493 (O_493,N_23574,N_23195);
and UO_494 (O_494,N_24534,N_24984);
or UO_495 (O_495,N_24453,N_22562);
and UO_496 (O_496,N_24788,N_24361);
xnor UO_497 (O_497,N_24277,N_23658);
or UO_498 (O_498,N_24641,N_24492);
xnor UO_499 (O_499,N_23773,N_23188);
nor UO_500 (O_500,N_23465,N_23071);
and UO_501 (O_501,N_23072,N_24037);
nand UO_502 (O_502,N_24753,N_23187);
or UO_503 (O_503,N_22696,N_24707);
and UO_504 (O_504,N_22773,N_23854);
nor UO_505 (O_505,N_24210,N_24270);
nor UO_506 (O_506,N_24147,N_22883);
xor UO_507 (O_507,N_23261,N_23660);
nor UO_508 (O_508,N_24214,N_22537);
xnor UO_509 (O_509,N_22516,N_22561);
nor UO_510 (O_510,N_23859,N_23376);
and UO_511 (O_511,N_23438,N_22752);
nor UO_512 (O_512,N_24215,N_24170);
and UO_513 (O_513,N_23951,N_24821);
and UO_514 (O_514,N_23278,N_24878);
nand UO_515 (O_515,N_23722,N_22837);
nand UO_516 (O_516,N_24292,N_24629);
xor UO_517 (O_517,N_23485,N_24722);
or UO_518 (O_518,N_24310,N_24041);
or UO_519 (O_519,N_24880,N_22653);
xor UO_520 (O_520,N_24571,N_23879);
and UO_521 (O_521,N_23315,N_22971);
xnor UO_522 (O_522,N_22563,N_24604);
xor UO_523 (O_523,N_23848,N_24636);
and UO_524 (O_524,N_24795,N_23838);
or UO_525 (O_525,N_24118,N_22599);
nand UO_526 (O_526,N_22839,N_22715);
nand UO_527 (O_527,N_23648,N_24507);
and UO_528 (O_528,N_23845,N_23265);
or UO_529 (O_529,N_24889,N_23214);
and UO_530 (O_530,N_24755,N_23818);
and UO_531 (O_531,N_22612,N_24671);
xnor UO_532 (O_532,N_23461,N_24324);
or UO_533 (O_533,N_24872,N_24030);
or UO_534 (O_534,N_23991,N_24286);
nor UO_535 (O_535,N_23877,N_24142);
nor UO_536 (O_536,N_24725,N_22935);
or UO_537 (O_537,N_24994,N_22697);
xor UO_538 (O_538,N_24803,N_23767);
nand UO_539 (O_539,N_24765,N_24869);
xor UO_540 (O_540,N_23891,N_22584);
nand UO_541 (O_541,N_22645,N_23517);
and UO_542 (O_542,N_24981,N_24208);
nand UO_543 (O_543,N_24632,N_23551);
and UO_544 (O_544,N_23912,N_24738);
or UO_545 (O_545,N_22589,N_23314);
nor UO_546 (O_546,N_22619,N_24742);
or UO_547 (O_547,N_24627,N_23855);
nand UO_548 (O_548,N_22995,N_23029);
or UO_549 (O_549,N_24782,N_23338);
and UO_550 (O_550,N_23824,N_22670);
nor UO_551 (O_551,N_24951,N_22716);
xor UO_552 (O_552,N_24894,N_23797);
or UO_553 (O_553,N_24300,N_23590);
nor UO_554 (O_554,N_24461,N_24731);
or UO_555 (O_555,N_24620,N_24345);
xnor UO_556 (O_556,N_23742,N_22791);
and UO_557 (O_557,N_23189,N_23789);
nor UO_558 (O_558,N_23162,N_23358);
or UO_559 (O_559,N_22681,N_24758);
or UO_560 (O_560,N_23496,N_24992);
or UO_561 (O_561,N_24135,N_24023);
nor UO_562 (O_562,N_23494,N_22769);
or UO_563 (O_563,N_23941,N_23568);
nand UO_564 (O_564,N_23980,N_22833);
nand UO_565 (O_565,N_24272,N_24585);
and UO_566 (O_566,N_24660,N_23906);
xor UO_567 (O_567,N_23695,N_22893);
xnor UO_568 (O_568,N_24055,N_23495);
xor UO_569 (O_569,N_24434,N_24687);
nand UO_570 (O_570,N_23349,N_24313);
and UO_571 (O_571,N_24163,N_23332);
xor UO_572 (O_572,N_24107,N_24776);
and UO_573 (O_573,N_24101,N_23624);
and UO_574 (O_574,N_23603,N_23711);
and UO_575 (O_575,N_22528,N_23451);
xor UO_576 (O_576,N_24008,N_23410);
and UO_577 (O_577,N_23378,N_24551);
nor UO_578 (O_578,N_23701,N_23639);
nand UO_579 (O_579,N_22841,N_22688);
xnor UO_580 (O_580,N_24908,N_23074);
xnor UO_581 (O_581,N_22755,N_23793);
nor UO_582 (O_582,N_24383,N_24370);
xor UO_583 (O_583,N_23325,N_23073);
xnor UO_584 (O_584,N_23521,N_23039);
nor UO_585 (O_585,N_23225,N_22604);
nand UO_586 (O_586,N_24820,N_23034);
xnor UO_587 (O_587,N_22781,N_24600);
nor UO_588 (O_588,N_24061,N_24295);
nor UO_589 (O_589,N_24194,N_24747);
nand UO_590 (O_590,N_23166,N_23285);
nor UO_591 (O_591,N_23131,N_22921);
nor UO_592 (O_592,N_24084,N_23835);
nand UO_593 (O_593,N_24563,N_24605);
xor UO_594 (O_594,N_24058,N_24420);
nor UO_595 (O_595,N_22501,N_24103);
or UO_596 (O_596,N_24656,N_23082);
nand UO_597 (O_597,N_23656,N_24791);
and UO_598 (O_598,N_22547,N_24457);
or UO_599 (O_599,N_23930,N_23807);
nor UO_600 (O_600,N_23121,N_23104);
or UO_601 (O_601,N_24275,N_24786);
or UO_602 (O_602,N_23958,N_23914);
or UO_603 (O_603,N_23146,N_24970);
and UO_604 (O_604,N_22700,N_23904);
or UO_605 (O_605,N_23777,N_23390);
and UO_606 (O_606,N_23035,N_23373);
xnor UO_607 (O_607,N_24177,N_23347);
nand UO_608 (O_608,N_23345,N_22786);
or UO_609 (O_609,N_24083,N_23880);
or UO_610 (O_610,N_24890,N_22651);
nor UO_611 (O_611,N_22875,N_24499);
and UO_612 (O_612,N_24745,N_23596);
nand UO_613 (O_613,N_23872,N_23101);
nand UO_614 (O_614,N_24005,N_23370);
or UO_615 (O_615,N_24288,N_23005);
nand UO_616 (O_616,N_23616,N_23222);
nand UO_617 (O_617,N_24131,N_22639);
xor UO_618 (O_618,N_23972,N_24912);
nor UO_619 (O_619,N_24657,N_23042);
nand UO_620 (O_620,N_23392,N_22573);
xor UO_621 (O_621,N_24393,N_23978);
and UO_622 (O_622,N_23963,N_22650);
and UO_623 (O_623,N_23700,N_24195);
nor UO_624 (O_624,N_22970,N_23106);
xnor UO_625 (O_625,N_22861,N_24257);
nand UO_626 (O_626,N_23622,N_23902);
or UO_627 (O_627,N_23552,N_23058);
nand UO_628 (O_628,N_23110,N_23446);
nand UO_629 (O_629,N_24097,N_24748);
and UO_630 (O_630,N_23709,N_24445);
nand UO_631 (O_631,N_23982,N_23821);
nand UO_632 (O_632,N_22556,N_23669);
xnor UO_633 (O_633,N_22504,N_23053);
xnor UO_634 (O_634,N_24573,N_22994);
or UO_635 (O_635,N_24836,N_22686);
and UO_636 (O_636,N_22739,N_23288);
xor UO_637 (O_637,N_24344,N_24678);
xnor UO_638 (O_638,N_23155,N_24610);
nand UO_639 (O_639,N_23509,N_24188);
nand UO_640 (O_640,N_24273,N_22912);
nor UO_641 (O_641,N_23524,N_22969);
nand UO_642 (O_642,N_24506,N_22932);
and UO_643 (O_643,N_22820,N_23098);
nor UO_644 (O_644,N_24428,N_24716);
xnor UO_645 (O_645,N_24792,N_22866);
xnor UO_646 (O_646,N_23570,N_23079);
nand UO_647 (O_647,N_23704,N_24104);
xnor UO_648 (O_648,N_24038,N_23422);
or UO_649 (O_649,N_22907,N_24827);
xor UO_650 (O_650,N_24355,N_23522);
xor UO_651 (O_651,N_22635,N_23786);
nand UO_652 (O_652,N_24220,N_22738);
and UO_653 (O_653,N_22643,N_22659);
xor UO_654 (O_654,N_22903,N_23617);
nor UO_655 (O_655,N_23343,N_24670);
nor UO_656 (O_656,N_22724,N_22742);
nand UO_657 (O_657,N_24033,N_24866);
or UO_658 (O_658,N_23530,N_24056);
nand UO_659 (O_659,N_24322,N_23748);
nand UO_660 (O_660,N_23721,N_22515);
nor UO_661 (O_661,N_23956,N_24959);
and UO_662 (O_662,N_23257,N_22719);
or UO_663 (O_663,N_24561,N_22945);
nor UO_664 (O_664,N_24592,N_24400);
or UO_665 (O_665,N_24070,N_24943);
or UO_666 (O_666,N_24105,N_24574);
or UO_667 (O_667,N_23132,N_23337);
and UO_668 (O_668,N_23028,N_22566);
or UO_669 (O_669,N_24153,N_23426);
nor UO_670 (O_670,N_24372,N_22731);
nand UO_671 (O_671,N_23710,N_22672);
nor UO_672 (O_672,N_24377,N_22674);
or UO_673 (O_673,N_24887,N_23460);
nor UO_674 (O_674,N_24854,N_22894);
xnor UO_675 (O_675,N_24192,N_23322);
and UO_676 (O_676,N_24213,N_22801);
xor UO_677 (O_677,N_24206,N_23056);
or UO_678 (O_678,N_23979,N_23575);
or UO_679 (O_679,N_24306,N_22904);
nand UO_680 (O_680,N_23323,N_23869);
nand UO_681 (O_681,N_23652,N_24897);
nand UO_682 (O_682,N_24997,N_23976);
xnor UO_683 (O_683,N_24914,N_23646);
nor UO_684 (O_684,N_23965,N_24556);
nor UO_685 (O_685,N_22965,N_24721);
xor UO_686 (O_686,N_24548,N_24018);
and UO_687 (O_687,N_23336,N_24078);
nand UO_688 (O_688,N_23678,N_24087);
xnor UO_689 (O_689,N_24366,N_22684);
or UO_690 (O_690,N_24472,N_22569);
and UO_691 (O_691,N_23752,N_24926);
or UO_692 (O_692,N_24814,N_23569);
or UO_693 (O_693,N_22579,N_23586);
or UO_694 (O_694,N_22749,N_24279);
or UO_695 (O_695,N_23180,N_24387);
and UO_696 (O_696,N_22677,N_22757);
and UO_697 (O_697,N_24109,N_22900);
nor UO_698 (O_698,N_23004,N_23740);
xor UO_699 (O_699,N_24602,N_24096);
or UO_700 (O_700,N_22575,N_24198);
or UO_701 (O_701,N_23734,N_24945);
and UO_702 (O_702,N_24614,N_23871);
nand UO_703 (O_703,N_23385,N_23116);
and UO_704 (O_704,N_24016,N_23822);
nor UO_705 (O_705,N_23237,N_22648);
or UO_706 (O_706,N_23741,N_23263);
and UO_707 (O_707,N_23966,N_24838);
nor UO_708 (O_708,N_24584,N_23040);
xnor UO_709 (O_709,N_24956,N_23017);
nand UO_710 (O_710,N_22624,N_22829);
or UO_711 (O_711,N_24983,N_23149);
or UO_712 (O_712,N_24046,N_24761);
and UO_713 (O_713,N_24471,N_23232);
nor UO_714 (O_714,N_23022,N_24332);
nand UO_715 (O_715,N_24510,N_24699);
and UO_716 (O_716,N_24057,N_24850);
nor UO_717 (O_717,N_23113,N_24157);
or UO_718 (O_718,N_22574,N_23894);
nand UO_719 (O_719,N_24537,N_24182);
nor UO_720 (O_720,N_23830,N_22502);
or UO_721 (O_721,N_24276,N_24993);
and UO_722 (O_722,N_23896,N_22661);
or UO_723 (O_723,N_23122,N_23086);
nand UO_724 (O_724,N_23199,N_22805);
xnor UO_725 (O_725,N_24542,N_24857);
nor UO_726 (O_726,N_24906,N_24704);
xnor UO_727 (O_727,N_24726,N_24336);
or UO_728 (O_728,N_23281,N_23749);
nor UO_729 (O_729,N_24496,N_22822);
nor UO_730 (O_730,N_24054,N_23313);
xnor UO_731 (O_731,N_24128,N_23255);
nor UO_732 (O_732,N_22592,N_24044);
and UO_733 (O_733,N_22795,N_23312);
nand UO_734 (O_734,N_24690,N_24001);
and UO_735 (O_735,N_24910,N_24532);
nand UO_736 (O_736,N_23463,N_24482);
xor UO_737 (O_737,N_22993,N_24121);
and UO_738 (O_738,N_24430,N_24454);
nor UO_739 (O_739,N_23756,N_23546);
nand UO_740 (O_740,N_23050,N_24833);
nor UO_741 (O_741,N_24264,N_24358);
or UO_742 (O_742,N_24235,N_23923);
and UO_743 (O_743,N_22953,N_23697);
or UO_744 (O_744,N_23601,N_23503);
xnor UO_745 (O_745,N_24710,N_23508);
xnor UO_746 (O_746,N_22884,N_24470);
and UO_747 (O_747,N_24117,N_24995);
or UO_748 (O_748,N_22913,N_24884);
xor UO_749 (O_749,N_23761,N_24953);
nor UO_750 (O_750,N_23834,N_24174);
nor UO_751 (O_751,N_23772,N_22794);
xor UO_752 (O_752,N_22500,N_24092);
nor UO_753 (O_753,N_23809,N_24065);
and UO_754 (O_754,N_23895,N_24567);
and UO_755 (O_755,N_23501,N_24354);
and UO_756 (O_756,N_24500,N_23927);
xnor UO_757 (O_757,N_23931,N_23226);
nand UO_758 (O_758,N_22872,N_23268);
nand UO_759 (O_759,N_24907,N_23037);
and UO_760 (O_760,N_24810,N_24359);
nor UO_761 (O_761,N_24543,N_23284);
or UO_762 (O_762,N_23466,N_23427);
nand UO_763 (O_763,N_24625,N_24972);
nor UO_764 (O_764,N_22879,N_23087);
or UO_765 (O_765,N_23957,N_22614);
or UO_766 (O_766,N_24628,N_24115);
nand UO_767 (O_767,N_22707,N_24694);
nand UO_768 (O_768,N_23000,N_22885);
nand UO_769 (O_769,N_22832,N_23383);
or UO_770 (O_770,N_22901,N_22981);
nor UO_771 (O_771,N_24896,N_22859);
nand UO_772 (O_772,N_24793,N_24328);
xnor UO_773 (O_773,N_24397,N_23380);
or UO_774 (O_774,N_24438,N_22863);
xor UO_775 (O_775,N_24465,N_24380);
nor UO_776 (O_776,N_24684,N_23434);
nor UO_777 (O_777,N_23641,N_23726);
nor UO_778 (O_778,N_23407,N_23990);
and UO_779 (O_779,N_22878,N_22714);
nor UO_780 (O_780,N_24314,N_23610);
nor UO_781 (O_781,N_23482,N_23729);
nand UO_782 (O_782,N_24925,N_24187);
xnor UO_783 (O_783,N_23959,N_22527);
and UO_784 (O_784,N_24942,N_23216);
xnor UO_785 (O_785,N_23310,N_23038);
or UO_786 (O_786,N_24069,N_22942);
nor UO_787 (O_787,N_24325,N_23264);
and UO_788 (O_788,N_23806,N_24822);
and UO_789 (O_789,N_23423,N_24911);
and UO_790 (O_790,N_22565,N_23273);
or UO_791 (O_791,N_22784,N_24560);
and UO_792 (O_792,N_22873,N_24750);
nand UO_793 (O_793,N_24252,N_23795);
nand UO_794 (O_794,N_24027,N_24154);
xor UO_795 (O_795,N_24184,N_24216);
nand UO_796 (O_796,N_24186,N_24780);
nand UO_797 (O_797,N_24528,N_24613);
nor UO_798 (O_798,N_22654,N_24373);
or UO_799 (O_799,N_23357,N_22868);
nor UO_800 (O_800,N_23269,N_22778);
nand UO_801 (O_801,N_24053,N_22554);
xor UO_802 (O_802,N_23449,N_23949);
nor UO_803 (O_803,N_23002,N_23961);
xor UO_804 (O_804,N_22967,N_22692);
nor UO_805 (O_805,N_23595,N_23382);
nand UO_806 (O_806,N_24265,N_23452);
and UO_807 (O_807,N_22888,N_24847);
xor UO_808 (O_808,N_23502,N_24374);
or UO_809 (O_809,N_23558,N_23750);
nor UO_810 (O_810,N_23488,N_24856);
xor UO_811 (O_811,N_23368,N_23565);
nand UO_812 (O_812,N_24654,N_23408);
or UO_813 (O_813,N_22792,N_23008);
nand UO_814 (O_814,N_23985,N_23388);
nand UO_815 (O_815,N_24785,N_24253);
nand UO_816 (O_816,N_24879,N_23506);
and UO_817 (O_817,N_22949,N_24954);
and UO_818 (O_818,N_24317,N_23191);
and UO_819 (O_819,N_22905,N_23197);
and UO_820 (O_820,N_24861,N_23812);
nand UO_821 (O_821,N_24301,N_23075);
or UO_822 (O_822,N_24164,N_23401);
xor UO_823 (O_823,N_23085,N_24243);
nand UO_824 (O_824,N_22818,N_24867);
nand UO_825 (O_825,N_24759,N_24502);
nor UO_826 (O_826,N_24824,N_23393);
nor UO_827 (O_827,N_24015,N_24948);
nand UO_828 (O_828,N_24988,N_24891);
nor UO_829 (O_829,N_24223,N_22934);
and UO_830 (O_830,N_24775,N_23778);
and UO_831 (O_831,N_23456,N_23230);
and UO_832 (O_832,N_24781,N_23201);
or UO_833 (O_833,N_23787,N_23399);
xnor UO_834 (O_834,N_24486,N_22622);
nand UO_835 (O_835,N_22706,N_23527);
xnor UO_836 (O_836,N_23013,N_23685);
and UO_837 (O_837,N_24166,N_24651);
nor UO_838 (O_838,N_24479,N_23290);
nor UO_839 (O_839,N_24662,N_23626);
nand UO_840 (O_840,N_23714,N_23905);
nor UO_841 (O_841,N_23707,N_24368);
and UO_842 (O_842,N_23716,N_22860);
xor UO_843 (O_843,N_24698,N_24073);
xnor UO_844 (O_844,N_22766,N_24835);
xor UO_845 (O_845,N_23816,N_23539);
or UO_846 (O_846,N_24508,N_24794);
nand UO_847 (O_847,N_24834,N_24934);
xor UO_848 (O_848,N_23174,N_22777);
and UO_849 (O_849,N_24017,N_22865);
and UO_850 (O_850,N_24570,N_24531);
or UO_851 (O_851,N_23505,N_23719);
xnor UO_852 (O_852,N_22652,N_22916);
or UO_853 (O_853,N_22748,N_24406);
nand UO_854 (O_854,N_24419,N_23684);
xnor UO_855 (O_855,N_23108,N_22896);
nand UO_856 (O_856,N_24080,N_24051);
xnor UO_857 (O_857,N_22754,N_23535);
nor UO_858 (O_858,N_24787,N_24920);
and UO_859 (O_859,N_24143,N_22668);
nand UO_860 (O_860,N_23960,N_23297);
and UO_861 (O_861,N_24979,N_23846);
nand UO_862 (O_862,N_23636,N_24568);
and UO_863 (O_863,N_24079,N_23318);
nor UO_864 (O_864,N_23119,N_23754);
or UO_865 (O_865,N_23954,N_24876);
nand UO_866 (O_866,N_23736,N_23964);
nand UO_867 (O_867,N_24338,N_24309);
or UO_868 (O_868,N_23469,N_24039);
nor UO_869 (O_869,N_22509,N_24477);
and UO_870 (O_870,N_24905,N_24848);
xnor UO_871 (O_871,N_22804,N_24971);
nor UO_872 (O_872,N_23346,N_22525);
or UO_873 (O_873,N_24071,N_23995);
nor UO_874 (O_874,N_24049,N_24525);
xor UO_875 (O_875,N_24132,N_22991);
xnor UO_876 (O_876,N_24562,N_24852);
or UO_877 (O_877,N_24519,N_22627);
xnor UO_878 (O_878,N_24588,N_24036);
nand UO_879 (O_879,N_22553,N_22533);
nor UO_880 (O_880,N_22638,N_23955);
nand UO_881 (O_881,N_23198,N_24774);
or UO_882 (O_882,N_23744,N_22989);
nand UO_883 (O_883,N_24148,N_23443);
or UO_884 (O_884,N_22824,N_23549);
and UO_885 (O_885,N_24982,N_23559);
nor UO_886 (O_886,N_23066,N_22678);
xor UO_887 (O_887,N_24196,N_24043);
nor UO_888 (O_888,N_23920,N_23989);
xnor UO_889 (O_889,N_23832,N_22939);
nand UO_890 (O_890,N_23305,N_24633);
nand UO_891 (O_891,N_22842,N_24767);
nand UO_892 (O_892,N_24236,N_24675);
xor UO_893 (O_893,N_23929,N_23100);
nor UO_894 (O_894,N_23173,N_24783);
and UO_895 (O_895,N_23298,N_23849);
nor UO_896 (O_896,N_23351,N_24715);
nor UO_897 (O_897,N_23142,N_22790);
nor UO_898 (O_898,N_23445,N_24855);
nand UO_899 (O_899,N_24973,N_24237);
xnor UO_900 (O_900,N_22621,N_23827);
xnor UO_901 (O_901,N_24189,N_23060);
nor UO_902 (O_902,N_24859,N_24175);
or UO_903 (O_903,N_23244,N_23289);
nand UO_904 (O_904,N_23207,N_23417);
or UO_905 (O_905,N_24801,N_24811);
and UO_906 (O_906,N_23157,N_23262);
and UO_907 (O_907,N_24111,N_22733);
xnor UO_908 (O_908,N_24558,N_23243);
nand UO_909 (O_909,N_24140,N_23511);
nor UO_910 (O_910,N_24550,N_24623);
xnor UO_911 (O_911,N_24649,N_24040);
and UO_912 (O_912,N_23212,N_24638);
nor UO_913 (O_913,N_24849,N_22728);
xor UO_914 (O_914,N_23492,N_23882);
and UO_915 (O_915,N_22761,N_24130);
or UO_916 (O_916,N_23200,N_22788);
and UO_917 (O_917,N_22800,N_22834);
nor UO_918 (O_918,N_22718,N_24930);
or UO_919 (O_919,N_24346,N_22810);
nor UO_920 (O_920,N_24045,N_24207);
nand UO_921 (O_921,N_23018,N_23554);
or UO_922 (O_922,N_24960,N_22524);
nor UO_923 (O_923,N_23842,N_23732);
xor UO_924 (O_924,N_23352,N_22920);
and UO_925 (O_925,N_24509,N_23883);
nor UO_926 (O_926,N_23766,N_23484);
nor UO_927 (O_927,N_22762,N_24809);
and UO_928 (O_928,N_22695,N_23910);
xor UO_929 (O_929,N_24727,N_22806);
or UO_930 (O_930,N_23942,N_24396);
or UO_931 (O_931,N_22765,N_24241);
xor UO_932 (O_932,N_23924,N_24564);
nor UO_933 (O_933,N_22631,N_24611);
xnor UO_934 (O_934,N_22943,N_24741);
nand UO_935 (O_935,N_23544,N_23365);
nor UO_936 (O_936,N_23588,N_23103);
nand UO_937 (O_937,N_24595,N_24371);
nor UO_938 (O_938,N_23655,N_24941);
or UO_939 (O_939,N_24842,N_22891);
or UO_940 (O_940,N_23384,N_23433);
xnor UO_941 (O_941,N_24009,N_24609);
xnor UO_942 (O_942,N_24032,N_22756);
nor UO_943 (O_943,N_22549,N_24034);
and UO_944 (O_944,N_24432,N_24048);
xnor UO_945 (O_945,N_23301,N_23396);
or UO_946 (O_946,N_24389,N_24647);
and UO_947 (O_947,N_24437,N_23145);
nand UO_948 (O_948,N_24365,N_23657);
xor UO_949 (O_949,N_22825,N_24224);
nand UO_950 (O_950,N_22555,N_23643);
and UO_951 (O_951,N_22782,N_24088);
and UO_952 (O_952,N_23580,N_22852);
and UO_953 (O_953,N_23168,N_22511);
nand UO_954 (O_954,N_24072,N_23183);
xnor UO_955 (O_955,N_24524,N_24494);
or UO_956 (O_956,N_22803,N_24841);
xor UO_957 (O_957,N_24768,N_23409);
or UO_958 (O_958,N_24766,N_23718);
nand UO_959 (O_959,N_22517,N_24596);
nor UO_960 (O_960,N_23046,N_23607);
or UO_961 (O_961,N_23210,N_24858);
nand UO_962 (O_962,N_22611,N_23780);
xor UO_963 (O_963,N_22960,N_22973);
nor UO_964 (O_964,N_24311,N_24004);
nand UO_965 (O_965,N_23275,N_24697);
nor UO_966 (O_966,N_24474,N_23791);
nand UO_967 (O_967,N_22703,N_23030);
xor UO_968 (O_968,N_22968,N_24095);
xor UO_969 (O_969,N_22821,N_24736);
nor UO_970 (O_970,N_22998,N_24090);
or UO_971 (O_971,N_23178,N_23940);
or UO_972 (O_972,N_23364,N_24155);
nand UO_973 (O_973,N_23374,N_23454);
xnor UO_974 (O_974,N_23339,N_23808);
nand UO_975 (O_975,N_24002,N_24617);
and UO_976 (O_976,N_23706,N_23582);
and UO_977 (O_977,N_24555,N_23317);
or UO_978 (O_978,N_23932,N_23928);
xor UO_979 (O_979,N_24580,N_23922);
xnor UO_980 (O_980,N_23913,N_23850);
nor UO_981 (O_981,N_23675,N_22671);
nand UO_982 (O_982,N_24688,N_23654);
and UO_983 (O_983,N_24417,N_22946);
nand UO_984 (O_984,N_22508,N_22626);
xnor UO_985 (O_985,N_22976,N_24388);
nand UO_986 (O_986,N_23689,N_23911);
nand UO_987 (O_987,N_22545,N_24025);
and UO_988 (O_988,N_22699,N_23540);
or UO_989 (O_989,N_23397,N_24760);
nor UO_990 (O_990,N_22552,N_23801);
xnor UO_991 (O_991,N_24347,N_24407);
nand UO_992 (O_992,N_24882,N_22734);
and UO_993 (O_993,N_24404,N_24172);
nor UO_994 (O_994,N_24291,N_22987);
nor UO_995 (O_995,N_23236,N_23480);
nor UO_996 (O_996,N_23640,N_22926);
and UO_997 (O_997,N_24764,N_23088);
nor UO_998 (O_998,N_23246,N_23874);
or UO_999 (O_999,N_23470,N_23865);
xnor UO_1000 (O_1000,N_24735,N_23286);
nand UO_1001 (O_1001,N_22507,N_24451);
nor UO_1002 (O_1002,N_24674,N_24873);
and UO_1003 (O_1003,N_23757,N_23324);
nand UO_1004 (O_1004,N_23092,N_22505);
nand UO_1005 (O_1005,N_24076,N_23708);
and UO_1006 (O_1006,N_24523,N_24935);
xnor UO_1007 (O_1007,N_24068,N_23802);
and UO_1008 (O_1008,N_23179,N_24197);
and UO_1009 (O_1009,N_24066,N_24226);
xnor UO_1010 (O_1010,N_22740,N_23418);
nor UO_1011 (O_1011,N_22690,N_23900);
nand UO_1012 (O_1012,N_24335,N_22520);
xor UO_1013 (O_1013,N_23843,N_23781);
and UO_1014 (O_1014,N_23623,N_24327);
or UO_1015 (O_1015,N_23436,N_23547);
or UO_1016 (O_1016,N_24957,N_23442);
nor UO_1017 (O_1017,N_23340,N_23350);
and UO_1018 (O_1018,N_24985,N_23986);
and UO_1019 (O_1019,N_24664,N_22958);
or UO_1020 (O_1020,N_24021,N_23703);
and UO_1021 (O_1021,N_22886,N_24769);
xor UO_1022 (O_1022,N_23306,N_23209);
or UO_1023 (O_1023,N_23478,N_24851);
nor UO_1024 (O_1024,N_24421,N_22951);
nand UO_1025 (O_1025,N_24391,N_22526);
and UO_1026 (O_1026,N_23873,N_23015);
or UO_1027 (O_1027,N_23202,N_24818);
or UO_1028 (O_1028,N_23238,N_24922);
nor UO_1029 (O_1029,N_24789,N_22521);
and UO_1030 (O_1030,N_22914,N_22632);
and UO_1031 (O_1031,N_24190,N_23693);
or UO_1032 (O_1032,N_23276,N_24597);
and UO_1033 (O_1033,N_24150,N_23829);
nand UO_1034 (O_1034,N_23147,N_22922);
or UO_1035 (O_1035,N_24411,N_24114);
nand UO_1036 (O_1036,N_24149,N_23720);
or UO_1037 (O_1037,N_22664,N_23938);
nor UO_1038 (O_1038,N_23934,N_24517);
xor UO_1039 (O_1039,N_24491,N_22610);
nand UO_1040 (O_1040,N_23759,N_23462);
nor UO_1041 (O_1041,N_22694,N_24655);
or UO_1042 (O_1042,N_24165,N_23021);
nand UO_1043 (O_1043,N_23153,N_22940);
xor UO_1044 (O_1044,N_23398,N_24378);
nor UO_1045 (O_1045,N_24204,N_23642);
xor UO_1046 (O_1046,N_24763,N_24892);
nor UO_1047 (O_1047,N_23686,N_23097);
nor UO_1048 (O_1048,N_23836,N_24642);
nand UO_1049 (O_1049,N_23974,N_22854);
and UO_1050 (O_1050,N_23084,N_23514);
xor UO_1051 (O_1051,N_23672,N_24513);
and UO_1052 (O_1052,N_23860,N_23775);
and UO_1053 (O_1053,N_24062,N_23948);
xnor UO_1054 (O_1054,N_22753,N_22827);
nand UO_1055 (O_1055,N_24720,N_22763);
xnor UO_1056 (O_1056,N_23414,N_23065);
nor UO_1057 (O_1057,N_23645,N_23602);
and UO_1058 (O_1058,N_24974,N_24085);
nor UO_1059 (O_1059,N_22846,N_24778);
nand UO_1060 (O_1060,N_24127,N_22902);
and UO_1061 (O_1061,N_24089,N_22797);
nor UO_1062 (O_1062,N_23839,N_24724);
and UO_1063 (O_1063,N_24159,N_24547);
nand UO_1064 (O_1064,N_23486,N_22587);
nand UO_1065 (O_1065,N_24191,N_23453);
and UO_1066 (O_1066,N_22557,N_24501);
nor UO_1067 (O_1067,N_24996,N_22608);
nand UO_1068 (O_1068,N_23429,N_22809);
or UO_1069 (O_1069,N_24512,N_24893);
nor UO_1070 (O_1070,N_24334,N_24622);
and UO_1071 (O_1071,N_22737,N_22980);
or UO_1072 (O_1072,N_23862,N_23629);
xnor UO_1073 (O_1073,N_24616,N_22845);
nor UO_1074 (O_1074,N_22702,N_22689);
nor UO_1075 (O_1075,N_23059,N_24050);
xor UO_1076 (O_1076,N_22577,N_23240);
or UO_1077 (O_1077,N_22510,N_23881);
or UO_1078 (O_1078,N_22807,N_22864);
and UO_1079 (O_1079,N_23676,N_22657);
nor UO_1080 (O_1080,N_22955,N_23992);
or UO_1081 (O_1081,N_24297,N_22735);
nand UO_1082 (O_1082,N_24466,N_24116);
nor UO_1083 (O_1083,N_24000,N_24784);
and UO_1084 (O_1084,N_23249,N_24961);
or UO_1085 (O_1085,N_24807,N_23796);
nor UO_1086 (O_1086,N_22658,N_22876);
nor UO_1087 (O_1087,N_23887,N_23571);
and UO_1088 (O_1088,N_23561,N_23229);
nor UO_1089 (O_1089,N_24446,N_23144);
nor UO_1090 (O_1090,N_23099,N_24952);
nor UO_1091 (O_1091,N_23083,N_22578);
nor UO_1092 (O_1092,N_24705,N_24081);
or UO_1093 (O_1093,N_24737,N_24003);
and UO_1094 (O_1094,N_24441,N_23457);
or UO_1095 (O_1095,N_24799,N_24659);
or UO_1096 (O_1096,N_24546,N_23677);
nand UO_1097 (O_1097,N_23727,N_23387);
and UO_1098 (O_1098,N_23464,N_24545);
and UO_1099 (O_1099,N_24539,N_23128);
nor UO_1100 (O_1100,N_23782,N_22640);
nor UO_1101 (O_1101,N_23673,N_23130);
xnor UO_1102 (O_1102,N_24183,N_23428);
and UO_1103 (O_1103,N_23557,N_23717);
nor UO_1104 (O_1104,N_22710,N_24376);
or UO_1105 (O_1105,N_22514,N_24899);
nor UO_1106 (O_1106,N_24138,N_23975);
xor UO_1107 (O_1107,N_23252,N_24917);
xnor UO_1108 (O_1108,N_23765,N_22623);
xor UO_1109 (O_1109,N_23068,N_23355);
and UO_1110 (O_1110,N_23129,N_23593);
and UO_1111 (O_1111,N_23858,N_22988);
nor UO_1112 (O_1112,N_23300,N_24577);
nand UO_1113 (O_1113,N_24618,N_24816);
nand UO_1114 (O_1114,N_23528,N_23971);
xor UO_1115 (O_1115,N_24673,N_23481);
and UO_1116 (O_1116,N_23769,N_24644);
nand UO_1117 (O_1117,N_24193,N_24732);
nor UO_1118 (O_1118,N_24110,N_23770);
or UO_1119 (O_1119,N_23556,N_24020);
nand UO_1120 (O_1120,N_23280,N_23831);
nor UO_1121 (O_1121,N_24958,N_23448);
and UO_1122 (O_1122,N_23327,N_22609);
nand UO_1123 (O_1123,N_24931,N_23592);
xor UO_1124 (O_1124,N_22917,N_22855);
or UO_1125 (O_1125,N_23291,N_24619);
xor UO_1126 (O_1126,N_24886,N_22743);
xor UO_1127 (O_1127,N_24860,N_23632);
or UO_1128 (O_1128,N_23006,N_24806);
or UO_1129 (O_1129,N_23447,N_24488);
or UO_1130 (O_1130,N_24615,N_23604);
xnor UO_1131 (O_1131,N_24485,N_24321);
and UO_1132 (O_1132,N_22529,N_23788);
and UO_1133 (O_1133,N_23585,N_24669);
and UO_1134 (O_1134,N_22948,N_23043);
xor UO_1135 (O_1135,N_23510,N_24977);
nor UO_1136 (O_1136,N_24691,N_23233);
nand UO_1137 (O_1137,N_23776,N_23953);
xnor UO_1138 (O_1138,N_23745,N_24093);
or UO_1139 (O_1139,N_22625,N_22617);
and UO_1140 (O_1140,N_23526,N_22783);
and UO_1141 (O_1141,N_24955,N_22634);
and UO_1142 (O_1142,N_23319,N_23536);
or UO_1143 (O_1143,N_24805,N_23023);
xnor UO_1144 (O_1144,N_22745,N_24229);
nor UO_1145 (O_1145,N_24650,N_24752);
nor UO_1146 (O_1146,N_24639,N_24442);
and UO_1147 (O_1147,N_24151,N_24804);
nand UO_1148 (O_1148,N_23283,N_24635);
xnor UO_1149 (O_1149,N_24227,N_23828);
nand UO_1150 (O_1150,N_23371,N_22603);
and UO_1151 (O_1151,N_24262,N_23926);
nand UO_1152 (O_1152,N_23304,N_22667);
nand UO_1153 (O_1153,N_24360,N_22816);
nor UO_1154 (O_1154,N_23628,N_23968);
nand UO_1155 (O_1155,N_24904,N_24624);
xor UO_1156 (O_1156,N_23599,N_23739);
nand UO_1157 (O_1157,N_24762,N_22974);
nand UO_1158 (O_1158,N_23001,N_24530);
and UO_1159 (O_1159,N_23055,N_24819);
xnor UO_1160 (O_1160,N_23499,N_24280);
nand UO_1161 (O_1161,N_23361,N_24123);
and UO_1162 (O_1162,N_22576,N_23061);
or UO_1163 (O_1163,N_22898,N_22683);
nand UO_1164 (O_1164,N_23192,N_24287);
or UO_1165 (O_1165,N_24790,N_22856);
nand UO_1166 (O_1166,N_23578,N_22572);
and UO_1167 (O_1167,N_24357,N_24459);
nand UO_1168 (O_1168,N_23331,N_23497);
and UO_1169 (O_1169,N_22567,N_23794);
xor UO_1170 (O_1170,N_23048,N_23783);
and UO_1171 (O_1171,N_23591,N_22767);
nor UO_1172 (O_1172,N_23841,N_23014);
and UO_1173 (O_1173,N_24593,N_24829);
and UO_1174 (O_1174,N_23901,N_22598);
nand UO_1175 (O_1175,N_23994,N_24415);
xnor UO_1176 (O_1176,N_23751,N_24696);
and UO_1177 (O_1177,N_22817,N_22814);
or UO_1178 (O_1178,N_24394,N_23983);
nand UO_1179 (O_1179,N_23458,N_22982);
nor UO_1180 (O_1180,N_22911,N_23114);
nor UO_1181 (O_1181,N_22523,N_24950);
or UO_1182 (O_1182,N_23952,N_23833);
nor UO_1183 (O_1183,N_22544,N_22568);
nor UO_1184 (O_1184,N_22906,N_22662);
nor UO_1185 (O_1185,N_24364,N_24504);
nor UO_1186 (O_1186,N_23589,N_24141);
nand UO_1187 (O_1187,N_23386,N_24589);
nand UO_1188 (O_1188,N_23164,N_23919);
xnor UO_1189 (O_1189,N_24634,N_23335);
or UO_1190 (O_1190,N_24250,N_24312);
or UO_1191 (O_1191,N_23962,N_24343);
and UO_1192 (O_1192,N_24777,N_23329);
or UO_1193 (O_1193,N_23944,N_23705);
nor UO_1194 (O_1194,N_22538,N_22759);
xnor UO_1195 (O_1195,N_23688,N_24221);
or UO_1196 (O_1196,N_22828,N_23169);
xnor UO_1197 (O_1197,N_24231,N_23538);
and UO_1198 (O_1198,N_23402,N_24756);
and UO_1199 (O_1199,N_23814,N_24582);
or UO_1200 (O_1200,N_23026,N_23915);
and UO_1201 (O_1201,N_23158,N_22596);
nand UO_1202 (O_1202,N_23999,N_23533);
nand UO_1203 (O_1203,N_23138,N_23421);
xnor UO_1204 (O_1204,N_23746,N_23251);
or UO_1205 (O_1205,N_22682,N_24963);
nand UO_1206 (O_1206,N_24575,N_23545);
xor UO_1207 (O_1207,N_23476,N_24443);
or UO_1208 (O_1208,N_22513,N_24399);
and UO_1209 (O_1209,N_24382,N_24962);
and UO_1210 (O_1210,N_23790,N_24652);
xor UO_1211 (O_1211,N_24772,N_23851);
or UO_1212 (O_1212,N_23430,N_23095);
or UO_1213 (O_1213,N_23052,N_23647);
or UO_1214 (O_1214,N_22950,N_24211);
nand UO_1215 (O_1215,N_24412,N_23117);
and UO_1216 (O_1216,N_22698,N_22535);
nand UO_1217 (O_1217,N_24251,N_23738);
xor UO_1218 (O_1218,N_24167,N_24267);
and UO_1219 (O_1219,N_23532,N_23217);
xnor UO_1220 (O_1220,N_24489,N_24514);
or UO_1221 (O_1221,N_24901,N_24682);
and UO_1222 (O_1222,N_22889,N_24082);
xnor UO_1223 (O_1223,N_24238,N_23635);
or UO_1224 (O_1224,N_23577,N_23069);
xor UO_1225 (O_1225,N_22954,N_23627);
nand UO_1226 (O_1226,N_22819,N_23221);
nor UO_1227 (O_1227,N_24540,N_23044);
nor UO_1228 (O_1228,N_23356,N_23112);
and UO_1229 (O_1229,N_23267,N_24511);
and UO_1230 (O_1230,N_22522,N_23011);
and UO_1231 (O_1231,N_24522,N_24064);
nand UO_1232 (O_1232,N_23171,N_24319);
nor UO_1233 (O_1233,N_22704,N_22996);
and UO_1234 (O_1234,N_22744,N_24591);
nand UO_1235 (O_1235,N_23344,N_24552);
nor UO_1236 (O_1236,N_22908,N_24939);
or UO_1237 (O_1237,N_22850,N_24830);
or UO_1238 (O_1238,N_24843,N_24469);
and UO_1239 (O_1239,N_23659,N_24516);
and UO_1240 (O_1240,N_24423,N_23223);
nor UO_1241 (O_1241,N_24458,N_24483);
nor UO_1242 (O_1242,N_22564,N_22774);
or UO_1243 (O_1243,N_23473,N_23819);
or UO_1244 (O_1244,N_22947,N_22601);
xnor UO_1245 (O_1245,N_24683,N_24863);
nor UO_1246 (O_1246,N_23513,N_24518);
and UO_1247 (O_1247,N_23431,N_24481);
xor UO_1248 (O_1248,N_23472,N_23621);
xnor UO_1249 (O_1249,N_24498,N_22897);
or UO_1250 (O_1250,N_23070,N_23856);
and UO_1251 (O_1251,N_24969,N_22895);
xor UO_1252 (O_1252,N_24200,N_24619);
nor UO_1253 (O_1253,N_24592,N_24940);
or UO_1254 (O_1254,N_23306,N_23927);
or UO_1255 (O_1255,N_23063,N_23087);
nand UO_1256 (O_1256,N_24172,N_23414);
nor UO_1257 (O_1257,N_23650,N_24318);
or UO_1258 (O_1258,N_23318,N_24585);
and UO_1259 (O_1259,N_23809,N_23645);
nor UO_1260 (O_1260,N_22547,N_24333);
and UO_1261 (O_1261,N_24854,N_24818);
nand UO_1262 (O_1262,N_23912,N_24483);
and UO_1263 (O_1263,N_22582,N_23541);
or UO_1264 (O_1264,N_23397,N_24125);
and UO_1265 (O_1265,N_23330,N_24039);
nand UO_1266 (O_1266,N_23358,N_23495);
or UO_1267 (O_1267,N_23329,N_24367);
nor UO_1268 (O_1268,N_22729,N_22532);
or UO_1269 (O_1269,N_23220,N_23368);
nor UO_1270 (O_1270,N_24544,N_24166);
nor UO_1271 (O_1271,N_22995,N_23550);
and UO_1272 (O_1272,N_23915,N_24623);
xor UO_1273 (O_1273,N_24384,N_24436);
nor UO_1274 (O_1274,N_23071,N_23178);
xnor UO_1275 (O_1275,N_22839,N_23612);
xnor UO_1276 (O_1276,N_24719,N_23412);
xnor UO_1277 (O_1277,N_22742,N_24058);
nor UO_1278 (O_1278,N_23639,N_23912);
nor UO_1279 (O_1279,N_23341,N_24395);
nand UO_1280 (O_1280,N_23546,N_22760);
or UO_1281 (O_1281,N_24977,N_24324);
nand UO_1282 (O_1282,N_24663,N_24348);
or UO_1283 (O_1283,N_22775,N_22778);
nor UO_1284 (O_1284,N_23981,N_24419);
nand UO_1285 (O_1285,N_24957,N_22591);
and UO_1286 (O_1286,N_24367,N_23384);
and UO_1287 (O_1287,N_24841,N_24778);
xnor UO_1288 (O_1288,N_24124,N_24617);
or UO_1289 (O_1289,N_23016,N_22990);
nor UO_1290 (O_1290,N_23395,N_23584);
and UO_1291 (O_1291,N_24962,N_24713);
and UO_1292 (O_1292,N_24738,N_23798);
and UO_1293 (O_1293,N_23776,N_23605);
nor UO_1294 (O_1294,N_23718,N_24242);
nand UO_1295 (O_1295,N_24267,N_24191);
or UO_1296 (O_1296,N_23417,N_23553);
nor UO_1297 (O_1297,N_23875,N_23186);
or UO_1298 (O_1298,N_23766,N_24683);
nand UO_1299 (O_1299,N_23987,N_23210);
xor UO_1300 (O_1300,N_23409,N_24904);
or UO_1301 (O_1301,N_23325,N_23204);
and UO_1302 (O_1302,N_24515,N_24709);
and UO_1303 (O_1303,N_23764,N_23887);
nand UO_1304 (O_1304,N_24953,N_23724);
xor UO_1305 (O_1305,N_24115,N_24071);
xor UO_1306 (O_1306,N_23470,N_24686);
xnor UO_1307 (O_1307,N_24228,N_24690);
nor UO_1308 (O_1308,N_22563,N_23605);
nand UO_1309 (O_1309,N_22717,N_24250);
or UO_1310 (O_1310,N_24001,N_24748);
or UO_1311 (O_1311,N_24560,N_23841);
and UO_1312 (O_1312,N_23931,N_23073);
nor UO_1313 (O_1313,N_23765,N_23669);
and UO_1314 (O_1314,N_23682,N_23396);
nand UO_1315 (O_1315,N_22887,N_24024);
nor UO_1316 (O_1316,N_24148,N_23050);
xor UO_1317 (O_1317,N_24352,N_23542);
or UO_1318 (O_1318,N_24080,N_24148);
nor UO_1319 (O_1319,N_22836,N_22634);
and UO_1320 (O_1320,N_22564,N_24986);
or UO_1321 (O_1321,N_22660,N_22869);
and UO_1322 (O_1322,N_23828,N_24538);
xor UO_1323 (O_1323,N_23616,N_24649);
nand UO_1324 (O_1324,N_23659,N_24020);
nand UO_1325 (O_1325,N_24364,N_24371);
or UO_1326 (O_1326,N_24002,N_23803);
or UO_1327 (O_1327,N_24061,N_23312);
nand UO_1328 (O_1328,N_23234,N_24518);
or UO_1329 (O_1329,N_22858,N_24565);
nand UO_1330 (O_1330,N_24472,N_22786);
xor UO_1331 (O_1331,N_24393,N_23242);
or UO_1332 (O_1332,N_22543,N_22758);
and UO_1333 (O_1333,N_24951,N_22919);
and UO_1334 (O_1334,N_24626,N_24268);
and UO_1335 (O_1335,N_22562,N_22994);
nor UO_1336 (O_1336,N_22607,N_22826);
or UO_1337 (O_1337,N_22697,N_24914);
and UO_1338 (O_1338,N_23376,N_22987);
or UO_1339 (O_1339,N_23048,N_22741);
nand UO_1340 (O_1340,N_24205,N_23295);
xor UO_1341 (O_1341,N_22977,N_22572);
or UO_1342 (O_1342,N_22503,N_23011);
or UO_1343 (O_1343,N_24646,N_24033);
nor UO_1344 (O_1344,N_22529,N_22507);
nor UO_1345 (O_1345,N_23719,N_24902);
nand UO_1346 (O_1346,N_23504,N_22541);
nand UO_1347 (O_1347,N_24594,N_24668);
xor UO_1348 (O_1348,N_22519,N_23350);
and UO_1349 (O_1349,N_24228,N_24392);
nand UO_1350 (O_1350,N_23175,N_22864);
and UO_1351 (O_1351,N_24780,N_22567);
or UO_1352 (O_1352,N_22827,N_23148);
nand UO_1353 (O_1353,N_23075,N_23383);
and UO_1354 (O_1354,N_22671,N_24813);
and UO_1355 (O_1355,N_23433,N_23759);
or UO_1356 (O_1356,N_22850,N_23610);
or UO_1357 (O_1357,N_22995,N_24773);
xor UO_1358 (O_1358,N_24695,N_23113);
and UO_1359 (O_1359,N_23146,N_24737);
and UO_1360 (O_1360,N_22738,N_24711);
or UO_1361 (O_1361,N_22997,N_24650);
or UO_1362 (O_1362,N_24985,N_22765);
and UO_1363 (O_1363,N_24103,N_23886);
and UO_1364 (O_1364,N_24889,N_24461);
nor UO_1365 (O_1365,N_22620,N_24328);
or UO_1366 (O_1366,N_24086,N_23058);
nand UO_1367 (O_1367,N_23083,N_23424);
or UO_1368 (O_1368,N_24586,N_24706);
xor UO_1369 (O_1369,N_24386,N_23971);
nand UO_1370 (O_1370,N_24005,N_22682);
or UO_1371 (O_1371,N_23313,N_24077);
or UO_1372 (O_1372,N_24356,N_24624);
nor UO_1373 (O_1373,N_24618,N_24576);
or UO_1374 (O_1374,N_24333,N_24488);
or UO_1375 (O_1375,N_24338,N_22518);
nor UO_1376 (O_1376,N_24515,N_22526);
nor UO_1377 (O_1377,N_24654,N_24737);
or UO_1378 (O_1378,N_23730,N_23018);
xnor UO_1379 (O_1379,N_23466,N_22750);
or UO_1380 (O_1380,N_24078,N_23396);
nand UO_1381 (O_1381,N_24099,N_24982);
or UO_1382 (O_1382,N_23282,N_24554);
nor UO_1383 (O_1383,N_22927,N_23613);
or UO_1384 (O_1384,N_23614,N_24532);
nor UO_1385 (O_1385,N_23745,N_23437);
xnor UO_1386 (O_1386,N_22584,N_22881);
or UO_1387 (O_1387,N_22818,N_24057);
xor UO_1388 (O_1388,N_24485,N_24600);
and UO_1389 (O_1389,N_22834,N_23034);
nor UO_1390 (O_1390,N_23373,N_24093);
and UO_1391 (O_1391,N_23038,N_22655);
nand UO_1392 (O_1392,N_23921,N_24325);
nor UO_1393 (O_1393,N_24075,N_22756);
xnor UO_1394 (O_1394,N_24251,N_24973);
or UO_1395 (O_1395,N_24520,N_23531);
xnor UO_1396 (O_1396,N_24780,N_23255);
nor UO_1397 (O_1397,N_23859,N_23035);
xnor UO_1398 (O_1398,N_24642,N_24152);
nor UO_1399 (O_1399,N_23589,N_22689);
nor UO_1400 (O_1400,N_24063,N_24830);
and UO_1401 (O_1401,N_24657,N_24191);
and UO_1402 (O_1402,N_23368,N_24644);
and UO_1403 (O_1403,N_23502,N_22669);
nor UO_1404 (O_1404,N_24902,N_24752);
nand UO_1405 (O_1405,N_23533,N_23273);
or UO_1406 (O_1406,N_23899,N_24945);
nand UO_1407 (O_1407,N_24570,N_22721);
nand UO_1408 (O_1408,N_24389,N_24011);
or UO_1409 (O_1409,N_24984,N_23427);
and UO_1410 (O_1410,N_24301,N_24957);
or UO_1411 (O_1411,N_23714,N_23187);
and UO_1412 (O_1412,N_23706,N_23896);
nand UO_1413 (O_1413,N_23920,N_22562);
nor UO_1414 (O_1414,N_24585,N_24024);
nor UO_1415 (O_1415,N_22724,N_23788);
nand UO_1416 (O_1416,N_23290,N_22558);
nand UO_1417 (O_1417,N_24964,N_23296);
xor UO_1418 (O_1418,N_23444,N_23534);
and UO_1419 (O_1419,N_24183,N_24216);
xnor UO_1420 (O_1420,N_24612,N_23661);
nor UO_1421 (O_1421,N_24654,N_24458);
xor UO_1422 (O_1422,N_22526,N_23121);
nor UO_1423 (O_1423,N_23369,N_24837);
xnor UO_1424 (O_1424,N_24924,N_24255);
nor UO_1425 (O_1425,N_23517,N_24021);
nand UO_1426 (O_1426,N_23574,N_23345);
nor UO_1427 (O_1427,N_22841,N_23669);
xor UO_1428 (O_1428,N_22704,N_24356);
and UO_1429 (O_1429,N_24262,N_24459);
nor UO_1430 (O_1430,N_22621,N_23109);
xor UO_1431 (O_1431,N_23987,N_23522);
nor UO_1432 (O_1432,N_22560,N_24580);
xnor UO_1433 (O_1433,N_23987,N_24746);
nand UO_1434 (O_1434,N_23062,N_23885);
xor UO_1435 (O_1435,N_23734,N_24294);
nand UO_1436 (O_1436,N_22669,N_23350);
nand UO_1437 (O_1437,N_24609,N_23317);
xor UO_1438 (O_1438,N_22850,N_22676);
nand UO_1439 (O_1439,N_23338,N_22701);
or UO_1440 (O_1440,N_24922,N_23086);
nand UO_1441 (O_1441,N_24482,N_24176);
nor UO_1442 (O_1442,N_23303,N_22857);
or UO_1443 (O_1443,N_24782,N_24230);
nand UO_1444 (O_1444,N_23802,N_22844);
or UO_1445 (O_1445,N_24867,N_22935);
or UO_1446 (O_1446,N_24192,N_23948);
and UO_1447 (O_1447,N_24817,N_23645);
and UO_1448 (O_1448,N_23648,N_23866);
nor UO_1449 (O_1449,N_23861,N_23830);
and UO_1450 (O_1450,N_23255,N_23050);
nand UO_1451 (O_1451,N_22584,N_24139);
xnor UO_1452 (O_1452,N_24289,N_24838);
nand UO_1453 (O_1453,N_23950,N_23599);
nor UO_1454 (O_1454,N_22619,N_24831);
nor UO_1455 (O_1455,N_22577,N_22877);
and UO_1456 (O_1456,N_23105,N_22882);
and UO_1457 (O_1457,N_22636,N_23286);
nand UO_1458 (O_1458,N_22818,N_24086);
nand UO_1459 (O_1459,N_24520,N_23788);
nor UO_1460 (O_1460,N_24239,N_24580);
xor UO_1461 (O_1461,N_24045,N_22602);
xor UO_1462 (O_1462,N_23241,N_23310);
xor UO_1463 (O_1463,N_22739,N_24270);
xnor UO_1464 (O_1464,N_23792,N_24023);
xnor UO_1465 (O_1465,N_24282,N_23559);
nor UO_1466 (O_1466,N_23020,N_24659);
or UO_1467 (O_1467,N_23905,N_23965);
xnor UO_1468 (O_1468,N_24543,N_22651);
and UO_1469 (O_1469,N_23383,N_22650);
and UO_1470 (O_1470,N_24928,N_23200);
nand UO_1471 (O_1471,N_23791,N_22854);
nand UO_1472 (O_1472,N_24199,N_24490);
or UO_1473 (O_1473,N_24641,N_23097);
nor UO_1474 (O_1474,N_24573,N_24493);
or UO_1475 (O_1475,N_24224,N_23616);
nand UO_1476 (O_1476,N_24945,N_22932);
nand UO_1477 (O_1477,N_24568,N_23690);
nand UO_1478 (O_1478,N_23436,N_24443);
nor UO_1479 (O_1479,N_23625,N_24269);
nor UO_1480 (O_1480,N_23541,N_24065);
nand UO_1481 (O_1481,N_24545,N_22629);
nor UO_1482 (O_1482,N_24449,N_22787);
nand UO_1483 (O_1483,N_22515,N_24477);
and UO_1484 (O_1484,N_24555,N_22862);
xor UO_1485 (O_1485,N_24367,N_24040);
nor UO_1486 (O_1486,N_23731,N_24581);
or UO_1487 (O_1487,N_24339,N_24354);
nand UO_1488 (O_1488,N_24202,N_24934);
xor UO_1489 (O_1489,N_24620,N_22874);
xor UO_1490 (O_1490,N_23959,N_24054);
nor UO_1491 (O_1491,N_23936,N_23506);
xnor UO_1492 (O_1492,N_23711,N_24601);
or UO_1493 (O_1493,N_23064,N_22638);
or UO_1494 (O_1494,N_24425,N_23175);
or UO_1495 (O_1495,N_24020,N_24571);
nor UO_1496 (O_1496,N_23393,N_22548);
or UO_1497 (O_1497,N_23006,N_23427);
nand UO_1498 (O_1498,N_22833,N_22975);
and UO_1499 (O_1499,N_24170,N_24950);
and UO_1500 (O_1500,N_24904,N_24380);
xnor UO_1501 (O_1501,N_23620,N_23614);
or UO_1502 (O_1502,N_22737,N_23947);
nand UO_1503 (O_1503,N_22975,N_23547);
nand UO_1504 (O_1504,N_23345,N_23894);
or UO_1505 (O_1505,N_24478,N_23872);
or UO_1506 (O_1506,N_24854,N_24557);
nand UO_1507 (O_1507,N_24110,N_24323);
nand UO_1508 (O_1508,N_23362,N_24792);
xor UO_1509 (O_1509,N_24789,N_24021);
nand UO_1510 (O_1510,N_22671,N_24612);
nor UO_1511 (O_1511,N_24700,N_23589);
and UO_1512 (O_1512,N_24705,N_24679);
xnor UO_1513 (O_1513,N_23941,N_23577);
or UO_1514 (O_1514,N_23437,N_24747);
xor UO_1515 (O_1515,N_22648,N_24937);
xor UO_1516 (O_1516,N_22504,N_22770);
nor UO_1517 (O_1517,N_23912,N_24967);
nand UO_1518 (O_1518,N_24093,N_24195);
or UO_1519 (O_1519,N_23328,N_22765);
nand UO_1520 (O_1520,N_24888,N_24593);
nor UO_1521 (O_1521,N_23843,N_23884);
xor UO_1522 (O_1522,N_23684,N_23166);
nor UO_1523 (O_1523,N_22886,N_24649);
and UO_1524 (O_1524,N_23067,N_24982);
xnor UO_1525 (O_1525,N_22717,N_24494);
nand UO_1526 (O_1526,N_24675,N_23092);
nand UO_1527 (O_1527,N_24505,N_23883);
nand UO_1528 (O_1528,N_23189,N_24012);
nor UO_1529 (O_1529,N_24664,N_22643);
nor UO_1530 (O_1530,N_24709,N_24678);
nor UO_1531 (O_1531,N_22840,N_24080);
xor UO_1532 (O_1532,N_22707,N_23669);
nand UO_1533 (O_1533,N_22994,N_22527);
or UO_1534 (O_1534,N_24957,N_22535);
and UO_1535 (O_1535,N_24031,N_23966);
xor UO_1536 (O_1536,N_23466,N_22505);
or UO_1537 (O_1537,N_22912,N_23281);
xnor UO_1538 (O_1538,N_24369,N_23054);
xnor UO_1539 (O_1539,N_23040,N_22766);
nand UO_1540 (O_1540,N_23380,N_23144);
xor UO_1541 (O_1541,N_24668,N_24623);
nand UO_1542 (O_1542,N_24906,N_23965);
nand UO_1543 (O_1543,N_24967,N_24578);
and UO_1544 (O_1544,N_23751,N_23261);
and UO_1545 (O_1545,N_22576,N_23831);
and UO_1546 (O_1546,N_24296,N_24849);
nand UO_1547 (O_1547,N_23461,N_24261);
xor UO_1548 (O_1548,N_24001,N_23348);
nor UO_1549 (O_1549,N_24216,N_24462);
or UO_1550 (O_1550,N_23416,N_24419);
nor UO_1551 (O_1551,N_24137,N_22720);
nand UO_1552 (O_1552,N_24744,N_22838);
nand UO_1553 (O_1553,N_22859,N_23544);
or UO_1554 (O_1554,N_24708,N_24792);
nor UO_1555 (O_1555,N_22517,N_24155);
or UO_1556 (O_1556,N_23071,N_24536);
and UO_1557 (O_1557,N_24648,N_23220);
or UO_1558 (O_1558,N_23162,N_24672);
or UO_1559 (O_1559,N_24622,N_23491);
xnor UO_1560 (O_1560,N_24757,N_24103);
nand UO_1561 (O_1561,N_23951,N_23880);
or UO_1562 (O_1562,N_23226,N_22533);
nand UO_1563 (O_1563,N_22796,N_22650);
xor UO_1564 (O_1564,N_24748,N_23759);
and UO_1565 (O_1565,N_24581,N_24845);
and UO_1566 (O_1566,N_24303,N_22511);
nor UO_1567 (O_1567,N_24085,N_23604);
nand UO_1568 (O_1568,N_24335,N_24180);
or UO_1569 (O_1569,N_23577,N_24840);
or UO_1570 (O_1570,N_23125,N_24108);
or UO_1571 (O_1571,N_23643,N_22836);
and UO_1572 (O_1572,N_22563,N_24137);
and UO_1573 (O_1573,N_22875,N_23841);
or UO_1574 (O_1574,N_24819,N_24975);
nor UO_1575 (O_1575,N_23874,N_24640);
xnor UO_1576 (O_1576,N_22616,N_23001);
nor UO_1577 (O_1577,N_22662,N_24857);
and UO_1578 (O_1578,N_23290,N_23556);
and UO_1579 (O_1579,N_22943,N_23017);
and UO_1580 (O_1580,N_24705,N_22944);
nand UO_1581 (O_1581,N_24438,N_23389);
nor UO_1582 (O_1582,N_23436,N_24911);
nand UO_1583 (O_1583,N_23178,N_23073);
and UO_1584 (O_1584,N_23001,N_23018);
nand UO_1585 (O_1585,N_24905,N_24281);
or UO_1586 (O_1586,N_23195,N_22557);
and UO_1587 (O_1587,N_24483,N_23877);
nor UO_1588 (O_1588,N_23091,N_23461);
and UO_1589 (O_1589,N_23925,N_24504);
or UO_1590 (O_1590,N_23555,N_23026);
and UO_1591 (O_1591,N_23369,N_23610);
or UO_1592 (O_1592,N_24203,N_23442);
nand UO_1593 (O_1593,N_24364,N_23134);
and UO_1594 (O_1594,N_23978,N_24153);
and UO_1595 (O_1595,N_24242,N_24215);
xnor UO_1596 (O_1596,N_23353,N_22886);
and UO_1597 (O_1597,N_24843,N_24857);
nor UO_1598 (O_1598,N_23676,N_23050);
xnor UO_1599 (O_1599,N_24013,N_24248);
and UO_1600 (O_1600,N_24845,N_24349);
nor UO_1601 (O_1601,N_24158,N_23471);
xor UO_1602 (O_1602,N_24346,N_23920);
or UO_1603 (O_1603,N_23713,N_22698);
xnor UO_1604 (O_1604,N_22673,N_24090);
and UO_1605 (O_1605,N_23554,N_23442);
nand UO_1606 (O_1606,N_24205,N_23008);
and UO_1607 (O_1607,N_22638,N_23641);
or UO_1608 (O_1608,N_22660,N_23412);
xor UO_1609 (O_1609,N_24160,N_23829);
and UO_1610 (O_1610,N_24502,N_24867);
nand UO_1611 (O_1611,N_24721,N_23648);
or UO_1612 (O_1612,N_24882,N_23399);
and UO_1613 (O_1613,N_23932,N_23936);
and UO_1614 (O_1614,N_22608,N_24788);
and UO_1615 (O_1615,N_23732,N_23939);
and UO_1616 (O_1616,N_23901,N_23436);
nor UO_1617 (O_1617,N_23441,N_23705);
nand UO_1618 (O_1618,N_23279,N_23536);
nor UO_1619 (O_1619,N_22559,N_23285);
nor UO_1620 (O_1620,N_23279,N_22538);
nand UO_1621 (O_1621,N_22761,N_23183);
nand UO_1622 (O_1622,N_23460,N_23480);
nand UO_1623 (O_1623,N_22669,N_24610);
and UO_1624 (O_1624,N_23509,N_23641);
nor UO_1625 (O_1625,N_22816,N_24701);
and UO_1626 (O_1626,N_24585,N_23148);
nor UO_1627 (O_1627,N_23326,N_22883);
nor UO_1628 (O_1628,N_22806,N_23957);
and UO_1629 (O_1629,N_23274,N_24329);
nand UO_1630 (O_1630,N_23959,N_23499);
nand UO_1631 (O_1631,N_22579,N_22767);
and UO_1632 (O_1632,N_22535,N_23133);
or UO_1633 (O_1633,N_23085,N_24159);
and UO_1634 (O_1634,N_24814,N_23787);
nor UO_1635 (O_1635,N_23852,N_24058);
nor UO_1636 (O_1636,N_24911,N_22604);
or UO_1637 (O_1637,N_24023,N_23891);
xor UO_1638 (O_1638,N_23209,N_24273);
xor UO_1639 (O_1639,N_23869,N_24893);
xor UO_1640 (O_1640,N_23059,N_22827);
nand UO_1641 (O_1641,N_23471,N_22758);
or UO_1642 (O_1642,N_22573,N_23311);
nor UO_1643 (O_1643,N_24282,N_23465);
and UO_1644 (O_1644,N_23937,N_23007);
xnor UO_1645 (O_1645,N_24391,N_22850);
nor UO_1646 (O_1646,N_24398,N_24446);
and UO_1647 (O_1647,N_23350,N_24817);
nor UO_1648 (O_1648,N_23954,N_24034);
or UO_1649 (O_1649,N_23215,N_24037);
or UO_1650 (O_1650,N_24279,N_24673);
nand UO_1651 (O_1651,N_24919,N_22881);
and UO_1652 (O_1652,N_22925,N_23973);
or UO_1653 (O_1653,N_23728,N_22832);
or UO_1654 (O_1654,N_22559,N_24342);
nand UO_1655 (O_1655,N_24186,N_24029);
nor UO_1656 (O_1656,N_24061,N_24798);
and UO_1657 (O_1657,N_23103,N_24902);
and UO_1658 (O_1658,N_24543,N_24794);
xor UO_1659 (O_1659,N_23146,N_22558);
and UO_1660 (O_1660,N_23145,N_24638);
or UO_1661 (O_1661,N_23088,N_22752);
nor UO_1662 (O_1662,N_22866,N_23812);
nand UO_1663 (O_1663,N_23635,N_23802);
nand UO_1664 (O_1664,N_24902,N_24054);
nor UO_1665 (O_1665,N_24043,N_24552);
nand UO_1666 (O_1666,N_23702,N_23422);
nor UO_1667 (O_1667,N_24243,N_23383);
nor UO_1668 (O_1668,N_22669,N_24269);
nor UO_1669 (O_1669,N_24544,N_23327);
and UO_1670 (O_1670,N_24268,N_22670);
xnor UO_1671 (O_1671,N_24748,N_23514);
xor UO_1672 (O_1672,N_23393,N_24917);
or UO_1673 (O_1673,N_24525,N_22725);
and UO_1674 (O_1674,N_23925,N_23035);
or UO_1675 (O_1675,N_24372,N_22533);
nor UO_1676 (O_1676,N_23714,N_24770);
nor UO_1677 (O_1677,N_24695,N_23015);
nor UO_1678 (O_1678,N_24984,N_23586);
and UO_1679 (O_1679,N_22989,N_23910);
nor UO_1680 (O_1680,N_23796,N_24231);
or UO_1681 (O_1681,N_23074,N_24472);
nor UO_1682 (O_1682,N_23818,N_24270);
and UO_1683 (O_1683,N_23582,N_23723);
nor UO_1684 (O_1684,N_23847,N_23284);
or UO_1685 (O_1685,N_24748,N_23228);
nor UO_1686 (O_1686,N_24211,N_23388);
and UO_1687 (O_1687,N_24952,N_24584);
xor UO_1688 (O_1688,N_22958,N_24401);
nor UO_1689 (O_1689,N_23378,N_23584);
xor UO_1690 (O_1690,N_22621,N_24709);
or UO_1691 (O_1691,N_23613,N_24462);
xor UO_1692 (O_1692,N_22590,N_23705);
nor UO_1693 (O_1693,N_22578,N_24515);
nor UO_1694 (O_1694,N_24554,N_23836);
or UO_1695 (O_1695,N_23988,N_22634);
nor UO_1696 (O_1696,N_24969,N_24734);
or UO_1697 (O_1697,N_24359,N_24785);
or UO_1698 (O_1698,N_23069,N_23397);
xnor UO_1699 (O_1699,N_23960,N_22887);
or UO_1700 (O_1700,N_23647,N_24269);
xor UO_1701 (O_1701,N_24541,N_23175);
nand UO_1702 (O_1702,N_24409,N_24193);
xnor UO_1703 (O_1703,N_24323,N_22500);
nor UO_1704 (O_1704,N_24798,N_23153);
and UO_1705 (O_1705,N_23959,N_24791);
nor UO_1706 (O_1706,N_24956,N_22770);
or UO_1707 (O_1707,N_23503,N_22612);
nor UO_1708 (O_1708,N_24856,N_24494);
nand UO_1709 (O_1709,N_23444,N_23505);
xor UO_1710 (O_1710,N_23279,N_23940);
and UO_1711 (O_1711,N_24426,N_22990);
nor UO_1712 (O_1712,N_23123,N_24467);
nand UO_1713 (O_1713,N_22684,N_23217);
nor UO_1714 (O_1714,N_22617,N_23889);
or UO_1715 (O_1715,N_24451,N_23815);
nor UO_1716 (O_1716,N_24834,N_24391);
xnor UO_1717 (O_1717,N_23492,N_23985);
and UO_1718 (O_1718,N_23762,N_23246);
nor UO_1719 (O_1719,N_23706,N_24888);
or UO_1720 (O_1720,N_23606,N_22941);
nand UO_1721 (O_1721,N_22840,N_23535);
and UO_1722 (O_1722,N_24230,N_24383);
or UO_1723 (O_1723,N_22831,N_22693);
nand UO_1724 (O_1724,N_23264,N_23809);
nand UO_1725 (O_1725,N_23676,N_23468);
or UO_1726 (O_1726,N_23099,N_24784);
nand UO_1727 (O_1727,N_24103,N_23865);
nand UO_1728 (O_1728,N_24318,N_22571);
nand UO_1729 (O_1729,N_24422,N_22669);
xnor UO_1730 (O_1730,N_23214,N_23346);
xor UO_1731 (O_1731,N_24008,N_22903);
xnor UO_1732 (O_1732,N_23121,N_23035);
or UO_1733 (O_1733,N_23444,N_23263);
nand UO_1734 (O_1734,N_23646,N_24224);
or UO_1735 (O_1735,N_23339,N_23479);
nor UO_1736 (O_1736,N_23896,N_22652);
nor UO_1737 (O_1737,N_23632,N_24268);
and UO_1738 (O_1738,N_22600,N_24949);
nand UO_1739 (O_1739,N_22701,N_24046);
or UO_1740 (O_1740,N_24712,N_24227);
nor UO_1741 (O_1741,N_24159,N_22666);
nor UO_1742 (O_1742,N_23707,N_23218);
and UO_1743 (O_1743,N_23052,N_22794);
xor UO_1744 (O_1744,N_22645,N_24201);
nand UO_1745 (O_1745,N_24545,N_24600);
or UO_1746 (O_1746,N_22905,N_23535);
and UO_1747 (O_1747,N_23697,N_22522);
nor UO_1748 (O_1748,N_23998,N_24857);
and UO_1749 (O_1749,N_23900,N_23017);
xnor UO_1750 (O_1750,N_23118,N_24851);
or UO_1751 (O_1751,N_24273,N_23401);
xnor UO_1752 (O_1752,N_24105,N_23773);
nand UO_1753 (O_1753,N_23499,N_23045);
nand UO_1754 (O_1754,N_24146,N_23813);
and UO_1755 (O_1755,N_24989,N_24772);
nand UO_1756 (O_1756,N_23307,N_23884);
or UO_1757 (O_1757,N_23853,N_24203);
nand UO_1758 (O_1758,N_23872,N_23436);
xor UO_1759 (O_1759,N_23999,N_23678);
nand UO_1760 (O_1760,N_24283,N_24987);
xor UO_1761 (O_1761,N_24054,N_24141);
nor UO_1762 (O_1762,N_23619,N_22907);
xnor UO_1763 (O_1763,N_24523,N_23720);
nor UO_1764 (O_1764,N_24087,N_23150);
nand UO_1765 (O_1765,N_22964,N_23202);
nand UO_1766 (O_1766,N_23389,N_23764);
nor UO_1767 (O_1767,N_22664,N_22591);
xor UO_1768 (O_1768,N_24168,N_23819);
and UO_1769 (O_1769,N_23192,N_22639);
nand UO_1770 (O_1770,N_23032,N_24960);
xor UO_1771 (O_1771,N_24424,N_23908);
or UO_1772 (O_1772,N_22954,N_22529);
xnor UO_1773 (O_1773,N_23377,N_22945);
nand UO_1774 (O_1774,N_22992,N_24965);
or UO_1775 (O_1775,N_22798,N_24085);
or UO_1776 (O_1776,N_22881,N_23022);
nor UO_1777 (O_1777,N_23320,N_23765);
xor UO_1778 (O_1778,N_22569,N_23716);
or UO_1779 (O_1779,N_24638,N_24139);
nor UO_1780 (O_1780,N_23905,N_22787);
xor UO_1781 (O_1781,N_23023,N_22818);
xnor UO_1782 (O_1782,N_24181,N_24201);
and UO_1783 (O_1783,N_24564,N_22612);
xnor UO_1784 (O_1784,N_22726,N_23055);
and UO_1785 (O_1785,N_24202,N_23178);
nor UO_1786 (O_1786,N_24393,N_24248);
and UO_1787 (O_1787,N_24478,N_23757);
and UO_1788 (O_1788,N_23229,N_24262);
or UO_1789 (O_1789,N_23317,N_23830);
and UO_1790 (O_1790,N_22592,N_22542);
nor UO_1791 (O_1791,N_24208,N_23652);
or UO_1792 (O_1792,N_24289,N_23178);
or UO_1793 (O_1793,N_23003,N_22885);
and UO_1794 (O_1794,N_22803,N_23164);
and UO_1795 (O_1795,N_23433,N_23864);
nand UO_1796 (O_1796,N_23384,N_23024);
or UO_1797 (O_1797,N_23213,N_22527);
or UO_1798 (O_1798,N_23233,N_22586);
nor UO_1799 (O_1799,N_23380,N_24340);
xor UO_1800 (O_1800,N_24037,N_23698);
nor UO_1801 (O_1801,N_22806,N_23038);
and UO_1802 (O_1802,N_22591,N_24336);
nand UO_1803 (O_1803,N_22732,N_23159);
nor UO_1804 (O_1804,N_22678,N_23918);
nor UO_1805 (O_1805,N_24375,N_23353);
and UO_1806 (O_1806,N_22692,N_22757);
nor UO_1807 (O_1807,N_23903,N_22621);
and UO_1808 (O_1808,N_24523,N_24085);
xor UO_1809 (O_1809,N_24920,N_22708);
xnor UO_1810 (O_1810,N_24634,N_24346);
xnor UO_1811 (O_1811,N_23643,N_23313);
and UO_1812 (O_1812,N_23282,N_24246);
and UO_1813 (O_1813,N_24173,N_23982);
nor UO_1814 (O_1814,N_22630,N_24879);
nor UO_1815 (O_1815,N_24353,N_24281);
xnor UO_1816 (O_1816,N_24057,N_23547);
or UO_1817 (O_1817,N_24250,N_23685);
nand UO_1818 (O_1818,N_22732,N_23192);
nor UO_1819 (O_1819,N_24890,N_23279);
and UO_1820 (O_1820,N_24324,N_22822);
or UO_1821 (O_1821,N_22695,N_22761);
or UO_1822 (O_1822,N_23516,N_22541);
xnor UO_1823 (O_1823,N_24799,N_24271);
xnor UO_1824 (O_1824,N_24492,N_22866);
or UO_1825 (O_1825,N_22504,N_23342);
or UO_1826 (O_1826,N_22842,N_22784);
and UO_1827 (O_1827,N_23120,N_24901);
or UO_1828 (O_1828,N_24130,N_24102);
nand UO_1829 (O_1829,N_24698,N_24543);
nor UO_1830 (O_1830,N_22700,N_23906);
or UO_1831 (O_1831,N_23144,N_22887);
and UO_1832 (O_1832,N_24310,N_24535);
nand UO_1833 (O_1833,N_24274,N_23299);
or UO_1834 (O_1834,N_23376,N_24553);
and UO_1835 (O_1835,N_22663,N_24894);
or UO_1836 (O_1836,N_23117,N_23135);
and UO_1837 (O_1837,N_23437,N_23829);
and UO_1838 (O_1838,N_23086,N_24074);
xnor UO_1839 (O_1839,N_24754,N_24895);
or UO_1840 (O_1840,N_24839,N_23526);
or UO_1841 (O_1841,N_23445,N_24441);
or UO_1842 (O_1842,N_23891,N_24511);
or UO_1843 (O_1843,N_23665,N_23081);
nor UO_1844 (O_1844,N_24756,N_24531);
nor UO_1845 (O_1845,N_23047,N_24206);
nand UO_1846 (O_1846,N_23053,N_24438);
and UO_1847 (O_1847,N_23248,N_24972);
nand UO_1848 (O_1848,N_23512,N_23552);
and UO_1849 (O_1849,N_23969,N_23768);
or UO_1850 (O_1850,N_24975,N_24202);
nand UO_1851 (O_1851,N_24505,N_23999);
nand UO_1852 (O_1852,N_24373,N_24724);
nand UO_1853 (O_1853,N_24630,N_24322);
nand UO_1854 (O_1854,N_22927,N_24241);
xnor UO_1855 (O_1855,N_24743,N_24631);
nor UO_1856 (O_1856,N_23488,N_22745);
nor UO_1857 (O_1857,N_23089,N_23086);
or UO_1858 (O_1858,N_24002,N_23604);
xor UO_1859 (O_1859,N_23095,N_23418);
and UO_1860 (O_1860,N_24524,N_23285);
xor UO_1861 (O_1861,N_23243,N_22795);
or UO_1862 (O_1862,N_22857,N_23413);
and UO_1863 (O_1863,N_24911,N_23931);
or UO_1864 (O_1864,N_23897,N_23867);
nand UO_1865 (O_1865,N_24460,N_24794);
and UO_1866 (O_1866,N_24064,N_23672);
and UO_1867 (O_1867,N_22954,N_23576);
xnor UO_1868 (O_1868,N_23672,N_23915);
nand UO_1869 (O_1869,N_24450,N_24593);
or UO_1870 (O_1870,N_23239,N_24306);
or UO_1871 (O_1871,N_23800,N_22829);
and UO_1872 (O_1872,N_24023,N_23698);
xor UO_1873 (O_1873,N_24038,N_24833);
nor UO_1874 (O_1874,N_22581,N_22790);
nor UO_1875 (O_1875,N_24310,N_24867);
nor UO_1876 (O_1876,N_24986,N_23433);
nand UO_1877 (O_1877,N_23153,N_23452);
xor UO_1878 (O_1878,N_23817,N_24609);
nand UO_1879 (O_1879,N_24660,N_23509);
nand UO_1880 (O_1880,N_22927,N_24544);
xnor UO_1881 (O_1881,N_23706,N_24112);
and UO_1882 (O_1882,N_23198,N_22590);
or UO_1883 (O_1883,N_22979,N_24470);
or UO_1884 (O_1884,N_22837,N_24637);
xor UO_1885 (O_1885,N_23837,N_22788);
nor UO_1886 (O_1886,N_22970,N_22586);
xnor UO_1887 (O_1887,N_22818,N_24055);
and UO_1888 (O_1888,N_24224,N_24636);
xnor UO_1889 (O_1889,N_23195,N_24250);
and UO_1890 (O_1890,N_24133,N_23526);
or UO_1891 (O_1891,N_23353,N_24938);
xnor UO_1892 (O_1892,N_23590,N_23975);
nor UO_1893 (O_1893,N_24715,N_24987);
or UO_1894 (O_1894,N_22878,N_23623);
nor UO_1895 (O_1895,N_24151,N_23512);
or UO_1896 (O_1896,N_23425,N_23407);
nand UO_1897 (O_1897,N_23493,N_24668);
and UO_1898 (O_1898,N_23034,N_24441);
nor UO_1899 (O_1899,N_22535,N_24138);
or UO_1900 (O_1900,N_23755,N_23542);
xor UO_1901 (O_1901,N_23058,N_24958);
or UO_1902 (O_1902,N_24969,N_22939);
xor UO_1903 (O_1903,N_23901,N_22993);
or UO_1904 (O_1904,N_24224,N_24548);
nor UO_1905 (O_1905,N_23471,N_24261);
xnor UO_1906 (O_1906,N_22748,N_22709);
nand UO_1907 (O_1907,N_24680,N_23836);
and UO_1908 (O_1908,N_23502,N_24187);
and UO_1909 (O_1909,N_22828,N_22548);
xor UO_1910 (O_1910,N_23990,N_22629);
nand UO_1911 (O_1911,N_24775,N_23649);
xor UO_1912 (O_1912,N_23064,N_24313);
nand UO_1913 (O_1913,N_22731,N_24640);
or UO_1914 (O_1914,N_22597,N_24441);
xor UO_1915 (O_1915,N_22802,N_23291);
or UO_1916 (O_1916,N_23086,N_23451);
or UO_1917 (O_1917,N_24168,N_24606);
xor UO_1918 (O_1918,N_24801,N_22529);
and UO_1919 (O_1919,N_24373,N_23241);
and UO_1920 (O_1920,N_23814,N_23959);
nand UO_1921 (O_1921,N_24758,N_24051);
and UO_1922 (O_1922,N_22774,N_24913);
or UO_1923 (O_1923,N_23708,N_24906);
or UO_1924 (O_1924,N_24242,N_24693);
nor UO_1925 (O_1925,N_24817,N_22505);
or UO_1926 (O_1926,N_24718,N_22519);
xnor UO_1927 (O_1927,N_22814,N_24936);
nand UO_1928 (O_1928,N_23394,N_22859);
or UO_1929 (O_1929,N_23418,N_22559);
xnor UO_1930 (O_1930,N_24989,N_23463);
and UO_1931 (O_1931,N_22750,N_24321);
and UO_1932 (O_1932,N_22616,N_24700);
and UO_1933 (O_1933,N_23803,N_24647);
nor UO_1934 (O_1934,N_24640,N_23674);
nor UO_1935 (O_1935,N_24311,N_22550);
nor UO_1936 (O_1936,N_24943,N_22569);
xnor UO_1937 (O_1937,N_23802,N_23790);
nand UO_1938 (O_1938,N_23086,N_24474);
xnor UO_1939 (O_1939,N_23824,N_24274);
and UO_1940 (O_1940,N_22850,N_24587);
nor UO_1941 (O_1941,N_24782,N_23421);
or UO_1942 (O_1942,N_22593,N_23595);
and UO_1943 (O_1943,N_22738,N_22966);
and UO_1944 (O_1944,N_23978,N_22898);
or UO_1945 (O_1945,N_22868,N_22863);
nor UO_1946 (O_1946,N_24744,N_24925);
or UO_1947 (O_1947,N_23036,N_23771);
and UO_1948 (O_1948,N_23393,N_24180);
nand UO_1949 (O_1949,N_23432,N_24492);
nand UO_1950 (O_1950,N_24629,N_24416);
and UO_1951 (O_1951,N_23986,N_24724);
or UO_1952 (O_1952,N_23419,N_24228);
nor UO_1953 (O_1953,N_24246,N_24406);
and UO_1954 (O_1954,N_24043,N_24056);
nor UO_1955 (O_1955,N_22842,N_24437);
nand UO_1956 (O_1956,N_22883,N_22872);
or UO_1957 (O_1957,N_22692,N_24707);
xnor UO_1958 (O_1958,N_24089,N_24874);
nand UO_1959 (O_1959,N_23930,N_23215);
nor UO_1960 (O_1960,N_23596,N_22829);
or UO_1961 (O_1961,N_23091,N_23924);
nand UO_1962 (O_1962,N_23132,N_22623);
xor UO_1963 (O_1963,N_24534,N_23743);
xnor UO_1964 (O_1964,N_23119,N_22923);
or UO_1965 (O_1965,N_23540,N_23205);
nand UO_1966 (O_1966,N_23811,N_23493);
nor UO_1967 (O_1967,N_23741,N_24112);
xor UO_1968 (O_1968,N_24306,N_22627);
xor UO_1969 (O_1969,N_22942,N_23870);
and UO_1970 (O_1970,N_23352,N_24661);
nand UO_1971 (O_1971,N_22936,N_23723);
nand UO_1972 (O_1972,N_24708,N_23497);
nand UO_1973 (O_1973,N_22500,N_24616);
and UO_1974 (O_1974,N_23765,N_22761);
nand UO_1975 (O_1975,N_23752,N_22647);
nand UO_1976 (O_1976,N_23169,N_24778);
and UO_1977 (O_1977,N_22502,N_23019);
and UO_1978 (O_1978,N_24297,N_24331);
and UO_1979 (O_1979,N_23285,N_23722);
and UO_1980 (O_1980,N_24772,N_23214);
and UO_1981 (O_1981,N_24380,N_22900);
xnor UO_1982 (O_1982,N_24567,N_24886);
and UO_1983 (O_1983,N_24609,N_23781);
nand UO_1984 (O_1984,N_22924,N_24589);
or UO_1985 (O_1985,N_23889,N_24846);
or UO_1986 (O_1986,N_22508,N_23331);
or UO_1987 (O_1987,N_22606,N_24344);
and UO_1988 (O_1988,N_24738,N_24291);
nand UO_1989 (O_1989,N_23279,N_24947);
nand UO_1990 (O_1990,N_24060,N_23609);
and UO_1991 (O_1991,N_22572,N_23909);
nand UO_1992 (O_1992,N_23661,N_24479);
xor UO_1993 (O_1993,N_22568,N_24679);
xnor UO_1994 (O_1994,N_24674,N_23724);
xor UO_1995 (O_1995,N_23424,N_23403);
or UO_1996 (O_1996,N_22777,N_24821);
nor UO_1997 (O_1997,N_24178,N_24923);
nor UO_1998 (O_1998,N_24333,N_22560);
or UO_1999 (O_1999,N_23952,N_23256);
nor UO_2000 (O_2000,N_23935,N_23414);
and UO_2001 (O_2001,N_23298,N_23807);
and UO_2002 (O_2002,N_23177,N_22589);
and UO_2003 (O_2003,N_23184,N_24145);
and UO_2004 (O_2004,N_22721,N_24832);
nand UO_2005 (O_2005,N_22766,N_22585);
xnor UO_2006 (O_2006,N_24419,N_23023);
nand UO_2007 (O_2007,N_24638,N_24478);
nand UO_2008 (O_2008,N_22690,N_24152);
nand UO_2009 (O_2009,N_23432,N_22759);
nand UO_2010 (O_2010,N_23471,N_24686);
xor UO_2011 (O_2011,N_23605,N_24964);
or UO_2012 (O_2012,N_24121,N_22737);
nand UO_2013 (O_2013,N_24046,N_24356);
and UO_2014 (O_2014,N_23596,N_23862);
nand UO_2015 (O_2015,N_23210,N_22929);
and UO_2016 (O_2016,N_23953,N_22906);
nor UO_2017 (O_2017,N_23345,N_23652);
and UO_2018 (O_2018,N_23439,N_23851);
and UO_2019 (O_2019,N_24566,N_23326);
nor UO_2020 (O_2020,N_24893,N_23935);
xor UO_2021 (O_2021,N_24961,N_23215);
or UO_2022 (O_2022,N_24058,N_23981);
or UO_2023 (O_2023,N_24424,N_22623);
nor UO_2024 (O_2024,N_23040,N_23242);
nor UO_2025 (O_2025,N_22810,N_24890);
or UO_2026 (O_2026,N_23407,N_23012);
xnor UO_2027 (O_2027,N_22799,N_22534);
nand UO_2028 (O_2028,N_24685,N_23466);
and UO_2029 (O_2029,N_23995,N_24011);
nor UO_2030 (O_2030,N_24417,N_24309);
nand UO_2031 (O_2031,N_22765,N_22672);
nand UO_2032 (O_2032,N_24616,N_24506);
xor UO_2033 (O_2033,N_24833,N_22626);
or UO_2034 (O_2034,N_23934,N_22883);
xnor UO_2035 (O_2035,N_22836,N_23514);
and UO_2036 (O_2036,N_22505,N_24683);
nand UO_2037 (O_2037,N_24907,N_23712);
and UO_2038 (O_2038,N_22677,N_23241);
and UO_2039 (O_2039,N_22646,N_23441);
xor UO_2040 (O_2040,N_23768,N_22743);
nand UO_2041 (O_2041,N_23302,N_23025);
xnor UO_2042 (O_2042,N_22800,N_24012);
xor UO_2043 (O_2043,N_23011,N_22985);
or UO_2044 (O_2044,N_23356,N_23706);
and UO_2045 (O_2045,N_22742,N_23754);
nor UO_2046 (O_2046,N_24433,N_23487);
nor UO_2047 (O_2047,N_24513,N_22965);
xnor UO_2048 (O_2048,N_24755,N_22864);
or UO_2049 (O_2049,N_24994,N_23881);
and UO_2050 (O_2050,N_24984,N_24452);
and UO_2051 (O_2051,N_23749,N_23690);
nand UO_2052 (O_2052,N_23562,N_23095);
and UO_2053 (O_2053,N_24953,N_23733);
or UO_2054 (O_2054,N_23267,N_24850);
xnor UO_2055 (O_2055,N_22603,N_23409);
nand UO_2056 (O_2056,N_22623,N_24201);
and UO_2057 (O_2057,N_24735,N_24557);
xnor UO_2058 (O_2058,N_22775,N_23515);
and UO_2059 (O_2059,N_24497,N_24150);
nor UO_2060 (O_2060,N_23552,N_23236);
nand UO_2061 (O_2061,N_22782,N_24180);
xor UO_2062 (O_2062,N_24270,N_22912);
xor UO_2063 (O_2063,N_22506,N_23877);
and UO_2064 (O_2064,N_24721,N_23947);
or UO_2065 (O_2065,N_23493,N_24807);
or UO_2066 (O_2066,N_24782,N_23252);
or UO_2067 (O_2067,N_22659,N_23724);
xnor UO_2068 (O_2068,N_22894,N_23366);
nand UO_2069 (O_2069,N_23952,N_23909);
nor UO_2070 (O_2070,N_24997,N_22737);
nand UO_2071 (O_2071,N_24741,N_22629);
nor UO_2072 (O_2072,N_23987,N_23404);
xnor UO_2073 (O_2073,N_22650,N_24092);
or UO_2074 (O_2074,N_23128,N_23634);
nor UO_2075 (O_2075,N_24789,N_22954);
and UO_2076 (O_2076,N_22572,N_23322);
xnor UO_2077 (O_2077,N_22569,N_24956);
xor UO_2078 (O_2078,N_22958,N_23912);
nand UO_2079 (O_2079,N_23796,N_24166);
and UO_2080 (O_2080,N_24030,N_24547);
and UO_2081 (O_2081,N_22556,N_24544);
nor UO_2082 (O_2082,N_24084,N_23497);
nand UO_2083 (O_2083,N_23072,N_23551);
nand UO_2084 (O_2084,N_24088,N_24531);
or UO_2085 (O_2085,N_24821,N_24868);
xor UO_2086 (O_2086,N_24389,N_23843);
nand UO_2087 (O_2087,N_23161,N_23817);
nor UO_2088 (O_2088,N_23149,N_24078);
nor UO_2089 (O_2089,N_23819,N_24513);
or UO_2090 (O_2090,N_24330,N_22812);
or UO_2091 (O_2091,N_23003,N_23529);
nor UO_2092 (O_2092,N_22746,N_24484);
or UO_2093 (O_2093,N_24865,N_24585);
and UO_2094 (O_2094,N_23677,N_22578);
nor UO_2095 (O_2095,N_24306,N_24853);
nor UO_2096 (O_2096,N_23958,N_23103);
xor UO_2097 (O_2097,N_24214,N_23150);
xor UO_2098 (O_2098,N_24891,N_22762);
and UO_2099 (O_2099,N_22830,N_22610);
or UO_2100 (O_2100,N_23359,N_23234);
and UO_2101 (O_2101,N_23140,N_24982);
and UO_2102 (O_2102,N_24209,N_23439);
and UO_2103 (O_2103,N_23976,N_24602);
or UO_2104 (O_2104,N_22956,N_22729);
nand UO_2105 (O_2105,N_24205,N_23435);
and UO_2106 (O_2106,N_24784,N_22708);
or UO_2107 (O_2107,N_23155,N_22527);
nand UO_2108 (O_2108,N_23654,N_23163);
xnor UO_2109 (O_2109,N_24894,N_22745);
and UO_2110 (O_2110,N_23993,N_23055);
nor UO_2111 (O_2111,N_22957,N_23506);
nor UO_2112 (O_2112,N_23495,N_23009);
xnor UO_2113 (O_2113,N_23884,N_23397);
nor UO_2114 (O_2114,N_23331,N_23259);
nand UO_2115 (O_2115,N_23110,N_23261);
or UO_2116 (O_2116,N_23751,N_22840);
xor UO_2117 (O_2117,N_24831,N_22790);
xor UO_2118 (O_2118,N_23740,N_23102);
or UO_2119 (O_2119,N_23240,N_22564);
nand UO_2120 (O_2120,N_23886,N_23262);
or UO_2121 (O_2121,N_23944,N_22894);
xor UO_2122 (O_2122,N_23043,N_23342);
nor UO_2123 (O_2123,N_24253,N_23779);
xor UO_2124 (O_2124,N_22529,N_24204);
nor UO_2125 (O_2125,N_24577,N_24104);
or UO_2126 (O_2126,N_23231,N_24405);
nand UO_2127 (O_2127,N_23498,N_24226);
nand UO_2128 (O_2128,N_22995,N_24702);
or UO_2129 (O_2129,N_24317,N_23978);
nand UO_2130 (O_2130,N_22789,N_24471);
nand UO_2131 (O_2131,N_23666,N_24233);
and UO_2132 (O_2132,N_24509,N_23826);
and UO_2133 (O_2133,N_24379,N_24413);
nand UO_2134 (O_2134,N_24443,N_24166);
or UO_2135 (O_2135,N_24299,N_23628);
xnor UO_2136 (O_2136,N_22627,N_23376);
or UO_2137 (O_2137,N_24388,N_22846);
and UO_2138 (O_2138,N_22951,N_23487);
nor UO_2139 (O_2139,N_22977,N_22804);
xnor UO_2140 (O_2140,N_24494,N_24934);
or UO_2141 (O_2141,N_23590,N_24597);
xnor UO_2142 (O_2142,N_24324,N_22747);
xor UO_2143 (O_2143,N_24244,N_22921);
nand UO_2144 (O_2144,N_22620,N_22676);
nand UO_2145 (O_2145,N_23507,N_23753);
xnor UO_2146 (O_2146,N_24541,N_24997);
and UO_2147 (O_2147,N_23017,N_23212);
nand UO_2148 (O_2148,N_23193,N_22775);
nand UO_2149 (O_2149,N_23148,N_24386);
or UO_2150 (O_2150,N_23647,N_24369);
xnor UO_2151 (O_2151,N_22863,N_22587);
xor UO_2152 (O_2152,N_24018,N_23888);
xnor UO_2153 (O_2153,N_24149,N_22801);
nand UO_2154 (O_2154,N_23230,N_24806);
nand UO_2155 (O_2155,N_22863,N_24687);
nor UO_2156 (O_2156,N_22617,N_23250);
nand UO_2157 (O_2157,N_23081,N_23834);
or UO_2158 (O_2158,N_24696,N_24925);
nand UO_2159 (O_2159,N_24165,N_22923);
xor UO_2160 (O_2160,N_24457,N_24433);
xnor UO_2161 (O_2161,N_24912,N_23675);
nand UO_2162 (O_2162,N_22873,N_24840);
and UO_2163 (O_2163,N_24582,N_22811);
nand UO_2164 (O_2164,N_24641,N_23569);
and UO_2165 (O_2165,N_23878,N_22754);
xor UO_2166 (O_2166,N_22634,N_24736);
and UO_2167 (O_2167,N_22868,N_22661);
or UO_2168 (O_2168,N_22790,N_22938);
nand UO_2169 (O_2169,N_24843,N_22636);
nor UO_2170 (O_2170,N_24050,N_22714);
xnor UO_2171 (O_2171,N_23420,N_24352);
nand UO_2172 (O_2172,N_24778,N_24861);
or UO_2173 (O_2173,N_23944,N_23781);
nor UO_2174 (O_2174,N_24024,N_23240);
and UO_2175 (O_2175,N_23861,N_22731);
or UO_2176 (O_2176,N_22786,N_24473);
or UO_2177 (O_2177,N_24477,N_24719);
xor UO_2178 (O_2178,N_24305,N_23891);
xor UO_2179 (O_2179,N_22670,N_24083);
nor UO_2180 (O_2180,N_24103,N_23428);
xnor UO_2181 (O_2181,N_23959,N_24681);
and UO_2182 (O_2182,N_24633,N_23080);
and UO_2183 (O_2183,N_23292,N_24744);
nand UO_2184 (O_2184,N_24300,N_23586);
nor UO_2185 (O_2185,N_24256,N_22994);
and UO_2186 (O_2186,N_22800,N_22914);
nand UO_2187 (O_2187,N_24047,N_24628);
nand UO_2188 (O_2188,N_23656,N_23667);
xor UO_2189 (O_2189,N_22586,N_24298);
nand UO_2190 (O_2190,N_24038,N_24854);
and UO_2191 (O_2191,N_24361,N_23193);
xnor UO_2192 (O_2192,N_24961,N_23669);
and UO_2193 (O_2193,N_23783,N_22910);
or UO_2194 (O_2194,N_22785,N_22961);
nor UO_2195 (O_2195,N_24626,N_24140);
or UO_2196 (O_2196,N_24145,N_23280);
nand UO_2197 (O_2197,N_23370,N_22985);
xor UO_2198 (O_2198,N_24240,N_23915);
or UO_2199 (O_2199,N_22967,N_24912);
xnor UO_2200 (O_2200,N_24496,N_22797);
or UO_2201 (O_2201,N_24281,N_24124);
xnor UO_2202 (O_2202,N_22702,N_24044);
xor UO_2203 (O_2203,N_24102,N_22728);
and UO_2204 (O_2204,N_24815,N_22615);
or UO_2205 (O_2205,N_24708,N_23358);
nor UO_2206 (O_2206,N_22533,N_22974);
xor UO_2207 (O_2207,N_22927,N_22640);
or UO_2208 (O_2208,N_23402,N_24731);
and UO_2209 (O_2209,N_23725,N_24462);
nand UO_2210 (O_2210,N_24554,N_23380);
xnor UO_2211 (O_2211,N_22728,N_24446);
nor UO_2212 (O_2212,N_24424,N_22501);
and UO_2213 (O_2213,N_22739,N_23748);
or UO_2214 (O_2214,N_23732,N_23591);
nand UO_2215 (O_2215,N_23778,N_22790);
and UO_2216 (O_2216,N_23416,N_24142);
nand UO_2217 (O_2217,N_24949,N_24265);
nand UO_2218 (O_2218,N_24858,N_23903);
nand UO_2219 (O_2219,N_23861,N_24730);
nand UO_2220 (O_2220,N_23312,N_23177);
nor UO_2221 (O_2221,N_24551,N_24054);
xor UO_2222 (O_2222,N_24634,N_24746);
or UO_2223 (O_2223,N_24652,N_24386);
xor UO_2224 (O_2224,N_23819,N_22523);
nor UO_2225 (O_2225,N_23402,N_22963);
nor UO_2226 (O_2226,N_23547,N_23980);
nor UO_2227 (O_2227,N_22579,N_24511);
and UO_2228 (O_2228,N_23664,N_22850);
and UO_2229 (O_2229,N_23965,N_24690);
xnor UO_2230 (O_2230,N_23795,N_24751);
and UO_2231 (O_2231,N_24906,N_23887);
and UO_2232 (O_2232,N_23692,N_24377);
or UO_2233 (O_2233,N_23937,N_22676);
and UO_2234 (O_2234,N_23149,N_24843);
nor UO_2235 (O_2235,N_24481,N_22952);
xnor UO_2236 (O_2236,N_23439,N_23753);
xnor UO_2237 (O_2237,N_22833,N_24616);
xor UO_2238 (O_2238,N_23552,N_22849);
or UO_2239 (O_2239,N_23354,N_22587);
xor UO_2240 (O_2240,N_23957,N_22932);
nand UO_2241 (O_2241,N_24420,N_23391);
xor UO_2242 (O_2242,N_23441,N_24323);
or UO_2243 (O_2243,N_23054,N_24334);
xnor UO_2244 (O_2244,N_24076,N_23646);
xor UO_2245 (O_2245,N_24027,N_24905);
xnor UO_2246 (O_2246,N_23369,N_24078);
or UO_2247 (O_2247,N_22507,N_24137);
nor UO_2248 (O_2248,N_22564,N_23886);
and UO_2249 (O_2249,N_22686,N_23590);
xnor UO_2250 (O_2250,N_22903,N_23989);
and UO_2251 (O_2251,N_23881,N_23137);
nor UO_2252 (O_2252,N_23545,N_23375);
nor UO_2253 (O_2253,N_23423,N_23300);
xor UO_2254 (O_2254,N_24650,N_23975);
or UO_2255 (O_2255,N_23332,N_24852);
or UO_2256 (O_2256,N_24031,N_24898);
or UO_2257 (O_2257,N_23598,N_23631);
and UO_2258 (O_2258,N_24680,N_23806);
xor UO_2259 (O_2259,N_23391,N_23613);
xor UO_2260 (O_2260,N_24339,N_22669);
or UO_2261 (O_2261,N_23461,N_24033);
and UO_2262 (O_2262,N_24029,N_23028);
and UO_2263 (O_2263,N_22915,N_23705);
or UO_2264 (O_2264,N_23847,N_24847);
nor UO_2265 (O_2265,N_24935,N_22853);
or UO_2266 (O_2266,N_24092,N_23326);
or UO_2267 (O_2267,N_23447,N_23089);
nor UO_2268 (O_2268,N_24318,N_23077);
xnor UO_2269 (O_2269,N_23488,N_23252);
nor UO_2270 (O_2270,N_22924,N_24250);
and UO_2271 (O_2271,N_23758,N_22935);
nand UO_2272 (O_2272,N_24006,N_24382);
nand UO_2273 (O_2273,N_23779,N_23721);
nor UO_2274 (O_2274,N_23344,N_23835);
xnor UO_2275 (O_2275,N_24419,N_22608);
or UO_2276 (O_2276,N_23006,N_23242);
and UO_2277 (O_2277,N_23523,N_22901);
nand UO_2278 (O_2278,N_22912,N_24734);
xnor UO_2279 (O_2279,N_24719,N_24993);
nor UO_2280 (O_2280,N_22564,N_24486);
nand UO_2281 (O_2281,N_23921,N_23278);
nand UO_2282 (O_2282,N_23767,N_24508);
nor UO_2283 (O_2283,N_22632,N_23782);
or UO_2284 (O_2284,N_24235,N_23184);
nor UO_2285 (O_2285,N_24175,N_22853);
nor UO_2286 (O_2286,N_23213,N_23720);
and UO_2287 (O_2287,N_24320,N_24227);
or UO_2288 (O_2288,N_23576,N_22718);
nor UO_2289 (O_2289,N_23486,N_22651);
xnor UO_2290 (O_2290,N_24679,N_23514);
nand UO_2291 (O_2291,N_23291,N_22723);
and UO_2292 (O_2292,N_24318,N_23122);
or UO_2293 (O_2293,N_23705,N_24144);
or UO_2294 (O_2294,N_22895,N_22859);
nand UO_2295 (O_2295,N_23050,N_24106);
xnor UO_2296 (O_2296,N_24459,N_23207);
xnor UO_2297 (O_2297,N_24412,N_23493);
xor UO_2298 (O_2298,N_23964,N_23705);
or UO_2299 (O_2299,N_22657,N_23085);
xnor UO_2300 (O_2300,N_23987,N_23489);
and UO_2301 (O_2301,N_23125,N_24537);
or UO_2302 (O_2302,N_22567,N_23855);
and UO_2303 (O_2303,N_23623,N_23417);
and UO_2304 (O_2304,N_22839,N_23307);
or UO_2305 (O_2305,N_22868,N_23802);
xnor UO_2306 (O_2306,N_24431,N_24568);
and UO_2307 (O_2307,N_23686,N_22727);
and UO_2308 (O_2308,N_24158,N_23643);
and UO_2309 (O_2309,N_24478,N_23118);
and UO_2310 (O_2310,N_24029,N_23754);
or UO_2311 (O_2311,N_22960,N_22677);
and UO_2312 (O_2312,N_23581,N_23272);
nor UO_2313 (O_2313,N_23440,N_23293);
nand UO_2314 (O_2314,N_23609,N_24476);
and UO_2315 (O_2315,N_22708,N_23991);
and UO_2316 (O_2316,N_24720,N_24036);
or UO_2317 (O_2317,N_23123,N_24053);
xnor UO_2318 (O_2318,N_23098,N_23748);
nand UO_2319 (O_2319,N_24313,N_24334);
xor UO_2320 (O_2320,N_22924,N_23532);
nor UO_2321 (O_2321,N_24403,N_24543);
nor UO_2322 (O_2322,N_23537,N_23929);
nand UO_2323 (O_2323,N_23952,N_24079);
nand UO_2324 (O_2324,N_23758,N_24517);
nor UO_2325 (O_2325,N_23937,N_22506);
or UO_2326 (O_2326,N_22857,N_23366);
and UO_2327 (O_2327,N_23828,N_24713);
or UO_2328 (O_2328,N_24051,N_22679);
or UO_2329 (O_2329,N_23797,N_22618);
or UO_2330 (O_2330,N_23487,N_23540);
or UO_2331 (O_2331,N_23619,N_22620);
and UO_2332 (O_2332,N_23323,N_24101);
nor UO_2333 (O_2333,N_23827,N_23116);
or UO_2334 (O_2334,N_23041,N_23451);
and UO_2335 (O_2335,N_24074,N_22822);
or UO_2336 (O_2336,N_24712,N_23906);
or UO_2337 (O_2337,N_23180,N_23779);
xnor UO_2338 (O_2338,N_23429,N_23716);
nand UO_2339 (O_2339,N_22782,N_22810);
and UO_2340 (O_2340,N_23072,N_23894);
and UO_2341 (O_2341,N_23140,N_23142);
and UO_2342 (O_2342,N_23632,N_24792);
or UO_2343 (O_2343,N_24217,N_24622);
nand UO_2344 (O_2344,N_22647,N_23276);
and UO_2345 (O_2345,N_22964,N_24104);
nand UO_2346 (O_2346,N_24177,N_23922);
or UO_2347 (O_2347,N_23733,N_24062);
or UO_2348 (O_2348,N_24635,N_24845);
and UO_2349 (O_2349,N_24079,N_24318);
or UO_2350 (O_2350,N_22587,N_22521);
or UO_2351 (O_2351,N_24309,N_22817);
nor UO_2352 (O_2352,N_24785,N_24586);
nand UO_2353 (O_2353,N_23158,N_24310);
or UO_2354 (O_2354,N_24433,N_24080);
and UO_2355 (O_2355,N_23933,N_22583);
nand UO_2356 (O_2356,N_23797,N_22808);
or UO_2357 (O_2357,N_24602,N_24555);
nor UO_2358 (O_2358,N_23326,N_23952);
xor UO_2359 (O_2359,N_23819,N_22678);
nor UO_2360 (O_2360,N_23268,N_24077);
and UO_2361 (O_2361,N_23917,N_22724);
or UO_2362 (O_2362,N_24097,N_24536);
or UO_2363 (O_2363,N_23586,N_23283);
and UO_2364 (O_2364,N_24488,N_23765);
xor UO_2365 (O_2365,N_24365,N_24924);
and UO_2366 (O_2366,N_24395,N_24907);
and UO_2367 (O_2367,N_22744,N_24027);
nor UO_2368 (O_2368,N_22787,N_24339);
nand UO_2369 (O_2369,N_22824,N_23627);
and UO_2370 (O_2370,N_24877,N_23547);
nor UO_2371 (O_2371,N_23044,N_24814);
or UO_2372 (O_2372,N_24401,N_22648);
nor UO_2373 (O_2373,N_24754,N_22830);
or UO_2374 (O_2374,N_23060,N_23486);
xnor UO_2375 (O_2375,N_24069,N_23816);
nor UO_2376 (O_2376,N_22730,N_23293);
nor UO_2377 (O_2377,N_23841,N_23633);
or UO_2378 (O_2378,N_23641,N_23053);
or UO_2379 (O_2379,N_22716,N_23008);
nand UO_2380 (O_2380,N_23566,N_24296);
or UO_2381 (O_2381,N_24138,N_24391);
xor UO_2382 (O_2382,N_24097,N_22824);
and UO_2383 (O_2383,N_22980,N_23238);
nor UO_2384 (O_2384,N_23463,N_24171);
nand UO_2385 (O_2385,N_24724,N_22888);
or UO_2386 (O_2386,N_23222,N_23858);
and UO_2387 (O_2387,N_24301,N_24289);
nor UO_2388 (O_2388,N_23897,N_24896);
and UO_2389 (O_2389,N_24350,N_23306);
and UO_2390 (O_2390,N_23743,N_24386);
and UO_2391 (O_2391,N_23158,N_22602);
or UO_2392 (O_2392,N_22796,N_23517);
or UO_2393 (O_2393,N_24593,N_24332);
and UO_2394 (O_2394,N_22701,N_22985);
nand UO_2395 (O_2395,N_24978,N_23399);
nor UO_2396 (O_2396,N_22964,N_22954);
nor UO_2397 (O_2397,N_22851,N_23293);
and UO_2398 (O_2398,N_23889,N_24577);
or UO_2399 (O_2399,N_22542,N_22506);
or UO_2400 (O_2400,N_23667,N_24509);
nand UO_2401 (O_2401,N_22930,N_24289);
nand UO_2402 (O_2402,N_23775,N_23106);
nand UO_2403 (O_2403,N_23694,N_23366);
nand UO_2404 (O_2404,N_24184,N_23364);
nand UO_2405 (O_2405,N_22757,N_22948);
and UO_2406 (O_2406,N_22784,N_23794);
or UO_2407 (O_2407,N_24575,N_22752);
nor UO_2408 (O_2408,N_22959,N_24477);
or UO_2409 (O_2409,N_23299,N_23752);
nand UO_2410 (O_2410,N_24405,N_24194);
nand UO_2411 (O_2411,N_22531,N_24148);
xor UO_2412 (O_2412,N_23837,N_23533);
xor UO_2413 (O_2413,N_22744,N_22923);
nand UO_2414 (O_2414,N_24507,N_22638);
nand UO_2415 (O_2415,N_23367,N_24902);
xnor UO_2416 (O_2416,N_23048,N_24344);
nor UO_2417 (O_2417,N_24632,N_24446);
nor UO_2418 (O_2418,N_24327,N_22885);
and UO_2419 (O_2419,N_22758,N_22530);
xor UO_2420 (O_2420,N_23789,N_24812);
or UO_2421 (O_2421,N_23121,N_24126);
xor UO_2422 (O_2422,N_23170,N_22748);
nor UO_2423 (O_2423,N_23995,N_24517);
or UO_2424 (O_2424,N_22840,N_24901);
or UO_2425 (O_2425,N_23144,N_24444);
xor UO_2426 (O_2426,N_23785,N_24656);
xor UO_2427 (O_2427,N_23668,N_24182);
nor UO_2428 (O_2428,N_22800,N_23267);
nand UO_2429 (O_2429,N_22691,N_22819);
xor UO_2430 (O_2430,N_22918,N_24179);
or UO_2431 (O_2431,N_23390,N_22708);
xnor UO_2432 (O_2432,N_24494,N_23572);
nor UO_2433 (O_2433,N_23403,N_23263);
nor UO_2434 (O_2434,N_24156,N_24957);
nand UO_2435 (O_2435,N_22736,N_24900);
or UO_2436 (O_2436,N_23276,N_24596);
nand UO_2437 (O_2437,N_24902,N_22842);
and UO_2438 (O_2438,N_22755,N_23242);
or UO_2439 (O_2439,N_22501,N_22571);
nor UO_2440 (O_2440,N_24078,N_22900);
xnor UO_2441 (O_2441,N_23116,N_23681);
and UO_2442 (O_2442,N_23449,N_23725);
or UO_2443 (O_2443,N_24355,N_22720);
and UO_2444 (O_2444,N_24530,N_23178);
xor UO_2445 (O_2445,N_24882,N_23800);
nand UO_2446 (O_2446,N_22853,N_24732);
xnor UO_2447 (O_2447,N_24090,N_22701);
and UO_2448 (O_2448,N_23284,N_22713);
or UO_2449 (O_2449,N_23570,N_23878);
or UO_2450 (O_2450,N_23560,N_23850);
or UO_2451 (O_2451,N_23244,N_22962);
and UO_2452 (O_2452,N_23920,N_22772);
and UO_2453 (O_2453,N_24894,N_22753);
and UO_2454 (O_2454,N_23142,N_23874);
nand UO_2455 (O_2455,N_23588,N_23790);
nor UO_2456 (O_2456,N_23315,N_23038);
nand UO_2457 (O_2457,N_23660,N_24817);
nand UO_2458 (O_2458,N_23943,N_23843);
nor UO_2459 (O_2459,N_24822,N_22597);
nor UO_2460 (O_2460,N_22516,N_23405);
or UO_2461 (O_2461,N_24982,N_24403);
or UO_2462 (O_2462,N_24052,N_22526);
nand UO_2463 (O_2463,N_22757,N_23406);
or UO_2464 (O_2464,N_23868,N_24703);
nor UO_2465 (O_2465,N_24181,N_23541);
and UO_2466 (O_2466,N_24310,N_22963);
and UO_2467 (O_2467,N_23259,N_23130);
and UO_2468 (O_2468,N_24354,N_23507);
xnor UO_2469 (O_2469,N_22695,N_23602);
nor UO_2470 (O_2470,N_24808,N_23016);
nor UO_2471 (O_2471,N_23475,N_23147);
nand UO_2472 (O_2472,N_22905,N_23246);
and UO_2473 (O_2473,N_22939,N_22541);
xnor UO_2474 (O_2474,N_22859,N_23781);
nor UO_2475 (O_2475,N_22768,N_22846);
nand UO_2476 (O_2476,N_23744,N_24276);
or UO_2477 (O_2477,N_22907,N_22971);
xor UO_2478 (O_2478,N_23341,N_23044);
nor UO_2479 (O_2479,N_22965,N_24022);
nor UO_2480 (O_2480,N_22598,N_24836);
xor UO_2481 (O_2481,N_23029,N_23851);
xor UO_2482 (O_2482,N_24490,N_23279);
or UO_2483 (O_2483,N_22543,N_24976);
nand UO_2484 (O_2484,N_24439,N_23490);
nor UO_2485 (O_2485,N_23180,N_23248);
xnor UO_2486 (O_2486,N_22788,N_24971);
or UO_2487 (O_2487,N_23100,N_24280);
nor UO_2488 (O_2488,N_24641,N_23447);
nor UO_2489 (O_2489,N_24056,N_23307);
or UO_2490 (O_2490,N_24408,N_23308);
nor UO_2491 (O_2491,N_24117,N_22503);
nand UO_2492 (O_2492,N_24678,N_24943);
nor UO_2493 (O_2493,N_23305,N_23069);
nand UO_2494 (O_2494,N_23223,N_24960);
xnor UO_2495 (O_2495,N_22722,N_22910);
nand UO_2496 (O_2496,N_24494,N_24424);
or UO_2497 (O_2497,N_24124,N_22527);
and UO_2498 (O_2498,N_24739,N_23894);
nor UO_2499 (O_2499,N_23100,N_23594);
or UO_2500 (O_2500,N_24494,N_22557);
or UO_2501 (O_2501,N_24487,N_23993);
and UO_2502 (O_2502,N_23516,N_24167);
nand UO_2503 (O_2503,N_24709,N_23944);
nand UO_2504 (O_2504,N_24075,N_23475);
nand UO_2505 (O_2505,N_22662,N_23660);
or UO_2506 (O_2506,N_22503,N_23468);
nand UO_2507 (O_2507,N_24275,N_24421);
xnor UO_2508 (O_2508,N_23308,N_22975);
xnor UO_2509 (O_2509,N_24122,N_24513);
or UO_2510 (O_2510,N_24792,N_22561);
and UO_2511 (O_2511,N_24317,N_24353);
and UO_2512 (O_2512,N_23820,N_23314);
or UO_2513 (O_2513,N_23568,N_23211);
nor UO_2514 (O_2514,N_24000,N_24095);
nor UO_2515 (O_2515,N_24597,N_23707);
and UO_2516 (O_2516,N_24891,N_23444);
nand UO_2517 (O_2517,N_24392,N_23737);
nand UO_2518 (O_2518,N_23566,N_22879);
xor UO_2519 (O_2519,N_24265,N_23326);
xnor UO_2520 (O_2520,N_24942,N_22517);
or UO_2521 (O_2521,N_23378,N_23538);
nor UO_2522 (O_2522,N_24209,N_22962);
xnor UO_2523 (O_2523,N_24010,N_23700);
nor UO_2524 (O_2524,N_24806,N_22722);
nand UO_2525 (O_2525,N_23753,N_24112);
nor UO_2526 (O_2526,N_23186,N_23239);
nor UO_2527 (O_2527,N_24881,N_23072);
and UO_2528 (O_2528,N_23312,N_24458);
or UO_2529 (O_2529,N_23578,N_24575);
and UO_2530 (O_2530,N_24760,N_23581);
or UO_2531 (O_2531,N_23490,N_23594);
nand UO_2532 (O_2532,N_23823,N_22702);
or UO_2533 (O_2533,N_23502,N_24134);
xor UO_2534 (O_2534,N_22999,N_24455);
nor UO_2535 (O_2535,N_24420,N_22621);
nor UO_2536 (O_2536,N_24107,N_22529);
or UO_2537 (O_2537,N_23970,N_24805);
or UO_2538 (O_2538,N_24377,N_23214);
nor UO_2539 (O_2539,N_24601,N_24619);
nor UO_2540 (O_2540,N_24285,N_23743);
nand UO_2541 (O_2541,N_23359,N_24210);
nand UO_2542 (O_2542,N_24753,N_24861);
xor UO_2543 (O_2543,N_22779,N_23655);
and UO_2544 (O_2544,N_24718,N_22563);
nand UO_2545 (O_2545,N_22626,N_22882);
and UO_2546 (O_2546,N_23496,N_24776);
nor UO_2547 (O_2547,N_24256,N_23747);
nor UO_2548 (O_2548,N_24342,N_22963);
and UO_2549 (O_2549,N_24663,N_23848);
or UO_2550 (O_2550,N_23527,N_22804);
nor UO_2551 (O_2551,N_22843,N_23793);
nor UO_2552 (O_2552,N_22671,N_23863);
or UO_2553 (O_2553,N_24305,N_23080);
or UO_2554 (O_2554,N_22673,N_23356);
xnor UO_2555 (O_2555,N_23614,N_24887);
nor UO_2556 (O_2556,N_24743,N_23701);
nand UO_2557 (O_2557,N_23592,N_23263);
nand UO_2558 (O_2558,N_22599,N_23827);
nor UO_2559 (O_2559,N_22569,N_23978);
or UO_2560 (O_2560,N_24822,N_23213);
xnor UO_2561 (O_2561,N_24075,N_24506);
or UO_2562 (O_2562,N_22625,N_23194);
xor UO_2563 (O_2563,N_23084,N_23827);
and UO_2564 (O_2564,N_22585,N_24544);
and UO_2565 (O_2565,N_23772,N_23551);
or UO_2566 (O_2566,N_24192,N_23573);
and UO_2567 (O_2567,N_23380,N_22794);
or UO_2568 (O_2568,N_24395,N_23934);
nand UO_2569 (O_2569,N_23270,N_22941);
nand UO_2570 (O_2570,N_22514,N_23196);
or UO_2571 (O_2571,N_24510,N_24915);
nor UO_2572 (O_2572,N_23959,N_22543);
nor UO_2573 (O_2573,N_24697,N_24505);
or UO_2574 (O_2574,N_23633,N_24734);
nor UO_2575 (O_2575,N_24550,N_23854);
xnor UO_2576 (O_2576,N_23072,N_22700);
or UO_2577 (O_2577,N_23456,N_24434);
and UO_2578 (O_2578,N_22609,N_23886);
nor UO_2579 (O_2579,N_23167,N_24917);
nor UO_2580 (O_2580,N_24395,N_22989);
xnor UO_2581 (O_2581,N_23783,N_23661);
or UO_2582 (O_2582,N_23794,N_23460);
nand UO_2583 (O_2583,N_24973,N_22554);
nor UO_2584 (O_2584,N_24968,N_24587);
or UO_2585 (O_2585,N_22943,N_22698);
nand UO_2586 (O_2586,N_22695,N_23127);
and UO_2587 (O_2587,N_23008,N_24823);
nor UO_2588 (O_2588,N_24865,N_24258);
xor UO_2589 (O_2589,N_23006,N_24117);
and UO_2590 (O_2590,N_23621,N_23202);
nand UO_2591 (O_2591,N_23466,N_22677);
xor UO_2592 (O_2592,N_24568,N_23581);
nor UO_2593 (O_2593,N_22585,N_23716);
xor UO_2594 (O_2594,N_23190,N_23559);
or UO_2595 (O_2595,N_24413,N_24882);
or UO_2596 (O_2596,N_22824,N_23615);
xnor UO_2597 (O_2597,N_24755,N_24076);
xor UO_2598 (O_2598,N_24476,N_23843);
and UO_2599 (O_2599,N_24705,N_24531);
nor UO_2600 (O_2600,N_23461,N_22903);
xor UO_2601 (O_2601,N_24144,N_24908);
and UO_2602 (O_2602,N_22988,N_23483);
and UO_2603 (O_2603,N_23556,N_23465);
xor UO_2604 (O_2604,N_23848,N_23446);
and UO_2605 (O_2605,N_24883,N_24885);
nand UO_2606 (O_2606,N_23420,N_24524);
nor UO_2607 (O_2607,N_23119,N_22828);
nor UO_2608 (O_2608,N_22932,N_24914);
nor UO_2609 (O_2609,N_24977,N_23527);
and UO_2610 (O_2610,N_23968,N_24444);
xor UO_2611 (O_2611,N_24594,N_23800);
or UO_2612 (O_2612,N_23777,N_24437);
and UO_2613 (O_2613,N_24950,N_23281);
or UO_2614 (O_2614,N_23188,N_22631);
or UO_2615 (O_2615,N_22749,N_23510);
or UO_2616 (O_2616,N_23007,N_24586);
xor UO_2617 (O_2617,N_22958,N_24442);
xor UO_2618 (O_2618,N_23888,N_24174);
xnor UO_2619 (O_2619,N_22849,N_24757);
xnor UO_2620 (O_2620,N_24488,N_23426);
xor UO_2621 (O_2621,N_23472,N_23806);
or UO_2622 (O_2622,N_24083,N_22663);
or UO_2623 (O_2623,N_24735,N_22785);
or UO_2624 (O_2624,N_22534,N_24209);
or UO_2625 (O_2625,N_23173,N_23669);
nor UO_2626 (O_2626,N_22750,N_24306);
nand UO_2627 (O_2627,N_23056,N_24330);
or UO_2628 (O_2628,N_23144,N_24801);
xnor UO_2629 (O_2629,N_24414,N_22875);
nor UO_2630 (O_2630,N_23047,N_23118);
and UO_2631 (O_2631,N_23350,N_22848);
and UO_2632 (O_2632,N_23319,N_23654);
or UO_2633 (O_2633,N_23416,N_22842);
and UO_2634 (O_2634,N_22565,N_22746);
xor UO_2635 (O_2635,N_22744,N_23280);
nand UO_2636 (O_2636,N_23397,N_24316);
or UO_2637 (O_2637,N_24139,N_24237);
or UO_2638 (O_2638,N_22976,N_24657);
nand UO_2639 (O_2639,N_23077,N_24162);
or UO_2640 (O_2640,N_24322,N_22984);
xor UO_2641 (O_2641,N_24046,N_23208);
nand UO_2642 (O_2642,N_22646,N_23946);
and UO_2643 (O_2643,N_24552,N_23531);
nor UO_2644 (O_2644,N_23799,N_23969);
nand UO_2645 (O_2645,N_23060,N_24022);
nand UO_2646 (O_2646,N_24280,N_24000);
xnor UO_2647 (O_2647,N_23827,N_24829);
nand UO_2648 (O_2648,N_22523,N_23875);
xnor UO_2649 (O_2649,N_23800,N_24752);
xor UO_2650 (O_2650,N_22845,N_22864);
and UO_2651 (O_2651,N_22718,N_23362);
xor UO_2652 (O_2652,N_24776,N_23695);
xnor UO_2653 (O_2653,N_24150,N_22607);
or UO_2654 (O_2654,N_22750,N_24848);
nor UO_2655 (O_2655,N_24092,N_23778);
nor UO_2656 (O_2656,N_24077,N_23415);
xor UO_2657 (O_2657,N_23154,N_22695);
or UO_2658 (O_2658,N_23397,N_24853);
and UO_2659 (O_2659,N_23385,N_24616);
nor UO_2660 (O_2660,N_24501,N_24272);
nor UO_2661 (O_2661,N_24242,N_24193);
and UO_2662 (O_2662,N_23479,N_24564);
nand UO_2663 (O_2663,N_23763,N_24867);
or UO_2664 (O_2664,N_24327,N_24715);
nor UO_2665 (O_2665,N_24060,N_24447);
nand UO_2666 (O_2666,N_23116,N_23187);
nand UO_2667 (O_2667,N_23403,N_22939);
nand UO_2668 (O_2668,N_24226,N_24608);
nor UO_2669 (O_2669,N_23416,N_23887);
and UO_2670 (O_2670,N_24849,N_24433);
or UO_2671 (O_2671,N_22607,N_24789);
nand UO_2672 (O_2672,N_23297,N_24787);
xnor UO_2673 (O_2673,N_23504,N_23421);
nor UO_2674 (O_2674,N_22932,N_22855);
or UO_2675 (O_2675,N_24118,N_24534);
nand UO_2676 (O_2676,N_23520,N_23098);
or UO_2677 (O_2677,N_23867,N_23136);
and UO_2678 (O_2678,N_24376,N_23951);
xnor UO_2679 (O_2679,N_24126,N_24082);
nor UO_2680 (O_2680,N_24038,N_24620);
nand UO_2681 (O_2681,N_22751,N_22966);
or UO_2682 (O_2682,N_24764,N_22693);
nand UO_2683 (O_2683,N_24381,N_22847);
and UO_2684 (O_2684,N_23130,N_23612);
nor UO_2685 (O_2685,N_22792,N_23892);
and UO_2686 (O_2686,N_24157,N_24091);
or UO_2687 (O_2687,N_22699,N_24338);
nand UO_2688 (O_2688,N_23578,N_23345);
or UO_2689 (O_2689,N_24985,N_23759);
xor UO_2690 (O_2690,N_23780,N_24619);
nand UO_2691 (O_2691,N_24709,N_23728);
nand UO_2692 (O_2692,N_23013,N_23356);
and UO_2693 (O_2693,N_23082,N_24090);
xor UO_2694 (O_2694,N_23867,N_23387);
and UO_2695 (O_2695,N_24739,N_22750);
or UO_2696 (O_2696,N_24081,N_23741);
xor UO_2697 (O_2697,N_24384,N_24169);
nand UO_2698 (O_2698,N_22748,N_24311);
and UO_2699 (O_2699,N_22623,N_24740);
nand UO_2700 (O_2700,N_24749,N_24253);
or UO_2701 (O_2701,N_24726,N_22958);
and UO_2702 (O_2702,N_22509,N_23640);
or UO_2703 (O_2703,N_24245,N_23059);
nand UO_2704 (O_2704,N_24278,N_22849);
nor UO_2705 (O_2705,N_24063,N_24075);
nor UO_2706 (O_2706,N_22813,N_24556);
nand UO_2707 (O_2707,N_24661,N_22508);
nand UO_2708 (O_2708,N_24658,N_22559);
nor UO_2709 (O_2709,N_23813,N_23388);
nand UO_2710 (O_2710,N_23989,N_22851);
nor UO_2711 (O_2711,N_23274,N_23767);
and UO_2712 (O_2712,N_23496,N_22945);
and UO_2713 (O_2713,N_24785,N_24892);
xor UO_2714 (O_2714,N_24795,N_23554);
xnor UO_2715 (O_2715,N_24549,N_24144);
nand UO_2716 (O_2716,N_23438,N_23923);
nor UO_2717 (O_2717,N_22880,N_22667);
and UO_2718 (O_2718,N_23037,N_24378);
nand UO_2719 (O_2719,N_24113,N_23179);
nor UO_2720 (O_2720,N_24339,N_23837);
nor UO_2721 (O_2721,N_23229,N_24403);
and UO_2722 (O_2722,N_23593,N_24345);
nor UO_2723 (O_2723,N_24614,N_24009);
xor UO_2724 (O_2724,N_22619,N_23746);
nand UO_2725 (O_2725,N_22734,N_24078);
and UO_2726 (O_2726,N_22820,N_24692);
or UO_2727 (O_2727,N_23830,N_24271);
nor UO_2728 (O_2728,N_24660,N_22964);
nor UO_2729 (O_2729,N_24482,N_23797);
and UO_2730 (O_2730,N_22745,N_24265);
nor UO_2731 (O_2731,N_24737,N_24034);
nor UO_2732 (O_2732,N_24025,N_24252);
nand UO_2733 (O_2733,N_24076,N_24026);
nand UO_2734 (O_2734,N_24849,N_24674);
and UO_2735 (O_2735,N_22514,N_23494);
nand UO_2736 (O_2736,N_24062,N_24692);
or UO_2737 (O_2737,N_24901,N_24288);
or UO_2738 (O_2738,N_24954,N_23946);
xnor UO_2739 (O_2739,N_24667,N_22821);
and UO_2740 (O_2740,N_22719,N_23482);
or UO_2741 (O_2741,N_24274,N_24081);
xnor UO_2742 (O_2742,N_24076,N_23444);
xnor UO_2743 (O_2743,N_24486,N_24652);
nand UO_2744 (O_2744,N_24049,N_23256);
and UO_2745 (O_2745,N_22970,N_24118);
or UO_2746 (O_2746,N_24698,N_23855);
xor UO_2747 (O_2747,N_24623,N_22932);
nor UO_2748 (O_2748,N_24741,N_22622);
xnor UO_2749 (O_2749,N_23806,N_23125);
xnor UO_2750 (O_2750,N_22628,N_24752);
nor UO_2751 (O_2751,N_24482,N_24475);
and UO_2752 (O_2752,N_22851,N_22607);
xor UO_2753 (O_2753,N_24764,N_23707);
nand UO_2754 (O_2754,N_22793,N_23875);
nand UO_2755 (O_2755,N_22529,N_24624);
nor UO_2756 (O_2756,N_23496,N_24184);
and UO_2757 (O_2757,N_23609,N_24877);
xnor UO_2758 (O_2758,N_23813,N_23955);
nand UO_2759 (O_2759,N_22686,N_23882);
nand UO_2760 (O_2760,N_23793,N_24417);
or UO_2761 (O_2761,N_23438,N_24923);
xor UO_2762 (O_2762,N_24411,N_23517);
and UO_2763 (O_2763,N_23386,N_23729);
nand UO_2764 (O_2764,N_22522,N_22776);
and UO_2765 (O_2765,N_24992,N_23929);
nand UO_2766 (O_2766,N_24971,N_23593);
or UO_2767 (O_2767,N_23155,N_22595);
nor UO_2768 (O_2768,N_24064,N_22755);
nor UO_2769 (O_2769,N_24568,N_23352);
and UO_2770 (O_2770,N_24663,N_23271);
xnor UO_2771 (O_2771,N_23690,N_24885);
and UO_2772 (O_2772,N_22549,N_23216);
xor UO_2773 (O_2773,N_23607,N_24473);
and UO_2774 (O_2774,N_23708,N_22551);
nand UO_2775 (O_2775,N_22515,N_24089);
xor UO_2776 (O_2776,N_23554,N_24973);
nand UO_2777 (O_2777,N_24433,N_23207);
nand UO_2778 (O_2778,N_23339,N_23365);
or UO_2779 (O_2779,N_23983,N_24063);
nor UO_2780 (O_2780,N_24071,N_24615);
xor UO_2781 (O_2781,N_22527,N_23064);
xor UO_2782 (O_2782,N_22620,N_23766);
or UO_2783 (O_2783,N_24787,N_23550);
or UO_2784 (O_2784,N_22771,N_24319);
or UO_2785 (O_2785,N_22916,N_22570);
xnor UO_2786 (O_2786,N_22536,N_23186);
nor UO_2787 (O_2787,N_24363,N_24029);
or UO_2788 (O_2788,N_23148,N_24487);
xor UO_2789 (O_2789,N_23970,N_23539);
nor UO_2790 (O_2790,N_24880,N_23098);
nand UO_2791 (O_2791,N_22824,N_24074);
xnor UO_2792 (O_2792,N_22751,N_23016);
and UO_2793 (O_2793,N_24386,N_24137);
nor UO_2794 (O_2794,N_23829,N_24463);
and UO_2795 (O_2795,N_22606,N_23511);
nand UO_2796 (O_2796,N_24793,N_24919);
nor UO_2797 (O_2797,N_24988,N_24325);
nand UO_2798 (O_2798,N_24004,N_24278);
nor UO_2799 (O_2799,N_23269,N_23107);
nor UO_2800 (O_2800,N_23436,N_24949);
nor UO_2801 (O_2801,N_23096,N_23658);
and UO_2802 (O_2802,N_24298,N_24759);
nand UO_2803 (O_2803,N_22988,N_24518);
and UO_2804 (O_2804,N_24265,N_22850);
nand UO_2805 (O_2805,N_24900,N_22975);
xor UO_2806 (O_2806,N_23441,N_24153);
and UO_2807 (O_2807,N_23148,N_23753);
nand UO_2808 (O_2808,N_24170,N_24619);
nor UO_2809 (O_2809,N_24666,N_23546);
nor UO_2810 (O_2810,N_22794,N_22849);
and UO_2811 (O_2811,N_22968,N_22743);
xnor UO_2812 (O_2812,N_22778,N_23938);
xor UO_2813 (O_2813,N_23638,N_22784);
or UO_2814 (O_2814,N_24325,N_24689);
or UO_2815 (O_2815,N_23587,N_24343);
xnor UO_2816 (O_2816,N_22822,N_23068);
or UO_2817 (O_2817,N_24420,N_24978);
or UO_2818 (O_2818,N_24613,N_22902);
nor UO_2819 (O_2819,N_24546,N_23475);
or UO_2820 (O_2820,N_23965,N_22825);
xor UO_2821 (O_2821,N_24238,N_24626);
nor UO_2822 (O_2822,N_22616,N_24298);
and UO_2823 (O_2823,N_23161,N_22802);
xnor UO_2824 (O_2824,N_24993,N_24266);
or UO_2825 (O_2825,N_23942,N_24576);
nand UO_2826 (O_2826,N_24560,N_23659);
nand UO_2827 (O_2827,N_24291,N_24826);
nand UO_2828 (O_2828,N_23538,N_23460);
nor UO_2829 (O_2829,N_24722,N_23105);
nand UO_2830 (O_2830,N_24390,N_23210);
nor UO_2831 (O_2831,N_24434,N_23283);
and UO_2832 (O_2832,N_22535,N_24026);
nor UO_2833 (O_2833,N_23952,N_23901);
nand UO_2834 (O_2834,N_24864,N_23852);
xnor UO_2835 (O_2835,N_24805,N_22752);
xnor UO_2836 (O_2836,N_23450,N_22643);
xor UO_2837 (O_2837,N_23219,N_23721);
nand UO_2838 (O_2838,N_24714,N_23558);
or UO_2839 (O_2839,N_23843,N_23127);
or UO_2840 (O_2840,N_24608,N_23056);
xnor UO_2841 (O_2841,N_23195,N_23292);
nand UO_2842 (O_2842,N_23304,N_24531);
xor UO_2843 (O_2843,N_23638,N_24835);
or UO_2844 (O_2844,N_24351,N_24851);
or UO_2845 (O_2845,N_23145,N_24454);
nand UO_2846 (O_2846,N_23821,N_22995);
xnor UO_2847 (O_2847,N_22959,N_24097);
or UO_2848 (O_2848,N_24539,N_22846);
nand UO_2849 (O_2849,N_24335,N_23769);
or UO_2850 (O_2850,N_22674,N_24243);
and UO_2851 (O_2851,N_24514,N_24263);
or UO_2852 (O_2852,N_24599,N_22634);
and UO_2853 (O_2853,N_23868,N_22943);
nand UO_2854 (O_2854,N_24509,N_24466);
nand UO_2855 (O_2855,N_22516,N_23189);
nor UO_2856 (O_2856,N_24439,N_24684);
xnor UO_2857 (O_2857,N_24261,N_24179);
xor UO_2858 (O_2858,N_24998,N_24148);
xnor UO_2859 (O_2859,N_22989,N_24913);
nor UO_2860 (O_2860,N_23143,N_23545);
or UO_2861 (O_2861,N_23434,N_24162);
nor UO_2862 (O_2862,N_23895,N_24039);
xor UO_2863 (O_2863,N_22910,N_23373);
nand UO_2864 (O_2864,N_24123,N_24406);
xnor UO_2865 (O_2865,N_22524,N_24665);
or UO_2866 (O_2866,N_24551,N_23832);
nand UO_2867 (O_2867,N_24173,N_23583);
or UO_2868 (O_2868,N_23074,N_22806);
xor UO_2869 (O_2869,N_23372,N_22882);
or UO_2870 (O_2870,N_22609,N_22884);
and UO_2871 (O_2871,N_23183,N_24812);
nor UO_2872 (O_2872,N_24713,N_22899);
or UO_2873 (O_2873,N_23161,N_24494);
nand UO_2874 (O_2874,N_24056,N_24681);
and UO_2875 (O_2875,N_24368,N_23568);
and UO_2876 (O_2876,N_23777,N_24694);
and UO_2877 (O_2877,N_22996,N_24021);
and UO_2878 (O_2878,N_24277,N_24002);
and UO_2879 (O_2879,N_24772,N_24229);
xor UO_2880 (O_2880,N_23943,N_23698);
and UO_2881 (O_2881,N_24505,N_24211);
xnor UO_2882 (O_2882,N_22662,N_23524);
and UO_2883 (O_2883,N_22824,N_24284);
or UO_2884 (O_2884,N_23919,N_23869);
nor UO_2885 (O_2885,N_23164,N_24653);
nand UO_2886 (O_2886,N_24687,N_23600);
nor UO_2887 (O_2887,N_24151,N_23112);
and UO_2888 (O_2888,N_24973,N_24036);
and UO_2889 (O_2889,N_23520,N_24234);
and UO_2890 (O_2890,N_24042,N_24306);
nand UO_2891 (O_2891,N_22670,N_23549);
and UO_2892 (O_2892,N_23011,N_24769);
and UO_2893 (O_2893,N_23309,N_24556);
nor UO_2894 (O_2894,N_23533,N_22899);
and UO_2895 (O_2895,N_23433,N_22757);
and UO_2896 (O_2896,N_22597,N_23451);
nand UO_2897 (O_2897,N_22610,N_23424);
and UO_2898 (O_2898,N_23957,N_23445);
or UO_2899 (O_2899,N_24872,N_23072);
and UO_2900 (O_2900,N_24228,N_23524);
nor UO_2901 (O_2901,N_24924,N_24802);
xor UO_2902 (O_2902,N_22537,N_24921);
xnor UO_2903 (O_2903,N_24974,N_24832);
xnor UO_2904 (O_2904,N_24808,N_23833);
xnor UO_2905 (O_2905,N_23591,N_24772);
xor UO_2906 (O_2906,N_23977,N_22646);
nand UO_2907 (O_2907,N_22994,N_23589);
nand UO_2908 (O_2908,N_24495,N_23271);
xnor UO_2909 (O_2909,N_24642,N_22824);
xnor UO_2910 (O_2910,N_22798,N_23879);
or UO_2911 (O_2911,N_23167,N_24227);
and UO_2912 (O_2912,N_23992,N_22819);
and UO_2913 (O_2913,N_22611,N_22836);
and UO_2914 (O_2914,N_23708,N_23422);
nand UO_2915 (O_2915,N_23119,N_23666);
and UO_2916 (O_2916,N_23604,N_23642);
or UO_2917 (O_2917,N_24721,N_23676);
nor UO_2918 (O_2918,N_23703,N_24353);
nor UO_2919 (O_2919,N_23095,N_23127);
and UO_2920 (O_2920,N_24911,N_23762);
xnor UO_2921 (O_2921,N_23997,N_24429);
nor UO_2922 (O_2922,N_24469,N_24770);
nor UO_2923 (O_2923,N_22655,N_24799);
nor UO_2924 (O_2924,N_22806,N_22934);
nand UO_2925 (O_2925,N_22873,N_23767);
nand UO_2926 (O_2926,N_23063,N_23525);
nand UO_2927 (O_2927,N_23292,N_24266);
nor UO_2928 (O_2928,N_24409,N_24165);
xor UO_2929 (O_2929,N_24576,N_23793);
nor UO_2930 (O_2930,N_22642,N_24977);
or UO_2931 (O_2931,N_23243,N_24759);
nor UO_2932 (O_2932,N_22647,N_24397);
and UO_2933 (O_2933,N_24462,N_23570);
nor UO_2934 (O_2934,N_24155,N_24154);
nor UO_2935 (O_2935,N_22981,N_23171);
xnor UO_2936 (O_2936,N_23094,N_23811);
or UO_2937 (O_2937,N_22629,N_23536);
nand UO_2938 (O_2938,N_23574,N_24563);
nor UO_2939 (O_2939,N_23659,N_23106);
nor UO_2940 (O_2940,N_23330,N_24176);
xnor UO_2941 (O_2941,N_23361,N_23755);
nor UO_2942 (O_2942,N_24010,N_23623);
and UO_2943 (O_2943,N_24807,N_23327);
nand UO_2944 (O_2944,N_24932,N_24110);
nand UO_2945 (O_2945,N_23561,N_24816);
and UO_2946 (O_2946,N_22879,N_23385);
and UO_2947 (O_2947,N_24003,N_24330);
and UO_2948 (O_2948,N_24650,N_23678);
nor UO_2949 (O_2949,N_22901,N_24461);
nor UO_2950 (O_2950,N_24887,N_24031);
nand UO_2951 (O_2951,N_23151,N_24979);
or UO_2952 (O_2952,N_24679,N_24214);
nor UO_2953 (O_2953,N_24812,N_24682);
nand UO_2954 (O_2954,N_24329,N_24039);
or UO_2955 (O_2955,N_22986,N_23194);
xor UO_2956 (O_2956,N_22936,N_22815);
and UO_2957 (O_2957,N_22898,N_24034);
or UO_2958 (O_2958,N_24503,N_22921);
nand UO_2959 (O_2959,N_22811,N_24325);
nand UO_2960 (O_2960,N_22665,N_24671);
and UO_2961 (O_2961,N_23292,N_23118);
nor UO_2962 (O_2962,N_22988,N_24307);
and UO_2963 (O_2963,N_23004,N_24919);
nor UO_2964 (O_2964,N_24033,N_24258);
and UO_2965 (O_2965,N_23010,N_23346);
nand UO_2966 (O_2966,N_23861,N_24943);
xor UO_2967 (O_2967,N_24376,N_24412);
or UO_2968 (O_2968,N_23339,N_23058);
and UO_2969 (O_2969,N_24134,N_23005);
nand UO_2970 (O_2970,N_24216,N_23817);
or UO_2971 (O_2971,N_24429,N_23682);
xor UO_2972 (O_2972,N_23128,N_23178);
or UO_2973 (O_2973,N_23958,N_22611);
xor UO_2974 (O_2974,N_23338,N_23835);
or UO_2975 (O_2975,N_22893,N_24220);
and UO_2976 (O_2976,N_23617,N_22602);
nor UO_2977 (O_2977,N_22946,N_24324);
or UO_2978 (O_2978,N_24309,N_22761);
nand UO_2979 (O_2979,N_24789,N_22801);
xnor UO_2980 (O_2980,N_22826,N_22857);
nor UO_2981 (O_2981,N_24228,N_23665);
and UO_2982 (O_2982,N_23001,N_23924);
xnor UO_2983 (O_2983,N_24161,N_23315);
nand UO_2984 (O_2984,N_22698,N_23702);
nand UO_2985 (O_2985,N_24107,N_23386);
and UO_2986 (O_2986,N_23106,N_22694);
and UO_2987 (O_2987,N_23082,N_23288);
xor UO_2988 (O_2988,N_24895,N_24053);
and UO_2989 (O_2989,N_22711,N_23621);
nor UO_2990 (O_2990,N_24409,N_24309);
nor UO_2991 (O_2991,N_23076,N_24675);
or UO_2992 (O_2992,N_23629,N_24826);
and UO_2993 (O_2993,N_22994,N_24494);
or UO_2994 (O_2994,N_23914,N_24855);
xnor UO_2995 (O_2995,N_23601,N_23807);
nor UO_2996 (O_2996,N_24325,N_22935);
and UO_2997 (O_2997,N_23882,N_24125);
or UO_2998 (O_2998,N_23010,N_23930);
and UO_2999 (O_2999,N_23325,N_24670);
endmodule