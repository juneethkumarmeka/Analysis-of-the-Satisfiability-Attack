module basic_1000_10000_1500_10_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_672,In_55);
or U1 (N_1,In_392,In_382);
xnor U2 (N_2,In_77,In_297);
nor U3 (N_3,In_847,In_659);
or U4 (N_4,In_461,In_12);
xor U5 (N_5,In_264,In_887);
xor U6 (N_6,In_548,In_124);
or U7 (N_7,In_222,In_832);
and U8 (N_8,In_941,In_924);
or U9 (N_9,In_667,In_391);
nand U10 (N_10,In_572,In_878);
nand U11 (N_11,In_576,In_266);
xor U12 (N_12,In_870,In_165);
nor U13 (N_13,In_670,In_387);
xnor U14 (N_14,In_444,In_351);
nor U15 (N_15,In_738,In_586);
or U16 (N_16,In_317,In_554);
nor U17 (N_17,In_830,In_495);
nor U18 (N_18,In_637,In_268);
and U19 (N_19,In_557,In_766);
nand U20 (N_20,In_919,In_189);
and U21 (N_21,In_947,In_786);
nor U22 (N_22,In_997,In_530);
and U23 (N_23,In_730,In_904);
nor U24 (N_24,In_58,In_826);
nor U25 (N_25,In_771,In_116);
nor U26 (N_26,In_521,In_54);
xor U27 (N_27,In_109,In_419);
xnor U28 (N_28,In_307,In_599);
or U29 (N_29,In_596,In_203);
or U30 (N_30,In_200,In_843);
and U31 (N_31,In_119,In_75);
xnor U32 (N_32,In_519,In_6);
nor U33 (N_33,In_179,In_410);
nand U34 (N_34,In_618,In_312);
nand U35 (N_35,In_629,In_964);
xor U36 (N_36,In_68,In_793);
or U37 (N_37,In_885,In_675);
and U38 (N_38,In_676,In_489);
and U39 (N_39,In_161,In_220);
xnor U40 (N_40,In_588,In_398);
nand U41 (N_41,In_869,In_320);
or U42 (N_42,In_17,In_753);
nand U43 (N_43,In_851,In_270);
xnor U44 (N_44,In_673,In_842);
nand U45 (N_45,In_816,In_577);
nand U46 (N_46,In_412,In_810);
xor U47 (N_47,In_978,In_550);
xnor U48 (N_48,In_875,In_132);
nor U49 (N_49,In_634,In_286);
and U50 (N_50,In_206,In_556);
xor U51 (N_51,In_397,In_769);
or U52 (N_52,In_3,In_473);
nand U53 (N_53,In_196,In_724);
nand U54 (N_54,In_224,In_115);
nand U55 (N_55,In_920,In_140);
or U56 (N_56,In_526,In_963);
nor U57 (N_57,In_788,In_815);
nand U58 (N_58,In_479,In_233);
nor U59 (N_59,In_937,In_299);
and U60 (N_60,In_945,In_239);
and U61 (N_61,In_67,In_414);
and U62 (N_62,In_825,In_544);
nand U63 (N_63,In_925,In_765);
and U64 (N_64,In_632,In_418);
nor U65 (N_65,In_462,In_631);
nor U66 (N_66,In_693,In_562);
xnor U67 (N_67,In_610,In_591);
or U68 (N_68,In_792,In_31);
and U69 (N_69,In_638,In_421);
nor U70 (N_70,In_61,In_865);
nand U71 (N_71,In_844,In_368);
nor U72 (N_72,In_129,In_219);
xor U73 (N_73,In_511,In_501);
nor U74 (N_74,In_492,In_290);
nand U75 (N_75,In_982,In_779);
xnor U76 (N_76,In_898,In_147);
nand U77 (N_77,In_795,In_746);
or U78 (N_78,In_587,In_799);
xor U79 (N_79,In_447,In_737);
and U80 (N_80,In_961,In_98);
nor U81 (N_81,In_522,In_893);
and U82 (N_82,In_120,In_274);
nand U83 (N_83,In_452,In_575);
xor U84 (N_84,In_767,In_783);
xnor U85 (N_85,In_278,In_74);
xnor U86 (N_86,In_697,In_62);
nor U87 (N_87,In_143,In_755);
or U88 (N_88,In_190,In_101);
and U89 (N_89,In_216,In_43);
or U90 (N_90,In_326,In_431);
nor U91 (N_91,In_34,In_329);
nor U92 (N_92,In_177,In_877);
nor U93 (N_93,In_87,In_872);
nor U94 (N_94,In_440,In_531);
nand U95 (N_95,In_370,In_520);
nand U96 (N_96,In_926,In_666);
or U97 (N_97,In_929,In_22);
xor U98 (N_98,In_135,In_229);
or U99 (N_99,In_646,In_118);
nand U100 (N_100,In_958,In_453);
nand U101 (N_101,In_623,In_487);
or U102 (N_102,In_363,In_818);
nand U103 (N_103,In_477,In_27);
nand U104 (N_104,In_288,In_934);
or U105 (N_105,In_938,In_366);
nand U106 (N_106,In_959,In_225);
and U107 (N_107,In_51,In_772);
nand U108 (N_108,In_295,In_604);
nor U109 (N_109,In_78,In_207);
or U110 (N_110,In_181,In_498);
and U111 (N_111,In_123,In_867);
and U112 (N_112,In_966,In_99);
xnor U113 (N_113,In_617,In_652);
or U114 (N_114,In_41,In_517);
or U115 (N_115,In_327,In_237);
xor U116 (N_116,In_256,In_324);
or U117 (N_117,In_852,In_968);
or U118 (N_118,In_19,In_45);
xnor U119 (N_119,In_801,In_940);
nor U120 (N_120,In_460,In_349);
nand U121 (N_121,In_276,In_361);
or U122 (N_122,In_267,In_735);
nor U123 (N_123,In_969,In_726);
xor U124 (N_124,In_113,In_60);
nand U125 (N_125,In_86,In_261);
nor U126 (N_126,In_450,In_791);
and U127 (N_127,In_745,In_967);
xnor U128 (N_128,In_987,In_829);
nor U129 (N_129,In_653,In_390);
or U130 (N_130,In_689,In_794);
xor U131 (N_131,In_175,In_752);
or U132 (N_132,In_465,In_640);
nor U133 (N_133,In_664,In_65);
nand U134 (N_134,In_809,In_305);
nand U135 (N_135,In_403,In_104);
nor U136 (N_136,In_152,In_743);
nor U137 (N_137,In_907,In_892);
nor U138 (N_138,In_608,In_992);
or U139 (N_139,In_611,In_525);
xor U140 (N_140,In_318,In_146);
nor U141 (N_141,In_142,In_401);
and U142 (N_142,In_955,In_476);
nor U143 (N_143,In_908,In_499);
or U144 (N_144,In_989,In_407);
xnor U145 (N_145,In_339,In_80);
nor U146 (N_146,In_425,In_536);
nor U147 (N_147,In_985,In_137);
nor U148 (N_148,In_8,In_930);
and U149 (N_149,In_943,In_680);
xor U150 (N_150,In_72,In_448);
and U151 (N_151,In_262,In_645);
xnor U152 (N_152,In_367,In_706);
xor U153 (N_153,In_127,In_903);
or U154 (N_154,In_381,In_833);
xor U155 (N_155,In_580,In_626);
or U156 (N_156,In_770,In_9);
or U157 (N_157,In_496,In_215);
and U158 (N_158,In_131,In_413);
or U159 (N_159,In_861,In_121);
xnor U160 (N_160,In_551,In_927);
nand U161 (N_161,In_889,In_117);
nor U162 (N_162,In_111,In_600);
or U163 (N_163,In_897,In_373);
or U164 (N_164,In_47,In_917);
or U165 (N_165,In_641,In_708);
nand U166 (N_166,In_973,In_26);
xnor U167 (N_167,In_70,In_931);
nand U168 (N_168,In_841,In_506);
nand U169 (N_169,In_356,In_674);
nand U170 (N_170,In_654,In_837);
xor U171 (N_171,In_406,In_376);
and U172 (N_172,In_319,In_482);
nor U173 (N_173,In_516,In_178);
nor U174 (N_174,In_480,In_658);
or U175 (N_175,In_125,In_909);
nor U176 (N_176,In_707,In_911);
and U177 (N_177,In_923,In_56);
nor U178 (N_178,In_170,In_294);
nand U179 (N_179,In_173,In_928);
or U180 (N_180,In_375,In_630);
nand U181 (N_181,In_429,In_221);
and U182 (N_182,In_97,In_729);
xor U183 (N_183,In_463,In_609);
nor U184 (N_184,In_838,In_508);
and U185 (N_185,In_823,In_95);
or U186 (N_186,In_896,In_972);
nand U187 (N_187,In_71,In_570);
nand U188 (N_188,In_628,In_559);
and U189 (N_189,In_773,In_249);
and U190 (N_190,In_332,In_154);
nor U191 (N_191,In_252,In_248);
or U192 (N_192,In_379,In_106);
or U193 (N_193,In_85,In_651);
nor U194 (N_194,In_728,In_820);
or U195 (N_195,In_245,In_979);
nand U196 (N_196,In_643,In_272);
nor U197 (N_197,In_227,In_183);
or U198 (N_198,In_775,In_939);
nor U199 (N_199,In_633,In_824);
or U200 (N_200,In_714,In_442);
nand U201 (N_201,In_310,In_990);
or U202 (N_202,In_690,In_597);
or U203 (N_203,In_991,In_474);
and U204 (N_204,In_731,In_749);
nand U205 (N_205,In_33,In_199);
or U206 (N_206,In_814,In_565);
nand U207 (N_207,In_112,In_141);
xnor U208 (N_208,In_352,In_936);
nand U209 (N_209,In_571,In_157);
nor U210 (N_210,In_662,In_504);
xnor U211 (N_211,In_420,In_529);
and U212 (N_212,In_93,In_204);
nand U213 (N_213,In_346,In_894);
nand U214 (N_214,In_443,In_828);
xnor U215 (N_215,In_144,In_321);
and U216 (N_216,In_541,In_218);
and U217 (N_217,In_136,In_685);
nor U218 (N_218,In_612,In_345);
nor U219 (N_219,In_408,In_343);
or U220 (N_220,In_21,In_171);
and U221 (N_221,In_918,In_0);
or U222 (N_222,In_411,In_754);
and U223 (N_223,In_895,In_426);
or U224 (N_224,In_347,In_240);
or U225 (N_225,In_24,In_478);
and U226 (N_226,In_246,In_621);
xnor U227 (N_227,In_607,In_856);
nor U228 (N_228,In_899,In_291);
nor U229 (N_229,In_946,In_205);
or U230 (N_230,In_732,In_883);
or U231 (N_231,In_836,In_306);
nand U232 (N_232,In_579,In_960);
or U233 (N_233,In_90,In_542);
xnor U234 (N_234,In_874,In_789);
nand U235 (N_235,In_108,In_405);
xor U236 (N_236,In_718,In_581);
nor U237 (N_237,In_563,In_624);
nand U238 (N_238,In_721,In_970);
or U239 (N_239,In_778,In_890);
xnor U240 (N_240,In_153,In_293);
xnor U241 (N_241,In_49,In_906);
nor U242 (N_242,In_300,In_988);
or U243 (N_243,In_255,In_507);
xnor U244 (N_244,In_168,In_20);
and U245 (N_245,In_549,In_176);
nor U246 (N_246,In_759,In_649);
xor U247 (N_247,In_81,In_932);
and U248 (N_248,In_311,In_415);
or U249 (N_249,In_337,In_59);
and U250 (N_250,In_701,In_213);
and U251 (N_251,In_762,In_493);
nor U252 (N_252,In_438,In_423);
nand U253 (N_253,In_582,In_96);
and U254 (N_254,In_601,In_717);
and U255 (N_255,In_271,In_134);
or U256 (N_256,In_314,In_359);
and U257 (N_257,In_226,In_705);
nor U258 (N_258,In_962,In_914);
nor U259 (N_259,In_130,In_469);
xor U260 (N_260,In_921,In_342);
and U261 (N_261,In_558,In_540);
xor U262 (N_262,In_569,In_458);
nor U263 (N_263,In_313,In_485);
xnor U264 (N_264,In_433,In_751);
nand U265 (N_265,In_486,In_163);
or U266 (N_266,In_533,In_302);
xor U267 (N_267,In_583,In_719);
nor U268 (N_268,In_790,In_491);
xor U269 (N_269,In_148,In_845);
or U270 (N_270,In_965,In_949);
nand U271 (N_271,In_538,In_527);
nand U272 (N_272,In_957,In_798);
and U273 (N_273,In_360,In_807);
nor U274 (N_274,In_528,In_364);
xor U275 (N_275,In_287,In_292);
and U276 (N_276,In_734,In_358);
or U277 (N_277,In_275,In_235);
nor U278 (N_278,In_393,In_602);
xnor U279 (N_279,In_615,In_513);
or U280 (N_280,In_396,In_211);
nand U281 (N_281,In_635,In_301);
or U282 (N_282,In_739,In_547);
or U283 (N_283,In_677,In_922);
nand U284 (N_284,In_866,In_644);
xnor U285 (N_285,In_372,In_386);
nor U286 (N_286,In_277,In_518);
nand U287 (N_287,In_912,In_627);
and U288 (N_288,In_834,In_30);
or U289 (N_289,In_683,In_787);
xor U290 (N_290,In_325,In_995);
nor U291 (N_291,In_840,In_999);
or U292 (N_292,In_891,In_150);
or U293 (N_293,In_57,In_503);
nor U294 (N_294,In_819,In_455);
or U295 (N_295,In_354,In_122);
and U296 (N_296,In_915,In_663);
or U297 (N_297,In_335,In_243);
or U298 (N_298,In_484,In_910);
nand U299 (N_299,In_715,In_44);
nor U300 (N_300,In_510,In_858);
and U301 (N_301,In_328,In_155);
or U302 (N_302,In_524,In_13);
nor U303 (N_303,In_839,In_192);
nand U304 (N_304,In_209,In_539);
xnor U305 (N_305,In_811,In_696);
and U306 (N_306,In_91,In_552);
or U307 (N_307,In_713,In_523);
or U308 (N_308,In_172,In_669);
xor U309 (N_309,In_281,In_954);
and U310 (N_310,In_956,In_280);
nand U311 (N_311,In_441,In_747);
and U312 (N_312,In_971,In_258);
nor U313 (N_313,In_863,In_201);
nand U314 (N_314,In_574,In_802);
nor U315 (N_315,In_699,In_813);
and U316 (N_316,In_848,In_232);
xor U317 (N_317,In_236,In_880);
and U318 (N_318,In_590,In_993);
nand U319 (N_319,In_1,In_107);
or U320 (N_320,In_388,In_736);
or U321 (N_321,In_38,In_193);
nor U322 (N_322,In_636,In_468);
and U323 (N_323,In_682,In_244);
nand U324 (N_324,In_620,In_812);
nand U325 (N_325,In_402,In_534);
and U326 (N_326,In_7,In_905);
and U327 (N_327,In_174,In_126);
xor U328 (N_328,In_437,In_944);
nand U329 (N_329,In_350,In_83);
xor U330 (N_330,In_14,In_716);
nand U331 (N_331,In_39,In_29);
and U332 (N_332,In_665,In_785);
xnor U333 (N_333,In_876,In_756);
xor U334 (N_334,In_92,In_76);
nand U335 (N_335,In_849,In_532);
xnor U336 (N_336,In_191,In_854);
nand U337 (N_337,In_254,In_512);
nand U338 (N_338,In_688,In_916);
or U339 (N_339,In_614,In_449);
nor U340 (N_340,In_821,In_657);
nand U341 (N_341,In_166,In_862);
nand U342 (N_342,In_727,In_763);
or U343 (N_343,In_723,In_333);
or U344 (N_344,In_709,In_208);
nand U345 (N_345,In_592,In_758);
or U346 (N_346,In_257,In_655);
nor U347 (N_347,In_984,In_598);
nor U348 (N_348,In_5,In_284);
nand U349 (N_349,In_871,In_500);
and U350 (N_350,In_11,In_231);
and U351 (N_351,In_336,In_416);
xor U352 (N_352,In_855,In_804);
xnor U353 (N_353,In_198,In_975);
nor U354 (N_354,In_377,In_289);
nor U355 (N_355,In_241,In_385);
nor U356 (N_356,In_578,In_466);
nor U357 (N_357,In_269,In_341);
nor U358 (N_358,In_555,In_40);
and U359 (N_359,In_860,In_744);
and U360 (N_360,In_711,In_900);
or U361 (N_361,In_454,In_760);
xor U362 (N_362,In_545,In_774);
and U363 (N_363,In_757,In_502);
nand U364 (N_364,In_330,In_948);
and U365 (N_365,In_102,In_202);
xor U366 (N_366,In_432,In_399);
nand U367 (N_367,In_296,In_2);
nand U368 (N_368,In_355,In_933);
nand U369 (N_369,In_66,In_186);
nand U370 (N_370,In_285,In_681);
nor U371 (N_371,In_668,In_303);
nand U372 (N_372,In_671,In_994);
or U373 (N_373,In_167,In_430);
and U374 (N_374,In_648,In_23);
or U375 (N_375,In_642,In_553);
nor U376 (N_376,In_82,In_457);
nor U377 (N_377,In_700,In_725);
nand U378 (N_378,In_656,In_194);
or U379 (N_379,In_52,In_369);
nand U380 (N_380,In_234,In_253);
xor U381 (N_381,In_451,In_494);
and U382 (N_382,In_589,In_986);
or U383 (N_383,In_846,In_446);
and U384 (N_384,In_230,In_162);
nor U385 (N_385,In_260,In_394);
nand U386 (N_386,In_282,In_365);
or U387 (N_387,In_564,In_384);
xnor U388 (N_388,In_472,In_835);
nor U389 (N_389,In_195,In_800);
or U390 (N_390,In_84,In_263);
xor U391 (N_391,In_981,In_16);
or U392 (N_392,In_537,In_214);
nor U393 (N_393,In_951,In_505);
xor U394 (N_394,In_535,In_470);
or U395 (N_395,In_400,In_187);
xnor U396 (N_396,In_94,In_348);
nor U397 (N_397,In_128,In_691);
nor U398 (N_398,In_395,In_622);
or U399 (N_399,In_831,In_584);
and U400 (N_400,In_10,In_561);
or U401 (N_401,In_996,In_362);
xor U402 (N_402,In_942,In_764);
or U403 (N_403,In_606,In_650);
or U404 (N_404,In_712,In_546);
xnor U405 (N_405,In_315,In_156);
nand U406 (N_406,In_509,In_164);
xor U407 (N_407,In_188,In_103);
nand U408 (N_408,In_619,In_741);
or U409 (N_409,In_265,In_567);
and U410 (N_410,In_661,In_250);
and U411 (N_411,In_417,In_273);
xor U412 (N_412,In_445,In_692);
nor U413 (N_413,In_702,In_777);
or U414 (N_414,In_238,In_976);
and U415 (N_415,In_69,In_902);
and U416 (N_416,In_89,In_340);
xor U417 (N_417,In_776,In_710);
or U418 (N_418,In_853,In_114);
or U419 (N_419,In_748,In_679);
nor U420 (N_420,In_768,In_827);
and U421 (N_421,In_464,In_138);
nor U422 (N_422,In_805,In_338);
nand U423 (N_423,In_4,In_595);
xnor U424 (N_424,In_378,In_145);
xnor U425 (N_425,In_316,In_404);
or U426 (N_426,In_46,In_782);
nor U427 (N_427,In_901,In_42);
nor U428 (N_428,In_63,In_139);
nand U429 (N_429,In_424,In_158);
or U430 (N_430,In_88,In_953);
nand U431 (N_431,In_977,In_873);
nand U432 (N_432,In_822,In_881);
nand U433 (N_433,In_490,In_952);
xnor U434 (N_434,In_180,In_568);
or U435 (N_435,In_497,In_684);
or U436 (N_436,In_488,In_371);
xnor U437 (N_437,In_409,In_616);
or U438 (N_438,In_603,In_110);
xor U439 (N_439,In_344,In_25);
nand U440 (N_440,In_308,In_247);
or U441 (N_441,In_15,In_428);
nand U442 (N_442,In_36,In_475);
nor U443 (N_443,In_722,In_647);
nand U444 (N_444,In_212,In_259);
or U445 (N_445,In_35,In_435);
nor U446 (N_446,In_808,In_456);
and U447 (N_447,In_331,In_18);
xor U448 (N_448,In_251,In_309);
nand U449 (N_449,In_100,In_733);
nand U450 (N_450,In_639,In_687);
and U451 (N_451,In_298,In_228);
or U452 (N_452,In_483,In_471);
or U453 (N_453,In_380,In_913);
nand U454 (N_454,In_37,In_374);
nand U455 (N_455,In_210,In_159);
and U456 (N_456,In_560,In_323);
nor U457 (N_457,In_850,In_283);
or U458 (N_458,In_750,In_864);
or U459 (N_459,In_857,In_720);
xnor U460 (N_460,In_28,In_434);
and U461 (N_461,In_660,In_797);
nand U462 (N_462,In_704,In_151);
or U463 (N_463,In_781,In_703);
or U464 (N_464,In_422,In_879);
nand U465 (N_465,In_980,In_223);
xor U466 (N_466,In_182,In_935);
nor U467 (N_467,In_304,In_439);
nand U468 (N_468,In_48,In_868);
nor U469 (N_469,In_436,In_197);
nor U470 (N_470,In_459,In_73);
nor U471 (N_471,In_886,In_884);
nor U472 (N_472,In_950,In_467);
xor U473 (N_473,In_133,In_859);
or U474 (N_474,In_983,In_593);
nand U475 (N_475,In_796,In_585);
xor U476 (N_476,In_784,In_974);
or U477 (N_477,In_79,In_740);
nor U478 (N_478,In_105,In_698);
xor U479 (N_479,In_594,In_383);
or U480 (N_480,In_761,In_357);
xor U481 (N_481,In_50,In_573);
and U482 (N_482,In_334,In_481);
and U483 (N_483,In_322,In_806);
or U484 (N_484,In_353,In_678);
nor U485 (N_485,In_185,In_780);
or U486 (N_486,In_514,In_742);
or U487 (N_487,In_888,In_427);
or U488 (N_488,In_184,In_998);
xnor U489 (N_489,In_803,In_53);
and U490 (N_490,In_160,In_217);
or U491 (N_491,In_695,In_279);
and U492 (N_492,In_149,In_613);
xor U493 (N_493,In_169,In_389);
or U494 (N_494,In_817,In_625);
and U495 (N_495,In_64,In_694);
and U496 (N_496,In_242,In_882);
and U497 (N_497,In_32,In_686);
or U498 (N_498,In_605,In_566);
nand U499 (N_499,In_543,In_515);
nand U500 (N_500,In_889,In_89);
or U501 (N_501,In_663,In_988);
nor U502 (N_502,In_50,In_686);
and U503 (N_503,In_812,In_673);
nor U504 (N_504,In_274,In_854);
or U505 (N_505,In_38,In_745);
xor U506 (N_506,In_256,In_633);
nor U507 (N_507,In_573,In_877);
nand U508 (N_508,In_194,In_535);
nor U509 (N_509,In_833,In_773);
and U510 (N_510,In_519,In_580);
xor U511 (N_511,In_622,In_880);
or U512 (N_512,In_866,In_522);
and U513 (N_513,In_612,In_930);
nand U514 (N_514,In_194,In_606);
xnor U515 (N_515,In_500,In_283);
nand U516 (N_516,In_451,In_137);
nor U517 (N_517,In_502,In_392);
nor U518 (N_518,In_856,In_451);
nor U519 (N_519,In_370,In_778);
nand U520 (N_520,In_306,In_275);
and U521 (N_521,In_345,In_37);
xnor U522 (N_522,In_970,In_774);
nand U523 (N_523,In_433,In_667);
or U524 (N_524,In_781,In_314);
xor U525 (N_525,In_885,In_719);
nand U526 (N_526,In_573,In_808);
and U527 (N_527,In_972,In_377);
and U528 (N_528,In_219,In_463);
and U529 (N_529,In_29,In_701);
nand U530 (N_530,In_114,In_794);
xor U531 (N_531,In_823,In_608);
and U532 (N_532,In_696,In_619);
nand U533 (N_533,In_407,In_766);
xor U534 (N_534,In_902,In_951);
xnor U535 (N_535,In_211,In_893);
nand U536 (N_536,In_821,In_138);
or U537 (N_537,In_705,In_747);
nand U538 (N_538,In_992,In_24);
and U539 (N_539,In_497,In_6);
nor U540 (N_540,In_28,In_368);
nor U541 (N_541,In_687,In_999);
or U542 (N_542,In_811,In_841);
nor U543 (N_543,In_961,In_894);
nand U544 (N_544,In_362,In_371);
xnor U545 (N_545,In_812,In_654);
nor U546 (N_546,In_757,In_484);
or U547 (N_547,In_325,In_737);
nor U548 (N_548,In_128,In_69);
xnor U549 (N_549,In_26,In_50);
nand U550 (N_550,In_804,In_352);
and U551 (N_551,In_506,In_631);
nor U552 (N_552,In_820,In_781);
nand U553 (N_553,In_38,In_483);
and U554 (N_554,In_744,In_416);
nand U555 (N_555,In_671,In_770);
or U556 (N_556,In_665,In_849);
and U557 (N_557,In_333,In_550);
and U558 (N_558,In_476,In_691);
nor U559 (N_559,In_415,In_765);
xnor U560 (N_560,In_698,In_774);
nand U561 (N_561,In_571,In_371);
nor U562 (N_562,In_572,In_665);
or U563 (N_563,In_154,In_211);
xor U564 (N_564,In_833,In_148);
xor U565 (N_565,In_950,In_993);
and U566 (N_566,In_665,In_550);
nand U567 (N_567,In_190,In_223);
xor U568 (N_568,In_334,In_805);
or U569 (N_569,In_974,In_710);
and U570 (N_570,In_971,In_722);
nor U571 (N_571,In_461,In_96);
or U572 (N_572,In_281,In_628);
nor U573 (N_573,In_712,In_887);
nor U574 (N_574,In_708,In_533);
and U575 (N_575,In_765,In_232);
xnor U576 (N_576,In_712,In_627);
or U577 (N_577,In_952,In_436);
and U578 (N_578,In_86,In_611);
nor U579 (N_579,In_276,In_56);
or U580 (N_580,In_383,In_325);
or U581 (N_581,In_741,In_494);
nand U582 (N_582,In_58,In_57);
and U583 (N_583,In_195,In_163);
nor U584 (N_584,In_6,In_747);
and U585 (N_585,In_964,In_840);
nand U586 (N_586,In_279,In_658);
and U587 (N_587,In_846,In_553);
nor U588 (N_588,In_854,In_448);
or U589 (N_589,In_540,In_332);
nand U590 (N_590,In_445,In_218);
nor U591 (N_591,In_388,In_564);
and U592 (N_592,In_871,In_775);
and U593 (N_593,In_684,In_252);
or U594 (N_594,In_68,In_128);
nor U595 (N_595,In_374,In_113);
nand U596 (N_596,In_51,In_0);
nand U597 (N_597,In_118,In_44);
xnor U598 (N_598,In_366,In_801);
nor U599 (N_599,In_681,In_846);
nand U600 (N_600,In_581,In_690);
and U601 (N_601,In_251,In_457);
nand U602 (N_602,In_208,In_408);
and U603 (N_603,In_426,In_795);
and U604 (N_604,In_344,In_239);
nand U605 (N_605,In_621,In_195);
and U606 (N_606,In_145,In_913);
xor U607 (N_607,In_861,In_607);
xor U608 (N_608,In_702,In_271);
xnor U609 (N_609,In_8,In_818);
xnor U610 (N_610,In_599,In_687);
nor U611 (N_611,In_12,In_247);
xor U612 (N_612,In_633,In_963);
xor U613 (N_613,In_394,In_741);
nor U614 (N_614,In_48,In_730);
and U615 (N_615,In_890,In_433);
nor U616 (N_616,In_391,In_470);
and U617 (N_617,In_516,In_676);
nor U618 (N_618,In_517,In_196);
and U619 (N_619,In_839,In_693);
xnor U620 (N_620,In_796,In_991);
nand U621 (N_621,In_415,In_33);
or U622 (N_622,In_527,In_761);
or U623 (N_623,In_967,In_776);
nand U624 (N_624,In_233,In_702);
xnor U625 (N_625,In_816,In_370);
and U626 (N_626,In_911,In_609);
nand U627 (N_627,In_734,In_920);
and U628 (N_628,In_651,In_441);
xnor U629 (N_629,In_527,In_390);
and U630 (N_630,In_708,In_828);
xnor U631 (N_631,In_491,In_632);
or U632 (N_632,In_160,In_478);
or U633 (N_633,In_883,In_663);
nor U634 (N_634,In_544,In_727);
nand U635 (N_635,In_806,In_542);
or U636 (N_636,In_725,In_969);
xnor U637 (N_637,In_976,In_191);
or U638 (N_638,In_415,In_339);
nor U639 (N_639,In_299,In_837);
nand U640 (N_640,In_96,In_493);
and U641 (N_641,In_33,In_497);
xnor U642 (N_642,In_287,In_866);
and U643 (N_643,In_164,In_132);
and U644 (N_644,In_589,In_34);
or U645 (N_645,In_793,In_254);
xnor U646 (N_646,In_255,In_708);
nor U647 (N_647,In_592,In_567);
nor U648 (N_648,In_862,In_347);
xor U649 (N_649,In_509,In_260);
nand U650 (N_650,In_214,In_295);
nor U651 (N_651,In_694,In_650);
xor U652 (N_652,In_308,In_43);
xor U653 (N_653,In_232,In_750);
and U654 (N_654,In_465,In_875);
nand U655 (N_655,In_50,In_230);
or U656 (N_656,In_426,In_397);
nor U657 (N_657,In_490,In_393);
or U658 (N_658,In_402,In_806);
nor U659 (N_659,In_585,In_446);
xnor U660 (N_660,In_88,In_741);
or U661 (N_661,In_31,In_344);
or U662 (N_662,In_259,In_115);
nand U663 (N_663,In_160,In_193);
and U664 (N_664,In_944,In_82);
nand U665 (N_665,In_271,In_261);
or U666 (N_666,In_824,In_409);
or U667 (N_667,In_715,In_181);
nand U668 (N_668,In_794,In_938);
nor U669 (N_669,In_304,In_276);
xnor U670 (N_670,In_439,In_640);
and U671 (N_671,In_113,In_389);
and U672 (N_672,In_173,In_251);
or U673 (N_673,In_44,In_460);
or U674 (N_674,In_287,In_517);
xor U675 (N_675,In_235,In_872);
nor U676 (N_676,In_208,In_713);
or U677 (N_677,In_463,In_537);
nor U678 (N_678,In_575,In_662);
xnor U679 (N_679,In_813,In_696);
nand U680 (N_680,In_15,In_844);
nor U681 (N_681,In_835,In_420);
xor U682 (N_682,In_606,In_384);
and U683 (N_683,In_836,In_307);
and U684 (N_684,In_489,In_469);
and U685 (N_685,In_536,In_201);
or U686 (N_686,In_720,In_260);
and U687 (N_687,In_998,In_558);
nand U688 (N_688,In_631,In_94);
or U689 (N_689,In_889,In_295);
xor U690 (N_690,In_729,In_928);
nand U691 (N_691,In_684,In_982);
xor U692 (N_692,In_93,In_253);
xor U693 (N_693,In_698,In_298);
nor U694 (N_694,In_503,In_739);
xnor U695 (N_695,In_679,In_766);
or U696 (N_696,In_361,In_596);
and U697 (N_697,In_211,In_964);
nand U698 (N_698,In_866,In_549);
and U699 (N_699,In_98,In_290);
xnor U700 (N_700,In_67,In_671);
xor U701 (N_701,In_338,In_799);
or U702 (N_702,In_256,In_847);
nand U703 (N_703,In_924,In_454);
and U704 (N_704,In_530,In_214);
or U705 (N_705,In_91,In_173);
nor U706 (N_706,In_51,In_510);
and U707 (N_707,In_603,In_666);
and U708 (N_708,In_845,In_164);
nor U709 (N_709,In_556,In_221);
or U710 (N_710,In_264,In_808);
nor U711 (N_711,In_742,In_472);
and U712 (N_712,In_177,In_465);
and U713 (N_713,In_881,In_889);
nor U714 (N_714,In_487,In_695);
nand U715 (N_715,In_615,In_601);
nor U716 (N_716,In_453,In_932);
xor U717 (N_717,In_239,In_381);
xnor U718 (N_718,In_865,In_99);
xnor U719 (N_719,In_765,In_598);
or U720 (N_720,In_946,In_724);
and U721 (N_721,In_382,In_141);
nand U722 (N_722,In_601,In_595);
nand U723 (N_723,In_221,In_202);
or U724 (N_724,In_27,In_991);
nand U725 (N_725,In_622,In_429);
nand U726 (N_726,In_797,In_759);
nor U727 (N_727,In_154,In_829);
or U728 (N_728,In_367,In_64);
and U729 (N_729,In_865,In_912);
nand U730 (N_730,In_234,In_79);
and U731 (N_731,In_461,In_188);
nand U732 (N_732,In_880,In_566);
and U733 (N_733,In_588,In_106);
xnor U734 (N_734,In_209,In_187);
and U735 (N_735,In_651,In_293);
or U736 (N_736,In_783,In_19);
nor U737 (N_737,In_848,In_268);
and U738 (N_738,In_800,In_260);
xnor U739 (N_739,In_438,In_469);
or U740 (N_740,In_887,In_726);
or U741 (N_741,In_659,In_336);
nand U742 (N_742,In_867,In_655);
nand U743 (N_743,In_159,In_372);
xnor U744 (N_744,In_956,In_118);
or U745 (N_745,In_970,In_675);
and U746 (N_746,In_306,In_86);
nor U747 (N_747,In_577,In_366);
xnor U748 (N_748,In_514,In_409);
xnor U749 (N_749,In_678,In_448);
nor U750 (N_750,In_572,In_902);
or U751 (N_751,In_894,In_483);
xor U752 (N_752,In_970,In_294);
or U753 (N_753,In_877,In_673);
xnor U754 (N_754,In_900,In_92);
xor U755 (N_755,In_755,In_6);
xnor U756 (N_756,In_264,In_15);
nor U757 (N_757,In_961,In_441);
nor U758 (N_758,In_917,In_800);
xnor U759 (N_759,In_514,In_903);
nor U760 (N_760,In_521,In_689);
nand U761 (N_761,In_454,In_209);
and U762 (N_762,In_415,In_422);
xor U763 (N_763,In_118,In_128);
and U764 (N_764,In_743,In_260);
nand U765 (N_765,In_436,In_144);
and U766 (N_766,In_279,In_898);
or U767 (N_767,In_130,In_547);
nand U768 (N_768,In_694,In_771);
or U769 (N_769,In_504,In_184);
or U770 (N_770,In_627,In_601);
xnor U771 (N_771,In_349,In_939);
nor U772 (N_772,In_982,In_921);
xor U773 (N_773,In_88,In_224);
nand U774 (N_774,In_992,In_787);
nor U775 (N_775,In_110,In_570);
and U776 (N_776,In_474,In_609);
nor U777 (N_777,In_337,In_370);
xor U778 (N_778,In_531,In_261);
nand U779 (N_779,In_949,In_243);
and U780 (N_780,In_918,In_248);
nor U781 (N_781,In_252,In_264);
and U782 (N_782,In_170,In_902);
and U783 (N_783,In_529,In_557);
or U784 (N_784,In_214,In_191);
xnor U785 (N_785,In_778,In_414);
nand U786 (N_786,In_304,In_399);
nor U787 (N_787,In_315,In_133);
xnor U788 (N_788,In_106,In_547);
or U789 (N_789,In_681,In_88);
or U790 (N_790,In_797,In_0);
xor U791 (N_791,In_244,In_993);
nor U792 (N_792,In_418,In_172);
xnor U793 (N_793,In_24,In_232);
xor U794 (N_794,In_75,In_558);
nand U795 (N_795,In_132,In_778);
xor U796 (N_796,In_866,In_887);
nor U797 (N_797,In_549,In_153);
xnor U798 (N_798,In_514,In_95);
nor U799 (N_799,In_865,In_485);
or U800 (N_800,In_873,In_635);
nor U801 (N_801,In_943,In_942);
xnor U802 (N_802,In_610,In_243);
and U803 (N_803,In_257,In_296);
and U804 (N_804,In_955,In_770);
or U805 (N_805,In_694,In_71);
or U806 (N_806,In_51,In_687);
and U807 (N_807,In_608,In_876);
and U808 (N_808,In_548,In_136);
nand U809 (N_809,In_509,In_630);
or U810 (N_810,In_518,In_324);
or U811 (N_811,In_570,In_5);
nand U812 (N_812,In_89,In_608);
nand U813 (N_813,In_724,In_871);
or U814 (N_814,In_387,In_490);
xor U815 (N_815,In_237,In_640);
or U816 (N_816,In_685,In_462);
xnor U817 (N_817,In_286,In_100);
or U818 (N_818,In_908,In_887);
or U819 (N_819,In_726,In_947);
and U820 (N_820,In_659,In_500);
and U821 (N_821,In_795,In_535);
nand U822 (N_822,In_58,In_427);
xor U823 (N_823,In_159,In_628);
nand U824 (N_824,In_407,In_90);
nor U825 (N_825,In_235,In_198);
nor U826 (N_826,In_62,In_833);
nand U827 (N_827,In_355,In_776);
or U828 (N_828,In_407,In_192);
or U829 (N_829,In_374,In_121);
nand U830 (N_830,In_579,In_138);
xor U831 (N_831,In_503,In_293);
nor U832 (N_832,In_271,In_818);
or U833 (N_833,In_336,In_392);
or U834 (N_834,In_125,In_450);
xor U835 (N_835,In_72,In_934);
or U836 (N_836,In_306,In_24);
xor U837 (N_837,In_224,In_728);
xnor U838 (N_838,In_293,In_484);
nand U839 (N_839,In_231,In_62);
or U840 (N_840,In_8,In_85);
nand U841 (N_841,In_795,In_105);
or U842 (N_842,In_369,In_443);
xor U843 (N_843,In_661,In_802);
xnor U844 (N_844,In_606,In_802);
and U845 (N_845,In_19,In_797);
nand U846 (N_846,In_651,In_570);
and U847 (N_847,In_953,In_236);
xor U848 (N_848,In_181,In_253);
and U849 (N_849,In_449,In_296);
or U850 (N_850,In_243,In_356);
nor U851 (N_851,In_231,In_744);
nand U852 (N_852,In_100,In_517);
nand U853 (N_853,In_133,In_613);
or U854 (N_854,In_274,In_410);
or U855 (N_855,In_260,In_144);
and U856 (N_856,In_264,In_920);
xnor U857 (N_857,In_119,In_980);
nor U858 (N_858,In_116,In_119);
and U859 (N_859,In_231,In_805);
nor U860 (N_860,In_838,In_144);
xor U861 (N_861,In_45,In_98);
nand U862 (N_862,In_598,In_621);
and U863 (N_863,In_103,In_1);
nor U864 (N_864,In_233,In_318);
nand U865 (N_865,In_43,In_413);
or U866 (N_866,In_982,In_351);
xor U867 (N_867,In_83,In_668);
nor U868 (N_868,In_780,In_978);
nand U869 (N_869,In_448,In_731);
or U870 (N_870,In_256,In_400);
nor U871 (N_871,In_826,In_18);
nand U872 (N_872,In_442,In_126);
or U873 (N_873,In_193,In_547);
nand U874 (N_874,In_54,In_70);
or U875 (N_875,In_401,In_422);
xor U876 (N_876,In_503,In_613);
or U877 (N_877,In_314,In_665);
nor U878 (N_878,In_555,In_435);
nor U879 (N_879,In_791,In_935);
or U880 (N_880,In_595,In_46);
nand U881 (N_881,In_737,In_766);
nor U882 (N_882,In_942,In_886);
nor U883 (N_883,In_572,In_414);
and U884 (N_884,In_663,In_751);
xor U885 (N_885,In_336,In_431);
nor U886 (N_886,In_640,In_723);
nor U887 (N_887,In_945,In_972);
nand U888 (N_888,In_168,In_398);
nor U889 (N_889,In_793,In_918);
and U890 (N_890,In_983,In_943);
nor U891 (N_891,In_674,In_837);
or U892 (N_892,In_60,In_186);
xnor U893 (N_893,In_966,In_499);
nor U894 (N_894,In_279,In_110);
or U895 (N_895,In_597,In_546);
xnor U896 (N_896,In_297,In_712);
xor U897 (N_897,In_790,In_967);
and U898 (N_898,In_984,In_506);
nand U899 (N_899,In_636,In_707);
xor U900 (N_900,In_258,In_547);
nor U901 (N_901,In_103,In_536);
nand U902 (N_902,In_442,In_554);
or U903 (N_903,In_497,In_555);
nand U904 (N_904,In_274,In_218);
and U905 (N_905,In_177,In_307);
xor U906 (N_906,In_28,In_77);
nor U907 (N_907,In_697,In_190);
or U908 (N_908,In_556,In_291);
nand U909 (N_909,In_104,In_768);
nor U910 (N_910,In_460,In_134);
nor U911 (N_911,In_217,In_966);
nor U912 (N_912,In_644,In_169);
or U913 (N_913,In_643,In_410);
xnor U914 (N_914,In_495,In_343);
or U915 (N_915,In_38,In_217);
or U916 (N_916,In_240,In_793);
nand U917 (N_917,In_891,In_248);
nand U918 (N_918,In_653,In_890);
nand U919 (N_919,In_782,In_512);
and U920 (N_920,In_518,In_457);
nor U921 (N_921,In_441,In_785);
nor U922 (N_922,In_487,In_269);
xor U923 (N_923,In_420,In_643);
nor U924 (N_924,In_215,In_84);
xnor U925 (N_925,In_948,In_276);
xnor U926 (N_926,In_802,In_524);
nor U927 (N_927,In_141,In_356);
and U928 (N_928,In_941,In_870);
and U929 (N_929,In_968,In_22);
nand U930 (N_930,In_314,In_985);
nand U931 (N_931,In_886,In_283);
nor U932 (N_932,In_339,In_337);
xor U933 (N_933,In_827,In_776);
and U934 (N_934,In_869,In_0);
nor U935 (N_935,In_572,In_875);
or U936 (N_936,In_97,In_206);
and U937 (N_937,In_316,In_617);
or U938 (N_938,In_201,In_727);
and U939 (N_939,In_775,In_95);
nand U940 (N_940,In_66,In_403);
or U941 (N_941,In_30,In_303);
nand U942 (N_942,In_714,In_879);
or U943 (N_943,In_87,In_844);
nand U944 (N_944,In_49,In_44);
nor U945 (N_945,In_849,In_540);
nand U946 (N_946,In_372,In_530);
nand U947 (N_947,In_607,In_424);
nor U948 (N_948,In_593,In_406);
and U949 (N_949,In_189,In_697);
nand U950 (N_950,In_819,In_378);
and U951 (N_951,In_404,In_488);
xor U952 (N_952,In_257,In_43);
nor U953 (N_953,In_237,In_510);
xnor U954 (N_954,In_325,In_579);
nor U955 (N_955,In_797,In_365);
and U956 (N_956,In_235,In_584);
or U957 (N_957,In_524,In_760);
nor U958 (N_958,In_23,In_714);
nand U959 (N_959,In_693,In_44);
xor U960 (N_960,In_109,In_954);
nand U961 (N_961,In_594,In_294);
and U962 (N_962,In_424,In_984);
xor U963 (N_963,In_233,In_140);
nand U964 (N_964,In_625,In_623);
nor U965 (N_965,In_153,In_203);
xnor U966 (N_966,In_165,In_183);
or U967 (N_967,In_382,In_299);
or U968 (N_968,In_547,In_926);
nand U969 (N_969,In_200,In_831);
or U970 (N_970,In_716,In_431);
xor U971 (N_971,In_898,In_511);
and U972 (N_972,In_611,In_223);
xnor U973 (N_973,In_415,In_961);
nor U974 (N_974,In_496,In_347);
nor U975 (N_975,In_806,In_844);
xor U976 (N_976,In_534,In_941);
nor U977 (N_977,In_63,In_730);
or U978 (N_978,In_321,In_271);
nor U979 (N_979,In_322,In_353);
nor U980 (N_980,In_487,In_536);
xnor U981 (N_981,In_513,In_542);
or U982 (N_982,In_269,In_271);
nand U983 (N_983,In_221,In_273);
and U984 (N_984,In_143,In_549);
xor U985 (N_985,In_314,In_315);
or U986 (N_986,In_296,In_840);
or U987 (N_987,In_658,In_900);
or U988 (N_988,In_211,In_749);
nand U989 (N_989,In_592,In_533);
nor U990 (N_990,In_752,In_385);
xnor U991 (N_991,In_407,In_517);
nand U992 (N_992,In_686,In_777);
nand U993 (N_993,In_168,In_799);
nor U994 (N_994,In_457,In_137);
nand U995 (N_995,In_881,In_972);
nor U996 (N_996,In_975,In_850);
nand U997 (N_997,In_827,In_294);
nand U998 (N_998,In_702,In_285);
nor U999 (N_999,In_577,In_131);
xor U1000 (N_1000,N_984,N_634);
and U1001 (N_1001,N_346,N_792);
nor U1002 (N_1002,N_130,N_712);
or U1003 (N_1003,N_994,N_217);
xnor U1004 (N_1004,N_100,N_564);
xnor U1005 (N_1005,N_832,N_575);
nand U1006 (N_1006,N_589,N_967);
nand U1007 (N_1007,N_696,N_656);
xor U1008 (N_1008,N_170,N_443);
or U1009 (N_1009,N_401,N_242);
and U1010 (N_1010,N_464,N_509);
and U1011 (N_1011,N_680,N_688);
or U1012 (N_1012,N_337,N_156);
nand U1013 (N_1013,N_183,N_639);
or U1014 (N_1014,N_459,N_442);
nor U1015 (N_1015,N_216,N_798);
or U1016 (N_1016,N_79,N_512);
nor U1017 (N_1017,N_264,N_610);
or U1018 (N_1018,N_387,N_775);
nand U1019 (N_1019,N_43,N_434);
or U1020 (N_1020,N_840,N_996);
and U1021 (N_1021,N_326,N_966);
nor U1022 (N_1022,N_621,N_578);
and U1023 (N_1023,N_152,N_882);
and U1024 (N_1024,N_803,N_470);
nor U1025 (N_1025,N_647,N_222);
and U1026 (N_1026,N_486,N_674);
and U1027 (N_1027,N_925,N_403);
xnor U1028 (N_1028,N_192,N_899);
nor U1029 (N_1029,N_884,N_672);
and U1030 (N_1030,N_394,N_953);
or U1031 (N_1031,N_576,N_719);
nor U1032 (N_1032,N_502,N_633);
and U1033 (N_1033,N_200,N_123);
nor U1034 (N_1034,N_777,N_67);
nor U1035 (N_1035,N_587,N_377);
nor U1036 (N_1036,N_223,N_140);
xnor U1037 (N_1037,N_157,N_51);
or U1038 (N_1038,N_344,N_530);
and U1039 (N_1039,N_112,N_56);
xor U1040 (N_1040,N_304,N_641);
nor U1041 (N_1041,N_848,N_262);
and U1042 (N_1042,N_661,N_833);
xor U1043 (N_1043,N_109,N_684);
or U1044 (N_1044,N_824,N_513);
nor U1045 (N_1045,N_335,N_700);
xnor U1046 (N_1046,N_711,N_350);
nand U1047 (N_1047,N_26,N_16);
or U1048 (N_1048,N_707,N_323);
xnor U1049 (N_1049,N_59,N_106);
and U1050 (N_1050,N_36,N_131);
nand U1051 (N_1051,N_797,N_664);
nor U1052 (N_1052,N_506,N_355);
xnor U1053 (N_1053,N_504,N_657);
or U1054 (N_1054,N_806,N_354);
or U1055 (N_1055,N_207,N_336);
or U1056 (N_1056,N_312,N_908);
nor U1057 (N_1057,N_245,N_5);
or U1058 (N_1058,N_975,N_616);
and U1059 (N_1059,N_545,N_758);
nor U1060 (N_1060,N_97,N_760);
or U1061 (N_1061,N_776,N_930);
xnor U1062 (N_1062,N_801,N_821);
nand U1063 (N_1063,N_72,N_944);
and U1064 (N_1064,N_116,N_698);
nand U1065 (N_1065,N_198,N_46);
xnor U1066 (N_1066,N_255,N_583);
or U1067 (N_1067,N_640,N_121);
xor U1068 (N_1068,N_615,N_514);
and U1069 (N_1069,N_3,N_98);
nor U1070 (N_1070,N_909,N_7);
xor U1071 (N_1071,N_400,N_722);
or U1072 (N_1072,N_381,N_324);
or U1073 (N_1073,N_503,N_710);
nand U1074 (N_1074,N_208,N_148);
and U1075 (N_1075,N_213,N_817);
or U1076 (N_1076,N_297,N_340);
nand U1077 (N_1077,N_667,N_359);
xnor U1078 (N_1078,N_463,N_628);
xnor U1079 (N_1079,N_706,N_124);
nor U1080 (N_1080,N_126,N_597);
and U1081 (N_1081,N_37,N_224);
and U1082 (N_1082,N_138,N_870);
nand U1083 (N_1083,N_220,N_643);
nand U1084 (N_1084,N_972,N_168);
nand U1085 (N_1085,N_412,N_648);
nor U1086 (N_1086,N_181,N_869);
nand U1087 (N_1087,N_609,N_416);
nor U1088 (N_1088,N_982,N_219);
and U1089 (N_1089,N_0,N_136);
xnor U1090 (N_1090,N_475,N_890);
or U1091 (N_1091,N_21,N_726);
and U1092 (N_1092,N_270,N_291);
xnor U1093 (N_1093,N_493,N_604);
or U1094 (N_1094,N_283,N_841);
nand U1095 (N_1095,N_686,N_250);
or U1096 (N_1096,N_742,N_831);
xnor U1097 (N_1097,N_339,N_511);
or U1098 (N_1098,N_483,N_497);
nor U1099 (N_1099,N_836,N_741);
xnor U1100 (N_1100,N_665,N_863);
nor U1101 (N_1101,N_693,N_215);
nor U1102 (N_1102,N_781,N_997);
and U1103 (N_1103,N_613,N_101);
xnor U1104 (N_1104,N_602,N_888);
xnor U1105 (N_1105,N_375,N_286);
nor U1106 (N_1106,N_714,N_951);
or U1107 (N_1107,N_795,N_364);
nor U1108 (N_1108,N_800,N_537);
nor U1109 (N_1109,N_857,N_135);
xnor U1110 (N_1110,N_622,N_662);
or U1111 (N_1111,N_744,N_763);
and U1112 (N_1112,N_63,N_757);
nand U1113 (N_1113,N_180,N_977);
nor U1114 (N_1114,N_269,N_980);
xnor U1115 (N_1115,N_808,N_432);
xor U1116 (N_1116,N_425,N_499);
and U1117 (N_1117,N_729,N_179);
nand U1118 (N_1118,N_391,N_654);
nor U1119 (N_1119,N_60,N_382);
nor U1120 (N_1120,N_221,N_469);
nand U1121 (N_1121,N_644,N_64);
and U1122 (N_1122,N_747,N_592);
or U1123 (N_1123,N_68,N_995);
nor U1124 (N_1124,N_663,N_551);
xor U1125 (N_1125,N_823,N_19);
or U1126 (N_1126,N_931,N_186);
nor U1127 (N_1127,N_93,N_30);
nand U1128 (N_1128,N_118,N_778);
nand U1129 (N_1129,N_73,N_393);
xnor U1130 (N_1130,N_174,N_708);
xnor U1131 (N_1131,N_251,N_531);
or U1132 (N_1132,N_471,N_331);
xnor U1133 (N_1133,N_791,N_383);
nor U1134 (N_1134,N_399,N_13);
and U1135 (N_1135,N_415,N_92);
nor U1136 (N_1136,N_133,N_86);
nor U1137 (N_1137,N_411,N_128);
and U1138 (N_1138,N_683,N_709);
or U1139 (N_1139,N_608,N_164);
xnor U1140 (N_1140,N_84,N_827);
nand U1141 (N_1141,N_548,N_958);
nand U1142 (N_1142,N_986,N_992);
or U1143 (N_1143,N_182,N_178);
or U1144 (N_1144,N_750,N_771);
nand U1145 (N_1145,N_756,N_856);
xnor U1146 (N_1146,N_449,N_723);
or U1147 (N_1147,N_435,N_272);
or U1148 (N_1148,N_906,N_161);
or U1149 (N_1149,N_851,N_745);
and U1150 (N_1150,N_48,N_41);
xor U1151 (N_1151,N_11,N_993);
nand U1152 (N_1152,N_860,N_488);
or U1153 (N_1153,N_322,N_99);
and U1154 (N_1154,N_386,N_636);
or U1155 (N_1155,N_102,N_185);
nand U1156 (N_1156,N_838,N_959);
nor U1157 (N_1157,N_27,N_642);
and U1158 (N_1158,N_839,N_85);
xor U1159 (N_1159,N_794,N_914);
xnor U1160 (N_1160,N_158,N_507);
nand U1161 (N_1161,N_211,N_38);
nor U1162 (N_1162,N_120,N_630);
and U1163 (N_1163,N_385,N_467);
nand U1164 (N_1164,N_34,N_873);
or U1165 (N_1165,N_414,N_457);
nor U1166 (N_1166,N_897,N_834);
nor U1167 (N_1167,N_976,N_704);
or U1168 (N_1168,N_881,N_47);
and U1169 (N_1169,N_886,N_751);
or U1170 (N_1170,N_292,N_594);
and U1171 (N_1171,N_482,N_302);
and U1172 (N_1172,N_74,N_214);
nand U1173 (N_1173,N_490,N_405);
and U1174 (N_1174,N_212,N_903);
nand U1175 (N_1175,N_713,N_61);
or U1176 (N_1176,N_562,N_22);
xor U1177 (N_1177,N_352,N_934);
xnor U1178 (N_1178,N_943,N_620);
or U1179 (N_1179,N_572,N_783);
and U1180 (N_1180,N_240,N_521);
nor U1181 (N_1181,N_969,N_259);
xor U1182 (N_1182,N_445,N_261);
or U1183 (N_1183,N_252,N_165);
nor U1184 (N_1184,N_32,N_404);
nor U1185 (N_1185,N_24,N_308);
nor U1186 (N_1186,N_735,N_885);
or U1187 (N_1187,N_388,N_438);
nand U1188 (N_1188,N_44,N_358);
nand U1189 (N_1189,N_968,N_962);
and U1190 (N_1190,N_299,N_600);
or U1191 (N_1191,N_188,N_727);
nor U1192 (N_1192,N_289,N_205);
and U1193 (N_1193,N_380,N_96);
or U1194 (N_1194,N_139,N_901);
nand U1195 (N_1195,N_671,N_916);
nand U1196 (N_1196,N_522,N_111);
or U1197 (N_1197,N_384,N_920);
nand U1198 (N_1198,N_424,N_366);
or U1199 (N_1199,N_544,N_867);
or U1200 (N_1200,N_847,N_612);
xnor U1201 (N_1201,N_108,N_586);
xnor U1202 (N_1202,N_618,N_941);
nor U1203 (N_1203,N_721,N_942);
nor U1204 (N_1204,N_496,N_309);
nand U1205 (N_1205,N_439,N_787);
nor U1206 (N_1206,N_50,N_703);
or U1207 (N_1207,N_281,N_447);
nand U1208 (N_1208,N_12,N_517);
nand U1209 (N_1209,N_25,N_45);
nand U1210 (N_1210,N_154,N_638);
xnor U1211 (N_1211,N_601,N_440);
xnor U1212 (N_1212,N_317,N_9);
nand U1213 (N_1213,N_278,N_103);
nand U1214 (N_1214,N_265,N_476);
and U1215 (N_1215,N_441,N_244);
xor U1216 (N_1216,N_534,N_598);
xor U1217 (N_1217,N_753,N_226);
and U1218 (N_1218,N_546,N_955);
and U1219 (N_1219,N_311,N_117);
or U1220 (N_1220,N_973,N_631);
xnor U1221 (N_1221,N_614,N_347);
xor U1222 (N_1222,N_320,N_949);
and U1223 (N_1223,N_859,N_957);
and U1224 (N_1224,N_49,N_861);
nor U1225 (N_1225,N_591,N_162);
and U1226 (N_1226,N_367,N_649);
and U1227 (N_1227,N_327,N_66);
or U1228 (N_1228,N_846,N_538);
and U1229 (N_1229,N_623,N_501);
nor U1230 (N_1230,N_396,N_6);
or U1231 (N_1231,N_720,N_65);
or U1232 (N_1232,N_237,N_176);
nand U1233 (N_1233,N_734,N_875);
and U1234 (N_1234,N_369,N_257);
xor U1235 (N_1235,N_189,N_256);
or U1236 (N_1236,N_236,N_451);
and U1237 (N_1237,N_985,N_845);
nor U1238 (N_1238,N_754,N_738);
nor U1239 (N_1239,N_844,N_670);
or U1240 (N_1240,N_933,N_351);
xnor U1241 (N_1241,N_809,N_596);
xor U1242 (N_1242,N_605,N_196);
nand U1243 (N_1243,N_807,N_632);
and U1244 (N_1244,N_516,N_202);
nand U1245 (N_1245,N_762,N_853);
or U1246 (N_1246,N_107,N_915);
xor U1247 (N_1247,N_390,N_990);
or U1248 (N_1248,N_611,N_149);
nand U1249 (N_1249,N_487,N_203);
nor U1250 (N_1250,N_987,N_62);
nor U1251 (N_1251,N_782,N_767);
and U1252 (N_1252,N_498,N_479);
and U1253 (N_1253,N_816,N_728);
xnor U1254 (N_1254,N_260,N_279);
nor U1255 (N_1255,N_417,N_82);
xnor U1256 (N_1256,N_235,N_166);
and U1257 (N_1257,N_550,N_389);
nand U1258 (N_1258,N_91,N_129);
nand U1259 (N_1259,N_519,N_779);
nand U1260 (N_1260,N_746,N_796);
and U1261 (N_1261,N_280,N_561);
nand U1262 (N_1262,N_132,N_360);
and U1263 (N_1263,N_76,N_733);
nand U1264 (N_1264,N_150,N_828);
nor U1265 (N_1265,N_898,N_716);
nand U1266 (N_1266,N_134,N_419);
nand U1267 (N_1267,N_685,N_454);
xor U1268 (N_1268,N_105,N_427);
nor U1269 (N_1269,N_81,N_887);
xor U1270 (N_1270,N_558,N_141);
xor U1271 (N_1271,N_790,N_268);
nand U1272 (N_1272,N_876,N_406);
xnor U1273 (N_1273,N_617,N_749);
or U1274 (N_1274,N_811,N_936);
xnor U1275 (N_1275,N_55,N_374);
xnor U1276 (N_1276,N_581,N_568);
or U1277 (N_1277,N_619,N_330);
and U1278 (N_1278,N_912,N_536);
nand U1279 (N_1279,N_878,N_625);
and U1280 (N_1280,N_159,N_338);
xnor U1281 (N_1281,N_199,N_288);
xnor U1282 (N_1282,N_563,N_655);
or U1283 (N_1283,N_231,N_33);
and U1284 (N_1284,N_379,N_18);
nand U1285 (N_1285,N_239,N_892);
or U1286 (N_1286,N_145,N_542);
nand U1287 (N_1287,N_195,N_349);
and U1288 (N_1288,N_812,N_83);
nand U1289 (N_1289,N_879,N_209);
and U1290 (N_1290,N_724,N_458);
xor U1291 (N_1291,N_784,N_277);
or U1292 (N_1292,N_554,N_306);
nor U1293 (N_1293,N_42,N_789);
xor U1294 (N_1294,N_225,N_919);
nor U1295 (N_1295,N_187,N_820);
nand U1296 (N_1296,N_325,N_14);
xnor U1297 (N_1297,N_436,N_478);
xor U1298 (N_1298,N_263,N_314);
xor U1299 (N_1299,N_201,N_410);
or U1300 (N_1300,N_902,N_319);
or U1301 (N_1301,N_510,N_880);
xnor U1302 (N_1302,N_210,N_691);
nand U1303 (N_1303,N_635,N_173);
or U1304 (N_1304,N_917,N_296);
nand U1305 (N_1305,N_167,N_547);
or U1306 (N_1306,N_271,N_448);
or U1307 (N_1307,N_8,N_193);
xor U1308 (N_1308,N_249,N_543);
xor U1309 (N_1309,N_10,N_426);
nand U1310 (N_1310,N_155,N_151);
and U1311 (N_1311,N_570,N_153);
or U1312 (N_1312,N_541,N_190);
nor U1313 (N_1313,N_491,N_333);
nand U1314 (N_1314,N_921,N_893);
nor U1315 (N_1315,N_392,N_343);
xnor U1316 (N_1316,N_692,N_669);
and U1317 (N_1317,N_194,N_368);
and U1318 (N_1318,N_956,N_793);
nor U1319 (N_1319,N_687,N_705);
and U1320 (N_1320,N_465,N_298);
or U1321 (N_1321,N_730,N_676);
and U1322 (N_1322,N_287,N_577);
and U1323 (N_1323,N_370,N_765);
xor U1324 (N_1324,N_922,N_20);
and U1325 (N_1325,N_874,N_926);
nor U1326 (N_1326,N_739,N_571);
nand U1327 (N_1327,N_549,N_492);
nor U1328 (N_1328,N_595,N_815);
and U1329 (N_1329,N_865,N_755);
and U1330 (N_1330,N_918,N_275);
nor U1331 (N_1331,N_533,N_829);
nand U1332 (N_1332,N_57,N_764);
nand U1333 (N_1333,N_864,N_518);
nand U1334 (N_1334,N_715,N_247);
nor U1335 (N_1335,N_946,N_660);
nor U1336 (N_1336,N_607,N_206);
xnor U1337 (N_1337,N_637,N_998);
or U1338 (N_1338,N_31,N_842);
or U1339 (N_1339,N_588,N_446);
nor U1340 (N_1340,N_629,N_243);
and U1341 (N_1341,N_357,N_71);
nor U1342 (N_1342,N_160,N_565);
nand U1343 (N_1343,N_110,N_835);
and U1344 (N_1344,N_850,N_307);
or U1345 (N_1345,N_456,N_485);
xnor U1346 (N_1346,N_673,N_474);
nor U1347 (N_1347,N_520,N_295);
nand U1348 (N_1348,N_163,N_814);
xor U1349 (N_1349,N_768,N_114);
xnor U1350 (N_1350,N_29,N_653);
and U1351 (N_1351,N_54,N_408);
nand U1352 (N_1352,N_938,N_785);
nor U1353 (N_1353,N_172,N_627);
xnor U1354 (N_1354,N_378,N_737);
and U1355 (N_1355,N_87,N_274);
xnor U1356 (N_1356,N_332,N_780);
xor U1357 (N_1357,N_39,N_462);
or U1358 (N_1358,N_489,N_119);
nand U1359 (N_1359,N_500,N_896);
xor U1360 (N_1360,N_895,N_774);
nor U1361 (N_1361,N_675,N_238);
or U1362 (N_1362,N_4,N_80);
and U1363 (N_1363,N_788,N_70);
nand U1364 (N_1364,N_313,N_645);
nor U1365 (N_1365,N_695,N_566);
and U1366 (N_1366,N_862,N_1);
nand U1367 (N_1367,N_528,N_58);
and U1368 (N_1368,N_227,N_285);
and U1369 (N_1369,N_363,N_413);
nand U1370 (N_1370,N_420,N_246);
or U1371 (N_1371,N_127,N_699);
nor U1372 (N_1372,N_843,N_697);
or U1373 (N_1373,N_689,N_197);
nor U1374 (N_1374,N_428,N_477);
xnor U1375 (N_1375,N_433,N_813);
xor U1376 (N_1376,N_293,N_871);
or U1377 (N_1377,N_593,N_567);
and U1378 (N_1378,N_254,N_316);
nor U1379 (N_1379,N_321,N_125);
nor U1380 (N_1380,N_361,N_267);
or U1381 (N_1381,N_574,N_849);
xnor U1382 (N_1382,N_988,N_983);
xor U1383 (N_1383,N_342,N_113);
nor U1384 (N_1384,N_15,N_725);
and U1385 (N_1385,N_104,N_822);
nand U1386 (N_1386,N_52,N_266);
or U1387 (N_1387,N_95,N_184);
or U1388 (N_1388,N_830,N_866);
xor U1389 (N_1389,N_455,N_523);
nor U1390 (N_1390,N_234,N_229);
and U1391 (N_1391,N_772,N_315);
xor U1392 (N_1392,N_329,N_947);
and U1393 (N_1393,N_253,N_395);
xor U1394 (N_1394,N_883,N_872);
nor U1395 (N_1395,N_981,N_868);
and U1396 (N_1396,N_484,N_603);
or U1397 (N_1397,N_472,N_175);
and U1398 (N_1398,N_17,N_819);
xnor U1399 (N_1399,N_556,N_35);
xor U1400 (N_1400,N_748,N_171);
nand U1401 (N_1401,N_328,N_854);
xnor U1402 (N_1402,N_423,N_89);
nor U1403 (N_1403,N_891,N_461);
nand U1404 (N_1404,N_28,N_144);
and U1405 (N_1405,N_964,N_553);
nand U1406 (N_1406,N_804,N_421);
and U1407 (N_1407,N_569,N_429);
xor U1408 (N_1408,N_948,N_204);
or U1409 (N_1409,N_539,N_241);
and U1410 (N_1410,N_23,N_904);
xnor U1411 (N_1411,N_950,N_143);
xor U1412 (N_1412,N_353,N_2);
nor U1413 (N_1413,N_646,N_590);
nand U1414 (N_1414,N_481,N_422);
xor U1415 (N_1415,N_362,N_230);
or U1416 (N_1416,N_532,N_529);
and U1417 (N_1417,N_233,N_137);
nor U1418 (N_1418,N_651,N_398);
xnor U1419 (N_1419,N_606,N_894);
nand U1420 (N_1420,N_960,N_802);
xor U1421 (N_1421,N_770,N_923);
xnor U1422 (N_1422,N_584,N_90);
and U1423 (N_1423,N_122,N_855);
xnor U1424 (N_1424,N_626,N_284);
and U1425 (N_1425,N_397,N_371);
or U1426 (N_1426,N_345,N_248);
nand U1427 (N_1427,N_557,N_177);
and U1428 (N_1428,N_954,N_701);
and U1429 (N_1429,N_495,N_524);
xor U1430 (N_1430,N_658,N_69);
nand U1431 (N_1431,N_147,N_668);
or U1432 (N_1432,N_971,N_468);
xor U1433 (N_1433,N_852,N_560);
nor U1434 (N_1434,N_305,N_142);
or U1435 (N_1435,N_818,N_978);
xor U1436 (N_1436,N_961,N_678);
nor U1437 (N_1437,N_407,N_718);
xnor U1438 (N_1438,N_766,N_535);
nand U1439 (N_1439,N_473,N_582);
and U1440 (N_1440,N_907,N_540);
nor U1441 (N_1441,N_232,N_515);
or U1442 (N_1442,N_505,N_555);
or U1443 (N_1443,N_945,N_965);
and U1444 (N_1444,N_258,N_939);
nand U1445 (N_1445,N_282,N_430);
or U1446 (N_1446,N_679,N_759);
and U1447 (N_1447,N_940,N_373);
and U1448 (N_1448,N_273,N_666);
and U1449 (N_1449,N_999,N_677);
nor U1450 (N_1450,N_702,N_905);
xor U1451 (N_1451,N_480,N_743);
or U1452 (N_1452,N_334,N_372);
or U1453 (N_1453,N_889,N_526);
or U1454 (N_1454,N_228,N_952);
xor U1455 (N_1455,N_301,N_752);
and U1456 (N_1456,N_431,N_78);
or U1457 (N_1457,N_979,N_731);
or U1458 (N_1458,N_928,N_88);
xor U1459 (N_1459,N_682,N_573);
nor U1460 (N_1460,N_732,N_376);
xnor U1461 (N_1461,N_659,N_75);
or U1462 (N_1462,N_310,N_690);
nor U1463 (N_1463,N_911,N_927);
nand U1464 (N_1464,N_935,N_694);
nand U1465 (N_1465,N_599,N_508);
or U1466 (N_1466,N_466,N_169);
and U1467 (N_1467,N_810,N_527);
xnor U1468 (N_1468,N_799,N_991);
or U1469 (N_1469,N_769,N_494);
or U1470 (N_1470,N_318,N_453);
nor U1471 (N_1471,N_218,N_624);
and U1472 (N_1472,N_525,N_826);
or U1473 (N_1473,N_303,N_437);
nand U1474 (N_1474,N_740,N_356);
or U1475 (N_1475,N_452,N_409);
xnor U1476 (N_1476,N_579,N_932);
xor U1477 (N_1477,N_937,N_418);
xnor U1478 (N_1478,N_650,N_858);
nor U1479 (N_1479,N_40,N_348);
and U1480 (N_1480,N_929,N_460);
xor U1481 (N_1481,N_94,N_963);
and U1482 (N_1482,N_341,N_191);
nor U1483 (N_1483,N_717,N_53);
xnor U1484 (N_1484,N_294,N_146);
xor U1485 (N_1485,N_585,N_773);
and U1486 (N_1486,N_974,N_900);
xnor U1487 (N_1487,N_681,N_444);
and U1488 (N_1488,N_805,N_115);
or U1489 (N_1489,N_989,N_877);
and U1490 (N_1490,N_786,N_276);
or U1491 (N_1491,N_652,N_300);
nand U1492 (N_1492,N_761,N_450);
or U1493 (N_1493,N_924,N_290);
xnor U1494 (N_1494,N_559,N_910);
nand U1495 (N_1495,N_825,N_837);
nand U1496 (N_1496,N_736,N_552);
xnor U1497 (N_1497,N_365,N_580);
xor U1498 (N_1498,N_913,N_970);
nand U1499 (N_1499,N_77,N_402);
or U1500 (N_1500,N_480,N_56);
xor U1501 (N_1501,N_235,N_188);
xnor U1502 (N_1502,N_339,N_110);
or U1503 (N_1503,N_95,N_974);
nand U1504 (N_1504,N_978,N_253);
or U1505 (N_1505,N_939,N_414);
nand U1506 (N_1506,N_119,N_878);
nand U1507 (N_1507,N_961,N_111);
nor U1508 (N_1508,N_12,N_334);
and U1509 (N_1509,N_697,N_58);
xor U1510 (N_1510,N_688,N_239);
xor U1511 (N_1511,N_156,N_245);
and U1512 (N_1512,N_484,N_400);
nor U1513 (N_1513,N_31,N_796);
nand U1514 (N_1514,N_410,N_406);
and U1515 (N_1515,N_83,N_214);
xor U1516 (N_1516,N_430,N_971);
xnor U1517 (N_1517,N_888,N_367);
xor U1518 (N_1518,N_696,N_712);
nand U1519 (N_1519,N_57,N_236);
and U1520 (N_1520,N_897,N_750);
xor U1521 (N_1521,N_759,N_650);
nand U1522 (N_1522,N_264,N_619);
and U1523 (N_1523,N_797,N_340);
nor U1524 (N_1524,N_322,N_791);
or U1525 (N_1525,N_749,N_969);
or U1526 (N_1526,N_818,N_870);
nand U1527 (N_1527,N_789,N_507);
nor U1528 (N_1528,N_355,N_572);
nand U1529 (N_1529,N_763,N_946);
or U1530 (N_1530,N_136,N_253);
xor U1531 (N_1531,N_629,N_411);
nor U1532 (N_1532,N_819,N_493);
nor U1533 (N_1533,N_102,N_163);
and U1534 (N_1534,N_740,N_102);
xnor U1535 (N_1535,N_512,N_101);
nor U1536 (N_1536,N_366,N_801);
nor U1537 (N_1537,N_461,N_362);
and U1538 (N_1538,N_290,N_582);
nand U1539 (N_1539,N_236,N_282);
xnor U1540 (N_1540,N_844,N_948);
and U1541 (N_1541,N_880,N_198);
xor U1542 (N_1542,N_495,N_465);
nor U1543 (N_1543,N_210,N_826);
and U1544 (N_1544,N_340,N_757);
xor U1545 (N_1545,N_820,N_390);
nand U1546 (N_1546,N_846,N_845);
nor U1547 (N_1547,N_933,N_724);
nand U1548 (N_1548,N_327,N_359);
nor U1549 (N_1549,N_398,N_865);
or U1550 (N_1550,N_446,N_944);
or U1551 (N_1551,N_425,N_144);
nand U1552 (N_1552,N_826,N_492);
nor U1553 (N_1553,N_40,N_654);
xor U1554 (N_1554,N_556,N_463);
xnor U1555 (N_1555,N_719,N_857);
nand U1556 (N_1556,N_345,N_560);
and U1557 (N_1557,N_137,N_885);
nand U1558 (N_1558,N_63,N_947);
xor U1559 (N_1559,N_827,N_463);
and U1560 (N_1560,N_991,N_869);
or U1561 (N_1561,N_4,N_393);
nand U1562 (N_1562,N_673,N_989);
and U1563 (N_1563,N_651,N_775);
or U1564 (N_1564,N_408,N_12);
and U1565 (N_1565,N_856,N_110);
nand U1566 (N_1566,N_507,N_470);
nand U1567 (N_1567,N_59,N_296);
xnor U1568 (N_1568,N_475,N_741);
or U1569 (N_1569,N_201,N_903);
or U1570 (N_1570,N_300,N_669);
xnor U1571 (N_1571,N_370,N_26);
or U1572 (N_1572,N_132,N_463);
or U1573 (N_1573,N_722,N_445);
nand U1574 (N_1574,N_544,N_49);
xnor U1575 (N_1575,N_188,N_145);
nor U1576 (N_1576,N_312,N_188);
and U1577 (N_1577,N_938,N_901);
xnor U1578 (N_1578,N_177,N_299);
or U1579 (N_1579,N_461,N_92);
xnor U1580 (N_1580,N_492,N_356);
xor U1581 (N_1581,N_925,N_285);
or U1582 (N_1582,N_793,N_229);
xnor U1583 (N_1583,N_456,N_335);
nor U1584 (N_1584,N_379,N_773);
or U1585 (N_1585,N_839,N_931);
nor U1586 (N_1586,N_960,N_425);
nand U1587 (N_1587,N_606,N_16);
or U1588 (N_1588,N_818,N_701);
xor U1589 (N_1589,N_869,N_975);
xnor U1590 (N_1590,N_726,N_491);
and U1591 (N_1591,N_927,N_859);
or U1592 (N_1592,N_499,N_474);
and U1593 (N_1593,N_427,N_620);
xnor U1594 (N_1594,N_543,N_442);
xnor U1595 (N_1595,N_965,N_553);
and U1596 (N_1596,N_694,N_47);
xor U1597 (N_1597,N_420,N_522);
and U1598 (N_1598,N_25,N_366);
xor U1599 (N_1599,N_201,N_318);
and U1600 (N_1600,N_570,N_649);
or U1601 (N_1601,N_745,N_20);
xor U1602 (N_1602,N_126,N_627);
or U1603 (N_1603,N_218,N_473);
or U1604 (N_1604,N_128,N_303);
or U1605 (N_1605,N_876,N_526);
and U1606 (N_1606,N_95,N_629);
xor U1607 (N_1607,N_196,N_992);
nand U1608 (N_1608,N_718,N_206);
or U1609 (N_1609,N_136,N_142);
and U1610 (N_1610,N_710,N_719);
xor U1611 (N_1611,N_513,N_536);
or U1612 (N_1612,N_794,N_931);
nand U1613 (N_1613,N_156,N_601);
and U1614 (N_1614,N_571,N_668);
and U1615 (N_1615,N_488,N_544);
and U1616 (N_1616,N_140,N_996);
xor U1617 (N_1617,N_849,N_98);
and U1618 (N_1618,N_512,N_706);
or U1619 (N_1619,N_450,N_97);
xnor U1620 (N_1620,N_707,N_819);
and U1621 (N_1621,N_38,N_950);
xor U1622 (N_1622,N_361,N_156);
nand U1623 (N_1623,N_13,N_595);
nand U1624 (N_1624,N_307,N_346);
nand U1625 (N_1625,N_817,N_460);
nor U1626 (N_1626,N_353,N_509);
nor U1627 (N_1627,N_531,N_210);
nand U1628 (N_1628,N_904,N_952);
nor U1629 (N_1629,N_186,N_152);
or U1630 (N_1630,N_87,N_567);
xor U1631 (N_1631,N_196,N_512);
and U1632 (N_1632,N_227,N_117);
and U1633 (N_1633,N_429,N_780);
nand U1634 (N_1634,N_332,N_951);
xor U1635 (N_1635,N_553,N_570);
nand U1636 (N_1636,N_102,N_417);
nand U1637 (N_1637,N_372,N_37);
nand U1638 (N_1638,N_703,N_791);
xnor U1639 (N_1639,N_535,N_340);
xor U1640 (N_1640,N_720,N_360);
or U1641 (N_1641,N_759,N_602);
xor U1642 (N_1642,N_289,N_514);
nor U1643 (N_1643,N_159,N_889);
and U1644 (N_1644,N_927,N_888);
xnor U1645 (N_1645,N_936,N_841);
xor U1646 (N_1646,N_507,N_352);
xor U1647 (N_1647,N_76,N_910);
nor U1648 (N_1648,N_512,N_218);
or U1649 (N_1649,N_794,N_502);
xor U1650 (N_1650,N_840,N_890);
and U1651 (N_1651,N_274,N_122);
or U1652 (N_1652,N_807,N_309);
nor U1653 (N_1653,N_750,N_186);
xnor U1654 (N_1654,N_575,N_160);
or U1655 (N_1655,N_63,N_304);
or U1656 (N_1656,N_598,N_232);
or U1657 (N_1657,N_782,N_923);
and U1658 (N_1658,N_253,N_225);
nand U1659 (N_1659,N_268,N_93);
nor U1660 (N_1660,N_48,N_536);
nor U1661 (N_1661,N_688,N_725);
and U1662 (N_1662,N_906,N_343);
xor U1663 (N_1663,N_799,N_290);
and U1664 (N_1664,N_286,N_799);
and U1665 (N_1665,N_40,N_294);
nand U1666 (N_1666,N_949,N_82);
or U1667 (N_1667,N_411,N_566);
or U1668 (N_1668,N_344,N_952);
and U1669 (N_1669,N_397,N_516);
xnor U1670 (N_1670,N_748,N_49);
xor U1671 (N_1671,N_914,N_65);
or U1672 (N_1672,N_950,N_167);
or U1673 (N_1673,N_149,N_170);
xor U1674 (N_1674,N_830,N_35);
xnor U1675 (N_1675,N_142,N_462);
xnor U1676 (N_1676,N_609,N_152);
xor U1677 (N_1677,N_837,N_522);
nand U1678 (N_1678,N_433,N_672);
nand U1679 (N_1679,N_183,N_4);
or U1680 (N_1680,N_555,N_658);
or U1681 (N_1681,N_856,N_727);
nand U1682 (N_1682,N_416,N_540);
nor U1683 (N_1683,N_589,N_170);
and U1684 (N_1684,N_949,N_156);
nor U1685 (N_1685,N_404,N_148);
nand U1686 (N_1686,N_893,N_389);
and U1687 (N_1687,N_368,N_708);
or U1688 (N_1688,N_365,N_784);
or U1689 (N_1689,N_390,N_797);
nor U1690 (N_1690,N_805,N_167);
or U1691 (N_1691,N_276,N_185);
nor U1692 (N_1692,N_280,N_408);
or U1693 (N_1693,N_576,N_57);
and U1694 (N_1694,N_895,N_358);
or U1695 (N_1695,N_758,N_780);
nor U1696 (N_1696,N_585,N_839);
xnor U1697 (N_1697,N_108,N_556);
nand U1698 (N_1698,N_849,N_50);
or U1699 (N_1699,N_977,N_634);
nor U1700 (N_1700,N_725,N_689);
and U1701 (N_1701,N_758,N_753);
xor U1702 (N_1702,N_904,N_300);
or U1703 (N_1703,N_588,N_232);
or U1704 (N_1704,N_499,N_875);
and U1705 (N_1705,N_953,N_889);
xnor U1706 (N_1706,N_512,N_937);
nand U1707 (N_1707,N_199,N_160);
or U1708 (N_1708,N_571,N_321);
xnor U1709 (N_1709,N_279,N_195);
and U1710 (N_1710,N_988,N_154);
or U1711 (N_1711,N_937,N_126);
nand U1712 (N_1712,N_236,N_490);
or U1713 (N_1713,N_659,N_814);
and U1714 (N_1714,N_378,N_999);
xor U1715 (N_1715,N_180,N_332);
and U1716 (N_1716,N_528,N_340);
and U1717 (N_1717,N_526,N_696);
or U1718 (N_1718,N_735,N_775);
nor U1719 (N_1719,N_151,N_517);
and U1720 (N_1720,N_110,N_72);
and U1721 (N_1721,N_458,N_355);
xor U1722 (N_1722,N_250,N_204);
or U1723 (N_1723,N_650,N_440);
nand U1724 (N_1724,N_367,N_858);
nor U1725 (N_1725,N_215,N_898);
or U1726 (N_1726,N_92,N_445);
and U1727 (N_1727,N_949,N_880);
and U1728 (N_1728,N_502,N_293);
nor U1729 (N_1729,N_225,N_891);
and U1730 (N_1730,N_415,N_245);
nand U1731 (N_1731,N_664,N_882);
nand U1732 (N_1732,N_27,N_672);
nand U1733 (N_1733,N_733,N_876);
nand U1734 (N_1734,N_316,N_874);
or U1735 (N_1735,N_332,N_947);
and U1736 (N_1736,N_754,N_392);
nand U1737 (N_1737,N_136,N_563);
and U1738 (N_1738,N_18,N_636);
xor U1739 (N_1739,N_174,N_180);
or U1740 (N_1740,N_537,N_386);
nor U1741 (N_1741,N_77,N_179);
xor U1742 (N_1742,N_879,N_307);
xor U1743 (N_1743,N_772,N_431);
and U1744 (N_1744,N_348,N_289);
or U1745 (N_1745,N_365,N_644);
nand U1746 (N_1746,N_641,N_520);
or U1747 (N_1747,N_411,N_464);
and U1748 (N_1748,N_602,N_28);
nand U1749 (N_1749,N_176,N_837);
and U1750 (N_1750,N_623,N_393);
xnor U1751 (N_1751,N_119,N_265);
and U1752 (N_1752,N_739,N_243);
nor U1753 (N_1753,N_144,N_504);
nand U1754 (N_1754,N_689,N_385);
nand U1755 (N_1755,N_452,N_2);
nand U1756 (N_1756,N_148,N_532);
xor U1757 (N_1757,N_258,N_883);
and U1758 (N_1758,N_188,N_209);
and U1759 (N_1759,N_326,N_907);
nand U1760 (N_1760,N_309,N_330);
nor U1761 (N_1761,N_842,N_456);
or U1762 (N_1762,N_232,N_255);
xnor U1763 (N_1763,N_269,N_628);
nor U1764 (N_1764,N_646,N_79);
nor U1765 (N_1765,N_657,N_190);
and U1766 (N_1766,N_685,N_299);
nand U1767 (N_1767,N_188,N_822);
nor U1768 (N_1768,N_315,N_649);
xor U1769 (N_1769,N_610,N_375);
xor U1770 (N_1770,N_893,N_705);
and U1771 (N_1771,N_396,N_554);
or U1772 (N_1772,N_764,N_251);
and U1773 (N_1773,N_162,N_529);
nor U1774 (N_1774,N_578,N_296);
nor U1775 (N_1775,N_757,N_543);
nor U1776 (N_1776,N_573,N_527);
xor U1777 (N_1777,N_511,N_102);
nor U1778 (N_1778,N_140,N_867);
xnor U1779 (N_1779,N_13,N_868);
nor U1780 (N_1780,N_4,N_10);
nor U1781 (N_1781,N_74,N_395);
xor U1782 (N_1782,N_440,N_833);
or U1783 (N_1783,N_922,N_752);
and U1784 (N_1784,N_652,N_13);
or U1785 (N_1785,N_681,N_512);
xor U1786 (N_1786,N_871,N_229);
nor U1787 (N_1787,N_260,N_979);
nand U1788 (N_1788,N_661,N_92);
or U1789 (N_1789,N_665,N_383);
nand U1790 (N_1790,N_98,N_980);
nor U1791 (N_1791,N_461,N_536);
and U1792 (N_1792,N_365,N_649);
nand U1793 (N_1793,N_740,N_256);
and U1794 (N_1794,N_46,N_387);
nand U1795 (N_1795,N_615,N_642);
xnor U1796 (N_1796,N_766,N_324);
nor U1797 (N_1797,N_748,N_356);
and U1798 (N_1798,N_246,N_216);
xor U1799 (N_1799,N_578,N_800);
xor U1800 (N_1800,N_972,N_288);
and U1801 (N_1801,N_861,N_416);
nand U1802 (N_1802,N_576,N_493);
xor U1803 (N_1803,N_255,N_373);
and U1804 (N_1804,N_147,N_785);
nand U1805 (N_1805,N_583,N_536);
and U1806 (N_1806,N_906,N_254);
and U1807 (N_1807,N_738,N_829);
nor U1808 (N_1808,N_231,N_97);
xnor U1809 (N_1809,N_732,N_786);
nor U1810 (N_1810,N_737,N_950);
nor U1811 (N_1811,N_711,N_291);
nand U1812 (N_1812,N_500,N_143);
and U1813 (N_1813,N_89,N_687);
or U1814 (N_1814,N_874,N_954);
nand U1815 (N_1815,N_791,N_821);
nand U1816 (N_1816,N_561,N_606);
nand U1817 (N_1817,N_700,N_780);
xnor U1818 (N_1818,N_989,N_539);
nand U1819 (N_1819,N_366,N_278);
nor U1820 (N_1820,N_984,N_714);
xnor U1821 (N_1821,N_733,N_815);
xor U1822 (N_1822,N_696,N_920);
and U1823 (N_1823,N_992,N_395);
or U1824 (N_1824,N_667,N_253);
xor U1825 (N_1825,N_981,N_147);
nor U1826 (N_1826,N_393,N_251);
nor U1827 (N_1827,N_998,N_283);
xnor U1828 (N_1828,N_205,N_582);
nand U1829 (N_1829,N_291,N_97);
and U1830 (N_1830,N_352,N_713);
or U1831 (N_1831,N_950,N_55);
nand U1832 (N_1832,N_828,N_163);
nor U1833 (N_1833,N_717,N_706);
nand U1834 (N_1834,N_652,N_966);
or U1835 (N_1835,N_680,N_331);
xnor U1836 (N_1836,N_121,N_738);
and U1837 (N_1837,N_364,N_183);
xnor U1838 (N_1838,N_215,N_60);
nor U1839 (N_1839,N_308,N_33);
nor U1840 (N_1840,N_322,N_409);
nand U1841 (N_1841,N_833,N_289);
and U1842 (N_1842,N_418,N_160);
nor U1843 (N_1843,N_697,N_194);
or U1844 (N_1844,N_354,N_562);
xor U1845 (N_1845,N_784,N_525);
nor U1846 (N_1846,N_32,N_792);
xnor U1847 (N_1847,N_346,N_411);
nand U1848 (N_1848,N_595,N_423);
xor U1849 (N_1849,N_46,N_2);
xor U1850 (N_1850,N_662,N_957);
or U1851 (N_1851,N_589,N_597);
or U1852 (N_1852,N_627,N_235);
nor U1853 (N_1853,N_961,N_844);
and U1854 (N_1854,N_841,N_495);
nor U1855 (N_1855,N_978,N_646);
nor U1856 (N_1856,N_228,N_615);
nand U1857 (N_1857,N_894,N_690);
or U1858 (N_1858,N_164,N_958);
nand U1859 (N_1859,N_161,N_66);
xor U1860 (N_1860,N_163,N_769);
nor U1861 (N_1861,N_730,N_342);
and U1862 (N_1862,N_445,N_434);
or U1863 (N_1863,N_500,N_982);
xnor U1864 (N_1864,N_896,N_382);
nand U1865 (N_1865,N_316,N_230);
nand U1866 (N_1866,N_318,N_716);
and U1867 (N_1867,N_864,N_251);
xnor U1868 (N_1868,N_185,N_941);
xor U1869 (N_1869,N_212,N_782);
nor U1870 (N_1870,N_968,N_119);
or U1871 (N_1871,N_802,N_190);
or U1872 (N_1872,N_556,N_773);
xor U1873 (N_1873,N_388,N_592);
or U1874 (N_1874,N_384,N_834);
xor U1875 (N_1875,N_146,N_325);
or U1876 (N_1876,N_909,N_725);
nand U1877 (N_1877,N_397,N_223);
or U1878 (N_1878,N_846,N_936);
or U1879 (N_1879,N_879,N_594);
and U1880 (N_1880,N_898,N_797);
nand U1881 (N_1881,N_870,N_303);
xnor U1882 (N_1882,N_287,N_714);
and U1883 (N_1883,N_143,N_606);
or U1884 (N_1884,N_112,N_232);
nor U1885 (N_1885,N_664,N_633);
nor U1886 (N_1886,N_482,N_435);
xor U1887 (N_1887,N_451,N_126);
nand U1888 (N_1888,N_786,N_859);
or U1889 (N_1889,N_429,N_438);
nor U1890 (N_1890,N_870,N_62);
nor U1891 (N_1891,N_261,N_412);
xor U1892 (N_1892,N_188,N_75);
and U1893 (N_1893,N_666,N_2);
xor U1894 (N_1894,N_130,N_5);
xnor U1895 (N_1895,N_381,N_316);
or U1896 (N_1896,N_379,N_671);
xnor U1897 (N_1897,N_214,N_447);
nand U1898 (N_1898,N_101,N_438);
xor U1899 (N_1899,N_591,N_12);
nor U1900 (N_1900,N_532,N_933);
xor U1901 (N_1901,N_112,N_733);
or U1902 (N_1902,N_55,N_36);
nor U1903 (N_1903,N_601,N_845);
nor U1904 (N_1904,N_519,N_829);
nand U1905 (N_1905,N_177,N_132);
nand U1906 (N_1906,N_140,N_884);
xor U1907 (N_1907,N_210,N_698);
or U1908 (N_1908,N_10,N_226);
and U1909 (N_1909,N_189,N_127);
or U1910 (N_1910,N_935,N_307);
or U1911 (N_1911,N_276,N_484);
xnor U1912 (N_1912,N_817,N_137);
xor U1913 (N_1913,N_901,N_330);
nand U1914 (N_1914,N_896,N_556);
nand U1915 (N_1915,N_838,N_837);
and U1916 (N_1916,N_204,N_888);
and U1917 (N_1917,N_447,N_833);
and U1918 (N_1918,N_134,N_828);
nor U1919 (N_1919,N_400,N_883);
or U1920 (N_1920,N_275,N_72);
nand U1921 (N_1921,N_154,N_493);
nand U1922 (N_1922,N_779,N_917);
or U1923 (N_1923,N_281,N_317);
xor U1924 (N_1924,N_857,N_657);
nand U1925 (N_1925,N_448,N_281);
nand U1926 (N_1926,N_251,N_708);
xnor U1927 (N_1927,N_874,N_228);
nand U1928 (N_1928,N_678,N_667);
nor U1929 (N_1929,N_462,N_780);
nor U1930 (N_1930,N_994,N_361);
and U1931 (N_1931,N_427,N_195);
nand U1932 (N_1932,N_966,N_617);
xor U1933 (N_1933,N_965,N_488);
nor U1934 (N_1934,N_449,N_905);
or U1935 (N_1935,N_399,N_266);
or U1936 (N_1936,N_997,N_618);
nor U1937 (N_1937,N_758,N_168);
or U1938 (N_1938,N_444,N_373);
nor U1939 (N_1939,N_978,N_555);
xnor U1940 (N_1940,N_804,N_488);
and U1941 (N_1941,N_338,N_995);
or U1942 (N_1942,N_734,N_298);
or U1943 (N_1943,N_481,N_894);
nand U1944 (N_1944,N_464,N_441);
or U1945 (N_1945,N_726,N_667);
and U1946 (N_1946,N_645,N_688);
or U1947 (N_1947,N_12,N_759);
nand U1948 (N_1948,N_634,N_817);
nor U1949 (N_1949,N_986,N_837);
or U1950 (N_1950,N_831,N_908);
nand U1951 (N_1951,N_457,N_84);
and U1952 (N_1952,N_451,N_694);
xnor U1953 (N_1953,N_341,N_164);
nor U1954 (N_1954,N_740,N_985);
nor U1955 (N_1955,N_426,N_683);
and U1956 (N_1956,N_285,N_977);
xor U1957 (N_1957,N_611,N_214);
nand U1958 (N_1958,N_940,N_532);
and U1959 (N_1959,N_864,N_640);
nand U1960 (N_1960,N_851,N_13);
or U1961 (N_1961,N_216,N_718);
or U1962 (N_1962,N_572,N_772);
and U1963 (N_1963,N_473,N_351);
xnor U1964 (N_1964,N_973,N_58);
xnor U1965 (N_1965,N_605,N_294);
and U1966 (N_1966,N_263,N_3);
nand U1967 (N_1967,N_366,N_275);
xor U1968 (N_1968,N_553,N_824);
nand U1969 (N_1969,N_615,N_833);
nor U1970 (N_1970,N_83,N_912);
and U1971 (N_1971,N_906,N_948);
or U1972 (N_1972,N_965,N_567);
xnor U1973 (N_1973,N_939,N_612);
xor U1974 (N_1974,N_831,N_541);
and U1975 (N_1975,N_546,N_618);
nor U1976 (N_1976,N_666,N_22);
or U1977 (N_1977,N_762,N_872);
nand U1978 (N_1978,N_947,N_70);
or U1979 (N_1979,N_374,N_953);
and U1980 (N_1980,N_860,N_853);
nand U1981 (N_1981,N_463,N_619);
and U1982 (N_1982,N_541,N_201);
nand U1983 (N_1983,N_590,N_52);
nor U1984 (N_1984,N_297,N_983);
and U1985 (N_1985,N_695,N_558);
nand U1986 (N_1986,N_371,N_405);
nor U1987 (N_1987,N_737,N_316);
nand U1988 (N_1988,N_285,N_730);
nor U1989 (N_1989,N_771,N_948);
xor U1990 (N_1990,N_655,N_646);
nor U1991 (N_1991,N_373,N_852);
nor U1992 (N_1992,N_327,N_124);
xnor U1993 (N_1993,N_391,N_468);
nand U1994 (N_1994,N_71,N_746);
or U1995 (N_1995,N_605,N_239);
nand U1996 (N_1996,N_499,N_899);
or U1997 (N_1997,N_330,N_254);
nand U1998 (N_1998,N_268,N_519);
or U1999 (N_1999,N_240,N_408);
nor U2000 (N_2000,N_1511,N_1918);
and U2001 (N_2001,N_1464,N_1973);
nor U2002 (N_2002,N_1446,N_1099);
and U2003 (N_2003,N_1055,N_1080);
nor U2004 (N_2004,N_1359,N_1412);
xnor U2005 (N_2005,N_1350,N_1500);
and U2006 (N_2006,N_1279,N_1353);
and U2007 (N_2007,N_1823,N_1104);
nand U2008 (N_2008,N_1056,N_1959);
nor U2009 (N_2009,N_1836,N_1762);
xnor U2010 (N_2010,N_1872,N_1127);
xnor U2011 (N_2011,N_1969,N_1718);
and U2012 (N_2012,N_1401,N_1999);
and U2013 (N_2013,N_1803,N_1314);
nor U2014 (N_2014,N_1981,N_1114);
nand U2015 (N_2015,N_1727,N_1550);
nor U2016 (N_2016,N_1186,N_1273);
and U2017 (N_2017,N_1945,N_1675);
nand U2018 (N_2018,N_1863,N_1925);
nand U2019 (N_2019,N_1492,N_1691);
xnor U2020 (N_2020,N_1032,N_1924);
xor U2021 (N_2021,N_1684,N_1390);
or U2022 (N_2022,N_1790,N_1749);
and U2023 (N_2023,N_1028,N_1225);
xnor U2024 (N_2024,N_1392,N_1816);
nand U2025 (N_2025,N_1929,N_1571);
nor U2026 (N_2026,N_1797,N_1370);
nor U2027 (N_2027,N_1341,N_1011);
nor U2028 (N_2028,N_1449,N_1840);
nand U2029 (N_2029,N_1319,N_1021);
nand U2030 (N_2030,N_1564,N_1502);
nand U2031 (N_2031,N_1213,N_1951);
nand U2032 (N_2032,N_1156,N_1327);
and U2033 (N_2033,N_1996,N_1100);
nand U2034 (N_2034,N_1585,N_1263);
and U2035 (N_2035,N_1133,N_1938);
or U2036 (N_2036,N_1381,N_1421);
nand U2037 (N_2037,N_1905,N_1636);
xnor U2038 (N_2038,N_1754,N_1694);
xnor U2039 (N_2039,N_1722,N_1460);
or U2040 (N_2040,N_1639,N_1185);
or U2041 (N_2041,N_1909,N_1025);
nand U2042 (N_2042,N_1868,N_1683);
xnor U2043 (N_2043,N_1424,N_1656);
xnor U2044 (N_2044,N_1833,N_1807);
nand U2045 (N_2045,N_1997,N_1526);
or U2046 (N_2046,N_1497,N_1117);
nand U2047 (N_2047,N_1400,N_1804);
and U2048 (N_2048,N_1292,N_1869);
and U2049 (N_2049,N_1825,N_1129);
and U2050 (N_2050,N_1619,N_1020);
xor U2051 (N_2051,N_1461,N_1196);
nor U2052 (N_2052,N_1764,N_1053);
nor U2053 (N_2053,N_1766,N_1626);
nand U2054 (N_2054,N_1422,N_1706);
or U2055 (N_2055,N_1544,N_1321);
and U2056 (N_2056,N_1465,N_1037);
nand U2057 (N_2057,N_1463,N_1505);
or U2058 (N_2058,N_1955,N_1111);
xnor U2059 (N_2059,N_1010,N_1264);
xor U2060 (N_2060,N_1972,N_1148);
and U2061 (N_2061,N_1748,N_1160);
xor U2062 (N_2062,N_1176,N_1587);
nor U2063 (N_2063,N_1755,N_1235);
or U2064 (N_2064,N_1128,N_1313);
and U2065 (N_2065,N_1956,N_1533);
and U2066 (N_2066,N_1077,N_1954);
or U2067 (N_2067,N_1680,N_1495);
and U2068 (N_2068,N_1480,N_1678);
xnor U2069 (N_2069,N_1976,N_1658);
xnor U2070 (N_2070,N_1700,N_1499);
or U2071 (N_2071,N_1484,N_1509);
xnor U2072 (N_2072,N_1591,N_1510);
xnor U2073 (N_2073,N_1805,N_1512);
xnor U2074 (N_2074,N_1076,N_1543);
xor U2075 (N_2075,N_1130,N_1625);
nor U2076 (N_2076,N_1473,N_1328);
nand U2077 (N_2077,N_1476,N_1709);
nand U2078 (N_2078,N_1151,N_1962);
nor U2079 (N_2079,N_1781,N_1627);
nand U2080 (N_2080,N_1751,N_1245);
nand U2081 (N_2081,N_1851,N_1943);
and U2082 (N_2082,N_1802,N_1087);
xnor U2083 (N_2083,N_1306,N_1758);
and U2084 (N_2084,N_1887,N_1047);
nor U2085 (N_2085,N_1072,N_1848);
nand U2086 (N_2086,N_1173,N_1960);
nor U2087 (N_2087,N_1197,N_1092);
and U2088 (N_2088,N_1271,N_1368);
xor U2089 (N_2089,N_1190,N_1578);
nand U2090 (N_2090,N_1682,N_1144);
nand U2091 (N_2091,N_1489,N_1435);
xor U2092 (N_2092,N_1559,N_1064);
xor U2093 (N_2093,N_1853,N_1702);
nor U2094 (N_2094,N_1006,N_1791);
or U2095 (N_2095,N_1725,N_1763);
nor U2096 (N_2096,N_1407,N_1441);
and U2097 (N_2097,N_1599,N_1039);
or U2098 (N_2098,N_1134,N_1685);
and U2099 (N_2099,N_1756,N_1590);
or U2100 (N_2100,N_1583,N_1004);
nor U2101 (N_2101,N_1681,N_1646);
nor U2102 (N_2102,N_1813,N_1101);
nor U2103 (N_2103,N_1574,N_1944);
or U2104 (N_2104,N_1601,N_1112);
nand U2105 (N_2105,N_1613,N_1908);
nand U2106 (N_2106,N_1082,N_1164);
nor U2107 (N_2107,N_1847,N_1491);
or U2108 (N_2108,N_1062,N_1690);
nor U2109 (N_2109,N_1671,N_1695);
xnor U2110 (N_2110,N_1391,N_1961);
xor U2111 (N_2111,N_1124,N_1881);
nor U2112 (N_2112,N_1211,N_1467);
xor U2113 (N_2113,N_1565,N_1913);
or U2114 (N_2114,N_1459,N_1462);
xnor U2115 (N_2115,N_1146,N_1677);
nand U2116 (N_2116,N_1261,N_1323);
nor U2117 (N_2117,N_1631,N_1773);
nand U2118 (N_2118,N_1102,N_1934);
nand U2119 (N_2119,N_1482,N_1882);
and U2120 (N_2120,N_1902,N_1932);
xor U2121 (N_2121,N_1079,N_1257);
nor U2122 (N_2122,N_1411,N_1380);
nand U2123 (N_2123,N_1324,N_1107);
nor U2124 (N_2124,N_1483,N_1506);
or U2125 (N_2125,N_1428,N_1985);
xor U2126 (N_2126,N_1771,N_1921);
and U2127 (N_2127,N_1720,N_1369);
nor U2128 (N_2128,N_1494,N_1209);
and U2129 (N_2129,N_1942,N_1545);
or U2130 (N_2130,N_1238,N_1255);
and U2131 (N_2131,N_1439,N_1230);
xor U2132 (N_2132,N_1356,N_1674);
xnor U2133 (N_2133,N_1901,N_1745);
and U2134 (N_2134,N_1995,N_1721);
or U2135 (N_2135,N_1679,N_1811);
or U2136 (N_2136,N_1325,N_1534);
and U2137 (N_2137,N_1384,N_1457);
xor U2138 (N_2138,N_1864,N_1360);
nand U2139 (N_2139,N_1192,N_1315);
nor U2140 (N_2140,N_1689,N_1701);
or U2141 (N_2141,N_1715,N_1386);
xor U2142 (N_2142,N_1178,N_1793);
and U2143 (N_2143,N_1195,N_1531);
xnor U2144 (N_2144,N_1644,N_1774);
or U2145 (N_2145,N_1275,N_1983);
and U2146 (N_2146,N_1091,N_1598);
and U2147 (N_2147,N_1856,N_1068);
or U2148 (N_2148,N_1686,N_1035);
nor U2149 (N_2149,N_1903,N_1635);
nor U2150 (N_2150,N_1189,N_1661);
or U2151 (N_2151,N_1251,N_1885);
and U2152 (N_2152,N_1865,N_1736);
xor U2153 (N_2153,N_1085,N_1937);
xnor U2154 (N_2154,N_1719,N_1743);
nor U2155 (N_2155,N_1294,N_1249);
and U2156 (N_2156,N_1078,N_1979);
and U2157 (N_2157,N_1479,N_1474);
nor U2158 (N_2158,N_1866,N_1377);
nor U2159 (N_2159,N_1397,N_1002);
and U2160 (N_2160,N_1224,N_1250);
xor U2161 (N_2161,N_1917,N_1567);
xor U2162 (N_2162,N_1334,N_1330);
xor U2163 (N_2163,N_1931,N_1054);
xnor U2164 (N_2164,N_1606,N_1270);
nor U2165 (N_2165,N_1935,N_1241);
xor U2166 (N_2166,N_1783,N_1012);
nor U2167 (N_2167,N_1001,N_1450);
nand U2168 (N_2168,N_1883,N_1592);
xnor U2169 (N_2169,N_1523,N_1553);
xor U2170 (N_2170,N_1824,N_1466);
xnor U2171 (N_2171,N_1285,N_1729);
xnor U2172 (N_2172,N_1974,N_1304);
nor U2173 (N_2173,N_1637,N_1288);
xnor U2174 (N_2174,N_1896,N_1005);
or U2175 (N_2175,N_1501,N_1308);
or U2176 (N_2176,N_1726,N_1141);
nand U2177 (N_2177,N_1894,N_1958);
and U2178 (N_2178,N_1967,N_1094);
and U2179 (N_2179,N_1916,N_1303);
and U2180 (N_2180,N_1546,N_1535);
xor U2181 (N_2181,N_1188,N_1788);
nor U2182 (N_2182,N_1207,N_1723);
and U2183 (N_2183,N_1612,N_1216);
nand U2184 (N_2184,N_1222,N_1815);
nor U2185 (N_2185,N_1965,N_1800);
nor U2186 (N_2186,N_1568,N_1518);
xnor U2187 (N_2187,N_1529,N_1109);
nand U2188 (N_2188,N_1968,N_1456);
or U2189 (N_2189,N_1915,N_1414);
or U2190 (N_2190,N_1507,N_1427);
and U2191 (N_2191,N_1106,N_1821);
nor U2192 (N_2192,N_1110,N_1817);
nor U2193 (N_2193,N_1605,N_1317);
xnor U2194 (N_2194,N_1859,N_1069);
and U2195 (N_2195,N_1454,N_1268);
and U2196 (N_2196,N_1448,N_1750);
xnor U2197 (N_2197,N_1152,N_1378);
nor U2198 (N_2198,N_1581,N_1738);
and U2199 (N_2199,N_1071,N_1322);
and U2200 (N_2200,N_1551,N_1346);
nor U2201 (N_2201,N_1367,N_1597);
nand U2202 (N_2202,N_1073,N_1044);
nand U2203 (N_2203,N_1170,N_1858);
xnor U2204 (N_2204,N_1385,N_1291);
xnor U2205 (N_2205,N_1589,N_1892);
or U2206 (N_2206,N_1794,N_1237);
and U2207 (N_2207,N_1352,N_1003);
nor U2208 (N_2208,N_1812,N_1120);
or U2209 (N_2209,N_1329,N_1052);
and U2210 (N_2210,N_1880,N_1277);
and U2211 (N_2211,N_1066,N_1673);
or U2212 (N_2212,N_1042,N_1991);
nor U2213 (N_2213,N_1232,N_1137);
or U2214 (N_2214,N_1978,N_1442);
nand U2215 (N_2215,N_1218,N_1150);
nand U2216 (N_2216,N_1014,N_1452);
nor U2217 (N_2217,N_1017,N_1900);
xor U2218 (N_2218,N_1373,N_1946);
xor U2219 (N_2219,N_1734,N_1179);
nor U2220 (N_2220,N_1493,N_1552);
nand U2221 (N_2221,N_1579,N_1286);
nor U2222 (N_2222,N_1714,N_1787);
nand U2223 (N_2223,N_1132,N_1970);
nand U2224 (N_2224,N_1167,N_1349);
xor U2225 (N_2225,N_1547,N_1065);
or U2226 (N_2226,N_1784,N_1290);
nor U2227 (N_2227,N_1418,N_1514);
xor U2228 (N_2228,N_1486,N_1562);
xor U2229 (N_2229,N_1116,N_1074);
xnor U2230 (N_2230,N_1844,N_1839);
nor U2231 (N_2231,N_1202,N_1095);
and U2232 (N_2232,N_1036,N_1363);
nor U2233 (N_2233,N_1398,N_1712);
and U2234 (N_2234,N_1532,N_1335);
xor U2235 (N_2235,N_1309,N_1382);
xor U2236 (N_2236,N_1860,N_1366);
and U2237 (N_2237,N_1050,N_1650);
nand U2238 (N_2238,N_1785,N_1301);
and U2239 (N_2239,N_1582,N_1379);
or U2240 (N_2240,N_1293,N_1469);
nand U2241 (N_2241,N_1888,N_1159);
or U2242 (N_2242,N_1737,N_1830);
xnor U2243 (N_2243,N_1283,N_1707);
xor U2244 (N_2244,N_1478,N_1402);
nand U2245 (N_2245,N_1242,N_1394);
xor U2246 (N_2246,N_1419,N_1410);
nand U2247 (N_2247,N_1770,N_1776);
nand U2248 (N_2248,N_1539,N_1375);
and U2249 (N_2249,N_1549,N_1862);
nand U2250 (N_2250,N_1267,N_1614);
nor U2251 (N_2251,N_1618,N_1593);
or U2252 (N_2252,N_1098,N_1113);
or U2253 (N_2253,N_1557,N_1229);
and U2254 (N_2254,N_1697,N_1563);
or U2255 (N_2255,N_1090,N_1395);
or U2256 (N_2256,N_1498,N_1611);
and U2257 (N_2257,N_1698,N_1822);
or U2258 (N_2258,N_1140,N_1629);
or U2259 (N_2259,N_1947,N_1259);
and U2260 (N_2260,N_1520,N_1300);
nor U2261 (N_2261,N_1121,N_1299);
or U2262 (N_2262,N_1119,N_1425);
or U2263 (N_2263,N_1759,N_1655);
and U2264 (N_2264,N_1841,N_1540);
or U2265 (N_2265,N_1354,N_1772);
nor U2266 (N_2266,N_1873,N_1302);
and U2267 (N_2267,N_1244,N_1818);
and U2268 (N_2268,N_1857,N_1835);
or U2269 (N_2269,N_1215,N_1051);
or U2270 (N_2270,N_1657,N_1024);
and U2271 (N_2271,N_1645,N_1846);
and U2272 (N_2272,N_1886,N_1716);
nor U2273 (N_2273,N_1827,N_1345);
nand U2274 (N_2274,N_1515,N_1573);
nor U2275 (N_2275,N_1084,N_1408);
nor U2276 (N_2276,N_1426,N_1634);
nand U2277 (N_2277,N_1168,N_1642);
nor U2278 (N_2278,N_1941,N_1537);
nand U2279 (N_2279,N_1747,N_1871);
and U2280 (N_2280,N_1984,N_1029);
nor U2281 (N_2281,N_1198,N_1855);
nand U2282 (N_2282,N_1409,N_1138);
xor U2283 (N_2283,N_1775,N_1096);
and U2284 (N_2284,N_1624,N_1554);
nand U2285 (N_2285,N_1210,N_1236);
nor U2286 (N_2286,N_1849,N_1383);
nor U2287 (N_2287,N_1240,N_1861);
nand U2288 (N_2288,N_1490,N_1992);
nor U2289 (N_2289,N_1633,N_1342);
and U2290 (N_2290,N_1687,N_1027);
or U2291 (N_2291,N_1513,N_1994);
or U2292 (N_2292,N_1212,N_1975);
nand U2293 (N_2293,N_1699,N_1193);
and U2294 (N_2294,N_1374,N_1870);
and U2295 (N_2295,N_1089,N_1522);
and U2296 (N_2296,N_1744,N_1971);
and U2297 (N_2297,N_1911,N_1423);
xnor U2298 (N_2298,N_1157,N_1337);
or U2299 (N_2299,N_1045,N_1149);
and U2300 (N_2300,N_1060,N_1226);
nor U2301 (N_2301,N_1355,N_1191);
nor U2302 (N_2302,N_1664,N_1161);
and U2303 (N_2303,N_1019,N_1649);
and U2304 (N_2304,N_1906,N_1525);
nor U2305 (N_2305,N_1586,N_1013);
and U2306 (N_2306,N_1181,N_1757);
nand U2307 (N_2307,N_1158,N_1576);
and U2308 (N_2308,N_1524,N_1431);
nand U2309 (N_2309,N_1340,N_1284);
xnor U2310 (N_2310,N_1103,N_1575);
nand U2311 (N_2311,N_1007,N_1023);
xor U2312 (N_2312,N_1123,N_1852);
nor U2313 (N_2313,N_1993,N_1280);
nor U2314 (N_2314,N_1388,N_1980);
nand U2315 (N_2315,N_1753,N_1538);
nor U2316 (N_2316,N_1845,N_1708);
or U2317 (N_2317,N_1604,N_1171);
or U2318 (N_2318,N_1767,N_1075);
xnor U2319 (N_2319,N_1765,N_1227);
xnor U2320 (N_2320,N_1610,N_1620);
xor U2321 (N_2321,N_1086,N_1471);
and U2322 (N_2322,N_1405,N_1434);
nor U2323 (N_2323,N_1016,N_1221);
xnor U2324 (N_2324,N_1616,N_1806);
and U2325 (N_2325,N_1891,N_1070);
xnor U2326 (N_2326,N_1603,N_1049);
xor U2327 (N_2327,N_1752,N_1986);
and U2328 (N_2328,N_1258,N_1733);
xor U2329 (N_2329,N_1118,N_1820);
or U2330 (N_2330,N_1662,N_1663);
nand U2331 (N_2331,N_1436,N_1950);
nand U2332 (N_2332,N_1200,N_1541);
nand U2333 (N_2333,N_1332,N_1615);
nor U2334 (N_2334,N_1630,N_1939);
nand U2335 (N_2335,N_1338,N_1761);
nor U2336 (N_2336,N_1796,N_1348);
and U2337 (N_2337,N_1180,N_1415);
xor U2338 (N_2338,N_1711,N_1208);
or U2339 (N_2339,N_1728,N_1331);
nor U2340 (N_2340,N_1287,N_1632);
or U2341 (N_2341,N_1115,N_1289);
nor U2342 (N_2342,N_1654,N_1651);
nor U2343 (N_2343,N_1361,N_1399);
nand U2344 (N_2344,N_1808,N_1254);
nor U2345 (N_2345,N_1688,N_1162);
xnor U2346 (N_2346,N_1879,N_1081);
nand U2347 (N_2347,N_1187,N_1282);
nor U2348 (N_2348,N_1364,N_1488);
or U2349 (N_2349,N_1778,N_1219);
or U2350 (N_2350,N_1890,N_1949);
nor U2351 (N_2351,N_1878,N_1223);
nor U2352 (N_2352,N_1217,N_1204);
xnor U2353 (N_2353,N_1919,N_1247);
nand U2354 (N_2354,N_1713,N_1595);
or U2355 (N_2355,N_1233,N_1067);
or U2356 (N_2356,N_1740,N_1372);
nand U2357 (N_2357,N_1692,N_1622);
and U2358 (N_2358,N_1030,N_1310);
nand U2359 (N_2359,N_1147,N_1246);
xor U2360 (N_2360,N_1199,N_1169);
and U2361 (N_2361,N_1566,N_1000);
nand U2362 (N_2362,N_1730,N_1660);
or U2363 (N_2363,N_1362,N_1516);
nor U2364 (N_2364,N_1977,N_1026);
xnor U2365 (N_2365,N_1136,N_1819);
xor U2366 (N_2366,N_1311,N_1780);
nor U2367 (N_2367,N_1838,N_1628);
nor U2368 (N_2368,N_1305,N_1814);
nor U2369 (N_2369,N_1854,N_1357);
nor U2370 (N_2370,N_1703,N_1358);
or U2371 (N_2371,N_1899,N_1406);
and U2372 (N_2372,N_1850,N_1920);
or U2373 (N_2373,N_1952,N_1298);
or U2374 (N_2374,N_1470,N_1741);
or U2375 (N_2375,N_1307,N_1640);
and U2376 (N_2376,N_1269,N_1481);
or U2377 (N_2377,N_1059,N_1572);
or U2378 (N_2378,N_1966,N_1165);
xor U2379 (N_2379,N_1914,N_1867);
nand U2380 (N_2380,N_1046,N_1731);
and U2381 (N_2381,N_1989,N_1666);
nand U2382 (N_2382,N_1617,N_1982);
xor U2383 (N_2383,N_1875,N_1792);
nand U2384 (N_2384,N_1239,N_1953);
and U2385 (N_2385,N_1155,N_1536);
xnor U2386 (N_2386,N_1876,N_1560);
xnor U2387 (N_2387,N_1131,N_1668);
nand U2388 (N_2388,N_1496,N_1638);
xnor U2389 (N_2389,N_1710,N_1256);
xnor U2390 (N_2390,N_1834,N_1831);
or U2391 (N_2391,N_1561,N_1122);
xnor U2392 (N_2392,N_1600,N_1177);
nand U2393 (N_2393,N_1798,N_1445);
nor U2394 (N_2394,N_1214,N_1735);
nand U2395 (N_2395,N_1907,N_1503);
or U2396 (N_2396,N_1704,N_1588);
or U2397 (N_2397,N_1033,N_1556);
or U2398 (N_2398,N_1927,N_1607);
and U2399 (N_2399,N_1432,N_1904);
xor U2400 (N_2400,N_1444,N_1057);
nor U2401 (N_2401,N_1231,N_1933);
nand U2402 (N_2402,N_1438,N_1316);
nor U2403 (N_2403,N_1040,N_1205);
xnor U2404 (N_2404,N_1018,N_1829);
nand U2405 (N_2405,N_1504,N_1810);
xor U2406 (N_2406,N_1228,N_1570);
nand U2407 (N_2407,N_1458,N_1403);
xor U2408 (N_2408,N_1339,N_1542);
and U2409 (N_2409,N_1260,N_1670);
and U2410 (N_2410,N_1371,N_1837);
and U2411 (N_2411,N_1608,N_1125);
nand U2412 (N_2412,N_1468,N_1912);
xnor U2413 (N_2413,N_1295,N_1453);
xor U2414 (N_2414,N_1387,N_1987);
or U2415 (N_2415,N_1717,N_1786);
and U2416 (N_2416,N_1963,N_1889);
or U2417 (N_2417,N_1936,N_1031);
or U2418 (N_2418,N_1333,N_1577);
nand U2419 (N_2419,N_1347,N_1248);
nand U2420 (N_2420,N_1154,N_1182);
or U2421 (N_2421,N_1430,N_1376);
nor U2422 (N_2422,N_1009,N_1487);
nor U2423 (N_2423,N_1724,N_1093);
xnor U2424 (N_2424,N_1139,N_1326);
nand U2425 (N_2425,N_1665,N_1643);
or U2426 (N_2426,N_1143,N_1063);
or U2427 (N_2427,N_1022,N_1530);
nor U2428 (N_2428,N_1433,N_1455);
nor U2429 (N_2429,N_1884,N_1922);
nand U2430 (N_2430,N_1447,N_1647);
nand U2431 (N_2431,N_1548,N_1826);
nor U2432 (N_2432,N_1351,N_1343);
or U2433 (N_2433,N_1693,N_1517);
nor U2434 (N_2434,N_1153,N_1253);
and U2435 (N_2435,N_1083,N_1957);
nor U2436 (N_2436,N_1145,N_1404);
or U2437 (N_2437,N_1252,N_1088);
or U2438 (N_2438,N_1528,N_1194);
xnor U2439 (N_2439,N_1521,N_1344);
nor U2440 (N_2440,N_1653,N_1842);
nand U2441 (N_2441,N_1417,N_1440);
nand U2442 (N_2442,N_1206,N_1201);
nand U2443 (N_2443,N_1998,N_1281);
xor U2444 (N_2444,N_1895,N_1472);
nor U2445 (N_2445,N_1320,N_1061);
nand U2446 (N_2446,N_1832,N_1318);
nor U2447 (N_2447,N_1809,N_1243);
xor U2448 (N_2448,N_1964,N_1266);
or U2449 (N_2449,N_1746,N_1779);
xnor U2450 (N_2450,N_1527,N_1782);
nor U2451 (N_2451,N_1135,N_1166);
xor U2452 (N_2452,N_1940,N_1008);
xor U2453 (N_2453,N_1297,N_1659);
nand U2454 (N_2454,N_1183,N_1041);
and U2455 (N_2455,N_1203,N_1519);
nor U2456 (N_2456,N_1508,N_1108);
nor U2457 (N_2457,N_1485,N_1777);
nand U2458 (N_2458,N_1990,N_1828);
or U2459 (N_2459,N_1609,N_1877);
or U2460 (N_2460,N_1175,N_1555);
nand U2461 (N_2461,N_1843,N_1898);
or U2462 (N_2462,N_1789,N_1584);
nor U2463 (N_2463,N_1184,N_1477);
nand U2464 (N_2464,N_1893,N_1648);
nand U2465 (N_2465,N_1769,N_1163);
and U2466 (N_2466,N_1038,N_1897);
or U2467 (N_2467,N_1336,N_1274);
xnor U2468 (N_2468,N_1272,N_1278);
and U2469 (N_2469,N_1416,N_1652);
and U2470 (N_2470,N_1389,N_1437);
nor U2471 (N_2471,N_1928,N_1602);
nor U2472 (N_2472,N_1742,N_1234);
nor U2473 (N_2473,N_1558,N_1396);
and U2474 (N_2474,N_1451,N_1795);
xor U2475 (N_2475,N_1105,N_1594);
and U2476 (N_2476,N_1097,N_1569);
xor U2477 (N_2477,N_1174,N_1676);
and U2478 (N_2478,N_1799,N_1220);
and U2479 (N_2479,N_1596,N_1669);
nand U2480 (N_2480,N_1015,N_1296);
xnor U2481 (N_2481,N_1312,N_1475);
xnor U2482 (N_2482,N_1420,N_1988);
or U2483 (N_2483,N_1365,N_1948);
and U2484 (N_2484,N_1262,N_1265);
and U2485 (N_2485,N_1768,N_1923);
nand U2486 (N_2486,N_1621,N_1443);
nor U2487 (N_2487,N_1413,N_1760);
nor U2488 (N_2488,N_1034,N_1623);
nor U2489 (N_2489,N_1126,N_1732);
or U2490 (N_2490,N_1393,N_1739);
nand U2491 (N_2491,N_1801,N_1696);
or U2492 (N_2492,N_1641,N_1926);
nor U2493 (N_2493,N_1142,N_1910);
xnor U2494 (N_2494,N_1705,N_1580);
and U2495 (N_2495,N_1672,N_1058);
and U2496 (N_2496,N_1048,N_1874);
nand U2497 (N_2497,N_1667,N_1043);
or U2498 (N_2498,N_1429,N_1172);
or U2499 (N_2499,N_1930,N_1276);
or U2500 (N_2500,N_1699,N_1069);
nand U2501 (N_2501,N_1050,N_1332);
or U2502 (N_2502,N_1193,N_1520);
or U2503 (N_2503,N_1295,N_1264);
xor U2504 (N_2504,N_1263,N_1628);
xor U2505 (N_2505,N_1426,N_1073);
nand U2506 (N_2506,N_1768,N_1409);
nand U2507 (N_2507,N_1987,N_1130);
and U2508 (N_2508,N_1378,N_1734);
xor U2509 (N_2509,N_1424,N_1877);
xnor U2510 (N_2510,N_1732,N_1231);
nor U2511 (N_2511,N_1027,N_1309);
nor U2512 (N_2512,N_1007,N_1319);
and U2513 (N_2513,N_1526,N_1801);
or U2514 (N_2514,N_1485,N_1836);
nand U2515 (N_2515,N_1537,N_1973);
nor U2516 (N_2516,N_1301,N_1718);
nand U2517 (N_2517,N_1018,N_1435);
and U2518 (N_2518,N_1176,N_1444);
or U2519 (N_2519,N_1809,N_1992);
or U2520 (N_2520,N_1797,N_1276);
xor U2521 (N_2521,N_1934,N_1356);
xor U2522 (N_2522,N_1408,N_1232);
and U2523 (N_2523,N_1183,N_1491);
or U2524 (N_2524,N_1602,N_1674);
xor U2525 (N_2525,N_1319,N_1732);
xnor U2526 (N_2526,N_1064,N_1816);
nor U2527 (N_2527,N_1387,N_1682);
nor U2528 (N_2528,N_1164,N_1040);
xnor U2529 (N_2529,N_1523,N_1992);
nor U2530 (N_2530,N_1621,N_1922);
and U2531 (N_2531,N_1369,N_1737);
and U2532 (N_2532,N_1692,N_1841);
nand U2533 (N_2533,N_1250,N_1165);
or U2534 (N_2534,N_1125,N_1675);
or U2535 (N_2535,N_1056,N_1360);
and U2536 (N_2536,N_1454,N_1774);
or U2537 (N_2537,N_1806,N_1304);
and U2538 (N_2538,N_1503,N_1462);
nand U2539 (N_2539,N_1788,N_1484);
nand U2540 (N_2540,N_1574,N_1885);
or U2541 (N_2541,N_1826,N_1275);
and U2542 (N_2542,N_1667,N_1315);
and U2543 (N_2543,N_1094,N_1958);
xnor U2544 (N_2544,N_1419,N_1568);
and U2545 (N_2545,N_1490,N_1881);
or U2546 (N_2546,N_1229,N_1661);
xnor U2547 (N_2547,N_1317,N_1504);
nand U2548 (N_2548,N_1613,N_1389);
xor U2549 (N_2549,N_1769,N_1262);
nor U2550 (N_2550,N_1845,N_1137);
nand U2551 (N_2551,N_1940,N_1004);
nand U2552 (N_2552,N_1229,N_1399);
nand U2553 (N_2553,N_1023,N_1967);
xor U2554 (N_2554,N_1832,N_1647);
xor U2555 (N_2555,N_1723,N_1717);
xnor U2556 (N_2556,N_1559,N_1233);
xnor U2557 (N_2557,N_1381,N_1811);
and U2558 (N_2558,N_1630,N_1149);
nand U2559 (N_2559,N_1613,N_1825);
xor U2560 (N_2560,N_1479,N_1323);
nor U2561 (N_2561,N_1486,N_1003);
xnor U2562 (N_2562,N_1594,N_1275);
or U2563 (N_2563,N_1682,N_1497);
or U2564 (N_2564,N_1775,N_1628);
or U2565 (N_2565,N_1116,N_1786);
or U2566 (N_2566,N_1500,N_1123);
nand U2567 (N_2567,N_1497,N_1930);
xnor U2568 (N_2568,N_1992,N_1810);
nand U2569 (N_2569,N_1144,N_1130);
nor U2570 (N_2570,N_1570,N_1089);
and U2571 (N_2571,N_1839,N_1091);
nor U2572 (N_2572,N_1480,N_1525);
and U2573 (N_2573,N_1423,N_1833);
xnor U2574 (N_2574,N_1727,N_1865);
or U2575 (N_2575,N_1094,N_1442);
xnor U2576 (N_2576,N_1194,N_1357);
xor U2577 (N_2577,N_1135,N_1258);
nor U2578 (N_2578,N_1223,N_1010);
nand U2579 (N_2579,N_1429,N_1587);
nand U2580 (N_2580,N_1127,N_1923);
or U2581 (N_2581,N_1883,N_1329);
xor U2582 (N_2582,N_1693,N_1359);
nand U2583 (N_2583,N_1957,N_1362);
nand U2584 (N_2584,N_1938,N_1914);
nand U2585 (N_2585,N_1546,N_1126);
nor U2586 (N_2586,N_1113,N_1362);
nor U2587 (N_2587,N_1192,N_1752);
nand U2588 (N_2588,N_1216,N_1819);
or U2589 (N_2589,N_1481,N_1318);
xnor U2590 (N_2590,N_1337,N_1230);
or U2591 (N_2591,N_1126,N_1993);
or U2592 (N_2592,N_1664,N_1268);
nand U2593 (N_2593,N_1896,N_1751);
and U2594 (N_2594,N_1360,N_1805);
nand U2595 (N_2595,N_1215,N_1878);
xnor U2596 (N_2596,N_1662,N_1560);
nand U2597 (N_2597,N_1313,N_1261);
and U2598 (N_2598,N_1806,N_1531);
nand U2599 (N_2599,N_1806,N_1060);
xnor U2600 (N_2600,N_1067,N_1210);
xor U2601 (N_2601,N_1764,N_1066);
nand U2602 (N_2602,N_1860,N_1394);
or U2603 (N_2603,N_1241,N_1552);
nand U2604 (N_2604,N_1531,N_1983);
xnor U2605 (N_2605,N_1841,N_1126);
xor U2606 (N_2606,N_1993,N_1749);
nand U2607 (N_2607,N_1672,N_1786);
or U2608 (N_2608,N_1439,N_1371);
nor U2609 (N_2609,N_1628,N_1721);
xor U2610 (N_2610,N_1986,N_1583);
xor U2611 (N_2611,N_1287,N_1648);
and U2612 (N_2612,N_1655,N_1083);
or U2613 (N_2613,N_1660,N_1248);
and U2614 (N_2614,N_1627,N_1058);
nor U2615 (N_2615,N_1361,N_1677);
nor U2616 (N_2616,N_1207,N_1636);
nand U2617 (N_2617,N_1995,N_1560);
nand U2618 (N_2618,N_1675,N_1294);
xor U2619 (N_2619,N_1774,N_1991);
nand U2620 (N_2620,N_1650,N_1767);
and U2621 (N_2621,N_1577,N_1872);
nand U2622 (N_2622,N_1643,N_1710);
nand U2623 (N_2623,N_1869,N_1470);
nor U2624 (N_2624,N_1736,N_1989);
and U2625 (N_2625,N_1155,N_1178);
nand U2626 (N_2626,N_1130,N_1885);
nor U2627 (N_2627,N_1085,N_1017);
nand U2628 (N_2628,N_1070,N_1170);
nand U2629 (N_2629,N_1275,N_1782);
or U2630 (N_2630,N_1547,N_1488);
xnor U2631 (N_2631,N_1143,N_1710);
nand U2632 (N_2632,N_1918,N_1006);
or U2633 (N_2633,N_1177,N_1033);
and U2634 (N_2634,N_1783,N_1537);
xor U2635 (N_2635,N_1153,N_1374);
xor U2636 (N_2636,N_1149,N_1904);
nand U2637 (N_2637,N_1645,N_1458);
nor U2638 (N_2638,N_1691,N_1210);
xor U2639 (N_2639,N_1212,N_1110);
xor U2640 (N_2640,N_1867,N_1100);
and U2641 (N_2641,N_1279,N_1322);
nor U2642 (N_2642,N_1636,N_1977);
and U2643 (N_2643,N_1014,N_1752);
nand U2644 (N_2644,N_1831,N_1122);
nor U2645 (N_2645,N_1320,N_1902);
or U2646 (N_2646,N_1963,N_1342);
nand U2647 (N_2647,N_1771,N_1723);
nor U2648 (N_2648,N_1337,N_1678);
or U2649 (N_2649,N_1139,N_1213);
and U2650 (N_2650,N_1460,N_1172);
and U2651 (N_2651,N_1726,N_1273);
nor U2652 (N_2652,N_1094,N_1423);
or U2653 (N_2653,N_1737,N_1362);
nor U2654 (N_2654,N_1814,N_1432);
or U2655 (N_2655,N_1364,N_1346);
nor U2656 (N_2656,N_1114,N_1011);
xor U2657 (N_2657,N_1164,N_1760);
nor U2658 (N_2658,N_1288,N_1312);
nand U2659 (N_2659,N_1092,N_1273);
xor U2660 (N_2660,N_1109,N_1214);
or U2661 (N_2661,N_1300,N_1746);
xnor U2662 (N_2662,N_1498,N_1847);
nor U2663 (N_2663,N_1310,N_1822);
xnor U2664 (N_2664,N_1758,N_1678);
xnor U2665 (N_2665,N_1351,N_1467);
xor U2666 (N_2666,N_1488,N_1393);
and U2667 (N_2667,N_1131,N_1597);
or U2668 (N_2668,N_1797,N_1777);
nor U2669 (N_2669,N_1213,N_1581);
nand U2670 (N_2670,N_1362,N_1815);
and U2671 (N_2671,N_1761,N_1888);
nor U2672 (N_2672,N_1507,N_1069);
nand U2673 (N_2673,N_1880,N_1078);
nand U2674 (N_2674,N_1484,N_1136);
or U2675 (N_2675,N_1257,N_1859);
and U2676 (N_2676,N_1436,N_1975);
or U2677 (N_2677,N_1071,N_1076);
nand U2678 (N_2678,N_1330,N_1678);
nand U2679 (N_2679,N_1041,N_1478);
and U2680 (N_2680,N_1058,N_1178);
xor U2681 (N_2681,N_1595,N_1089);
nor U2682 (N_2682,N_1007,N_1999);
nor U2683 (N_2683,N_1864,N_1396);
or U2684 (N_2684,N_1728,N_1774);
nor U2685 (N_2685,N_1998,N_1058);
nor U2686 (N_2686,N_1428,N_1677);
and U2687 (N_2687,N_1319,N_1674);
nand U2688 (N_2688,N_1056,N_1795);
and U2689 (N_2689,N_1801,N_1764);
or U2690 (N_2690,N_1111,N_1241);
nor U2691 (N_2691,N_1040,N_1786);
nand U2692 (N_2692,N_1031,N_1796);
nand U2693 (N_2693,N_1845,N_1129);
xor U2694 (N_2694,N_1105,N_1937);
xnor U2695 (N_2695,N_1838,N_1131);
nand U2696 (N_2696,N_1169,N_1439);
or U2697 (N_2697,N_1561,N_1463);
or U2698 (N_2698,N_1990,N_1858);
xor U2699 (N_2699,N_1691,N_1246);
xor U2700 (N_2700,N_1461,N_1476);
nor U2701 (N_2701,N_1751,N_1661);
nand U2702 (N_2702,N_1379,N_1848);
nand U2703 (N_2703,N_1656,N_1114);
nand U2704 (N_2704,N_1987,N_1870);
nand U2705 (N_2705,N_1797,N_1535);
and U2706 (N_2706,N_1745,N_1909);
nand U2707 (N_2707,N_1642,N_1377);
xor U2708 (N_2708,N_1431,N_1378);
and U2709 (N_2709,N_1406,N_1496);
nand U2710 (N_2710,N_1437,N_1533);
nor U2711 (N_2711,N_1669,N_1359);
nor U2712 (N_2712,N_1276,N_1397);
xor U2713 (N_2713,N_1926,N_1855);
xnor U2714 (N_2714,N_1480,N_1869);
and U2715 (N_2715,N_1794,N_1690);
nor U2716 (N_2716,N_1982,N_1801);
nand U2717 (N_2717,N_1210,N_1520);
and U2718 (N_2718,N_1161,N_1311);
nand U2719 (N_2719,N_1520,N_1738);
xor U2720 (N_2720,N_1541,N_1387);
nor U2721 (N_2721,N_1417,N_1476);
nor U2722 (N_2722,N_1682,N_1430);
or U2723 (N_2723,N_1240,N_1992);
xnor U2724 (N_2724,N_1891,N_1248);
xor U2725 (N_2725,N_1340,N_1758);
nand U2726 (N_2726,N_1825,N_1591);
xnor U2727 (N_2727,N_1215,N_1118);
nand U2728 (N_2728,N_1675,N_1879);
nand U2729 (N_2729,N_1644,N_1803);
nand U2730 (N_2730,N_1714,N_1331);
or U2731 (N_2731,N_1677,N_1287);
and U2732 (N_2732,N_1947,N_1948);
nor U2733 (N_2733,N_1917,N_1963);
nor U2734 (N_2734,N_1157,N_1648);
xor U2735 (N_2735,N_1094,N_1956);
and U2736 (N_2736,N_1088,N_1281);
nor U2737 (N_2737,N_1024,N_1229);
or U2738 (N_2738,N_1328,N_1083);
and U2739 (N_2739,N_1856,N_1328);
nor U2740 (N_2740,N_1194,N_1145);
xnor U2741 (N_2741,N_1418,N_1573);
nand U2742 (N_2742,N_1507,N_1152);
or U2743 (N_2743,N_1002,N_1289);
or U2744 (N_2744,N_1099,N_1274);
nor U2745 (N_2745,N_1992,N_1767);
xnor U2746 (N_2746,N_1652,N_1881);
or U2747 (N_2747,N_1930,N_1201);
and U2748 (N_2748,N_1186,N_1289);
and U2749 (N_2749,N_1399,N_1075);
and U2750 (N_2750,N_1993,N_1495);
or U2751 (N_2751,N_1022,N_1052);
nand U2752 (N_2752,N_1037,N_1953);
nor U2753 (N_2753,N_1175,N_1983);
xor U2754 (N_2754,N_1868,N_1718);
xor U2755 (N_2755,N_1058,N_1800);
and U2756 (N_2756,N_1357,N_1698);
nand U2757 (N_2757,N_1368,N_1413);
xnor U2758 (N_2758,N_1598,N_1261);
or U2759 (N_2759,N_1969,N_1233);
or U2760 (N_2760,N_1751,N_1368);
or U2761 (N_2761,N_1060,N_1247);
and U2762 (N_2762,N_1173,N_1605);
xor U2763 (N_2763,N_1024,N_1227);
nor U2764 (N_2764,N_1266,N_1909);
or U2765 (N_2765,N_1542,N_1239);
xnor U2766 (N_2766,N_1805,N_1073);
and U2767 (N_2767,N_1383,N_1433);
xnor U2768 (N_2768,N_1028,N_1328);
nand U2769 (N_2769,N_1809,N_1047);
xnor U2770 (N_2770,N_1091,N_1023);
or U2771 (N_2771,N_1596,N_1358);
and U2772 (N_2772,N_1952,N_1887);
xor U2773 (N_2773,N_1678,N_1791);
xnor U2774 (N_2774,N_1556,N_1906);
or U2775 (N_2775,N_1412,N_1351);
nand U2776 (N_2776,N_1606,N_1368);
xnor U2777 (N_2777,N_1718,N_1631);
nand U2778 (N_2778,N_1001,N_1725);
nor U2779 (N_2779,N_1237,N_1123);
nor U2780 (N_2780,N_1724,N_1717);
or U2781 (N_2781,N_1006,N_1175);
or U2782 (N_2782,N_1538,N_1040);
or U2783 (N_2783,N_1980,N_1078);
and U2784 (N_2784,N_1288,N_1871);
and U2785 (N_2785,N_1393,N_1240);
nand U2786 (N_2786,N_1191,N_1952);
xnor U2787 (N_2787,N_1609,N_1203);
or U2788 (N_2788,N_1920,N_1685);
and U2789 (N_2789,N_1109,N_1296);
xor U2790 (N_2790,N_1609,N_1410);
xor U2791 (N_2791,N_1223,N_1571);
or U2792 (N_2792,N_1268,N_1624);
nor U2793 (N_2793,N_1615,N_1944);
nor U2794 (N_2794,N_1779,N_1879);
or U2795 (N_2795,N_1494,N_1803);
or U2796 (N_2796,N_1403,N_1786);
and U2797 (N_2797,N_1487,N_1026);
xnor U2798 (N_2798,N_1566,N_1992);
nor U2799 (N_2799,N_1364,N_1370);
or U2800 (N_2800,N_1095,N_1279);
nand U2801 (N_2801,N_1584,N_1781);
nand U2802 (N_2802,N_1528,N_1568);
and U2803 (N_2803,N_1338,N_1871);
and U2804 (N_2804,N_1549,N_1878);
nor U2805 (N_2805,N_1515,N_1958);
nor U2806 (N_2806,N_1847,N_1826);
nor U2807 (N_2807,N_1512,N_1839);
xnor U2808 (N_2808,N_1710,N_1116);
and U2809 (N_2809,N_1806,N_1506);
xor U2810 (N_2810,N_1120,N_1194);
or U2811 (N_2811,N_1049,N_1250);
nor U2812 (N_2812,N_1617,N_1312);
and U2813 (N_2813,N_1713,N_1736);
and U2814 (N_2814,N_1948,N_1343);
nor U2815 (N_2815,N_1948,N_1852);
nand U2816 (N_2816,N_1202,N_1050);
or U2817 (N_2817,N_1235,N_1633);
and U2818 (N_2818,N_1291,N_1388);
xnor U2819 (N_2819,N_1292,N_1859);
and U2820 (N_2820,N_1094,N_1957);
xor U2821 (N_2821,N_1680,N_1260);
nand U2822 (N_2822,N_1971,N_1789);
or U2823 (N_2823,N_1315,N_1945);
and U2824 (N_2824,N_1786,N_1359);
xor U2825 (N_2825,N_1388,N_1767);
nand U2826 (N_2826,N_1015,N_1388);
nor U2827 (N_2827,N_1646,N_1232);
or U2828 (N_2828,N_1780,N_1296);
and U2829 (N_2829,N_1978,N_1436);
nand U2830 (N_2830,N_1330,N_1340);
nand U2831 (N_2831,N_1192,N_1429);
nor U2832 (N_2832,N_1264,N_1152);
or U2833 (N_2833,N_1298,N_1999);
nor U2834 (N_2834,N_1220,N_1500);
nand U2835 (N_2835,N_1217,N_1456);
or U2836 (N_2836,N_1112,N_1012);
or U2837 (N_2837,N_1328,N_1811);
nand U2838 (N_2838,N_1744,N_1552);
nor U2839 (N_2839,N_1183,N_1784);
and U2840 (N_2840,N_1252,N_1746);
xor U2841 (N_2841,N_1444,N_1580);
nor U2842 (N_2842,N_1295,N_1519);
and U2843 (N_2843,N_1260,N_1265);
nor U2844 (N_2844,N_1329,N_1704);
and U2845 (N_2845,N_1216,N_1073);
xnor U2846 (N_2846,N_1454,N_1781);
nor U2847 (N_2847,N_1499,N_1575);
xor U2848 (N_2848,N_1870,N_1437);
nand U2849 (N_2849,N_1305,N_1513);
and U2850 (N_2850,N_1894,N_1832);
nand U2851 (N_2851,N_1005,N_1594);
xnor U2852 (N_2852,N_1518,N_1703);
or U2853 (N_2853,N_1420,N_1945);
or U2854 (N_2854,N_1790,N_1327);
xor U2855 (N_2855,N_1414,N_1316);
or U2856 (N_2856,N_1134,N_1274);
and U2857 (N_2857,N_1878,N_1551);
and U2858 (N_2858,N_1183,N_1133);
nand U2859 (N_2859,N_1959,N_1281);
and U2860 (N_2860,N_1642,N_1583);
nor U2861 (N_2861,N_1689,N_1778);
or U2862 (N_2862,N_1271,N_1288);
xnor U2863 (N_2863,N_1442,N_1437);
nor U2864 (N_2864,N_1566,N_1450);
xor U2865 (N_2865,N_1845,N_1758);
or U2866 (N_2866,N_1252,N_1631);
nand U2867 (N_2867,N_1306,N_1541);
and U2868 (N_2868,N_1860,N_1050);
nand U2869 (N_2869,N_1815,N_1360);
or U2870 (N_2870,N_1993,N_1471);
and U2871 (N_2871,N_1170,N_1220);
nand U2872 (N_2872,N_1857,N_1180);
and U2873 (N_2873,N_1181,N_1248);
nand U2874 (N_2874,N_1366,N_1743);
xnor U2875 (N_2875,N_1716,N_1890);
nand U2876 (N_2876,N_1098,N_1184);
nand U2877 (N_2877,N_1991,N_1791);
nor U2878 (N_2878,N_1405,N_1406);
and U2879 (N_2879,N_1473,N_1461);
xor U2880 (N_2880,N_1455,N_1111);
and U2881 (N_2881,N_1227,N_1239);
xnor U2882 (N_2882,N_1794,N_1830);
xor U2883 (N_2883,N_1572,N_1403);
nand U2884 (N_2884,N_1417,N_1204);
nand U2885 (N_2885,N_1094,N_1864);
and U2886 (N_2886,N_1961,N_1498);
xnor U2887 (N_2887,N_1712,N_1187);
nand U2888 (N_2888,N_1893,N_1959);
nand U2889 (N_2889,N_1674,N_1944);
xor U2890 (N_2890,N_1646,N_1850);
and U2891 (N_2891,N_1545,N_1531);
nand U2892 (N_2892,N_1293,N_1515);
nor U2893 (N_2893,N_1375,N_1827);
xor U2894 (N_2894,N_1808,N_1310);
or U2895 (N_2895,N_1083,N_1204);
or U2896 (N_2896,N_1944,N_1010);
and U2897 (N_2897,N_1886,N_1913);
or U2898 (N_2898,N_1478,N_1785);
and U2899 (N_2899,N_1347,N_1512);
nand U2900 (N_2900,N_1503,N_1184);
or U2901 (N_2901,N_1317,N_1168);
nand U2902 (N_2902,N_1520,N_1112);
or U2903 (N_2903,N_1393,N_1437);
nand U2904 (N_2904,N_1170,N_1288);
or U2905 (N_2905,N_1797,N_1384);
nand U2906 (N_2906,N_1487,N_1237);
nor U2907 (N_2907,N_1047,N_1298);
or U2908 (N_2908,N_1131,N_1601);
xor U2909 (N_2909,N_1207,N_1597);
nor U2910 (N_2910,N_1943,N_1419);
nor U2911 (N_2911,N_1087,N_1217);
or U2912 (N_2912,N_1792,N_1963);
nor U2913 (N_2913,N_1111,N_1042);
nand U2914 (N_2914,N_1650,N_1471);
nand U2915 (N_2915,N_1710,N_1751);
xnor U2916 (N_2916,N_1020,N_1321);
xor U2917 (N_2917,N_1522,N_1119);
and U2918 (N_2918,N_1558,N_1342);
nand U2919 (N_2919,N_1919,N_1453);
and U2920 (N_2920,N_1221,N_1680);
and U2921 (N_2921,N_1990,N_1206);
nor U2922 (N_2922,N_1835,N_1681);
xnor U2923 (N_2923,N_1348,N_1666);
and U2924 (N_2924,N_1721,N_1757);
or U2925 (N_2925,N_1206,N_1063);
xor U2926 (N_2926,N_1164,N_1819);
xnor U2927 (N_2927,N_1113,N_1278);
nand U2928 (N_2928,N_1861,N_1880);
or U2929 (N_2929,N_1339,N_1513);
nand U2930 (N_2930,N_1722,N_1395);
nand U2931 (N_2931,N_1178,N_1832);
xnor U2932 (N_2932,N_1849,N_1893);
or U2933 (N_2933,N_1316,N_1175);
and U2934 (N_2934,N_1265,N_1053);
and U2935 (N_2935,N_1035,N_1207);
xnor U2936 (N_2936,N_1532,N_1269);
xnor U2937 (N_2937,N_1807,N_1107);
nor U2938 (N_2938,N_1198,N_1586);
or U2939 (N_2939,N_1154,N_1099);
nand U2940 (N_2940,N_1581,N_1687);
or U2941 (N_2941,N_1958,N_1534);
and U2942 (N_2942,N_1115,N_1918);
nor U2943 (N_2943,N_1364,N_1671);
nor U2944 (N_2944,N_1708,N_1220);
or U2945 (N_2945,N_1511,N_1531);
nor U2946 (N_2946,N_1632,N_1587);
and U2947 (N_2947,N_1773,N_1435);
nor U2948 (N_2948,N_1683,N_1147);
nor U2949 (N_2949,N_1067,N_1879);
and U2950 (N_2950,N_1447,N_1483);
and U2951 (N_2951,N_1634,N_1529);
nand U2952 (N_2952,N_1689,N_1823);
and U2953 (N_2953,N_1905,N_1647);
and U2954 (N_2954,N_1926,N_1556);
nor U2955 (N_2955,N_1107,N_1922);
nor U2956 (N_2956,N_1159,N_1223);
xor U2957 (N_2957,N_1182,N_1456);
xnor U2958 (N_2958,N_1808,N_1558);
nor U2959 (N_2959,N_1279,N_1646);
nand U2960 (N_2960,N_1691,N_1896);
nand U2961 (N_2961,N_1905,N_1773);
and U2962 (N_2962,N_1725,N_1138);
nor U2963 (N_2963,N_1610,N_1702);
nor U2964 (N_2964,N_1306,N_1566);
and U2965 (N_2965,N_1617,N_1474);
or U2966 (N_2966,N_1071,N_1619);
or U2967 (N_2967,N_1069,N_1149);
or U2968 (N_2968,N_1044,N_1417);
nand U2969 (N_2969,N_1768,N_1170);
nand U2970 (N_2970,N_1649,N_1377);
nor U2971 (N_2971,N_1749,N_1801);
and U2972 (N_2972,N_1112,N_1535);
or U2973 (N_2973,N_1070,N_1296);
and U2974 (N_2974,N_1080,N_1924);
nand U2975 (N_2975,N_1408,N_1102);
or U2976 (N_2976,N_1291,N_1743);
and U2977 (N_2977,N_1986,N_1586);
nand U2978 (N_2978,N_1006,N_1626);
nand U2979 (N_2979,N_1238,N_1514);
nor U2980 (N_2980,N_1790,N_1611);
xor U2981 (N_2981,N_1409,N_1657);
nor U2982 (N_2982,N_1211,N_1464);
or U2983 (N_2983,N_1686,N_1345);
or U2984 (N_2984,N_1750,N_1628);
nor U2985 (N_2985,N_1464,N_1601);
and U2986 (N_2986,N_1187,N_1757);
xor U2987 (N_2987,N_1530,N_1895);
or U2988 (N_2988,N_1620,N_1256);
xnor U2989 (N_2989,N_1089,N_1730);
nand U2990 (N_2990,N_1185,N_1967);
xnor U2991 (N_2991,N_1285,N_1421);
or U2992 (N_2992,N_1202,N_1963);
nor U2993 (N_2993,N_1189,N_1503);
or U2994 (N_2994,N_1201,N_1736);
or U2995 (N_2995,N_1716,N_1585);
and U2996 (N_2996,N_1212,N_1728);
or U2997 (N_2997,N_1101,N_1644);
nor U2998 (N_2998,N_1108,N_1195);
nand U2999 (N_2999,N_1068,N_1866);
and U3000 (N_3000,N_2077,N_2438);
or U3001 (N_3001,N_2984,N_2141);
or U3002 (N_3002,N_2181,N_2944);
xor U3003 (N_3003,N_2857,N_2090);
or U3004 (N_3004,N_2232,N_2377);
nor U3005 (N_3005,N_2201,N_2165);
nor U3006 (N_3006,N_2818,N_2981);
xor U3007 (N_3007,N_2954,N_2744);
xor U3008 (N_3008,N_2621,N_2599);
or U3009 (N_3009,N_2014,N_2992);
or U3010 (N_3010,N_2749,N_2295);
and U3011 (N_3011,N_2568,N_2159);
nand U3012 (N_3012,N_2203,N_2590);
and U3013 (N_3013,N_2890,N_2188);
and U3014 (N_3014,N_2307,N_2782);
or U3015 (N_3015,N_2584,N_2688);
and U3016 (N_3016,N_2551,N_2013);
nand U3017 (N_3017,N_2597,N_2069);
xor U3018 (N_3018,N_2790,N_2375);
xnor U3019 (N_3019,N_2518,N_2112);
or U3020 (N_3020,N_2988,N_2824);
nand U3021 (N_3021,N_2022,N_2448);
and U3022 (N_3022,N_2481,N_2389);
nand U3023 (N_3023,N_2755,N_2603);
or U3024 (N_3024,N_2690,N_2631);
or U3025 (N_3025,N_2106,N_2542);
and U3026 (N_3026,N_2015,N_2155);
nand U3027 (N_3027,N_2003,N_2460);
and U3028 (N_3028,N_2239,N_2170);
nand U3029 (N_3029,N_2140,N_2515);
nand U3030 (N_3030,N_2317,N_2735);
and U3031 (N_3031,N_2175,N_2540);
xnor U3032 (N_3032,N_2932,N_2523);
or U3033 (N_3033,N_2913,N_2645);
nor U3034 (N_3034,N_2330,N_2017);
nand U3035 (N_3035,N_2624,N_2355);
xnor U3036 (N_3036,N_2304,N_2573);
nor U3037 (N_3037,N_2452,N_2627);
nand U3038 (N_3038,N_2537,N_2467);
nor U3039 (N_3039,N_2176,N_2081);
and U3040 (N_3040,N_2608,N_2921);
nor U3041 (N_3041,N_2530,N_2810);
nor U3042 (N_3042,N_2426,N_2216);
nor U3043 (N_3043,N_2822,N_2907);
nor U3044 (N_3044,N_2235,N_2629);
and U3045 (N_3045,N_2787,N_2403);
or U3046 (N_3046,N_2137,N_2314);
and U3047 (N_3047,N_2492,N_2634);
or U3048 (N_3048,N_2157,N_2870);
nand U3049 (N_3049,N_2335,N_2699);
nand U3050 (N_3050,N_2485,N_2423);
xor U3051 (N_3051,N_2497,N_2948);
nor U3052 (N_3052,N_2612,N_2343);
nand U3053 (N_3053,N_2904,N_2398);
xnor U3054 (N_3054,N_2328,N_2059);
nor U3055 (N_3055,N_2421,N_2034);
or U3056 (N_3056,N_2290,N_2287);
and U3057 (N_3057,N_2873,N_2943);
and U3058 (N_3058,N_2206,N_2358);
nand U3059 (N_3059,N_2698,N_2173);
or U3060 (N_3060,N_2115,N_2142);
xor U3061 (N_3061,N_2231,N_2549);
or U3062 (N_3062,N_2225,N_2522);
nor U3063 (N_3063,N_2102,N_2051);
xnor U3064 (N_3064,N_2779,N_2359);
nor U3065 (N_3065,N_2025,N_2647);
nand U3066 (N_3066,N_2630,N_2935);
nor U3067 (N_3067,N_2606,N_2392);
and U3068 (N_3068,N_2985,N_2361);
xor U3069 (N_3069,N_2980,N_2575);
nand U3070 (N_3070,N_2498,N_2710);
nor U3071 (N_3071,N_2427,N_2461);
nand U3072 (N_3072,N_2605,N_2373);
or U3073 (N_3073,N_2739,N_2070);
xnor U3074 (N_3074,N_2192,N_2742);
nor U3075 (N_3075,N_2660,N_2591);
nor U3076 (N_3076,N_2886,N_2973);
nand U3077 (N_3077,N_2585,N_2846);
or U3078 (N_3078,N_2422,N_2390);
and U3079 (N_3079,N_2505,N_2026);
and U3080 (N_3080,N_2833,N_2502);
nor U3081 (N_3081,N_2082,N_2756);
and U3082 (N_3082,N_2765,N_2995);
xor U3083 (N_3083,N_2487,N_2270);
nor U3084 (N_3084,N_2848,N_2190);
and U3085 (N_3085,N_2120,N_2956);
nand U3086 (N_3086,N_2587,N_2951);
nor U3087 (N_3087,N_2391,N_2506);
nor U3088 (N_3088,N_2387,N_2257);
and U3089 (N_3089,N_2879,N_2686);
nor U3090 (N_3090,N_2182,N_2702);
and U3091 (N_3091,N_2649,N_2315);
or U3092 (N_3092,N_2805,N_2644);
nand U3093 (N_3093,N_2926,N_2741);
and U3094 (N_3094,N_2029,N_2915);
and U3095 (N_3095,N_2899,N_2352);
nor U3096 (N_3096,N_2854,N_2967);
xnor U3097 (N_3097,N_2908,N_2039);
or U3098 (N_3098,N_2310,N_2404);
nand U3099 (N_3099,N_2222,N_2852);
or U3100 (N_3100,N_2368,N_2507);
or U3101 (N_3101,N_2910,N_2708);
xor U3102 (N_3102,N_2097,N_2292);
xor U3103 (N_3103,N_2254,N_2047);
or U3104 (N_3104,N_2085,N_2817);
nand U3105 (N_3105,N_2503,N_2925);
and U3106 (N_3106,N_2436,N_2867);
nor U3107 (N_3107,N_2840,N_2723);
or U3108 (N_3108,N_2950,N_2652);
xor U3109 (N_3109,N_2750,N_2774);
or U3110 (N_3110,N_2128,N_2564);
xor U3111 (N_3111,N_2882,N_2199);
nor U3112 (N_3112,N_2078,N_2341);
xor U3113 (N_3113,N_2999,N_2863);
and U3114 (N_3114,N_2156,N_2707);
nand U3115 (N_3115,N_2813,N_2303);
xor U3116 (N_3116,N_2826,N_2562);
and U3117 (N_3117,N_2246,N_2855);
or U3118 (N_3118,N_2365,N_2345);
and U3119 (N_3119,N_2145,N_2832);
or U3120 (N_3120,N_2903,N_2093);
nand U3121 (N_3121,N_2496,N_2226);
or U3122 (N_3122,N_2306,N_2610);
nand U3123 (N_3123,N_2527,N_2208);
or U3124 (N_3124,N_2125,N_2844);
and U3125 (N_3125,N_2348,N_2781);
nor U3126 (N_3126,N_2010,N_2062);
or U3127 (N_3127,N_2209,N_2185);
nor U3128 (N_3128,N_2520,N_2350);
and U3129 (N_3129,N_2119,N_2320);
nor U3130 (N_3130,N_2374,N_2730);
and U3131 (N_3131,N_2732,N_2224);
nor U3132 (N_3132,N_2117,N_2695);
and U3133 (N_3133,N_2743,N_2458);
xnor U3134 (N_3134,N_2964,N_2800);
or U3135 (N_3135,N_2114,N_2005);
xor U3136 (N_3136,N_2476,N_2164);
nor U3137 (N_3137,N_2417,N_2693);
or U3138 (N_3138,N_2576,N_2061);
nor U3139 (N_3139,N_2234,N_2463);
nand U3140 (N_3140,N_2200,N_2275);
or U3141 (N_3141,N_2768,N_2689);
nand U3142 (N_3142,N_2640,N_2443);
xor U3143 (N_3143,N_2979,N_2843);
nor U3144 (N_3144,N_2475,N_2472);
and U3145 (N_3145,N_2439,N_2301);
nand U3146 (N_3146,N_2991,N_2966);
nor U3147 (N_3147,N_2433,N_2938);
and U3148 (N_3148,N_2842,N_2703);
xnor U3149 (N_3149,N_2032,N_2207);
nand U3150 (N_3150,N_2037,N_2351);
nand U3151 (N_3151,N_2313,N_2924);
xor U3152 (N_3152,N_2018,N_2311);
nand U3153 (N_3153,N_2623,N_2717);
xor U3154 (N_3154,N_2508,N_2495);
xnor U3155 (N_3155,N_2602,N_2801);
or U3156 (N_3156,N_2588,N_2579);
and U3157 (N_3157,N_2978,N_2428);
and U3158 (N_3158,N_2278,N_2401);
or U3159 (N_3159,N_2521,N_2212);
and U3160 (N_3160,N_2131,N_2148);
nand U3161 (N_3161,N_2001,N_2135);
xor U3162 (N_3162,N_2132,N_2468);
or U3163 (N_3163,N_2546,N_2811);
nand U3164 (N_3164,N_2223,N_2764);
or U3165 (N_3165,N_2912,N_2930);
xor U3166 (N_3166,N_2796,N_2514);
xnor U3167 (N_3167,N_2883,N_2963);
and U3168 (N_3168,N_2598,N_2154);
nand U3169 (N_3169,N_2543,N_2663);
xnor U3170 (N_3170,N_2655,N_2672);
xor U3171 (N_3171,N_2607,N_2366);
or U3172 (N_3172,N_2676,N_2260);
nor U3173 (N_3173,N_2038,N_2785);
and U3174 (N_3174,N_2035,N_2734);
nand U3175 (N_3175,N_2477,N_2880);
xnor U3176 (N_3176,N_2194,N_2720);
nor U3177 (N_3177,N_2211,N_2828);
xor U3178 (N_3178,N_2681,N_2715);
nand U3179 (N_3179,N_2776,N_2339);
nor U3180 (N_3180,N_2751,N_2473);
nand U3181 (N_3181,N_2923,N_2936);
or U3182 (N_3182,N_2968,N_2264);
nand U3183 (N_3183,N_2321,N_2240);
xor U3184 (N_3184,N_2806,N_2529);
nor U3185 (N_3185,N_2896,N_2258);
nand U3186 (N_3186,N_2803,N_2658);
nor U3187 (N_3187,N_2040,N_2011);
and U3188 (N_3188,N_2583,N_2383);
or U3189 (N_3189,N_2911,N_2107);
nor U3190 (N_3190,N_2673,N_2074);
nand U3191 (N_3191,N_2356,N_2594);
and U3192 (N_3192,N_2332,N_2233);
xor U3193 (N_3193,N_2493,N_2531);
nor U3194 (N_3194,N_2198,N_2108);
nand U3195 (N_3195,N_2094,N_2110);
and U3196 (N_3196,N_2685,N_2550);
nand U3197 (N_3197,N_2628,N_2657);
or U3198 (N_3198,N_2816,N_2241);
nand U3199 (N_3199,N_2259,N_2449);
nand U3200 (N_3200,N_2380,N_2101);
and U3201 (N_3201,N_2126,N_2395);
nor U3202 (N_3202,N_2553,N_2087);
or U3203 (N_3203,N_2354,N_2318);
and U3204 (N_3204,N_2268,N_2041);
xnor U3205 (N_3205,N_2626,N_2280);
xnor U3206 (N_3206,N_2186,N_2180);
xnor U3207 (N_3207,N_2152,N_2281);
nor U3208 (N_3208,N_2976,N_2856);
and U3209 (N_3209,N_2788,N_2946);
and U3210 (N_3210,N_2949,N_2648);
or U3211 (N_3211,N_2678,N_2456);
xor U3212 (N_3212,N_2016,N_2794);
nor U3213 (N_3213,N_2319,N_2396);
and U3214 (N_3214,N_2592,N_2308);
and U3215 (N_3215,N_2197,N_2172);
nor U3216 (N_3216,N_2958,N_2369);
nand U3217 (N_3217,N_2277,N_2641);
xor U3218 (N_3218,N_2725,N_2849);
and U3219 (N_3219,N_2048,N_2600);
xor U3220 (N_3220,N_2722,N_2033);
or U3221 (N_3221,N_2272,N_2651);
or U3222 (N_3222,N_2429,N_2837);
and U3223 (N_3223,N_2334,N_2885);
nor U3224 (N_3224,N_2831,N_2793);
or U3225 (N_3225,N_2009,N_2916);
and U3226 (N_3226,N_2002,N_2312);
nand U3227 (N_3227,N_2664,N_2215);
or U3228 (N_3228,N_2073,N_2763);
xnor U3229 (N_3229,N_2454,N_2299);
xor U3230 (N_3230,N_2884,N_2163);
nand U3231 (N_3231,N_2516,N_2970);
or U3232 (N_3232,N_2525,N_2929);
nand U3233 (N_3233,N_2245,N_2044);
nand U3234 (N_3234,N_2187,N_2242);
or U3235 (N_3235,N_2006,N_2795);
nand U3236 (N_3236,N_2563,N_2758);
or U3237 (N_3237,N_2213,N_2363);
nand U3238 (N_3238,N_2571,N_2736);
xor U3239 (N_3239,N_2284,N_2836);
nand U3240 (N_3240,N_2791,N_2559);
and U3241 (N_3241,N_2441,N_2451);
or U3242 (N_3242,N_2920,N_2298);
nor U3243 (N_3243,N_2166,N_2953);
or U3244 (N_3244,N_2065,N_2323);
or U3245 (N_3245,N_2766,N_2344);
and U3246 (N_3246,N_2174,N_2668);
and U3247 (N_3247,N_2305,N_2850);
xor U3248 (N_3248,N_2545,N_2394);
nor U3249 (N_3249,N_2459,N_2705);
and U3250 (N_3250,N_2068,N_2536);
xor U3251 (N_3251,N_2731,N_2060);
xnor U3252 (N_3252,N_2614,N_2079);
nor U3253 (N_3253,N_2983,N_2748);
nor U3254 (N_3254,N_2021,N_2269);
and U3255 (N_3255,N_2729,N_2711);
xnor U3256 (N_3256,N_2121,N_2990);
or U3257 (N_3257,N_2236,N_2043);
nand U3258 (N_3258,N_2092,N_2214);
or U3259 (N_3259,N_2918,N_2020);
nor U3260 (N_3260,N_2414,N_2229);
nand U3261 (N_3261,N_2113,N_2362);
nor U3262 (N_3262,N_2595,N_2249);
nor U3263 (N_3263,N_2679,N_2397);
and U3264 (N_3264,N_2385,N_2819);
nand U3265 (N_3265,N_2195,N_2388);
nor U3266 (N_3266,N_2478,N_2757);
or U3267 (N_3267,N_2581,N_2063);
and U3268 (N_3268,N_2099,N_2682);
nor U3269 (N_3269,N_2453,N_2419);
nand U3270 (N_3270,N_2513,N_2760);
or U3271 (N_3271,N_2875,N_2871);
nand U3272 (N_3272,N_2567,N_2490);
nor U3273 (N_3273,N_2815,N_2480);
or U3274 (N_3274,N_2372,N_2248);
xor U3275 (N_3275,N_2302,N_2000);
nand U3276 (N_3276,N_2639,N_2338);
xnor U3277 (N_3277,N_2413,N_2609);
or U3278 (N_3278,N_2894,N_2792);
nor U3279 (N_3279,N_2799,N_2718);
nand U3280 (N_3280,N_2130,N_2075);
nand U3281 (N_3281,N_2704,N_2965);
or U3282 (N_3282,N_2998,N_2928);
nor U3283 (N_3283,N_2619,N_2820);
nor U3284 (N_3284,N_2694,N_2737);
xnor U3285 (N_3285,N_2892,N_2408);
nand U3286 (N_3286,N_2118,N_2738);
nand U3287 (N_3287,N_2726,N_2510);
nand U3288 (N_3288,N_2191,N_2556);
or U3289 (N_3289,N_2777,N_2960);
nand U3290 (N_3290,N_2469,N_2582);
nor U3291 (N_3291,N_2905,N_2642);
or U3292 (N_3292,N_2489,N_2210);
nand U3293 (N_3293,N_2237,N_2446);
xor U3294 (N_3294,N_2346,N_2888);
xor U3295 (N_3295,N_2127,N_2019);
nand U3296 (N_3296,N_2504,N_2656);
nand U3297 (N_3297,N_2218,N_2294);
nor U3298 (N_3298,N_2544,N_2784);
nor U3299 (N_3299,N_2716,N_2895);
or U3300 (N_3300,N_2430,N_2378);
or U3301 (N_3301,N_2511,N_2901);
xor U3302 (N_3302,N_2296,N_2752);
or U3303 (N_3303,N_2045,N_2116);
nor U3304 (N_3304,N_2286,N_2570);
or U3305 (N_3305,N_2067,N_2547);
nor U3306 (N_3306,N_2560,N_2667);
nand U3307 (N_3307,N_2728,N_2691);
or U3308 (N_3308,N_2031,N_2144);
nor U3309 (N_3309,N_2007,N_2227);
xnor U3310 (N_3310,N_2578,N_2219);
or U3311 (N_3311,N_2786,N_2465);
or U3312 (N_3312,N_2196,N_2534);
xor U3313 (N_3313,N_2517,N_2637);
nand U3314 (N_3314,N_2812,N_2569);
nand U3315 (N_3315,N_2986,N_2593);
and U3316 (N_3316,N_2959,N_2288);
and U3317 (N_3317,N_2424,N_2555);
or U3318 (N_3318,N_2941,N_2162);
and U3319 (N_3319,N_2376,N_2046);
nand U3320 (N_3320,N_2080,N_2807);
xnor U3321 (N_3321,N_2860,N_2158);
and U3322 (N_3322,N_2088,N_2989);
nand U3323 (N_3323,N_2474,N_2384);
nand U3324 (N_3324,N_2701,N_2444);
and U3325 (N_3325,N_2221,N_2266);
xor U3326 (N_3326,N_2431,N_2761);
nor U3327 (N_3327,N_2975,N_2122);
nand U3328 (N_3328,N_2399,N_2851);
or U3329 (N_3329,N_2798,N_2541);
nor U3330 (N_3330,N_2036,N_2412);
and U3331 (N_3331,N_2675,N_2434);
nand U3332 (N_3332,N_2974,N_2909);
nor U3333 (N_3333,N_2084,N_2111);
and U3334 (N_3334,N_2494,N_2053);
and U3335 (N_3335,N_2291,N_2276);
or U3336 (N_3336,N_2572,N_2835);
and U3337 (N_3337,N_2753,N_2382);
and U3338 (N_3338,N_2872,N_2643);
nand U3339 (N_3339,N_2055,N_2866);
nor U3340 (N_3340,N_2309,N_2861);
xnor U3341 (N_3341,N_2220,N_2838);
xnor U3342 (N_3342,N_2149,N_2184);
nand U3343 (N_3343,N_2435,N_2906);
and U3344 (N_3344,N_2865,N_2405);
nand U3345 (N_3345,N_2406,N_2635);
nor U3346 (N_3346,N_2706,N_2049);
or U3347 (N_3347,N_2680,N_2877);
or U3348 (N_3348,N_2747,N_2847);
nor U3349 (N_3349,N_2322,N_2178);
nand U3350 (N_3350,N_2876,N_2654);
and U3351 (N_3351,N_2153,N_2586);
xor U3352 (N_3352,N_2931,N_2252);
or U3353 (N_3353,N_2420,N_2283);
xnor U3354 (N_3354,N_2827,N_2804);
xor U3355 (N_3355,N_2379,N_2971);
xnor U3356 (N_3356,N_2289,N_2071);
or U3357 (N_3357,N_2917,N_2274);
xor U3358 (N_3358,N_2267,N_2169);
or U3359 (N_3359,N_2927,N_2409);
and U3360 (N_3360,N_2168,N_2066);
xor U3361 (N_3361,N_2808,N_2393);
xnor U3362 (N_3362,N_2650,N_2618);
and U3363 (N_3363,N_2724,N_2324);
xnor U3364 (N_3364,N_2633,N_2615);
xnor U3365 (N_3365,N_2228,N_2823);
and U3366 (N_3366,N_2004,N_2410);
xnor U3367 (N_3367,N_2416,N_2133);
xnor U3368 (N_3368,N_2042,N_2919);
xnor U3369 (N_3369,N_2349,N_2889);
xor U3370 (N_3370,N_2740,N_2969);
and U3371 (N_3371,N_2887,N_2342);
and U3372 (N_3372,N_2357,N_2337);
nand U3373 (N_3373,N_2447,N_2329);
or U3374 (N_3374,N_2577,N_2440);
and U3375 (N_3375,N_2509,N_2136);
and U3376 (N_3376,N_2402,N_2947);
xor U3377 (N_3377,N_2669,N_2217);
and U3378 (N_3378,N_2364,N_2072);
nor U3379 (N_3379,N_2205,N_2483);
xnor U3380 (N_3380,N_2557,N_2662);
or U3381 (N_3381,N_2432,N_2809);
nand U3382 (N_3382,N_2881,N_2962);
xnor U3383 (N_3383,N_2386,N_2625);
or U3384 (N_3384,N_2437,N_2745);
xnor U3385 (N_3385,N_2442,N_2052);
nor U3386 (N_3386,N_2982,N_2620);
and U3387 (N_3387,N_2780,N_2891);
nor U3388 (N_3388,N_2407,N_2054);
nor U3389 (N_3389,N_2367,N_2957);
and U3390 (N_3390,N_2255,N_2696);
and U3391 (N_3391,N_2008,N_2940);
or U3392 (N_3392,N_2105,N_2251);
nor U3393 (N_3393,N_2499,N_2589);
nand U3394 (N_3394,N_2580,N_2922);
xor U3395 (N_3395,N_2353,N_2727);
or U3396 (N_3396,N_2138,N_2874);
nor U3397 (N_3397,N_2955,N_2261);
or U3398 (N_3398,N_2189,N_2646);
nor U3399 (N_3399,N_2900,N_2400);
or U3400 (N_3400,N_2653,N_2746);
nand U3401 (N_3401,N_2134,N_2665);
or U3402 (N_3402,N_2972,N_2772);
or U3403 (N_3403,N_2622,N_2247);
nor U3404 (N_3404,N_2825,N_2554);
nand U3405 (N_3405,N_2297,N_2023);
and U3406 (N_3406,N_2347,N_2450);
nor U3407 (N_3407,N_2095,N_2566);
or U3408 (N_3408,N_2933,N_2789);
xor U3409 (N_3409,N_2762,N_2057);
xnor U3410 (N_3410,N_2096,N_2243);
nand U3411 (N_3411,N_2687,N_2491);
nor U3412 (N_3412,N_2488,N_2336);
nor U3413 (N_3413,N_2845,N_2325);
or U3414 (N_3414,N_2370,N_2230);
nand U3415 (N_3415,N_2611,N_2331);
or U3416 (N_3416,N_2411,N_2617);
nor U3417 (N_3417,N_2471,N_2869);
xnor U3418 (N_3418,N_2129,N_2661);
xnor U3419 (N_3419,N_2538,N_2482);
and U3420 (N_3420,N_2455,N_2512);
and U3421 (N_3421,N_2632,N_2671);
nor U3422 (N_3422,N_2193,N_2853);
or U3423 (N_3423,N_2552,N_2273);
and U3424 (N_3424,N_2942,N_2802);
or U3425 (N_3425,N_2778,N_2697);
and U3426 (N_3426,N_2937,N_2300);
and U3427 (N_3427,N_2479,N_2714);
and U3428 (N_3428,N_2770,N_2466);
xor U3429 (N_3429,N_2532,N_2028);
nand U3430 (N_3430,N_2841,N_2445);
xor U3431 (N_3431,N_2558,N_2076);
nand U3432 (N_3432,N_2056,N_2997);
nand U3433 (N_3433,N_2179,N_2457);
and U3434 (N_3434,N_2098,N_2548);
and U3435 (N_3435,N_2202,N_2464);
nand U3436 (N_3436,N_2151,N_2616);
xor U3437 (N_3437,N_2265,N_2183);
and U3438 (N_3438,N_2700,N_2027);
and U3439 (N_3439,N_2058,N_2994);
nor U3440 (N_3440,N_2147,N_2719);
xor U3441 (N_3441,N_2143,N_2271);
nand U3442 (N_3442,N_2316,N_2987);
and U3443 (N_3443,N_2462,N_2238);
and U3444 (N_3444,N_2326,N_2961);
and U3445 (N_3445,N_2500,N_2683);
nor U3446 (N_3446,N_2371,N_2425);
and U3447 (N_3447,N_2160,N_2996);
or U3448 (N_3448,N_2759,N_2692);
or U3449 (N_3449,N_2528,N_2898);
nor U3450 (N_3450,N_2109,N_2327);
and U3451 (N_3451,N_2263,N_2821);
and U3452 (N_3452,N_2754,N_2333);
nor U3453 (N_3453,N_2535,N_2100);
and U3454 (N_3454,N_2712,N_2415);
nand U3455 (N_3455,N_2279,N_2524);
or U3456 (N_3456,N_2083,N_2868);
nor U3457 (N_3457,N_2470,N_2659);
xor U3458 (N_3458,N_2123,N_2285);
or U3459 (N_3459,N_2596,N_2171);
nor U3460 (N_3460,N_2360,N_2945);
or U3461 (N_3461,N_2859,N_2839);
xnor U3462 (N_3462,N_2858,N_2574);
and U3463 (N_3463,N_2993,N_2666);
nand U3464 (N_3464,N_2381,N_2709);
and U3465 (N_3465,N_2934,N_2684);
xor U3466 (N_3466,N_2561,N_2104);
nor U3467 (N_3467,N_2721,N_2167);
xor U3468 (N_3468,N_2893,N_2565);
or U3469 (N_3469,N_2064,N_2834);
or U3470 (N_3470,N_2024,N_2030);
nand U3471 (N_3471,N_2878,N_2091);
and U3472 (N_3472,N_2601,N_2733);
nor U3473 (N_3473,N_2862,N_2638);
nor U3474 (N_3474,N_2713,N_2769);
and U3475 (N_3475,N_2864,N_2012);
xor U3476 (N_3476,N_2797,N_2244);
nand U3477 (N_3477,N_2830,N_2526);
or U3478 (N_3478,N_2293,N_2902);
nor U3479 (N_3479,N_2146,N_2282);
nor U3480 (N_3480,N_2089,N_2262);
or U3481 (N_3481,N_2139,N_2418);
or U3482 (N_3482,N_2677,N_2636);
xor U3483 (N_3483,N_2814,N_2501);
xor U3484 (N_3484,N_2829,N_2539);
nor U3485 (N_3485,N_2939,N_2124);
nor U3486 (N_3486,N_2486,N_2783);
xor U3487 (N_3487,N_2977,N_2161);
nor U3488 (N_3488,N_2340,N_2775);
nand U3489 (N_3489,N_2253,N_2897);
xor U3490 (N_3490,N_2604,N_2256);
and U3491 (N_3491,N_2519,N_2103);
xnor U3492 (N_3492,N_2484,N_2914);
xnor U3493 (N_3493,N_2771,N_2533);
xor U3494 (N_3494,N_2952,N_2670);
nor U3495 (N_3495,N_2086,N_2150);
and U3496 (N_3496,N_2613,N_2050);
nand U3497 (N_3497,N_2767,N_2773);
nand U3498 (N_3498,N_2177,N_2204);
nor U3499 (N_3499,N_2674,N_2250);
nor U3500 (N_3500,N_2544,N_2208);
nor U3501 (N_3501,N_2908,N_2222);
or U3502 (N_3502,N_2435,N_2693);
xnor U3503 (N_3503,N_2378,N_2528);
and U3504 (N_3504,N_2962,N_2194);
or U3505 (N_3505,N_2546,N_2131);
and U3506 (N_3506,N_2313,N_2881);
nand U3507 (N_3507,N_2501,N_2432);
or U3508 (N_3508,N_2329,N_2787);
xnor U3509 (N_3509,N_2610,N_2423);
and U3510 (N_3510,N_2965,N_2126);
or U3511 (N_3511,N_2142,N_2303);
and U3512 (N_3512,N_2624,N_2742);
nand U3513 (N_3513,N_2804,N_2553);
and U3514 (N_3514,N_2522,N_2026);
or U3515 (N_3515,N_2477,N_2257);
and U3516 (N_3516,N_2049,N_2445);
nor U3517 (N_3517,N_2906,N_2390);
and U3518 (N_3518,N_2635,N_2800);
nand U3519 (N_3519,N_2464,N_2665);
and U3520 (N_3520,N_2545,N_2823);
or U3521 (N_3521,N_2686,N_2622);
and U3522 (N_3522,N_2434,N_2031);
xnor U3523 (N_3523,N_2283,N_2525);
xor U3524 (N_3524,N_2262,N_2766);
nand U3525 (N_3525,N_2810,N_2501);
or U3526 (N_3526,N_2566,N_2631);
or U3527 (N_3527,N_2186,N_2613);
nand U3528 (N_3528,N_2303,N_2354);
and U3529 (N_3529,N_2165,N_2420);
or U3530 (N_3530,N_2180,N_2021);
and U3531 (N_3531,N_2480,N_2419);
nand U3532 (N_3532,N_2820,N_2853);
nand U3533 (N_3533,N_2931,N_2451);
xor U3534 (N_3534,N_2794,N_2126);
and U3535 (N_3535,N_2085,N_2460);
and U3536 (N_3536,N_2196,N_2990);
or U3537 (N_3537,N_2842,N_2934);
xnor U3538 (N_3538,N_2856,N_2070);
nor U3539 (N_3539,N_2882,N_2207);
nand U3540 (N_3540,N_2784,N_2422);
and U3541 (N_3541,N_2010,N_2370);
or U3542 (N_3542,N_2907,N_2297);
nand U3543 (N_3543,N_2961,N_2502);
or U3544 (N_3544,N_2775,N_2189);
and U3545 (N_3545,N_2278,N_2848);
or U3546 (N_3546,N_2105,N_2777);
xnor U3547 (N_3547,N_2569,N_2754);
nand U3548 (N_3548,N_2896,N_2212);
nand U3549 (N_3549,N_2827,N_2700);
nor U3550 (N_3550,N_2619,N_2758);
nor U3551 (N_3551,N_2596,N_2527);
and U3552 (N_3552,N_2851,N_2248);
and U3553 (N_3553,N_2997,N_2722);
nor U3554 (N_3554,N_2639,N_2965);
xnor U3555 (N_3555,N_2916,N_2017);
or U3556 (N_3556,N_2247,N_2027);
and U3557 (N_3557,N_2564,N_2305);
nor U3558 (N_3558,N_2193,N_2412);
nand U3559 (N_3559,N_2200,N_2092);
nor U3560 (N_3560,N_2621,N_2880);
nand U3561 (N_3561,N_2639,N_2177);
xor U3562 (N_3562,N_2483,N_2442);
nor U3563 (N_3563,N_2304,N_2504);
and U3564 (N_3564,N_2369,N_2919);
and U3565 (N_3565,N_2667,N_2236);
nand U3566 (N_3566,N_2539,N_2920);
and U3567 (N_3567,N_2927,N_2262);
nand U3568 (N_3568,N_2045,N_2041);
or U3569 (N_3569,N_2377,N_2838);
nand U3570 (N_3570,N_2859,N_2379);
and U3571 (N_3571,N_2418,N_2970);
nor U3572 (N_3572,N_2611,N_2347);
nor U3573 (N_3573,N_2069,N_2295);
or U3574 (N_3574,N_2597,N_2841);
or U3575 (N_3575,N_2688,N_2669);
nand U3576 (N_3576,N_2345,N_2142);
nand U3577 (N_3577,N_2441,N_2139);
or U3578 (N_3578,N_2288,N_2120);
or U3579 (N_3579,N_2923,N_2058);
nor U3580 (N_3580,N_2322,N_2407);
xnor U3581 (N_3581,N_2547,N_2245);
and U3582 (N_3582,N_2782,N_2840);
nor U3583 (N_3583,N_2309,N_2435);
xor U3584 (N_3584,N_2865,N_2406);
nor U3585 (N_3585,N_2476,N_2486);
and U3586 (N_3586,N_2854,N_2161);
or U3587 (N_3587,N_2159,N_2855);
and U3588 (N_3588,N_2791,N_2636);
or U3589 (N_3589,N_2077,N_2512);
or U3590 (N_3590,N_2744,N_2524);
nand U3591 (N_3591,N_2722,N_2880);
nor U3592 (N_3592,N_2514,N_2891);
xor U3593 (N_3593,N_2898,N_2323);
or U3594 (N_3594,N_2752,N_2083);
nand U3595 (N_3595,N_2873,N_2131);
and U3596 (N_3596,N_2390,N_2879);
xor U3597 (N_3597,N_2178,N_2927);
nand U3598 (N_3598,N_2170,N_2854);
nor U3599 (N_3599,N_2210,N_2694);
nor U3600 (N_3600,N_2759,N_2953);
or U3601 (N_3601,N_2475,N_2868);
nand U3602 (N_3602,N_2570,N_2110);
and U3603 (N_3603,N_2073,N_2607);
xor U3604 (N_3604,N_2836,N_2027);
xnor U3605 (N_3605,N_2175,N_2478);
nor U3606 (N_3606,N_2521,N_2981);
and U3607 (N_3607,N_2947,N_2988);
and U3608 (N_3608,N_2358,N_2463);
nor U3609 (N_3609,N_2308,N_2980);
or U3610 (N_3610,N_2467,N_2941);
and U3611 (N_3611,N_2915,N_2061);
or U3612 (N_3612,N_2164,N_2148);
nor U3613 (N_3613,N_2535,N_2798);
and U3614 (N_3614,N_2936,N_2652);
nand U3615 (N_3615,N_2076,N_2768);
nor U3616 (N_3616,N_2102,N_2447);
xnor U3617 (N_3617,N_2466,N_2001);
nand U3618 (N_3618,N_2710,N_2852);
or U3619 (N_3619,N_2274,N_2569);
nand U3620 (N_3620,N_2223,N_2660);
and U3621 (N_3621,N_2653,N_2801);
and U3622 (N_3622,N_2654,N_2217);
xnor U3623 (N_3623,N_2506,N_2796);
nand U3624 (N_3624,N_2707,N_2534);
xor U3625 (N_3625,N_2023,N_2642);
nand U3626 (N_3626,N_2773,N_2068);
and U3627 (N_3627,N_2527,N_2757);
and U3628 (N_3628,N_2510,N_2719);
xor U3629 (N_3629,N_2755,N_2789);
or U3630 (N_3630,N_2507,N_2250);
xor U3631 (N_3631,N_2373,N_2464);
xor U3632 (N_3632,N_2200,N_2054);
or U3633 (N_3633,N_2673,N_2987);
xnor U3634 (N_3634,N_2429,N_2093);
and U3635 (N_3635,N_2205,N_2553);
or U3636 (N_3636,N_2169,N_2897);
nand U3637 (N_3637,N_2488,N_2035);
and U3638 (N_3638,N_2200,N_2325);
nor U3639 (N_3639,N_2548,N_2830);
xor U3640 (N_3640,N_2864,N_2790);
or U3641 (N_3641,N_2284,N_2722);
nand U3642 (N_3642,N_2435,N_2874);
or U3643 (N_3643,N_2823,N_2419);
or U3644 (N_3644,N_2040,N_2409);
or U3645 (N_3645,N_2473,N_2188);
or U3646 (N_3646,N_2364,N_2281);
nor U3647 (N_3647,N_2255,N_2520);
xnor U3648 (N_3648,N_2274,N_2060);
xnor U3649 (N_3649,N_2673,N_2403);
and U3650 (N_3650,N_2183,N_2661);
nor U3651 (N_3651,N_2886,N_2850);
and U3652 (N_3652,N_2779,N_2593);
and U3653 (N_3653,N_2363,N_2820);
xor U3654 (N_3654,N_2695,N_2225);
nor U3655 (N_3655,N_2335,N_2935);
nand U3656 (N_3656,N_2272,N_2723);
nor U3657 (N_3657,N_2408,N_2541);
or U3658 (N_3658,N_2134,N_2703);
nor U3659 (N_3659,N_2308,N_2266);
nand U3660 (N_3660,N_2530,N_2458);
nor U3661 (N_3661,N_2150,N_2826);
and U3662 (N_3662,N_2686,N_2373);
nand U3663 (N_3663,N_2741,N_2322);
nand U3664 (N_3664,N_2217,N_2805);
nor U3665 (N_3665,N_2586,N_2076);
or U3666 (N_3666,N_2235,N_2677);
or U3667 (N_3667,N_2526,N_2127);
and U3668 (N_3668,N_2637,N_2266);
or U3669 (N_3669,N_2280,N_2427);
xor U3670 (N_3670,N_2287,N_2691);
or U3671 (N_3671,N_2434,N_2335);
or U3672 (N_3672,N_2246,N_2959);
or U3673 (N_3673,N_2263,N_2505);
xnor U3674 (N_3674,N_2456,N_2411);
xor U3675 (N_3675,N_2726,N_2201);
and U3676 (N_3676,N_2330,N_2904);
or U3677 (N_3677,N_2915,N_2031);
nand U3678 (N_3678,N_2811,N_2172);
xor U3679 (N_3679,N_2999,N_2378);
nand U3680 (N_3680,N_2271,N_2987);
and U3681 (N_3681,N_2898,N_2000);
nand U3682 (N_3682,N_2226,N_2828);
and U3683 (N_3683,N_2996,N_2014);
nand U3684 (N_3684,N_2887,N_2097);
xnor U3685 (N_3685,N_2005,N_2397);
or U3686 (N_3686,N_2421,N_2650);
nand U3687 (N_3687,N_2978,N_2198);
xor U3688 (N_3688,N_2000,N_2606);
nor U3689 (N_3689,N_2210,N_2065);
and U3690 (N_3690,N_2331,N_2799);
and U3691 (N_3691,N_2800,N_2910);
nand U3692 (N_3692,N_2564,N_2574);
xor U3693 (N_3693,N_2596,N_2089);
or U3694 (N_3694,N_2662,N_2192);
nand U3695 (N_3695,N_2967,N_2474);
xor U3696 (N_3696,N_2595,N_2517);
or U3697 (N_3697,N_2415,N_2052);
or U3698 (N_3698,N_2098,N_2636);
or U3699 (N_3699,N_2488,N_2399);
nand U3700 (N_3700,N_2719,N_2906);
nand U3701 (N_3701,N_2149,N_2053);
nor U3702 (N_3702,N_2307,N_2333);
and U3703 (N_3703,N_2876,N_2556);
or U3704 (N_3704,N_2105,N_2595);
nand U3705 (N_3705,N_2215,N_2947);
nand U3706 (N_3706,N_2146,N_2070);
nor U3707 (N_3707,N_2198,N_2777);
and U3708 (N_3708,N_2495,N_2455);
xor U3709 (N_3709,N_2654,N_2102);
nand U3710 (N_3710,N_2536,N_2465);
and U3711 (N_3711,N_2555,N_2599);
nor U3712 (N_3712,N_2087,N_2672);
and U3713 (N_3713,N_2668,N_2852);
or U3714 (N_3714,N_2328,N_2017);
nand U3715 (N_3715,N_2294,N_2537);
and U3716 (N_3716,N_2473,N_2223);
nor U3717 (N_3717,N_2714,N_2255);
nor U3718 (N_3718,N_2090,N_2009);
or U3719 (N_3719,N_2948,N_2736);
xor U3720 (N_3720,N_2558,N_2886);
nor U3721 (N_3721,N_2054,N_2036);
or U3722 (N_3722,N_2659,N_2952);
xnor U3723 (N_3723,N_2627,N_2138);
or U3724 (N_3724,N_2087,N_2344);
and U3725 (N_3725,N_2784,N_2932);
xor U3726 (N_3726,N_2510,N_2272);
and U3727 (N_3727,N_2894,N_2686);
or U3728 (N_3728,N_2509,N_2693);
or U3729 (N_3729,N_2158,N_2411);
xor U3730 (N_3730,N_2407,N_2247);
nor U3731 (N_3731,N_2942,N_2254);
or U3732 (N_3732,N_2482,N_2234);
or U3733 (N_3733,N_2748,N_2608);
or U3734 (N_3734,N_2292,N_2153);
or U3735 (N_3735,N_2325,N_2288);
and U3736 (N_3736,N_2471,N_2205);
nor U3737 (N_3737,N_2441,N_2572);
xnor U3738 (N_3738,N_2486,N_2437);
xnor U3739 (N_3739,N_2443,N_2607);
nand U3740 (N_3740,N_2313,N_2944);
nor U3741 (N_3741,N_2228,N_2402);
nor U3742 (N_3742,N_2960,N_2108);
and U3743 (N_3743,N_2784,N_2554);
or U3744 (N_3744,N_2860,N_2212);
nor U3745 (N_3745,N_2392,N_2341);
or U3746 (N_3746,N_2307,N_2790);
nand U3747 (N_3747,N_2969,N_2428);
nor U3748 (N_3748,N_2072,N_2471);
xor U3749 (N_3749,N_2796,N_2784);
and U3750 (N_3750,N_2955,N_2455);
or U3751 (N_3751,N_2273,N_2966);
nand U3752 (N_3752,N_2195,N_2125);
nand U3753 (N_3753,N_2358,N_2579);
nand U3754 (N_3754,N_2552,N_2571);
xnor U3755 (N_3755,N_2576,N_2565);
nand U3756 (N_3756,N_2039,N_2360);
nand U3757 (N_3757,N_2602,N_2479);
xor U3758 (N_3758,N_2745,N_2736);
nor U3759 (N_3759,N_2627,N_2719);
nor U3760 (N_3760,N_2095,N_2572);
or U3761 (N_3761,N_2346,N_2337);
xnor U3762 (N_3762,N_2721,N_2448);
and U3763 (N_3763,N_2883,N_2057);
or U3764 (N_3764,N_2922,N_2908);
or U3765 (N_3765,N_2002,N_2456);
nand U3766 (N_3766,N_2900,N_2243);
or U3767 (N_3767,N_2233,N_2610);
or U3768 (N_3768,N_2352,N_2758);
or U3769 (N_3769,N_2864,N_2731);
nand U3770 (N_3770,N_2314,N_2260);
xnor U3771 (N_3771,N_2711,N_2807);
and U3772 (N_3772,N_2118,N_2362);
and U3773 (N_3773,N_2164,N_2268);
nor U3774 (N_3774,N_2795,N_2761);
or U3775 (N_3775,N_2968,N_2326);
nor U3776 (N_3776,N_2357,N_2482);
nor U3777 (N_3777,N_2462,N_2676);
nand U3778 (N_3778,N_2377,N_2950);
xnor U3779 (N_3779,N_2813,N_2907);
xor U3780 (N_3780,N_2732,N_2412);
or U3781 (N_3781,N_2506,N_2276);
or U3782 (N_3782,N_2195,N_2039);
nand U3783 (N_3783,N_2522,N_2878);
xnor U3784 (N_3784,N_2606,N_2526);
nand U3785 (N_3785,N_2964,N_2024);
and U3786 (N_3786,N_2291,N_2970);
or U3787 (N_3787,N_2160,N_2791);
nor U3788 (N_3788,N_2546,N_2791);
and U3789 (N_3789,N_2065,N_2175);
and U3790 (N_3790,N_2054,N_2766);
nor U3791 (N_3791,N_2331,N_2419);
nor U3792 (N_3792,N_2617,N_2038);
and U3793 (N_3793,N_2495,N_2489);
or U3794 (N_3794,N_2346,N_2243);
xnor U3795 (N_3795,N_2211,N_2257);
or U3796 (N_3796,N_2120,N_2583);
and U3797 (N_3797,N_2315,N_2011);
and U3798 (N_3798,N_2292,N_2964);
and U3799 (N_3799,N_2218,N_2959);
and U3800 (N_3800,N_2025,N_2676);
or U3801 (N_3801,N_2432,N_2574);
xnor U3802 (N_3802,N_2509,N_2206);
nand U3803 (N_3803,N_2038,N_2053);
nand U3804 (N_3804,N_2746,N_2293);
xnor U3805 (N_3805,N_2816,N_2805);
nand U3806 (N_3806,N_2221,N_2393);
nand U3807 (N_3807,N_2433,N_2750);
nor U3808 (N_3808,N_2147,N_2887);
nand U3809 (N_3809,N_2653,N_2463);
nor U3810 (N_3810,N_2894,N_2549);
xnor U3811 (N_3811,N_2408,N_2178);
xnor U3812 (N_3812,N_2304,N_2808);
nor U3813 (N_3813,N_2367,N_2015);
nor U3814 (N_3814,N_2290,N_2621);
nor U3815 (N_3815,N_2899,N_2539);
nand U3816 (N_3816,N_2522,N_2482);
nor U3817 (N_3817,N_2901,N_2142);
and U3818 (N_3818,N_2533,N_2198);
xor U3819 (N_3819,N_2924,N_2112);
xnor U3820 (N_3820,N_2948,N_2112);
or U3821 (N_3821,N_2133,N_2369);
nor U3822 (N_3822,N_2452,N_2762);
or U3823 (N_3823,N_2650,N_2430);
xor U3824 (N_3824,N_2506,N_2727);
nand U3825 (N_3825,N_2209,N_2868);
xor U3826 (N_3826,N_2168,N_2161);
nand U3827 (N_3827,N_2685,N_2809);
xnor U3828 (N_3828,N_2432,N_2518);
nor U3829 (N_3829,N_2005,N_2036);
xnor U3830 (N_3830,N_2393,N_2614);
or U3831 (N_3831,N_2863,N_2374);
and U3832 (N_3832,N_2332,N_2907);
or U3833 (N_3833,N_2296,N_2440);
and U3834 (N_3834,N_2209,N_2004);
or U3835 (N_3835,N_2631,N_2061);
or U3836 (N_3836,N_2592,N_2418);
nor U3837 (N_3837,N_2035,N_2168);
xnor U3838 (N_3838,N_2848,N_2841);
xnor U3839 (N_3839,N_2530,N_2037);
xnor U3840 (N_3840,N_2642,N_2077);
and U3841 (N_3841,N_2961,N_2036);
nand U3842 (N_3842,N_2965,N_2005);
xor U3843 (N_3843,N_2028,N_2231);
xnor U3844 (N_3844,N_2963,N_2996);
xnor U3845 (N_3845,N_2269,N_2756);
xor U3846 (N_3846,N_2637,N_2563);
or U3847 (N_3847,N_2633,N_2684);
nand U3848 (N_3848,N_2573,N_2821);
nand U3849 (N_3849,N_2973,N_2791);
and U3850 (N_3850,N_2774,N_2678);
xnor U3851 (N_3851,N_2940,N_2647);
or U3852 (N_3852,N_2313,N_2108);
and U3853 (N_3853,N_2601,N_2653);
and U3854 (N_3854,N_2910,N_2714);
nor U3855 (N_3855,N_2403,N_2964);
or U3856 (N_3856,N_2375,N_2874);
and U3857 (N_3857,N_2458,N_2504);
xor U3858 (N_3858,N_2424,N_2654);
nand U3859 (N_3859,N_2889,N_2066);
and U3860 (N_3860,N_2575,N_2203);
nor U3861 (N_3861,N_2912,N_2695);
xnor U3862 (N_3862,N_2096,N_2175);
nor U3863 (N_3863,N_2382,N_2703);
and U3864 (N_3864,N_2617,N_2760);
or U3865 (N_3865,N_2863,N_2135);
xnor U3866 (N_3866,N_2097,N_2525);
xor U3867 (N_3867,N_2201,N_2802);
nand U3868 (N_3868,N_2117,N_2304);
xnor U3869 (N_3869,N_2100,N_2841);
and U3870 (N_3870,N_2287,N_2166);
nor U3871 (N_3871,N_2384,N_2912);
xor U3872 (N_3872,N_2610,N_2405);
xor U3873 (N_3873,N_2434,N_2574);
or U3874 (N_3874,N_2015,N_2329);
and U3875 (N_3875,N_2042,N_2401);
nand U3876 (N_3876,N_2426,N_2453);
and U3877 (N_3877,N_2264,N_2248);
xnor U3878 (N_3878,N_2842,N_2470);
and U3879 (N_3879,N_2801,N_2585);
xor U3880 (N_3880,N_2078,N_2928);
xnor U3881 (N_3881,N_2023,N_2785);
nand U3882 (N_3882,N_2638,N_2216);
nor U3883 (N_3883,N_2436,N_2986);
nor U3884 (N_3884,N_2761,N_2302);
or U3885 (N_3885,N_2684,N_2902);
nand U3886 (N_3886,N_2813,N_2123);
or U3887 (N_3887,N_2070,N_2057);
and U3888 (N_3888,N_2214,N_2355);
xnor U3889 (N_3889,N_2572,N_2940);
xnor U3890 (N_3890,N_2149,N_2412);
xor U3891 (N_3891,N_2963,N_2230);
nor U3892 (N_3892,N_2314,N_2146);
nand U3893 (N_3893,N_2319,N_2192);
and U3894 (N_3894,N_2078,N_2456);
and U3895 (N_3895,N_2051,N_2396);
and U3896 (N_3896,N_2170,N_2836);
and U3897 (N_3897,N_2865,N_2325);
or U3898 (N_3898,N_2554,N_2466);
xor U3899 (N_3899,N_2574,N_2925);
xor U3900 (N_3900,N_2453,N_2191);
nor U3901 (N_3901,N_2664,N_2960);
nor U3902 (N_3902,N_2410,N_2671);
xnor U3903 (N_3903,N_2354,N_2938);
nor U3904 (N_3904,N_2685,N_2051);
or U3905 (N_3905,N_2098,N_2456);
xor U3906 (N_3906,N_2638,N_2720);
and U3907 (N_3907,N_2885,N_2243);
xor U3908 (N_3908,N_2560,N_2653);
or U3909 (N_3909,N_2238,N_2945);
nor U3910 (N_3910,N_2231,N_2821);
nand U3911 (N_3911,N_2080,N_2165);
nand U3912 (N_3912,N_2302,N_2835);
and U3913 (N_3913,N_2963,N_2420);
or U3914 (N_3914,N_2983,N_2079);
and U3915 (N_3915,N_2259,N_2814);
nor U3916 (N_3916,N_2805,N_2090);
nand U3917 (N_3917,N_2283,N_2841);
and U3918 (N_3918,N_2946,N_2079);
nand U3919 (N_3919,N_2719,N_2391);
xnor U3920 (N_3920,N_2279,N_2166);
and U3921 (N_3921,N_2718,N_2389);
xnor U3922 (N_3922,N_2464,N_2035);
xor U3923 (N_3923,N_2629,N_2305);
nor U3924 (N_3924,N_2934,N_2309);
nor U3925 (N_3925,N_2814,N_2914);
nand U3926 (N_3926,N_2656,N_2928);
and U3927 (N_3927,N_2059,N_2036);
nand U3928 (N_3928,N_2365,N_2427);
nor U3929 (N_3929,N_2799,N_2686);
or U3930 (N_3930,N_2749,N_2836);
xor U3931 (N_3931,N_2073,N_2542);
or U3932 (N_3932,N_2585,N_2981);
nor U3933 (N_3933,N_2132,N_2782);
nand U3934 (N_3934,N_2034,N_2181);
xnor U3935 (N_3935,N_2192,N_2539);
and U3936 (N_3936,N_2741,N_2791);
nand U3937 (N_3937,N_2033,N_2634);
and U3938 (N_3938,N_2056,N_2017);
xnor U3939 (N_3939,N_2255,N_2169);
and U3940 (N_3940,N_2534,N_2246);
nor U3941 (N_3941,N_2645,N_2213);
and U3942 (N_3942,N_2495,N_2639);
and U3943 (N_3943,N_2604,N_2170);
and U3944 (N_3944,N_2592,N_2890);
and U3945 (N_3945,N_2702,N_2900);
nand U3946 (N_3946,N_2751,N_2316);
and U3947 (N_3947,N_2104,N_2914);
and U3948 (N_3948,N_2711,N_2245);
nor U3949 (N_3949,N_2375,N_2425);
nand U3950 (N_3950,N_2271,N_2675);
nand U3951 (N_3951,N_2005,N_2242);
or U3952 (N_3952,N_2197,N_2394);
xnor U3953 (N_3953,N_2115,N_2898);
and U3954 (N_3954,N_2634,N_2570);
and U3955 (N_3955,N_2860,N_2942);
xor U3956 (N_3956,N_2111,N_2265);
nor U3957 (N_3957,N_2863,N_2291);
xnor U3958 (N_3958,N_2548,N_2861);
xor U3959 (N_3959,N_2128,N_2225);
and U3960 (N_3960,N_2067,N_2330);
nor U3961 (N_3961,N_2045,N_2154);
nand U3962 (N_3962,N_2918,N_2722);
and U3963 (N_3963,N_2567,N_2139);
and U3964 (N_3964,N_2220,N_2317);
or U3965 (N_3965,N_2766,N_2398);
nor U3966 (N_3966,N_2184,N_2864);
nor U3967 (N_3967,N_2817,N_2206);
and U3968 (N_3968,N_2035,N_2482);
xnor U3969 (N_3969,N_2313,N_2544);
nor U3970 (N_3970,N_2399,N_2085);
and U3971 (N_3971,N_2460,N_2105);
xor U3972 (N_3972,N_2527,N_2670);
nor U3973 (N_3973,N_2586,N_2098);
nor U3974 (N_3974,N_2925,N_2671);
or U3975 (N_3975,N_2968,N_2106);
or U3976 (N_3976,N_2326,N_2746);
nor U3977 (N_3977,N_2141,N_2214);
nand U3978 (N_3978,N_2809,N_2923);
nor U3979 (N_3979,N_2703,N_2731);
nor U3980 (N_3980,N_2701,N_2012);
nand U3981 (N_3981,N_2439,N_2069);
nor U3982 (N_3982,N_2930,N_2242);
xnor U3983 (N_3983,N_2300,N_2482);
and U3984 (N_3984,N_2679,N_2714);
and U3985 (N_3985,N_2800,N_2350);
or U3986 (N_3986,N_2336,N_2393);
nand U3987 (N_3987,N_2868,N_2148);
or U3988 (N_3988,N_2538,N_2294);
nand U3989 (N_3989,N_2521,N_2192);
nor U3990 (N_3990,N_2770,N_2890);
xnor U3991 (N_3991,N_2352,N_2026);
xnor U3992 (N_3992,N_2743,N_2467);
nor U3993 (N_3993,N_2715,N_2419);
and U3994 (N_3994,N_2975,N_2592);
nand U3995 (N_3995,N_2218,N_2021);
and U3996 (N_3996,N_2010,N_2792);
xor U3997 (N_3997,N_2077,N_2573);
and U3998 (N_3998,N_2319,N_2699);
nor U3999 (N_3999,N_2542,N_2547);
or U4000 (N_4000,N_3789,N_3573);
xnor U4001 (N_4001,N_3864,N_3575);
xor U4002 (N_4002,N_3736,N_3879);
or U4003 (N_4003,N_3241,N_3987);
xnor U4004 (N_4004,N_3989,N_3658);
nand U4005 (N_4005,N_3451,N_3534);
and U4006 (N_4006,N_3279,N_3657);
and U4007 (N_4007,N_3321,N_3886);
or U4008 (N_4008,N_3353,N_3191);
nand U4009 (N_4009,N_3696,N_3154);
nand U4010 (N_4010,N_3731,N_3602);
xor U4011 (N_4011,N_3294,N_3666);
and U4012 (N_4012,N_3040,N_3904);
or U4013 (N_4013,N_3887,N_3601);
nand U4014 (N_4014,N_3084,N_3101);
nor U4015 (N_4015,N_3242,N_3867);
or U4016 (N_4016,N_3512,N_3803);
xnor U4017 (N_4017,N_3131,N_3942);
nand U4018 (N_4018,N_3029,N_3516);
or U4019 (N_4019,N_3151,N_3769);
and U4020 (N_4020,N_3930,N_3238);
xnor U4021 (N_4021,N_3617,N_3269);
nand U4022 (N_4022,N_3903,N_3665);
nand U4023 (N_4023,N_3061,N_3290);
nor U4024 (N_4024,N_3271,N_3206);
and U4025 (N_4025,N_3068,N_3328);
xor U4026 (N_4026,N_3137,N_3664);
xnor U4027 (N_4027,N_3459,N_3087);
nor U4028 (N_4028,N_3521,N_3950);
or U4029 (N_4029,N_3817,N_3729);
and U4030 (N_4030,N_3974,N_3161);
or U4031 (N_4031,N_3750,N_3311);
or U4032 (N_4032,N_3509,N_3334);
xnor U4033 (N_4033,N_3198,N_3035);
nor U4034 (N_4034,N_3868,N_3452);
nand U4035 (N_4035,N_3285,N_3225);
and U4036 (N_4036,N_3663,N_3562);
or U4037 (N_4037,N_3286,N_3089);
and U4038 (N_4038,N_3860,N_3259);
or U4039 (N_4039,N_3100,N_3614);
nor U4040 (N_4040,N_3515,N_3183);
nor U4041 (N_4041,N_3379,N_3944);
or U4042 (N_4042,N_3160,N_3110);
xnor U4043 (N_4043,N_3656,N_3484);
nand U4044 (N_4044,N_3976,N_3244);
nand U4045 (N_4045,N_3468,N_3966);
nand U4046 (N_4046,N_3184,N_3748);
and U4047 (N_4047,N_3999,N_3098);
nor U4048 (N_4048,N_3308,N_3755);
nand U4049 (N_4049,N_3994,N_3367);
and U4050 (N_4050,N_3991,N_3365);
xnor U4051 (N_4051,N_3243,N_3037);
or U4052 (N_4052,N_3827,N_3275);
and U4053 (N_4053,N_3996,N_3090);
nor U4054 (N_4054,N_3929,N_3466);
and U4055 (N_4055,N_3413,N_3165);
nand U4056 (N_4056,N_3292,N_3371);
nor U4057 (N_4057,N_3687,N_3185);
nand U4058 (N_4058,N_3517,N_3266);
nor U4059 (N_4059,N_3073,N_3020);
nor U4060 (N_4060,N_3473,N_3431);
nor U4061 (N_4061,N_3938,N_3965);
and U4062 (N_4062,N_3680,N_3103);
xor U4063 (N_4063,N_3044,N_3799);
nand U4064 (N_4064,N_3193,N_3257);
nor U4065 (N_4065,N_3390,N_3757);
and U4066 (N_4066,N_3215,N_3033);
nand U4067 (N_4067,N_3330,N_3897);
nand U4068 (N_4068,N_3577,N_3447);
nand U4069 (N_4069,N_3756,N_3690);
or U4070 (N_4070,N_3639,N_3995);
and U4071 (N_4071,N_3941,N_3706);
nor U4072 (N_4072,N_3122,N_3915);
or U4073 (N_4073,N_3806,N_3818);
and U4074 (N_4074,N_3310,N_3300);
xnor U4075 (N_4075,N_3071,N_3004);
nand U4076 (N_4076,N_3946,N_3104);
nor U4077 (N_4077,N_3545,N_3564);
or U4078 (N_4078,N_3091,N_3066);
nor U4079 (N_4079,N_3819,N_3256);
xor U4080 (N_4080,N_3219,N_3265);
nand U4081 (N_4081,N_3895,N_3661);
xnor U4082 (N_4082,N_3503,N_3600);
nand U4083 (N_4083,N_3496,N_3546);
or U4084 (N_4084,N_3309,N_3357);
xor U4085 (N_4085,N_3507,N_3912);
and U4086 (N_4086,N_3060,N_3724);
xnor U4087 (N_4087,N_3423,N_3003);
nand U4088 (N_4088,N_3253,N_3366);
xor U4089 (N_4089,N_3030,N_3906);
or U4090 (N_4090,N_3607,N_3597);
and U4091 (N_4091,N_3524,N_3914);
xor U4092 (N_4092,N_3199,N_3155);
nand U4093 (N_4093,N_3361,N_3947);
and U4094 (N_4094,N_3857,N_3398);
nand U4095 (N_4095,N_3832,N_3646);
or U4096 (N_4096,N_3172,N_3691);
and U4097 (N_4097,N_3634,N_3475);
nor U4098 (N_4098,N_3758,N_3847);
and U4099 (N_4099,N_3317,N_3316);
and U4100 (N_4100,N_3149,N_3717);
nor U4101 (N_4101,N_3862,N_3686);
or U4102 (N_4102,N_3234,N_3877);
xor U4103 (N_4103,N_3523,N_3069);
nand U4104 (N_4104,N_3108,N_3982);
xnor U4105 (N_4105,N_3025,N_3583);
or U4106 (N_4106,N_3802,N_3402);
nand U4107 (N_4107,N_3192,N_3032);
xnor U4108 (N_4108,N_3822,N_3718);
nor U4109 (N_4109,N_3435,N_3625);
nand U4110 (N_4110,N_3767,N_3450);
xnor U4111 (N_4111,N_3418,N_3981);
and U4112 (N_4112,N_3063,N_3815);
or U4113 (N_4113,N_3039,N_3045);
xnor U4114 (N_4114,N_3074,N_3107);
or U4115 (N_4115,N_3386,N_3943);
nand U4116 (N_4116,N_3843,N_3358);
nor U4117 (N_4117,N_3760,N_3627);
and U4118 (N_4118,N_3732,N_3624);
and U4119 (N_4119,N_3099,N_3223);
or U4120 (N_4120,N_3688,N_3824);
and U4121 (N_4121,N_3430,N_3407);
and U4122 (N_4122,N_3791,N_3931);
nand U4123 (N_4123,N_3636,N_3876);
and U4124 (N_4124,N_3884,N_3700);
nor U4125 (N_4125,N_3499,N_3383);
nand U4126 (N_4126,N_3412,N_3428);
nor U4127 (N_4127,N_3844,N_3477);
and U4128 (N_4128,N_3923,N_3293);
nor U4129 (N_4129,N_3740,N_3894);
or U4130 (N_4130,N_3980,N_3917);
nand U4131 (N_4131,N_3124,N_3227);
nor U4132 (N_4132,N_3526,N_3725);
nor U4133 (N_4133,N_3962,N_3299);
nand U4134 (N_4134,N_3993,N_3853);
xnor U4135 (N_4135,N_3111,N_3608);
xor U4136 (N_4136,N_3631,N_3341);
nand U4137 (N_4137,N_3217,N_3434);
nand U4138 (N_4138,N_3081,N_3404);
or U4139 (N_4139,N_3618,N_3382);
or U4140 (N_4140,N_3850,N_3247);
and U4141 (N_4141,N_3008,N_3319);
or U4142 (N_4142,N_3659,N_3220);
nand U4143 (N_4143,N_3010,N_3694);
nor U4144 (N_4144,N_3922,N_3555);
nor U4145 (N_4145,N_3539,N_3650);
xnor U4146 (N_4146,N_3851,N_3798);
or U4147 (N_4147,N_3814,N_3504);
or U4148 (N_4148,N_3653,N_3830);
or U4149 (N_4149,N_3992,N_3533);
or U4150 (N_4150,N_3394,N_3861);
and U4151 (N_4151,N_3716,N_3576);
nor U4152 (N_4152,N_3261,N_3056);
xnor U4153 (N_4153,N_3405,N_3115);
or U4154 (N_4154,N_3794,N_3538);
nor U4155 (N_4155,N_3296,N_3479);
xor U4156 (N_4156,N_3465,N_3239);
nand U4157 (N_4157,N_3076,N_3537);
nand U4158 (N_4158,N_3342,N_3644);
nand U4159 (N_4159,N_3859,N_3273);
nor U4160 (N_4160,N_3753,N_3858);
nor U4161 (N_4161,N_3399,N_3442);
or U4162 (N_4162,N_3977,N_3018);
nor U4163 (N_4163,N_3335,N_3188);
or U4164 (N_4164,N_3514,N_3871);
nand U4165 (N_4165,N_3594,N_3128);
and U4166 (N_4166,N_3331,N_3795);
and U4167 (N_4167,N_3359,N_3648);
and U4168 (N_4168,N_3591,N_3505);
or U4169 (N_4169,N_3351,N_3488);
nor U4170 (N_4170,N_3167,N_3547);
xnor U4171 (N_4171,N_3751,N_3826);
and U4172 (N_4172,N_3936,N_3939);
xor U4173 (N_4173,N_3143,N_3774);
or U4174 (N_4174,N_3449,N_3727);
xor U4175 (N_4175,N_3375,N_3743);
or U4176 (N_4176,N_3440,N_3554);
and U4177 (N_4177,N_3508,N_3142);
or U4178 (N_4178,N_3189,N_3157);
xor U4179 (N_4179,N_3834,N_3264);
and U4180 (N_4180,N_3780,N_3667);
nor U4181 (N_4181,N_3113,N_3381);
or U4182 (N_4182,N_3338,N_3204);
and U4183 (N_4183,N_3775,N_3377);
and U4184 (N_4184,N_3721,N_3118);
or U4185 (N_4185,N_3820,N_3675);
nor U4186 (N_4186,N_3967,N_3001);
nand U4187 (N_4187,N_3075,N_3628);
nand U4188 (N_4188,N_3454,N_3590);
xnor U4189 (N_4189,N_3248,N_3368);
nor U4190 (N_4190,N_3570,N_3920);
and U4191 (N_4191,N_3043,N_3426);
and U4192 (N_4192,N_3322,N_3722);
and U4193 (N_4193,N_3875,N_3749);
nand U4194 (N_4194,N_3222,N_3782);
and U4195 (N_4195,N_3121,N_3582);
and U4196 (N_4196,N_3747,N_3000);
xnor U4197 (N_4197,N_3948,N_3202);
nor U4198 (N_4198,N_3211,N_3878);
xor U4199 (N_4199,N_3811,N_3671);
xor U4200 (N_4200,N_3134,N_3494);
xor U4201 (N_4201,N_3699,N_3096);
or U4202 (N_4202,N_3986,N_3112);
xor U4203 (N_4203,N_3541,N_3138);
nand U4204 (N_4204,N_3051,N_3865);
xnor U4205 (N_4205,N_3622,N_3072);
nor U4206 (N_4206,N_3088,N_3543);
nor U4207 (N_4207,N_3120,N_3070);
nor U4208 (N_4208,N_3179,N_3606);
and U4209 (N_4209,N_3026,N_3848);
and U4210 (N_4210,N_3762,N_3422);
or U4211 (N_4211,N_3017,N_3506);
or U4212 (N_4212,N_3298,N_3781);
nand U4213 (N_4213,N_3733,N_3899);
nand U4214 (N_4214,N_3773,N_3563);
nor U4215 (N_4215,N_3136,N_3233);
and U4216 (N_4216,N_3809,N_3208);
nand U4217 (N_4217,N_3352,N_3194);
or U4218 (N_4218,N_3683,N_3693);
nand U4219 (N_4219,N_3280,N_3821);
and U4220 (N_4220,N_3277,N_3937);
nor U4221 (N_4221,N_3015,N_3713);
nor U4222 (N_4222,N_3905,N_3370);
xnor U4223 (N_4223,N_3985,N_3196);
xnor U4224 (N_4224,N_3307,N_3213);
nand U4225 (N_4225,N_3954,N_3093);
and U4226 (N_4226,N_3129,N_3633);
nand U4227 (N_4227,N_3882,N_3957);
nor U4228 (N_4228,N_3489,N_3162);
or U4229 (N_4229,N_3778,N_3953);
nand U4230 (N_4230,N_3552,N_3487);
nor U4231 (N_4231,N_3355,N_3140);
nor U4232 (N_4232,N_3707,N_3510);
or U4233 (N_4233,N_3356,N_3186);
nor U4234 (N_4234,N_3260,N_3079);
xnor U4235 (N_4235,N_3497,N_3949);
xnor U4236 (N_4236,N_3152,N_3741);
xnor U4237 (N_4237,N_3491,N_3175);
or U4238 (N_4238,N_3952,N_3840);
and U4239 (N_4239,N_3207,N_3393);
xnor U4240 (N_4240,N_3963,N_3800);
or U4241 (N_4241,N_3187,N_3349);
nand U4242 (N_4242,N_3893,N_3150);
nor U4243 (N_4243,N_3173,N_3770);
nand U4244 (N_4244,N_3086,N_3205);
nor U4245 (N_4245,N_3889,N_3908);
nor U4246 (N_4246,N_3461,N_3444);
nand U4247 (N_4247,N_3472,N_3574);
nor U4248 (N_4248,N_3182,N_3542);
and U4249 (N_4249,N_3346,N_3610);
xnor U4250 (N_4250,N_3527,N_3869);
nand U4251 (N_4251,N_3347,N_3270);
nand U4252 (N_4252,N_3153,N_3710);
or U4253 (N_4253,N_3492,N_3525);
nor U4254 (N_4254,N_3805,N_3679);
or U4255 (N_4255,N_3522,N_3964);
nor U4256 (N_4256,N_3654,N_3998);
nor U4257 (N_4257,N_3097,N_3560);
nand U4258 (N_4258,N_3643,N_3655);
xor U4259 (N_4259,N_3326,N_3587);
nor U4260 (N_4260,N_3835,N_3652);
or U4261 (N_4261,N_3304,N_3973);
and U4262 (N_4262,N_3924,N_3870);
and U4263 (N_4263,N_3117,N_3336);
nor U4264 (N_4264,N_3268,N_3388);
nand U4265 (N_4265,N_3305,N_3518);
and U4266 (N_4266,N_3932,N_3839);
nand U4267 (N_4267,N_3578,N_3038);
and U4268 (N_4268,N_3016,N_3885);
or U4269 (N_4269,N_3284,N_3055);
or U4270 (N_4270,N_3580,N_3144);
xnor U4271 (N_4271,N_3050,N_3856);
nor U4272 (N_4272,N_3647,N_3984);
and U4273 (N_4273,N_3325,N_3776);
nand U4274 (N_4274,N_3469,N_3282);
and U4275 (N_4275,N_3500,N_3561);
and U4276 (N_4276,N_3586,N_3453);
nand U4277 (N_4277,N_3267,N_3888);
and U4278 (N_4278,N_3105,N_3312);
nand U4279 (N_4279,N_3171,N_3082);
xor U4280 (N_4280,N_3148,N_3866);
or U4281 (N_4281,N_3478,N_3232);
or U4282 (N_4282,N_3005,N_3119);
and U4283 (N_4283,N_3429,N_3988);
and U4284 (N_4284,N_3329,N_3302);
and U4285 (N_4285,N_3409,N_3909);
nand U4286 (N_4286,N_3406,N_3697);
nand U4287 (N_4287,N_3841,N_3180);
or U4288 (N_4288,N_3969,N_3918);
nand U4289 (N_4289,N_3557,N_3604);
nand U4290 (N_4290,N_3896,N_3880);
and U4291 (N_4291,N_3058,N_3723);
and U4292 (N_4292,N_3968,N_3881);
and U4293 (N_4293,N_3672,N_3703);
nand U4294 (N_4294,N_3961,N_3761);
and U4295 (N_4295,N_3786,N_3645);
xnor U4296 (N_4296,N_3024,N_3619);
nand U4297 (N_4297,N_3544,N_3983);
or U4298 (N_4298,N_3419,N_3139);
and U4299 (N_4299,N_3689,N_3460);
or U4300 (N_4300,N_3771,N_3616);
or U4301 (N_4301,N_3734,N_3380);
nand U4302 (N_4302,N_3065,N_3759);
nand U4303 (N_4303,N_3439,N_3021);
and U4304 (N_4304,N_3106,N_3599);
nand U4305 (N_4305,N_3629,N_3588);
or U4306 (N_4306,N_3258,N_3474);
and U4307 (N_4307,N_3972,N_3314);
nand U4308 (N_4308,N_3495,N_3907);
and U4309 (N_4309,N_3313,N_3945);
or U4310 (N_4310,N_3615,N_3642);
xor U4311 (N_4311,N_3958,N_3197);
or U4312 (N_4312,N_3739,N_3772);
nor U4313 (N_4313,N_3702,N_3513);
or U4314 (N_4314,N_3651,N_3009);
and U4315 (N_4315,N_3047,N_3788);
nand U4316 (N_4316,N_3558,N_3420);
or U4317 (N_4317,N_3480,N_3446);
and U4318 (N_4318,N_3324,N_3080);
nor U4319 (N_4319,N_3763,N_3414);
and U4320 (N_4320,N_3228,N_3842);
or U4321 (N_4321,N_3549,N_3064);
or U4322 (N_4322,N_3813,N_3333);
or U4323 (N_4323,N_3528,N_3530);
nor U4324 (N_4324,N_3014,N_3002);
xor U4325 (N_4325,N_3332,N_3318);
nand U4326 (N_4326,N_3415,N_3471);
and U4327 (N_4327,N_3400,N_3123);
nor U4328 (N_4328,N_3742,N_3910);
nor U4329 (N_4329,N_3873,N_3754);
nand U4330 (N_4330,N_3094,N_3410);
xor U4331 (N_4331,N_3274,N_3054);
or U4332 (N_4332,N_3927,N_3156);
and U4333 (N_4333,N_3837,N_3596);
and U4334 (N_4334,N_3956,N_3372);
nor U4335 (N_4335,N_3768,N_3236);
xnor U4336 (N_4336,N_3281,N_3166);
nor U4337 (N_4337,N_3396,N_3362);
xor U4338 (N_4338,N_3612,N_3456);
or U4339 (N_4339,N_3891,N_3833);
xnor U4340 (N_4340,N_3951,N_3845);
nor U4341 (N_4341,N_3935,N_3593);
nor U4342 (N_4342,N_3135,N_3458);
or U4343 (N_4343,N_3448,N_3603);
or U4344 (N_4344,N_3598,N_3417);
xnor U4345 (N_4345,N_3708,N_3221);
or U4346 (N_4346,N_3662,N_3291);
xnor U4347 (N_4347,N_3823,N_3323);
and U4348 (N_4348,N_3801,N_3674);
or U4349 (N_4349,N_3049,N_3676);
and U4350 (N_4350,N_3934,N_3462);
or U4351 (N_4351,N_3397,N_3632);
and U4352 (N_4352,N_3085,N_3787);
xnor U4353 (N_4353,N_3416,N_3289);
xor U4354 (N_4354,N_3395,N_3476);
or U4355 (N_4355,N_3637,N_3752);
nor U4356 (N_4356,N_3012,N_3036);
nand U4357 (N_4357,N_3023,N_3605);
nand U4358 (N_4358,N_3373,N_3433);
nor U4359 (N_4359,N_3490,N_3535);
nor U4360 (N_4360,N_3540,N_3116);
or U4361 (N_4361,N_3216,N_3295);
and U4362 (N_4362,N_3203,N_3872);
or U4363 (N_4363,N_3568,N_3581);
or U4364 (N_4364,N_3401,N_3337);
and U4365 (N_4365,N_3250,N_3831);
and U4366 (N_4366,N_3158,N_3933);
nand U4367 (N_4367,N_3997,N_3551);
and U4368 (N_4368,N_3793,N_3132);
nand U4369 (N_4369,N_3146,N_3125);
xnor U4370 (N_4370,N_3441,N_3874);
or U4371 (N_4371,N_3970,N_3031);
and U4372 (N_4372,N_3854,N_3916);
or U4373 (N_4373,N_3744,N_3481);
and U4374 (N_4374,N_3214,N_3251);
nand U4375 (N_4375,N_3765,N_3306);
and U4376 (N_4376,N_3836,N_3678);
xor U4377 (N_4377,N_3384,N_3437);
nor U4378 (N_4378,N_3684,N_3224);
nor U4379 (N_4379,N_3838,N_3053);
or U4380 (N_4380,N_3457,N_3272);
or U4381 (N_4381,N_3195,N_3249);
nor U4382 (N_4382,N_3519,N_3766);
and U4383 (N_4383,N_3403,N_3013);
or U4384 (N_4384,N_3901,N_3348);
nor U4385 (N_4385,N_3520,N_3387);
or U4386 (N_4386,N_3681,N_3254);
nand U4387 (N_4387,N_3719,N_3011);
xor U4388 (N_4388,N_3229,N_3320);
nand U4389 (N_4389,N_3237,N_3531);
and U4390 (N_4390,N_3720,N_3052);
nor U4391 (N_4391,N_3572,N_3231);
nor U4392 (N_4392,N_3502,N_3940);
and U4393 (N_4393,N_3159,N_3898);
nor U4394 (N_4394,N_3566,N_3092);
xnor U4395 (N_4395,N_3698,N_3746);
nor U4396 (N_4396,N_3640,N_3432);
and U4397 (N_4397,N_3925,N_3548);
nand U4398 (N_4398,N_3485,N_3609);
xnor U4399 (N_4399,N_3677,N_3133);
xor U4400 (N_4400,N_3921,N_3455);
or U4401 (N_4401,N_3042,N_3252);
nor U4402 (N_4402,N_3579,N_3621);
or U4403 (N_4403,N_3584,N_3670);
xnor U4404 (N_4404,N_3668,N_3028);
and U4405 (N_4405,N_3467,N_3190);
nand U4406 (N_4406,N_3493,N_3701);
nand U4407 (N_4407,N_3571,N_3245);
nand U4408 (N_4408,N_3164,N_3711);
nor U4409 (N_4409,N_3764,N_3630);
nor U4410 (N_4410,N_3246,N_3623);
or U4411 (N_4411,N_3620,N_3059);
or U4412 (N_4412,N_3804,N_3979);
or U4413 (N_4413,N_3178,N_3673);
or U4414 (N_4414,N_3436,N_3287);
nor U4415 (N_4415,N_3592,N_3235);
xnor U4416 (N_4416,N_3709,N_3852);
nor U4417 (N_4417,N_3807,N_3181);
nor U4418 (N_4418,N_3532,N_3790);
nor U4419 (N_4419,N_3738,N_3201);
and U4420 (N_4420,N_3212,N_3501);
and U4421 (N_4421,N_3726,N_3808);
xor U4422 (N_4422,N_3408,N_3470);
nand U4423 (N_4423,N_3048,N_3240);
or U4424 (N_4424,N_3890,N_3913);
xnor U4425 (N_4425,N_3177,N_3170);
nor U4426 (N_4426,N_3127,N_3559);
nor U4427 (N_4427,N_3883,N_3595);
nor U4428 (N_4428,N_3464,N_3218);
and U4429 (N_4429,N_3483,N_3785);
nand U4430 (N_4430,N_3263,N_3825);
xnor U4431 (N_4431,N_3041,N_3443);
or U4432 (N_4432,N_3130,N_3425);
and U4433 (N_4433,N_3209,N_3569);
nand U4434 (N_4434,N_3919,N_3169);
or U4435 (N_4435,N_3019,N_3421);
and U4436 (N_4436,N_3855,N_3445);
and U4437 (N_4437,N_3730,N_3463);
nor U4438 (N_4438,N_3482,N_3796);
xor U4439 (N_4439,N_3990,N_3354);
and U4440 (N_4440,N_3685,N_3168);
nand U4441 (N_4441,N_3062,N_3846);
nand U4442 (N_4442,N_3797,N_3392);
or U4443 (N_4443,N_3255,N_3278);
nand U4444 (N_4444,N_3391,N_3364);
nand U4445 (N_4445,N_3163,N_3034);
or U4446 (N_4446,N_3262,N_3565);
and U4447 (N_4447,N_3486,N_3057);
nor U4448 (N_4448,N_3109,N_3067);
xnor U4449 (N_4449,N_3550,N_3660);
nor U4450 (N_4450,N_3828,N_3682);
xor U4451 (N_4451,N_3378,N_3585);
nand U4452 (N_4452,N_3046,N_3369);
xnor U4453 (N_4453,N_3210,N_3340);
xor U4454 (N_4454,N_3900,N_3230);
nor U4455 (N_4455,N_3301,N_3200);
nand U4456 (N_4456,N_3892,N_3376);
nor U4457 (N_4457,N_3374,N_3626);
nor U4458 (N_4458,N_3692,N_3145);
nor U4459 (N_4459,N_3638,N_3816);
nand U4460 (N_4460,N_3735,N_3928);
nand U4461 (N_4461,N_3567,N_3360);
nor U4462 (N_4462,N_3078,N_3960);
and U4463 (N_4463,N_3955,N_3315);
nand U4464 (N_4464,N_3849,N_3705);
or U4465 (N_4465,N_3863,N_3728);
nand U4466 (N_4466,N_3327,N_3704);
nand U4467 (N_4467,N_3147,N_3812);
and U4468 (N_4468,N_3792,N_3344);
xnor U4469 (N_4469,N_3714,N_3810);
nand U4470 (N_4470,N_3737,N_3641);
or U4471 (N_4471,N_3427,N_3715);
xnor U4472 (N_4472,N_3926,N_3339);
and U4473 (N_4473,N_3649,N_3102);
xnor U4474 (N_4474,N_3613,N_3971);
or U4475 (N_4475,N_3779,N_3022);
nand U4476 (N_4476,N_3635,N_3297);
and U4477 (N_4477,N_3095,N_3745);
nor U4478 (N_4478,N_3411,N_3276);
nor U4479 (N_4479,N_3385,N_3176);
nand U4480 (N_4480,N_3027,N_3345);
nor U4481 (N_4481,N_3389,N_3784);
nor U4482 (N_4482,N_3226,N_3006);
nor U4483 (N_4483,N_3902,N_3303);
or U4484 (N_4484,N_3611,N_3114);
and U4485 (N_4485,N_3589,N_3083);
or U4486 (N_4486,N_3975,N_3126);
nor U4487 (N_4487,N_3959,N_3288);
and U4488 (N_4488,N_3536,N_3174);
or U4489 (N_4489,N_3695,N_3978);
or U4490 (N_4490,N_3498,N_3669);
and U4491 (N_4491,N_3343,N_3911);
nor U4492 (N_4492,N_3829,N_3077);
nand U4493 (N_4493,N_3350,N_3363);
or U4494 (N_4494,N_3783,N_3511);
nor U4495 (N_4495,N_3712,N_3141);
xor U4496 (N_4496,N_3438,N_3556);
xnor U4497 (N_4497,N_3283,N_3553);
nor U4498 (N_4498,N_3529,N_3007);
nor U4499 (N_4499,N_3777,N_3424);
xor U4500 (N_4500,N_3220,N_3704);
xnor U4501 (N_4501,N_3392,N_3547);
nand U4502 (N_4502,N_3704,N_3924);
and U4503 (N_4503,N_3916,N_3177);
nor U4504 (N_4504,N_3017,N_3309);
nand U4505 (N_4505,N_3871,N_3559);
xor U4506 (N_4506,N_3245,N_3110);
nor U4507 (N_4507,N_3519,N_3842);
xnor U4508 (N_4508,N_3238,N_3699);
nand U4509 (N_4509,N_3678,N_3573);
nand U4510 (N_4510,N_3368,N_3990);
nand U4511 (N_4511,N_3181,N_3866);
and U4512 (N_4512,N_3977,N_3679);
nor U4513 (N_4513,N_3197,N_3972);
or U4514 (N_4514,N_3066,N_3661);
nand U4515 (N_4515,N_3492,N_3022);
and U4516 (N_4516,N_3685,N_3867);
or U4517 (N_4517,N_3772,N_3504);
nand U4518 (N_4518,N_3933,N_3909);
nand U4519 (N_4519,N_3277,N_3321);
or U4520 (N_4520,N_3412,N_3437);
and U4521 (N_4521,N_3897,N_3104);
nor U4522 (N_4522,N_3825,N_3457);
xnor U4523 (N_4523,N_3756,N_3008);
or U4524 (N_4524,N_3212,N_3401);
or U4525 (N_4525,N_3792,N_3922);
nor U4526 (N_4526,N_3570,N_3870);
or U4527 (N_4527,N_3618,N_3714);
xnor U4528 (N_4528,N_3285,N_3763);
or U4529 (N_4529,N_3327,N_3422);
or U4530 (N_4530,N_3135,N_3487);
nor U4531 (N_4531,N_3485,N_3154);
nand U4532 (N_4532,N_3021,N_3469);
nor U4533 (N_4533,N_3061,N_3962);
xor U4534 (N_4534,N_3230,N_3597);
nor U4535 (N_4535,N_3870,N_3331);
nor U4536 (N_4536,N_3284,N_3406);
nand U4537 (N_4537,N_3986,N_3879);
nand U4538 (N_4538,N_3268,N_3846);
nand U4539 (N_4539,N_3311,N_3752);
nand U4540 (N_4540,N_3851,N_3522);
nor U4541 (N_4541,N_3826,N_3062);
xnor U4542 (N_4542,N_3035,N_3684);
nor U4543 (N_4543,N_3767,N_3650);
or U4544 (N_4544,N_3208,N_3248);
nand U4545 (N_4545,N_3699,N_3423);
and U4546 (N_4546,N_3645,N_3547);
nor U4547 (N_4547,N_3487,N_3646);
nor U4548 (N_4548,N_3209,N_3985);
xnor U4549 (N_4549,N_3682,N_3801);
nand U4550 (N_4550,N_3206,N_3088);
nand U4551 (N_4551,N_3291,N_3297);
and U4552 (N_4552,N_3485,N_3649);
or U4553 (N_4553,N_3562,N_3314);
and U4554 (N_4554,N_3701,N_3860);
nor U4555 (N_4555,N_3788,N_3069);
nand U4556 (N_4556,N_3394,N_3009);
nand U4557 (N_4557,N_3762,N_3320);
or U4558 (N_4558,N_3861,N_3895);
or U4559 (N_4559,N_3312,N_3168);
or U4560 (N_4560,N_3686,N_3693);
or U4561 (N_4561,N_3777,N_3526);
or U4562 (N_4562,N_3549,N_3771);
and U4563 (N_4563,N_3236,N_3584);
nand U4564 (N_4564,N_3962,N_3636);
xor U4565 (N_4565,N_3020,N_3633);
xor U4566 (N_4566,N_3535,N_3428);
xnor U4567 (N_4567,N_3159,N_3228);
and U4568 (N_4568,N_3222,N_3466);
xnor U4569 (N_4569,N_3609,N_3465);
nand U4570 (N_4570,N_3961,N_3027);
and U4571 (N_4571,N_3329,N_3227);
nor U4572 (N_4572,N_3075,N_3927);
or U4573 (N_4573,N_3761,N_3641);
nor U4574 (N_4574,N_3708,N_3843);
xnor U4575 (N_4575,N_3036,N_3576);
nand U4576 (N_4576,N_3764,N_3908);
nor U4577 (N_4577,N_3309,N_3396);
xor U4578 (N_4578,N_3001,N_3940);
and U4579 (N_4579,N_3367,N_3179);
and U4580 (N_4580,N_3266,N_3619);
or U4581 (N_4581,N_3274,N_3183);
nand U4582 (N_4582,N_3464,N_3066);
xor U4583 (N_4583,N_3507,N_3288);
or U4584 (N_4584,N_3379,N_3254);
and U4585 (N_4585,N_3857,N_3454);
nor U4586 (N_4586,N_3225,N_3520);
and U4587 (N_4587,N_3358,N_3215);
nand U4588 (N_4588,N_3072,N_3902);
or U4589 (N_4589,N_3156,N_3477);
xnor U4590 (N_4590,N_3347,N_3497);
and U4591 (N_4591,N_3287,N_3820);
nand U4592 (N_4592,N_3832,N_3300);
xnor U4593 (N_4593,N_3161,N_3016);
xnor U4594 (N_4594,N_3116,N_3114);
or U4595 (N_4595,N_3041,N_3885);
or U4596 (N_4596,N_3485,N_3580);
xor U4597 (N_4597,N_3138,N_3424);
nand U4598 (N_4598,N_3071,N_3872);
nor U4599 (N_4599,N_3462,N_3793);
xor U4600 (N_4600,N_3131,N_3510);
nand U4601 (N_4601,N_3881,N_3267);
or U4602 (N_4602,N_3417,N_3238);
and U4603 (N_4603,N_3760,N_3648);
xnor U4604 (N_4604,N_3359,N_3271);
and U4605 (N_4605,N_3258,N_3788);
and U4606 (N_4606,N_3054,N_3710);
xnor U4607 (N_4607,N_3025,N_3074);
nor U4608 (N_4608,N_3768,N_3454);
nand U4609 (N_4609,N_3051,N_3150);
nor U4610 (N_4610,N_3005,N_3905);
xor U4611 (N_4611,N_3234,N_3692);
nor U4612 (N_4612,N_3544,N_3794);
or U4613 (N_4613,N_3938,N_3741);
nor U4614 (N_4614,N_3390,N_3858);
or U4615 (N_4615,N_3519,N_3251);
and U4616 (N_4616,N_3380,N_3462);
xor U4617 (N_4617,N_3677,N_3988);
nand U4618 (N_4618,N_3350,N_3980);
nand U4619 (N_4619,N_3630,N_3012);
nand U4620 (N_4620,N_3517,N_3572);
xor U4621 (N_4621,N_3852,N_3180);
nor U4622 (N_4622,N_3015,N_3364);
xor U4623 (N_4623,N_3088,N_3984);
and U4624 (N_4624,N_3258,N_3703);
and U4625 (N_4625,N_3403,N_3889);
nand U4626 (N_4626,N_3445,N_3075);
or U4627 (N_4627,N_3625,N_3392);
nor U4628 (N_4628,N_3303,N_3350);
or U4629 (N_4629,N_3298,N_3560);
xor U4630 (N_4630,N_3408,N_3193);
or U4631 (N_4631,N_3631,N_3501);
nand U4632 (N_4632,N_3001,N_3665);
xnor U4633 (N_4633,N_3420,N_3606);
and U4634 (N_4634,N_3614,N_3146);
nand U4635 (N_4635,N_3434,N_3541);
and U4636 (N_4636,N_3571,N_3660);
and U4637 (N_4637,N_3357,N_3097);
xor U4638 (N_4638,N_3260,N_3098);
and U4639 (N_4639,N_3339,N_3688);
and U4640 (N_4640,N_3130,N_3347);
xnor U4641 (N_4641,N_3821,N_3007);
and U4642 (N_4642,N_3893,N_3705);
nor U4643 (N_4643,N_3832,N_3622);
or U4644 (N_4644,N_3935,N_3336);
xor U4645 (N_4645,N_3655,N_3984);
and U4646 (N_4646,N_3849,N_3057);
or U4647 (N_4647,N_3048,N_3056);
nand U4648 (N_4648,N_3547,N_3365);
or U4649 (N_4649,N_3787,N_3205);
nor U4650 (N_4650,N_3649,N_3595);
nor U4651 (N_4651,N_3148,N_3874);
xor U4652 (N_4652,N_3580,N_3373);
or U4653 (N_4653,N_3608,N_3222);
nor U4654 (N_4654,N_3158,N_3284);
or U4655 (N_4655,N_3070,N_3662);
and U4656 (N_4656,N_3937,N_3856);
nor U4657 (N_4657,N_3669,N_3808);
and U4658 (N_4658,N_3889,N_3439);
and U4659 (N_4659,N_3863,N_3843);
and U4660 (N_4660,N_3290,N_3815);
nor U4661 (N_4661,N_3920,N_3470);
and U4662 (N_4662,N_3569,N_3984);
nand U4663 (N_4663,N_3926,N_3808);
xor U4664 (N_4664,N_3984,N_3245);
and U4665 (N_4665,N_3000,N_3940);
and U4666 (N_4666,N_3377,N_3413);
nand U4667 (N_4667,N_3175,N_3331);
xnor U4668 (N_4668,N_3114,N_3184);
and U4669 (N_4669,N_3872,N_3488);
xor U4670 (N_4670,N_3132,N_3925);
nor U4671 (N_4671,N_3077,N_3630);
or U4672 (N_4672,N_3267,N_3744);
xor U4673 (N_4673,N_3063,N_3248);
xor U4674 (N_4674,N_3999,N_3250);
and U4675 (N_4675,N_3222,N_3472);
nor U4676 (N_4676,N_3054,N_3221);
nor U4677 (N_4677,N_3714,N_3109);
and U4678 (N_4678,N_3837,N_3879);
and U4679 (N_4679,N_3527,N_3037);
nand U4680 (N_4680,N_3870,N_3339);
and U4681 (N_4681,N_3053,N_3716);
xor U4682 (N_4682,N_3343,N_3265);
or U4683 (N_4683,N_3204,N_3868);
nor U4684 (N_4684,N_3800,N_3316);
and U4685 (N_4685,N_3739,N_3956);
nand U4686 (N_4686,N_3716,N_3179);
xor U4687 (N_4687,N_3365,N_3924);
or U4688 (N_4688,N_3833,N_3362);
xnor U4689 (N_4689,N_3428,N_3055);
or U4690 (N_4690,N_3911,N_3734);
nand U4691 (N_4691,N_3152,N_3176);
nor U4692 (N_4692,N_3070,N_3749);
xor U4693 (N_4693,N_3936,N_3466);
nor U4694 (N_4694,N_3692,N_3208);
or U4695 (N_4695,N_3821,N_3278);
nor U4696 (N_4696,N_3436,N_3260);
xor U4697 (N_4697,N_3204,N_3166);
and U4698 (N_4698,N_3970,N_3813);
nand U4699 (N_4699,N_3939,N_3475);
xnor U4700 (N_4700,N_3287,N_3021);
or U4701 (N_4701,N_3611,N_3927);
nor U4702 (N_4702,N_3252,N_3327);
xor U4703 (N_4703,N_3485,N_3162);
nor U4704 (N_4704,N_3154,N_3028);
xor U4705 (N_4705,N_3537,N_3484);
xor U4706 (N_4706,N_3074,N_3784);
nor U4707 (N_4707,N_3808,N_3106);
nand U4708 (N_4708,N_3973,N_3987);
nand U4709 (N_4709,N_3477,N_3496);
xor U4710 (N_4710,N_3947,N_3973);
and U4711 (N_4711,N_3524,N_3648);
xor U4712 (N_4712,N_3351,N_3787);
xnor U4713 (N_4713,N_3980,N_3203);
and U4714 (N_4714,N_3700,N_3119);
or U4715 (N_4715,N_3492,N_3344);
nand U4716 (N_4716,N_3578,N_3553);
nand U4717 (N_4717,N_3626,N_3341);
or U4718 (N_4718,N_3049,N_3270);
or U4719 (N_4719,N_3650,N_3591);
xor U4720 (N_4720,N_3829,N_3859);
or U4721 (N_4721,N_3136,N_3178);
nor U4722 (N_4722,N_3281,N_3976);
xnor U4723 (N_4723,N_3753,N_3813);
and U4724 (N_4724,N_3767,N_3792);
nand U4725 (N_4725,N_3159,N_3341);
and U4726 (N_4726,N_3205,N_3418);
and U4727 (N_4727,N_3452,N_3702);
or U4728 (N_4728,N_3855,N_3641);
nor U4729 (N_4729,N_3692,N_3589);
nand U4730 (N_4730,N_3391,N_3040);
nor U4731 (N_4731,N_3500,N_3910);
and U4732 (N_4732,N_3362,N_3505);
nor U4733 (N_4733,N_3603,N_3466);
nor U4734 (N_4734,N_3291,N_3226);
nand U4735 (N_4735,N_3869,N_3719);
nand U4736 (N_4736,N_3611,N_3701);
nor U4737 (N_4737,N_3707,N_3251);
and U4738 (N_4738,N_3718,N_3173);
xor U4739 (N_4739,N_3793,N_3447);
nor U4740 (N_4740,N_3697,N_3945);
or U4741 (N_4741,N_3570,N_3730);
xnor U4742 (N_4742,N_3555,N_3282);
or U4743 (N_4743,N_3011,N_3770);
or U4744 (N_4744,N_3578,N_3284);
and U4745 (N_4745,N_3939,N_3248);
nor U4746 (N_4746,N_3683,N_3769);
or U4747 (N_4747,N_3541,N_3299);
nand U4748 (N_4748,N_3827,N_3531);
or U4749 (N_4749,N_3471,N_3448);
xnor U4750 (N_4750,N_3298,N_3266);
or U4751 (N_4751,N_3999,N_3783);
xor U4752 (N_4752,N_3625,N_3049);
xor U4753 (N_4753,N_3165,N_3898);
and U4754 (N_4754,N_3222,N_3922);
or U4755 (N_4755,N_3174,N_3348);
nor U4756 (N_4756,N_3260,N_3873);
xnor U4757 (N_4757,N_3030,N_3578);
xnor U4758 (N_4758,N_3150,N_3456);
or U4759 (N_4759,N_3975,N_3540);
nand U4760 (N_4760,N_3263,N_3990);
nand U4761 (N_4761,N_3818,N_3572);
xnor U4762 (N_4762,N_3435,N_3789);
nor U4763 (N_4763,N_3657,N_3133);
nand U4764 (N_4764,N_3366,N_3558);
nor U4765 (N_4765,N_3602,N_3027);
or U4766 (N_4766,N_3165,N_3773);
nand U4767 (N_4767,N_3686,N_3594);
and U4768 (N_4768,N_3424,N_3720);
or U4769 (N_4769,N_3155,N_3905);
xnor U4770 (N_4770,N_3055,N_3700);
nand U4771 (N_4771,N_3827,N_3687);
nand U4772 (N_4772,N_3611,N_3925);
nor U4773 (N_4773,N_3795,N_3267);
xnor U4774 (N_4774,N_3501,N_3473);
or U4775 (N_4775,N_3054,N_3114);
xnor U4776 (N_4776,N_3454,N_3537);
or U4777 (N_4777,N_3343,N_3160);
xor U4778 (N_4778,N_3614,N_3436);
nor U4779 (N_4779,N_3116,N_3167);
xor U4780 (N_4780,N_3355,N_3998);
or U4781 (N_4781,N_3705,N_3709);
nor U4782 (N_4782,N_3876,N_3279);
or U4783 (N_4783,N_3783,N_3434);
or U4784 (N_4784,N_3828,N_3485);
and U4785 (N_4785,N_3939,N_3511);
or U4786 (N_4786,N_3778,N_3214);
or U4787 (N_4787,N_3385,N_3075);
nor U4788 (N_4788,N_3312,N_3956);
and U4789 (N_4789,N_3239,N_3689);
or U4790 (N_4790,N_3576,N_3683);
nand U4791 (N_4791,N_3859,N_3432);
nor U4792 (N_4792,N_3728,N_3044);
and U4793 (N_4793,N_3485,N_3297);
nor U4794 (N_4794,N_3755,N_3437);
nand U4795 (N_4795,N_3902,N_3979);
nor U4796 (N_4796,N_3266,N_3647);
xnor U4797 (N_4797,N_3454,N_3684);
or U4798 (N_4798,N_3303,N_3814);
xnor U4799 (N_4799,N_3082,N_3464);
nor U4800 (N_4800,N_3853,N_3906);
or U4801 (N_4801,N_3717,N_3436);
xnor U4802 (N_4802,N_3729,N_3621);
or U4803 (N_4803,N_3641,N_3038);
nand U4804 (N_4804,N_3605,N_3636);
xnor U4805 (N_4805,N_3542,N_3167);
nor U4806 (N_4806,N_3130,N_3301);
or U4807 (N_4807,N_3891,N_3766);
and U4808 (N_4808,N_3587,N_3734);
nand U4809 (N_4809,N_3332,N_3566);
nand U4810 (N_4810,N_3532,N_3876);
nor U4811 (N_4811,N_3785,N_3782);
nor U4812 (N_4812,N_3887,N_3150);
nor U4813 (N_4813,N_3307,N_3525);
and U4814 (N_4814,N_3820,N_3749);
xor U4815 (N_4815,N_3909,N_3590);
nand U4816 (N_4816,N_3462,N_3127);
nor U4817 (N_4817,N_3973,N_3591);
nor U4818 (N_4818,N_3639,N_3897);
and U4819 (N_4819,N_3264,N_3976);
nor U4820 (N_4820,N_3711,N_3511);
and U4821 (N_4821,N_3791,N_3738);
and U4822 (N_4822,N_3998,N_3314);
xnor U4823 (N_4823,N_3350,N_3923);
nand U4824 (N_4824,N_3772,N_3717);
xor U4825 (N_4825,N_3501,N_3779);
xor U4826 (N_4826,N_3504,N_3507);
xnor U4827 (N_4827,N_3623,N_3114);
xor U4828 (N_4828,N_3291,N_3346);
or U4829 (N_4829,N_3894,N_3046);
xnor U4830 (N_4830,N_3470,N_3585);
and U4831 (N_4831,N_3197,N_3561);
xnor U4832 (N_4832,N_3797,N_3939);
nand U4833 (N_4833,N_3697,N_3925);
nand U4834 (N_4834,N_3343,N_3330);
or U4835 (N_4835,N_3581,N_3747);
and U4836 (N_4836,N_3183,N_3791);
xnor U4837 (N_4837,N_3097,N_3553);
nor U4838 (N_4838,N_3254,N_3441);
or U4839 (N_4839,N_3805,N_3375);
nor U4840 (N_4840,N_3982,N_3679);
and U4841 (N_4841,N_3600,N_3536);
xnor U4842 (N_4842,N_3319,N_3712);
xor U4843 (N_4843,N_3131,N_3296);
and U4844 (N_4844,N_3191,N_3712);
and U4845 (N_4845,N_3602,N_3343);
xor U4846 (N_4846,N_3566,N_3105);
or U4847 (N_4847,N_3696,N_3880);
nand U4848 (N_4848,N_3037,N_3857);
and U4849 (N_4849,N_3128,N_3345);
xor U4850 (N_4850,N_3553,N_3152);
nand U4851 (N_4851,N_3975,N_3916);
nand U4852 (N_4852,N_3264,N_3409);
and U4853 (N_4853,N_3181,N_3789);
nor U4854 (N_4854,N_3385,N_3522);
or U4855 (N_4855,N_3916,N_3139);
or U4856 (N_4856,N_3627,N_3885);
nand U4857 (N_4857,N_3799,N_3275);
xor U4858 (N_4858,N_3061,N_3933);
or U4859 (N_4859,N_3710,N_3256);
xnor U4860 (N_4860,N_3425,N_3807);
and U4861 (N_4861,N_3772,N_3056);
or U4862 (N_4862,N_3817,N_3584);
or U4863 (N_4863,N_3042,N_3139);
nor U4864 (N_4864,N_3281,N_3899);
or U4865 (N_4865,N_3218,N_3037);
xnor U4866 (N_4866,N_3718,N_3473);
and U4867 (N_4867,N_3712,N_3746);
nand U4868 (N_4868,N_3203,N_3132);
xnor U4869 (N_4869,N_3130,N_3001);
and U4870 (N_4870,N_3669,N_3956);
or U4871 (N_4871,N_3229,N_3817);
xor U4872 (N_4872,N_3085,N_3531);
nor U4873 (N_4873,N_3737,N_3480);
or U4874 (N_4874,N_3092,N_3048);
or U4875 (N_4875,N_3230,N_3883);
nor U4876 (N_4876,N_3106,N_3240);
nor U4877 (N_4877,N_3175,N_3337);
nand U4878 (N_4878,N_3178,N_3645);
xnor U4879 (N_4879,N_3913,N_3216);
and U4880 (N_4880,N_3241,N_3408);
nor U4881 (N_4881,N_3450,N_3427);
or U4882 (N_4882,N_3356,N_3738);
or U4883 (N_4883,N_3095,N_3492);
or U4884 (N_4884,N_3298,N_3508);
nand U4885 (N_4885,N_3079,N_3546);
or U4886 (N_4886,N_3112,N_3903);
and U4887 (N_4887,N_3813,N_3745);
or U4888 (N_4888,N_3918,N_3190);
and U4889 (N_4889,N_3077,N_3014);
xor U4890 (N_4890,N_3288,N_3116);
nand U4891 (N_4891,N_3881,N_3701);
and U4892 (N_4892,N_3731,N_3033);
xnor U4893 (N_4893,N_3143,N_3732);
xnor U4894 (N_4894,N_3356,N_3352);
or U4895 (N_4895,N_3956,N_3069);
nand U4896 (N_4896,N_3228,N_3683);
and U4897 (N_4897,N_3989,N_3314);
nand U4898 (N_4898,N_3913,N_3694);
nand U4899 (N_4899,N_3808,N_3364);
nand U4900 (N_4900,N_3437,N_3669);
xor U4901 (N_4901,N_3640,N_3630);
xor U4902 (N_4902,N_3215,N_3239);
nand U4903 (N_4903,N_3292,N_3074);
nand U4904 (N_4904,N_3607,N_3008);
and U4905 (N_4905,N_3126,N_3056);
or U4906 (N_4906,N_3330,N_3293);
nor U4907 (N_4907,N_3231,N_3165);
xnor U4908 (N_4908,N_3212,N_3295);
nand U4909 (N_4909,N_3676,N_3579);
xnor U4910 (N_4910,N_3484,N_3008);
or U4911 (N_4911,N_3869,N_3903);
and U4912 (N_4912,N_3216,N_3742);
nor U4913 (N_4913,N_3111,N_3294);
and U4914 (N_4914,N_3855,N_3371);
or U4915 (N_4915,N_3709,N_3841);
xor U4916 (N_4916,N_3274,N_3867);
or U4917 (N_4917,N_3597,N_3111);
nor U4918 (N_4918,N_3136,N_3608);
and U4919 (N_4919,N_3871,N_3902);
xor U4920 (N_4920,N_3537,N_3814);
or U4921 (N_4921,N_3027,N_3957);
nand U4922 (N_4922,N_3329,N_3919);
nand U4923 (N_4923,N_3664,N_3414);
nor U4924 (N_4924,N_3162,N_3033);
or U4925 (N_4925,N_3238,N_3914);
xnor U4926 (N_4926,N_3284,N_3719);
nor U4927 (N_4927,N_3032,N_3135);
and U4928 (N_4928,N_3628,N_3649);
nor U4929 (N_4929,N_3223,N_3329);
and U4930 (N_4930,N_3324,N_3000);
or U4931 (N_4931,N_3380,N_3648);
nor U4932 (N_4932,N_3915,N_3954);
or U4933 (N_4933,N_3650,N_3865);
and U4934 (N_4934,N_3514,N_3763);
or U4935 (N_4935,N_3508,N_3814);
xnor U4936 (N_4936,N_3397,N_3280);
and U4937 (N_4937,N_3499,N_3570);
nand U4938 (N_4938,N_3757,N_3908);
or U4939 (N_4939,N_3332,N_3420);
or U4940 (N_4940,N_3291,N_3947);
nand U4941 (N_4941,N_3947,N_3424);
nand U4942 (N_4942,N_3486,N_3024);
xnor U4943 (N_4943,N_3258,N_3153);
or U4944 (N_4944,N_3104,N_3789);
and U4945 (N_4945,N_3584,N_3747);
nor U4946 (N_4946,N_3248,N_3226);
or U4947 (N_4947,N_3767,N_3797);
xnor U4948 (N_4948,N_3104,N_3144);
xnor U4949 (N_4949,N_3488,N_3826);
and U4950 (N_4950,N_3016,N_3997);
nand U4951 (N_4951,N_3940,N_3936);
xnor U4952 (N_4952,N_3717,N_3527);
nor U4953 (N_4953,N_3961,N_3497);
xnor U4954 (N_4954,N_3139,N_3780);
and U4955 (N_4955,N_3916,N_3649);
nand U4956 (N_4956,N_3182,N_3337);
and U4957 (N_4957,N_3613,N_3643);
nor U4958 (N_4958,N_3996,N_3250);
nand U4959 (N_4959,N_3131,N_3496);
xor U4960 (N_4960,N_3062,N_3889);
and U4961 (N_4961,N_3177,N_3145);
or U4962 (N_4962,N_3451,N_3152);
xnor U4963 (N_4963,N_3384,N_3363);
nand U4964 (N_4964,N_3392,N_3533);
xor U4965 (N_4965,N_3865,N_3358);
or U4966 (N_4966,N_3929,N_3977);
xor U4967 (N_4967,N_3378,N_3250);
nand U4968 (N_4968,N_3324,N_3561);
xor U4969 (N_4969,N_3793,N_3337);
or U4970 (N_4970,N_3843,N_3043);
nor U4971 (N_4971,N_3047,N_3747);
and U4972 (N_4972,N_3628,N_3657);
or U4973 (N_4973,N_3058,N_3216);
nor U4974 (N_4974,N_3646,N_3039);
nor U4975 (N_4975,N_3171,N_3927);
xnor U4976 (N_4976,N_3446,N_3645);
and U4977 (N_4977,N_3310,N_3262);
xor U4978 (N_4978,N_3442,N_3409);
nor U4979 (N_4979,N_3401,N_3308);
xor U4980 (N_4980,N_3272,N_3963);
and U4981 (N_4981,N_3722,N_3308);
xnor U4982 (N_4982,N_3701,N_3817);
and U4983 (N_4983,N_3253,N_3038);
and U4984 (N_4984,N_3032,N_3040);
or U4985 (N_4985,N_3497,N_3047);
nand U4986 (N_4986,N_3602,N_3180);
xor U4987 (N_4987,N_3333,N_3780);
nor U4988 (N_4988,N_3533,N_3812);
or U4989 (N_4989,N_3080,N_3304);
and U4990 (N_4990,N_3405,N_3053);
or U4991 (N_4991,N_3452,N_3154);
nand U4992 (N_4992,N_3545,N_3758);
xor U4993 (N_4993,N_3354,N_3366);
nor U4994 (N_4994,N_3278,N_3620);
nor U4995 (N_4995,N_3338,N_3464);
xnor U4996 (N_4996,N_3655,N_3332);
xor U4997 (N_4997,N_3126,N_3384);
and U4998 (N_4998,N_3933,N_3838);
xnor U4999 (N_4999,N_3625,N_3354);
and U5000 (N_5000,N_4347,N_4201);
nand U5001 (N_5001,N_4662,N_4616);
nand U5002 (N_5002,N_4134,N_4003);
nor U5003 (N_5003,N_4868,N_4219);
nor U5004 (N_5004,N_4486,N_4230);
and U5005 (N_5005,N_4456,N_4323);
and U5006 (N_5006,N_4995,N_4862);
nand U5007 (N_5007,N_4790,N_4850);
and U5008 (N_5008,N_4966,N_4770);
xor U5009 (N_5009,N_4418,N_4047);
nor U5010 (N_5010,N_4700,N_4978);
nand U5011 (N_5011,N_4358,N_4648);
xnor U5012 (N_5012,N_4322,N_4196);
xnor U5013 (N_5013,N_4617,N_4619);
and U5014 (N_5014,N_4846,N_4774);
xnor U5015 (N_5015,N_4404,N_4021);
or U5016 (N_5016,N_4389,N_4559);
nor U5017 (N_5017,N_4656,N_4841);
and U5018 (N_5018,N_4124,N_4554);
nor U5019 (N_5019,N_4688,N_4419);
xnor U5020 (N_5020,N_4765,N_4275);
nand U5021 (N_5021,N_4414,N_4571);
xor U5022 (N_5022,N_4564,N_4232);
nand U5023 (N_5023,N_4484,N_4033);
xnor U5024 (N_5024,N_4173,N_4022);
nand U5025 (N_5025,N_4535,N_4977);
xor U5026 (N_5026,N_4953,N_4589);
and U5027 (N_5027,N_4899,N_4957);
or U5028 (N_5028,N_4244,N_4032);
or U5029 (N_5029,N_4821,N_4290);
nand U5030 (N_5030,N_4476,N_4982);
and U5031 (N_5031,N_4612,N_4380);
nand U5032 (N_5032,N_4624,N_4939);
and U5033 (N_5033,N_4509,N_4601);
nand U5034 (N_5034,N_4831,N_4144);
nand U5035 (N_5035,N_4822,N_4816);
xnor U5036 (N_5036,N_4042,N_4407);
xor U5037 (N_5037,N_4713,N_4704);
nand U5038 (N_5038,N_4209,N_4179);
nand U5039 (N_5039,N_4193,N_4689);
xnor U5040 (N_5040,N_4388,N_4257);
xor U5041 (N_5041,N_4718,N_4216);
and U5042 (N_5042,N_4326,N_4263);
nor U5043 (N_5043,N_4301,N_4349);
xnor U5044 (N_5044,N_4408,N_4789);
nor U5045 (N_5045,N_4670,N_4501);
xor U5046 (N_5046,N_4307,N_4299);
nor U5047 (N_5047,N_4884,N_4062);
or U5048 (N_5048,N_4383,N_4785);
xor U5049 (N_5049,N_4231,N_4956);
xnor U5050 (N_5050,N_4182,N_4321);
nor U5051 (N_5051,N_4190,N_4373);
and U5052 (N_5052,N_4056,N_4813);
nor U5053 (N_5053,N_4129,N_4611);
and U5054 (N_5054,N_4253,N_4127);
nand U5055 (N_5055,N_4563,N_4913);
and U5056 (N_5056,N_4236,N_4744);
or U5057 (N_5057,N_4360,N_4210);
or U5058 (N_5058,N_4767,N_4641);
or U5059 (N_5059,N_4803,N_4320);
xor U5060 (N_5060,N_4459,N_4396);
xnor U5061 (N_5061,N_4833,N_4748);
nor U5062 (N_5062,N_4630,N_4946);
or U5063 (N_5063,N_4101,N_4915);
and U5064 (N_5064,N_4663,N_4994);
nor U5065 (N_5065,N_4806,N_4306);
and U5066 (N_5066,N_4660,N_4010);
or U5067 (N_5067,N_4579,N_4989);
nor U5068 (N_5068,N_4628,N_4873);
and U5069 (N_5069,N_4123,N_4963);
xnor U5070 (N_5070,N_4737,N_4421);
or U5071 (N_5071,N_4200,N_4888);
or U5072 (N_5072,N_4066,N_4541);
nand U5073 (N_5073,N_4023,N_4233);
xnor U5074 (N_5074,N_4511,N_4118);
or U5075 (N_5075,N_4731,N_4649);
and U5076 (N_5076,N_4981,N_4696);
xor U5077 (N_5077,N_4519,N_4657);
nand U5078 (N_5078,N_4286,N_4222);
and U5079 (N_5079,N_4152,N_4268);
and U5080 (N_5080,N_4925,N_4083);
and U5081 (N_5081,N_4131,N_4111);
nand U5082 (N_5082,N_4933,N_4531);
nand U5083 (N_5083,N_4264,N_4202);
or U5084 (N_5084,N_4712,N_4271);
nor U5085 (N_5085,N_4654,N_4824);
nor U5086 (N_5086,N_4020,N_4410);
and U5087 (N_5087,N_4783,N_4635);
xor U5088 (N_5088,N_4935,N_4413);
and U5089 (N_5089,N_4430,N_4666);
xnor U5090 (N_5090,N_4922,N_4968);
or U5091 (N_5091,N_4613,N_4415);
nor U5092 (N_5092,N_4428,N_4431);
or U5093 (N_5093,N_4840,N_4191);
or U5094 (N_5094,N_4087,N_4034);
nand U5095 (N_5095,N_4401,N_4874);
xnor U5096 (N_5096,N_4581,N_4603);
nand U5097 (N_5097,N_4221,N_4308);
xor U5098 (N_5098,N_4171,N_4830);
xor U5099 (N_5099,N_4909,N_4084);
or U5100 (N_5100,N_4183,N_4949);
and U5101 (N_5101,N_4885,N_4256);
or U5102 (N_5102,N_4204,N_4262);
nor U5103 (N_5103,N_4681,N_4335);
nor U5104 (N_5104,N_4629,N_4461);
or U5105 (N_5105,N_4610,N_4908);
or U5106 (N_5106,N_4446,N_4961);
or U5107 (N_5107,N_4467,N_4241);
and U5108 (N_5108,N_4512,N_4902);
nor U5109 (N_5109,N_4569,N_4544);
or U5110 (N_5110,N_4618,N_4832);
xor U5111 (N_5111,N_4690,N_4365);
or U5112 (N_5112,N_4845,N_4153);
and U5113 (N_5113,N_4435,N_4403);
nor U5114 (N_5114,N_4378,N_4823);
xnor U5115 (N_5115,N_4565,N_4941);
nand U5116 (N_5116,N_4354,N_4987);
nor U5117 (N_5117,N_4778,N_4776);
or U5118 (N_5118,N_4602,N_4267);
xor U5119 (N_5119,N_4441,N_4574);
and U5120 (N_5120,N_4433,N_4324);
or U5121 (N_5121,N_4537,N_4522);
xor U5122 (N_5122,N_4107,N_4856);
and U5123 (N_5123,N_4983,N_4787);
or U5124 (N_5124,N_4504,N_4438);
or U5125 (N_5125,N_4483,N_4572);
and U5126 (N_5126,N_4714,N_4515);
nor U5127 (N_5127,N_4086,N_4288);
and U5128 (N_5128,N_4708,N_4252);
or U5129 (N_5129,N_4112,N_4758);
nand U5130 (N_5130,N_4600,N_4639);
and U5131 (N_5131,N_4959,N_4283);
and U5132 (N_5132,N_4235,N_4142);
nor U5133 (N_5133,N_4854,N_4063);
or U5134 (N_5134,N_4447,N_4916);
nor U5135 (N_5135,N_4595,N_4036);
nand U5136 (N_5136,N_4679,N_4992);
or U5137 (N_5137,N_4474,N_4097);
or U5138 (N_5138,N_4647,N_4310);
nor U5139 (N_5139,N_4820,N_4234);
and U5140 (N_5140,N_4543,N_4351);
or U5141 (N_5141,N_4952,N_4008);
or U5142 (N_5142,N_4811,N_4672);
nor U5143 (N_5143,N_4353,N_4702);
nor U5144 (N_5144,N_4085,N_4105);
nor U5145 (N_5145,N_4212,N_4178);
and U5146 (N_5146,N_4181,N_4497);
xor U5147 (N_5147,N_4099,N_4895);
nand U5148 (N_5148,N_4440,N_4137);
xnor U5149 (N_5149,N_4550,N_4586);
nor U5150 (N_5150,N_4312,N_4297);
and U5151 (N_5151,N_4742,N_4710);
and U5152 (N_5152,N_4014,N_4067);
or U5153 (N_5153,N_4168,N_4214);
or U5154 (N_5154,N_4120,N_4962);
nor U5155 (N_5155,N_4694,N_4606);
xor U5156 (N_5156,N_4675,N_4109);
and U5157 (N_5157,N_4059,N_4761);
or U5158 (N_5158,N_4882,N_4701);
or U5159 (N_5159,N_4028,N_4521);
or U5160 (N_5160,N_4130,N_4429);
or U5161 (N_5161,N_4805,N_4155);
and U5162 (N_5162,N_4043,N_4526);
xnor U5163 (N_5163,N_4492,N_4398);
xnor U5164 (N_5164,N_4000,N_4457);
xnor U5165 (N_5165,N_4637,N_4905);
nand U5166 (N_5166,N_4277,N_4875);
or U5167 (N_5167,N_4402,N_4687);
or U5168 (N_5168,N_4927,N_4809);
xnor U5169 (N_5169,N_4012,N_4334);
and U5170 (N_5170,N_4692,N_4273);
and U5171 (N_5171,N_4625,N_4529);
or U5172 (N_5172,N_4919,N_4049);
or U5173 (N_5173,N_4197,N_4432);
nor U5174 (N_5174,N_4655,N_4065);
xnor U5175 (N_5175,N_4638,N_4685);
nand U5176 (N_5176,N_4923,N_4327);
nor U5177 (N_5177,N_4620,N_4242);
nand U5178 (N_5178,N_4141,N_4229);
or U5179 (N_5179,N_4169,N_4091);
nand U5180 (N_5180,N_4294,N_4355);
and U5181 (N_5181,N_4132,N_4829);
or U5182 (N_5182,N_4582,N_4548);
or U5183 (N_5183,N_4050,N_4914);
or U5184 (N_5184,N_4732,N_4186);
xor U5185 (N_5185,N_4801,N_4707);
xnor U5186 (N_5186,N_4540,N_4549);
and U5187 (N_5187,N_4160,N_4266);
or U5188 (N_5188,N_4330,N_4976);
and U5189 (N_5189,N_4860,N_4004);
and U5190 (N_5190,N_4458,N_4468);
nand U5191 (N_5191,N_4017,N_4779);
nand U5192 (N_5192,N_4979,N_4305);
nand U5193 (N_5193,N_4376,N_4937);
nand U5194 (N_5194,N_4460,N_4487);
nor U5195 (N_5195,N_4715,N_4920);
xor U5196 (N_5196,N_4117,N_4090);
or U5197 (N_5197,N_4400,N_4317);
nor U5198 (N_5198,N_4348,N_4172);
or U5199 (N_5199,N_4369,N_4735);
nand U5200 (N_5200,N_4969,N_4073);
nor U5201 (N_5201,N_4967,N_4578);
and U5202 (N_5202,N_4651,N_4652);
or U5203 (N_5203,N_4157,N_4103);
nor U5204 (N_5204,N_4743,N_4005);
nand U5205 (N_5205,N_4081,N_4680);
nor U5206 (N_5206,N_4048,N_4760);
or U5207 (N_5207,N_4886,N_4557);
nand U5208 (N_5208,N_4552,N_4673);
and U5209 (N_5209,N_4208,N_4819);
nor U5210 (N_5210,N_4339,N_4771);
nand U5211 (N_5211,N_4300,N_4836);
nand U5212 (N_5212,N_4782,N_4590);
and U5213 (N_5213,N_4146,N_4745);
nor U5214 (N_5214,N_4812,N_4009);
nor U5215 (N_5215,N_4532,N_4736);
and U5216 (N_5216,N_4449,N_4561);
or U5217 (N_5217,N_4167,N_4072);
nor U5218 (N_5218,N_4955,N_4839);
and U5219 (N_5219,N_4807,N_4553);
or U5220 (N_5220,N_4721,N_4071);
nand U5221 (N_5221,N_4855,N_4577);
xnor U5222 (N_5222,N_4795,N_4954);
xor U5223 (N_5223,N_4653,N_4313);
or U5224 (N_5224,N_4808,N_4942);
xor U5225 (N_5225,N_4848,N_4986);
nand U5226 (N_5226,N_4716,N_4929);
or U5227 (N_5227,N_4074,N_4027);
and U5228 (N_5228,N_4045,N_4261);
and U5229 (N_5229,N_4255,N_4724);
and U5230 (N_5230,N_4536,N_4108);
or U5231 (N_5231,N_4135,N_4523);
nand U5232 (N_5232,N_4671,N_4211);
and U5233 (N_5233,N_4272,N_4597);
and U5234 (N_5234,N_4040,N_4876);
xnor U5235 (N_5235,N_4165,N_4930);
or U5236 (N_5236,N_4910,N_4426);
and U5237 (N_5237,N_4871,N_4781);
xnor U5238 (N_5238,N_4102,N_4149);
nand U5239 (N_5239,N_4406,N_4901);
nand U5240 (N_5240,N_4451,N_4082);
nor U5241 (N_5241,N_4912,N_4974);
nor U5242 (N_5242,N_4371,N_4281);
nand U5243 (N_5243,N_4057,N_4826);
or U5244 (N_5244,N_4566,N_4213);
nor U5245 (N_5245,N_4650,N_4605);
nand U5246 (N_5246,N_4733,N_4298);
nand U5247 (N_5247,N_4906,N_4517);
nand U5248 (N_5248,N_4316,N_4594);
and U5249 (N_5249,N_4883,N_4070);
and U5250 (N_5250,N_4644,N_4678);
nand U5251 (N_5251,N_4176,N_4897);
and U5252 (N_5252,N_4366,N_4016);
xor U5253 (N_5253,N_4293,N_4238);
and U5254 (N_5254,N_4188,N_4239);
or U5255 (N_5255,N_4342,N_4089);
nor U5256 (N_5256,N_4391,N_4999);
xor U5257 (N_5257,N_4058,N_4174);
nor U5258 (N_5258,N_4194,N_4865);
or U5259 (N_5259,N_4104,N_4343);
or U5260 (N_5260,N_4844,N_4198);
and U5261 (N_5261,N_4280,N_4251);
nand U5262 (N_5262,N_4437,N_4469);
and U5263 (N_5263,N_4508,N_4296);
nor U5264 (N_5264,N_4729,N_4125);
xor U5265 (N_5265,N_4698,N_4029);
nand U5266 (N_5266,N_4887,N_4228);
and U5267 (N_5267,N_4363,N_4061);
xor U5268 (N_5268,N_4480,N_4872);
or U5269 (N_5269,N_4800,N_4470);
xor U5270 (N_5270,N_4409,N_4417);
nand U5271 (N_5271,N_4037,N_4691);
nand U5272 (N_5272,N_4717,N_4659);
xor U5273 (N_5273,N_4434,N_4940);
xnor U5274 (N_5274,N_4356,N_4799);
or U5275 (N_5275,N_4834,N_4325);
nor U5276 (N_5276,N_4627,N_4113);
nand U5277 (N_5277,N_4412,N_4060);
and U5278 (N_5278,N_4265,N_4924);
nand U5279 (N_5279,N_4907,N_4847);
or U5280 (N_5280,N_4730,N_4423);
nor U5281 (N_5281,N_4911,N_4001);
nor U5282 (N_5282,N_4094,N_4815);
nand U5283 (N_5283,N_4555,N_4857);
xnor U5284 (N_5284,N_4709,N_4562);
nand U5285 (N_5285,N_4755,N_4524);
xnor U5286 (N_5286,N_4970,N_4533);
xor U5287 (N_5287,N_4436,N_4128);
nor U5288 (N_5288,N_4495,N_4362);
xor U5289 (N_5289,N_4077,N_4393);
nor U5290 (N_5290,N_4493,N_4151);
xor U5291 (N_5291,N_4175,N_4545);
nor U5292 (N_5292,N_4530,N_4180);
nor U5293 (N_5293,N_4161,N_4479);
or U5294 (N_5294,N_4534,N_4279);
nor U5295 (N_5295,N_4359,N_4943);
nor U5296 (N_5296,N_4051,N_4757);
or U5297 (N_5297,N_4187,N_4777);
xor U5298 (N_5298,N_4780,N_4665);
xnor U5299 (N_5299,N_4686,N_4706);
nand U5300 (N_5300,N_4773,N_4386);
nor U5301 (N_5301,N_4794,N_4722);
or U5302 (N_5302,N_4703,N_4585);
nand U5303 (N_5303,N_4684,N_4998);
or U5304 (N_5304,N_4934,N_4215);
or U5305 (N_5305,N_4642,N_4973);
nor U5306 (N_5306,N_4024,N_4747);
or U5307 (N_5307,N_4282,N_4921);
nand U5308 (N_5308,N_4122,N_4772);
nor U5309 (N_5309,N_4473,N_4139);
or U5310 (N_5310,N_4505,N_4006);
or U5311 (N_5311,N_4471,N_4598);
and U5312 (N_5312,N_4329,N_4226);
nand U5313 (N_5313,N_4568,N_4903);
nand U5314 (N_5314,N_4053,N_4560);
or U5315 (N_5315,N_4250,N_4972);
and U5316 (N_5316,N_4311,N_4333);
or U5317 (N_5317,N_4587,N_4879);
nand U5318 (N_5318,N_4835,N_4643);
nor U5319 (N_5319,N_4038,N_4990);
and U5320 (N_5320,N_4633,N_4240);
nor U5321 (N_5321,N_4945,N_4520);
xnor U5322 (N_5322,N_4516,N_4859);
and U5323 (N_5323,N_4140,N_4424);
xnor U5324 (N_5324,N_4192,N_4588);
nand U5325 (N_5325,N_4491,N_4177);
nand U5326 (N_5326,N_4898,N_4466);
and U5327 (N_5327,N_4258,N_4614);
xnor U5328 (N_5328,N_4950,N_4810);
or U5329 (N_5329,N_4502,N_4853);
xor U5330 (N_5330,N_4900,N_4331);
or U5331 (N_5331,N_4669,N_4041);
xnor U5332 (N_5332,N_4368,N_4858);
xnor U5333 (N_5333,N_4098,N_4607);
or U5334 (N_5334,N_4503,N_4754);
nor U5335 (N_5335,N_4926,N_4866);
and U5336 (N_5336,N_4318,N_4965);
xor U5337 (N_5337,N_4525,N_4749);
xor U5338 (N_5338,N_4890,N_4889);
xnor U5339 (N_5339,N_4891,N_4218);
nand U5340 (N_5340,N_4340,N_4547);
and U5341 (N_5341,N_4971,N_4793);
nor U5342 (N_5342,N_4797,N_4500);
nand U5343 (N_5343,N_4427,N_4851);
xnor U5344 (N_5344,N_4775,N_4792);
nand U5345 (N_5345,N_4740,N_4997);
or U5346 (N_5346,N_4576,N_4392);
and U5347 (N_5347,N_4079,N_4944);
nor U5348 (N_5348,N_4119,N_4013);
or U5349 (N_5349,N_4928,N_4078);
nor U5350 (N_5350,N_4158,N_4189);
xnor U5351 (N_5351,N_4695,N_4475);
nor U5352 (N_5352,N_4015,N_4092);
and U5353 (N_5353,N_4031,N_4843);
or U5354 (N_5354,N_4025,N_4110);
xor U5355 (N_5355,N_4439,N_4828);
xnor U5356 (N_5356,N_4917,N_4224);
xor U5357 (N_5357,N_4615,N_4938);
or U5358 (N_5358,N_4881,N_4287);
and U5359 (N_5359,N_4076,N_4150);
and U5360 (N_5360,N_4260,N_4247);
xnor U5361 (N_5361,N_4304,N_4817);
nand U5362 (N_5362,N_4556,N_4482);
nor U5363 (N_5363,N_4372,N_4636);
nand U5364 (N_5364,N_4245,N_4784);
or U5365 (N_5365,N_4626,N_4720);
nand U5366 (N_5366,N_4465,N_4126);
or U5367 (N_5367,N_4518,N_4870);
nand U5368 (N_5368,N_4217,N_4682);
or U5369 (N_5369,N_4075,N_4677);
nor U5370 (N_5370,N_4768,N_4632);
or U5371 (N_5371,N_4095,N_4039);
xnor U5372 (N_5372,N_4007,N_4115);
nor U5373 (N_5373,N_4207,N_4878);
or U5374 (N_5374,N_4507,N_4496);
xor U5375 (N_5375,N_4199,N_4416);
nor U5376 (N_5376,N_4462,N_4880);
xnor U5377 (N_5377,N_4044,N_4384);
nor U5378 (N_5378,N_4162,N_4405);
xor U5379 (N_5379,N_4542,N_4584);
or U5380 (N_5380,N_4804,N_4592);
and U5381 (N_5381,N_4206,N_4489);
nor U5382 (N_5382,N_4759,N_4727);
or U5383 (N_5383,N_4464,N_4454);
nand U5384 (N_5384,N_4237,N_4445);
nor U5385 (N_5385,N_4551,N_4975);
and U5386 (N_5386,N_4580,N_4646);
and U5387 (N_5387,N_4996,N_4148);
or U5388 (N_5388,N_4763,N_4528);
nor U5389 (N_5389,N_4932,N_4738);
or U5390 (N_5390,N_4184,N_4002);
nand U5391 (N_5391,N_4711,N_4463);
nand U5392 (N_5392,N_4947,N_4752);
nand U5393 (N_5393,N_4667,N_4270);
nand U5394 (N_5394,N_4159,N_4145);
or U5395 (N_5395,N_4621,N_4904);
and U5396 (N_5396,N_4225,N_4668);
nand U5397 (N_5397,N_4751,N_4018);
and U5398 (N_5398,N_4332,N_4499);
nor U5399 (N_5399,N_4370,N_4609);
or U5400 (N_5400,N_4227,N_4259);
nor U5401 (N_5401,N_4964,N_4220);
and U5402 (N_5402,N_4116,N_4345);
nand U5403 (N_5403,N_4593,N_4699);
xnor U5404 (N_5404,N_4814,N_4849);
nand U5405 (N_5405,N_4026,N_4399);
nand U5406 (N_5406,N_4030,N_4842);
nand U5407 (N_5407,N_4309,N_4106);
or U5408 (N_5408,N_4422,N_4068);
xor U5409 (N_5409,N_4506,N_4477);
xnor U5410 (N_5410,N_4052,N_4640);
and U5411 (N_5411,N_4136,N_4510);
and U5412 (N_5412,N_4693,N_4269);
nor U5413 (N_5413,N_4278,N_4664);
xor U5414 (N_5414,N_4725,N_4527);
or U5415 (N_5415,N_4302,N_4705);
or U5416 (N_5416,N_4364,N_4357);
or U5417 (N_5417,N_4988,N_4170);
nand U5418 (N_5418,N_4756,N_4993);
nor U5419 (N_5419,N_4674,N_4753);
and U5420 (N_5420,N_4093,N_4893);
nand U5421 (N_5421,N_4723,N_4490);
and U5422 (N_5422,N_4156,N_4802);
nor U5423 (N_5423,N_4285,N_4991);
or U5424 (N_5424,N_4303,N_4825);
and U5425 (N_5425,N_4344,N_4337);
nand U5426 (N_5426,N_4918,N_4539);
and U5427 (N_5427,N_4166,N_4390);
nand U5428 (N_5428,N_4798,N_4960);
or U5429 (N_5429,N_4948,N_4596);
or U5430 (N_5430,N_4382,N_4154);
nand U5431 (N_5431,N_4623,N_4444);
or U5432 (N_5432,N_4538,N_4573);
nor U5433 (N_5433,N_4734,N_4608);
nor U5434 (N_5434,N_4488,N_4138);
or U5435 (N_5435,N_4728,N_4494);
and U5436 (N_5436,N_4604,N_4837);
and U5437 (N_5437,N_4838,N_4455);
or U5438 (N_5438,N_4514,N_4425);
and U5439 (N_5439,N_4069,N_4223);
or U5440 (N_5440,N_4080,N_4634);
xnor U5441 (N_5441,N_4254,N_4591);
and U5442 (N_5442,N_4739,N_4676);
nand U5443 (N_5443,N_4863,N_4661);
nand U5444 (N_5444,N_4096,N_4011);
nand U5445 (N_5445,N_4448,N_4367);
xor U5446 (N_5446,N_4896,N_4361);
nor U5447 (N_5447,N_4645,N_4478);
or U5448 (N_5448,N_4791,N_4350);
or U5449 (N_5449,N_4246,N_4599);
nand U5450 (N_5450,N_4064,N_4315);
xor U5451 (N_5451,N_4786,N_4381);
nand U5452 (N_5452,N_4284,N_4248);
or U5453 (N_5453,N_4249,N_4243);
nand U5454 (N_5454,N_4485,N_4377);
xor U5455 (N_5455,N_4764,N_4796);
xor U5456 (N_5456,N_4035,N_4289);
or U5457 (N_5457,N_4443,N_4726);
and U5458 (N_5458,N_4513,N_4395);
xor U5459 (N_5459,N_4861,N_4719);
nor U5460 (N_5460,N_4546,N_4319);
and U5461 (N_5461,N_4827,N_4147);
or U5462 (N_5462,N_4788,N_4984);
nand U5463 (N_5463,N_4387,N_4314);
nand U5464 (N_5464,N_4411,N_4762);
xor U5465 (N_5465,N_4143,N_4452);
nand U5466 (N_5466,N_4274,N_4951);
xnor U5467 (N_5467,N_4980,N_4328);
and U5468 (N_5468,N_4054,N_4877);
nor U5469 (N_5469,N_4631,N_4766);
or U5470 (N_5470,N_4385,N_4397);
nor U5471 (N_5471,N_4869,N_4203);
or U5472 (N_5472,N_4394,N_4818);
nand U5473 (N_5473,N_4338,N_4088);
xor U5474 (N_5474,N_4019,N_4958);
nand U5475 (N_5475,N_4570,N_4498);
xnor U5476 (N_5476,N_4100,N_4276);
xor U5477 (N_5477,N_4336,N_4450);
or U5478 (N_5478,N_4769,N_4985);
and U5479 (N_5479,N_4658,N_4697);
and U5480 (N_5480,N_4055,N_4746);
and U5481 (N_5481,N_4114,N_4931);
nor U5482 (N_5482,N_4453,N_4346);
or U5483 (N_5483,N_4121,N_4575);
and U5484 (N_5484,N_4185,N_4894);
or U5485 (N_5485,N_4622,N_4472);
or U5486 (N_5486,N_4341,N_4750);
and U5487 (N_5487,N_4352,N_4558);
and U5488 (N_5488,N_4292,N_4133);
and U5489 (N_5489,N_4892,N_4164);
xnor U5490 (N_5490,N_4442,N_4567);
and U5491 (N_5491,N_4379,N_4205);
xnor U5492 (N_5492,N_4163,N_4864);
xnor U5493 (N_5493,N_4375,N_4295);
nor U5494 (N_5494,N_4195,N_4374);
nor U5495 (N_5495,N_4046,N_4291);
xnor U5496 (N_5496,N_4936,N_4741);
or U5497 (N_5497,N_4583,N_4683);
nand U5498 (N_5498,N_4867,N_4852);
or U5499 (N_5499,N_4420,N_4481);
or U5500 (N_5500,N_4220,N_4645);
or U5501 (N_5501,N_4445,N_4522);
and U5502 (N_5502,N_4998,N_4873);
nor U5503 (N_5503,N_4970,N_4337);
nor U5504 (N_5504,N_4422,N_4221);
or U5505 (N_5505,N_4039,N_4510);
nand U5506 (N_5506,N_4004,N_4407);
or U5507 (N_5507,N_4344,N_4663);
xnor U5508 (N_5508,N_4789,N_4911);
xnor U5509 (N_5509,N_4617,N_4248);
and U5510 (N_5510,N_4005,N_4627);
or U5511 (N_5511,N_4497,N_4633);
nor U5512 (N_5512,N_4794,N_4301);
nand U5513 (N_5513,N_4154,N_4489);
nor U5514 (N_5514,N_4914,N_4383);
nor U5515 (N_5515,N_4585,N_4809);
or U5516 (N_5516,N_4191,N_4955);
xor U5517 (N_5517,N_4010,N_4862);
and U5518 (N_5518,N_4211,N_4031);
or U5519 (N_5519,N_4306,N_4107);
and U5520 (N_5520,N_4866,N_4037);
nand U5521 (N_5521,N_4863,N_4816);
xnor U5522 (N_5522,N_4232,N_4723);
nor U5523 (N_5523,N_4231,N_4773);
nor U5524 (N_5524,N_4207,N_4962);
xor U5525 (N_5525,N_4695,N_4985);
xor U5526 (N_5526,N_4070,N_4860);
xor U5527 (N_5527,N_4177,N_4309);
nand U5528 (N_5528,N_4144,N_4790);
nand U5529 (N_5529,N_4099,N_4270);
or U5530 (N_5530,N_4103,N_4235);
nand U5531 (N_5531,N_4892,N_4156);
xor U5532 (N_5532,N_4352,N_4048);
and U5533 (N_5533,N_4091,N_4064);
and U5534 (N_5534,N_4877,N_4397);
or U5535 (N_5535,N_4456,N_4354);
xor U5536 (N_5536,N_4029,N_4787);
nor U5537 (N_5537,N_4287,N_4190);
nor U5538 (N_5538,N_4585,N_4893);
or U5539 (N_5539,N_4299,N_4681);
and U5540 (N_5540,N_4636,N_4533);
or U5541 (N_5541,N_4132,N_4486);
xnor U5542 (N_5542,N_4434,N_4715);
nand U5543 (N_5543,N_4390,N_4578);
xnor U5544 (N_5544,N_4826,N_4724);
and U5545 (N_5545,N_4553,N_4048);
and U5546 (N_5546,N_4636,N_4383);
and U5547 (N_5547,N_4510,N_4591);
nor U5548 (N_5548,N_4626,N_4541);
xnor U5549 (N_5549,N_4073,N_4003);
nor U5550 (N_5550,N_4128,N_4702);
or U5551 (N_5551,N_4211,N_4894);
nor U5552 (N_5552,N_4104,N_4315);
xor U5553 (N_5553,N_4589,N_4092);
nor U5554 (N_5554,N_4076,N_4605);
and U5555 (N_5555,N_4283,N_4382);
and U5556 (N_5556,N_4958,N_4467);
xor U5557 (N_5557,N_4772,N_4753);
nor U5558 (N_5558,N_4495,N_4441);
and U5559 (N_5559,N_4222,N_4897);
xor U5560 (N_5560,N_4983,N_4914);
and U5561 (N_5561,N_4324,N_4209);
or U5562 (N_5562,N_4870,N_4777);
xnor U5563 (N_5563,N_4824,N_4334);
or U5564 (N_5564,N_4883,N_4642);
and U5565 (N_5565,N_4129,N_4403);
nor U5566 (N_5566,N_4550,N_4415);
xor U5567 (N_5567,N_4560,N_4813);
nor U5568 (N_5568,N_4122,N_4538);
nor U5569 (N_5569,N_4852,N_4642);
nand U5570 (N_5570,N_4074,N_4333);
xor U5571 (N_5571,N_4765,N_4245);
and U5572 (N_5572,N_4810,N_4057);
xor U5573 (N_5573,N_4469,N_4297);
and U5574 (N_5574,N_4158,N_4173);
nor U5575 (N_5575,N_4275,N_4210);
xor U5576 (N_5576,N_4839,N_4431);
xnor U5577 (N_5577,N_4659,N_4620);
nor U5578 (N_5578,N_4265,N_4179);
xor U5579 (N_5579,N_4439,N_4435);
nor U5580 (N_5580,N_4299,N_4310);
and U5581 (N_5581,N_4505,N_4117);
and U5582 (N_5582,N_4296,N_4848);
or U5583 (N_5583,N_4247,N_4411);
or U5584 (N_5584,N_4463,N_4548);
nor U5585 (N_5585,N_4021,N_4950);
nand U5586 (N_5586,N_4849,N_4390);
xnor U5587 (N_5587,N_4023,N_4404);
nand U5588 (N_5588,N_4630,N_4137);
and U5589 (N_5589,N_4701,N_4919);
xnor U5590 (N_5590,N_4326,N_4982);
and U5591 (N_5591,N_4826,N_4937);
and U5592 (N_5592,N_4989,N_4958);
or U5593 (N_5593,N_4703,N_4245);
or U5594 (N_5594,N_4173,N_4189);
and U5595 (N_5595,N_4641,N_4134);
or U5596 (N_5596,N_4059,N_4024);
or U5597 (N_5597,N_4113,N_4107);
or U5598 (N_5598,N_4491,N_4778);
nand U5599 (N_5599,N_4488,N_4988);
xnor U5600 (N_5600,N_4208,N_4573);
nor U5601 (N_5601,N_4040,N_4597);
or U5602 (N_5602,N_4517,N_4985);
nand U5603 (N_5603,N_4123,N_4862);
xnor U5604 (N_5604,N_4912,N_4939);
and U5605 (N_5605,N_4079,N_4480);
nor U5606 (N_5606,N_4191,N_4761);
xnor U5607 (N_5607,N_4491,N_4550);
nand U5608 (N_5608,N_4188,N_4271);
or U5609 (N_5609,N_4989,N_4525);
or U5610 (N_5610,N_4407,N_4441);
or U5611 (N_5611,N_4813,N_4931);
nand U5612 (N_5612,N_4480,N_4978);
xor U5613 (N_5613,N_4096,N_4205);
nand U5614 (N_5614,N_4036,N_4964);
or U5615 (N_5615,N_4196,N_4868);
nor U5616 (N_5616,N_4208,N_4529);
nand U5617 (N_5617,N_4565,N_4431);
xor U5618 (N_5618,N_4465,N_4210);
or U5619 (N_5619,N_4487,N_4474);
or U5620 (N_5620,N_4956,N_4636);
or U5621 (N_5621,N_4494,N_4770);
nand U5622 (N_5622,N_4105,N_4447);
or U5623 (N_5623,N_4649,N_4697);
nor U5624 (N_5624,N_4501,N_4547);
xor U5625 (N_5625,N_4643,N_4648);
or U5626 (N_5626,N_4981,N_4484);
nand U5627 (N_5627,N_4654,N_4498);
and U5628 (N_5628,N_4379,N_4892);
xnor U5629 (N_5629,N_4562,N_4522);
and U5630 (N_5630,N_4698,N_4575);
nor U5631 (N_5631,N_4283,N_4446);
and U5632 (N_5632,N_4589,N_4991);
xnor U5633 (N_5633,N_4652,N_4139);
nand U5634 (N_5634,N_4494,N_4852);
nor U5635 (N_5635,N_4990,N_4594);
and U5636 (N_5636,N_4181,N_4923);
and U5637 (N_5637,N_4193,N_4444);
nand U5638 (N_5638,N_4711,N_4975);
xnor U5639 (N_5639,N_4777,N_4540);
and U5640 (N_5640,N_4591,N_4891);
xor U5641 (N_5641,N_4292,N_4833);
nor U5642 (N_5642,N_4104,N_4310);
or U5643 (N_5643,N_4519,N_4783);
and U5644 (N_5644,N_4967,N_4891);
or U5645 (N_5645,N_4133,N_4409);
nand U5646 (N_5646,N_4352,N_4880);
xor U5647 (N_5647,N_4691,N_4114);
nor U5648 (N_5648,N_4066,N_4349);
xnor U5649 (N_5649,N_4893,N_4073);
or U5650 (N_5650,N_4287,N_4252);
nand U5651 (N_5651,N_4394,N_4967);
xor U5652 (N_5652,N_4229,N_4824);
and U5653 (N_5653,N_4009,N_4089);
nand U5654 (N_5654,N_4410,N_4023);
xor U5655 (N_5655,N_4194,N_4880);
xnor U5656 (N_5656,N_4142,N_4132);
nand U5657 (N_5657,N_4377,N_4064);
nor U5658 (N_5658,N_4238,N_4721);
or U5659 (N_5659,N_4177,N_4885);
xnor U5660 (N_5660,N_4690,N_4562);
and U5661 (N_5661,N_4412,N_4181);
xnor U5662 (N_5662,N_4120,N_4739);
nand U5663 (N_5663,N_4949,N_4712);
nor U5664 (N_5664,N_4210,N_4678);
and U5665 (N_5665,N_4282,N_4049);
xor U5666 (N_5666,N_4002,N_4605);
nand U5667 (N_5667,N_4755,N_4003);
or U5668 (N_5668,N_4003,N_4262);
nor U5669 (N_5669,N_4494,N_4269);
xor U5670 (N_5670,N_4847,N_4062);
nor U5671 (N_5671,N_4086,N_4746);
or U5672 (N_5672,N_4573,N_4703);
nand U5673 (N_5673,N_4562,N_4644);
nor U5674 (N_5674,N_4908,N_4308);
or U5675 (N_5675,N_4408,N_4186);
xor U5676 (N_5676,N_4316,N_4562);
and U5677 (N_5677,N_4537,N_4891);
xnor U5678 (N_5678,N_4035,N_4222);
xnor U5679 (N_5679,N_4083,N_4578);
nor U5680 (N_5680,N_4506,N_4213);
xnor U5681 (N_5681,N_4448,N_4270);
or U5682 (N_5682,N_4740,N_4147);
nor U5683 (N_5683,N_4570,N_4138);
and U5684 (N_5684,N_4581,N_4831);
xor U5685 (N_5685,N_4757,N_4024);
or U5686 (N_5686,N_4390,N_4546);
xnor U5687 (N_5687,N_4279,N_4077);
nor U5688 (N_5688,N_4403,N_4743);
xnor U5689 (N_5689,N_4665,N_4836);
nand U5690 (N_5690,N_4462,N_4291);
or U5691 (N_5691,N_4079,N_4725);
xnor U5692 (N_5692,N_4699,N_4407);
nand U5693 (N_5693,N_4244,N_4998);
nor U5694 (N_5694,N_4468,N_4344);
xor U5695 (N_5695,N_4314,N_4042);
nand U5696 (N_5696,N_4424,N_4326);
and U5697 (N_5697,N_4232,N_4579);
xor U5698 (N_5698,N_4770,N_4885);
nor U5699 (N_5699,N_4379,N_4439);
nor U5700 (N_5700,N_4782,N_4965);
and U5701 (N_5701,N_4622,N_4816);
nand U5702 (N_5702,N_4556,N_4602);
and U5703 (N_5703,N_4276,N_4486);
nor U5704 (N_5704,N_4735,N_4840);
xor U5705 (N_5705,N_4429,N_4452);
nand U5706 (N_5706,N_4696,N_4308);
and U5707 (N_5707,N_4546,N_4554);
xnor U5708 (N_5708,N_4574,N_4107);
xnor U5709 (N_5709,N_4304,N_4505);
or U5710 (N_5710,N_4345,N_4594);
and U5711 (N_5711,N_4567,N_4639);
or U5712 (N_5712,N_4193,N_4253);
xor U5713 (N_5713,N_4439,N_4821);
nor U5714 (N_5714,N_4417,N_4957);
xnor U5715 (N_5715,N_4887,N_4812);
nor U5716 (N_5716,N_4008,N_4767);
nand U5717 (N_5717,N_4015,N_4507);
xor U5718 (N_5718,N_4760,N_4553);
or U5719 (N_5719,N_4719,N_4592);
nor U5720 (N_5720,N_4637,N_4370);
xor U5721 (N_5721,N_4004,N_4631);
xor U5722 (N_5722,N_4847,N_4299);
and U5723 (N_5723,N_4504,N_4008);
and U5724 (N_5724,N_4814,N_4799);
or U5725 (N_5725,N_4915,N_4374);
xor U5726 (N_5726,N_4346,N_4255);
nor U5727 (N_5727,N_4722,N_4678);
nand U5728 (N_5728,N_4325,N_4593);
and U5729 (N_5729,N_4623,N_4197);
nor U5730 (N_5730,N_4126,N_4923);
or U5731 (N_5731,N_4458,N_4325);
nor U5732 (N_5732,N_4227,N_4841);
and U5733 (N_5733,N_4791,N_4424);
or U5734 (N_5734,N_4825,N_4008);
or U5735 (N_5735,N_4582,N_4173);
nand U5736 (N_5736,N_4211,N_4364);
or U5737 (N_5737,N_4312,N_4802);
nand U5738 (N_5738,N_4529,N_4695);
nand U5739 (N_5739,N_4495,N_4112);
nor U5740 (N_5740,N_4093,N_4791);
or U5741 (N_5741,N_4102,N_4909);
and U5742 (N_5742,N_4673,N_4737);
or U5743 (N_5743,N_4193,N_4657);
or U5744 (N_5744,N_4786,N_4567);
nand U5745 (N_5745,N_4840,N_4141);
nor U5746 (N_5746,N_4376,N_4700);
and U5747 (N_5747,N_4806,N_4122);
and U5748 (N_5748,N_4792,N_4253);
xor U5749 (N_5749,N_4988,N_4400);
or U5750 (N_5750,N_4597,N_4972);
xor U5751 (N_5751,N_4381,N_4299);
nand U5752 (N_5752,N_4719,N_4965);
nand U5753 (N_5753,N_4874,N_4778);
and U5754 (N_5754,N_4742,N_4557);
xnor U5755 (N_5755,N_4041,N_4643);
and U5756 (N_5756,N_4870,N_4509);
or U5757 (N_5757,N_4002,N_4412);
nand U5758 (N_5758,N_4502,N_4160);
and U5759 (N_5759,N_4015,N_4320);
or U5760 (N_5760,N_4835,N_4713);
xor U5761 (N_5761,N_4109,N_4749);
nor U5762 (N_5762,N_4756,N_4185);
or U5763 (N_5763,N_4378,N_4348);
and U5764 (N_5764,N_4161,N_4418);
or U5765 (N_5765,N_4141,N_4725);
nand U5766 (N_5766,N_4535,N_4356);
or U5767 (N_5767,N_4629,N_4664);
nand U5768 (N_5768,N_4944,N_4542);
or U5769 (N_5769,N_4009,N_4595);
nor U5770 (N_5770,N_4732,N_4599);
xor U5771 (N_5771,N_4532,N_4672);
and U5772 (N_5772,N_4469,N_4744);
nor U5773 (N_5773,N_4334,N_4474);
nand U5774 (N_5774,N_4738,N_4172);
nor U5775 (N_5775,N_4727,N_4000);
nor U5776 (N_5776,N_4463,N_4718);
xor U5777 (N_5777,N_4037,N_4486);
and U5778 (N_5778,N_4721,N_4680);
and U5779 (N_5779,N_4524,N_4740);
xor U5780 (N_5780,N_4856,N_4897);
or U5781 (N_5781,N_4413,N_4305);
or U5782 (N_5782,N_4125,N_4630);
nand U5783 (N_5783,N_4275,N_4983);
or U5784 (N_5784,N_4512,N_4005);
nand U5785 (N_5785,N_4889,N_4970);
nand U5786 (N_5786,N_4862,N_4014);
or U5787 (N_5787,N_4822,N_4842);
and U5788 (N_5788,N_4621,N_4594);
nor U5789 (N_5789,N_4792,N_4330);
xor U5790 (N_5790,N_4422,N_4605);
xnor U5791 (N_5791,N_4262,N_4949);
and U5792 (N_5792,N_4601,N_4758);
nand U5793 (N_5793,N_4087,N_4245);
xor U5794 (N_5794,N_4646,N_4175);
nor U5795 (N_5795,N_4016,N_4918);
nor U5796 (N_5796,N_4400,N_4554);
or U5797 (N_5797,N_4964,N_4195);
nand U5798 (N_5798,N_4636,N_4300);
or U5799 (N_5799,N_4699,N_4803);
and U5800 (N_5800,N_4132,N_4291);
nor U5801 (N_5801,N_4507,N_4131);
xnor U5802 (N_5802,N_4134,N_4797);
nor U5803 (N_5803,N_4320,N_4490);
or U5804 (N_5804,N_4080,N_4292);
and U5805 (N_5805,N_4622,N_4793);
nand U5806 (N_5806,N_4103,N_4516);
or U5807 (N_5807,N_4323,N_4823);
nor U5808 (N_5808,N_4677,N_4706);
nor U5809 (N_5809,N_4537,N_4771);
nand U5810 (N_5810,N_4102,N_4105);
or U5811 (N_5811,N_4009,N_4885);
nor U5812 (N_5812,N_4552,N_4782);
nand U5813 (N_5813,N_4591,N_4540);
xor U5814 (N_5814,N_4697,N_4864);
or U5815 (N_5815,N_4119,N_4091);
and U5816 (N_5816,N_4113,N_4246);
xor U5817 (N_5817,N_4256,N_4351);
or U5818 (N_5818,N_4010,N_4129);
nor U5819 (N_5819,N_4068,N_4592);
nand U5820 (N_5820,N_4463,N_4100);
and U5821 (N_5821,N_4373,N_4206);
and U5822 (N_5822,N_4104,N_4902);
nor U5823 (N_5823,N_4325,N_4485);
xor U5824 (N_5824,N_4052,N_4943);
or U5825 (N_5825,N_4363,N_4131);
and U5826 (N_5826,N_4652,N_4870);
nand U5827 (N_5827,N_4523,N_4750);
nand U5828 (N_5828,N_4892,N_4339);
or U5829 (N_5829,N_4798,N_4156);
xnor U5830 (N_5830,N_4206,N_4951);
and U5831 (N_5831,N_4982,N_4070);
xor U5832 (N_5832,N_4022,N_4991);
nor U5833 (N_5833,N_4517,N_4632);
or U5834 (N_5834,N_4706,N_4642);
nand U5835 (N_5835,N_4726,N_4610);
and U5836 (N_5836,N_4580,N_4271);
and U5837 (N_5837,N_4092,N_4776);
xnor U5838 (N_5838,N_4881,N_4705);
or U5839 (N_5839,N_4230,N_4113);
and U5840 (N_5840,N_4273,N_4716);
and U5841 (N_5841,N_4794,N_4400);
nor U5842 (N_5842,N_4835,N_4878);
xnor U5843 (N_5843,N_4930,N_4764);
nor U5844 (N_5844,N_4956,N_4317);
and U5845 (N_5845,N_4037,N_4821);
and U5846 (N_5846,N_4582,N_4149);
nor U5847 (N_5847,N_4263,N_4411);
nor U5848 (N_5848,N_4987,N_4640);
nor U5849 (N_5849,N_4514,N_4421);
xor U5850 (N_5850,N_4782,N_4538);
and U5851 (N_5851,N_4381,N_4594);
nor U5852 (N_5852,N_4183,N_4933);
nor U5853 (N_5853,N_4345,N_4869);
xor U5854 (N_5854,N_4669,N_4093);
xnor U5855 (N_5855,N_4861,N_4490);
nor U5856 (N_5856,N_4957,N_4473);
or U5857 (N_5857,N_4098,N_4639);
nand U5858 (N_5858,N_4687,N_4344);
nor U5859 (N_5859,N_4086,N_4768);
xor U5860 (N_5860,N_4694,N_4789);
or U5861 (N_5861,N_4540,N_4453);
and U5862 (N_5862,N_4035,N_4296);
and U5863 (N_5863,N_4830,N_4794);
and U5864 (N_5864,N_4369,N_4764);
xnor U5865 (N_5865,N_4255,N_4584);
or U5866 (N_5866,N_4669,N_4934);
nand U5867 (N_5867,N_4814,N_4704);
nor U5868 (N_5868,N_4144,N_4599);
xnor U5869 (N_5869,N_4494,N_4870);
nor U5870 (N_5870,N_4055,N_4661);
and U5871 (N_5871,N_4941,N_4893);
and U5872 (N_5872,N_4713,N_4321);
nand U5873 (N_5873,N_4314,N_4286);
and U5874 (N_5874,N_4941,N_4949);
xor U5875 (N_5875,N_4039,N_4760);
nor U5876 (N_5876,N_4176,N_4096);
nor U5877 (N_5877,N_4426,N_4404);
nand U5878 (N_5878,N_4222,N_4577);
nand U5879 (N_5879,N_4577,N_4401);
nor U5880 (N_5880,N_4324,N_4750);
nand U5881 (N_5881,N_4289,N_4783);
or U5882 (N_5882,N_4728,N_4991);
nand U5883 (N_5883,N_4146,N_4134);
xnor U5884 (N_5884,N_4935,N_4992);
or U5885 (N_5885,N_4382,N_4895);
or U5886 (N_5886,N_4587,N_4591);
nor U5887 (N_5887,N_4624,N_4354);
nor U5888 (N_5888,N_4455,N_4830);
nand U5889 (N_5889,N_4403,N_4588);
and U5890 (N_5890,N_4922,N_4892);
nor U5891 (N_5891,N_4060,N_4345);
nor U5892 (N_5892,N_4573,N_4942);
nor U5893 (N_5893,N_4312,N_4286);
or U5894 (N_5894,N_4568,N_4097);
or U5895 (N_5895,N_4697,N_4462);
or U5896 (N_5896,N_4222,N_4180);
nor U5897 (N_5897,N_4932,N_4492);
and U5898 (N_5898,N_4551,N_4304);
xor U5899 (N_5899,N_4983,N_4472);
xnor U5900 (N_5900,N_4468,N_4356);
xnor U5901 (N_5901,N_4781,N_4233);
nand U5902 (N_5902,N_4844,N_4089);
xor U5903 (N_5903,N_4207,N_4533);
and U5904 (N_5904,N_4092,N_4456);
nand U5905 (N_5905,N_4450,N_4184);
nand U5906 (N_5906,N_4259,N_4343);
or U5907 (N_5907,N_4093,N_4165);
nand U5908 (N_5908,N_4504,N_4309);
or U5909 (N_5909,N_4530,N_4606);
xor U5910 (N_5910,N_4311,N_4462);
nor U5911 (N_5911,N_4125,N_4668);
nand U5912 (N_5912,N_4542,N_4120);
nand U5913 (N_5913,N_4337,N_4526);
nand U5914 (N_5914,N_4889,N_4102);
nand U5915 (N_5915,N_4612,N_4167);
or U5916 (N_5916,N_4520,N_4982);
nor U5917 (N_5917,N_4707,N_4683);
and U5918 (N_5918,N_4071,N_4858);
nand U5919 (N_5919,N_4617,N_4687);
nor U5920 (N_5920,N_4749,N_4061);
or U5921 (N_5921,N_4742,N_4832);
nor U5922 (N_5922,N_4442,N_4983);
xnor U5923 (N_5923,N_4426,N_4051);
xor U5924 (N_5924,N_4046,N_4339);
nor U5925 (N_5925,N_4207,N_4338);
nand U5926 (N_5926,N_4218,N_4249);
xor U5927 (N_5927,N_4706,N_4232);
and U5928 (N_5928,N_4386,N_4809);
or U5929 (N_5929,N_4189,N_4267);
and U5930 (N_5930,N_4468,N_4557);
nand U5931 (N_5931,N_4954,N_4162);
nor U5932 (N_5932,N_4256,N_4248);
or U5933 (N_5933,N_4433,N_4704);
and U5934 (N_5934,N_4942,N_4642);
or U5935 (N_5935,N_4087,N_4095);
or U5936 (N_5936,N_4393,N_4663);
or U5937 (N_5937,N_4030,N_4910);
and U5938 (N_5938,N_4944,N_4717);
nor U5939 (N_5939,N_4579,N_4063);
nand U5940 (N_5940,N_4374,N_4082);
nand U5941 (N_5941,N_4490,N_4112);
or U5942 (N_5942,N_4036,N_4597);
nand U5943 (N_5943,N_4996,N_4178);
xnor U5944 (N_5944,N_4283,N_4873);
nand U5945 (N_5945,N_4237,N_4761);
xor U5946 (N_5946,N_4656,N_4264);
xnor U5947 (N_5947,N_4082,N_4691);
or U5948 (N_5948,N_4535,N_4904);
xnor U5949 (N_5949,N_4693,N_4403);
nor U5950 (N_5950,N_4226,N_4334);
or U5951 (N_5951,N_4431,N_4426);
xor U5952 (N_5952,N_4925,N_4495);
nor U5953 (N_5953,N_4705,N_4976);
nor U5954 (N_5954,N_4660,N_4987);
nor U5955 (N_5955,N_4225,N_4050);
nor U5956 (N_5956,N_4897,N_4347);
and U5957 (N_5957,N_4815,N_4048);
xnor U5958 (N_5958,N_4975,N_4330);
and U5959 (N_5959,N_4588,N_4729);
and U5960 (N_5960,N_4075,N_4086);
xor U5961 (N_5961,N_4693,N_4592);
or U5962 (N_5962,N_4688,N_4501);
or U5963 (N_5963,N_4300,N_4675);
nand U5964 (N_5964,N_4698,N_4996);
and U5965 (N_5965,N_4607,N_4977);
or U5966 (N_5966,N_4145,N_4972);
xnor U5967 (N_5967,N_4939,N_4547);
nand U5968 (N_5968,N_4391,N_4094);
or U5969 (N_5969,N_4938,N_4973);
nand U5970 (N_5970,N_4395,N_4938);
and U5971 (N_5971,N_4337,N_4371);
nand U5972 (N_5972,N_4684,N_4345);
or U5973 (N_5973,N_4899,N_4633);
nand U5974 (N_5974,N_4607,N_4512);
nand U5975 (N_5975,N_4958,N_4911);
xnor U5976 (N_5976,N_4140,N_4861);
or U5977 (N_5977,N_4345,N_4399);
xnor U5978 (N_5978,N_4099,N_4878);
nand U5979 (N_5979,N_4286,N_4340);
nand U5980 (N_5980,N_4359,N_4961);
xnor U5981 (N_5981,N_4068,N_4766);
or U5982 (N_5982,N_4433,N_4150);
xnor U5983 (N_5983,N_4536,N_4476);
xnor U5984 (N_5984,N_4903,N_4391);
and U5985 (N_5985,N_4287,N_4221);
and U5986 (N_5986,N_4527,N_4018);
nand U5987 (N_5987,N_4767,N_4210);
and U5988 (N_5988,N_4576,N_4568);
and U5989 (N_5989,N_4544,N_4233);
xnor U5990 (N_5990,N_4425,N_4986);
nand U5991 (N_5991,N_4039,N_4540);
nor U5992 (N_5992,N_4417,N_4472);
xnor U5993 (N_5993,N_4243,N_4011);
xor U5994 (N_5994,N_4563,N_4417);
nand U5995 (N_5995,N_4964,N_4782);
or U5996 (N_5996,N_4593,N_4944);
nand U5997 (N_5997,N_4104,N_4991);
xnor U5998 (N_5998,N_4086,N_4121);
or U5999 (N_5999,N_4504,N_4546);
or U6000 (N_6000,N_5419,N_5213);
nor U6001 (N_6001,N_5851,N_5017);
nand U6002 (N_6002,N_5471,N_5308);
nor U6003 (N_6003,N_5075,N_5840);
xor U6004 (N_6004,N_5722,N_5614);
and U6005 (N_6005,N_5378,N_5904);
xnor U6006 (N_6006,N_5374,N_5372);
nand U6007 (N_6007,N_5117,N_5223);
or U6008 (N_6008,N_5058,N_5038);
nand U6009 (N_6009,N_5777,N_5275);
nand U6010 (N_6010,N_5617,N_5499);
and U6011 (N_6011,N_5476,N_5636);
xnor U6012 (N_6012,N_5850,N_5100);
and U6013 (N_6013,N_5911,N_5009);
xor U6014 (N_6014,N_5122,N_5628);
xnor U6015 (N_6015,N_5907,N_5989);
or U6016 (N_6016,N_5504,N_5229);
and U6017 (N_6017,N_5800,N_5875);
xor U6018 (N_6018,N_5257,N_5558);
xnor U6019 (N_6019,N_5666,N_5055);
nor U6020 (N_6020,N_5649,N_5693);
or U6021 (N_6021,N_5979,N_5268);
and U6022 (N_6022,N_5940,N_5891);
or U6023 (N_6023,N_5852,N_5143);
nand U6024 (N_6024,N_5113,N_5067);
and U6025 (N_6025,N_5166,N_5252);
nor U6026 (N_6026,N_5464,N_5365);
and U6027 (N_6027,N_5924,N_5262);
and U6028 (N_6028,N_5084,N_5239);
nor U6029 (N_6029,N_5236,N_5848);
xor U6030 (N_6030,N_5659,N_5463);
or U6031 (N_6031,N_5644,N_5887);
nand U6032 (N_6032,N_5266,N_5221);
or U6033 (N_6033,N_5358,N_5178);
xnor U6034 (N_6034,N_5235,N_5453);
and U6035 (N_6035,N_5844,N_5602);
nor U6036 (N_6036,N_5623,N_5783);
and U6037 (N_6037,N_5707,N_5838);
nand U6038 (N_6038,N_5658,N_5801);
nand U6039 (N_6039,N_5396,N_5615);
and U6040 (N_6040,N_5879,N_5081);
nor U6041 (N_6041,N_5402,N_5789);
and U6042 (N_6042,N_5509,N_5151);
nand U6043 (N_6043,N_5170,N_5949);
xnor U6044 (N_6044,N_5926,N_5206);
xnor U6045 (N_6045,N_5336,N_5026);
or U6046 (N_6046,N_5281,N_5973);
nor U6047 (N_6047,N_5467,N_5642);
nor U6048 (N_6048,N_5123,N_5534);
nor U6049 (N_6049,N_5836,N_5042);
xor U6050 (N_6050,N_5885,N_5234);
xnor U6051 (N_6051,N_5595,N_5005);
nand U6052 (N_6052,N_5002,N_5457);
or U6053 (N_6053,N_5124,N_5757);
nand U6054 (N_6054,N_5695,N_5580);
xor U6055 (N_6055,N_5568,N_5766);
xnor U6056 (N_6056,N_5125,N_5134);
or U6057 (N_6057,N_5047,N_5027);
or U6058 (N_6058,N_5812,N_5790);
and U6059 (N_6059,N_5043,N_5622);
xor U6060 (N_6060,N_5974,N_5962);
nand U6061 (N_6061,N_5461,N_5512);
and U6062 (N_6062,N_5046,N_5715);
xor U6063 (N_6063,N_5380,N_5231);
or U6064 (N_6064,N_5684,N_5128);
nand U6065 (N_6065,N_5746,N_5906);
and U6066 (N_6066,N_5525,N_5687);
xnor U6067 (N_6067,N_5408,N_5846);
or U6068 (N_6068,N_5246,N_5630);
and U6069 (N_6069,N_5720,N_5604);
nand U6070 (N_6070,N_5390,N_5277);
and U6071 (N_6071,N_5218,N_5621);
nor U6072 (N_6072,N_5954,N_5528);
xnor U6073 (N_6073,N_5352,N_5116);
xnor U6074 (N_6074,N_5028,N_5226);
xnor U6075 (N_6075,N_5379,N_5893);
xnor U6076 (N_6076,N_5347,N_5708);
xor U6077 (N_6077,N_5016,N_5322);
or U6078 (N_6078,N_5425,N_5514);
or U6079 (N_6079,N_5288,N_5925);
or U6080 (N_6080,N_5943,N_5792);
xor U6081 (N_6081,N_5176,N_5824);
and U6082 (N_6082,N_5340,N_5173);
nor U6083 (N_6083,N_5329,N_5874);
nor U6084 (N_6084,N_5227,N_5552);
nor U6085 (N_6085,N_5302,N_5270);
nor U6086 (N_6086,N_5803,N_5039);
or U6087 (N_6087,N_5169,N_5983);
or U6088 (N_6088,N_5353,N_5489);
xnor U6089 (N_6089,N_5426,N_5035);
xnor U6090 (N_6090,N_5115,N_5423);
nor U6091 (N_6091,N_5496,N_5758);
xnor U6092 (N_6092,N_5465,N_5019);
nor U6093 (N_6093,N_5383,N_5245);
xnor U6094 (N_6094,N_5008,N_5003);
nand U6095 (N_6095,N_5742,N_5348);
nor U6096 (N_6096,N_5669,N_5418);
nand U6097 (N_6097,N_5110,N_5401);
and U6098 (N_6098,N_5267,N_5936);
and U6099 (N_6099,N_5272,N_5431);
xor U6100 (N_6100,N_5540,N_5806);
xor U6101 (N_6101,N_5572,N_5769);
nand U6102 (N_6102,N_5505,N_5053);
and U6103 (N_6103,N_5247,N_5705);
nor U6104 (N_6104,N_5845,N_5085);
nor U6105 (N_6105,N_5611,N_5204);
or U6106 (N_6106,N_5560,N_5459);
or U6107 (N_6107,N_5037,N_5564);
nand U6108 (N_6108,N_5620,N_5307);
and U6109 (N_6109,N_5212,N_5886);
xnor U6110 (N_6110,N_5819,N_5503);
xnor U6111 (N_6111,N_5698,N_5590);
and U6112 (N_6112,N_5316,N_5146);
nor U6113 (N_6113,N_5474,N_5955);
nand U6114 (N_6114,N_5843,N_5916);
or U6115 (N_6115,N_5051,N_5538);
xor U6116 (N_6116,N_5969,N_5452);
xor U6117 (N_6117,N_5325,N_5424);
nand U6118 (N_6118,N_5385,N_5565);
nor U6119 (N_6119,N_5784,N_5036);
xor U6120 (N_6120,N_5119,N_5738);
or U6121 (N_6121,N_5144,N_5205);
or U6122 (N_6122,N_5967,N_5873);
or U6123 (N_6123,N_5631,N_5980);
and U6124 (N_6124,N_5359,N_5948);
or U6125 (N_6125,N_5902,N_5935);
nand U6126 (N_6126,N_5567,N_5716);
nand U6127 (N_6127,N_5177,N_5068);
or U6128 (N_6128,N_5287,N_5928);
or U6129 (N_6129,N_5683,N_5090);
nor U6130 (N_6130,N_5208,N_5473);
nand U6131 (N_6131,N_5972,N_5183);
nor U6132 (N_6132,N_5121,N_5888);
or U6133 (N_6133,N_5711,N_5289);
nor U6134 (N_6134,N_5398,N_5368);
xor U6135 (N_6135,N_5399,N_5938);
nor U6136 (N_6136,N_5071,N_5482);
nor U6137 (N_6137,N_5070,N_5576);
xnor U6138 (N_6138,N_5545,N_5317);
nor U6139 (N_6139,N_5571,N_5515);
and U6140 (N_6140,N_5010,N_5826);
nand U6141 (N_6141,N_5569,N_5494);
nor U6142 (N_6142,N_5714,N_5394);
or U6143 (N_6143,N_5422,N_5781);
or U6144 (N_6144,N_5518,N_5646);
and U6145 (N_6145,N_5349,N_5686);
nor U6146 (N_6146,N_5248,N_5430);
nor U6147 (N_6147,N_5500,N_5153);
or U6148 (N_6148,N_5581,N_5040);
nor U6149 (N_6149,N_5921,N_5673);
xor U6150 (N_6150,N_5855,N_5914);
xor U6151 (N_6151,N_5295,N_5409);
nor U6152 (N_6152,N_5727,N_5250);
or U6153 (N_6153,N_5154,N_5472);
xnor U6154 (N_6154,N_5296,N_5030);
and U6155 (N_6155,N_5158,N_5098);
or U6156 (N_6156,N_5999,N_5774);
xor U6157 (N_6157,N_5355,N_5253);
nand U6158 (N_6158,N_5920,N_5148);
xor U6159 (N_6159,N_5061,N_5141);
nand U6160 (N_6160,N_5201,N_5961);
xor U6161 (N_6161,N_5913,N_5458);
or U6162 (N_6162,N_5324,N_5435);
xor U6163 (N_6163,N_5701,N_5563);
and U6164 (N_6164,N_5788,N_5662);
or U6165 (N_6165,N_5754,N_5388);
xor U6166 (N_6166,N_5413,N_5910);
and U6167 (N_6167,N_5444,N_5917);
xor U6168 (N_6168,N_5432,N_5326);
or U6169 (N_6169,N_5450,N_5335);
xnor U6170 (N_6170,N_5041,N_5541);
nand U6171 (N_6171,N_5439,N_5650);
or U6172 (N_6172,N_5403,N_5895);
xnor U6173 (N_6173,N_5543,N_5735);
nor U6174 (N_6174,N_5607,N_5438);
nor U6175 (N_6175,N_5069,N_5164);
or U6176 (N_6176,N_5127,N_5510);
or U6177 (N_6177,N_5995,N_5020);
nand U6178 (N_6178,N_5680,N_5606);
and U6179 (N_6179,N_5209,N_5837);
nor U6180 (N_6180,N_5918,N_5480);
or U6181 (N_6181,N_5729,N_5798);
or U6182 (N_6182,N_5670,N_5958);
nor U6183 (N_6183,N_5062,N_5537);
and U6184 (N_6184,N_5187,N_5185);
and U6185 (N_6185,N_5933,N_5109);
xnor U6186 (N_6186,N_5282,N_5199);
or U6187 (N_6187,N_5136,N_5618);
or U6188 (N_6188,N_5884,N_5878);
nor U6189 (N_6189,N_5997,N_5544);
xor U6190 (N_6190,N_5807,N_5842);
and U6191 (N_6191,N_5978,N_5276);
and U6192 (N_6192,N_5006,N_5702);
and U6193 (N_6193,N_5321,N_5782);
nand U6194 (N_6194,N_5147,N_5330);
nor U6195 (N_6195,N_5584,N_5072);
or U6196 (N_6196,N_5377,N_5951);
xor U6197 (N_6197,N_5853,N_5101);
or U6198 (N_6198,N_5106,N_5114);
xor U6199 (N_6199,N_5696,N_5832);
nor U6200 (N_6200,N_5883,N_5214);
xor U6201 (N_6201,N_5271,N_5896);
and U6202 (N_6202,N_5847,N_5486);
or U6203 (N_6203,N_5033,N_5478);
or U6204 (N_6204,N_5493,N_5905);
xnor U6205 (N_6205,N_5140,N_5290);
nor U6206 (N_6206,N_5095,N_5507);
or U6207 (N_6207,N_5600,N_5303);
nor U6208 (N_6208,N_5533,N_5025);
nor U6209 (N_6209,N_5909,N_5343);
and U6210 (N_6210,N_5490,N_5987);
nor U6211 (N_6211,N_5386,N_5404);
nand U6212 (N_6212,N_5815,N_5759);
nor U6213 (N_6213,N_5021,N_5096);
nor U6214 (N_6214,N_5491,N_5653);
or U6215 (N_6215,N_5014,N_5249);
and U6216 (N_6216,N_5532,N_5104);
and U6217 (N_6217,N_5718,N_5172);
xor U6218 (N_6218,N_5313,N_5655);
nor U6219 (N_6219,N_5341,N_5744);
or U6220 (N_6220,N_5286,N_5859);
nor U6221 (N_6221,N_5120,N_5880);
and U6222 (N_6222,N_5188,N_5138);
nor U6223 (N_6223,N_5864,N_5274);
or U6224 (N_6224,N_5566,N_5334);
xor U6225 (N_6225,N_5992,N_5672);
nand U6226 (N_6226,N_5203,N_5721);
nor U6227 (N_6227,N_5548,N_5079);
and U6228 (N_6228,N_5640,N_5497);
nand U6229 (N_6229,N_5823,N_5179);
or U6230 (N_6230,N_5501,N_5901);
nor U6231 (N_6231,N_5743,N_5381);
or U6232 (N_6232,N_5944,N_5354);
nor U6233 (N_6233,N_5829,N_5656);
and U6234 (N_6234,N_5828,N_5389);
and U6235 (N_6235,N_5311,N_5778);
nor U6236 (N_6236,N_5470,N_5258);
nand U6237 (N_6237,N_5261,N_5004);
or U6238 (N_6238,N_5054,N_5191);
xnor U6239 (N_6239,N_5112,N_5882);
xnor U6240 (N_6240,N_5269,N_5132);
xor U6241 (N_6241,N_5217,N_5719);
nand U6242 (N_6242,N_5369,N_5495);
xnor U6243 (N_6243,N_5919,N_5947);
nand U6244 (N_6244,N_5741,N_5001);
nand U6245 (N_6245,N_5050,N_5159);
or U6246 (N_6246,N_5671,N_5278);
nand U6247 (N_6247,N_5899,N_5157);
and U6248 (N_6248,N_5481,N_5866);
and U6249 (N_6249,N_5263,N_5007);
xor U6250 (N_6250,N_5562,N_5156);
or U6251 (N_6251,N_5991,N_5256);
xnor U6252 (N_6252,N_5542,N_5894);
and U6253 (N_6253,N_5160,N_5820);
and U6254 (N_6254,N_5023,N_5596);
nand U6255 (N_6255,N_5968,N_5858);
xor U6256 (N_6256,N_5900,N_5092);
and U6257 (N_6257,N_5180,N_5877);
nand U6258 (N_6258,N_5592,N_5485);
xor U6259 (N_6259,N_5225,N_5796);
nand U6260 (N_6260,N_5787,N_5661);
or U6261 (N_6261,N_5391,N_5626);
nand U6262 (N_6262,N_5700,N_5049);
and U6263 (N_6263,N_5243,N_5076);
and U6264 (N_6264,N_5551,N_5387);
or U6265 (N_6265,N_5315,N_5802);
or U6266 (N_6266,N_5797,N_5416);
xor U6267 (N_6267,N_5810,N_5657);
and U6268 (N_6268,N_5415,N_5927);
or U6269 (N_6269,N_5097,N_5632);
nand U6270 (N_6270,N_5254,N_5469);
or U6271 (N_6271,N_5454,N_5080);
or U6272 (N_6272,N_5956,N_5908);
xnor U6273 (N_6273,N_5970,N_5216);
or U6274 (N_6274,N_5594,N_5857);
nand U6275 (N_6275,N_5000,N_5665);
xnor U6276 (N_6276,N_5728,N_5182);
nor U6277 (N_6277,N_5570,N_5346);
or U6278 (N_6278,N_5255,N_5530);
and U6279 (N_6279,N_5984,N_5821);
nand U6280 (N_6280,N_5641,N_5706);
and U6281 (N_6281,N_5678,N_5407);
nor U6282 (N_6282,N_5427,N_5445);
and U6283 (N_6283,N_5367,N_5129);
xor U6284 (N_6284,N_5616,N_5867);
xor U6285 (N_6285,N_5405,N_5816);
or U6286 (N_6286,N_5161,N_5152);
or U6287 (N_6287,N_5804,N_5118);
nand U6288 (N_6288,N_5344,N_5664);
nor U6289 (N_6289,N_5291,N_5220);
xnor U6290 (N_6290,N_5400,N_5811);
and U6291 (N_6291,N_5609,N_5959);
xor U6292 (N_6292,N_5103,N_5342);
or U6293 (N_6293,N_5310,N_5064);
nand U6294 (N_6294,N_5523,N_5610);
or U6295 (N_6295,N_5306,N_5710);
nor U6296 (N_6296,N_5487,N_5760);
or U6297 (N_6297,N_5436,N_5163);
nor U6298 (N_6298,N_5950,N_5192);
or U6299 (N_6299,N_5745,N_5215);
nor U6300 (N_6300,N_5056,N_5207);
or U6301 (N_6301,N_5304,N_5704);
nand U6302 (N_6302,N_5421,N_5145);
xnor U6303 (N_6303,N_5554,N_5597);
and U6304 (N_6304,N_5210,N_5516);
nand U6305 (N_6305,N_5668,N_5625);
xnor U6306 (N_6306,N_5773,N_5652);
nand U6307 (N_6307,N_5111,N_5939);
nor U6308 (N_6308,N_5517,N_5863);
or U6309 (N_6309,N_5559,N_5638);
nand U6310 (N_6310,N_5251,N_5734);
and U6311 (N_6311,N_5382,N_5692);
xnor U6312 (N_6312,N_5726,N_5107);
and U6313 (N_6313,N_5181,N_5605);
xor U6314 (N_6314,N_5839,N_5946);
and U6315 (N_6315,N_5603,N_5589);
or U6316 (N_6316,N_5725,N_5361);
xor U6317 (N_6317,N_5360,N_5976);
or U6318 (N_6318,N_5189,N_5395);
nor U6319 (N_6319,N_5593,N_5637);
or U6320 (N_6320,N_5780,N_5015);
nor U6321 (N_6321,N_5747,N_5446);
nor U6322 (N_6322,N_5860,N_5032);
xnor U6323 (N_6323,N_5338,N_5550);
and U6324 (N_6324,N_5724,N_5674);
nand U6325 (N_6325,N_5856,N_5198);
nand U6326 (N_6326,N_5498,N_5048);
and U6327 (N_6327,N_5332,N_5393);
or U6328 (N_6328,N_5553,N_5817);
or U6329 (N_6329,N_5135,N_5193);
xnor U6330 (N_6330,N_5772,N_5447);
xnor U6331 (N_6331,N_5849,N_5608);
xor U6332 (N_6332,N_5078,N_5539);
and U6333 (N_6333,N_5945,N_5868);
nor U6334 (N_6334,N_5162,N_5786);
nor U6335 (N_6335,N_5292,N_5619);
nor U6336 (N_6336,N_5676,N_5685);
nor U6337 (N_6337,N_5331,N_5371);
nor U6338 (N_6338,N_5966,N_5126);
nand U6339 (N_6339,N_5663,N_5732);
xnor U6340 (N_6340,N_5733,N_5155);
nand U6341 (N_6341,N_5579,N_5799);
and U6342 (N_6342,N_5953,N_5294);
nand U6343 (N_6343,N_5133,N_5511);
nand U6344 (N_6344,N_5770,N_5598);
and U6345 (N_6345,N_5351,N_5065);
and U6346 (N_6346,N_5522,N_5627);
nor U6347 (N_6347,N_5988,N_5131);
nor U6348 (N_6348,N_5280,N_5869);
or U6349 (N_6349,N_5736,N_5755);
or U6350 (N_6350,N_5779,N_5876);
and U6351 (N_6351,N_5519,N_5767);
or U6352 (N_6352,N_5975,N_5690);
nand U6353 (N_6353,N_5813,N_5751);
xor U6354 (N_6354,N_5309,N_5283);
xor U6355 (N_6355,N_5437,N_5406);
and U6356 (N_6356,N_5184,N_5822);
nand U6357 (N_6357,N_5297,N_5689);
and U6358 (N_6358,N_5996,N_5808);
xnor U6359 (N_6359,N_5750,N_5224);
and U6360 (N_6360,N_5083,N_5362);
nor U6361 (N_6361,N_5529,N_5264);
and U6362 (N_6362,N_5284,N_5763);
or U6363 (N_6363,N_5230,N_5034);
nand U6364 (N_6364,N_5682,N_5105);
xor U6365 (N_6365,N_5197,N_5073);
or U6366 (N_6366,N_5488,N_5872);
nor U6367 (N_6367,N_5577,N_5578);
and U6368 (N_6368,N_5202,N_5881);
xnor U6369 (N_6369,N_5862,N_5479);
nor U6370 (N_6370,N_5323,N_5314);
nand U6371 (N_6371,N_5645,N_5357);
or U6372 (N_6372,N_5149,N_5433);
xor U6373 (N_6373,N_5827,N_5265);
nand U6374 (N_6374,N_5468,N_5492);
nor U6375 (N_6375,N_5587,N_5775);
or U6376 (N_6376,N_5586,N_5740);
nor U6377 (N_6377,N_5934,N_5318);
nand U6378 (N_6378,N_5228,N_5993);
and U6379 (N_6379,N_5694,N_5521);
nor U6380 (N_6380,N_5086,N_5764);
and U6381 (N_6381,N_5376,N_5417);
nor U6382 (N_6382,N_5892,N_5449);
nand U6383 (N_6383,N_5923,N_5865);
nand U6384 (N_6384,N_5561,N_5455);
nor U6385 (N_6385,N_5462,N_5793);
nand U6386 (N_6386,N_5585,N_5889);
or U6387 (N_6387,N_5613,N_5599);
xnor U6388 (N_6388,N_5903,N_5765);
and U6389 (N_6389,N_5441,N_5013);
xor U6390 (N_6390,N_5524,N_5713);
xnor U6391 (N_6391,N_5526,N_5660);
nor U6392 (N_6392,N_5709,N_5679);
and U6393 (N_6393,N_5981,N_5977);
nand U6394 (N_6394,N_5434,N_5273);
and U6395 (N_6395,N_5477,N_5871);
xor U6396 (N_6396,N_5174,N_5363);
xor U6397 (N_6397,N_5731,N_5633);
xnor U6398 (N_6398,N_5691,N_5410);
xnor U6399 (N_6399,N_5285,N_5366);
nor U6400 (N_6400,N_5932,N_5535);
xor U6401 (N_6401,N_5861,N_5739);
nor U6402 (N_6402,N_5484,N_5712);
nand U6403 (N_6403,N_5167,N_5384);
nand U6404 (N_6404,N_5912,N_5536);
and U6405 (N_6405,N_5574,N_5942);
nand U6406 (N_6406,N_5299,N_5794);
and U6407 (N_6407,N_5506,N_5791);
and U6408 (N_6408,N_5483,N_5527);
or U6409 (N_6409,N_5089,N_5142);
or U6410 (N_6410,N_5730,N_5588);
and U6411 (N_6411,N_5029,N_5897);
nand U6412 (N_6412,N_5186,N_5688);
or U6413 (N_6413,N_5168,N_5094);
nand U6414 (N_6414,N_5108,N_5240);
nand U6415 (N_6415,N_5677,N_5200);
and U6416 (N_6416,N_5531,N_5411);
xor U6417 (N_6417,N_5091,N_5238);
and U6418 (N_6418,N_5082,N_5024);
or U6419 (N_6419,N_5320,N_5088);
nand U6420 (N_6420,N_5963,N_5260);
nand U6421 (N_6421,N_5964,N_5737);
nor U6422 (N_6422,N_5830,N_5077);
nor U6423 (N_6423,N_5546,N_5356);
xor U6424 (N_6424,N_5634,N_5044);
xor U6425 (N_6425,N_5573,N_5150);
and U6426 (N_6426,N_5412,N_5647);
nor U6427 (N_6427,N_5965,N_5937);
xor U6428 (N_6428,N_5957,N_5898);
nor U6429 (N_6429,N_5440,N_5748);
nor U6430 (N_6430,N_5931,N_5971);
and U6431 (N_6431,N_5854,N_5339);
nor U6432 (N_6432,N_5752,N_5699);
or U6433 (N_6433,N_5241,N_5137);
nand U6434 (N_6434,N_5831,N_5675);
nor U6435 (N_6435,N_5749,N_5375);
and U6436 (N_6436,N_5635,N_5756);
xnor U6437 (N_6437,N_5194,N_5312);
xor U6438 (N_6438,N_5319,N_5451);
nand U6439 (N_6439,N_5429,N_5443);
or U6440 (N_6440,N_5219,N_5591);
nand U6441 (N_6441,N_5428,N_5612);
xor U6442 (N_6442,N_5460,N_5795);
or U6443 (N_6443,N_5717,N_5814);
or U6444 (N_6444,N_5990,N_5952);
and U6445 (N_6445,N_5420,N_5762);
nor U6446 (N_6446,N_5809,N_5475);
nor U6447 (N_6447,N_5761,N_5930);
or U6448 (N_6448,N_5350,N_5300);
xor U6449 (N_6449,N_5557,N_5196);
or U6450 (N_6450,N_5703,N_5575);
or U6451 (N_6451,N_5244,N_5011);
or U6452 (N_6452,N_5982,N_5045);
nand U6453 (N_6453,N_5785,N_5059);
and U6454 (N_6454,N_5442,N_5654);
xnor U6455 (N_6455,N_5986,N_5998);
nand U6456 (N_6456,N_5629,N_5502);
nand U6457 (N_6457,N_5237,N_5651);
or U6458 (N_6458,N_5681,N_5643);
and U6459 (N_6459,N_5834,N_5060);
xor U6460 (N_6460,N_5345,N_5520);
or U6461 (N_6461,N_5583,N_5922);
nor U6462 (N_6462,N_5305,N_5508);
xor U6463 (N_6463,N_5171,N_5985);
nand U6464 (N_6464,N_5624,N_5556);
or U6465 (N_6465,N_5211,N_5370);
or U6466 (N_6466,N_5392,N_5298);
or U6467 (N_6467,N_5232,N_5242);
and U6468 (N_6468,N_5994,N_5841);
nor U6469 (N_6469,N_5031,N_5753);
nand U6470 (N_6470,N_5087,N_5648);
or U6471 (N_6471,N_5547,N_5328);
xnor U6472 (N_6472,N_5052,N_5456);
xnor U6473 (N_6473,N_5639,N_5582);
and U6474 (N_6474,N_5102,N_5337);
nor U6475 (N_6475,N_5139,N_5175);
and U6476 (N_6476,N_5233,N_5929);
or U6477 (N_6477,N_5818,N_5941);
nand U6478 (N_6478,N_5513,N_5018);
nor U6479 (N_6479,N_5397,N_5333);
and U6480 (N_6480,N_5301,N_5130);
nor U6481 (N_6481,N_5012,N_5555);
nand U6482 (N_6482,N_5915,N_5723);
nor U6483 (N_6483,N_5093,N_5099);
xnor U6484 (N_6484,N_5466,N_5222);
and U6485 (N_6485,N_5835,N_5259);
nor U6486 (N_6486,N_5601,N_5667);
or U6487 (N_6487,N_5165,N_5448);
and U6488 (N_6488,N_5833,N_5549);
or U6489 (N_6489,N_5890,N_5414);
or U6490 (N_6490,N_5364,N_5870);
nor U6491 (N_6491,N_5195,N_5022);
xor U6492 (N_6492,N_5373,N_5960);
or U6493 (N_6493,N_5776,N_5825);
and U6494 (N_6494,N_5279,N_5057);
or U6495 (N_6495,N_5768,N_5063);
xnor U6496 (N_6496,N_5293,N_5771);
or U6497 (N_6497,N_5074,N_5066);
nor U6498 (N_6498,N_5697,N_5190);
xnor U6499 (N_6499,N_5805,N_5327);
nor U6500 (N_6500,N_5084,N_5157);
or U6501 (N_6501,N_5170,N_5209);
nor U6502 (N_6502,N_5085,N_5800);
or U6503 (N_6503,N_5511,N_5708);
nand U6504 (N_6504,N_5890,N_5243);
nor U6505 (N_6505,N_5455,N_5092);
nor U6506 (N_6506,N_5627,N_5953);
or U6507 (N_6507,N_5115,N_5862);
nand U6508 (N_6508,N_5402,N_5464);
nand U6509 (N_6509,N_5145,N_5144);
nand U6510 (N_6510,N_5141,N_5453);
nor U6511 (N_6511,N_5494,N_5793);
xnor U6512 (N_6512,N_5283,N_5727);
nor U6513 (N_6513,N_5211,N_5094);
and U6514 (N_6514,N_5644,N_5287);
or U6515 (N_6515,N_5806,N_5603);
and U6516 (N_6516,N_5413,N_5537);
nand U6517 (N_6517,N_5791,N_5730);
nand U6518 (N_6518,N_5608,N_5123);
nand U6519 (N_6519,N_5035,N_5613);
xor U6520 (N_6520,N_5772,N_5500);
nand U6521 (N_6521,N_5785,N_5745);
xor U6522 (N_6522,N_5982,N_5454);
xor U6523 (N_6523,N_5062,N_5779);
xnor U6524 (N_6524,N_5417,N_5332);
nor U6525 (N_6525,N_5678,N_5351);
nor U6526 (N_6526,N_5537,N_5763);
and U6527 (N_6527,N_5181,N_5393);
nand U6528 (N_6528,N_5260,N_5644);
nor U6529 (N_6529,N_5003,N_5043);
or U6530 (N_6530,N_5586,N_5297);
and U6531 (N_6531,N_5194,N_5376);
nand U6532 (N_6532,N_5199,N_5952);
or U6533 (N_6533,N_5578,N_5057);
and U6534 (N_6534,N_5798,N_5623);
nand U6535 (N_6535,N_5561,N_5132);
nand U6536 (N_6536,N_5605,N_5737);
and U6537 (N_6537,N_5561,N_5644);
or U6538 (N_6538,N_5907,N_5235);
nor U6539 (N_6539,N_5466,N_5762);
xnor U6540 (N_6540,N_5169,N_5815);
nor U6541 (N_6541,N_5092,N_5209);
or U6542 (N_6542,N_5147,N_5122);
nor U6543 (N_6543,N_5810,N_5473);
xnor U6544 (N_6544,N_5967,N_5903);
or U6545 (N_6545,N_5149,N_5926);
and U6546 (N_6546,N_5353,N_5906);
or U6547 (N_6547,N_5544,N_5398);
nand U6548 (N_6548,N_5852,N_5760);
nand U6549 (N_6549,N_5231,N_5826);
and U6550 (N_6550,N_5604,N_5307);
nor U6551 (N_6551,N_5120,N_5875);
or U6552 (N_6552,N_5545,N_5640);
nor U6553 (N_6553,N_5375,N_5461);
and U6554 (N_6554,N_5271,N_5979);
xnor U6555 (N_6555,N_5263,N_5367);
and U6556 (N_6556,N_5868,N_5334);
nand U6557 (N_6557,N_5968,N_5771);
nor U6558 (N_6558,N_5167,N_5836);
nand U6559 (N_6559,N_5918,N_5365);
or U6560 (N_6560,N_5253,N_5588);
nor U6561 (N_6561,N_5832,N_5662);
xnor U6562 (N_6562,N_5815,N_5103);
and U6563 (N_6563,N_5437,N_5829);
nor U6564 (N_6564,N_5253,N_5830);
nand U6565 (N_6565,N_5043,N_5082);
or U6566 (N_6566,N_5703,N_5396);
nand U6567 (N_6567,N_5699,N_5841);
nand U6568 (N_6568,N_5655,N_5961);
nand U6569 (N_6569,N_5456,N_5454);
and U6570 (N_6570,N_5884,N_5294);
nand U6571 (N_6571,N_5226,N_5902);
and U6572 (N_6572,N_5872,N_5345);
and U6573 (N_6573,N_5887,N_5682);
xnor U6574 (N_6574,N_5866,N_5010);
and U6575 (N_6575,N_5937,N_5255);
or U6576 (N_6576,N_5702,N_5695);
nand U6577 (N_6577,N_5920,N_5931);
nand U6578 (N_6578,N_5697,N_5027);
or U6579 (N_6579,N_5674,N_5861);
nand U6580 (N_6580,N_5980,N_5372);
or U6581 (N_6581,N_5786,N_5907);
nor U6582 (N_6582,N_5832,N_5553);
nand U6583 (N_6583,N_5251,N_5097);
xnor U6584 (N_6584,N_5135,N_5654);
nand U6585 (N_6585,N_5855,N_5259);
or U6586 (N_6586,N_5438,N_5430);
nor U6587 (N_6587,N_5227,N_5123);
xor U6588 (N_6588,N_5294,N_5523);
xnor U6589 (N_6589,N_5711,N_5250);
nor U6590 (N_6590,N_5120,N_5648);
nor U6591 (N_6591,N_5257,N_5120);
and U6592 (N_6592,N_5949,N_5766);
and U6593 (N_6593,N_5205,N_5531);
and U6594 (N_6594,N_5872,N_5469);
nand U6595 (N_6595,N_5629,N_5362);
nor U6596 (N_6596,N_5325,N_5298);
xnor U6597 (N_6597,N_5942,N_5806);
xor U6598 (N_6598,N_5269,N_5148);
nand U6599 (N_6599,N_5450,N_5665);
or U6600 (N_6600,N_5596,N_5265);
nor U6601 (N_6601,N_5157,N_5803);
xor U6602 (N_6602,N_5150,N_5265);
and U6603 (N_6603,N_5558,N_5747);
or U6604 (N_6604,N_5058,N_5493);
nand U6605 (N_6605,N_5104,N_5966);
nor U6606 (N_6606,N_5606,N_5356);
and U6607 (N_6607,N_5704,N_5326);
and U6608 (N_6608,N_5368,N_5069);
nor U6609 (N_6609,N_5498,N_5604);
and U6610 (N_6610,N_5248,N_5063);
and U6611 (N_6611,N_5397,N_5594);
nand U6612 (N_6612,N_5463,N_5122);
nand U6613 (N_6613,N_5264,N_5319);
xor U6614 (N_6614,N_5572,N_5629);
or U6615 (N_6615,N_5190,N_5557);
or U6616 (N_6616,N_5118,N_5823);
nand U6617 (N_6617,N_5419,N_5288);
or U6618 (N_6618,N_5500,N_5529);
or U6619 (N_6619,N_5875,N_5886);
xor U6620 (N_6620,N_5690,N_5804);
nor U6621 (N_6621,N_5518,N_5858);
or U6622 (N_6622,N_5753,N_5997);
xnor U6623 (N_6623,N_5787,N_5234);
xor U6624 (N_6624,N_5284,N_5515);
nor U6625 (N_6625,N_5602,N_5937);
and U6626 (N_6626,N_5723,N_5765);
and U6627 (N_6627,N_5361,N_5281);
and U6628 (N_6628,N_5592,N_5461);
or U6629 (N_6629,N_5582,N_5066);
xor U6630 (N_6630,N_5656,N_5388);
xor U6631 (N_6631,N_5574,N_5872);
and U6632 (N_6632,N_5226,N_5536);
and U6633 (N_6633,N_5363,N_5952);
xnor U6634 (N_6634,N_5388,N_5172);
nand U6635 (N_6635,N_5746,N_5137);
and U6636 (N_6636,N_5968,N_5772);
and U6637 (N_6637,N_5621,N_5118);
nor U6638 (N_6638,N_5577,N_5503);
or U6639 (N_6639,N_5847,N_5950);
and U6640 (N_6640,N_5514,N_5529);
and U6641 (N_6641,N_5934,N_5552);
nand U6642 (N_6642,N_5829,N_5595);
xor U6643 (N_6643,N_5313,N_5632);
or U6644 (N_6644,N_5833,N_5945);
nor U6645 (N_6645,N_5493,N_5236);
or U6646 (N_6646,N_5226,N_5623);
and U6647 (N_6647,N_5945,N_5646);
and U6648 (N_6648,N_5448,N_5113);
and U6649 (N_6649,N_5715,N_5036);
nand U6650 (N_6650,N_5570,N_5651);
nor U6651 (N_6651,N_5304,N_5028);
and U6652 (N_6652,N_5447,N_5759);
nand U6653 (N_6653,N_5928,N_5375);
or U6654 (N_6654,N_5473,N_5773);
nand U6655 (N_6655,N_5556,N_5257);
nor U6656 (N_6656,N_5202,N_5100);
xnor U6657 (N_6657,N_5604,N_5532);
and U6658 (N_6658,N_5489,N_5281);
xnor U6659 (N_6659,N_5398,N_5891);
xnor U6660 (N_6660,N_5326,N_5274);
nor U6661 (N_6661,N_5574,N_5465);
or U6662 (N_6662,N_5893,N_5131);
nand U6663 (N_6663,N_5944,N_5955);
xnor U6664 (N_6664,N_5361,N_5962);
xor U6665 (N_6665,N_5581,N_5468);
or U6666 (N_6666,N_5987,N_5374);
nand U6667 (N_6667,N_5550,N_5747);
nor U6668 (N_6668,N_5914,N_5123);
and U6669 (N_6669,N_5815,N_5985);
and U6670 (N_6670,N_5390,N_5487);
and U6671 (N_6671,N_5188,N_5102);
nor U6672 (N_6672,N_5778,N_5494);
nor U6673 (N_6673,N_5787,N_5579);
nor U6674 (N_6674,N_5803,N_5114);
xnor U6675 (N_6675,N_5048,N_5546);
xnor U6676 (N_6676,N_5196,N_5346);
nand U6677 (N_6677,N_5009,N_5047);
or U6678 (N_6678,N_5369,N_5787);
nor U6679 (N_6679,N_5113,N_5421);
nand U6680 (N_6680,N_5392,N_5635);
nand U6681 (N_6681,N_5531,N_5017);
nand U6682 (N_6682,N_5191,N_5354);
nor U6683 (N_6683,N_5365,N_5939);
and U6684 (N_6684,N_5186,N_5448);
or U6685 (N_6685,N_5051,N_5261);
xnor U6686 (N_6686,N_5703,N_5765);
xor U6687 (N_6687,N_5350,N_5403);
nand U6688 (N_6688,N_5122,N_5380);
or U6689 (N_6689,N_5741,N_5330);
and U6690 (N_6690,N_5630,N_5327);
or U6691 (N_6691,N_5616,N_5757);
nor U6692 (N_6692,N_5477,N_5688);
and U6693 (N_6693,N_5108,N_5649);
nor U6694 (N_6694,N_5820,N_5141);
nor U6695 (N_6695,N_5893,N_5624);
and U6696 (N_6696,N_5631,N_5550);
and U6697 (N_6697,N_5213,N_5337);
and U6698 (N_6698,N_5122,N_5373);
nor U6699 (N_6699,N_5286,N_5148);
xnor U6700 (N_6700,N_5817,N_5487);
xnor U6701 (N_6701,N_5048,N_5759);
nand U6702 (N_6702,N_5531,N_5064);
nand U6703 (N_6703,N_5767,N_5708);
nand U6704 (N_6704,N_5980,N_5378);
xnor U6705 (N_6705,N_5053,N_5675);
and U6706 (N_6706,N_5047,N_5100);
xnor U6707 (N_6707,N_5930,N_5825);
and U6708 (N_6708,N_5213,N_5176);
and U6709 (N_6709,N_5518,N_5911);
and U6710 (N_6710,N_5519,N_5724);
nor U6711 (N_6711,N_5149,N_5697);
nand U6712 (N_6712,N_5527,N_5579);
nor U6713 (N_6713,N_5017,N_5741);
nor U6714 (N_6714,N_5792,N_5375);
nand U6715 (N_6715,N_5122,N_5081);
or U6716 (N_6716,N_5945,N_5006);
nor U6717 (N_6717,N_5941,N_5228);
nor U6718 (N_6718,N_5393,N_5025);
xor U6719 (N_6719,N_5129,N_5042);
or U6720 (N_6720,N_5464,N_5727);
or U6721 (N_6721,N_5917,N_5244);
xor U6722 (N_6722,N_5660,N_5579);
or U6723 (N_6723,N_5045,N_5494);
nor U6724 (N_6724,N_5738,N_5125);
nand U6725 (N_6725,N_5626,N_5734);
xnor U6726 (N_6726,N_5760,N_5783);
nand U6727 (N_6727,N_5161,N_5971);
nand U6728 (N_6728,N_5018,N_5692);
nor U6729 (N_6729,N_5103,N_5715);
xnor U6730 (N_6730,N_5023,N_5494);
nor U6731 (N_6731,N_5372,N_5542);
nor U6732 (N_6732,N_5188,N_5166);
nor U6733 (N_6733,N_5599,N_5645);
or U6734 (N_6734,N_5206,N_5533);
or U6735 (N_6735,N_5431,N_5008);
nand U6736 (N_6736,N_5555,N_5299);
or U6737 (N_6737,N_5219,N_5637);
nand U6738 (N_6738,N_5276,N_5449);
nand U6739 (N_6739,N_5252,N_5513);
nand U6740 (N_6740,N_5423,N_5481);
nor U6741 (N_6741,N_5628,N_5406);
nand U6742 (N_6742,N_5057,N_5293);
and U6743 (N_6743,N_5592,N_5840);
xnor U6744 (N_6744,N_5284,N_5726);
and U6745 (N_6745,N_5964,N_5771);
xor U6746 (N_6746,N_5674,N_5444);
or U6747 (N_6747,N_5208,N_5790);
nor U6748 (N_6748,N_5806,N_5447);
or U6749 (N_6749,N_5733,N_5702);
and U6750 (N_6750,N_5120,N_5770);
nor U6751 (N_6751,N_5463,N_5539);
xnor U6752 (N_6752,N_5064,N_5125);
nor U6753 (N_6753,N_5738,N_5309);
nand U6754 (N_6754,N_5764,N_5107);
or U6755 (N_6755,N_5966,N_5047);
and U6756 (N_6756,N_5126,N_5437);
nand U6757 (N_6757,N_5597,N_5239);
or U6758 (N_6758,N_5693,N_5917);
and U6759 (N_6759,N_5568,N_5840);
nor U6760 (N_6760,N_5641,N_5749);
and U6761 (N_6761,N_5847,N_5014);
nand U6762 (N_6762,N_5588,N_5564);
nor U6763 (N_6763,N_5160,N_5915);
xor U6764 (N_6764,N_5111,N_5873);
and U6765 (N_6765,N_5422,N_5527);
nand U6766 (N_6766,N_5298,N_5748);
and U6767 (N_6767,N_5939,N_5535);
or U6768 (N_6768,N_5881,N_5806);
and U6769 (N_6769,N_5908,N_5280);
and U6770 (N_6770,N_5855,N_5015);
and U6771 (N_6771,N_5773,N_5842);
xnor U6772 (N_6772,N_5604,N_5100);
nor U6773 (N_6773,N_5659,N_5235);
nor U6774 (N_6774,N_5020,N_5023);
or U6775 (N_6775,N_5611,N_5665);
nand U6776 (N_6776,N_5120,N_5635);
nor U6777 (N_6777,N_5455,N_5071);
nor U6778 (N_6778,N_5660,N_5538);
or U6779 (N_6779,N_5951,N_5668);
or U6780 (N_6780,N_5695,N_5086);
nand U6781 (N_6781,N_5564,N_5753);
and U6782 (N_6782,N_5151,N_5920);
nand U6783 (N_6783,N_5222,N_5577);
nand U6784 (N_6784,N_5256,N_5281);
nor U6785 (N_6785,N_5747,N_5553);
xor U6786 (N_6786,N_5214,N_5603);
nor U6787 (N_6787,N_5807,N_5423);
nor U6788 (N_6788,N_5856,N_5808);
and U6789 (N_6789,N_5110,N_5162);
and U6790 (N_6790,N_5771,N_5378);
and U6791 (N_6791,N_5558,N_5867);
and U6792 (N_6792,N_5981,N_5258);
and U6793 (N_6793,N_5191,N_5431);
nand U6794 (N_6794,N_5084,N_5633);
and U6795 (N_6795,N_5497,N_5622);
or U6796 (N_6796,N_5264,N_5702);
xnor U6797 (N_6797,N_5471,N_5078);
nand U6798 (N_6798,N_5525,N_5916);
or U6799 (N_6799,N_5090,N_5182);
nand U6800 (N_6800,N_5430,N_5336);
or U6801 (N_6801,N_5910,N_5296);
nor U6802 (N_6802,N_5442,N_5385);
nor U6803 (N_6803,N_5277,N_5835);
nor U6804 (N_6804,N_5111,N_5962);
nor U6805 (N_6805,N_5086,N_5645);
xor U6806 (N_6806,N_5023,N_5338);
and U6807 (N_6807,N_5341,N_5643);
and U6808 (N_6808,N_5634,N_5016);
nor U6809 (N_6809,N_5306,N_5122);
nand U6810 (N_6810,N_5906,N_5027);
xor U6811 (N_6811,N_5677,N_5342);
xnor U6812 (N_6812,N_5398,N_5495);
nand U6813 (N_6813,N_5013,N_5415);
nand U6814 (N_6814,N_5763,N_5583);
nand U6815 (N_6815,N_5560,N_5159);
xnor U6816 (N_6816,N_5846,N_5732);
nor U6817 (N_6817,N_5667,N_5751);
or U6818 (N_6818,N_5734,N_5133);
nand U6819 (N_6819,N_5509,N_5828);
xnor U6820 (N_6820,N_5403,N_5908);
xnor U6821 (N_6821,N_5460,N_5765);
xnor U6822 (N_6822,N_5181,N_5777);
or U6823 (N_6823,N_5360,N_5711);
or U6824 (N_6824,N_5938,N_5506);
nor U6825 (N_6825,N_5598,N_5750);
and U6826 (N_6826,N_5242,N_5499);
xor U6827 (N_6827,N_5018,N_5151);
and U6828 (N_6828,N_5884,N_5123);
xnor U6829 (N_6829,N_5670,N_5927);
nand U6830 (N_6830,N_5833,N_5857);
and U6831 (N_6831,N_5032,N_5873);
and U6832 (N_6832,N_5127,N_5696);
or U6833 (N_6833,N_5122,N_5343);
or U6834 (N_6834,N_5135,N_5544);
nand U6835 (N_6835,N_5999,N_5976);
xnor U6836 (N_6836,N_5802,N_5239);
xnor U6837 (N_6837,N_5277,N_5068);
nor U6838 (N_6838,N_5513,N_5870);
nor U6839 (N_6839,N_5771,N_5572);
and U6840 (N_6840,N_5570,N_5614);
or U6841 (N_6841,N_5199,N_5841);
nor U6842 (N_6842,N_5750,N_5975);
or U6843 (N_6843,N_5069,N_5261);
or U6844 (N_6844,N_5634,N_5275);
xor U6845 (N_6845,N_5150,N_5775);
or U6846 (N_6846,N_5900,N_5300);
nand U6847 (N_6847,N_5379,N_5335);
nand U6848 (N_6848,N_5661,N_5579);
nand U6849 (N_6849,N_5625,N_5779);
or U6850 (N_6850,N_5811,N_5926);
xor U6851 (N_6851,N_5866,N_5531);
nand U6852 (N_6852,N_5294,N_5696);
and U6853 (N_6853,N_5350,N_5453);
or U6854 (N_6854,N_5751,N_5925);
and U6855 (N_6855,N_5576,N_5353);
nand U6856 (N_6856,N_5787,N_5838);
nor U6857 (N_6857,N_5866,N_5553);
nand U6858 (N_6858,N_5782,N_5537);
and U6859 (N_6859,N_5688,N_5564);
xnor U6860 (N_6860,N_5721,N_5129);
and U6861 (N_6861,N_5307,N_5323);
nor U6862 (N_6862,N_5488,N_5711);
xor U6863 (N_6863,N_5566,N_5614);
and U6864 (N_6864,N_5125,N_5223);
xnor U6865 (N_6865,N_5244,N_5024);
nor U6866 (N_6866,N_5934,N_5891);
xor U6867 (N_6867,N_5943,N_5315);
or U6868 (N_6868,N_5438,N_5474);
or U6869 (N_6869,N_5646,N_5014);
xnor U6870 (N_6870,N_5332,N_5541);
xnor U6871 (N_6871,N_5077,N_5977);
and U6872 (N_6872,N_5980,N_5557);
nor U6873 (N_6873,N_5393,N_5473);
nand U6874 (N_6874,N_5622,N_5036);
and U6875 (N_6875,N_5275,N_5014);
xnor U6876 (N_6876,N_5135,N_5015);
and U6877 (N_6877,N_5482,N_5853);
nand U6878 (N_6878,N_5303,N_5988);
xor U6879 (N_6879,N_5224,N_5232);
or U6880 (N_6880,N_5736,N_5560);
nor U6881 (N_6881,N_5544,N_5440);
nor U6882 (N_6882,N_5142,N_5631);
nand U6883 (N_6883,N_5160,N_5391);
or U6884 (N_6884,N_5534,N_5803);
or U6885 (N_6885,N_5440,N_5099);
xor U6886 (N_6886,N_5053,N_5907);
or U6887 (N_6887,N_5764,N_5620);
nand U6888 (N_6888,N_5680,N_5060);
or U6889 (N_6889,N_5187,N_5986);
or U6890 (N_6890,N_5746,N_5890);
nor U6891 (N_6891,N_5988,N_5320);
or U6892 (N_6892,N_5042,N_5281);
nand U6893 (N_6893,N_5727,N_5531);
nand U6894 (N_6894,N_5387,N_5069);
nand U6895 (N_6895,N_5519,N_5805);
nand U6896 (N_6896,N_5543,N_5613);
or U6897 (N_6897,N_5686,N_5073);
or U6898 (N_6898,N_5793,N_5472);
xnor U6899 (N_6899,N_5532,N_5246);
nand U6900 (N_6900,N_5439,N_5628);
and U6901 (N_6901,N_5030,N_5144);
xor U6902 (N_6902,N_5105,N_5384);
nand U6903 (N_6903,N_5503,N_5282);
nand U6904 (N_6904,N_5065,N_5030);
or U6905 (N_6905,N_5372,N_5056);
and U6906 (N_6906,N_5876,N_5735);
or U6907 (N_6907,N_5609,N_5924);
or U6908 (N_6908,N_5506,N_5079);
nor U6909 (N_6909,N_5075,N_5288);
or U6910 (N_6910,N_5489,N_5302);
nor U6911 (N_6911,N_5217,N_5425);
nor U6912 (N_6912,N_5394,N_5763);
nor U6913 (N_6913,N_5128,N_5188);
xnor U6914 (N_6914,N_5525,N_5348);
nand U6915 (N_6915,N_5981,N_5420);
nor U6916 (N_6916,N_5004,N_5648);
nor U6917 (N_6917,N_5059,N_5679);
xnor U6918 (N_6918,N_5013,N_5928);
or U6919 (N_6919,N_5962,N_5617);
xor U6920 (N_6920,N_5104,N_5812);
or U6921 (N_6921,N_5145,N_5673);
xor U6922 (N_6922,N_5651,N_5967);
nand U6923 (N_6923,N_5947,N_5401);
nand U6924 (N_6924,N_5324,N_5760);
and U6925 (N_6925,N_5190,N_5143);
or U6926 (N_6926,N_5223,N_5053);
nand U6927 (N_6927,N_5138,N_5067);
and U6928 (N_6928,N_5796,N_5705);
xnor U6929 (N_6929,N_5492,N_5571);
and U6930 (N_6930,N_5054,N_5996);
nand U6931 (N_6931,N_5598,N_5951);
xor U6932 (N_6932,N_5625,N_5770);
xor U6933 (N_6933,N_5706,N_5502);
and U6934 (N_6934,N_5601,N_5086);
or U6935 (N_6935,N_5959,N_5098);
and U6936 (N_6936,N_5611,N_5515);
or U6937 (N_6937,N_5893,N_5669);
nand U6938 (N_6938,N_5982,N_5978);
xor U6939 (N_6939,N_5481,N_5247);
nor U6940 (N_6940,N_5761,N_5979);
and U6941 (N_6941,N_5423,N_5899);
nand U6942 (N_6942,N_5051,N_5123);
or U6943 (N_6943,N_5793,N_5413);
or U6944 (N_6944,N_5537,N_5475);
or U6945 (N_6945,N_5639,N_5852);
or U6946 (N_6946,N_5328,N_5457);
and U6947 (N_6947,N_5539,N_5187);
nand U6948 (N_6948,N_5949,N_5139);
or U6949 (N_6949,N_5587,N_5107);
or U6950 (N_6950,N_5059,N_5566);
nor U6951 (N_6951,N_5038,N_5406);
nor U6952 (N_6952,N_5641,N_5530);
and U6953 (N_6953,N_5981,N_5845);
or U6954 (N_6954,N_5334,N_5588);
nand U6955 (N_6955,N_5504,N_5439);
xnor U6956 (N_6956,N_5606,N_5495);
nor U6957 (N_6957,N_5675,N_5912);
or U6958 (N_6958,N_5574,N_5812);
or U6959 (N_6959,N_5529,N_5197);
nand U6960 (N_6960,N_5718,N_5771);
nand U6961 (N_6961,N_5924,N_5017);
or U6962 (N_6962,N_5295,N_5529);
and U6963 (N_6963,N_5220,N_5505);
or U6964 (N_6964,N_5143,N_5628);
xor U6965 (N_6965,N_5740,N_5239);
xor U6966 (N_6966,N_5421,N_5149);
and U6967 (N_6967,N_5845,N_5245);
and U6968 (N_6968,N_5469,N_5294);
xor U6969 (N_6969,N_5790,N_5374);
xor U6970 (N_6970,N_5914,N_5120);
and U6971 (N_6971,N_5868,N_5675);
nor U6972 (N_6972,N_5395,N_5293);
nand U6973 (N_6973,N_5864,N_5919);
or U6974 (N_6974,N_5255,N_5405);
xnor U6975 (N_6975,N_5915,N_5024);
nand U6976 (N_6976,N_5765,N_5774);
nor U6977 (N_6977,N_5581,N_5181);
nand U6978 (N_6978,N_5396,N_5976);
nand U6979 (N_6979,N_5887,N_5469);
nor U6980 (N_6980,N_5892,N_5502);
and U6981 (N_6981,N_5156,N_5839);
and U6982 (N_6982,N_5004,N_5334);
nand U6983 (N_6983,N_5797,N_5868);
and U6984 (N_6984,N_5402,N_5287);
xnor U6985 (N_6985,N_5914,N_5597);
nor U6986 (N_6986,N_5750,N_5684);
or U6987 (N_6987,N_5139,N_5215);
and U6988 (N_6988,N_5337,N_5289);
or U6989 (N_6989,N_5295,N_5352);
xnor U6990 (N_6990,N_5639,N_5076);
and U6991 (N_6991,N_5951,N_5081);
nand U6992 (N_6992,N_5878,N_5695);
nor U6993 (N_6993,N_5386,N_5214);
xor U6994 (N_6994,N_5065,N_5792);
xnor U6995 (N_6995,N_5549,N_5000);
nor U6996 (N_6996,N_5978,N_5310);
or U6997 (N_6997,N_5488,N_5201);
xor U6998 (N_6998,N_5478,N_5069);
xor U6999 (N_6999,N_5323,N_5876);
nand U7000 (N_7000,N_6222,N_6583);
nand U7001 (N_7001,N_6199,N_6787);
and U7002 (N_7002,N_6759,N_6336);
nor U7003 (N_7003,N_6897,N_6414);
or U7004 (N_7004,N_6916,N_6044);
or U7005 (N_7005,N_6821,N_6774);
or U7006 (N_7006,N_6520,N_6541);
nand U7007 (N_7007,N_6797,N_6272);
and U7008 (N_7008,N_6205,N_6179);
and U7009 (N_7009,N_6572,N_6319);
nand U7010 (N_7010,N_6437,N_6038);
or U7011 (N_7011,N_6534,N_6650);
or U7012 (N_7012,N_6761,N_6428);
nand U7013 (N_7013,N_6213,N_6555);
and U7014 (N_7014,N_6031,N_6683);
xnor U7015 (N_7015,N_6106,N_6218);
and U7016 (N_7016,N_6411,N_6753);
and U7017 (N_7017,N_6508,N_6907);
nor U7018 (N_7018,N_6851,N_6206);
nand U7019 (N_7019,N_6515,N_6030);
and U7020 (N_7020,N_6754,N_6283);
nor U7021 (N_7021,N_6624,N_6450);
nand U7022 (N_7022,N_6798,N_6826);
nand U7023 (N_7023,N_6169,N_6291);
nor U7024 (N_7024,N_6153,N_6101);
nand U7025 (N_7025,N_6945,N_6524);
nand U7026 (N_7026,N_6873,N_6081);
xor U7027 (N_7027,N_6785,N_6056);
nand U7028 (N_7028,N_6965,N_6117);
and U7029 (N_7029,N_6582,N_6440);
nor U7030 (N_7030,N_6167,N_6870);
xnor U7031 (N_7031,N_6055,N_6135);
nor U7032 (N_7032,N_6111,N_6337);
or U7033 (N_7033,N_6773,N_6838);
nor U7034 (N_7034,N_6015,N_6629);
and U7035 (N_7035,N_6180,N_6615);
nand U7036 (N_7036,N_6090,N_6721);
nor U7037 (N_7037,N_6995,N_6365);
or U7038 (N_7038,N_6134,N_6751);
xnor U7039 (N_7039,N_6538,N_6128);
nor U7040 (N_7040,N_6045,N_6529);
nand U7041 (N_7041,N_6458,N_6631);
xor U7042 (N_7042,N_6516,N_6221);
nand U7043 (N_7043,N_6509,N_6868);
nand U7044 (N_7044,N_6547,N_6843);
xnor U7045 (N_7045,N_6560,N_6522);
or U7046 (N_7046,N_6658,N_6715);
and U7047 (N_7047,N_6493,N_6014);
xnor U7048 (N_7048,N_6284,N_6643);
xnor U7049 (N_7049,N_6289,N_6392);
nand U7050 (N_7050,N_6967,N_6871);
nand U7051 (N_7051,N_6640,N_6404);
nor U7052 (N_7052,N_6766,N_6910);
nand U7053 (N_7053,N_6237,N_6489);
nand U7054 (N_7054,N_6905,N_6588);
nand U7055 (N_7055,N_6646,N_6723);
nor U7056 (N_7056,N_6926,N_6184);
and U7057 (N_7057,N_6784,N_6394);
or U7058 (N_7058,N_6755,N_6164);
nand U7059 (N_7059,N_6756,N_6483);
and U7060 (N_7060,N_6687,N_6035);
xor U7061 (N_7061,N_6518,N_6811);
nand U7062 (N_7062,N_6147,N_6636);
nand U7063 (N_7063,N_6098,N_6127);
nand U7064 (N_7064,N_6660,N_6827);
xnor U7065 (N_7065,N_6338,N_6924);
nor U7066 (N_7066,N_6677,N_6885);
nand U7067 (N_7067,N_6341,N_6302);
nor U7068 (N_7068,N_6920,N_6275);
nor U7069 (N_7069,N_6079,N_6639);
or U7070 (N_7070,N_6463,N_6674);
xnor U7071 (N_7071,N_6514,N_6653);
nand U7072 (N_7072,N_6500,N_6625);
xor U7073 (N_7073,N_6412,N_6681);
or U7074 (N_7074,N_6857,N_6778);
nor U7075 (N_7075,N_6737,N_6672);
or U7076 (N_7076,N_6110,N_6919);
nand U7077 (N_7077,N_6542,N_6148);
or U7078 (N_7078,N_6251,N_6570);
or U7079 (N_7079,N_6379,N_6280);
nand U7080 (N_7080,N_6068,N_6757);
and U7081 (N_7081,N_6490,N_6353);
or U7082 (N_7082,N_6256,N_6861);
or U7083 (N_7083,N_6507,N_6913);
nand U7084 (N_7084,N_6259,N_6896);
xor U7085 (N_7085,N_6791,N_6510);
and U7086 (N_7086,N_6075,N_6113);
and U7087 (N_7087,N_6427,N_6977);
nand U7088 (N_7088,N_6480,N_6645);
nor U7089 (N_7089,N_6479,N_6799);
or U7090 (N_7090,N_6354,N_6026);
and U7091 (N_7091,N_6496,N_6579);
nand U7092 (N_7092,N_6183,N_6501);
and U7093 (N_7093,N_6462,N_6215);
xnor U7094 (N_7094,N_6065,N_6929);
xnor U7095 (N_7095,N_6904,N_6159);
nor U7096 (N_7096,N_6264,N_6422);
or U7097 (N_7097,N_6123,N_6989);
or U7098 (N_7098,N_6220,N_6714);
xnor U7099 (N_7099,N_6842,N_6959);
nor U7100 (N_7100,N_6602,N_6418);
or U7101 (N_7101,N_6066,N_6409);
and U7102 (N_7102,N_6670,N_6953);
or U7103 (N_7103,N_6832,N_6362);
and U7104 (N_7104,N_6062,N_6740);
nor U7105 (N_7105,N_6387,N_6684);
or U7106 (N_7106,N_6777,N_6049);
or U7107 (N_7107,N_6342,N_6494);
and U7108 (N_7108,N_6266,N_6517);
and U7109 (N_7109,N_6734,N_6241);
or U7110 (N_7110,N_6344,N_6512);
nand U7111 (N_7111,N_6425,N_6872);
and U7112 (N_7112,N_6020,N_6545);
xor U7113 (N_7113,N_6993,N_6285);
nor U7114 (N_7114,N_6277,N_6688);
nor U7115 (N_7115,N_6532,N_6188);
or U7116 (N_7116,N_6381,N_6162);
nor U7117 (N_7117,N_6760,N_6890);
xor U7118 (N_7118,N_6617,N_6958);
and U7119 (N_7119,N_6722,N_6423);
or U7120 (N_7120,N_6666,N_6887);
xor U7121 (N_7121,N_6587,N_6668);
xor U7122 (N_7122,N_6018,N_6004);
nor U7123 (N_7123,N_6611,N_6007);
or U7124 (N_7124,N_6836,N_6185);
nor U7125 (N_7125,N_6380,N_6013);
and U7126 (N_7126,N_6499,N_6738);
nor U7127 (N_7127,N_6306,N_6553);
nor U7128 (N_7128,N_6008,N_6828);
xor U7129 (N_7129,N_6069,N_6996);
and U7130 (N_7130,N_6519,N_6361);
nand U7131 (N_7131,N_6969,N_6772);
and U7132 (N_7132,N_6096,N_6983);
or U7133 (N_7133,N_6824,N_6957);
or U7134 (N_7134,N_6936,N_6619);
nand U7135 (N_7135,N_6589,N_6931);
xor U7136 (N_7136,N_6009,N_6837);
nor U7137 (N_7137,N_6476,N_6024);
xor U7138 (N_7138,N_6349,N_6248);
and U7139 (N_7139,N_6895,N_6716);
or U7140 (N_7140,N_6933,N_6922);
and U7141 (N_7141,N_6229,N_6961);
nand U7142 (N_7142,N_6002,N_6810);
or U7143 (N_7143,N_6234,N_6955);
xnor U7144 (N_7144,N_6119,N_6097);
xor U7145 (N_7145,N_6564,N_6999);
nand U7146 (N_7146,N_6987,N_6276);
nand U7147 (N_7147,N_6825,N_6161);
nand U7148 (N_7148,N_6556,N_6962);
nand U7149 (N_7149,N_6432,N_6847);
and U7150 (N_7150,N_6892,N_6511);
or U7151 (N_7151,N_6858,N_6051);
xnor U7152 (N_7152,N_6224,N_6889);
or U7153 (N_7153,N_6917,N_6431);
xnor U7154 (N_7154,N_6976,N_6124);
and U7155 (N_7155,N_6930,N_6357);
or U7156 (N_7156,N_6840,N_6614);
and U7157 (N_7157,N_6800,N_6523);
nand U7158 (N_7158,N_6401,N_6765);
xor U7159 (N_7159,N_6731,N_6782);
xnor U7160 (N_7160,N_6654,N_6152);
nand U7161 (N_7161,N_6769,N_6807);
and U7162 (N_7162,N_6812,N_6239);
and U7163 (N_7163,N_6621,N_6442);
and U7164 (N_7164,N_6963,N_6537);
nand U7165 (N_7165,N_6574,N_6292);
or U7166 (N_7166,N_6893,N_6728);
or U7167 (N_7167,N_6464,N_6622);
nand U7168 (N_7168,N_6763,N_6703);
nor U7169 (N_7169,N_6439,N_6181);
xnor U7170 (N_7170,N_6371,N_6059);
nor U7171 (N_7171,N_6941,N_6375);
or U7172 (N_7172,N_6042,N_6567);
xnor U7173 (N_7173,N_6290,N_6313);
xor U7174 (N_7174,N_6656,N_6608);
nor U7175 (N_7175,N_6942,N_6938);
xor U7176 (N_7176,N_6947,N_6638);
xor U7177 (N_7177,N_6350,N_6746);
nand U7178 (N_7178,N_6815,N_6869);
xor U7179 (N_7179,N_6407,N_6103);
nor U7180 (N_7180,N_6317,N_6637);
and U7181 (N_7181,N_6690,N_6804);
and U7182 (N_7182,N_6084,N_6443);
xor U7183 (N_7183,N_6590,N_6813);
and U7184 (N_7184,N_6005,N_6664);
xor U7185 (N_7185,N_6258,N_6633);
and U7186 (N_7186,N_6894,N_6487);
and U7187 (N_7187,N_6729,N_6793);
or U7188 (N_7188,N_6739,N_6197);
nor U7189 (N_7189,N_6121,N_6415);
xor U7190 (N_7190,N_6441,N_6707);
nand U7191 (N_7191,N_6540,N_6378);
nand U7192 (N_7192,N_6484,N_6974);
and U7193 (N_7193,N_6328,N_6805);
and U7194 (N_7194,N_6448,N_6054);
nand U7195 (N_7195,N_6607,N_6166);
or U7196 (N_7196,N_6300,N_6599);
and U7197 (N_7197,N_6486,N_6543);
nand U7198 (N_7198,N_6446,N_6419);
nor U7199 (N_7199,N_6359,N_6549);
and U7200 (N_7200,N_6454,N_6834);
nor U7201 (N_7201,N_6250,N_6318);
nor U7202 (N_7202,N_6899,N_6597);
nand U7203 (N_7203,N_6029,N_6456);
nand U7204 (N_7204,N_6485,N_6087);
or U7205 (N_7205,N_6080,N_6309);
xor U7206 (N_7206,N_6665,N_6100);
xor U7207 (N_7207,N_6848,N_6841);
or U7208 (N_7208,N_6600,N_6470);
and U7209 (N_7209,N_6860,N_6240);
nand U7210 (N_7210,N_6612,N_6606);
nor U7211 (N_7211,N_6023,N_6028);
or U7212 (N_7212,N_6770,N_6580);
xor U7213 (N_7213,N_6880,N_6434);
xnor U7214 (N_7214,N_6742,N_6189);
or U7215 (N_7215,N_6286,N_6488);
and U7216 (N_7216,N_6498,N_6705);
nor U7217 (N_7217,N_6390,N_6964);
nand U7218 (N_7218,N_6946,N_6561);
or U7219 (N_7219,N_6471,N_6844);
and U7220 (N_7220,N_6634,N_6943);
nor U7221 (N_7221,N_6830,N_6596);
nand U7222 (N_7222,N_6850,N_6505);
nand U7223 (N_7223,N_6262,N_6326);
or U7224 (N_7224,N_6058,N_6203);
nand U7225 (N_7225,N_6720,N_6991);
nor U7226 (N_7226,N_6116,N_6376);
xor U7227 (N_7227,N_6822,N_6748);
nor U7228 (N_7228,N_6649,N_6829);
and U7229 (N_7229,N_6346,N_6339);
xnor U7230 (N_7230,N_6052,N_6254);
nand U7231 (N_7231,N_6806,N_6244);
nand U7232 (N_7232,N_6741,N_6403);
nor U7233 (N_7233,N_6017,N_6710);
or U7234 (N_7234,N_6122,N_6576);
nand U7235 (N_7235,N_6949,N_6261);
or U7236 (N_7236,N_6492,N_6037);
or U7237 (N_7237,N_6584,N_6466);
xnor U7238 (N_7238,N_6310,N_6544);
nand U7239 (N_7239,N_6662,N_6077);
nand U7240 (N_7240,N_6709,N_6695);
nand U7241 (N_7241,N_6546,N_6884);
and U7242 (N_7242,N_6420,N_6182);
nor U7243 (N_7243,N_6652,N_6565);
nor U7244 (N_7244,N_6104,N_6911);
or U7245 (N_7245,N_6444,N_6789);
xor U7246 (N_7246,N_6736,N_6112);
nand U7247 (N_7247,N_6973,N_6503);
nand U7248 (N_7248,N_6475,N_6552);
or U7249 (N_7249,N_6726,N_6201);
xor U7250 (N_7250,N_6831,N_6330);
nand U7251 (N_7251,N_6360,N_6253);
nor U7252 (N_7252,N_6853,N_6088);
xor U7253 (N_7253,N_6718,N_6998);
or U7254 (N_7254,N_6156,N_6732);
nor U7255 (N_7255,N_6818,N_6495);
nand U7256 (N_7256,N_6888,N_6143);
and U7257 (N_7257,N_6416,N_6061);
or U7258 (N_7258,N_6385,N_6078);
nand U7259 (N_7259,N_6288,N_6591);
or U7260 (N_7260,N_6956,N_6796);
nand U7261 (N_7261,N_6136,N_6814);
nand U7262 (N_7262,N_6655,N_6735);
xnor U7263 (N_7263,N_6578,N_6883);
and U7264 (N_7264,N_6083,N_6165);
or U7265 (N_7265,N_6265,N_6295);
nand U7266 (N_7266,N_6041,N_6954);
nor U7267 (N_7267,N_6010,N_6238);
nand U7268 (N_7268,N_6725,N_6208);
xnor U7269 (N_7269,N_6391,N_6314);
nor U7270 (N_7270,N_6383,N_6388);
and U7271 (N_7271,N_6355,N_6610);
nor U7272 (N_7272,N_6481,N_6193);
nand U7273 (N_7273,N_6105,N_6115);
and U7274 (N_7274,N_6630,N_6327);
nor U7275 (N_7275,N_6712,N_6866);
or U7276 (N_7276,N_6173,N_6025);
nand U7277 (N_7277,N_6170,N_6150);
nand U7278 (N_7278,N_6747,N_6141);
xnor U7279 (N_7279,N_6781,N_6790);
and U7280 (N_7280,N_6076,N_6269);
nand U7281 (N_7281,N_6698,N_6303);
nor U7282 (N_7282,N_6803,N_6794);
xor U7283 (N_7283,N_6278,N_6347);
nand U7284 (N_7284,N_6348,N_6859);
xnor U7285 (N_7285,N_6990,N_6363);
or U7286 (N_7286,N_6909,N_6155);
and U7287 (N_7287,N_6377,N_6396);
or U7288 (N_7288,N_6569,N_6095);
nand U7289 (N_7289,N_6089,N_6114);
xor U7290 (N_7290,N_6242,N_6163);
or U7291 (N_7291,N_6226,N_6981);
nor U7292 (N_7292,N_6057,N_6594);
xor U7293 (N_7293,N_6281,N_6006);
and U7294 (N_7294,N_6701,N_6219);
nor U7295 (N_7295,N_6408,N_6764);
or U7296 (N_7296,N_6533,N_6817);
and U7297 (N_7297,N_6642,N_6568);
and U7298 (N_7298,N_6539,N_6675);
or U7299 (N_7299,N_6724,N_6273);
and U7300 (N_7300,N_6255,N_6146);
nor U7301 (N_7301,N_6863,N_6072);
nand U7302 (N_7302,N_6762,N_6648);
xor U7303 (N_7303,N_6506,N_6340);
xnor U7304 (N_7304,N_6073,N_6384);
and U7305 (N_7305,N_6557,N_6074);
or U7306 (N_7306,N_6875,N_6249);
nand U7307 (N_7307,N_6216,N_6329);
or U7308 (N_7308,N_6985,N_6402);
nor U7309 (N_7309,N_6585,N_6345);
nand U7310 (N_7310,N_6022,N_6187);
or U7311 (N_7311,N_6382,N_6433);
xnor U7312 (N_7312,N_6852,N_6477);
or U7313 (N_7313,N_6039,N_6521);
nor U7314 (N_7314,N_6043,N_6680);
or U7315 (N_7315,N_6125,N_6914);
nor U7316 (N_7316,N_6616,N_6154);
nor U7317 (N_7317,N_6386,N_6951);
and U7318 (N_7318,N_6398,N_6268);
or U7319 (N_7319,N_6823,N_6944);
and U7320 (N_7320,N_6536,N_6312);
and U7321 (N_7321,N_6000,N_6050);
and U7322 (N_7322,N_6700,N_6228);
or U7323 (N_7323,N_6697,N_6053);
and U7324 (N_7324,N_6373,N_6935);
nand U7325 (N_7325,N_6708,N_6535);
xnor U7326 (N_7326,N_6632,N_6177);
xnor U7327 (N_7327,N_6395,N_6595);
and U7328 (N_7328,N_6145,N_6118);
or U7329 (N_7329,N_6452,N_6877);
nor U7330 (N_7330,N_6623,N_6855);
and U7331 (N_7331,N_6711,N_6635);
xor U7332 (N_7332,N_6968,N_6603);
xor U7333 (N_7333,N_6468,N_6676);
nor U7334 (N_7334,N_6093,N_6399);
or U7335 (N_7335,N_6601,N_6862);
nand U7336 (N_7336,N_6370,N_6997);
nor U7337 (N_7337,N_6129,N_6333);
or U7338 (N_7338,N_6369,N_6270);
xnor U7339 (N_7339,N_6912,N_6232);
nand U7340 (N_7340,N_6527,N_6036);
nor U7341 (N_7341,N_6854,N_6451);
and U7342 (N_7342,N_6316,N_6694);
nand U7343 (N_7343,N_6194,N_6245);
xor U7344 (N_7344,N_6592,N_6801);
and U7345 (N_7345,N_6727,N_6984);
and U7346 (N_7346,N_6667,N_6663);
xor U7347 (N_7347,N_6651,N_6372);
xor U7348 (N_7348,N_6882,N_6358);
xnor U7349 (N_7349,N_6192,N_6833);
nand U7350 (N_7350,N_6158,N_6323);
nor U7351 (N_7351,N_6246,N_6641);
and U7352 (N_7352,N_6932,N_6461);
nand U7353 (N_7353,N_6906,N_6478);
xor U7354 (N_7354,N_6299,N_6132);
nor U7355 (N_7355,N_6693,N_6048);
xor U7356 (N_7356,N_6332,N_6881);
and U7357 (N_7357,N_6139,N_6012);
nor U7358 (N_7358,N_6502,N_6260);
xnor U7359 (N_7359,N_6575,N_6469);
or U7360 (N_7360,N_6436,N_6356);
xnor U7361 (N_7361,N_6702,N_6294);
nand U7362 (N_7362,N_6067,N_6898);
or U7363 (N_7363,N_6447,N_6682);
xor U7364 (N_7364,N_6421,N_6138);
xnor U7365 (N_7365,N_6032,N_6657);
xnor U7366 (N_7366,N_6678,N_6927);
or U7367 (N_7367,N_6047,N_6768);
nand U7368 (N_7368,N_6178,N_6426);
and U7369 (N_7369,N_6952,N_6343);
nor U7370 (N_7370,N_6970,N_6168);
and U7371 (N_7371,N_6472,N_6424);
and U7372 (N_7372,N_6978,N_6788);
or U7373 (N_7373,N_6429,N_6324);
or U7374 (N_7374,N_6525,N_6878);
or U7375 (N_7375,N_6200,N_6752);
or U7376 (N_7376,N_6779,N_6107);
nor U7377 (N_7377,N_6235,N_6937);
nor U7378 (N_7378,N_6802,N_6971);
or U7379 (N_7379,N_6460,N_6367);
xnor U7380 (N_7380,N_6102,N_6467);
nor U7381 (N_7381,N_6186,N_6531);
or U7382 (N_7382,N_6749,N_6322);
or U7383 (N_7383,N_6679,N_6389);
nand U7384 (N_7384,N_6795,N_6307);
or U7385 (N_7385,N_6070,N_6659);
nand U7386 (N_7386,N_6001,N_6271);
nor U7387 (N_7387,N_6819,N_6435);
nand U7388 (N_7388,N_6689,N_6016);
xor U7389 (N_7389,N_6172,N_6717);
nand U7390 (N_7390,N_6282,N_6413);
nand U7391 (N_7391,N_6923,N_6417);
and U7392 (N_7392,N_6366,N_6157);
xor U7393 (N_7393,N_6808,N_6120);
nand U7394 (N_7394,N_6975,N_6247);
xnor U7395 (N_7395,N_6513,N_6928);
nor U7396 (N_7396,N_6939,N_6331);
nor U7397 (N_7397,N_6966,N_6647);
nor U7398 (N_7398,N_6046,N_6982);
nor U7399 (N_7399,N_6559,N_6609);
or U7400 (N_7400,N_6236,N_6845);
nor U7401 (N_7401,N_6085,N_6335);
nand U7402 (N_7402,N_6325,N_6233);
and U7403 (N_7403,N_6142,N_6207);
xnor U7404 (N_7404,N_6992,N_6699);
or U7405 (N_7405,N_6204,N_6554);
nand U7406 (N_7406,N_6908,N_6465);
nor U7407 (N_7407,N_6151,N_6550);
or U7408 (N_7408,N_6252,N_6867);
xnor U7409 (N_7409,N_6526,N_6202);
nand U7410 (N_7410,N_6980,N_6225);
nor U7411 (N_7411,N_6321,N_6820);
xnor U7412 (N_7412,N_6071,N_6308);
and U7413 (N_7413,N_6528,N_6430);
nand U7414 (N_7414,N_6750,N_6856);
xnor U7415 (N_7415,N_6033,N_6003);
xor U7416 (N_7416,N_6210,N_6979);
xor U7417 (N_7417,N_6839,N_6713);
or U7418 (N_7418,N_6160,N_6792);
nand U7419 (N_7419,N_6130,N_6783);
nand U7420 (N_7420,N_6628,N_6243);
xnor U7421 (N_7421,N_6835,N_6620);
nor U7422 (N_7422,N_6405,N_6950);
nand U7423 (N_7423,N_6459,N_6445);
and U7424 (N_7424,N_6940,N_6126);
nand U7425 (N_7425,N_6091,N_6393);
and U7426 (N_7426,N_6175,N_6733);
and U7427 (N_7427,N_6864,N_6704);
xor U7428 (N_7428,N_6972,N_6482);
nand U7429 (N_7429,N_6581,N_6315);
nor U7430 (N_7430,N_6915,N_6196);
or U7431 (N_7431,N_6562,N_6334);
xor U7432 (N_7432,N_6457,N_6902);
or U7433 (N_7433,N_6776,N_6876);
xor U7434 (N_7434,N_6780,N_6231);
nor U7435 (N_7435,N_6497,N_6530);
and U7436 (N_7436,N_6174,N_6696);
xnor U7437 (N_7437,N_6627,N_6060);
or U7438 (N_7438,N_6986,N_6176);
and U7439 (N_7439,N_6744,N_6925);
nor U7440 (N_7440,N_6137,N_6267);
nand U7441 (N_7441,N_6274,N_6691);
nand U7442 (N_7442,N_6198,N_6661);
and U7443 (N_7443,N_6563,N_6669);
and U7444 (N_7444,N_6287,N_6211);
or U7445 (N_7445,N_6673,N_6613);
or U7446 (N_7446,N_6758,N_6571);
nor U7447 (N_7447,N_6586,N_6311);
nor U7448 (N_7448,N_6809,N_6410);
xnor U7449 (N_7449,N_6685,N_6293);
nor U7450 (N_7450,N_6368,N_6548);
or U7451 (N_7451,N_6297,N_6598);
nand U7452 (N_7452,N_6296,N_6577);
nor U7453 (N_7453,N_6364,N_6604);
nor U7454 (N_7454,N_6767,N_6019);
or U7455 (N_7455,N_6397,N_6891);
xor U7456 (N_7456,N_6305,N_6092);
nor U7457 (N_7457,N_6021,N_6879);
xor U7458 (N_7458,N_6743,N_6719);
nor U7459 (N_7459,N_6209,N_6900);
nand U7460 (N_7460,N_6217,N_6094);
or U7461 (N_7461,N_6406,N_6191);
and U7462 (N_7462,N_6605,N_6374);
nand U7463 (N_7463,N_6573,N_6988);
or U7464 (N_7464,N_6190,N_6109);
nand U7465 (N_7465,N_6918,N_6133);
nand U7466 (N_7466,N_6400,N_6771);
nor U7467 (N_7467,N_6257,N_6040);
or U7468 (N_7468,N_6849,N_6706);
or U7469 (N_7469,N_6108,N_6865);
or U7470 (N_7470,N_6027,N_6455);
xnor U7471 (N_7471,N_6223,N_6901);
and U7472 (N_7472,N_6064,N_6692);
or U7473 (N_7473,N_6263,N_6745);
xor U7474 (N_7474,N_6011,N_6566);
nand U7475 (N_7475,N_6934,N_6846);
nand U7476 (N_7476,N_6352,N_6504);
nand U7477 (N_7477,N_6473,N_6082);
and U7478 (N_7478,N_6140,N_6816);
nand U7479 (N_7479,N_6034,N_6304);
nor U7480 (N_7480,N_6474,N_6558);
nand U7481 (N_7481,N_6960,N_6438);
or U7482 (N_7482,N_6131,N_6644);
or U7483 (N_7483,N_6149,N_6214);
nand U7484 (N_7484,N_6730,N_6063);
nor U7485 (N_7485,N_6099,N_6449);
nor U7486 (N_7486,N_6686,N_6618);
or U7487 (N_7487,N_6786,N_6301);
nor U7488 (N_7488,N_6298,N_6144);
and U7489 (N_7489,N_6551,N_6775);
xor U7490 (N_7490,N_6320,N_6593);
and U7491 (N_7491,N_6230,N_6453);
nand U7492 (N_7492,N_6903,N_6491);
nor U7493 (N_7493,N_6921,N_6351);
nor U7494 (N_7494,N_6874,N_6086);
xor U7495 (N_7495,N_6227,N_6626);
and U7496 (N_7496,N_6212,N_6886);
nand U7497 (N_7497,N_6195,N_6948);
nor U7498 (N_7498,N_6671,N_6994);
nand U7499 (N_7499,N_6171,N_6279);
nand U7500 (N_7500,N_6842,N_6778);
or U7501 (N_7501,N_6905,N_6507);
and U7502 (N_7502,N_6929,N_6013);
nor U7503 (N_7503,N_6421,N_6397);
and U7504 (N_7504,N_6526,N_6194);
xor U7505 (N_7505,N_6744,N_6879);
nor U7506 (N_7506,N_6000,N_6886);
and U7507 (N_7507,N_6692,N_6176);
xor U7508 (N_7508,N_6944,N_6578);
nor U7509 (N_7509,N_6231,N_6536);
nor U7510 (N_7510,N_6349,N_6243);
xor U7511 (N_7511,N_6530,N_6438);
and U7512 (N_7512,N_6455,N_6932);
and U7513 (N_7513,N_6178,N_6698);
or U7514 (N_7514,N_6856,N_6128);
and U7515 (N_7515,N_6294,N_6767);
or U7516 (N_7516,N_6955,N_6004);
nor U7517 (N_7517,N_6178,N_6125);
nor U7518 (N_7518,N_6213,N_6463);
and U7519 (N_7519,N_6695,N_6104);
xor U7520 (N_7520,N_6504,N_6633);
nor U7521 (N_7521,N_6145,N_6174);
nor U7522 (N_7522,N_6592,N_6257);
and U7523 (N_7523,N_6891,N_6479);
nor U7524 (N_7524,N_6995,N_6050);
nor U7525 (N_7525,N_6441,N_6969);
and U7526 (N_7526,N_6229,N_6669);
or U7527 (N_7527,N_6296,N_6324);
nor U7528 (N_7528,N_6000,N_6893);
nand U7529 (N_7529,N_6046,N_6922);
nor U7530 (N_7530,N_6320,N_6290);
xnor U7531 (N_7531,N_6605,N_6042);
nand U7532 (N_7532,N_6741,N_6151);
xor U7533 (N_7533,N_6546,N_6263);
and U7534 (N_7534,N_6913,N_6574);
nand U7535 (N_7535,N_6088,N_6492);
or U7536 (N_7536,N_6116,N_6471);
nor U7537 (N_7537,N_6944,N_6837);
nand U7538 (N_7538,N_6908,N_6636);
xor U7539 (N_7539,N_6990,N_6873);
and U7540 (N_7540,N_6289,N_6792);
or U7541 (N_7541,N_6560,N_6960);
xnor U7542 (N_7542,N_6805,N_6372);
or U7543 (N_7543,N_6040,N_6601);
nand U7544 (N_7544,N_6581,N_6353);
and U7545 (N_7545,N_6251,N_6360);
or U7546 (N_7546,N_6189,N_6176);
nor U7547 (N_7547,N_6422,N_6712);
xor U7548 (N_7548,N_6994,N_6612);
xor U7549 (N_7549,N_6704,N_6011);
xnor U7550 (N_7550,N_6589,N_6993);
or U7551 (N_7551,N_6409,N_6565);
or U7552 (N_7552,N_6426,N_6514);
nor U7553 (N_7553,N_6423,N_6810);
nor U7554 (N_7554,N_6748,N_6216);
xnor U7555 (N_7555,N_6163,N_6545);
and U7556 (N_7556,N_6705,N_6847);
nor U7557 (N_7557,N_6833,N_6497);
nor U7558 (N_7558,N_6084,N_6701);
and U7559 (N_7559,N_6396,N_6325);
nor U7560 (N_7560,N_6521,N_6730);
or U7561 (N_7561,N_6858,N_6007);
nor U7562 (N_7562,N_6590,N_6057);
nor U7563 (N_7563,N_6193,N_6153);
or U7564 (N_7564,N_6096,N_6057);
nor U7565 (N_7565,N_6134,N_6310);
nand U7566 (N_7566,N_6522,N_6941);
xnor U7567 (N_7567,N_6027,N_6898);
or U7568 (N_7568,N_6857,N_6994);
and U7569 (N_7569,N_6729,N_6206);
and U7570 (N_7570,N_6240,N_6865);
or U7571 (N_7571,N_6267,N_6318);
nor U7572 (N_7572,N_6916,N_6129);
nand U7573 (N_7573,N_6498,N_6695);
and U7574 (N_7574,N_6784,N_6208);
nand U7575 (N_7575,N_6040,N_6263);
or U7576 (N_7576,N_6295,N_6856);
xor U7577 (N_7577,N_6054,N_6797);
and U7578 (N_7578,N_6041,N_6185);
nor U7579 (N_7579,N_6950,N_6144);
and U7580 (N_7580,N_6756,N_6269);
or U7581 (N_7581,N_6897,N_6329);
nand U7582 (N_7582,N_6833,N_6811);
and U7583 (N_7583,N_6398,N_6832);
nor U7584 (N_7584,N_6576,N_6511);
nand U7585 (N_7585,N_6227,N_6144);
nand U7586 (N_7586,N_6479,N_6681);
or U7587 (N_7587,N_6064,N_6632);
and U7588 (N_7588,N_6527,N_6578);
nand U7589 (N_7589,N_6786,N_6251);
and U7590 (N_7590,N_6057,N_6065);
xnor U7591 (N_7591,N_6920,N_6497);
nor U7592 (N_7592,N_6918,N_6760);
xnor U7593 (N_7593,N_6156,N_6022);
and U7594 (N_7594,N_6019,N_6302);
nand U7595 (N_7595,N_6254,N_6102);
nand U7596 (N_7596,N_6762,N_6377);
or U7597 (N_7597,N_6133,N_6856);
or U7598 (N_7598,N_6915,N_6291);
and U7599 (N_7599,N_6243,N_6067);
nand U7600 (N_7600,N_6748,N_6023);
nand U7601 (N_7601,N_6874,N_6041);
or U7602 (N_7602,N_6036,N_6494);
xor U7603 (N_7603,N_6145,N_6543);
or U7604 (N_7604,N_6323,N_6145);
nand U7605 (N_7605,N_6908,N_6064);
or U7606 (N_7606,N_6270,N_6829);
xnor U7607 (N_7607,N_6552,N_6819);
nor U7608 (N_7608,N_6968,N_6632);
and U7609 (N_7609,N_6190,N_6904);
and U7610 (N_7610,N_6330,N_6401);
or U7611 (N_7611,N_6052,N_6860);
xor U7612 (N_7612,N_6509,N_6398);
or U7613 (N_7613,N_6379,N_6783);
and U7614 (N_7614,N_6843,N_6993);
nor U7615 (N_7615,N_6015,N_6921);
and U7616 (N_7616,N_6658,N_6023);
nand U7617 (N_7617,N_6256,N_6501);
nand U7618 (N_7618,N_6574,N_6315);
and U7619 (N_7619,N_6741,N_6054);
xor U7620 (N_7620,N_6762,N_6258);
nand U7621 (N_7621,N_6749,N_6360);
and U7622 (N_7622,N_6526,N_6766);
nor U7623 (N_7623,N_6554,N_6007);
nor U7624 (N_7624,N_6798,N_6019);
nor U7625 (N_7625,N_6156,N_6788);
nor U7626 (N_7626,N_6466,N_6906);
or U7627 (N_7627,N_6619,N_6365);
nand U7628 (N_7628,N_6013,N_6357);
xor U7629 (N_7629,N_6803,N_6432);
xnor U7630 (N_7630,N_6600,N_6252);
nand U7631 (N_7631,N_6525,N_6628);
xor U7632 (N_7632,N_6289,N_6400);
nand U7633 (N_7633,N_6177,N_6694);
xnor U7634 (N_7634,N_6002,N_6770);
nand U7635 (N_7635,N_6233,N_6742);
and U7636 (N_7636,N_6271,N_6065);
or U7637 (N_7637,N_6362,N_6775);
and U7638 (N_7638,N_6899,N_6053);
or U7639 (N_7639,N_6239,N_6921);
xor U7640 (N_7640,N_6564,N_6814);
xnor U7641 (N_7641,N_6489,N_6684);
xor U7642 (N_7642,N_6516,N_6044);
xnor U7643 (N_7643,N_6210,N_6725);
nor U7644 (N_7644,N_6738,N_6609);
nor U7645 (N_7645,N_6900,N_6992);
nor U7646 (N_7646,N_6538,N_6288);
nor U7647 (N_7647,N_6428,N_6665);
nor U7648 (N_7648,N_6712,N_6780);
nand U7649 (N_7649,N_6887,N_6169);
nand U7650 (N_7650,N_6749,N_6287);
and U7651 (N_7651,N_6817,N_6243);
or U7652 (N_7652,N_6339,N_6566);
nand U7653 (N_7653,N_6239,N_6380);
nand U7654 (N_7654,N_6009,N_6583);
xnor U7655 (N_7655,N_6387,N_6928);
or U7656 (N_7656,N_6399,N_6711);
and U7657 (N_7657,N_6625,N_6907);
nand U7658 (N_7658,N_6346,N_6760);
nand U7659 (N_7659,N_6952,N_6745);
nor U7660 (N_7660,N_6351,N_6120);
nor U7661 (N_7661,N_6286,N_6428);
nand U7662 (N_7662,N_6371,N_6217);
nand U7663 (N_7663,N_6913,N_6272);
and U7664 (N_7664,N_6217,N_6333);
xor U7665 (N_7665,N_6428,N_6885);
and U7666 (N_7666,N_6702,N_6085);
nor U7667 (N_7667,N_6120,N_6053);
nor U7668 (N_7668,N_6819,N_6397);
and U7669 (N_7669,N_6820,N_6568);
and U7670 (N_7670,N_6685,N_6404);
nor U7671 (N_7671,N_6504,N_6605);
and U7672 (N_7672,N_6803,N_6731);
xor U7673 (N_7673,N_6422,N_6507);
or U7674 (N_7674,N_6411,N_6835);
and U7675 (N_7675,N_6624,N_6801);
xnor U7676 (N_7676,N_6947,N_6030);
and U7677 (N_7677,N_6854,N_6418);
nor U7678 (N_7678,N_6716,N_6275);
and U7679 (N_7679,N_6314,N_6612);
nand U7680 (N_7680,N_6192,N_6968);
nor U7681 (N_7681,N_6878,N_6805);
nor U7682 (N_7682,N_6662,N_6514);
nand U7683 (N_7683,N_6901,N_6978);
xor U7684 (N_7684,N_6036,N_6334);
and U7685 (N_7685,N_6680,N_6212);
nor U7686 (N_7686,N_6334,N_6431);
nand U7687 (N_7687,N_6492,N_6787);
nand U7688 (N_7688,N_6148,N_6650);
nand U7689 (N_7689,N_6567,N_6238);
or U7690 (N_7690,N_6423,N_6035);
or U7691 (N_7691,N_6351,N_6730);
xnor U7692 (N_7692,N_6051,N_6096);
and U7693 (N_7693,N_6484,N_6001);
xnor U7694 (N_7694,N_6368,N_6874);
and U7695 (N_7695,N_6947,N_6674);
nand U7696 (N_7696,N_6927,N_6040);
xor U7697 (N_7697,N_6922,N_6466);
xor U7698 (N_7698,N_6904,N_6202);
xnor U7699 (N_7699,N_6844,N_6715);
or U7700 (N_7700,N_6346,N_6483);
and U7701 (N_7701,N_6671,N_6117);
nand U7702 (N_7702,N_6305,N_6166);
or U7703 (N_7703,N_6542,N_6630);
and U7704 (N_7704,N_6059,N_6987);
nand U7705 (N_7705,N_6729,N_6470);
xnor U7706 (N_7706,N_6194,N_6636);
and U7707 (N_7707,N_6336,N_6383);
or U7708 (N_7708,N_6508,N_6056);
xnor U7709 (N_7709,N_6683,N_6870);
nor U7710 (N_7710,N_6675,N_6034);
nor U7711 (N_7711,N_6868,N_6535);
xor U7712 (N_7712,N_6959,N_6445);
and U7713 (N_7713,N_6501,N_6165);
nor U7714 (N_7714,N_6493,N_6348);
nand U7715 (N_7715,N_6163,N_6270);
and U7716 (N_7716,N_6822,N_6162);
and U7717 (N_7717,N_6218,N_6311);
xor U7718 (N_7718,N_6596,N_6700);
or U7719 (N_7719,N_6360,N_6399);
nor U7720 (N_7720,N_6428,N_6485);
nand U7721 (N_7721,N_6404,N_6707);
xor U7722 (N_7722,N_6494,N_6842);
or U7723 (N_7723,N_6211,N_6296);
xor U7724 (N_7724,N_6413,N_6077);
or U7725 (N_7725,N_6402,N_6562);
nand U7726 (N_7726,N_6146,N_6170);
nor U7727 (N_7727,N_6704,N_6472);
nor U7728 (N_7728,N_6551,N_6872);
nor U7729 (N_7729,N_6252,N_6180);
xnor U7730 (N_7730,N_6445,N_6931);
or U7731 (N_7731,N_6532,N_6809);
or U7732 (N_7732,N_6614,N_6566);
nand U7733 (N_7733,N_6341,N_6786);
nor U7734 (N_7734,N_6403,N_6168);
and U7735 (N_7735,N_6093,N_6802);
xnor U7736 (N_7736,N_6473,N_6441);
and U7737 (N_7737,N_6990,N_6376);
or U7738 (N_7738,N_6068,N_6417);
and U7739 (N_7739,N_6724,N_6410);
xor U7740 (N_7740,N_6610,N_6991);
nand U7741 (N_7741,N_6802,N_6766);
nand U7742 (N_7742,N_6253,N_6408);
or U7743 (N_7743,N_6673,N_6000);
xnor U7744 (N_7744,N_6955,N_6949);
and U7745 (N_7745,N_6697,N_6618);
and U7746 (N_7746,N_6487,N_6550);
nor U7747 (N_7747,N_6133,N_6531);
xnor U7748 (N_7748,N_6830,N_6827);
nor U7749 (N_7749,N_6987,N_6499);
xor U7750 (N_7750,N_6937,N_6024);
and U7751 (N_7751,N_6588,N_6568);
and U7752 (N_7752,N_6657,N_6340);
nand U7753 (N_7753,N_6784,N_6417);
nand U7754 (N_7754,N_6684,N_6843);
and U7755 (N_7755,N_6405,N_6610);
nand U7756 (N_7756,N_6380,N_6998);
nand U7757 (N_7757,N_6033,N_6465);
and U7758 (N_7758,N_6107,N_6130);
xor U7759 (N_7759,N_6932,N_6195);
nand U7760 (N_7760,N_6412,N_6984);
nor U7761 (N_7761,N_6081,N_6476);
xor U7762 (N_7762,N_6043,N_6468);
and U7763 (N_7763,N_6437,N_6921);
or U7764 (N_7764,N_6018,N_6396);
nand U7765 (N_7765,N_6571,N_6212);
xnor U7766 (N_7766,N_6830,N_6543);
and U7767 (N_7767,N_6312,N_6317);
xnor U7768 (N_7768,N_6944,N_6233);
xnor U7769 (N_7769,N_6835,N_6697);
nand U7770 (N_7770,N_6427,N_6321);
and U7771 (N_7771,N_6958,N_6998);
nor U7772 (N_7772,N_6845,N_6251);
nor U7773 (N_7773,N_6774,N_6603);
xor U7774 (N_7774,N_6543,N_6887);
xnor U7775 (N_7775,N_6030,N_6840);
nand U7776 (N_7776,N_6356,N_6058);
xnor U7777 (N_7777,N_6216,N_6983);
nor U7778 (N_7778,N_6374,N_6858);
or U7779 (N_7779,N_6636,N_6023);
xor U7780 (N_7780,N_6520,N_6421);
and U7781 (N_7781,N_6595,N_6587);
nor U7782 (N_7782,N_6599,N_6536);
and U7783 (N_7783,N_6616,N_6461);
nand U7784 (N_7784,N_6532,N_6206);
and U7785 (N_7785,N_6848,N_6780);
and U7786 (N_7786,N_6831,N_6432);
nand U7787 (N_7787,N_6293,N_6583);
nor U7788 (N_7788,N_6649,N_6540);
nor U7789 (N_7789,N_6717,N_6590);
nor U7790 (N_7790,N_6596,N_6699);
and U7791 (N_7791,N_6749,N_6822);
nand U7792 (N_7792,N_6162,N_6693);
or U7793 (N_7793,N_6041,N_6550);
and U7794 (N_7794,N_6125,N_6901);
nand U7795 (N_7795,N_6915,N_6631);
and U7796 (N_7796,N_6093,N_6699);
nor U7797 (N_7797,N_6070,N_6136);
or U7798 (N_7798,N_6560,N_6928);
nor U7799 (N_7799,N_6104,N_6111);
or U7800 (N_7800,N_6923,N_6623);
or U7801 (N_7801,N_6661,N_6125);
nor U7802 (N_7802,N_6947,N_6371);
xor U7803 (N_7803,N_6987,N_6813);
nor U7804 (N_7804,N_6997,N_6316);
and U7805 (N_7805,N_6109,N_6465);
or U7806 (N_7806,N_6037,N_6459);
nor U7807 (N_7807,N_6705,N_6127);
or U7808 (N_7808,N_6717,N_6014);
nor U7809 (N_7809,N_6852,N_6283);
nand U7810 (N_7810,N_6374,N_6509);
nand U7811 (N_7811,N_6316,N_6017);
or U7812 (N_7812,N_6697,N_6363);
nand U7813 (N_7813,N_6155,N_6335);
nand U7814 (N_7814,N_6220,N_6076);
and U7815 (N_7815,N_6063,N_6855);
nor U7816 (N_7816,N_6314,N_6155);
or U7817 (N_7817,N_6716,N_6033);
nand U7818 (N_7818,N_6843,N_6081);
xnor U7819 (N_7819,N_6644,N_6508);
xor U7820 (N_7820,N_6050,N_6092);
nor U7821 (N_7821,N_6058,N_6915);
nor U7822 (N_7822,N_6722,N_6353);
and U7823 (N_7823,N_6799,N_6617);
and U7824 (N_7824,N_6553,N_6392);
or U7825 (N_7825,N_6135,N_6442);
and U7826 (N_7826,N_6492,N_6699);
and U7827 (N_7827,N_6620,N_6450);
and U7828 (N_7828,N_6337,N_6765);
or U7829 (N_7829,N_6237,N_6869);
or U7830 (N_7830,N_6541,N_6122);
nor U7831 (N_7831,N_6919,N_6791);
nor U7832 (N_7832,N_6019,N_6705);
and U7833 (N_7833,N_6206,N_6136);
nor U7834 (N_7834,N_6516,N_6559);
xor U7835 (N_7835,N_6840,N_6453);
nand U7836 (N_7836,N_6376,N_6331);
nor U7837 (N_7837,N_6369,N_6516);
xnor U7838 (N_7838,N_6103,N_6788);
xor U7839 (N_7839,N_6004,N_6709);
nor U7840 (N_7840,N_6593,N_6636);
nor U7841 (N_7841,N_6311,N_6787);
nor U7842 (N_7842,N_6635,N_6237);
or U7843 (N_7843,N_6420,N_6215);
nand U7844 (N_7844,N_6091,N_6120);
nor U7845 (N_7845,N_6565,N_6150);
nor U7846 (N_7846,N_6157,N_6806);
nand U7847 (N_7847,N_6133,N_6767);
or U7848 (N_7848,N_6796,N_6294);
nor U7849 (N_7849,N_6872,N_6768);
nor U7850 (N_7850,N_6553,N_6251);
nand U7851 (N_7851,N_6352,N_6633);
and U7852 (N_7852,N_6713,N_6239);
xor U7853 (N_7853,N_6953,N_6825);
and U7854 (N_7854,N_6869,N_6969);
and U7855 (N_7855,N_6581,N_6736);
or U7856 (N_7856,N_6832,N_6383);
nand U7857 (N_7857,N_6316,N_6444);
or U7858 (N_7858,N_6396,N_6766);
nand U7859 (N_7859,N_6447,N_6162);
xor U7860 (N_7860,N_6274,N_6710);
xor U7861 (N_7861,N_6202,N_6529);
nand U7862 (N_7862,N_6295,N_6888);
nor U7863 (N_7863,N_6683,N_6145);
nand U7864 (N_7864,N_6677,N_6091);
or U7865 (N_7865,N_6148,N_6659);
or U7866 (N_7866,N_6661,N_6585);
xor U7867 (N_7867,N_6232,N_6814);
or U7868 (N_7868,N_6557,N_6570);
nor U7869 (N_7869,N_6683,N_6163);
nor U7870 (N_7870,N_6597,N_6275);
nor U7871 (N_7871,N_6826,N_6472);
xnor U7872 (N_7872,N_6929,N_6792);
xor U7873 (N_7873,N_6218,N_6593);
nor U7874 (N_7874,N_6391,N_6399);
or U7875 (N_7875,N_6968,N_6442);
and U7876 (N_7876,N_6399,N_6803);
xor U7877 (N_7877,N_6751,N_6616);
xor U7878 (N_7878,N_6406,N_6959);
and U7879 (N_7879,N_6405,N_6231);
or U7880 (N_7880,N_6653,N_6954);
xor U7881 (N_7881,N_6188,N_6114);
nor U7882 (N_7882,N_6427,N_6667);
nand U7883 (N_7883,N_6593,N_6621);
nor U7884 (N_7884,N_6573,N_6863);
nor U7885 (N_7885,N_6929,N_6949);
and U7886 (N_7886,N_6086,N_6051);
or U7887 (N_7887,N_6898,N_6666);
or U7888 (N_7888,N_6714,N_6585);
or U7889 (N_7889,N_6173,N_6098);
xnor U7890 (N_7890,N_6461,N_6712);
xor U7891 (N_7891,N_6134,N_6403);
and U7892 (N_7892,N_6052,N_6977);
and U7893 (N_7893,N_6933,N_6588);
nor U7894 (N_7894,N_6405,N_6521);
xor U7895 (N_7895,N_6238,N_6030);
nand U7896 (N_7896,N_6017,N_6988);
and U7897 (N_7897,N_6538,N_6910);
xnor U7898 (N_7898,N_6105,N_6292);
and U7899 (N_7899,N_6598,N_6634);
and U7900 (N_7900,N_6018,N_6567);
xnor U7901 (N_7901,N_6424,N_6645);
xor U7902 (N_7902,N_6466,N_6687);
nand U7903 (N_7903,N_6580,N_6521);
nor U7904 (N_7904,N_6919,N_6777);
or U7905 (N_7905,N_6470,N_6518);
xor U7906 (N_7906,N_6444,N_6735);
nor U7907 (N_7907,N_6499,N_6288);
or U7908 (N_7908,N_6869,N_6831);
and U7909 (N_7909,N_6231,N_6560);
xor U7910 (N_7910,N_6045,N_6838);
nor U7911 (N_7911,N_6666,N_6347);
and U7912 (N_7912,N_6448,N_6895);
and U7913 (N_7913,N_6872,N_6823);
xor U7914 (N_7914,N_6048,N_6080);
xor U7915 (N_7915,N_6003,N_6171);
nand U7916 (N_7916,N_6670,N_6969);
and U7917 (N_7917,N_6840,N_6827);
nor U7918 (N_7918,N_6613,N_6284);
nor U7919 (N_7919,N_6797,N_6462);
xor U7920 (N_7920,N_6762,N_6254);
nand U7921 (N_7921,N_6101,N_6407);
xor U7922 (N_7922,N_6173,N_6276);
nand U7923 (N_7923,N_6586,N_6680);
nand U7924 (N_7924,N_6920,N_6266);
nor U7925 (N_7925,N_6213,N_6215);
nor U7926 (N_7926,N_6445,N_6587);
nand U7927 (N_7927,N_6216,N_6238);
nor U7928 (N_7928,N_6167,N_6464);
nor U7929 (N_7929,N_6728,N_6028);
and U7930 (N_7930,N_6142,N_6185);
xor U7931 (N_7931,N_6125,N_6911);
nand U7932 (N_7932,N_6398,N_6165);
xnor U7933 (N_7933,N_6500,N_6536);
and U7934 (N_7934,N_6121,N_6565);
xor U7935 (N_7935,N_6675,N_6921);
xnor U7936 (N_7936,N_6262,N_6381);
and U7937 (N_7937,N_6762,N_6787);
or U7938 (N_7938,N_6018,N_6629);
and U7939 (N_7939,N_6968,N_6068);
nand U7940 (N_7940,N_6186,N_6559);
and U7941 (N_7941,N_6086,N_6301);
or U7942 (N_7942,N_6263,N_6728);
nor U7943 (N_7943,N_6595,N_6017);
and U7944 (N_7944,N_6051,N_6625);
nor U7945 (N_7945,N_6529,N_6125);
nand U7946 (N_7946,N_6630,N_6789);
and U7947 (N_7947,N_6259,N_6949);
and U7948 (N_7948,N_6517,N_6243);
xnor U7949 (N_7949,N_6134,N_6007);
or U7950 (N_7950,N_6075,N_6497);
xor U7951 (N_7951,N_6829,N_6885);
nand U7952 (N_7952,N_6595,N_6657);
nand U7953 (N_7953,N_6557,N_6437);
or U7954 (N_7954,N_6717,N_6350);
nand U7955 (N_7955,N_6692,N_6694);
or U7956 (N_7956,N_6571,N_6960);
or U7957 (N_7957,N_6147,N_6640);
xnor U7958 (N_7958,N_6066,N_6987);
and U7959 (N_7959,N_6667,N_6371);
or U7960 (N_7960,N_6488,N_6589);
nand U7961 (N_7961,N_6526,N_6003);
nand U7962 (N_7962,N_6584,N_6325);
or U7963 (N_7963,N_6979,N_6294);
and U7964 (N_7964,N_6091,N_6568);
nor U7965 (N_7965,N_6253,N_6708);
or U7966 (N_7966,N_6279,N_6834);
xnor U7967 (N_7967,N_6863,N_6858);
and U7968 (N_7968,N_6533,N_6725);
nand U7969 (N_7969,N_6821,N_6104);
and U7970 (N_7970,N_6302,N_6580);
xor U7971 (N_7971,N_6039,N_6348);
nand U7972 (N_7972,N_6797,N_6983);
nor U7973 (N_7973,N_6409,N_6220);
or U7974 (N_7974,N_6687,N_6292);
xor U7975 (N_7975,N_6147,N_6218);
xnor U7976 (N_7976,N_6692,N_6431);
xnor U7977 (N_7977,N_6953,N_6994);
xor U7978 (N_7978,N_6456,N_6405);
nor U7979 (N_7979,N_6186,N_6078);
xor U7980 (N_7980,N_6284,N_6877);
and U7981 (N_7981,N_6158,N_6297);
xor U7982 (N_7982,N_6326,N_6101);
and U7983 (N_7983,N_6108,N_6641);
xor U7984 (N_7984,N_6141,N_6999);
nand U7985 (N_7985,N_6865,N_6522);
xor U7986 (N_7986,N_6171,N_6688);
or U7987 (N_7987,N_6696,N_6656);
nand U7988 (N_7988,N_6555,N_6084);
and U7989 (N_7989,N_6588,N_6349);
nand U7990 (N_7990,N_6494,N_6845);
nor U7991 (N_7991,N_6093,N_6026);
nand U7992 (N_7992,N_6922,N_6425);
nand U7993 (N_7993,N_6356,N_6691);
nand U7994 (N_7994,N_6495,N_6416);
and U7995 (N_7995,N_6395,N_6696);
and U7996 (N_7996,N_6474,N_6531);
nand U7997 (N_7997,N_6306,N_6566);
nand U7998 (N_7998,N_6398,N_6991);
and U7999 (N_7999,N_6580,N_6624);
nand U8000 (N_8000,N_7467,N_7523);
nor U8001 (N_8001,N_7706,N_7740);
nor U8002 (N_8002,N_7159,N_7533);
nor U8003 (N_8003,N_7911,N_7526);
xor U8004 (N_8004,N_7953,N_7046);
xor U8005 (N_8005,N_7906,N_7466);
xor U8006 (N_8006,N_7468,N_7516);
or U8007 (N_8007,N_7388,N_7960);
nor U8008 (N_8008,N_7107,N_7549);
xor U8009 (N_8009,N_7835,N_7202);
or U8010 (N_8010,N_7044,N_7238);
and U8011 (N_8011,N_7180,N_7934);
nor U8012 (N_8012,N_7479,N_7597);
and U8013 (N_8013,N_7700,N_7945);
xnor U8014 (N_8014,N_7478,N_7949);
xor U8015 (N_8015,N_7299,N_7635);
nor U8016 (N_8016,N_7722,N_7903);
and U8017 (N_8017,N_7900,N_7561);
nand U8018 (N_8018,N_7755,N_7551);
and U8019 (N_8019,N_7333,N_7752);
nand U8020 (N_8020,N_7637,N_7422);
nor U8021 (N_8021,N_7131,N_7286);
nor U8022 (N_8022,N_7718,N_7730);
nor U8023 (N_8023,N_7449,N_7263);
nor U8024 (N_8024,N_7772,N_7611);
xnor U8025 (N_8025,N_7552,N_7653);
or U8026 (N_8026,N_7307,N_7062);
or U8027 (N_8027,N_7398,N_7465);
or U8028 (N_8028,N_7072,N_7432);
nor U8029 (N_8029,N_7066,N_7117);
or U8030 (N_8030,N_7091,N_7486);
or U8031 (N_8031,N_7330,N_7183);
nand U8032 (N_8032,N_7578,N_7227);
and U8033 (N_8033,N_7579,N_7636);
nand U8034 (N_8034,N_7827,N_7356);
and U8035 (N_8035,N_7562,N_7677);
xnor U8036 (N_8036,N_7296,N_7801);
and U8037 (N_8037,N_7712,N_7867);
nor U8038 (N_8038,N_7645,N_7147);
or U8039 (N_8039,N_7993,N_7111);
and U8040 (N_8040,N_7010,N_7918);
and U8041 (N_8041,N_7493,N_7018);
nand U8042 (N_8042,N_7361,N_7698);
xnor U8043 (N_8043,N_7992,N_7774);
nand U8044 (N_8044,N_7097,N_7223);
nor U8045 (N_8045,N_7986,N_7259);
nand U8046 (N_8046,N_7825,N_7198);
nor U8047 (N_8047,N_7373,N_7112);
xor U8048 (N_8048,N_7309,N_7882);
and U8049 (N_8049,N_7028,N_7914);
nand U8050 (N_8050,N_7065,N_7424);
xnor U8051 (N_8051,N_7406,N_7931);
and U8052 (N_8052,N_7411,N_7646);
or U8053 (N_8053,N_7823,N_7342);
xor U8054 (N_8054,N_7474,N_7485);
or U8055 (N_8055,N_7345,N_7690);
xor U8056 (N_8056,N_7142,N_7996);
xor U8057 (N_8057,N_7125,N_7812);
nand U8058 (N_8058,N_7442,N_7007);
or U8059 (N_8059,N_7988,N_7761);
nor U8060 (N_8060,N_7572,N_7133);
xnor U8061 (N_8061,N_7505,N_7499);
or U8062 (N_8062,N_7366,N_7948);
and U8063 (N_8063,N_7257,N_7058);
nor U8064 (N_8064,N_7412,N_7494);
and U8065 (N_8065,N_7826,N_7910);
xor U8066 (N_8066,N_7195,N_7703);
and U8067 (N_8067,N_7976,N_7045);
xnor U8068 (N_8068,N_7952,N_7023);
nand U8069 (N_8069,N_7689,N_7215);
xnor U8070 (N_8070,N_7311,N_7222);
nor U8071 (N_8071,N_7460,N_7547);
and U8072 (N_8072,N_7425,N_7317);
or U8073 (N_8073,N_7355,N_7252);
or U8074 (N_8074,N_7265,N_7660);
nor U8075 (N_8075,N_7270,N_7435);
xor U8076 (N_8076,N_7266,N_7418);
nand U8077 (N_8077,N_7304,N_7370);
or U8078 (N_8078,N_7335,N_7121);
nor U8079 (N_8079,N_7648,N_7248);
and U8080 (N_8080,N_7544,N_7186);
nor U8081 (N_8081,N_7780,N_7742);
nor U8082 (N_8082,N_7741,N_7613);
nand U8083 (N_8083,N_7413,N_7497);
nor U8084 (N_8084,N_7175,N_7316);
nor U8085 (N_8085,N_7380,N_7577);
or U8086 (N_8086,N_7455,N_7429);
or U8087 (N_8087,N_7723,N_7278);
nor U8088 (N_8088,N_7093,N_7786);
nand U8089 (N_8089,N_7545,N_7255);
nand U8090 (N_8090,N_7433,N_7899);
nand U8091 (N_8091,N_7981,N_7804);
or U8092 (N_8092,N_7924,N_7284);
and U8093 (N_8093,N_7445,N_7793);
or U8094 (N_8094,N_7405,N_7515);
nor U8095 (N_8095,N_7922,N_7151);
and U8096 (N_8096,N_7353,N_7037);
or U8097 (N_8097,N_7947,N_7123);
nor U8098 (N_8098,N_7575,N_7365);
nor U8099 (N_8099,N_7074,N_7941);
or U8100 (N_8100,N_7052,N_7502);
nor U8101 (N_8101,N_7347,N_7077);
or U8102 (N_8102,N_7387,N_7165);
xor U8103 (N_8103,N_7861,N_7145);
nor U8104 (N_8104,N_7008,N_7878);
and U8105 (N_8105,N_7488,N_7068);
xnor U8106 (N_8106,N_7319,N_7492);
and U8107 (N_8107,N_7115,N_7854);
nand U8108 (N_8108,N_7399,N_7908);
nand U8109 (N_8109,N_7944,N_7003);
nor U8110 (N_8110,N_7546,N_7883);
or U8111 (N_8111,N_7113,N_7118);
xor U8112 (N_8112,N_7629,N_7616);
xor U8113 (N_8113,N_7391,N_7663);
nand U8114 (N_8114,N_7927,N_7079);
and U8115 (N_8115,N_7343,N_7846);
or U8116 (N_8116,N_7171,N_7651);
nand U8117 (N_8117,N_7098,N_7625);
or U8118 (N_8118,N_7315,N_7739);
nor U8119 (N_8119,N_7452,N_7354);
xor U8120 (N_8120,N_7961,N_7759);
and U8121 (N_8121,N_7288,N_7456);
or U8122 (N_8122,N_7129,N_7916);
or U8123 (N_8123,N_7135,N_7276);
and U8124 (N_8124,N_7674,N_7331);
and U8125 (N_8125,N_7682,N_7457);
xnor U8126 (N_8126,N_7870,N_7866);
nand U8127 (N_8127,N_7326,N_7576);
nand U8128 (N_8128,N_7753,N_7102);
nand U8129 (N_8129,N_7570,N_7235);
nand U8130 (N_8130,N_7737,N_7029);
nand U8131 (N_8131,N_7959,N_7713);
nand U8132 (N_8132,N_7390,N_7153);
and U8133 (N_8133,N_7231,N_7845);
xnor U8134 (N_8134,N_7218,N_7249);
xor U8135 (N_8135,N_7024,N_7427);
xnor U8136 (N_8136,N_7087,N_7940);
nand U8137 (N_8137,N_7053,N_7528);
nand U8138 (N_8138,N_7512,N_7314);
or U8139 (N_8139,N_7586,N_7704);
nand U8140 (N_8140,N_7969,N_7778);
xor U8141 (N_8141,N_7691,N_7621);
xnor U8142 (N_8142,N_7628,N_7438);
and U8143 (N_8143,N_7164,N_7243);
nand U8144 (N_8144,N_7876,N_7287);
nand U8145 (N_8145,N_7749,N_7396);
xor U8146 (N_8146,N_7915,N_7104);
xnor U8147 (N_8147,N_7401,N_7925);
nand U8148 (N_8148,N_7791,N_7094);
nand U8149 (N_8149,N_7206,N_7514);
or U8150 (N_8150,N_7828,N_7187);
xor U8151 (N_8151,N_7081,N_7001);
or U8152 (N_8152,N_7088,N_7855);
xor U8153 (N_8153,N_7064,N_7211);
xor U8154 (N_8154,N_7587,N_7824);
or U8155 (N_8155,N_7033,N_7178);
and U8156 (N_8156,N_7327,N_7728);
and U8157 (N_8157,N_7513,N_7848);
and U8158 (N_8158,N_7417,N_7606);
xnor U8159 (N_8159,N_7527,N_7693);
or U8160 (N_8160,N_7601,N_7734);
and U8161 (N_8161,N_7143,N_7303);
or U8162 (N_8162,N_7559,N_7108);
or U8163 (N_8163,N_7384,N_7638);
nand U8164 (N_8164,N_7950,N_7219);
xnor U8165 (N_8165,N_7995,N_7509);
nand U8166 (N_8166,N_7639,N_7926);
nor U8167 (N_8167,N_7262,N_7736);
nand U8168 (N_8168,N_7776,N_7285);
nor U8169 (N_8169,N_7536,N_7367);
nand U8170 (N_8170,N_7853,N_7894);
nor U8171 (N_8171,N_7834,N_7051);
or U8172 (N_8172,N_7710,N_7913);
or U8173 (N_8173,N_7884,N_7610);
xor U8174 (N_8174,N_7225,N_7763);
nand U8175 (N_8175,N_7671,N_7893);
or U8176 (N_8176,N_7747,N_7240);
and U8177 (N_8177,N_7122,N_7358);
or U8178 (N_8178,N_7082,N_7936);
and U8179 (N_8179,N_7128,N_7731);
or U8180 (N_8180,N_7043,N_7530);
xnor U8181 (N_8181,N_7328,N_7807);
or U8182 (N_8182,N_7683,N_7933);
or U8183 (N_8183,N_7658,N_7477);
and U8184 (N_8184,N_7084,N_7009);
xor U8185 (N_8185,N_7283,N_7932);
nor U8186 (N_8186,N_7800,N_7463);
nor U8187 (N_8187,N_7811,N_7817);
and U8188 (N_8188,N_7100,N_7055);
or U8189 (N_8189,N_7298,N_7831);
nor U8190 (N_8190,N_7869,N_7372);
and U8191 (N_8191,N_7224,N_7972);
nor U8192 (N_8192,N_7127,N_7034);
nand U8193 (N_8193,N_7738,N_7312);
and U8194 (N_8194,N_7404,N_7371);
xnor U8195 (N_8195,N_7631,N_7140);
nand U8196 (N_8196,N_7822,N_7144);
or U8197 (N_8197,N_7684,N_7888);
xnor U8198 (N_8198,N_7318,N_7428);
xor U8199 (N_8199,N_7350,N_7167);
or U8200 (N_8200,N_7771,N_7843);
and U8201 (N_8201,N_7919,N_7116);
xnor U8202 (N_8202,N_7538,N_7818);
or U8203 (N_8203,N_7274,N_7061);
xor U8204 (N_8204,N_7005,N_7419);
or U8205 (N_8205,N_7701,N_7634);
xnor U8206 (N_8206,N_7157,N_7733);
nor U8207 (N_8207,N_7607,N_7955);
nor U8208 (N_8208,N_7229,N_7099);
xor U8209 (N_8209,N_7168,N_7139);
nand U8210 (N_8210,N_7602,N_7381);
xnor U8211 (N_8211,N_7820,N_7132);
and U8212 (N_8212,N_7176,N_7770);
nor U8213 (N_8213,N_7439,N_7471);
and U8214 (N_8214,N_7756,N_7724);
nand U8215 (N_8215,N_7078,N_7650);
and U8216 (N_8216,N_7806,N_7850);
xor U8217 (N_8217,N_7320,N_7633);
nor U8218 (N_8218,N_7324,N_7434);
or U8219 (N_8219,N_7357,N_7500);
xor U8220 (N_8220,N_7310,N_7415);
xnor U8221 (N_8221,N_7160,N_7967);
and U8222 (N_8222,N_7185,N_7214);
and U8223 (N_8223,N_7872,N_7483);
xor U8224 (N_8224,N_7994,N_7885);
nor U8225 (N_8225,N_7448,N_7155);
xor U8226 (N_8226,N_7630,N_7879);
nor U8227 (N_8227,N_7194,N_7119);
xnor U8228 (N_8228,N_7340,N_7805);
or U8229 (N_8229,N_7745,N_7177);
nand U8230 (N_8230,N_7397,N_7569);
nor U8231 (N_8231,N_7138,N_7833);
nand U8232 (N_8232,N_7768,N_7858);
and U8233 (N_8233,N_7059,N_7360);
and U8234 (N_8234,N_7473,N_7989);
nand U8235 (N_8235,N_7203,N_7379);
xnor U8236 (N_8236,N_7930,N_7481);
xor U8237 (N_8237,N_7664,N_7661);
nor U8238 (N_8238,N_7622,N_7676);
xor U8239 (N_8239,N_7518,N_7431);
xnor U8240 (N_8240,N_7212,N_7732);
and U8241 (N_8241,N_7532,N_7714);
nor U8242 (N_8242,N_7294,N_7726);
and U8243 (N_8243,N_7902,N_7236);
xor U8244 (N_8244,N_7244,N_7459);
or U8245 (N_8245,N_7556,N_7260);
nor U8246 (N_8246,N_7120,N_7694);
or U8247 (N_8247,N_7443,N_7548);
nor U8248 (N_8248,N_7781,N_7348);
nand U8249 (N_8249,N_7070,N_7839);
nor U8250 (N_8250,N_7596,N_7654);
or U8251 (N_8251,N_7725,N_7624);
nand U8252 (N_8252,N_7234,N_7169);
xor U8253 (N_8253,N_7246,N_7554);
nand U8254 (N_8254,N_7782,N_7983);
nand U8255 (N_8255,N_7182,N_7537);
xnor U8256 (N_8256,N_7297,N_7997);
xnor U8257 (N_8257,N_7166,N_7662);
nand U8258 (N_8258,N_7400,N_7057);
nor U8259 (N_8259,N_7374,N_7787);
xor U8260 (N_8260,N_7364,N_7641);
nor U8261 (N_8261,N_7395,N_7280);
nor U8262 (N_8262,N_7598,N_7179);
nor U8263 (N_8263,N_7308,N_7541);
and U8264 (N_8264,N_7134,N_7040);
or U8265 (N_8265,N_7475,N_7668);
xnor U8266 (N_8266,N_7892,N_7574);
and U8267 (N_8267,N_7498,N_7810);
nand U8268 (N_8268,N_7764,N_7543);
or U8269 (N_8269,N_7232,N_7982);
and U8270 (N_8270,N_7069,N_7519);
nand U8271 (N_8271,N_7582,N_7279);
or U8272 (N_8272,N_7838,N_7815);
xnor U8273 (N_8273,N_7382,N_7670);
xnor U8274 (N_8274,N_7106,N_7482);
or U8275 (N_8275,N_7090,N_7349);
or U8276 (N_8276,N_7436,N_7321);
xor U8277 (N_8277,N_7016,N_7220);
or U8278 (N_8278,N_7665,N_7496);
or U8279 (N_8279,N_7808,N_7025);
and U8280 (N_8280,N_7453,N_7089);
nand U8281 (N_8281,N_7464,N_7440);
and U8282 (N_8282,N_7409,N_7256);
xor U8283 (N_8283,N_7623,N_7487);
and U8284 (N_8284,N_7666,N_7985);
or U8285 (N_8285,N_7696,N_7020);
xor U8286 (N_8286,N_7991,N_7857);
and U8287 (N_8287,N_7004,N_7291);
nor U8288 (N_8288,N_7375,N_7130);
nor U8289 (N_8289,N_7977,N_7385);
and U8290 (N_8290,N_7735,N_7697);
or U8291 (N_8291,N_7889,N_7184);
and U8292 (N_8292,N_7096,N_7531);
nand U8293 (N_8293,N_7612,N_7282);
nor U8294 (N_8294,N_7154,N_7011);
or U8295 (N_8295,N_7686,N_7788);
nor U8296 (N_8296,N_7501,N_7103);
nand U8297 (N_8297,N_7300,N_7821);
and U8298 (N_8298,N_7871,N_7192);
and U8299 (N_8299,N_7026,N_7588);
or U8300 (N_8300,N_7978,N_7362);
or U8301 (N_8301,N_7716,N_7659);
xor U8302 (N_8302,N_7715,N_7000);
xnor U8303 (N_8303,N_7346,N_7408);
nor U8304 (N_8304,N_7868,N_7794);
nand U8305 (N_8305,N_7403,N_7603);
or U8306 (N_8306,N_7273,N_7864);
and U8307 (N_8307,N_7942,N_7264);
or U8308 (N_8308,N_7840,N_7619);
nand U8309 (N_8309,N_7987,N_7880);
and U8310 (N_8310,N_7565,N_7454);
nor U8311 (N_8311,N_7517,N_7964);
and U8312 (N_8312,N_7150,N_7799);
xnor U8313 (N_8313,N_7054,N_7797);
or U8314 (N_8314,N_7954,N_7047);
xor U8315 (N_8315,N_7975,N_7002);
xor U8316 (N_8316,N_7490,N_7775);
xor U8317 (N_8317,N_7557,N_7522);
or U8318 (N_8318,N_7829,N_7277);
xor U8319 (N_8319,N_7874,N_7325);
nor U8320 (N_8320,N_7275,N_7237);
xnor U8321 (N_8321,N_7110,N_7251);
nand U8322 (N_8322,N_7743,N_7642);
nor U8323 (N_8323,N_7393,N_7525);
or U8324 (N_8324,N_7226,N_7784);
and U8325 (N_8325,N_7905,N_7216);
nand U8326 (N_8326,N_7254,N_7369);
nor U8327 (N_8327,N_7126,N_7250);
and U8328 (N_8328,N_7489,N_7149);
xnor U8329 (N_8329,N_7796,N_7935);
and U8330 (N_8330,N_7592,N_7594);
xor U8331 (N_8331,N_7377,N_7394);
xor U8332 (N_8332,N_7017,N_7208);
xnor U8333 (N_8333,N_7627,N_7476);
or U8334 (N_8334,N_7245,N_7553);
or U8335 (N_8335,N_7137,N_7708);
nand U8336 (N_8336,N_7887,N_7261);
xnor U8337 (N_8337,N_7550,N_7757);
xor U8338 (N_8338,N_7392,N_7205);
and U8339 (N_8339,N_7970,N_7890);
nor U8340 (N_8340,N_7067,N_7909);
or U8341 (N_8341,N_7063,N_7022);
and U8342 (N_8342,N_7920,N_7626);
nand U8343 (N_8343,N_7162,N_7599);
nand U8344 (N_8344,N_7241,N_7535);
or U8345 (N_8345,N_7785,N_7152);
or U8346 (N_8346,N_7938,N_7649);
xnor U8347 (N_8347,N_7253,N_7030);
or U8348 (N_8348,N_7056,N_7719);
and U8349 (N_8349,N_7711,N_7746);
xor U8350 (N_8350,N_7289,N_7109);
nor U8351 (N_8351,N_7727,N_7495);
and U8352 (N_8352,N_7458,N_7558);
xnor U8353 (N_8353,N_7114,N_7075);
xnor U8354 (N_8354,N_7792,N_7667);
or U8355 (N_8355,N_7656,N_7809);
nor U8356 (N_8356,N_7760,N_7181);
or U8357 (N_8357,N_7032,N_7695);
xor U8358 (N_8358,N_7966,N_7269);
or U8359 (N_8359,N_7600,N_7041);
and U8360 (N_8360,N_7563,N_7378);
or U8361 (N_8361,N_7595,N_7917);
or U8362 (N_8362,N_7873,N_7580);
nand U8363 (N_8363,N_7414,N_7086);
nand U8364 (N_8364,N_7451,N_7534);
or U8365 (N_8365,N_7707,N_7036);
xnor U8366 (N_8366,N_7640,N_7865);
and U8367 (N_8367,N_7213,N_7337);
or U8368 (N_8368,N_7407,N_7441);
and U8369 (N_8369,N_7672,N_7402);
nand U8370 (N_8370,N_7984,N_7416);
and U8371 (N_8371,N_7221,N_7830);
and U8372 (N_8372,N_7015,N_7907);
nor U8373 (N_8373,N_7173,N_7302);
nand U8374 (N_8374,N_7589,N_7779);
or U8375 (N_8375,N_7389,N_7951);
or U8376 (N_8376,N_7073,N_7912);
nand U8377 (N_8377,N_7124,N_7583);
nor U8378 (N_8378,N_7188,N_7762);
or U8379 (N_8379,N_7946,N_7963);
and U8380 (N_8380,N_7470,N_7146);
nor U8381 (N_8381,N_7161,N_7555);
and U8382 (N_8382,N_7156,N_7567);
xnor U8383 (N_8383,N_7614,N_7590);
or U8384 (N_8384,N_7744,N_7692);
xnor U8385 (N_8385,N_7189,N_7267);
nand U8386 (N_8386,N_7585,N_7242);
and U8387 (N_8387,N_7469,N_7174);
xor U8388 (N_8388,N_7617,N_7895);
xnor U8389 (N_8389,N_7201,N_7904);
and U8390 (N_8390,N_7573,N_7293);
xnor U8391 (N_8391,N_7301,N_7647);
nor U8392 (N_8392,N_7191,N_7856);
nor U8393 (N_8393,N_7632,N_7480);
nand U8394 (N_8394,N_7542,N_7038);
nand U8395 (N_8395,N_7620,N_7998);
and U8396 (N_8396,N_7844,N_7420);
xor U8397 (N_8397,N_7450,N_7957);
and U8398 (N_8398,N_7842,N_7973);
and U8399 (N_8399,N_7679,N_7790);
nor U8400 (N_8400,N_7281,N_7462);
nor U8401 (N_8401,N_7593,N_7604);
nor U8402 (N_8402,N_7341,N_7581);
and U8403 (N_8403,N_7897,N_7847);
xnor U8404 (N_8404,N_7272,N_7875);
xnor U8405 (N_8405,N_7886,N_7092);
xor U8406 (N_8406,N_7507,N_7750);
nor U8407 (N_8407,N_7437,N_7196);
nor U8408 (N_8408,N_7789,N_7506);
nand U8409 (N_8409,N_7083,N_7021);
or U8410 (N_8410,N_7271,N_7410);
and U8411 (N_8411,N_7295,N_7510);
nor U8412 (N_8412,N_7200,N_7748);
nor U8413 (N_8413,N_7031,N_7014);
nor U8414 (N_8414,N_7929,N_7773);
or U8415 (N_8415,N_7681,N_7209);
and U8416 (N_8416,N_7339,N_7896);
xnor U8417 (N_8417,N_7049,N_7539);
and U8418 (N_8418,N_7521,N_7334);
xnor U8419 (N_8419,N_7344,N_7172);
and U8420 (N_8420,N_7207,N_7447);
and U8421 (N_8421,N_7491,N_7305);
nor U8422 (N_8422,N_7901,N_7136);
nor U8423 (N_8423,N_7338,N_7444);
and U8424 (N_8424,N_7819,N_7657);
and U8425 (N_8425,N_7571,N_7190);
nor U8426 (N_8426,N_7841,N_7193);
nor U8427 (N_8427,N_7609,N_7247);
nand U8428 (N_8428,N_7859,N_7352);
nand U8429 (N_8429,N_7322,N_7877);
nand U8430 (N_8430,N_7956,N_7816);
nand U8431 (N_8431,N_7644,N_7678);
xnor U8432 (N_8432,N_7958,N_7979);
xor U8433 (N_8433,N_7085,N_7717);
or U8434 (N_8434,N_7446,N_7702);
or U8435 (N_8435,N_7540,N_7720);
nor U8436 (N_8436,N_7584,N_7363);
or U8437 (N_8437,N_7217,N_7329);
and U8438 (N_8438,N_7990,N_7351);
xor U8439 (N_8439,N_7891,N_7685);
and U8440 (N_8440,N_7675,N_7832);
nand U8441 (N_8441,N_7655,N_7268);
or U8442 (N_8442,N_7503,N_7836);
and U8443 (N_8443,N_7560,N_7921);
and U8444 (N_8444,N_7766,N_7430);
xor U8445 (N_8445,N_7204,N_7862);
xor U8446 (N_8446,N_7042,N_7669);
or U8447 (N_8447,N_7802,N_7013);
nand U8448 (N_8448,N_7060,N_7968);
xnor U8449 (N_8449,N_7368,N_7292);
and U8450 (N_8450,N_7306,N_7980);
or U8451 (N_8451,N_7939,N_7006);
nand U8452 (N_8452,N_7508,N_7965);
or U8453 (N_8453,N_7798,N_7472);
nor U8454 (N_8454,N_7524,N_7699);
or U8455 (N_8455,N_7751,N_7426);
and U8456 (N_8456,N_7199,N_7048);
or U8457 (N_8457,N_7758,N_7837);
nor U8458 (N_8458,N_7504,N_7050);
and U8459 (N_8459,N_7962,N_7148);
and U8460 (N_8460,N_7233,N_7313);
and U8461 (N_8461,N_7386,N_7795);
or U8462 (N_8462,N_7258,N_7928);
or U8463 (N_8463,N_7566,N_7643);
nor U8464 (N_8464,N_7336,N_7769);
and U8465 (N_8465,N_7852,N_7814);
xnor U8466 (N_8466,N_7511,N_7680);
or U8467 (N_8467,N_7618,N_7608);
or U8468 (N_8468,N_7461,N_7076);
xnor U8469 (N_8469,N_7359,N_7019);
xnor U8470 (N_8470,N_7851,N_7777);
and U8471 (N_8471,N_7898,N_7813);
xor U8472 (N_8472,N_7383,N_7721);
nor U8473 (N_8473,N_7323,N_7615);
and U8474 (N_8474,N_7376,N_7923);
nor U8475 (N_8475,N_7228,N_7673);
nor U8476 (N_8476,N_7095,N_7197);
nand U8477 (N_8477,N_7709,N_7688);
nor U8478 (N_8478,N_7101,N_7754);
and U8479 (N_8479,N_7765,N_7332);
nor U8480 (N_8480,N_7937,N_7210);
nand U8481 (N_8481,N_7999,N_7605);
nor U8482 (N_8482,N_7729,N_7974);
and U8483 (N_8483,N_7783,N_7012);
or U8484 (N_8484,N_7141,N_7105);
or U8485 (N_8485,N_7035,N_7230);
or U8486 (N_8486,N_7568,N_7529);
and U8487 (N_8487,N_7849,N_7170);
nand U8488 (N_8488,N_7158,N_7591);
xor U8489 (N_8489,N_7767,N_7484);
xnor U8490 (N_8490,N_7290,N_7239);
or U8491 (N_8491,N_7705,N_7687);
nor U8492 (N_8492,N_7803,N_7652);
nor U8493 (N_8493,N_7039,N_7423);
or U8494 (N_8494,N_7860,N_7520);
nand U8495 (N_8495,N_7421,N_7943);
and U8496 (N_8496,N_7071,N_7863);
xor U8497 (N_8497,N_7163,N_7080);
nand U8498 (N_8498,N_7881,N_7971);
nor U8499 (N_8499,N_7027,N_7564);
and U8500 (N_8500,N_7369,N_7900);
nand U8501 (N_8501,N_7097,N_7061);
nand U8502 (N_8502,N_7380,N_7867);
nor U8503 (N_8503,N_7605,N_7493);
nand U8504 (N_8504,N_7080,N_7955);
nor U8505 (N_8505,N_7473,N_7826);
and U8506 (N_8506,N_7157,N_7337);
nand U8507 (N_8507,N_7785,N_7437);
or U8508 (N_8508,N_7982,N_7597);
nand U8509 (N_8509,N_7709,N_7905);
or U8510 (N_8510,N_7107,N_7750);
xor U8511 (N_8511,N_7230,N_7382);
and U8512 (N_8512,N_7676,N_7482);
or U8513 (N_8513,N_7462,N_7187);
or U8514 (N_8514,N_7357,N_7338);
xor U8515 (N_8515,N_7434,N_7715);
xor U8516 (N_8516,N_7761,N_7535);
nand U8517 (N_8517,N_7437,N_7134);
and U8518 (N_8518,N_7225,N_7262);
or U8519 (N_8519,N_7695,N_7130);
nor U8520 (N_8520,N_7660,N_7187);
nor U8521 (N_8521,N_7112,N_7986);
nand U8522 (N_8522,N_7999,N_7629);
xnor U8523 (N_8523,N_7319,N_7902);
or U8524 (N_8524,N_7654,N_7788);
or U8525 (N_8525,N_7558,N_7692);
nor U8526 (N_8526,N_7658,N_7151);
nor U8527 (N_8527,N_7597,N_7305);
or U8528 (N_8528,N_7287,N_7959);
or U8529 (N_8529,N_7994,N_7809);
and U8530 (N_8530,N_7065,N_7072);
or U8531 (N_8531,N_7817,N_7513);
and U8532 (N_8532,N_7038,N_7611);
nor U8533 (N_8533,N_7664,N_7579);
or U8534 (N_8534,N_7103,N_7119);
xnor U8535 (N_8535,N_7116,N_7718);
or U8536 (N_8536,N_7027,N_7538);
or U8537 (N_8537,N_7918,N_7204);
nor U8538 (N_8538,N_7775,N_7703);
nor U8539 (N_8539,N_7721,N_7594);
nor U8540 (N_8540,N_7986,N_7110);
nor U8541 (N_8541,N_7849,N_7450);
nand U8542 (N_8542,N_7820,N_7007);
or U8543 (N_8543,N_7545,N_7631);
or U8544 (N_8544,N_7410,N_7022);
or U8545 (N_8545,N_7887,N_7910);
xnor U8546 (N_8546,N_7451,N_7186);
or U8547 (N_8547,N_7849,N_7263);
xnor U8548 (N_8548,N_7179,N_7251);
nor U8549 (N_8549,N_7366,N_7382);
nand U8550 (N_8550,N_7730,N_7423);
xnor U8551 (N_8551,N_7506,N_7151);
nand U8552 (N_8552,N_7036,N_7320);
nand U8553 (N_8553,N_7117,N_7996);
nand U8554 (N_8554,N_7949,N_7680);
nand U8555 (N_8555,N_7250,N_7074);
or U8556 (N_8556,N_7442,N_7195);
nor U8557 (N_8557,N_7673,N_7707);
and U8558 (N_8558,N_7966,N_7208);
nor U8559 (N_8559,N_7907,N_7745);
nor U8560 (N_8560,N_7023,N_7866);
and U8561 (N_8561,N_7761,N_7641);
or U8562 (N_8562,N_7106,N_7244);
xor U8563 (N_8563,N_7513,N_7546);
and U8564 (N_8564,N_7671,N_7023);
or U8565 (N_8565,N_7466,N_7756);
and U8566 (N_8566,N_7754,N_7117);
nor U8567 (N_8567,N_7116,N_7234);
and U8568 (N_8568,N_7847,N_7198);
nand U8569 (N_8569,N_7616,N_7675);
or U8570 (N_8570,N_7665,N_7980);
xor U8571 (N_8571,N_7903,N_7300);
nand U8572 (N_8572,N_7931,N_7788);
or U8573 (N_8573,N_7977,N_7075);
or U8574 (N_8574,N_7860,N_7589);
nand U8575 (N_8575,N_7880,N_7794);
and U8576 (N_8576,N_7632,N_7575);
nor U8577 (N_8577,N_7096,N_7185);
nor U8578 (N_8578,N_7022,N_7178);
xor U8579 (N_8579,N_7288,N_7981);
nor U8580 (N_8580,N_7555,N_7077);
nand U8581 (N_8581,N_7752,N_7274);
xnor U8582 (N_8582,N_7030,N_7396);
xnor U8583 (N_8583,N_7484,N_7926);
and U8584 (N_8584,N_7041,N_7971);
xor U8585 (N_8585,N_7390,N_7631);
nor U8586 (N_8586,N_7709,N_7350);
nor U8587 (N_8587,N_7035,N_7792);
xnor U8588 (N_8588,N_7747,N_7637);
xnor U8589 (N_8589,N_7687,N_7119);
and U8590 (N_8590,N_7350,N_7295);
nor U8591 (N_8591,N_7079,N_7298);
nor U8592 (N_8592,N_7209,N_7130);
xnor U8593 (N_8593,N_7344,N_7999);
or U8594 (N_8594,N_7687,N_7721);
and U8595 (N_8595,N_7648,N_7931);
and U8596 (N_8596,N_7333,N_7794);
nor U8597 (N_8597,N_7306,N_7264);
or U8598 (N_8598,N_7998,N_7596);
nor U8599 (N_8599,N_7401,N_7281);
and U8600 (N_8600,N_7435,N_7481);
nand U8601 (N_8601,N_7966,N_7383);
xor U8602 (N_8602,N_7547,N_7974);
and U8603 (N_8603,N_7470,N_7250);
nor U8604 (N_8604,N_7612,N_7461);
and U8605 (N_8605,N_7196,N_7394);
nand U8606 (N_8606,N_7038,N_7981);
xor U8607 (N_8607,N_7100,N_7847);
xor U8608 (N_8608,N_7111,N_7430);
and U8609 (N_8609,N_7695,N_7431);
and U8610 (N_8610,N_7090,N_7408);
nor U8611 (N_8611,N_7885,N_7417);
and U8612 (N_8612,N_7703,N_7095);
nand U8613 (N_8613,N_7522,N_7818);
nand U8614 (N_8614,N_7812,N_7786);
and U8615 (N_8615,N_7794,N_7885);
xnor U8616 (N_8616,N_7966,N_7620);
or U8617 (N_8617,N_7726,N_7799);
and U8618 (N_8618,N_7841,N_7075);
nor U8619 (N_8619,N_7896,N_7973);
or U8620 (N_8620,N_7911,N_7018);
xor U8621 (N_8621,N_7587,N_7962);
nor U8622 (N_8622,N_7379,N_7457);
and U8623 (N_8623,N_7873,N_7058);
xor U8624 (N_8624,N_7696,N_7819);
and U8625 (N_8625,N_7711,N_7781);
and U8626 (N_8626,N_7115,N_7321);
nor U8627 (N_8627,N_7050,N_7967);
xnor U8628 (N_8628,N_7837,N_7205);
or U8629 (N_8629,N_7912,N_7312);
nand U8630 (N_8630,N_7694,N_7934);
or U8631 (N_8631,N_7183,N_7953);
nand U8632 (N_8632,N_7081,N_7868);
and U8633 (N_8633,N_7496,N_7818);
xor U8634 (N_8634,N_7702,N_7337);
nand U8635 (N_8635,N_7499,N_7375);
and U8636 (N_8636,N_7570,N_7664);
nor U8637 (N_8637,N_7351,N_7720);
xor U8638 (N_8638,N_7566,N_7228);
or U8639 (N_8639,N_7278,N_7284);
nand U8640 (N_8640,N_7828,N_7403);
nand U8641 (N_8641,N_7637,N_7628);
and U8642 (N_8642,N_7711,N_7405);
nand U8643 (N_8643,N_7525,N_7362);
xor U8644 (N_8644,N_7353,N_7015);
or U8645 (N_8645,N_7486,N_7150);
nor U8646 (N_8646,N_7641,N_7251);
or U8647 (N_8647,N_7702,N_7680);
nor U8648 (N_8648,N_7592,N_7124);
or U8649 (N_8649,N_7770,N_7004);
nand U8650 (N_8650,N_7730,N_7967);
nand U8651 (N_8651,N_7984,N_7446);
nor U8652 (N_8652,N_7036,N_7301);
and U8653 (N_8653,N_7809,N_7067);
nand U8654 (N_8654,N_7552,N_7748);
xor U8655 (N_8655,N_7514,N_7664);
nor U8656 (N_8656,N_7089,N_7931);
nand U8657 (N_8657,N_7403,N_7874);
and U8658 (N_8658,N_7841,N_7340);
or U8659 (N_8659,N_7581,N_7685);
nand U8660 (N_8660,N_7208,N_7902);
and U8661 (N_8661,N_7110,N_7953);
nand U8662 (N_8662,N_7896,N_7230);
xnor U8663 (N_8663,N_7492,N_7138);
nor U8664 (N_8664,N_7686,N_7365);
or U8665 (N_8665,N_7888,N_7201);
nand U8666 (N_8666,N_7764,N_7959);
and U8667 (N_8667,N_7333,N_7036);
xnor U8668 (N_8668,N_7996,N_7152);
nor U8669 (N_8669,N_7202,N_7736);
nor U8670 (N_8670,N_7913,N_7210);
and U8671 (N_8671,N_7845,N_7681);
nand U8672 (N_8672,N_7261,N_7799);
and U8673 (N_8673,N_7790,N_7907);
or U8674 (N_8674,N_7544,N_7867);
nand U8675 (N_8675,N_7728,N_7269);
and U8676 (N_8676,N_7508,N_7235);
xnor U8677 (N_8677,N_7352,N_7687);
nor U8678 (N_8678,N_7441,N_7625);
nor U8679 (N_8679,N_7179,N_7762);
or U8680 (N_8680,N_7369,N_7203);
nand U8681 (N_8681,N_7618,N_7413);
nor U8682 (N_8682,N_7057,N_7737);
nor U8683 (N_8683,N_7874,N_7128);
or U8684 (N_8684,N_7333,N_7072);
and U8685 (N_8685,N_7472,N_7067);
or U8686 (N_8686,N_7154,N_7542);
and U8687 (N_8687,N_7190,N_7389);
nand U8688 (N_8688,N_7356,N_7893);
nand U8689 (N_8689,N_7692,N_7598);
xnor U8690 (N_8690,N_7854,N_7864);
xor U8691 (N_8691,N_7639,N_7370);
nor U8692 (N_8692,N_7135,N_7263);
nor U8693 (N_8693,N_7680,N_7419);
or U8694 (N_8694,N_7322,N_7515);
nand U8695 (N_8695,N_7382,N_7830);
or U8696 (N_8696,N_7983,N_7752);
nand U8697 (N_8697,N_7676,N_7696);
and U8698 (N_8698,N_7118,N_7768);
and U8699 (N_8699,N_7474,N_7957);
and U8700 (N_8700,N_7911,N_7628);
nand U8701 (N_8701,N_7672,N_7639);
nor U8702 (N_8702,N_7673,N_7007);
xor U8703 (N_8703,N_7132,N_7118);
or U8704 (N_8704,N_7166,N_7990);
and U8705 (N_8705,N_7580,N_7536);
or U8706 (N_8706,N_7091,N_7813);
nor U8707 (N_8707,N_7766,N_7041);
nand U8708 (N_8708,N_7986,N_7757);
or U8709 (N_8709,N_7124,N_7753);
and U8710 (N_8710,N_7903,N_7079);
xnor U8711 (N_8711,N_7776,N_7979);
and U8712 (N_8712,N_7766,N_7477);
xnor U8713 (N_8713,N_7314,N_7834);
xnor U8714 (N_8714,N_7832,N_7826);
and U8715 (N_8715,N_7624,N_7076);
nor U8716 (N_8716,N_7488,N_7691);
nor U8717 (N_8717,N_7112,N_7887);
nor U8718 (N_8718,N_7590,N_7679);
nand U8719 (N_8719,N_7877,N_7553);
and U8720 (N_8720,N_7430,N_7502);
nand U8721 (N_8721,N_7516,N_7771);
xor U8722 (N_8722,N_7893,N_7743);
or U8723 (N_8723,N_7922,N_7570);
nor U8724 (N_8724,N_7773,N_7055);
nor U8725 (N_8725,N_7753,N_7669);
xor U8726 (N_8726,N_7298,N_7378);
nor U8727 (N_8727,N_7546,N_7814);
or U8728 (N_8728,N_7609,N_7047);
nand U8729 (N_8729,N_7214,N_7213);
and U8730 (N_8730,N_7385,N_7091);
nand U8731 (N_8731,N_7816,N_7016);
nand U8732 (N_8732,N_7845,N_7091);
nand U8733 (N_8733,N_7667,N_7171);
nand U8734 (N_8734,N_7377,N_7320);
nor U8735 (N_8735,N_7090,N_7736);
nand U8736 (N_8736,N_7006,N_7748);
xnor U8737 (N_8737,N_7545,N_7168);
or U8738 (N_8738,N_7781,N_7677);
and U8739 (N_8739,N_7659,N_7107);
nand U8740 (N_8740,N_7138,N_7193);
and U8741 (N_8741,N_7380,N_7988);
xor U8742 (N_8742,N_7070,N_7535);
and U8743 (N_8743,N_7053,N_7381);
and U8744 (N_8744,N_7529,N_7249);
xor U8745 (N_8745,N_7143,N_7907);
xor U8746 (N_8746,N_7210,N_7880);
and U8747 (N_8747,N_7263,N_7294);
nand U8748 (N_8748,N_7377,N_7032);
nand U8749 (N_8749,N_7749,N_7969);
nor U8750 (N_8750,N_7254,N_7849);
nor U8751 (N_8751,N_7765,N_7930);
nand U8752 (N_8752,N_7238,N_7449);
and U8753 (N_8753,N_7677,N_7463);
nor U8754 (N_8754,N_7363,N_7572);
xor U8755 (N_8755,N_7757,N_7840);
nor U8756 (N_8756,N_7257,N_7887);
and U8757 (N_8757,N_7769,N_7026);
or U8758 (N_8758,N_7021,N_7309);
nand U8759 (N_8759,N_7431,N_7461);
and U8760 (N_8760,N_7138,N_7260);
xor U8761 (N_8761,N_7057,N_7144);
xnor U8762 (N_8762,N_7109,N_7901);
nand U8763 (N_8763,N_7703,N_7945);
and U8764 (N_8764,N_7052,N_7071);
nand U8765 (N_8765,N_7637,N_7729);
xnor U8766 (N_8766,N_7065,N_7100);
or U8767 (N_8767,N_7116,N_7595);
nand U8768 (N_8768,N_7696,N_7128);
or U8769 (N_8769,N_7160,N_7550);
xor U8770 (N_8770,N_7384,N_7004);
or U8771 (N_8771,N_7906,N_7735);
or U8772 (N_8772,N_7002,N_7294);
xnor U8773 (N_8773,N_7089,N_7348);
xor U8774 (N_8774,N_7928,N_7798);
nand U8775 (N_8775,N_7387,N_7097);
xor U8776 (N_8776,N_7302,N_7694);
or U8777 (N_8777,N_7964,N_7086);
xor U8778 (N_8778,N_7881,N_7104);
or U8779 (N_8779,N_7334,N_7386);
nand U8780 (N_8780,N_7093,N_7861);
and U8781 (N_8781,N_7367,N_7106);
or U8782 (N_8782,N_7903,N_7323);
and U8783 (N_8783,N_7238,N_7821);
nor U8784 (N_8784,N_7954,N_7601);
xnor U8785 (N_8785,N_7780,N_7642);
and U8786 (N_8786,N_7101,N_7321);
xor U8787 (N_8787,N_7823,N_7552);
nand U8788 (N_8788,N_7000,N_7890);
nand U8789 (N_8789,N_7640,N_7368);
nand U8790 (N_8790,N_7686,N_7225);
or U8791 (N_8791,N_7540,N_7139);
xnor U8792 (N_8792,N_7613,N_7063);
nand U8793 (N_8793,N_7502,N_7428);
nor U8794 (N_8794,N_7720,N_7175);
and U8795 (N_8795,N_7461,N_7547);
and U8796 (N_8796,N_7696,N_7833);
or U8797 (N_8797,N_7927,N_7949);
nand U8798 (N_8798,N_7683,N_7533);
and U8799 (N_8799,N_7709,N_7628);
xor U8800 (N_8800,N_7985,N_7128);
nor U8801 (N_8801,N_7193,N_7243);
nand U8802 (N_8802,N_7117,N_7167);
xnor U8803 (N_8803,N_7663,N_7234);
nand U8804 (N_8804,N_7236,N_7768);
xnor U8805 (N_8805,N_7806,N_7160);
or U8806 (N_8806,N_7341,N_7895);
and U8807 (N_8807,N_7174,N_7252);
nor U8808 (N_8808,N_7157,N_7811);
or U8809 (N_8809,N_7666,N_7589);
nor U8810 (N_8810,N_7654,N_7212);
xnor U8811 (N_8811,N_7214,N_7362);
and U8812 (N_8812,N_7132,N_7889);
xnor U8813 (N_8813,N_7962,N_7387);
nand U8814 (N_8814,N_7405,N_7790);
nor U8815 (N_8815,N_7564,N_7435);
nand U8816 (N_8816,N_7413,N_7115);
nand U8817 (N_8817,N_7149,N_7830);
nand U8818 (N_8818,N_7035,N_7582);
xor U8819 (N_8819,N_7907,N_7424);
xnor U8820 (N_8820,N_7555,N_7150);
nand U8821 (N_8821,N_7354,N_7062);
nor U8822 (N_8822,N_7832,N_7710);
nor U8823 (N_8823,N_7485,N_7947);
and U8824 (N_8824,N_7499,N_7885);
nor U8825 (N_8825,N_7815,N_7512);
and U8826 (N_8826,N_7039,N_7278);
and U8827 (N_8827,N_7623,N_7793);
and U8828 (N_8828,N_7149,N_7521);
nand U8829 (N_8829,N_7648,N_7704);
xnor U8830 (N_8830,N_7077,N_7948);
and U8831 (N_8831,N_7824,N_7162);
xor U8832 (N_8832,N_7618,N_7879);
and U8833 (N_8833,N_7085,N_7902);
xnor U8834 (N_8834,N_7321,N_7206);
xor U8835 (N_8835,N_7157,N_7277);
xor U8836 (N_8836,N_7742,N_7232);
xor U8837 (N_8837,N_7979,N_7694);
or U8838 (N_8838,N_7965,N_7541);
or U8839 (N_8839,N_7919,N_7901);
and U8840 (N_8840,N_7301,N_7141);
or U8841 (N_8841,N_7703,N_7534);
and U8842 (N_8842,N_7962,N_7814);
xnor U8843 (N_8843,N_7470,N_7211);
nor U8844 (N_8844,N_7676,N_7877);
xor U8845 (N_8845,N_7704,N_7183);
nand U8846 (N_8846,N_7523,N_7236);
xnor U8847 (N_8847,N_7390,N_7203);
and U8848 (N_8848,N_7840,N_7548);
or U8849 (N_8849,N_7011,N_7882);
or U8850 (N_8850,N_7164,N_7928);
nor U8851 (N_8851,N_7711,N_7639);
or U8852 (N_8852,N_7813,N_7317);
nand U8853 (N_8853,N_7551,N_7878);
and U8854 (N_8854,N_7549,N_7605);
nor U8855 (N_8855,N_7896,N_7586);
or U8856 (N_8856,N_7010,N_7543);
and U8857 (N_8857,N_7672,N_7466);
and U8858 (N_8858,N_7609,N_7817);
nand U8859 (N_8859,N_7174,N_7125);
or U8860 (N_8860,N_7818,N_7885);
or U8861 (N_8861,N_7901,N_7131);
xor U8862 (N_8862,N_7900,N_7224);
or U8863 (N_8863,N_7646,N_7241);
nand U8864 (N_8864,N_7352,N_7788);
nand U8865 (N_8865,N_7947,N_7461);
nor U8866 (N_8866,N_7041,N_7169);
nand U8867 (N_8867,N_7210,N_7409);
and U8868 (N_8868,N_7302,N_7130);
nand U8869 (N_8869,N_7110,N_7105);
nand U8870 (N_8870,N_7390,N_7886);
nor U8871 (N_8871,N_7965,N_7626);
xnor U8872 (N_8872,N_7702,N_7104);
xnor U8873 (N_8873,N_7248,N_7255);
nor U8874 (N_8874,N_7400,N_7856);
and U8875 (N_8875,N_7848,N_7797);
xnor U8876 (N_8876,N_7969,N_7926);
xnor U8877 (N_8877,N_7564,N_7770);
and U8878 (N_8878,N_7731,N_7738);
and U8879 (N_8879,N_7250,N_7711);
xnor U8880 (N_8880,N_7758,N_7507);
or U8881 (N_8881,N_7518,N_7077);
nand U8882 (N_8882,N_7755,N_7936);
nand U8883 (N_8883,N_7816,N_7904);
or U8884 (N_8884,N_7272,N_7957);
xor U8885 (N_8885,N_7394,N_7404);
nand U8886 (N_8886,N_7367,N_7073);
nor U8887 (N_8887,N_7755,N_7586);
xor U8888 (N_8888,N_7039,N_7587);
xnor U8889 (N_8889,N_7276,N_7459);
or U8890 (N_8890,N_7752,N_7228);
nor U8891 (N_8891,N_7327,N_7441);
nand U8892 (N_8892,N_7094,N_7351);
and U8893 (N_8893,N_7559,N_7085);
nand U8894 (N_8894,N_7358,N_7846);
and U8895 (N_8895,N_7876,N_7191);
nor U8896 (N_8896,N_7816,N_7489);
and U8897 (N_8897,N_7390,N_7463);
xnor U8898 (N_8898,N_7675,N_7529);
and U8899 (N_8899,N_7773,N_7634);
nor U8900 (N_8900,N_7645,N_7677);
and U8901 (N_8901,N_7895,N_7581);
xnor U8902 (N_8902,N_7577,N_7203);
nor U8903 (N_8903,N_7227,N_7728);
and U8904 (N_8904,N_7575,N_7562);
or U8905 (N_8905,N_7199,N_7021);
and U8906 (N_8906,N_7281,N_7024);
nor U8907 (N_8907,N_7956,N_7961);
or U8908 (N_8908,N_7724,N_7559);
nor U8909 (N_8909,N_7474,N_7396);
and U8910 (N_8910,N_7608,N_7692);
and U8911 (N_8911,N_7893,N_7895);
or U8912 (N_8912,N_7058,N_7971);
nand U8913 (N_8913,N_7326,N_7325);
or U8914 (N_8914,N_7752,N_7090);
or U8915 (N_8915,N_7080,N_7894);
or U8916 (N_8916,N_7119,N_7653);
nand U8917 (N_8917,N_7310,N_7863);
and U8918 (N_8918,N_7249,N_7879);
xor U8919 (N_8919,N_7249,N_7201);
or U8920 (N_8920,N_7381,N_7284);
xnor U8921 (N_8921,N_7591,N_7912);
xnor U8922 (N_8922,N_7332,N_7879);
and U8923 (N_8923,N_7991,N_7890);
nor U8924 (N_8924,N_7429,N_7293);
or U8925 (N_8925,N_7112,N_7020);
or U8926 (N_8926,N_7644,N_7978);
and U8927 (N_8927,N_7176,N_7678);
xor U8928 (N_8928,N_7513,N_7925);
nor U8929 (N_8929,N_7888,N_7331);
nand U8930 (N_8930,N_7470,N_7660);
nand U8931 (N_8931,N_7754,N_7546);
xnor U8932 (N_8932,N_7182,N_7663);
nor U8933 (N_8933,N_7688,N_7652);
or U8934 (N_8934,N_7998,N_7480);
and U8935 (N_8935,N_7806,N_7760);
xor U8936 (N_8936,N_7937,N_7790);
nor U8937 (N_8937,N_7171,N_7194);
nor U8938 (N_8938,N_7342,N_7627);
nor U8939 (N_8939,N_7001,N_7514);
or U8940 (N_8940,N_7770,N_7756);
and U8941 (N_8941,N_7674,N_7013);
xnor U8942 (N_8942,N_7142,N_7440);
or U8943 (N_8943,N_7509,N_7955);
nor U8944 (N_8944,N_7259,N_7605);
and U8945 (N_8945,N_7567,N_7664);
xnor U8946 (N_8946,N_7281,N_7736);
xnor U8947 (N_8947,N_7167,N_7755);
xor U8948 (N_8948,N_7660,N_7515);
nor U8949 (N_8949,N_7075,N_7902);
nor U8950 (N_8950,N_7114,N_7629);
or U8951 (N_8951,N_7823,N_7988);
or U8952 (N_8952,N_7218,N_7913);
nand U8953 (N_8953,N_7208,N_7592);
xor U8954 (N_8954,N_7071,N_7207);
nand U8955 (N_8955,N_7368,N_7906);
or U8956 (N_8956,N_7490,N_7569);
and U8957 (N_8957,N_7636,N_7088);
or U8958 (N_8958,N_7896,N_7953);
or U8959 (N_8959,N_7464,N_7264);
and U8960 (N_8960,N_7289,N_7453);
nand U8961 (N_8961,N_7389,N_7876);
nand U8962 (N_8962,N_7366,N_7259);
or U8963 (N_8963,N_7346,N_7106);
xor U8964 (N_8964,N_7292,N_7999);
and U8965 (N_8965,N_7279,N_7942);
and U8966 (N_8966,N_7175,N_7177);
xor U8967 (N_8967,N_7139,N_7274);
nand U8968 (N_8968,N_7071,N_7608);
xor U8969 (N_8969,N_7012,N_7379);
xor U8970 (N_8970,N_7504,N_7764);
and U8971 (N_8971,N_7173,N_7778);
or U8972 (N_8972,N_7507,N_7824);
xnor U8973 (N_8973,N_7691,N_7946);
xor U8974 (N_8974,N_7384,N_7875);
nand U8975 (N_8975,N_7252,N_7541);
and U8976 (N_8976,N_7934,N_7788);
xnor U8977 (N_8977,N_7903,N_7613);
or U8978 (N_8978,N_7140,N_7187);
nor U8979 (N_8979,N_7243,N_7935);
or U8980 (N_8980,N_7810,N_7078);
or U8981 (N_8981,N_7802,N_7839);
xor U8982 (N_8982,N_7688,N_7410);
nand U8983 (N_8983,N_7233,N_7143);
or U8984 (N_8984,N_7753,N_7288);
nor U8985 (N_8985,N_7076,N_7290);
nand U8986 (N_8986,N_7590,N_7843);
and U8987 (N_8987,N_7527,N_7669);
nand U8988 (N_8988,N_7003,N_7411);
and U8989 (N_8989,N_7470,N_7457);
nor U8990 (N_8990,N_7920,N_7986);
xnor U8991 (N_8991,N_7929,N_7855);
nor U8992 (N_8992,N_7252,N_7315);
xnor U8993 (N_8993,N_7200,N_7535);
nor U8994 (N_8994,N_7333,N_7339);
nor U8995 (N_8995,N_7038,N_7511);
and U8996 (N_8996,N_7753,N_7417);
nor U8997 (N_8997,N_7196,N_7932);
xor U8998 (N_8998,N_7012,N_7118);
xnor U8999 (N_8999,N_7827,N_7862);
xor U9000 (N_9000,N_8716,N_8015);
and U9001 (N_9001,N_8430,N_8740);
nor U9002 (N_9002,N_8018,N_8849);
xnor U9003 (N_9003,N_8904,N_8076);
and U9004 (N_9004,N_8847,N_8420);
and U9005 (N_9005,N_8379,N_8841);
and U9006 (N_9006,N_8127,N_8779);
xor U9007 (N_9007,N_8217,N_8378);
nand U9008 (N_9008,N_8570,N_8502);
and U9009 (N_9009,N_8343,N_8397);
xnor U9010 (N_9010,N_8968,N_8545);
nor U9011 (N_9011,N_8234,N_8265);
nor U9012 (N_9012,N_8592,N_8607);
nand U9013 (N_9013,N_8778,N_8578);
xor U9014 (N_9014,N_8083,N_8737);
nor U9015 (N_9015,N_8565,N_8838);
and U9016 (N_9016,N_8048,N_8673);
and U9017 (N_9017,N_8872,N_8605);
and U9018 (N_9018,N_8387,N_8562);
xor U9019 (N_9019,N_8577,N_8403);
xor U9020 (N_9020,N_8100,N_8254);
xor U9021 (N_9021,N_8734,N_8978);
nor U9022 (N_9022,N_8557,N_8334);
nor U9023 (N_9023,N_8257,N_8001);
nand U9024 (N_9024,N_8351,N_8161);
nor U9025 (N_9025,N_8029,N_8081);
nor U9026 (N_9026,N_8485,N_8896);
and U9027 (N_9027,N_8766,N_8741);
nand U9028 (N_9028,N_8560,N_8617);
and U9029 (N_9029,N_8452,N_8979);
and U9030 (N_9030,N_8493,N_8044);
nor U9031 (N_9031,N_8084,N_8692);
or U9032 (N_9032,N_8369,N_8456);
xor U9033 (N_9033,N_8394,N_8839);
and U9034 (N_9034,N_8145,N_8151);
nand U9035 (N_9035,N_8213,N_8209);
nand U9036 (N_9036,N_8416,N_8755);
xnor U9037 (N_9037,N_8264,N_8381);
xor U9038 (N_9038,N_8527,N_8666);
xnor U9039 (N_9039,N_8568,N_8763);
nor U9040 (N_9040,N_8431,N_8542);
xnor U9041 (N_9041,N_8694,N_8159);
nor U9042 (N_9042,N_8267,N_8965);
and U9043 (N_9043,N_8483,N_8616);
xor U9044 (N_9044,N_8093,N_8138);
xnor U9045 (N_9045,N_8111,N_8647);
or U9046 (N_9046,N_8762,N_8126);
nand U9047 (N_9047,N_8116,N_8897);
nor U9048 (N_9048,N_8061,N_8525);
nor U9049 (N_9049,N_8675,N_8386);
nor U9050 (N_9050,N_8025,N_8625);
nor U9051 (N_9051,N_8171,N_8890);
xor U9052 (N_9052,N_8406,N_8930);
nor U9053 (N_9053,N_8922,N_8412);
and U9054 (N_9054,N_8540,N_8239);
nor U9055 (N_9055,N_8306,N_8328);
and U9056 (N_9056,N_8595,N_8224);
and U9057 (N_9057,N_8732,N_8682);
or U9058 (N_9058,N_8992,N_8554);
or U9059 (N_9059,N_8150,N_8441);
nor U9060 (N_9060,N_8384,N_8942);
xnor U9061 (N_9061,N_8374,N_8255);
xnor U9062 (N_9062,N_8760,N_8697);
nor U9063 (N_9063,N_8191,N_8047);
nand U9064 (N_9064,N_8020,N_8080);
xor U9065 (N_9065,N_8283,N_8921);
nand U9066 (N_9066,N_8758,N_8098);
xor U9067 (N_9067,N_8569,N_8319);
xor U9068 (N_9068,N_8511,N_8396);
and U9069 (N_9069,N_8999,N_8472);
or U9070 (N_9070,N_8086,N_8726);
or U9071 (N_9071,N_8866,N_8027);
xor U9072 (N_9072,N_8749,N_8376);
or U9073 (N_9073,N_8082,N_8218);
xor U9074 (N_9074,N_8228,N_8411);
and U9075 (N_9075,N_8400,N_8284);
or U9076 (N_9076,N_8658,N_8277);
nand U9077 (N_9077,N_8959,N_8419);
nand U9078 (N_9078,N_8842,N_8413);
nor U9079 (N_9079,N_8193,N_8905);
and U9080 (N_9080,N_8085,N_8961);
or U9081 (N_9081,N_8977,N_8517);
nor U9082 (N_9082,N_8809,N_8855);
nor U9083 (N_9083,N_8674,N_8588);
or U9084 (N_9084,N_8782,N_8739);
and U9085 (N_9085,N_8122,N_8520);
nor U9086 (N_9086,N_8875,N_8314);
or U9087 (N_9087,N_8795,N_8365);
nor U9088 (N_9088,N_8070,N_8305);
or U9089 (N_9089,N_8055,N_8688);
xor U9090 (N_9090,N_8153,N_8745);
xor U9091 (N_9091,N_8280,N_8194);
or U9092 (N_9092,N_8719,N_8722);
or U9093 (N_9093,N_8933,N_8495);
or U9094 (N_9094,N_8884,N_8501);
nor U9095 (N_9095,N_8892,N_8623);
and U9096 (N_9096,N_8939,N_8160);
or U9097 (N_9097,N_8442,N_8183);
and U9098 (N_9098,N_8805,N_8765);
or U9099 (N_9099,N_8212,N_8405);
xor U9100 (N_9100,N_8832,N_8598);
and U9101 (N_9101,N_8259,N_8262);
nand U9102 (N_9102,N_8951,N_8993);
or U9103 (N_9103,N_8211,N_8059);
xnor U9104 (N_9104,N_8634,N_8561);
or U9105 (N_9105,N_8534,N_8974);
xnor U9106 (N_9106,N_8445,N_8702);
xor U9107 (N_9107,N_8465,N_8219);
xnor U9108 (N_9108,N_8862,N_8606);
xnor U9109 (N_9109,N_8712,N_8711);
nor U9110 (N_9110,N_8115,N_8476);
nand U9111 (N_9111,N_8898,N_8589);
or U9112 (N_9112,N_8332,N_8735);
nor U9113 (N_9113,N_8176,N_8834);
nand U9114 (N_9114,N_8601,N_8099);
nand U9115 (N_9115,N_8035,N_8507);
or U9116 (N_9116,N_8757,N_8482);
nor U9117 (N_9117,N_8192,N_8698);
nand U9118 (N_9118,N_8425,N_8915);
xnor U9119 (N_9119,N_8731,N_8621);
nor U9120 (N_9120,N_8162,N_8272);
and U9121 (N_9121,N_8117,N_8803);
nor U9122 (N_9122,N_8132,N_8137);
nand U9123 (N_9123,N_8541,N_8913);
or U9124 (N_9124,N_8944,N_8798);
nand U9125 (N_9125,N_8903,N_8889);
nand U9126 (N_9126,N_8355,N_8599);
and U9127 (N_9127,N_8934,N_8385);
nor U9128 (N_9128,N_8096,N_8492);
and U9129 (N_9129,N_8079,N_8244);
and U9130 (N_9130,N_8156,N_8268);
and U9131 (N_9131,N_8195,N_8134);
nor U9132 (N_9132,N_8208,N_8584);
and U9133 (N_9133,N_8651,N_8626);
xor U9134 (N_9134,N_8072,N_8349);
xor U9135 (N_9135,N_8490,N_8513);
and U9136 (N_9136,N_8278,N_8781);
xnor U9137 (N_9137,N_8670,N_8181);
or U9138 (N_9138,N_8235,N_8356);
xnor U9139 (N_9139,N_8914,N_8232);
nor U9140 (N_9140,N_8699,N_8609);
and U9141 (N_9141,N_8249,N_8346);
or U9142 (N_9142,N_8230,N_8457);
and U9143 (N_9143,N_8250,N_8243);
or U9144 (N_9144,N_8556,N_8170);
and U9145 (N_9145,N_8986,N_8147);
nand U9146 (N_9146,N_8375,N_8207);
xnor U9147 (N_9147,N_8019,N_8506);
and U9148 (N_9148,N_8016,N_8410);
nor U9149 (N_9149,N_8481,N_8290);
and U9150 (N_9150,N_8491,N_8748);
and U9151 (N_9151,N_8330,N_8891);
and U9152 (N_9152,N_8812,N_8754);
xnor U9153 (N_9153,N_8785,N_8987);
xnor U9154 (N_9154,N_8260,N_8409);
nor U9155 (N_9155,N_8367,N_8777);
and U9156 (N_9156,N_8045,N_8067);
nor U9157 (N_9157,N_8276,N_8215);
and U9158 (N_9158,N_8058,N_8401);
nand U9159 (N_9159,N_8868,N_8344);
and U9160 (N_9160,N_8470,N_8124);
nor U9161 (N_9161,N_8318,N_8037);
nand U9162 (N_9162,N_8475,N_8860);
and U9163 (N_9163,N_8449,N_8786);
xor U9164 (N_9164,N_8797,N_8389);
or U9165 (N_9165,N_8774,N_8919);
nand U9166 (N_9166,N_8043,N_8202);
and U9167 (N_9167,N_8662,N_8801);
nand U9168 (N_9168,N_8619,N_8908);
or U9169 (N_9169,N_8585,N_8256);
nor U9170 (N_9170,N_8825,N_8970);
xnor U9171 (N_9171,N_8246,N_8173);
xnor U9172 (N_9172,N_8929,N_8461);
nor U9173 (N_9173,N_8281,N_8627);
and U9174 (N_9174,N_8852,N_8382);
or U9175 (N_9175,N_8874,N_8336);
or U9176 (N_9176,N_8575,N_8509);
xnor U9177 (N_9177,N_8604,N_8247);
and U9178 (N_9178,N_8851,N_8972);
and U9179 (N_9179,N_8088,N_8291);
nor U9180 (N_9180,N_8845,N_8295);
and U9181 (N_9181,N_8856,N_8641);
xnor U9182 (N_9182,N_8225,N_8593);
xnor U9183 (N_9183,N_8166,N_8279);
xnor U9184 (N_9184,N_8148,N_8790);
or U9185 (N_9185,N_8678,N_8631);
and U9186 (N_9186,N_8667,N_8990);
and U9187 (N_9187,N_8187,N_8414);
and U9188 (N_9188,N_8340,N_8041);
or U9189 (N_9189,N_8530,N_8804);
xnor U9190 (N_9190,N_8120,N_8309);
nand U9191 (N_9191,N_8854,N_8690);
or U9192 (N_9192,N_8761,N_8206);
and U9193 (N_9193,N_8303,N_8971);
and U9194 (N_9194,N_8906,N_8912);
or U9195 (N_9195,N_8299,N_8301);
nor U9196 (N_9196,N_8700,N_8710);
and U9197 (N_9197,N_8582,N_8358);
nand U9198 (N_9198,N_8240,N_8338);
or U9199 (N_9199,N_8594,N_8819);
nor U9200 (N_9200,N_8065,N_8455);
nand U9201 (N_9201,N_8460,N_8214);
and U9202 (N_9202,N_8364,N_8848);
and U9203 (N_9203,N_8723,N_8097);
and U9204 (N_9204,N_8226,N_8251);
or U9205 (N_9205,N_8611,N_8973);
and U9206 (N_9206,N_8721,N_8200);
nand U9207 (N_9207,N_8300,N_8596);
or U9208 (N_9208,N_8069,N_8546);
or U9209 (N_9209,N_8636,N_8021);
nand U9210 (N_9210,N_8806,N_8885);
nor U9211 (N_9211,N_8931,N_8899);
xor U9212 (N_9212,N_8424,N_8927);
nor U9213 (N_9213,N_8229,N_8007);
xnor U9214 (N_9214,N_8529,N_8233);
nand U9215 (N_9215,N_8687,N_8826);
or U9216 (N_9216,N_8296,N_8288);
nor U9217 (N_9217,N_8574,N_8423);
or U9218 (N_9218,N_8821,N_8664);
nor U9219 (N_9219,N_8600,N_8454);
or U9220 (N_9220,N_8853,N_8026);
xnor U9221 (N_9221,N_8759,N_8579);
and U9222 (N_9222,N_8936,N_8946);
xor U9223 (N_9223,N_8926,N_8780);
xnor U9224 (N_9224,N_8962,N_8034);
xor U9225 (N_9225,N_8443,N_8293);
xnor U9226 (N_9226,N_8075,N_8348);
or U9227 (N_9227,N_8564,N_8652);
nand U9228 (N_9228,N_8677,N_8494);
nand U9229 (N_9229,N_8107,N_8354);
xnor U9230 (N_9230,N_8125,N_8695);
nor U9231 (N_9231,N_8738,N_8857);
xnor U9232 (N_9232,N_8222,N_8794);
nand U9233 (N_9233,N_8679,N_8121);
xnor U9234 (N_9234,N_8179,N_8660);
and U9235 (N_9235,N_8182,N_8508);
and U9236 (N_9236,N_8154,N_8656);
or U9237 (N_9237,N_8923,N_8516);
nand U9238 (N_9238,N_8373,N_8510);
xnor U9239 (N_9239,N_8633,N_8415);
nand U9240 (N_9240,N_8448,N_8101);
nor U9241 (N_9241,N_8713,N_8089);
nand U9242 (N_9242,N_8672,N_8129);
nand U9243 (N_9243,N_8966,N_8004);
nor U9244 (N_9244,N_8360,N_8064);
xor U9245 (N_9245,N_8357,N_8184);
nand U9246 (N_9246,N_8642,N_8325);
or U9247 (N_9247,N_8752,N_8074);
nor U9248 (N_9248,N_8196,N_8624);
nor U9249 (N_9249,N_8543,N_8012);
xnor U9250 (N_9250,N_8747,N_8649);
nor U9251 (N_9251,N_8985,N_8000);
and U9252 (N_9252,N_8808,N_8581);
and U9253 (N_9253,N_8684,N_8049);
or U9254 (N_9254,N_8143,N_8458);
and U9255 (N_9255,N_8705,N_8613);
or U9256 (N_9256,N_8522,N_8275);
xnor U9257 (N_9257,N_8864,N_8395);
xnor U9258 (N_9258,N_8105,N_8302);
nand U9259 (N_9259,N_8620,N_8453);
or U9260 (N_9260,N_8612,N_8789);
and U9261 (N_9261,N_8052,N_8450);
nor U9262 (N_9262,N_8879,N_8539);
nor U9263 (N_9263,N_8068,N_8109);
and U9264 (N_9264,N_8858,N_8062);
or U9265 (N_9265,N_8135,N_8665);
and U9266 (N_9266,N_8937,N_8887);
xor U9267 (N_9267,N_8422,N_8335);
nor U9268 (N_9268,N_8242,N_8066);
nand U9269 (N_9269,N_8133,N_8918);
xnor U9270 (N_9270,N_8210,N_8551);
nor U9271 (N_9271,N_8963,N_8307);
nand U9272 (N_9272,N_8727,N_8655);
and U9273 (N_9273,N_8880,N_8149);
nand U9274 (N_9274,N_8615,N_8438);
and U9275 (N_9275,N_8865,N_8653);
and U9276 (N_9276,N_8802,N_8185);
nand U9277 (N_9277,N_8751,N_8022);
and U9278 (N_9278,N_8683,N_8686);
nand U9279 (N_9279,N_8877,N_8590);
xor U9280 (N_9280,N_8547,N_8362);
and U9281 (N_9281,N_8644,N_8496);
nand U9282 (N_9282,N_8870,N_8515);
and U9283 (N_9283,N_8828,N_8746);
xnor U9284 (N_9284,N_8948,N_8040);
or U9285 (N_9285,N_8427,N_8767);
nor U9286 (N_9286,N_8800,N_8114);
nor U9287 (N_9287,N_8152,N_8622);
nand U9288 (N_9288,N_8289,N_8014);
nand U9289 (N_9289,N_8708,N_8843);
nand U9290 (N_9290,N_8404,N_8236);
and U9291 (N_9291,N_8363,N_8553);
or U9292 (N_9292,N_8544,N_8337);
and U9293 (N_9293,N_8635,N_8046);
nor U9294 (N_9294,N_8947,N_8638);
nand U9295 (N_9295,N_8417,N_8392);
nand U9296 (N_9296,N_8603,N_8042);
nand U9297 (N_9297,N_8324,N_8119);
xor U9298 (N_9298,N_8359,N_8102);
nor U9299 (N_9299,N_8178,N_8753);
and U9300 (N_9300,N_8964,N_8883);
xor U9301 (N_9301,N_8252,N_8792);
and U9302 (N_9302,N_8943,N_8108);
xnor U9303 (N_9303,N_8768,N_8555);
and U9304 (N_9304,N_8190,N_8571);
and U9305 (N_9305,N_8245,N_8796);
xor U9306 (N_9306,N_8463,N_8725);
or U9307 (N_9307,N_8112,N_8895);
or U9308 (N_9308,N_8533,N_8876);
nand U9309 (N_9309,N_8514,N_8432);
and U9310 (N_9310,N_8886,N_8353);
xnor U9311 (N_9311,N_8294,N_8050);
and U9312 (N_9312,N_8311,N_8982);
nand U9313 (N_9313,N_8822,N_8371);
nor U9314 (N_9314,N_8907,N_8459);
nor U9315 (N_9315,N_8051,N_8205);
nor U9316 (N_9316,N_8024,N_8038);
nand U9317 (N_9317,N_8270,N_8998);
xor U9318 (N_9318,N_8783,N_8994);
and U9319 (N_9319,N_8750,N_8715);
and U9320 (N_9320,N_8310,N_8558);
or U9321 (N_9321,N_8580,N_8830);
xor U9322 (N_9322,N_8477,N_8503);
xnor U9323 (N_9323,N_8550,N_8292);
xor U9324 (N_9324,N_8241,N_8984);
nand U9325 (N_9325,N_8691,N_8106);
and U9326 (N_9326,N_8703,N_8274);
and U9327 (N_9327,N_8499,N_8077);
or U9328 (N_9328,N_8057,N_8421);
xnor U9329 (N_9329,N_8816,N_8468);
xnor U9330 (N_9330,N_8981,N_8628);
nor U9331 (N_9331,N_8464,N_8092);
nand U9332 (N_9332,N_8742,N_8141);
nor U9333 (N_9333,N_8829,N_8498);
nor U9334 (N_9334,N_8881,N_8273);
xnor U9335 (N_9335,N_8248,N_8407);
nor U9336 (N_9336,N_8158,N_8017);
nand U9337 (N_9337,N_8435,N_8989);
or U9338 (N_9338,N_8960,N_8180);
xnor U9339 (N_9339,N_8317,N_8304);
nand U9340 (N_9340,N_8479,N_8733);
or U9341 (N_9341,N_8433,N_8439);
nand U9342 (N_9342,N_8380,N_8835);
nand U9343 (N_9343,N_8451,N_8618);
or U9344 (N_9344,N_8536,N_8188);
and U9345 (N_9345,N_8775,N_8039);
nor U9346 (N_9346,N_8429,N_8744);
xor U9347 (N_9347,N_8199,N_8953);
and U9348 (N_9348,N_8920,N_8949);
nand U9349 (N_9349,N_8028,N_8312);
or U9350 (N_9350,N_8729,N_8391);
nand U9351 (N_9351,N_8201,N_8071);
nor U9352 (N_9352,N_8689,N_8002);
or U9353 (N_9353,N_8323,N_8032);
or U9354 (N_9354,N_8011,N_8736);
xor U9355 (N_9355,N_8669,N_8398);
xor U9356 (N_9356,N_8060,N_8282);
nor U9357 (N_9357,N_8350,N_8146);
and U9358 (N_9358,N_8566,N_8900);
and U9359 (N_9359,N_8910,N_8706);
nand U9360 (N_9360,N_8131,N_8444);
and U9361 (N_9361,N_8446,N_8714);
xor U9362 (N_9362,N_8911,N_8950);
nand U9363 (N_9363,N_8873,N_8639);
nor U9364 (N_9364,N_8271,N_8559);
nor U9365 (N_9365,N_8709,N_8958);
nand U9366 (N_9366,N_8327,N_8342);
nand U9367 (N_9367,N_8932,N_8377);
xor U9368 (N_9368,N_8743,N_8637);
and U9369 (N_9369,N_8165,N_8078);
nor U9370 (N_9370,N_8787,N_8010);
or U9371 (N_9371,N_8552,N_8997);
nor U9372 (N_9372,N_8426,N_8013);
nor U9373 (N_9373,N_8928,N_8372);
nor U9374 (N_9374,N_8685,N_8583);
nor U9375 (N_9375,N_8654,N_8893);
nor U9376 (N_9376,N_8663,N_8587);
nor U9377 (N_9377,N_8956,N_8681);
xnor U9378 (N_9378,N_8297,N_8370);
nand U9379 (N_9379,N_8469,N_8693);
nor U9380 (N_9380,N_8103,N_8917);
and U9381 (N_9381,N_8286,N_8671);
nor U9382 (N_9382,N_8329,N_8532);
nand U9383 (N_9383,N_8537,N_8489);
and U9384 (N_9384,N_8473,N_8339);
nor U9385 (N_9385,N_8602,N_8434);
xnor U9386 (N_9386,N_8320,N_8197);
nand U9387 (N_9387,N_8036,N_8680);
xor U9388 (N_9388,N_8894,N_8009);
nor U9389 (N_9389,N_8771,N_8198);
nor U9390 (N_9390,N_8253,N_8823);
or U9391 (N_9391,N_8837,N_8650);
xor U9392 (N_9392,N_8646,N_8586);
nor U9393 (N_9393,N_8846,N_8390);
or U9394 (N_9394,N_8793,N_8844);
or U9395 (N_9395,N_8957,N_8063);
or U9396 (N_9396,N_8110,N_8980);
nand U9397 (N_9397,N_8186,N_8728);
nand U9398 (N_9398,N_8172,N_8478);
nor U9399 (N_9399,N_8231,N_8807);
nor U9400 (N_9400,N_8287,N_8399);
nand U9401 (N_9401,N_8091,N_8657);
nor U9402 (N_9402,N_8827,N_8952);
or U9403 (N_9403,N_8139,N_8720);
xnor U9404 (N_9404,N_8869,N_8563);
and U9405 (N_9405,N_8167,N_8487);
or U9406 (N_9406,N_8056,N_8128);
nand U9407 (N_9407,N_8861,N_8053);
nor U9408 (N_9408,N_8815,N_8704);
and U9409 (N_9409,N_8940,N_8177);
xnor U9410 (N_9410,N_8909,N_8095);
nand U9411 (N_9411,N_8175,N_8157);
nand U9412 (N_9412,N_8006,N_8090);
or U9413 (N_9413,N_8204,N_8155);
nand U9414 (N_9414,N_8203,N_8850);
nand U9415 (N_9415,N_8833,N_8975);
xnor U9416 (N_9416,N_8428,N_8776);
nand U9417 (N_9417,N_8867,N_8003);
nand U9418 (N_9418,N_8144,N_8661);
or U9419 (N_9419,N_8707,N_8811);
nor U9420 (N_9420,N_8189,N_8169);
nor U9421 (N_9421,N_8488,N_8824);
xor U9422 (N_9422,N_8769,N_8916);
and U9423 (N_9423,N_8724,N_8941);
xor U9424 (N_9424,N_8333,N_8368);
and U9425 (N_9425,N_8030,N_8437);
nand U9426 (N_9426,N_8269,N_8788);
and U9427 (N_9427,N_8518,N_8347);
nand U9428 (N_9428,N_8504,N_8174);
or U9429 (N_9429,N_8471,N_8220);
xnor U9430 (N_9430,N_8505,N_8216);
or U9431 (N_9431,N_8925,N_8321);
or U9432 (N_9432,N_8480,N_8447);
xnor U9433 (N_9433,N_8831,N_8954);
xnor U9434 (N_9434,N_8331,N_8466);
or U9435 (N_9435,N_8996,N_8266);
nor U9436 (N_9436,N_8440,N_8326);
and U9437 (N_9437,N_8366,N_8969);
and U9438 (N_9438,N_8770,N_8263);
nand U9439 (N_9439,N_8818,N_8005);
xnor U9440 (N_9440,N_8549,N_8474);
xor U9441 (N_9441,N_8938,N_8572);
and U9442 (N_9442,N_8995,N_8840);
or U9443 (N_9443,N_8967,N_8237);
or U9444 (N_9444,N_8361,N_8168);
xnor U9445 (N_9445,N_8608,N_8418);
or U9446 (N_9446,N_8902,N_8345);
and U9447 (N_9447,N_8227,N_8882);
nand U9448 (N_9448,N_8863,N_8073);
nand U9449 (N_9449,N_8261,N_8659);
xor U9450 (N_9450,N_8648,N_8535);
xor U9451 (N_9451,N_8523,N_8104);
xor U9452 (N_9452,N_8730,N_8526);
and U9453 (N_9453,N_8591,N_8859);
xnor U9454 (N_9454,N_8676,N_8238);
and U9455 (N_9455,N_8629,N_8810);
and U9456 (N_9456,N_8140,N_8988);
xor U9457 (N_9457,N_8772,N_8597);
and U9458 (N_9458,N_8258,N_8548);
and U9459 (N_9459,N_8341,N_8696);
nand U9460 (N_9460,N_8983,N_8576);
or U9461 (N_9461,N_8813,N_8791);
nand U9462 (N_9462,N_8645,N_8512);
nand U9463 (N_9463,N_8383,N_8764);
xor U9464 (N_9464,N_8773,N_8087);
xor U9465 (N_9465,N_8888,N_8130);
or U9466 (N_9466,N_8298,N_8352);
xnor U9467 (N_9467,N_8701,N_8640);
xnor U9468 (N_9468,N_8221,N_8901);
nor U9469 (N_9469,N_8538,N_8610);
xor U9470 (N_9470,N_8799,N_8023);
nand U9471 (N_9471,N_8113,N_8497);
nand U9472 (N_9472,N_8521,N_8313);
or U9473 (N_9473,N_8316,N_8717);
nand U9474 (N_9474,N_8467,N_8322);
and U9475 (N_9475,N_8524,N_8976);
nor U9476 (N_9476,N_8315,N_8123);
nor U9477 (N_9477,N_8462,N_8008);
nor U9478 (N_9478,N_8223,N_8784);
or U9479 (N_9479,N_8393,N_8118);
and U9480 (N_9480,N_8573,N_8614);
xor U9481 (N_9481,N_8285,N_8817);
and U9482 (N_9482,N_8402,N_8814);
nand U9483 (N_9483,N_8054,N_8632);
and U9484 (N_9484,N_8484,N_8388);
and U9485 (N_9485,N_8031,N_8567);
or U9486 (N_9486,N_8935,N_8991);
xor U9487 (N_9487,N_8142,N_8836);
nand U9488 (N_9488,N_8820,N_8955);
nor U9489 (N_9489,N_8871,N_8668);
xnor U9490 (N_9490,N_8308,N_8164);
and U9491 (N_9491,N_8528,N_8878);
xor U9492 (N_9492,N_8408,N_8436);
or U9493 (N_9493,N_8486,N_8033);
or U9494 (N_9494,N_8163,N_8519);
xnor U9495 (N_9495,N_8756,N_8094);
or U9496 (N_9496,N_8718,N_8945);
or U9497 (N_9497,N_8136,N_8630);
or U9498 (N_9498,N_8500,N_8531);
nor U9499 (N_9499,N_8643,N_8924);
or U9500 (N_9500,N_8922,N_8241);
nor U9501 (N_9501,N_8605,N_8541);
nand U9502 (N_9502,N_8409,N_8855);
and U9503 (N_9503,N_8825,N_8932);
xnor U9504 (N_9504,N_8143,N_8770);
xor U9505 (N_9505,N_8122,N_8024);
and U9506 (N_9506,N_8387,N_8324);
and U9507 (N_9507,N_8184,N_8182);
nand U9508 (N_9508,N_8072,N_8521);
or U9509 (N_9509,N_8532,N_8203);
or U9510 (N_9510,N_8505,N_8763);
xor U9511 (N_9511,N_8163,N_8041);
nand U9512 (N_9512,N_8357,N_8643);
xnor U9513 (N_9513,N_8213,N_8387);
xnor U9514 (N_9514,N_8120,N_8299);
and U9515 (N_9515,N_8158,N_8744);
or U9516 (N_9516,N_8460,N_8334);
nand U9517 (N_9517,N_8329,N_8426);
nand U9518 (N_9518,N_8791,N_8679);
nor U9519 (N_9519,N_8832,N_8344);
nor U9520 (N_9520,N_8916,N_8886);
xnor U9521 (N_9521,N_8962,N_8209);
and U9522 (N_9522,N_8721,N_8731);
or U9523 (N_9523,N_8839,N_8053);
xor U9524 (N_9524,N_8885,N_8286);
nor U9525 (N_9525,N_8976,N_8020);
nor U9526 (N_9526,N_8976,N_8044);
xor U9527 (N_9527,N_8729,N_8046);
nor U9528 (N_9528,N_8916,N_8108);
and U9529 (N_9529,N_8599,N_8130);
nand U9530 (N_9530,N_8275,N_8774);
nand U9531 (N_9531,N_8837,N_8288);
nor U9532 (N_9532,N_8802,N_8134);
or U9533 (N_9533,N_8245,N_8757);
or U9534 (N_9534,N_8242,N_8313);
and U9535 (N_9535,N_8482,N_8937);
xnor U9536 (N_9536,N_8933,N_8848);
xor U9537 (N_9537,N_8237,N_8166);
and U9538 (N_9538,N_8634,N_8428);
and U9539 (N_9539,N_8178,N_8876);
xnor U9540 (N_9540,N_8047,N_8214);
and U9541 (N_9541,N_8574,N_8548);
or U9542 (N_9542,N_8290,N_8670);
nand U9543 (N_9543,N_8760,N_8924);
nor U9544 (N_9544,N_8923,N_8402);
or U9545 (N_9545,N_8185,N_8596);
xnor U9546 (N_9546,N_8276,N_8160);
nor U9547 (N_9547,N_8935,N_8164);
nor U9548 (N_9548,N_8514,N_8745);
nor U9549 (N_9549,N_8434,N_8575);
or U9550 (N_9550,N_8493,N_8964);
and U9551 (N_9551,N_8158,N_8426);
or U9552 (N_9552,N_8806,N_8556);
xnor U9553 (N_9553,N_8564,N_8709);
xor U9554 (N_9554,N_8991,N_8875);
and U9555 (N_9555,N_8602,N_8212);
nand U9556 (N_9556,N_8649,N_8123);
nand U9557 (N_9557,N_8876,N_8831);
and U9558 (N_9558,N_8734,N_8442);
or U9559 (N_9559,N_8478,N_8777);
and U9560 (N_9560,N_8845,N_8783);
nor U9561 (N_9561,N_8147,N_8034);
and U9562 (N_9562,N_8460,N_8542);
and U9563 (N_9563,N_8723,N_8290);
nor U9564 (N_9564,N_8580,N_8663);
nand U9565 (N_9565,N_8050,N_8723);
xor U9566 (N_9566,N_8059,N_8563);
xnor U9567 (N_9567,N_8983,N_8180);
nor U9568 (N_9568,N_8475,N_8284);
nor U9569 (N_9569,N_8905,N_8291);
or U9570 (N_9570,N_8307,N_8803);
or U9571 (N_9571,N_8665,N_8047);
xor U9572 (N_9572,N_8374,N_8510);
or U9573 (N_9573,N_8957,N_8164);
nor U9574 (N_9574,N_8273,N_8382);
or U9575 (N_9575,N_8420,N_8607);
nand U9576 (N_9576,N_8651,N_8306);
or U9577 (N_9577,N_8724,N_8599);
xor U9578 (N_9578,N_8638,N_8485);
nor U9579 (N_9579,N_8029,N_8157);
xor U9580 (N_9580,N_8387,N_8805);
nand U9581 (N_9581,N_8764,N_8984);
or U9582 (N_9582,N_8999,N_8930);
nor U9583 (N_9583,N_8451,N_8455);
xor U9584 (N_9584,N_8605,N_8766);
nor U9585 (N_9585,N_8749,N_8083);
nand U9586 (N_9586,N_8869,N_8856);
xor U9587 (N_9587,N_8704,N_8087);
nor U9588 (N_9588,N_8614,N_8598);
nand U9589 (N_9589,N_8908,N_8068);
nor U9590 (N_9590,N_8905,N_8129);
or U9591 (N_9591,N_8743,N_8063);
nor U9592 (N_9592,N_8252,N_8665);
and U9593 (N_9593,N_8797,N_8029);
xor U9594 (N_9594,N_8293,N_8348);
nor U9595 (N_9595,N_8265,N_8425);
and U9596 (N_9596,N_8364,N_8720);
nand U9597 (N_9597,N_8191,N_8150);
or U9598 (N_9598,N_8729,N_8948);
nand U9599 (N_9599,N_8624,N_8383);
xnor U9600 (N_9600,N_8930,N_8135);
and U9601 (N_9601,N_8131,N_8910);
nor U9602 (N_9602,N_8849,N_8537);
nor U9603 (N_9603,N_8993,N_8227);
nor U9604 (N_9604,N_8148,N_8655);
nand U9605 (N_9605,N_8878,N_8468);
xor U9606 (N_9606,N_8781,N_8561);
nor U9607 (N_9607,N_8769,N_8788);
xnor U9608 (N_9608,N_8854,N_8500);
nor U9609 (N_9609,N_8436,N_8608);
and U9610 (N_9610,N_8376,N_8080);
or U9611 (N_9611,N_8857,N_8064);
and U9612 (N_9612,N_8469,N_8135);
or U9613 (N_9613,N_8069,N_8399);
xor U9614 (N_9614,N_8471,N_8653);
nor U9615 (N_9615,N_8075,N_8155);
nand U9616 (N_9616,N_8268,N_8143);
xor U9617 (N_9617,N_8006,N_8149);
xor U9618 (N_9618,N_8363,N_8100);
nor U9619 (N_9619,N_8093,N_8810);
and U9620 (N_9620,N_8691,N_8027);
nand U9621 (N_9621,N_8893,N_8141);
nand U9622 (N_9622,N_8509,N_8790);
nor U9623 (N_9623,N_8321,N_8791);
nor U9624 (N_9624,N_8672,N_8811);
or U9625 (N_9625,N_8694,N_8494);
or U9626 (N_9626,N_8066,N_8974);
xnor U9627 (N_9627,N_8927,N_8923);
nor U9628 (N_9628,N_8459,N_8719);
xnor U9629 (N_9629,N_8654,N_8245);
and U9630 (N_9630,N_8986,N_8174);
nor U9631 (N_9631,N_8546,N_8452);
or U9632 (N_9632,N_8914,N_8686);
nor U9633 (N_9633,N_8275,N_8270);
xor U9634 (N_9634,N_8307,N_8338);
xor U9635 (N_9635,N_8283,N_8854);
or U9636 (N_9636,N_8924,N_8671);
nand U9637 (N_9637,N_8710,N_8093);
nand U9638 (N_9638,N_8162,N_8615);
xor U9639 (N_9639,N_8578,N_8865);
nor U9640 (N_9640,N_8974,N_8364);
nor U9641 (N_9641,N_8267,N_8951);
xnor U9642 (N_9642,N_8636,N_8689);
and U9643 (N_9643,N_8957,N_8002);
nor U9644 (N_9644,N_8606,N_8700);
nor U9645 (N_9645,N_8114,N_8223);
or U9646 (N_9646,N_8185,N_8669);
nor U9647 (N_9647,N_8007,N_8471);
xnor U9648 (N_9648,N_8408,N_8207);
nor U9649 (N_9649,N_8494,N_8346);
and U9650 (N_9650,N_8624,N_8451);
nand U9651 (N_9651,N_8750,N_8338);
xor U9652 (N_9652,N_8402,N_8162);
or U9653 (N_9653,N_8030,N_8355);
xnor U9654 (N_9654,N_8167,N_8337);
or U9655 (N_9655,N_8493,N_8151);
nor U9656 (N_9656,N_8805,N_8605);
nor U9657 (N_9657,N_8132,N_8838);
or U9658 (N_9658,N_8680,N_8944);
xor U9659 (N_9659,N_8207,N_8564);
or U9660 (N_9660,N_8060,N_8886);
xnor U9661 (N_9661,N_8501,N_8302);
or U9662 (N_9662,N_8492,N_8021);
nand U9663 (N_9663,N_8075,N_8214);
or U9664 (N_9664,N_8972,N_8074);
xnor U9665 (N_9665,N_8855,N_8840);
nor U9666 (N_9666,N_8620,N_8322);
xor U9667 (N_9667,N_8482,N_8981);
nand U9668 (N_9668,N_8428,N_8904);
and U9669 (N_9669,N_8682,N_8826);
nand U9670 (N_9670,N_8955,N_8123);
xor U9671 (N_9671,N_8747,N_8796);
or U9672 (N_9672,N_8715,N_8368);
nand U9673 (N_9673,N_8948,N_8649);
nand U9674 (N_9674,N_8159,N_8944);
nor U9675 (N_9675,N_8751,N_8323);
or U9676 (N_9676,N_8703,N_8217);
or U9677 (N_9677,N_8976,N_8179);
nor U9678 (N_9678,N_8500,N_8149);
or U9679 (N_9679,N_8130,N_8251);
or U9680 (N_9680,N_8331,N_8695);
xnor U9681 (N_9681,N_8965,N_8353);
nor U9682 (N_9682,N_8007,N_8674);
xnor U9683 (N_9683,N_8142,N_8335);
nor U9684 (N_9684,N_8344,N_8471);
and U9685 (N_9685,N_8368,N_8042);
or U9686 (N_9686,N_8312,N_8773);
nor U9687 (N_9687,N_8728,N_8455);
nor U9688 (N_9688,N_8861,N_8878);
nand U9689 (N_9689,N_8631,N_8751);
xnor U9690 (N_9690,N_8850,N_8123);
nand U9691 (N_9691,N_8286,N_8723);
nand U9692 (N_9692,N_8262,N_8024);
and U9693 (N_9693,N_8225,N_8378);
or U9694 (N_9694,N_8045,N_8481);
nand U9695 (N_9695,N_8844,N_8466);
or U9696 (N_9696,N_8018,N_8947);
and U9697 (N_9697,N_8765,N_8105);
and U9698 (N_9698,N_8908,N_8590);
nor U9699 (N_9699,N_8328,N_8605);
nor U9700 (N_9700,N_8077,N_8125);
nor U9701 (N_9701,N_8419,N_8030);
and U9702 (N_9702,N_8780,N_8082);
or U9703 (N_9703,N_8765,N_8559);
or U9704 (N_9704,N_8959,N_8436);
nand U9705 (N_9705,N_8710,N_8872);
nand U9706 (N_9706,N_8726,N_8407);
xor U9707 (N_9707,N_8500,N_8894);
xnor U9708 (N_9708,N_8836,N_8440);
or U9709 (N_9709,N_8532,N_8969);
or U9710 (N_9710,N_8467,N_8758);
and U9711 (N_9711,N_8623,N_8819);
or U9712 (N_9712,N_8906,N_8667);
and U9713 (N_9713,N_8315,N_8717);
or U9714 (N_9714,N_8408,N_8834);
nand U9715 (N_9715,N_8218,N_8392);
and U9716 (N_9716,N_8278,N_8555);
nand U9717 (N_9717,N_8062,N_8112);
and U9718 (N_9718,N_8248,N_8583);
or U9719 (N_9719,N_8113,N_8294);
or U9720 (N_9720,N_8551,N_8839);
xnor U9721 (N_9721,N_8543,N_8753);
or U9722 (N_9722,N_8528,N_8894);
and U9723 (N_9723,N_8932,N_8581);
nand U9724 (N_9724,N_8715,N_8234);
xnor U9725 (N_9725,N_8860,N_8373);
and U9726 (N_9726,N_8639,N_8733);
and U9727 (N_9727,N_8452,N_8884);
xnor U9728 (N_9728,N_8651,N_8297);
xnor U9729 (N_9729,N_8306,N_8786);
and U9730 (N_9730,N_8850,N_8477);
and U9731 (N_9731,N_8948,N_8682);
nand U9732 (N_9732,N_8836,N_8428);
and U9733 (N_9733,N_8988,N_8045);
and U9734 (N_9734,N_8312,N_8014);
nand U9735 (N_9735,N_8227,N_8857);
or U9736 (N_9736,N_8711,N_8465);
and U9737 (N_9737,N_8450,N_8335);
and U9738 (N_9738,N_8983,N_8354);
xnor U9739 (N_9739,N_8855,N_8068);
xnor U9740 (N_9740,N_8513,N_8114);
or U9741 (N_9741,N_8480,N_8919);
nor U9742 (N_9742,N_8260,N_8773);
or U9743 (N_9743,N_8323,N_8300);
xnor U9744 (N_9744,N_8025,N_8421);
and U9745 (N_9745,N_8917,N_8216);
nand U9746 (N_9746,N_8248,N_8488);
nand U9747 (N_9747,N_8259,N_8115);
or U9748 (N_9748,N_8585,N_8116);
nand U9749 (N_9749,N_8831,N_8595);
nand U9750 (N_9750,N_8481,N_8465);
nor U9751 (N_9751,N_8075,N_8287);
or U9752 (N_9752,N_8884,N_8343);
nand U9753 (N_9753,N_8062,N_8172);
and U9754 (N_9754,N_8221,N_8544);
nor U9755 (N_9755,N_8174,N_8097);
nor U9756 (N_9756,N_8397,N_8607);
nand U9757 (N_9757,N_8867,N_8026);
xnor U9758 (N_9758,N_8210,N_8438);
xnor U9759 (N_9759,N_8839,N_8088);
xnor U9760 (N_9760,N_8662,N_8034);
and U9761 (N_9761,N_8463,N_8000);
or U9762 (N_9762,N_8515,N_8944);
or U9763 (N_9763,N_8296,N_8586);
nor U9764 (N_9764,N_8018,N_8109);
and U9765 (N_9765,N_8549,N_8319);
nor U9766 (N_9766,N_8863,N_8151);
and U9767 (N_9767,N_8946,N_8498);
xor U9768 (N_9768,N_8358,N_8044);
and U9769 (N_9769,N_8689,N_8823);
nor U9770 (N_9770,N_8365,N_8268);
or U9771 (N_9771,N_8739,N_8190);
xor U9772 (N_9772,N_8556,N_8697);
nand U9773 (N_9773,N_8517,N_8480);
xnor U9774 (N_9774,N_8689,N_8215);
xor U9775 (N_9775,N_8224,N_8832);
xor U9776 (N_9776,N_8232,N_8272);
nand U9777 (N_9777,N_8643,N_8637);
nor U9778 (N_9778,N_8224,N_8893);
and U9779 (N_9779,N_8939,N_8628);
or U9780 (N_9780,N_8932,N_8931);
or U9781 (N_9781,N_8074,N_8213);
xnor U9782 (N_9782,N_8820,N_8337);
nand U9783 (N_9783,N_8301,N_8247);
and U9784 (N_9784,N_8835,N_8813);
xor U9785 (N_9785,N_8798,N_8198);
and U9786 (N_9786,N_8098,N_8477);
or U9787 (N_9787,N_8916,N_8202);
and U9788 (N_9788,N_8953,N_8453);
and U9789 (N_9789,N_8056,N_8717);
xor U9790 (N_9790,N_8523,N_8006);
nor U9791 (N_9791,N_8442,N_8126);
or U9792 (N_9792,N_8374,N_8103);
or U9793 (N_9793,N_8436,N_8186);
xnor U9794 (N_9794,N_8047,N_8227);
nand U9795 (N_9795,N_8685,N_8847);
nand U9796 (N_9796,N_8863,N_8932);
nor U9797 (N_9797,N_8341,N_8885);
nand U9798 (N_9798,N_8661,N_8846);
or U9799 (N_9799,N_8868,N_8443);
nand U9800 (N_9800,N_8431,N_8418);
nor U9801 (N_9801,N_8145,N_8353);
and U9802 (N_9802,N_8184,N_8386);
xnor U9803 (N_9803,N_8089,N_8933);
xnor U9804 (N_9804,N_8411,N_8173);
nand U9805 (N_9805,N_8282,N_8620);
nand U9806 (N_9806,N_8996,N_8367);
nand U9807 (N_9807,N_8955,N_8021);
nand U9808 (N_9808,N_8269,N_8555);
nand U9809 (N_9809,N_8452,N_8209);
or U9810 (N_9810,N_8414,N_8444);
xor U9811 (N_9811,N_8481,N_8758);
xor U9812 (N_9812,N_8342,N_8641);
nor U9813 (N_9813,N_8611,N_8979);
nor U9814 (N_9814,N_8360,N_8068);
xnor U9815 (N_9815,N_8452,N_8230);
nand U9816 (N_9816,N_8045,N_8218);
nand U9817 (N_9817,N_8233,N_8765);
nand U9818 (N_9818,N_8931,N_8502);
and U9819 (N_9819,N_8156,N_8677);
nand U9820 (N_9820,N_8325,N_8390);
or U9821 (N_9821,N_8431,N_8731);
xnor U9822 (N_9822,N_8305,N_8118);
or U9823 (N_9823,N_8989,N_8227);
xnor U9824 (N_9824,N_8365,N_8133);
and U9825 (N_9825,N_8585,N_8066);
or U9826 (N_9826,N_8669,N_8055);
xor U9827 (N_9827,N_8100,N_8357);
xor U9828 (N_9828,N_8143,N_8431);
nor U9829 (N_9829,N_8955,N_8459);
nand U9830 (N_9830,N_8413,N_8845);
or U9831 (N_9831,N_8939,N_8925);
or U9832 (N_9832,N_8560,N_8610);
nand U9833 (N_9833,N_8649,N_8880);
nand U9834 (N_9834,N_8557,N_8097);
xnor U9835 (N_9835,N_8095,N_8368);
nor U9836 (N_9836,N_8114,N_8024);
or U9837 (N_9837,N_8752,N_8437);
xnor U9838 (N_9838,N_8276,N_8430);
and U9839 (N_9839,N_8493,N_8534);
and U9840 (N_9840,N_8215,N_8494);
xnor U9841 (N_9841,N_8574,N_8611);
nor U9842 (N_9842,N_8697,N_8261);
and U9843 (N_9843,N_8646,N_8520);
nor U9844 (N_9844,N_8965,N_8404);
nor U9845 (N_9845,N_8745,N_8022);
xor U9846 (N_9846,N_8327,N_8430);
nand U9847 (N_9847,N_8344,N_8845);
and U9848 (N_9848,N_8095,N_8418);
and U9849 (N_9849,N_8563,N_8755);
nor U9850 (N_9850,N_8881,N_8698);
xnor U9851 (N_9851,N_8586,N_8273);
nor U9852 (N_9852,N_8348,N_8824);
and U9853 (N_9853,N_8278,N_8751);
nor U9854 (N_9854,N_8866,N_8737);
and U9855 (N_9855,N_8395,N_8003);
nand U9856 (N_9856,N_8858,N_8937);
or U9857 (N_9857,N_8703,N_8757);
or U9858 (N_9858,N_8825,N_8216);
xnor U9859 (N_9859,N_8181,N_8306);
or U9860 (N_9860,N_8409,N_8296);
and U9861 (N_9861,N_8564,N_8350);
or U9862 (N_9862,N_8040,N_8524);
xor U9863 (N_9863,N_8599,N_8810);
nand U9864 (N_9864,N_8684,N_8719);
xor U9865 (N_9865,N_8610,N_8516);
nand U9866 (N_9866,N_8341,N_8311);
and U9867 (N_9867,N_8364,N_8470);
xor U9868 (N_9868,N_8347,N_8649);
nor U9869 (N_9869,N_8459,N_8701);
and U9870 (N_9870,N_8700,N_8656);
or U9871 (N_9871,N_8639,N_8936);
xnor U9872 (N_9872,N_8235,N_8678);
xor U9873 (N_9873,N_8622,N_8610);
nand U9874 (N_9874,N_8740,N_8829);
nor U9875 (N_9875,N_8517,N_8370);
nand U9876 (N_9876,N_8821,N_8289);
and U9877 (N_9877,N_8164,N_8817);
nor U9878 (N_9878,N_8895,N_8453);
xnor U9879 (N_9879,N_8672,N_8526);
xor U9880 (N_9880,N_8974,N_8954);
nand U9881 (N_9881,N_8026,N_8229);
xnor U9882 (N_9882,N_8904,N_8230);
or U9883 (N_9883,N_8915,N_8077);
or U9884 (N_9884,N_8402,N_8698);
and U9885 (N_9885,N_8054,N_8882);
xor U9886 (N_9886,N_8985,N_8618);
xnor U9887 (N_9887,N_8233,N_8408);
or U9888 (N_9888,N_8850,N_8024);
nor U9889 (N_9889,N_8973,N_8400);
or U9890 (N_9890,N_8302,N_8315);
nand U9891 (N_9891,N_8731,N_8154);
or U9892 (N_9892,N_8828,N_8972);
nand U9893 (N_9893,N_8827,N_8177);
nand U9894 (N_9894,N_8475,N_8756);
and U9895 (N_9895,N_8871,N_8794);
nand U9896 (N_9896,N_8294,N_8965);
nor U9897 (N_9897,N_8905,N_8328);
or U9898 (N_9898,N_8874,N_8345);
xnor U9899 (N_9899,N_8565,N_8221);
nand U9900 (N_9900,N_8735,N_8273);
nor U9901 (N_9901,N_8140,N_8261);
or U9902 (N_9902,N_8725,N_8183);
and U9903 (N_9903,N_8280,N_8646);
xnor U9904 (N_9904,N_8581,N_8894);
or U9905 (N_9905,N_8682,N_8006);
nor U9906 (N_9906,N_8938,N_8454);
and U9907 (N_9907,N_8965,N_8197);
or U9908 (N_9908,N_8160,N_8125);
nor U9909 (N_9909,N_8554,N_8286);
xnor U9910 (N_9910,N_8406,N_8078);
nor U9911 (N_9911,N_8771,N_8118);
and U9912 (N_9912,N_8000,N_8010);
and U9913 (N_9913,N_8616,N_8082);
and U9914 (N_9914,N_8928,N_8204);
nor U9915 (N_9915,N_8748,N_8643);
or U9916 (N_9916,N_8091,N_8639);
and U9917 (N_9917,N_8737,N_8103);
or U9918 (N_9918,N_8182,N_8208);
and U9919 (N_9919,N_8154,N_8629);
nand U9920 (N_9920,N_8413,N_8348);
nand U9921 (N_9921,N_8047,N_8609);
xnor U9922 (N_9922,N_8093,N_8910);
and U9923 (N_9923,N_8750,N_8927);
nand U9924 (N_9924,N_8782,N_8014);
xor U9925 (N_9925,N_8576,N_8289);
nand U9926 (N_9926,N_8526,N_8488);
or U9927 (N_9927,N_8823,N_8198);
or U9928 (N_9928,N_8302,N_8942);
nand U9929 (N_9929,N_8268,N_8251);
nand U9930 (N_9930,N_8729,N_8452);
or U9931 (N_9931,N_8214,N_8253);
nor U9932 (N_9932,N_8868,N_8957);
xor U9933 (N_9933,N_8509,N_8783);
nor U9934 (N_9934,N_8494,N_8127);
nor U9935 (N_9935,N_8940,N_8490);
and U9936 (N_9936,N_8101,N_8653);
or U9937 (N_9937,N_8045,N_8347);
nand U9938 (N_9938,N_8716,N_8738);
nand U9939 (N_9939,N_8635,N_8692);
and U9940 (N_9940,N_8527,N_8445);
nand U9941 (N_9941,N_8491,N_8939);
nor U9942 (N_9942,N_8216,N_8631);
nor U9943 (N_9943,N_8567,N_8396);
or U9944 (N_9944,N_8955,N_8748);
or U9945 (N_9945,N_8181,N_8270);
nand U9946 (N_9946,N_8842,N_8923);
nor U9947 (N_9947,N_8502,N_8777);
nor U9948 (N_9948,N_8634,N_8240);
or U9949 (N_9949,N_8529,N_8955);
nand U9950 (N_9950,N_8056,N_8839);
nor U9951 (N_9951,N_8752,N_8548);
xnor U9952 (N_9952,N_8497,N_8802);
nor U9953 (N_9953,N_8435,N_8450);
or U9954 (N_9954,N_8766,N_8573);
or U9955 (N_9955,N_8441,N_8722);
nor U9956 (N_9956,N_8882,N_8747);
nand U9957 (N_9957,N_8913,N_8115);
nor U9958 (N_9958,N_8099,N_8061);
or U9959 (N_9959,N_8666,N_8198);
nand U9960 (N_9960,N_8045,N_8380);
or U9961 (N_9961,N_8220,N_8500);
and U9962 (N_9962,N_8362,N_8175);
nor U9963 (N_9963,N_8367,N_8036);
or U9964 (N_9964,N_8665,N_8343);
or U9965 (N_9965,N_8511,N_8084);
nand U9966 (N_9966,N_8517,N_8591);
or U9967 (N_9967,N_8505,N_8841);
xnor U9968 (N_9968,N_8527,N_8337);
and U9969 (N_9969,N_8450,N_8724);
nand U9970 (N_9970,N_8262,N_8093);
xor U9971 (N_9971,N_8165,N_8179);
xnor U9972 (N_9972,N_8257,N_8694);
and U9973 (N_9973,N_8504,N_8266);
or U9974 (N_9974,N_8091,N_8234);
nand U9975 (N_9975,N_8924,N_8915);
or U9976 (N_9976,N_8424,N_8645);
xor U9977 (N_9977,N_8302,N_8065);
xnor U9978 (N_9978,N_8285,N_8270);
xor U9979 (N_9979,N_8485,N_8942);
xor U9980 (N_9980,N_8822,N_8272);
nor U9981 (N_9981,N_8534,N_8505);
nand U9982 (N_9982,N_8117,N_8616);
and U9983 (N_9983,N_8642,N_8991);
xor U9984 (N_9984,N_8027,N_8800);
xor U9985 (N_9985,N_8428,N_8553);
nand U9986 (N_9986,N_8810,N_8291);
nand U9987 (N_9987,N_8362,N_8243);
xor U9988 (N_9988,N_8153,N_8611);
or U9989 (N_9989,N_8840,N_8258);
nand U9990 (N_9990,N_8021,N_8659);
xnor U9991 (N_9991,N_8523,N_8200);
nor U9992 (N_9992,N_8035,N_8204);
nand U9993 (N_9993,N_8332,N_8327);
nor U9994 (N_9994,N_8591,N_8083);
and U9995 (N_9995,N_8785,N_8201);
or U9996 (N_9996,N_8956,N_8408);
and U9997 (N_9997,N_8767,N_8254);
or U9998 (N_9998,N_8616,N_8527);
xnor U9999 (N_9999,N_8715,N_8596);
nor UO_0 (O_0,N_9702,N_9994);
nand UO_1 (O_1,N_9492,N_9787);
nor UO_2 (O_2,N_9350,N_9860);
and UO_3 (O_3,N_9916,N_9739);
nor UO_4 (O_4,N_9871,N_9631);
nor UO_5 (O_5,N_9719,N_9093);
and UO_6 (O_6,N_9861,N_9896);
nand UO_7 (O_7,N_9346,N_9001);
or UO_8 (O_8,N_9008,N_9418);
nand UO_9 (O_9,N_9309,N_9666);
nand UO_10 (O_10,N_9813,N_9143);
or UO_11 (O_11,N_9943,N_9213);
xor UO_12 (O_12,N_9215,N_9433);
nand UO_13 (O_13,N_9645,N_9487);
nor UO_14 (O_14,N_9032,N_9048);
or UO_15 (O_15,N_9327,N_9180);
xor UO_16 (O_16,N_9133,N_9386);
or UO_17 (O_17,N_9512,N_9184);
nand UO_18 (O_18,N_9582,N_9162);
nand UO_19 (O_19,N_9108,N_9928);
nand UO_20 (O_20,N_9357,N_9091);
or UO_21 (O_21,N_9891,N_9892);
nand UO_22 (O_22,N_9971,N_9038);
or UO_23 (O_23,N_9681,N_9980);
xor UO_24 (O_24,N_9097,N_9769);
or UO_25 (O_25,N_9453,N_9991);
xnor UO_26 (O_26,N_9363,N_9583);
and UO_27 (O_27,N_9717,N_9584);
nand UO_28 (O_28,N_9572,N_9904);
or UO_29 (O_29,N_9339,N_9912);
and UO_30 (O_30,N_9560,N_9260);
and UO_31 (O_31,N_9706,N_9758);
and UO_32 (O_32,N_9555,N_9367);
nor UO_33 (O_33,N_9444,N_9765);
xor UO_34 (O_34,N_9039,N_9410);
xnor UO_35 (O_35,N_9018,N_9581);
xnor UO_36 (O_36,N_9428,N_9277);
and UO_37 (O_37,N_9158,N_9883);
and UO_38 (O_38,N_9882,N_9227);
xnor UO_39 (O_39,N_9297,N_9618);
nand UO_40 (O_40,N_9710,N_9520);
nand UO_41 (O_41,N_9399,N_9374);
or UO_42 (O_42,N_9165,N_9379);
nand UO_43 (O_43,N_9821,N_9562);
or UO_44 (O_44,N_9371,N_9960);
nand UO_45 (O_45,N_9142,N_9894);
nand UO_46 (O_46,N_9907,N_9089);
and UO_47 (O_47,N_9629,N_9154);
xor UO_48 (O_48,N_9647,N_9638);
and UO_49 (O_49,N_9836,N_9544);
nand UO_50 (O_50,N_9848,N_9785);
nand UO_51 (O_51,N_9347,N_9000);
nor UO_52 (O_52,N_9780,N_9847);
and UO_53 (O_53,N_9941,N_9221);
xnor UO_54 (O_54,N_9087,N_9147);
nor UO_55 (O_55,N_9470,N_9968);
xor UO_56 (O_56,N_9812,N_9875);
nand UO_57 (O_57,N_9569,N_9852);
nor UO_58 (O_58,N_9306,N_9380);
xnor UO_59 (O_59,N_9020,N_9494);
nand UO_60 (O_60,N_9263,N_9173);
nor UO_61 (O_61,N_9043,N_9876);
nand UO_62 (O_62,N_9974,N_9617);
nand UO_63 (O_63,N_9660,N_9778);
or UO_64 (O_64,N_9044,N_9767);
xnor UO_65 (O_65,N_9151,N_9519);
and UO_66 (O_66,N_9257,N_9217);
nand UO_67 (O_67,N_9922,N_9388);
xnor UO_68 (O_68,N_9612,N_9402);
nor UO_69 (O_69,N_9017,N_9712);
nor UO_70 (O_70,N_9908,N_9580);
or UO_71 (O_71,N_9952,N_9164);
and UO_72 (O_72,N_9823,N_9850);
and UO_73 (O_73,N_9329,N_9766);
nor UO_74 (O_74,N_9438,N_9851);
and UO_75 (O_75,N_9929,N_9226);
nor UO_76 (O_76,N_9536,N_9628);
nand UO_77 (O_77,N_9294,N_9935);
xnor UO_78 (O_78,N_9366,N_9268);
nor UO_79 (O_79,N_9969,N_9161);
xor UO_80 (O_80,N_9220,N_9101);
or UO_81 (O_81,N_9095,N_9579);
and UO_82 (O_82,N_9114,N_9381);
nor UO_83 (O_83,N_9116,N_9862);
and UO_84 (O_84,N_9118,N_9281);
xor UO_85 (O_85,N_9282,N_9689);
or UO_86 (O_86,N_9325,N_9256);
or UO_87 (O_87,N_9732,N_9255);
nor UO_88 (O_88,N_9878,N_9760);
or UO_89 (O_89,N_9564,N_9976);
or UO_90 (O_90,N_9066,N_9397);
or UO_91 (O_91,N_9063,N_9687);
or UO_92 (O_92,N_9547,N_9352);
nand UO_93 (O_93,N_9334,N_9978);
nor UO_94 (O_94,N_9696,N_9197);
xor UO_95 (O_95,N_9383,N_9167);
xnor UO_96 (O_96,N_9324,N_9214);
and UO_97 (O_97,N_9679,N_9201);
nor UO_98 (O_98,N_9231,N_9313);
nand UO_99 (O_99,N_9172,N_9182);
nand UO_100 (O_100,N_9648,N_9073);
nor UO_101 (O_101,N_9740,N_9503);
or UO_102 (O_102,N_9469,N_9678);
or UO_103 (O_103,N_9455,N_9665);
nor UO_104 (O_104,N_9387,N_9448);
or UO_105 (O_105,N_9736,N_9077);
nand UO_106 (O_106,N_9181,N_9975);
xnor UO_107 (O_107,N_9566,N_9450);
and UO_108 (O_108,N_9752,N_9734);
nand UO_109 (O_109,N_9274,N_9565);
or UO_110 (O_110,N_9844,N_9075);
xnor UO_111 (O_111,N_9651,N_9452);
or UO_112 (O_112,N_9152,N_9890);
and UO_113 (O_113,N_9989,N_9171);
nor UO_114 (O_114,N_9996,N_9559);
xor UO_115 (O_115,N_9859,N_9676);
xor UO_116 (O_116,N_9258,N_9131);
xnor UO_117 (O_117,N_9473,N_9576);
xor UO_118 (O_118,N_9528,N_9405);
or UO_119 (O_119,N_9065,N_9482);
nand UO_120 (O_120,N_9510,N_9998);
xor UO_121 (O_121,N_9385,N_9242);
nor UO_122 (O_122,N_9872,N_9749);
and UO_123 (O_123,N_9634,N_9834);
xnor UO_124 (O_124,N_9695,N_9003);
or UO_125 (O_125,N_9030,N_9360);
nor UO_126 (O_126,N_9982,N_9076);
or UO_127 (O_127,N_9772,N_9814);
nand UO_128 (O_128,N_9791,N_9499);
nor UO_129 (O_129,N_9977,N_9248);
nor UO_130 (O_130,N_9556,N_9625);
or UO_131 (O_131,N_9176,N_9301);
nor UO_132 (O_132,N_9642,N_9506);
and UO_133 (O_133,N_9323,N_9392);
xnor UO_134 (O_134,N_9445,N_9305);
and UO_135 (O_135,N_9016,N_9229);
nor UO_136 (O_136,N_9238,N_9831);
nor UO_137 (O_137,N_9285,N_9790);
nand UO_138 (O_138,N_9839,N_9720);
nor UO_139 (O_139,N_9303,N_9054);
and UO_140 (O_140,N_9315,N_9549);
xnor UO_141 (O_141,N_9004,N_9269);
nor UO_142 (O_142,N_9150,N_9902);
xor UO_143 (O_143,N_9080,N_9832);
and UO_144 (O_144,N_9110,N_9439);
nand UO_145 (O_145,N_9573,N_9022);
or UO_146 (O_146,N_9825,N_9403);
or UO_147 (O_147,N_9845,N_9531);
or UO_148 (O_148,N_9328,N_9125);
nor UO_149 (O_149,N_9391,N_9726);
nand UO_150 (O_150,N_9923,N_9465);
nor UO_151 (O_151,N_9613,N_9755);
nand UO_152 (O_152,N_9746,N_9295);
nor UO_153 (O_153,N_9225,N_9046);
xor UO_154 (O_154,N_9422,N_9062);
and UO_155 (O_155,N_9486,N_9762);
nand UO_156 (O_156,N_9824,N_9290);
xnor UO_157 (O_157,N_9965,N_9316);
xor UO_158 (O_158,N_9525,N_9098);
and UO_159 (O_159,N_9312,N_9743);
and UO_160 (O_160,N_9854,N_9219);
or UO_161 (O_161,N_9774,N_9731);
or UO_162 (O_162,N_9052,N_9885);
xnor UO_163 (O_163,N_9906,N_9668);
and UO_164 (O_164,N_9649,N_9079);
and UO_165 (O_165,N_9764,N_9588);
or UO_166 (O_166,N_9267,N_9788);
nand UO_167 (O_167,N_9619,N_9507);
or UO_168 (O_168,N_9136,N_9776);
and UO_169 (O_169,N_9443,N_9815);
xnor UO_170 (O_170,N_9050,N_9423);
and UO_171 (O_171,N_9139,N_9011);
and UO_172 (O_172,N_9659,N_9886);
and UO_173 (O_173,N_9345,N_9972);
and UO_174 (O_174,N_9092,N_9090);
or UO_175 (O_175,N_9128,N_9661);
and UO_176 (O_176,N_9500,N_9368);
nor UO_177 (O_177,N_9446,N_9840);
and UO_178 (O_178,N_9911,N_9930);
nand UO_179 (O_179,N_9343,N_9551);
nor UO_180 (O_180,N_9511,N_9479);
xnor UO_181 (O_181,N_9212,N_9468);
or UO_182 (O_182,N_9166,N_9817);
nor UO_183 (O_183,N_9207,N_9477);
or UO_184 (O_184,N_9460,N_9222);
xor UO_185 (O_185,N_9698,N_9396);
nand UO_186 (O_186,N_9624,N_9750);
xnor UO_187 (O_187,N_9027,N_9598);
and UO_188 (O_188,N_9157,N_9252);
and UO_189 (O_189,N_9957,N_9149);
nor UO_190 (O_190,N_9307,N_9849);
nand UO_191 (O_191,N_9447,N_9311);
or UO_192 (O_192,N_9250,N_9632);
nand UO_193 (O_193,N_9737,N_9842);
or UO_194 (O_194,N_9170,N_9120);
xor UO_195 (O_195,N_9714,N_9070);
or UO_196 (O_196,N_9072,N_9721);
xnor UO_197 (O_197,N_9300,N_9081);
nand UO_198 (O_198,N_9672,N_9763);
and UO_199 (O_199,N_9035,N_9026);
nand UO_200 (O_200,N_9915,N_9997);
nor UO_201 (O_201,N_9454,N_9199);
nand UO_202 (O_202,N_9057,N_9663);
nand UO_203 (O_203,N_9554,N_9987);
or UO_204 (O_204,N_9389,N_9354);
xnor UO_205 (O_205,N_9086,N_9241);
and UO_206 (O_206,N_9779,N_9570);
nor UO_207 (O_207,N_9270,N_9708);
nand UO_208 (O_208,N_9962,N_9140);
nor UO_209 (O_209,N_9798,N_9527);
and UO_210 (O_210,N_9693,N_9561);
or UO_211 (O_211,N_9761,N_9633);
xnor UO_212 (O_212,N_9053,N_9417);
nor UO_213 (O_213,N_9627,N_9349);
and UO_214 (O_214,N_9273,N_9811);
xnor UO_215 (O_215,N_9146,N_9456);
and UO_216 (O_216,N_9218,N_9266);
nor UO_217 (O_217,N_9203,N_9333);
nand UO_218 (O_218,N_9942,N_9833);
xor UO_219 (O_219,N_9803,N_9376);
or UO_220 (O_220,N_9276,N_9042);
xor UO_221 (O_221,N_9863,N_9424);
xnor UO_222 (O_222,N_9175,N_9014);
nand UO_223 (O_223,N_9132,N_9129);
and UO_224 (O_224,N_9567,N_9233);
and UO_225 (O_225,N_9759,N_9085);
nor UO_226 (O_226,N_9356,N_9185);
and UO_227 (O_227,N_9667,N_9918);
and UO_228 (O_228,N_9190,N_9684);
and UO_229 (O_229,N_9671,N_9488);
nor UO_230 (O_230,N_9464,N_9728);
and UO_231 (O_231,N_9459,N_9291);
xor UO_232 (O_232,N_9523,N_9010);
nand UO_233 (O_233,N_9186,N_9228);
nand UO_234 (O_234,N_9718,N_9864);
and UO_235 (O_235,N_9163,N_9279);
nand UO_236 (O_236,N_9262,N_9105);
and UO_237 (O_237,N_9202,N_9206);
and UO_238 (O_238,N_9375,N_9103);
and UO_239 (O_239,N_9783,N_9781);
nand UO_240 (O_240,N_9558,N_9489);
nor UO_241 (O_241,N_9112,N_9733);
xnor UO_242 (O_242,N_9571,N_9058);
xor UO_243 (O_243,N_9302,N_9292);
xor UO_244 (O_244,N_9934,N_9382);
xnor UO_245 (O_245,N_9881,N_9592);
nand UO_246 (O_246,N_9056,N_9594);
and UO_247 (O_247,N_9156,N_9115);
nand UO_248 (O_248,N_9611,N_9951);
xor UO_249 (O_249,N_9209,N_9111);
and UO_250 (O_250,N_9135,N_9589);
and UO_251 (O_251,N_9514,N_9694);
nand UO_252 (O_252,N_9153,N_9843);
and UO_253 (O_253,N_9947,N_9716);
nor UO_254 (O_254,N_9421,N_9137);
xor UO_255 (O_255,N_9546,N_9436);
nor UO_256 (O_256,N_9574,N_9770);
nand UO_257 (O_257,N_9378,N_9462);
xnor UO_258 (O_258,N_9361,N_9094);
nor UO_259 (O_259,N_9786,N_9853);
nand UO_260 (O_260,N_9705,N_9319);
nand UO_261 (O_261,N_9472,N_9330);
nor UO_262 (O_262,N_9401,N_9868);
xor UO_263 (O_263,N_9703,N_9419);
or UO_264 (O_264,N_9795,N_9837);
xor UO_265 (O_265,N_9099,N_9485);
nand UO_266 (O_266,N_9899,N_9901);
and UO_267 (O_267,N_9874,N_9995);
xor UO_268 (O_268,N_9529,N_9686);
nor UO_269 (O_269,N_9355,N_9800);
nand UO_270 (O_270,N_9299,N_9002);
and UO_271 (O_271,N_9920,N_9953);
nor UO_272 (O_272,N_9321,N_9078);
or UO_273 (O_273,N_9936,N_9502);
nor UO_274 (O_274,N_9068,N_9320);
xnor UO_275 (O_275,N_9964,N_9024);
and UO_276 (O_276,N_9169,N_9373);
and UO_277 (O_277,N_9365,N_9621);
xor UO_278 (O_278,N_9508,N_9289);
or UO_279 (O_279,N_9013,N_9816);
xnor UO_280 (O_280,N_9984,N_9753);
nand UO_281 (O_281,N_9545,N_9474);
and UO_282 (O_282,N_9318,N_9707);
nor UO_283 (O_283,N_9692,N_9557);
xnor UO_284 (O_284,N_9657,N_9272);
nor UO_285 (O_285,N_9775,N_9993);
nand UO_286 (O_286,N_9884,N_9496);
and UO_287 (O_287,N_9275,N_9516);
xor UO_288 (O_288,N_9467,N_9160);
xor UO_289 (O_289,N_9999,N_9005);
nand UO_290 (O_290,N_9799,N_9179);
nor UO_291 (O_291,N_9973,N_9449);
and UO_292 (O_292,N_9045,N_9603);
or UO_293 (O_293,N_9606,N_9709);
xnor UO_294 (O_294,N_9919,N_9533);
and UO_295 (O_295,N_9713,N_9015);
nand UO_296 (O_296,N_9988,N_9568);
nor UO_297 (O_297,N_9126,N_9623);
or UO_298 (O_298,N_9841,N_9521);
xnor UO_299 (O_299,N_9518,N_9096);
nand UO_300 (O_300,N_9959,N_9127);
xnor UO_301 (O_301,N_9548,N_9029);
xnor UO_302 (O_302,N_9602,N_9596);
nand UO_303 (O_303,N_9782,N_9827);
or UO_304 (O_304,N_9244,N_9264);
xnor UO_305 (O_305,N_9434,N_9283);
nand UO_306 (O_306,N_9425,N_9828);
and UO_307 (O_307,N_9682,N_9522);
and UO_308 (O_308,N_9019,N_9543);
and UO_309 (O_309,N_9240,N_9491);
xor UO_310 (O_310,N_9187,N_9051);
or UO_311 (O_311,N_9287,N_9517);
or UO_312 (O_312,N_9178,N_9654);
nor UO_313 (O_313,N_9061,N_9646);
and UO_314 (O_314,N_9441,N_9963);
and UO_315 (O_315,N_9278,N_9138);
or UO_316 (O_316,N_9806,N_9680);
or UO_317 (O_317,N_9622,N_9483);
or UO_318 (O_318,N_9513,N_9223);
or UO_319 (O_319,N_9009,N_9064);
nand UO_320 (O_320,N_9643,N_9747);
nor UO_321 (O_321,N_9829,N_9208);
nor UO_322 (O_322,N_9701,N_9107);
xor UO_323 (O_323,N_9802,N_9204);
nor UO_324 (O_324,N_9652,N_9322);
xnor UO_325 (O_325,N_9336,N_9990);
xor UO_326 (O_326,N_9249,N_9243);
nand UO_327 (O_327,N_9711,N_9630);
nand UO_328 (O_328,N_9025,N_9768);
nor UO_329 (O_329,N_9082,N_9910);
and UO_330 (O_330,N_9905,N_9605);
or UO_331 (O_331,N_9597,N_9192);
nand UO_332 (O_332,N_9950,N_9794);
nor UO_333 (O_333,N_9777,N_9420);
nor UO_334 (O_334,N_9461,N_9614);
xor UO_335 (O_335,N_9636,N_9535);
and UO_336 (O_336,N_9879,N_9286);
nand UO_337 (O_337,N_9463,N_9804);
or UO_338 (O_338,N_9432,N_9939);
nor UO_339 (O_339,N_9640,N_9235);
nor UO_340 (O_340,N_9563,N_9210);
and UO_341 (O_341,N_9577,N_9600);
xnor UO_342 (O_342,N_9189,N_9616);
nor UO_343 (O_343,N_9195,N_9741);
or UO_344 (O_344,N_9818,N_9801);
and UO_345 (O_345,N_9415,N_9900);
nor UO_346 (O_346,N_9855,N_9748);
or UO_347 (O_347,N_9877,N_9835);
nor UO_348 (O_348,N_9404,N_9261);
nand UO_349 (O_349,N_9917,N_9493);
nor UO_350 (O_350,N_9134,N_9384);
nand UO_351 (O_351,N_9954,N_9595);
and UO_352 (O_352,N_9615,N_9442);
xnor UO_353 (O_353,N_9590,N_9183);
nand UO_354 (O_354,N_9921,N_9955);
nand UO_355 (O_355,N_9610,N_9585);
nand UO_356 (O_356,N_9858,N_9067);
xor UO_357 (O_357,N_9124,N_9893);
nor UO_358 (O_358,N_9236,N_9427);
or UO_359 (O_359,N_9055,N_9807);
xnor UO_360 (O_360,N_9575,N_9887);
nor UO_361 (O_361,N_9604,N_9102);
or UO_362 (O_362,N_9414,N_9224);
nor UO_363 (O_363,N_9838,N_9792);
nand UO_364 (O_364,N_9377,N_9700);
or UO_365 (O_365,N_9898,N_9412);
nor UO_366 (O_366,N_9395,N_9370);
nor UO_367 (O_367,N_9234,N_9981);
nand UO_368 (O_368,N_9155,N_9451);
xor UO_369 (O_369,N_9476,N_9431);
or UO_370 (O_370,N_9498,N_9593);
nor UO_371 (O_371,N_9406,N_9239);
or UO_372 (O_372,N_9109,N_9515);
nor UO_373 (O_373,N_9819,N_9797);
and UO_374 (O_374,N_9599,N_9538);
nor UO_375 (O_375,N_9074,N_9756);
or UO_376 (O_376,N_9130,N_9541);
xnor UO_377 (O_377,N_9738,N_9314);
or UO_378 (O_378,N_9931,N_9552);
nor UO_379 (O_379,N_9369,N_9047);
nand UO_380 (O_380,N_9106,N_9232);
and UO_381 (O_381,N_9690,N_9344);
and UO_382 (O_382,N_9331,N_9673);
nand UO_383 (O_383,N_9724,N_9656);
nand UO_384 (O_384,N_9637,N_9036);
or UO_385 (O_385,N_9591,N_9730);
nor UO_386 (O_386,N_9337,N_9340);
and UO_387 (O_387,N_9495,N_9725);
and UO_388 (O_388,N_9644,N_9805);
nand UO_389 (O_389,N_9609,N_9587);
xnor UO_390 (O_390,N_9104,N_9037);
xor UO_391 (O_391,N_9359,N_9122);
nor UO_392 (O_392,N_9534,N_9946);
and UO_393 (O_393,N_9809,N_9254);
nor UO_394 (O_394,N_9196,N_9857);
nand UO_395 (O_395,N_9727,N_9177);
nand UO_396 (O_396,N_9967,N_9691);
nand UO_397 (O_397,N_9924,N_9413);
and UO_398 (O_398,N_9400,N_9826);
nor UO_399 (O_399,N_9174,N_9490);
xnor UO_400 (O_400,N_9932,N_9084);
nor UO_401 (O_401,N_9117,N_9230);
and UO_402 (O_402,N_9793,N_9251);
and UO_403 (O_403,N_9664,N_9237);
and UO_404 (O_404,N_9979,N_9856);
nand UO_405 (O_405,N_9144,N_9280);
and UO_406 (O_406,N_9754,N_9407);
xnor UO_407 (O_407,N_9437,N_9398);
xor UO_408 (O_408,N_9674,N_9944);
and UO_409 (O_409,N_9820,N_9509);
xnor UO_410 (O_410,N_9745,N_9986);
nor UO_411 (O_411,N_9430,N_9970);
xor UO_412 (O_412,N_9796,N_9478);
and UO_413 (O_413,N_9317,N_9296);
and UO_414 (O_414,N_9524,N_9586);
nor UO_415 (O_415,N_9480,N_9626);
nor UO_416 (O_416,N_9897,N_9246);
nand UO_417 (O_417,N_9332,N_9159);
and UO_418 (O_418,N_9466,N_9608);
nor UO_419 (O_419,N_9956,N_9961);
or UO_420 (O_420,N_9639,N_9675);
nor UO_421 (O_421,N_9945,N_9023);
nand UO_422 (O_422,N_9457,N_9688);
or UO_423 (O_423,N_9670,N_9537);
nand UO_424 (O_424,N_9416,N_9411);
nor UO_425 (O_425,N_9033,N_9992);
and UO_426 (O_426,N_9429,N_9677);
nand UO_427 (O_427,N_9723,N_9846);
or UO_428 (O_428,N_9088,N_9869);
nor UO_429 (O_429,N_9194,N_9685);
nand UO_430 (O_430,N_9007,N_9284);
nand UO_431 (O_431,N_9607,N_9650);
nor UO_432 (O_432,N_9168,N_9049);
nor UO_433 (O_433,N_9342,N_9658);
nand UO_434 (O_434,N_9578,N_9394);
nor UO_435 (O_435,N_9426,N_9071);
or UO_436 (O_436,N_9926,N_9259);
nand UO_437 (O_437,N_9867,N_9925);
xnor UO_438 (O_438,N_9504,N_9310);
or UO_439 (O_439,N_9123,N_9880);
and UO_440 (O_440,N_9913,N_9830);
nand UO_441 (O_441,N_9353,N_9505);
and UO_442 (O_442,N_9408,N_9021);
and UO_443 (O_443,N_9873,N_9784);
xnor UO_444 (O_444,N_9121,N_9532);
nor UO_445 (O_445,N_9245,N_9773);
nor UO_446 (O_446,N_9041,N_9810);
nor UO_447 (O_447,N_9949,N_9145);
nand UO_448 (O_448,N_9870,N_9440);
and UO_449 (O_449,N_9205,N_9966);
xor UO_450 (O_450,N_9895,N_9914);
nand UO_451 (O_451,N_9028,N_9715);
nor UO_452 (O_452,N_9100,N_9113);
xnor UO_453 (O_453,N_9553,N_9697);
xor UO_454 (O_454,N_9348,N_9662);
xor UO_455 (O_455,N_9435,N_9751);
xor UO_456 (O_456,N_9742,N_9338);
xnor UO_457 (O_457,N_9481,N_9484);
nor UO_458 (O_458,N_9034,N_9358);
nor UO_459 (O_459,N_9983,N_9308);
or UO_460 (O_460,N_9335,N_9635);
xor UO_461 (O_461,N_9069,N_9191);
nand UO_462 (O_462,N_9937,N_9958);
or UO_463 (O_463,N_9744,N_9542);
or UO_464 (O_464,N_9304,N_9940);
xnor UO_465 (O_465,N_9866,N_9059);
or UO_466 (O_466,N_9247,N_9735);
nand UO_467 (O_467,N_9550,N_9601);
nand UO_468 (O_468,N_9141,N_9471);
or UO_469 (O_469,N_9497,N_9351);
xnor UO_470 (O_470,N_9188,N_9148);
xnor UO_471 (O_471,N_9655,N_9409);
nor UO_472 (O_472,N_9539,N_9393);
nor UO_473 (O_473,N_9530,N_9933);
and UO_474 (O_474,N_9683,N_9757);
or UO_475 (O_475,N_9031,N_9641);
or UO_476 (O_476,N_9216,N_9501);
nand UO_477 (O_477,N_9006,N_9372);
nand UO_478 (O_478,N_9540,N_9200);
xor UO_479 (O_479,N_9364,N_9060);
nand UO_480 (O_480,N_9699,N_9704);
or UO_481 (O_481,N_9253,N_9458);
xor UO_482 (O_482,N_9822,N_9265);
or UO_483 (O_483,N_9865,N_9620);
or UO_484 (O_484,N_9903,N_9722);
nand UO_485 (O_485,N_9211,N_9669);
or UO_486 (O_486,N_9326,N_9771);
and UO_487 (O_487,N_9341,N_9293);
xor UO_488 (O_488,N_9948,N_9271);
nand UO_489 (O_489,N_9985,N_9888);
xnor UO_490 (O_490,N_9889,N_9653);
nand UO_491 (O_491,N_9288,N_9040);
nand UO_492 (O_492,N_9475,N_9729);
and UO_493 (O_493,N_9193,N_9083);
nand UO_494 (O_494,N_9390,N_9789);
or UO_495 (O_495,N_9198,N_9909);
and UO_496 (O_496,N_9526,N_9298);
and UO_497 (O_497,N_9927,N_9119);
xor UO_498 (O_498,N_9808,N_9938);
nor UO_499 (O_499,N_9362,N_9012);
or UO_500 (O_500,N_9128,N_9242);
nor UO_501 (O_501,N_9790,N_9490);
or UO_502 (O_502,N_9259,N_9843);
nor UO_503 (O_503,N_9148,N_9570);
nand UO_504 (O_504,N_9212,N_9494);
and UO_505 (O_505,N_9296,N_9629);
nor UO_506 (O_506,N_9115,N_9651);
and UO_507 (O_507,N_9586,N_9855);
or UO_508 (O_508,N_9930,N_9645);
or UO_509 (O_509,N_9806,N_9072);
nor UO_510 (O_510,N_9708,N_9598);
xor UO_511 (O_511,N_9975,N_9685);
xor UO_512 (O_512,N_9055,N_9066);
and UO_513 (O_513,N_9459,N_9709);
nand UO_514 (O_514,N_9511,N_9574);
nand UO_515 (O_515,N_9002,N_9799);
and UO_516 (O_516,N_9943,N_9651);
xnor UO_517 (O_517,N_9116,N_9929);
xor UO_518 (O_518,N_9848,N_9000);
or UO_519 (O_519,N_9725,N_9395);
xor UO_520 (O_520,N_9373,N_9820);
nor UO_521 (O_521,N_9286,N_9506);
nand UO_522 (O_522,N_9406,N_9489);
and UO_523 (O_523,N_9909,N_9240);
xnor UO_524 (O_524,N_9444,N_9976);
nor UO_525 (O_525,N_9819,N_9744);
and UO_526 (O_526,N_9330,N_9782);
or UO_527 (O_527,N_9976,N_9424);
xnor UO_528 (O_528,N_9110,N_9254);
and UO_529 (O_529,N_9587,N_9231);
or UO_530 (O_530,N_9076,N_9421);
and UO_531 (O_531,N_9892,N_9921);
nor UO_532 (O_532,N_9225,N_9910);
xor UO_533 (O_533,N_9158,N_9485);
nor UO_534 (O_534,N_9866,N_9715);
and UO_535 (O_535,N_9662,N_9002);
nand UO_536 (O_536,N_9393,N_9015);
and UO_537 (O_537,N_9012,N_9385);
or UO_538 (O_538,N_9899,N_9651);
or UO_539 (O_539,N_9632,N_9653);
nor UO_540 (O_540,N_9311,N_9741);
nor UO_541 (O_541,N_9500,N_9586);
xnor UO_542 (O_542,N_9455,N_9460);
xnor UO_543 (O_543,N_9119,N_9621);
xor UO_544 (O_544,N_9774,N_9140);
nor UO_545 (O_545,N_9021,N_9573);
and UO_546 (O_546,N_9196,N_9012);
xnor UO_547 (O_547,N_9621,N_9441);
or UO_548 (O_548,N_9857,N_9609);
nand UO_549 (O_549,N_9823,N_9361);
xnor UO_550 (O_550,N_9686,N_9259);
nor UO_551 (O_551,N_9616,N_9004);
or UO_552 (O_552,N_9539,N_9268);
xnor UO_553 (O_553,N_9908,N_9944);
and UO_554 (O_554,N_9805,N_9852);
nor UO_555 (O_555,N_9940,N_9368);
nor UO_556 (O_556,N_9685,N_9055);
nand UO_557 (O_557,N_9649,N_9354);
nor UO_558 (O_558,N_9054,N_9549);
xor UO_559 (O_559,N_9040,N_9194);
or UO_560 (O_560,N_9480,N_9911);
xor UO_561 (O_561,N_9913,N_9260);
and UO_562 (O_562,N_9232,N_9834);
and UO_563 (O_563,N_9702,N_9502);
and UO_564 (O_564,N_9803,N_9901);
or UO_565 (O_565,N_9634,N_9517);
and UO_566 (O_566,N_9503,N_9196);
nand UO_567 (O_567,N_9852,N_9601);
or UO_568 (O_568,N_9539,N_9170);
xor UO_569 (O_569,N_9453,N_9399);
and UO_570 (O_570,N_9427,N_9473);
nor UO_571 (O_571,N_9372,N_9165);
nor UO_572 (O_572,N_9854,N_9474);
nor UO_573 (O_573,N_9457,N_9855);
nor UO_574 (O_574,N_9108,N_9467);
and UO_575 (O_575,N_9875,N_9141);
or UO_576 (O_576,N_9011,N_9279);
or UO_577 (O_577,N_9262,N_9140);
xnor UO_578 (O_578,N_9577,N_9440);
nand UO_579 (O_579,N_9551,N_9089);
or UO_580 (O_580,N_9205,N_9605);
nor UO_581 (O_581,N_9285,N_9021);
or UO_582 (O_582,N_9131,N_9288);
and UO_583 (O_583,N_9027,N_9622);
nand UO_584 (O_584,N_9932,N_9902);
xnor UO_585 (O_585,N_9983,N_9957);
or UO_586 (O_586,N_9847,N_9427);
and UO_587 (O_587,N_9736,N_9758);
or UO_588 (O_588,N_9872,N_9416);
xnor UO_589 (O_589,N_9215,N_9635);
and UO_590 (O_590,N_9632,N_9133);
nand UO_591 (O_591,N_9856,N_9896);
xor UO_592 (O_592,N_9297,N_9430);
or UO_593 (O_593,N_9641,N_9567);
or UO_594 (O_594,N_9919,N_9653);
and UO_595 (O_595,N_9369,N_9568);
and UO_596 (O_596,N_9705,N_9019);
xnor UO_597 (O_597,N_9225,N_9228);
xor UO_598 (O_598,N_9382,N_9304);
nor UO_599 (O_599,N_9309,N_9626);
xnor UO_600 (O_600,N_9176,N_9943);
xor UO_601 (O_601,N_9297,N_9131);
nor UO_602 (O_602,N_9970,N_9820);
xnor UO_603 (O_603,N_9342,N_9554);
nor UO_604 (O_604,N_9480,N_9561);
xnor UO_605 (O_605,N_9415,N_9663);
and UO_606 (O_606,N_9583,N_9090);
and UO_607 (O_607,N_9721,N_9094);
or UO_608 (O_608,N_9287,N_9512);
or UO_609 (O_609,N_9377,N_9312);
or UO_610 (O_610,N_9669,N_9907);
and UO_611 (O_611,N_9454,N_9459);
xnor UO_612 (O_612,N_9645,N_9423);
nand UO_613 (O_613,N_9947,N_9061);
or UO_614 (O_614,N_9471,N_9478);
and UO_615 (O_615,N_9795,N_9483);
nor UO_616 (O_616,N_9949,N_9141);
and UO_617 (O_617,N_9705,N_9873);
nor UO_618 (O_618,N_9641,N_9121);
xor UO_619 (O_619,N_9949,N_9371);
nand UO_620 (O_620,N_9675,N_9896);
or UO_621 (O_621,N_9812,N_9262);
nand UO_622 (O_622,N_9677,N_9205);
nor UO_623 (O_623,N_9611,N_9380);
and UO_624 (O_624,N_9800,N_9183);
nand UO_625 (O_625,N_9859,N_9328);
and UO_626 (O_626,N_9846,N_9013);
or UO_627 (O_627,N_9399,N_9296);
nand UO_628 (O_628,N_9900,N_9757);
nor UO_629 (O_629,N_9686,N_9875);
and UO_630 (O_630,N_9402,N_9374);
or UO_631 (O_631,N_9325,N_9375);
xor UO_632 (O_632,N_9010,N_9607);
and UO_633 (O_633,N_9948,N_9743);
nand UO_634 (O_634,N_9148,N_9342);
nand UO_635 (O_635,N_9077,N_9441);
xnor UO_636 (O_636,N_9178,N_9064);
xor UO_637 (O_637,N_9924,N_9621);
and UO_638 (O_638,N_9669,N_9381);
nor UO_639 (O_639,N_9593,N_9948);
nor UO_640 (O_640,N_9782,N_9858);
or UO_641 (O_641,N_9145,N_9739);
nand UO_642 (O_642,N_9300,N_9041);
nand UO_643 (O_643,N_9250,N_9834);
and UO_644 (O_644,N_9329,N_9325);
and UO_645 (O_645,N_9571,N_9542);
or UO_646 (O_646,N_9614,N_9991);
xor UO_647 (O_647,N_9762,N_9680);
nand UO_648 (O_648,N_9999,N_9373);
and UO_649 (O_649,N_9402,N_9005);
xor UO_650 (O_650,N_9335,N_9600);
nor UO_651 (O_651,N_9091,N_9871);
nand UO_652 (O_652,N_9312,N_9441);
nor UO_653 (O_653,N_9952,N_9975);
and UO_654 (O_654,N_9977,N_9147);
or UO_655 (O_655,N_9470,N_9389);
and UO_656 (O_656,N_9337,N_9047);
or UO_657 (O_657,N_9087,N_9420);
nand UO_658 (O_658,N_9778,N_9400);
nand UO_659 (O_659,N_9321,N_9258);
xnor UO_660 (O_660,N_9604,N_9498);
xnor UO_661 (O_661,N_9999,N_9647);
nand UO_662 (O_662,N_9867,N_9917);
nor UO_663 (O_663,N_9439,N_9780);
and UO_664 (O_664,N_9823,N_9593);
xor UO_665 (O_665,N_9930,N_9146);
nor UO_666 (O_666,N_9495,N_9205);
and UO_667 (O_667,N_9946,N_9031);
and UO_668 (O_668,N_9435,N_9699);
nor UO_669 (O_669,N_9612,N_9133);
nor UO_670 (O_670,N_9672,N_9881);
nor UO_671 (O_671,N_9206,N_9273);
and UO_672 (O_672,N_9180,N_9977);
xor UO_673 (O_673,N_9504,N_9619);
xor UO_674 (O_674,N_9631,N_9103);
nand UO_675 (O_675,N_9934,N_9117);
xnor UO_676 (O_676,N_9518,N_9700);
and UO_677 (O_677,N_9395,N_9748);
nand UO_678 (O_678,N_9485,N_9615);
and UO_679 (O_679,N_9209,N_9497);
xnor UO_680 (O_680,N_9963,N_9245);
nor UO_681 (O_681,N_9324,N_9370);
xor UO_682 (O_682,N_9412,N_9861);
nor UO_683 (O_683,N_9032,N_9562);
or UO_684 (O_684,N_9338,N_9168);
or UO_685 (O_685,N_9174,N_9013);
and UO_686 (O_686,N_9753,N_9715);
nor UO_687 (O_687,N_9880,N_9257);
xor UO_688 (O_688,N_9317,N_9407);
or UO_689 (O_689,N_9280,N_9596);
nor UO_690 (O_690,N_9954,N_9995);
nand UO_691 (O_691,N_9852,N_9517);
or UO_692 (O_692,N_9246,N_9939);
and UO_693 (O_693,N_9710,N_9988);
or UO_694 (O_694,N_9674,N_9257);
xnor UO_695 (O_695,N_9861,N_9014);
xor UO_696 (O_696,N_9635,N_9381);
nand UO_697 (O_697,N_9643,N_9607);
or UO_698 (O_698,N_9891,N_9699);
and UO_699 (O_699,N_9705,N_9579);
or UO_700 (O_700,N_9998,N_9427);
xor UO_701 (O_701,N_9174,N_9413);
and UO_702 (O_702,N_9388,N_9989);
nor UO_703 (O_703,N_9110,N_9079);
xnor UO_704 (O_704,N_9081,N_9103);
or UO_705 (O_705,N_9777,N_9441);
or UO_706 (O_706,N_9572,N_9134);
and UO_707 (O_707,N_9445,N_9773);
and UO_708 (O_708,N_9159,N_9775);
xor UO_709 (O_709,N_9745,N_9055);
nor UO_710 (O_710,N_9334,N_9615);
or UO_711 (O_711,N_9682,N_9141);
xor UO_712 (O_712,N_9329,N_9489);
and UO_713 (O_713,N_9001,N_9652);
and UO_714 (O_714,N_9301,N_9915);
and UO_715 (O_715,N_9642,N_9209);
nand UO_716 (O_716,N_9526,N_9714);
xor UO_717 (O_717,N_9314,N_9843);
or UO_718 (O_718,N_9041,N_9096);
nand UO_719 (O_719,N_9615,N_9414);
nand UO_720 (O_720,N_9364,N_9415);
xnor UO_721 (O_721,N_9689,N_9901);
xor UO_722 (O_722,N_9930,N_9736);
nand UO_723 (O_723,N_9967,N_9944);
nor UO_724 (O_724,N_9789,N_9000);
nand UO_725 (O_725,N_9458,N_9464);
nor UO_726 (O_726,N_9634,N_9042);
xnor UO_727 (O_727,N_9713,N_9408);
nor UO_728 (O_728,N_9115,N_9775);
nand UO_729 (O_729,N_9748,N_9733);
or UO_730 (O_730,N_9773,N_9218);
and UO_731 (O_731,N_9279,N_9958);
xnor UO_732 (O_732,N_9459,N_9995);
and UO_733 (O_733,N_9415,N_9072);
xor UO_734 (O_734,N_9505,N_9340);
xnor UO_735 (O_735,N_9020,N_9935);
and UO_736 (O_736,N_9290,N_9014);
nand UO_737 (O_737,N_9757,N_9885);
nor UO_738 (O_738,N_9152,N_9759);
nand UO_739 (O_739,N_9292,N_9836);
and UO_740 (O_740,N_9207,N_9047);
and UO_741 (O_741,N_9086,N_9639);
nand UO_742 (O_742,N_9632,N_9065);
or UO_743 (O_743,N_9471,N_9822);
and UO_744 (O_744,N_9469,N_9966);
and UO_745 (O_745,N_9034,N_9949);
nor UO_746 (O_746,N_9575,N_9880);
xnor UO_747 (O_747,N_9587,N_9297);
nand UO_748 (O_748,N_9074,N_9032);
or UO_749 (O_749,N_9785,N_9964);
nor UO_750 (O_750,N_9079,N_9583);
nand UO_751 (O_751,N_9638,N_9745);
or UO_752 (O_752,N_9227,N_9163);
nand UO_753 (O_753,N_9654,N_9859);
and UO_754 (O_754,N_9345,N_9335);
xnor UO_755 (O_755,N_9189,N_9505);
xor UO_756 (O_756,N_9059,N_9296);
and UO_757 (O_757,N_9532,N_9282);
and UO_758 (O_758,N_9142,N_9077);
nand UO_759 (O_759,N_9386,N_9980);
xor UO_760 (O_760,N_9327,N_9625);
xnor UO_761 (O_761,N_9627,N_9168);
nor UO_762 (O_762,N_9426,N_9627);
xor UO_763 (O_763,N_9142,N_9213);
nand UO_764 (O_764,N_9777,N_9785);
nand UO_765 (O_765,N_9384,N_9175);
xnor UO_766 (O_766,N_9671,N_9000);
nand UO_767 (O_767,N_9879,N_9351);
nand UO_768 (O_768,N_9929,N_9094);
and UO_769 (O_769,N_9276,N_9579);
nor UO_770 (O_770,N_9264,N_9823);
or UO_771 (O_771,N_9553,N_9677);
and UO_772 (O_772,N_9084,N_9351);
xnor UO_773 (O_773,N_9697,N_9547);
nand UO_774 (O_774,N_9665,N_9181);
nand UO_775 (O_775,N_9208,N_9535);
nor UO_776 (O_776,N_9588,N_9971);
nand UO_777 (O_777,N_9237,N_9562);
nand UO_778 (O_778,N_9856,N_9373);
and UO_779 (O_779,N_9430,N_9789);
or UO_780 (O_780,N_9606,N_9834);
or UO_781 (O_781,N_9225,N_9857);
xnor UO_782 (O_782,N_9894,N_9069);
xor UO_783 (O_783,N_9089,N_9753);
and UO_784 (O_784,N_9695,N_9962);
or UO_785 (O_785,N_9363,N_9465);
and UO_786 (O_786,N_9587,N_9462);
xnor UO_787 (O_787,N_9737,N_9634);
and UO_788 (O_788,N_9493,N_9049);
nor UO_789 (O_789,N_9606,N_9478);
and UO_790 (O_790,N_9996,N_9205);
or UO_791 (O_791,N_9441,N_9759);
or UO_792 (O_792,N_9389,N_9753);
and UO_793 (O_793,N_9915,N_9847);
or UO_794 (O_794,N_9396,N_9855);
xor UO_795 (O_795,N_9100,N_9612);
xnor UO_796 (O_796,N_9829,N_9936);
nand UO_797 (O_797,N_9955,N_9788);
xnor UO_798 (O_798,N_9893,N_9724);
nor UO_799 (O_799,N_9756,N_9077);
nor UO_800 (O_800,N_9084,N_9687);
nor UO_801 (O_801,N_9883,N_9815);
xnor UO_802 (O_802,N_9013,N_9842);
and UO_803 (O_803,N_9965,N_9811);
or UO_804 (O_804,N_9281,N_9805);
or UO_805 (O_805,N_9438,N_9800);
nand UO_806 (O_806,N_9116,N_9216);
nor UO_807 (O_807,N_9702,N_9291);
nor UO_808 (O_808,N_9116,N_9130);
xor UO_809 (O_809,N_9035,N_9748);
nor UO_810 (O_810,N_9335,N_9633);
nand UO_811 (O_811,N_9192,N_9154);
nand UO_812 (O_812,N_9299,N_9170);
nor UO_813 (O_813,N_9695,N_9561);
xnor UO_814 (O_814,N_9939,N_9377);
nand UO_815 (O_815,N_9788,N_9514);
or UO_816 (O_816,N_9858,N_9253);
and UO_817 (O_817,N_9106,N_9251);
nor UO_818 (O_818,N_9053,N_9261);
and UO_819 (O_819,N_9125,N_9839);
and UO_820 (O_820,N_9545,N_9814);
and UO_821 (O_821,N_9535,N_9602);
xnor UO_822 (O_822,N_9245,N_9143);
nand UO_823 (O_823,N_9460,N_9348);
nand UO_824 (O_824,N_9813,N_9960);
xnor UO_825 (O_825,N_9892,N_9907);
or UO_826 (O_826,N_9392,N_9160);
nand UO_827 (O_827,N_9188,N_9894);
nand UO_828 (O_828,N_9651,N_9751);
or UO_829 (O_829,N_9814,N_9473);
and UO_830 (O_830,N_9647,N_9739);
xor UO_831 (O_831,N_9881,N_9408);
xnor UO_832 (O_832,N_9619,N_9422);
xor UO_833 (O_833,N_9425,N_9618);
or UO_834 (O_834,N_9259,N_9064);
or UO_835 (O_835,N_9041,N_9266);
nor UO_836 (O_836,N_9640,N_9232);
xor UO_837 (O_837,N_9159,N_9855);
nor UO_838 (O_838,N_9478,N_9298);
or UO_839 (O_839,N_9615,N_9633);
xnor UO_840 (O_840,N_9982,N_9522);
and UO_841 (O_841,N_9327,N_9481);
or UO_842 (O_842,N_9423,N_9514);
or UO_843 (O_843,N_9400,N_9381);
xnor UO_844 (O_844,N_9741,N_9026);
and UO_845 (O_845,N_9698,N_9574);
and UO_846 (O_846,N_9801,N_9197);
nor UO_847 (O_847,N_9226,N_9012);
and UO_848 (O_848,N_9154,N_9062);
nand UO_849 (O_849,N_9185,N_9429);
or UO_850 (O_850,N_9815,N_9091);
nor UO_851 (O_851,N_9219,N_9593);
and UO_852 (O_852,N_9219,N_9356);
nor UO_853 (O_853,N_9033,N_9316);
xnor UO_854 (O_854,N_9161,N_9334);
nand UO_855 (O_855,N_9003,N_9632);
xnor UO_856 (O_856,N_9077,N_9770);
nand UO_857 (O_857,N_9171,N_9421);
and UO_858 (O_858,N_9357,N_9441);
or UO_859 (O_859,N_9202,N_9004);
and UO_860 (O_860,N_9909,N_9607);
nor UO_861 (O_861,N_9170,N_9629);
and UO_862 (O_862,N_9954,N_9326);
and UO_863 (O_863,N_9586,N_9565);
or UO_864 (O_864,N_9059,N_9860);
nand UO_865 (O_865,N_9882,N_9184);
nor UO_866 (O_866,N_9337,N_9815);
xnor UO_867 (O_867,N_9132,N_9164);
nand UO_868 (O_868,N_9134,N_9251);
nor UO_869 (O_869,N_9622,N_9858);
xor UO_870 (O_870,N_9268,N_9021);
nand UO_871 (O_871,N_9491,N_9249);
nand UO_872 (O_872,N_9805,N_9835);
nor UO_873 (O_873,N_9587,N_9388);
or UO_874 (O_874,N_9559,N_9866);
or UO_875 (O_875,N_9184,N_9669);
and UO_876 (O_876,N_9538,N_9589);
and UO_877 (O_877,N_9233,N_9936);
xnor UO_878 (O_878,N_9953,N_9207);
xnor UO_879 (O_879,N_9346,N_9314);
or UO_880 (O_880,N_9813,N_9615);
nor UO_881 (O_881,N_9950,N_9603);
nand UO_882 (O_882,N_9190,N_9621);
nand UO_883 (O_883,N_9872,N_9938);
xnor UO_884 (O_884,N_9122,N_9876);
and UO_885 (O_885,N_9488,N_9212);
nor UO_886 (O_886,N_9099,N_9801);
or UO_887 (O_887,N_9616,N_9647);
and UO_888 (O_888,N_9582,N_9682);
and UO_889 (O_889,N_9446,N_9105);
or UO_890 (O_890,N_9068,N_9798);
or UO_891 (O_891,N_9914,N_9353);
and UO_892 (O_892,N_9544,N_9296);
nand UO_893 (O_893,N_9542,N_9349);
nand UO_894 (O_894,N_9970,N_9449);
xnor UO_895 (O_895,N_9345,N_9987);
nand UO_896 (O_896,N_9185,N_9378);
or UO_897 (O_897,N_9249,N_9998);
xnor UO_898 (O_898,N_9920,N_9796);
nor UO_899 (O_899,N_9627,N_9643);
or UO_900 (O_900,N_9931,N_9997);
or UO_901 (O_901,N_9623,N_9085);
xnor UO_902 (O_902,N_9624,N_9971);
nand UO_903 (O_903,N_9845,N_9006);
xor UO_904 (O_904,N_9163,N_9010);
or UO_905 (O_905,N_9809,N_9742);
xor UO_906 (O_906,N_9545,N_9393);
or UO_907 (O_907,N_9297,N_9088);
nand UO_908 (O_908,N_9246,N_9118);
nand UO_909 (O_909,N_9416,N_9485);
nor UO_910 (O_910,N_9616,N_9717);
nand UO_911 (O_911,N_9242,N_9586);
and UO_912 (O_912,N_9701,N_9411);
nand UO_913 (O_913,N_9650,N_9294);
xnor UO_914 (O_914,N_9351,N_9805);
and UO_915 (O_915,N_9812,N_9169);
nor UO_916 (O_916,N_9701,N_9122);
nand UO_917 (O_917,N_9989,N_9795);
or UO_918 (O_918,N_9830,N_9737);
nor UO_919 (O_919,N_9163,N_9640);
nor UO_920 (O_920,N_9418,N_9037);
and UO_921 (O_921,N_9811,N_9890);
or UO_922 (O_922,N_9989,N_9336);
and UO_923 (O_923,N_9134,N_9086);
and UO_924 (O_924,N_9848,N_9167);
and UO_925 (O_925,N_9670,N_9894);
nor UO_926 (O_926,N_9736,N_9409);
or UO_927 (O_927,N_9069,N_9184);
nand UO_928 (O_928,N_9070,N_9045);
xnor UO_929 (O_929,N_9658,N_9286);
nand UO_930 (O_930,N_9241,N_9766);
and UO_931 (O_931,N_9235,N_9298);
nand UO_932 (O_932,N_9150,N_9471);
xor UO_933 (O_933,N_9784,N_9047);
nand UO_934 (O_934,N_9360,N_9927);
xnor UO_935 (O_935,N_9012,N_9045);
xnor UO_936 (O_936,N_9731,N_9358);
nand UO_937 (O_937,N_9717,N_9213);
nand UO_938 (O_938,N_9017,N_9899);
xor UO_939 (O_939,N_9221,N_9030);
xor UO_940 (O_940,N_9231,N_9877);
or UO_941 (O_941,N_9752,N_9779);
nand UO_942 (O_942,N_9705,N_9897);
xor UO_943 (O_943,N_9921,N_9188);
nand UO_944 (O_944,N_9607,N_9633);
or UO_945 (O_945,N_9077,N_9594);
and UO_946 (O_946,N_9350,N_9115);
nand UO_947 (O_947,N_9133,N_9332);
nor UO_948 (O_948,N_9282,N_9388);
nand UO_949 (O_949,N_9589,N_9469);
or UO_950 (O_950,N_9974,N_9333);
nor UO_951 (O_951,N_9396,N_9898);
or UO_952 (O_952,N_9157,N_9286);
nand UO_953 (O_953,N_9926,N_9691);
or UO_954 (O_954,N_9577,N_9683);
nor UO_955 (O_955,N_9920,N_9969);
or UO_956 (O_956,N_9208,N_9087);
nor UO_957 (O_957,N_9591,N_9624);
nand UO_958 (O_958,N_9780,N_9206);
xnor UO_959 (O_959,N_9632,N_9686);
or UO_960 (O_960,N_9665,N_9795);
or UO_961 (O_961,N_9706,N_9415);
nor UO_962 (O_962,N_9303,N_9147);
and UO_963 (O_963,N_9676,N_9126);
xnor UO_964 (O_964,N_9788,N_9382);
and UO_965 (O_965,N_9664,N_9820);
nand UO_966 (O_966,N_9212,N_9717);
nor UO_967 (O_967,N_9468,N_9180);
nor UO_968 (O_968,N_9991,N_9743);
xnor UO_969 (O_969,N_9019,N_9443);
xor UO_970 (O_970,N_9477,N_9472);
or UO_971 (O_971,N_9396,N_9514);
nor UO_972 (O_972,N_9079,N_9872);
and UO_973 (O_973,N_9887,N_9265);
xnor UO_974 (O_974,N_9771,N_9756);
nor UO_975 (O_975,N_9215,N_9079);
and UO_976 (O_976,N_9456,N_9627);
or UO_977 (O_977,N_9036,N_9662);
nor UO_978 (O_978,N_9559,N_9050);
or UO_979 (O_979,N_9584,N_9344);
and UO_980 (O_980,N_9395,N_9673);
or UO_981 (O_981,N_9332,N_9983);
nand UO_982 (O_982,N_9538,N_9645);
xnor UO_983 (O_983,N_9832,N_9769);
xnor UO_984 (O_984,N_9198,N_9539);
nand UO_985 (O_985,N_9077,N_9378);
and UO_986 (O_986,N_9980,N_9918);
nand UO_987 (O_987,N_9197,N_9850);
nand UO_988 (O_988,N_9023,N_9998);
nor UO_989 (O_989,N_9022,N_9375);
nand UO_990 (O_990,N_9124,N_9146);
nor UO_991 (O_991,N_9371,N_9334);
and UO_992 (O_992,N_9971,N_9741);
nor UO_993 (O_993,N_9886,N_9810);
nor UO_994 (O_994,N_9234,N_9963);
and UO_995 (O_995,N_9863,N_9458);
nor UO_996 (O_996,N_9699,N_9316);
and UO_997 (O_997,N_9366,N_9208);
and UO_998 (O_998,N_9898,N_9538);
nand UO_999 (O_999,N_9201,N_9886);
xnor UO_1000 (O_1000,N_9265,N_9722);
and UO_1001 (O_1001,N_9976,N_9785);
nor UO_1002 (O_1002,N_9048,N_9170);
or UO_1003 (O_1003,N_9433,N_9278);
xnor UO_1004 (O_1004,N_9405,N_9476);
nor UO_1005 (O_1005,N_9063,N_9487);
or UO_1006 (O_1006,N_9958,N_9150);
xnor UO_1007 (O_1007,N_9502,N_9122);
or UO_1008 (O_1008,N_9436,N_9979);
xor UO_1009 (O_1009,N_9238,N_9592);
nand UO_1010 (O_1010,N_9271,N_9918);
nand UO_1011 (O_1011,N_9903,N_9530);
or UO_1012 (O_1012,N_9896,N_9237);
and UO_1013 (O_1013,N_9187,N_9123);
nand UO_1014 (O_1014,N_9566,N_9582);
xnor UO_1015 (O_1015,N_9478,N_9915);
or UO_1016 (O_1016,N_9568,N_9513);
nand UO_1017 (O_1017,N_9692,N_9299);
nand UO_1018 (O_1018,N_9910,N_9378);
nor UO_1019 (O_1019,N_9478,N_9900);
nand UO_1020 (O_1020,N_9538,N_9484);
nand UO_1021 (O_1021,N_9824,N_9270);
or UO_1022 (O_1022,N_9675,N_9687);
nand UO_1023 (O_1023,N_9930,N_9775);
nor UO_1024 (O_1024,N_9956,N_9660);
xor UO_1025 (O_1025,N_9661,N_9064);
xor UO_1026 (O_1026,N_9982,N_9858);
nor UO_1027 (O_1027,N_9961,N_9706);
or UO_1028 (O_1028,N_9286,N_9617);
and UO_1029 (O_1029,N_9374,N_9590);
nand UO_1030 (O_1030,N_9164,N_9661);
or UO_1031 (O_1031,N_9144,N_9660);
or UO_1032 (O_1032,N_9512,N_9822);
nand UO_1033 (O_1033,N_9890,N_9134);
xor UO_1034 (O_1034,N_9261,N_9256);
and UO_1035 (O_1035,N_9692,N_9839);
nand UO_1036 (O_1036,N_9003,N_9005);
nor UO_1037 (O_1037,N_9372,N_9033);
and UO_1038 (O_1038,N_9329,N_9739);
nor UO_1039 (O_1039,N_9667,N_9162);
or UO_1040 (O_1040,N_9086,N_9091);
and UO_1041 (O_1041,N_9907,N_9465);
or UO_1042 (O_1042,N_9305,N_9880);
and UO_1043 (O_1043,N_9160,N_9163);
nor UO_1044 (O_1044,N_9635,N_9439);
and UO_1045 (O_1045,N_9893,N_9763);
xor UO_1046 (O_1046,N_9000,N_9276);
xnor UO_1047 (O_1047,N_9704,N_9505);
and UO_1048 (O_1048,N_9853,N_9175);
xor UO_1049 (O_1049,N_9217,N_9916);
nand UO_1050 (O_1050,N_9400,N_9913);
and UO_1051 (O_1051,N_9654,N_9431);
and UO_1052 (O_1052,N_9879,N_9236);
nor UO_1053 (O_1053,N_9832,N_9961);
xnor UO_1054 (O_1054,N_9786,N_9952);
xor UO_1055 (O_1055,N_9055,N_9417);
nand UO_1056 (O_1056,N_9260,N_9024);
xor UO_1057 (O_1057,N_9565,N_9978);
and UO_1058 (O_1058,N_9991,N_9312);
or UO_1059 (O_1059,N_9453,N_9802);
or UO_1060 (O_1060,N_9493,N_9636);
and UO_1061 (O_1061,N_9150,N_9446);
nor UO_1062 (O_1062,N_9295,N_9442);
nor UO_1063 (O_1063,N_9773,N_9785);
or UO_1064 (O_1064,N_9981,N_9155);
nand UO_1065 (O_1065,N_9200,N_9018);
nor UO_1066 (O_1066,N_9294,N_9392);
nand UO_1067 (O_1067,N_9886,N_9663);
xnor UO_1068 (O_1068,N_9378,N_9847);
nand UO_1069 (O_1069,N_9882,N_9706);
nand UO_1070 (O_1070,N_9580,N_9358);
nor UO_1071 (O_1071,N_9774,N_9197);
xnor UO_1072 (O_1072,N_9189,N_9889);
or UO_1073 (O_1073,N_9609,N_9978);
nand UO_1074 (O_1074,N_9233,N_9331);
xor UO_1075 (O_1075,N_9648,N_9291);
and UO_1076 (O_1076,N_9029,N_9174);
and UO_1077 (O_1077,N_9904,N_9582);
or UO_1078 (O_1078,N_9490,N_9140);
nand UO_1079 (O_1079,N_9491,N_9877);
xnor UO_1080 (O_1080,N_9627,N_9922);
and UO_1081 (O_1081,N_9211,N_9652);
and UO_1082 (O_1082,N_9919,N_9788);
or UO_1083 (O_1083,N_9949,N_9522);
and UO_1084 (O_1084,N_9440,N_9303);
or UO_1085 (O_1085,N_9269,N_9873);
xor UO_1086 (O_1086,N_9275,N_9518);
xor UO_1087 (O_1087,N_9733,N_9413);
xor UO_1088 (O_1088,N_9826,N_9551);
nand UO_1089 (O_1089,N_9795,N_9216);
or UO_1090 (O_1090,N_9190,N_9470);
and UO_1091 (O_1091,N_9562,N_9119);
xnor UO_1092 (O_1092,N_9168,N_9987);
or UO_1093 (O_1093,N_9578,N_9069);
xnor UO_1094 (O_1094,N_9389,N_9551);
and UO_1095 (O_1095,N_9536,N_9538);
or UO_1096 (O_1096,N_9611,N_9467);
xnor UO_1097 (O_1097,N_9813,N_9421);
nand UO_1098 (O_1098,N_9966,N_9097);
xor UO_1099 (O_1099,N_9133,N_9027);
nand UO_1100 (O_1100,N_9950,N_9376);
and UO_1101 (O_1101,N_9496,N_9981);
xor UO_1102 (O_1102,N_9804,N_9958);
and UO_1103 (O_1103,N_9815,N_9813);
nand UO_1104 (O_1104,N_9875,N_9504);
nand UO_1105 (O_1105,N_9501,N_9277);
xnor UO_1106 (O_1106,N_9961,N_9068);
xnor UO_1107 (O_1107,N_9676,N_9536);
and UO_1108 (O_1108,N_9715,N_9421);
nand UO_1109 (O_1109,N_9068,N_9174);
nor UO_1110 (O_1110,N_9214,N_9982);
nand UO_1111 (O_1111,N_9217,N_9586);
or UO_1112 (O_1112,N_9359,N_9001);
xor UO_1113 (O_1113,N_9944,N_9225);
and UO_1114 (O_1114,N_9902,N_9959);
and UO_1115 (O_1115,N_9081,N_9609);
xor UO_1116 (O_1116,N_9313,N_9867);
nand UO_1117 (O_1117,N_9670,N_9592);
nor UO_1118 (O_1118,N_9434,N_9151);
or UO_1119 (O_1119,N_9553,N_9951);
xor UO_1120 (O_1120,N_9245,N_9128);
and UO_1121 (O_1121,N_9051,N_9886);
nand UO_1122 (O_1122,N_9282,N_9965);
nor UO_1123 (O_1123,N_9645,N_9765);
or UO_1124 (O_1124,N_9365,N_9943);
or UO_1125 (O_1125,N_9984,N_9516);
nor UO_1126 (O_1126,N_9275,N_9263);
nand UO_1127 (O_1127,N_9659,N_9707);
xnor UO_1128 (O_1128,N_9724,N_9451);
nand UO_1129 (O_1129,N_9069,N_9116);
xor UO_1130 (O_1130,N_9736,N_9318);
nor UO_1131 (O_1131,N_9840,N_9977);
and UO_1132 (O_1132,N_9286,N_9054);
or UO_1133 (O_1133,N_9251,N_9521);
nor UO_1134 (O_1134,N_9550,N_9270);
nand UO_1135 (O_1135,N_9763,N_9858);
and UO_1136 (O_1136,N_9070,N_9309);
xnor UO_1137 (O_1137,N_9297,N_9813);
nor UO_1138 (O_1138,N_9082,N_9937);
nand UO_1139 (O_1139,N_9255,N_9742);
xor UO_1140 (O_1140,N_9996,N_9188);
nand UO_1141 (O_1141,N_9750,N_9011);
and UO_1142 (O_1142,N_9533,N_9438);
xnor UO_1143 (O_1143,N_9418,N_9821);
xnor UO_1144 (O_1144,N_9947,N_9897);
and UO_1145 (O_1145,N_9332,N_9100);
or UO_1146 (O_1146,N_9461,N_9006);
or UO_1147 (O_1147,N_9415,N_9524);
xnor UO_1148 (O_1148,N_9819,N_9676);
nand UO_1149 (O_1149,N_9927,N_9063);
nand UO_1150 (O_1150,N_9163,N_9413);
or UO_1151 (O_1151,N_9586,N_9342);
nand UO_1152 (O_1152,N_9211,N_9003);
and UO_1153 (O_1153,N_9655,N_9707);
and UO_1154 (O_1154,N_9036,N_9706);
nand UO_1155 (O_1155,N_9501,N_9464);
nor UO_1156 (O_1156,N_9801,N_9327);
xor UO_1157 (O_1157,N_9017,N_9548);
nor UO_1158 (O_1158,N_9644,N_9112);
and UO_1159 (O_1159,N_9698,N_9696);
and UO_1160 (O_1160,N_9585,N_9141);
nor UO_1161 (O_1161,N_9384,N_9262);
nand UO_1162 (O_1162,N_9188,N_9258);
nand UO_1163 (O_1163,N_9199,N_9763);
or UO_1164 (O_1164,N_9402,N_9375);
xnor UO_1165 (O_1165,N_9956,N_9584);
and UO_1166 (O_1166,N_9430,N_9027);
nor UO_1167 (O_1167,N_9177,N_9698);
and UO_1168 (O_1168,N_9528,N_9127);
xor UO_1169 (O_1169,N_9683,N_9825);
nand UO_1170 (O_1170,N_9495,N_9285);
or UO_1171 (O_1171,N_9522,N_9256);
nand UO_1172 (O_1172,N_9580,N_9484);
xnor UO_1173 (O_1173,N_9684,N_9004);
and UO_1174 (O_1174,N_9461,N_9493);
xor UO_1175 (O_1175,N_9744,N_9537);
nor UO_1176 (O_1176,N_9032,N_9295);
xor UO_1177 (O_1177,N_9983,N_9185);
nor UO_1178 (O_1178,N_9420,N_9418);
xnor UO_1179 (O_1179,N_9852,N_9651);
and UO_1180 (O_1180,N_9794,N_9497);
nand UO_1181 (O_1181,N_9737,N_9516);
nand UO_1182 (O_1182,N_9489,N_9164);
and UO_1183 (O_1183,N_9621,N_9858);
nor UO_1184 (O_1184,N_9191,N_9899);
nand UO_1185 (O_1185,N_9485,N_9989);
xnor UO_1186 (O_1186,N_9935,N_9848);
xnor UO_1187 (O_1187,N_9736,N_9889);
nand UO_1188 (O_1188,N_9433,N_9036);
xor UO_1189 (O_1189,N_9501,N_9470);
xor UO_1190 (O_1190,N_9522,N_9666);
xor UO_1191 (O_1191,N_9149,N_9336);
or UO_1192 (O_1192,N_9686,N_9985);
and UO_1193 (O_1193,N_9364,N_9629);
xor UO_1194 (O_1194,N_9285,N_9979);
or UO_1195 (O_1195,N_9981,N_9904);
nor UO_1196 (O_1196,N_9606,N_9566);
or UO_1197 (O_1197,N_9002,N_9489);
xor UO_1198 (O_1198,N_9307,N_9616);
or UO_1199 (O_1199,N_9016,N_9868);
xor UO_1200 (O_1200,N_9718,N_9364);
and UO_1201 (O_1201,N_9567,N_9216);
and UO_1202 (O_1202,N_9694,N_9477);
nand UO_1203 (O_1203,N_9310,N_9189);
nor UO_1204 (O_1204,N_9024,N_9216);
and UO_1205 (O_1205,N_9982,N_9453);
or UO_1206 (O_1206,N_9691,N_9851);
and UO_1207 (O_1207,N_9244,N_9814);
nor UO_1208 (O_1208,N_9511,N_9194);
nand UO_1209 (O_1209,N_9467,N_9981);
nand UO_1210 (O_1210,N_9190,N_9980);
nor UO_1211 (O_1211,N_9392,N_9374);
xor UO_1212 (O_1212,N_9741,N_9897);
and UO_1213 (O_1213,N_9576,N_9525);
nand UO_1214 (O_1214,N_9607,N_9906);
nor UO_1215 (O_1215,N_9381,N_9618);
xnor UO_1216 (O_1216,N_9559,N_9307);
or UO_1217 (O_1217,N_9468,N_9991);
or UO_1218 (O_1218,N_9468,N_9346);
nand UO_1219 (O_1219,N_9811,N_9480);
or UO_1220 (O_1220,N_9653,N_9276);
or UO_1221 (O_1221,N_9851,N_9083);
or UO_1222 (O_1222,N_9478,N_9777);
nand UO_1223 (O_1223,N_9731,N_9577);
xor UO_1224 (O_1224,N_9635,N_9940);
nor UO_1225 (O_1225,N_9473,N_9581);
nor UO_1226 (O_1226,N_9945,N_9553);
nor UO_1227 (O_1227,N_9079,N_9695);
nand UO_1228 (O_1228,N_9054,N_9613);
nor UO_1229 (O_1229,N_9335,N_9211);
xnor UO_1230 (O_1230,N_9184,N_9526);
and UO_1231 (O_1231,N_9164,N_9485);
nand UO_1232 (O_1232,N_9109,N_9402);
nand UO_1233 (O_1233,N_9959,N_9326);
nand UO_1234 (O_1234,N_9231,N_9717);
nand UO_1235 (O_1235,N_9480,N_9629);
xnor UO_1236 (O_1236,N_9359,N_9818);
and UO_1237 (O_1237,N_9451,N_9138);
or UO_1238 (O_1238,N_9975,N_9307);
xnor UO_1239 (O_1239,N_9616,N_9350);
and UO_1240 (O_1240,N_9367,N_9813);
xnor UO_1241 (O_1241,N_9905,N_9595);
xor UO_1242 (O_1242,N_9248,N_9482);
or UO_1243 (O_1243,N_9937,N_9929);
xnor UO_1244 (O_1244,N_9071,N_9114);
nor UO_1245 (O_1245,N_9933,N_9636);
nor UO_1246 (O_1246,N_9225,N_9930);
nor UO_1247 (O_1247,N_9607,N_9776);
nor UO_1248 (O_1248,N_9341,N_9001);
nand UO_1249 (O_1249,N_9672,N_9670);
or UO_1250 (O_1250,N_9194,N_9877);
nor UO_1251 (O_1251,N_9962,N_9713);
nand UO_1252 (O_1252,N_9355,N_9595);
and UO_1253 (O_1253,N_9709,N_9622);
or UO_1254 (O_1254,N_9868,N_9231);
nor UO_1255 (O_1255,N_9814,N_9140);
and UO_1256 (O_1256,N_9828,N_9278);
or UO_1257 (O_1257,N_9656,N_9221);
xnor UO_1258 (O_1258,N_9766,N_9020);
nor UO_1259 (O_1259,N_9385,N_9124);
nand UO_1260 (O_1260,N_9486,N_9457);
and UO_1261 (O_1261,N_9153,N_9087);
or UO_1262 (O_1262,N_9107,N_9262);
or UO_1263 (O_1263,N_9467,N_9831);
nand UO_1264 (O_1264,N_9703,N_9630);
nand UO_1265 (O_1265,N_9217,N_9494);
and UO_1266 (O_1266,N_9759,N_9603);
nor UO_1267 (O_1267,N_9989,N_9300);
nor UO_1268 (O_1268,N_9114,N_9369);
and UO_1269 (O_1269,N_9542,N_9899);
nor UO_1270 (O_1270,N_9629,N_9118);
xnor UO_1271 (O_1271,N_9565,N_9910);
nand UO_1272 (O_1272,N_9846,N_9112);
xnor UO_1273 (O_1273,N_9203,N_9731);
xor UO_1274 (O_1274,N_9610,N_9315);
or UO_1275 (O_1275,N_9305,N_9599);
or UO_1276 (O_1276,N_9355,N_9656);
or UO_1277 (O_1277,N_9422,N_9874);
nor UO_1278 (O_1278,N_9815,N_9164);
xor UO_1279 (O_1279,N_9467,N_9442);
or UO_1280 (O_1280,N_9713,N_9119);
and UO_1281 (O_1281,N_9325,N_9608);
nand UO_1282 (O_1282,N_9808,N_9471);
or UO_1283 (O_1283,N_9971,N_9738);
or UO_1284 (O_1284,N_9429,N_9796);
nor UO_1285 (O_1285,N_9991,N_9160);
nand UO_1286 (O_1286,N_9082,N_9062);
and UO_1287 (O_1287,N_9147,N_9842);
or UO_1288 (O_1288,N_9248,N_9903);
and UO_1289 (O_1289,N_9633,N_9346);
or UO_1290 (O_1290,N_9326,N_9459);
nand UO_1291 (O_1291,N_9940,N_9257);
nand UO_1292 (O_1292,N_9991,N_9106);
nor UO_1293 (O_1293,N_9430,N_9784);
or UO_1294 (O_1294,N_9547,N_9824);
xor UO_1295 (O_1295,N_9362,N_9712);
and UO_1296 (O_1296,N_9731,N_9141);
and UO_1297 (O_1297,N_9634,N_9232);
or UO_1298 (O_1298,N_9041,N_9012);
nor UO_1299 (O_1299,N_9403,N_9232);
xor UO_1300 (O_1300,N_9423,N_9672);
or UO_1301 (O_1301,N_9136,N_9391);
or UO_1302 (O_1302,N_9350,N_9307);
and UO_1303 (O_1303,N_9829,N_9985);
and UO_1304 (O_1304,N_9037,N_9937);
xnor UO_1305 (O_1305,N_9638,N_9066);
nand UO_1306 (O_1306,N_9782,N_9395);
nor UO_1307 (O_1307,N_9659,N_9200);
nor UO_1308 (O_1308,N_9783,N_9693);
nand UO_1309 (O_1309,N_9720,N_9926);
nor UO_1310 (O_1310,N_9757,N_9756);
nand UO_1311 (O_1311,N_9923,N_9143);
and UO_1312 (O_1312,N_9395,N_9847);
nor UO_1313 (O_1313,N_9366,N_9790);
or UO_1314 (O_1314,N_9782,N_9786);
or UO_1315 (O_1315,N_9185,N_9895);
and UO_1316 (O_1316,N_9054,N_9764);
or UO_1317 (O_1317,N_9278,N_9773);
and UO_1318 (O_1318,N_9943,N_9765);
or UO_1319 (O_1319,N_9168,N_9220);
nand UO_1320 (O_1320,N_9844,N_9989);
and UO_1321 (O_1321,N_9730,N_9237);
nand UO_1322 (O_1322,N_9105,N_9172);
xnor UO_1323 (O_1323,N_9985,N_9982);
nor UO_1324 (O_1324,N_9534,N_9231);
or UO_1325 (O_1325,N_9794,N_9618);
and UO_1326 (O_1326,N_9522,N_9627);
or UO_1327 (O_1327,N_9599,N_9901);
nor UO_1328 (O_1328,N_9940,N_9611);
or UO_1329 (O_1329,N_9659,N_9106);
nor UO_1330 (O_1330,N_9935,N_9831);
xnor UO_1331 (O_1331,N_9269,N_9938);
nor UO_1332 (O_1332,N_9408,N_9590);
nor UO_1333 (O_1333,N_9259,N_9520);
nor UO_1334 (O_1334,N_9669,N_9609);
nor UO_1335 (O_1335,N_9912,N_9877);
or UO_1336 (O_1336,N_9985,N_9403);
xnor UO_1337 (O_1337,N_9867,N_9284);
nor UO_1338 (O_1338,N_9388,N_9267);
nand UO_1339 (O_1339,N_9318,N_9677);
or UO_1340 (O_1340,N_9137,N_9918);
nor UO_1341 (O_1341,N_9113,N_9585);
nor UO_1342 (O_1342,N_9383,N_9300);
nand UO_1343 (O_1343,N_9774,N_9534);
nor UO_1344 (O_1344,N_9792,N_9295);
and UO_1345 (O_1345,N_9593,N_9918);
xor UO_1346 (O_1346,N_9282,N_9981);
nor UO_1347 (O_1347,N_9879,N_9634);
nand UO_1348 (O_1348,N_9125,N_9626);
xor UO_1349 (O_1349,N_9954,N_9817);
nor UO_1350 (O_1350,N_9958,N_9570);
nand UO_1351 (O_1351,N_9386,N_9053);
xnor UO_1352 (O_1352,N_9377,N_9398);
and UO_1353 (O_1353,N_9824,N_9062);
nand UO_1354 (O_1354,N_9803,N_9903);
and UO_1355 (O_1355,N_9414,N_9104);
nor UO_1356 (O_1356,N_9440,N_9196);
nor UO_1357 (O_1357,N_9339,N_9032);
nor UO_1358 (O_1358,N_9771,N_9841);
and UO_1359 (O_1359,N_9117,N_9743);
and UO_1360 (O_1360,N_9191,N_9722);
and UO_1361 (O_1361,N_9376,N_9337);
and UO_1362 (O_1362,N_9380,N_9047);
nand UO_1363 (O_1363,N_9504,N_9676);
nand UO_1364 (O_1364,N_9579,N_9092);
nor UO_1365 (O_1365,N_9532,N_9500);
or UO_1366 (O_1366,N_9101,N_9511);
nand UO_1367 (O_1367,N_9019,N_9664);
xnor UO_1368 (O_1368,N_9742,N_9432);
or UO_1369 (O_1369,N_9941,N_9840);
xor UO_1370 (O_1370,N_9144,N_9859);
xnor UO_1371 (O_1371,N_9910,N_9728);
and UO_1372 (O_1372,N_9843,N_9404);
nor UO_1373 (O_1373,N_9129,N_9259);
or UO_1374 (O_1374,N_9656,N_9157);
nor UO_1375 (O_1375,N_9232,N_9296);
xnor UO_1376 (O_1376,N_9912,N_9747);
nand UO_1377 (O_1377,N_9516,N_9819);
nand UO_1378 (O_1378,N_9298,N_9418);
xnor UO_1379 (O_1379,N_9810,N_9489);
xor UO_1380 (O_1380,N_9828,N_9747);
and UO_1381 (O_1381,N_9037,N_9387);
or UO_1382 (O_1382,N_9962,N_9992);
nor UO_1383 (O_1383,N_9260,N_9729);
and UO_1384 (O_1384,N_9548,N_9092);
or UO_1385 (O_1385,N_9485,N_9165);
xnor UO_1386 (O_1386,N_9206,N_9776);
and UO_1387 (O_1387,N_9189,N_9412);
or UO_1388 (O_1388,N_9374,N_9793);
and UO_1389 (O_1389,N_9250,N_9930);
or UO_1390 (O_1390,N_9098,N_9618);
xnor UO_1391 (O_1391,N_9843,N_9167);
or UO_1392 (O_1392,N_9538,N_9522);
nand UO_1393 (O_1393,N_9994,N_9430);
xor UO_1394 (O_1394,N_9486,N_9570);
nand UO_1395 (O_1395,N_9294,N_9164);
nor UO_1396 (O_1396,N_9076,N_9584);
nor UO_1397 (O_1397,N_9304,N_9073);
nand UO_1398 (O_1398,N_9388,N_9071);
nand UO_1399 (O_1399,N_9957,N_9246);
nand UO_1400 (O_1400,N_9357,N_9377);
nand UO_1401 (O_1401,N_9966,N_9927);
nor UO_1402 (O_1402,N_9237,N_9278);
or UO_1403 (O_1403,N_9438,N_9479);
nand UO_1404 (O_1404,N_9742,N_9675);
xnor UO_1405 (O_1405,N_9526,N_9888);
xor UO_1406 (O_1406,N_9342,N_9061);
nand UO_1407 (O_1407,N_9967,N_9036);
xor UO_1408 (O_1408,N_9122,N_9065);
nand UO_1409 (O_1409,N_9461,N_9944);
xnor UO_1410 (O_1410,N_9269,N_9048);
xnor UO_1411 (O_1411,N_9339,N_9811);
nand UO_1412 (O_1412,N_9598,N_9525);
nor UO_1413 (O_1413,N_9785,N_9749);
and UO_1414 (O_1414,N_9267,N_9010);
or UO_1415 (O_1415,N_9201,N_9176);
xor UO_1416 (O_1416,N_9284,N_9067);
or UO_1417 (O_1417,N_9640,N_9830);
nor UO_1418 (O_1418,N_9967,N_9385);
or UO_1419 (O_1419,N_9451,N_9962);
xor UO_1420 (O_1420,N_9494,N_9716);
nor UO_1421 (O_1421,N_9139,N_9872);
nand UO_1422 (O_1422,N_9807,N_9675);
and UO_1423 (O_1423,N_9589,N_9953);
nand UO_1424 (O_1424,N_9307,N_9965);
and UO_1425 (O_1425,N_9123,N_9704);
nand UO_1426 (O_1426,N_9265,N_9160);
and UO_1427 (O_1427,N_9331,N_9284);
nand UO_1428 (O_1428,N_9673,N_9442);
and UO_1429 (O_1429,N_9185,N_9375);
nor UO_1430 (O_1430,N_9096,N_9015);
nand UO_1431 (O_1431,N_9858,N_9749);
xor UO_1432 (O_1432,N_9293,N_9642);
xnor UO_1433 (O_1433,N_9852,N_9274);
and UO_1434 (O_1434,N_9432,N_9405);
nor UO_1435 (O_1435,N_9728,N_9306);
or UO_1436 (O_1436,N_9619,N_9705);
and UO_1437 (O_1437,N_9902,N_9977);
and UO_1438 (O_1438,N_9141,N_9584);
xor UO_1439 (O_1439,N_9317,N_9120);
and UO_1440 (O_1440,N_9579,N_9694);
nor UO_1441 (O_1441,N_9390,N_9021);
nand UO_1442 (O_1442,N_9057,N_9620);
and UO_1443 (O_1443,N_9159,N_9772);
or UO_1444 (O_1444,N_9331,N_9681);
nor UO_1445 (O_1445,N_9371,N_9626);
xnor UO_1446 (O_1446,N_9898,N_9610);
nand UO_1447 (O_1447,N_9547,N_9882);
nand UO_1448 (O_1448,N_9201,N_9913);
and UO_1449 (O_1449,N_9221,N_9769);
or UO_1450 (O_1450,N_9639,N_9018);
and UO_1451 (O_1451,N_9728,N_9267);
or UO_1452 (O_1452,N_9268,N_9617);
and UO_1453 (O_1453,N_9264,N_9828);
xnor UO_1454 (O_1454,N_9247,N_9716);
nor UO_1455 (O_1455,N_9082,N_9795);
nand UO_1456 (O_1456,N_9224,N_9838);
nor UO_1457 (O_1457,N_9598,N_9000);
xnor UO_1458 (O_1458,N_9313,N_9224);
nand UO_1459 (O_1459,N_9600,N_9900);
xnor UO_1460 (O_1460,N_9432,N_9581);
and UO_1461 (O_1461,N_9201,N_9304);
xnor UO_1462 (O_1462,N_9489,N_9412);
and UO_1463 (O_1463,N_9760,N_9542);
xnor UO_1464 (O_1464,N_9797,N_9851);
or UO_1465 (O_1465,N_9346,N_9846);
nor UO_1466 (O_1466,N_9971,N_9706);
nand UO_1467 (O_1467,N_9701,N_9900);
nand UO_1468 (O_1468,N_9641,N_9297);
nor UO_1469 (O_1469,N_9510,N_9151);
and UO_1470 (O_1470,N_9436,N_9319);
or UO_1471 (O_1471,N_9627,N_9714);
nand UO_1472 (O_1472,N_9714,N_9291);
nor UO_1473 (O_1473,N_9391,N_9192);
and UO_1474 (O_1474,N_9508,N_9124);
xnor UO_1475 (O_1475,N_9584,N_9750);
nor UO_1476 (O_1476,N_9787,N_9368);
nand UO_1477 (O_1477,N_9795,N_9764);
nand UO_1478 (O_1478,N_9454,N_9353);
nor UO_1479 (O_1479,N_9223,N_9356);
xor UO_1480 (O_1480,N_9068,N_9574);
nor UO_1481 (O_1481,N_9483,N_9997);
nor UO_1482 (O_1482,N_9078,N_9367);
nand UO_1483 (O_1483,N_9221,N_9677);
nor UO_1484 (O_1484,N_9945,N_9972);
nand UO_1485 (O_1485,N_9359,N_9867);
nand UO_1486 (O_1486,N_9037,N_9036);
nor UO_1487 (O_1487,N_9763,N_9792);
nor UO_1488 (O_1488,N_9316,N_9775);
xnor UO_1489 (O_1489,N_9958,N_9173);
nand UO_1490 (O_1490,N_9633,N_9598);
xor UO_1491 (O_1491,N_9235,N_9666);
and UO_1492 (O_1492,N_9419,N_9065);
xor UO_1493 (O_1493,N_9444,N_9604);
and UO_1494 (O_1494,N_9383,N_9657);
or UO_1495 (O_1495,N_9072,N_9844);
nand UO_1496 (O_1496,N_9545,N_9148);
or UO_1497 (O_1497,N_9146,N_9691);
or UO_1498 (O_1498,N_9406,N_9590);
and UO_1499 (O_1499,N_9679,N_9124);
endmodule