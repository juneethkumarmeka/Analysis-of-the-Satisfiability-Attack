module basic_500_3000_500_4_levels_2xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_4,In_283);
nand U1 (N_1,In_99,In_329);
nand U2 (N_2,In_141,In_319);
and U3 (N_3,In_46,In_149);
or U4 (N_4,In_164,In_311);
xnor U5 (N_5,In_260,In_350);
nand U6 (N_6,In_72,In_43);
nor U7 (N_7,In_478,In_443);
nor U8 (N_8,In_61,In_40);
or U9 (N_9,In_381,In_460);
or U10 (N_10,In_363,In_490);
nor U11 (N_11,In_318,In_153);
nand U12 (N_12,In_102,In_232);
nand U13 (N_13,In_345,In_454);
or U14 (N_14,In_127,In_304);
nor U15 (N_15,In_261,In_45);
nor U16 (N_16,In_364,In_154);
and U17 (N_17,In_30,In_240);
nor U18 (N_18,In_90,In_208);
or U19 (N_19,In_359,In_385);
nand U20 (N_20,In_471,In_440);
or U21 (N_21,In_75,In_190);
or U22 (N_22,In_248,In_276);
nor U23 (N_23,In_353,In_308);
nand U24 (N_24,In_316,In_129);
or U25 (N_25,In_394,In_2);
nand U26 (N_26,In_122,In_134);
and U27 (N_27,In_230,In_81);
or U28 (N_28,In_335,In_312);
nand U29 (N_29,In_222,In_243);
nand U30 (N_30,In_60,In_26);
or U31 (N_31,In_412,In_136);
nand U32 (N_32,In_434,In_135);
or U33 (N_33,In_441,In_449);
nand U34 (N_34,In_325,In_196);
or U35 (N_35,In_194,In_10);
or U36 (N_36,In_373,In_302);
nand U37 (N_37,In_498,In_126);
nor U38 (N_38,In_27,In_74);
nor U39 (N_39,In_370,In_413);
and U40 (N_40,In_78,In_371);
and U41 (N_41,In_409,In_19);
or U42 (N_42,In_170,In_66);
nor U43 (N_43,In_200,In_417);
nor U44 (N_44,In_266,In_235);
and U45 (N_45,In_431,In_391);
or U46 (N_46,In_393,In_142);
xnor U47 (N_47,In_53,In_357);
nand U48 (N_48,In_201,In_55);
nand U49 (N_49,In_155,In_392);
and U50 (N_50,In_14,In_404);
nor U51 (N_51,In_94,In_267);
or U52 (N_52,In_48,In_207);
nand U53 (N_53,In_202,In_307);
nand U54 (N_54,In_133,In_405);
nand U55 (N_55,In_281,In_358);
nor U56 (N_56,In_263,In_317);
nand U57 (N_57,In_328,In_220);
xnor U58 (N_58,In_44,In_84);
and U59 (N_59,In_466,In_54);
nor U60 (N_60,In_420,In_96);
and U61 (N_61,In_474,In_470);
xnor U62 (N_62,In_477,In_484);
nor U63 (N_63,In_241,In_121);
nand U64 (N_64,In_379,In_303);
or U65 (N_65,In_402,In_425);
and U66 (N_66,In_269,In_157);
nand U67 (N_67,In_86,In_73);
and U68 (N_68,In_399,In_245);
and U69 (N_69,In_337,In_206);
nor U70 (N_70,In_197,In_77);
nor U71 (N_71,In_499,In_396);
and U72 (N_72,In_204,In_192);
and U73 (N_73,In_321,In_17);
and U74 (N_74,In_106,In_233);
nand U75 (N_75,In_16,In_69);
nor U76 (N_76,In_175,In_216);
nor U77 (N_77,In_58,In_25);
or U78 (N_78,In_231,In_429);
nand U79 (N_79,In_457,In_462);
nor U80 (N_80,In_101,In_252);
or U81 (N_81,In_3,In_117);
nand U82 (N_82,In_479,In_91);
nand U83 (N_83,In_18,In_343);
and U84 (N_84,In_287,In_451);
nand U85 (N_85,In_158,In_463);
nor U86 (N_86,In_56,In_298);
or U87 (N_87,In_223,In_377);
nand U88 (N_88,In_296,In_116);
and U89 (N_89,In_254,In_111);
xnor U90 (N_90,In_489,In_203);
and U91 (N_91,In_143,In_493);
nand U92 (N_92,In_182,In_28);
nor U93 (N_93,In_6,In_476);
and U94 (N_94,In_426,In_144);
nor U95 (N_95,In_34,In_124);
or U96 (N_96,In_293,In_218);
or U97 (N_97,In_229,In_76);
and U98 (N_98,In_277,In_137);
nand U99 (N_99,In_314,In_384);
nand U100 (N_100,In_390,In_262);
or U101 (N_101,In_297,In_160);
and U102 (N_102,In_195,In_150);
or U103 (N_103,In_268,In_221);
nand U104 (N_104,In_284,In_33);
nor U105 (N_105,In_369,In_453);
nand U106 (N_106,In_23,In_125);
nor U107 (N_107,In_105,In_423);
nor U108 (N_108,In_242,In_271);
nor U109 (N_109,In_186,In_109);
nand U110 (N_110,In_497,In_419);
or U111 (N_111,In_209,In_52);
or U112 (N_112,In_301,In_382);
nor U113 (N_113,In_225,In_475);
nor U114 (N_114,In_289,In_11);
nand U115 (N_115,In_35,In_20);
nand U116 (N_116,In_305,In_159);
nor U117 (N_117,In_176,In_64);
nor U118 (N_118,In_288,In_444);
xnor U119 (N_119,In_42,In_458);
nand U120 (N_120,In_459,In_187);
nor U121 (N_121,In_421,In_112);
or U122 (N_122,In_51,In_224);
nand U123 (N_123,In_483,In_188);
nor U124 (N_124,In_294,In_47);
or U125 (N_125,In_118,In_88);
or U126 (N_126,In_89,In_217);
nand U127 (N_127,In_146,In_244);
and U128 (N_128,In_342,In_488);
or U129 (N_129,In_5,In_495);
or U130 (N_130,In_180,In_9);
or U131 (N_131,In_67,In_87);
xnor U132 (N_132,In_435,In_279);
nor U133 (N_133,In_171,In_332);
nor U134 (N_134,In_214,In_372);
nor U135 (N_135,In_465,In_278);
nor U136 (N_136,In_226,In_415);
or U137 (N_137,In_433,In_210);
xnor U138 (N_138,In_92,In_388);
nand U139 (N_139,In_365,In_411);
xor U140 (N_140,In_427,In_398);
nand U141 (N_141,In_165,In_8);
nor U142 (N_142,In_0,In_108);
nor U143 (N_143,In_32,In_15);
nand U144 (N_144,In_151,In_185);
nor U145 (N_145,In_336,In_322);
nand U146 (N_146,In_82,In_492);
nor U147 (N_147,In_290,In_383);
and U148 (N_148,In_464,In_401);
or U149 (N_149,In_39,In_324);
or U150 (N_150,In_270,In_282);
nand U151 (N_151,In_424,In_344);
nor U152 (N_152,In_215,In_323);
and U153 (N_153,In_445,In_50);
or U154 (N_154,In_41,In_339);
and U155 (N_155,In_148,In_178);
or U156 (N_156,In_286,In_237);
or U157 (N_157,In_456,In_114);
xnor U158 (N_158,In_367,In_494);
nor U159 (N_159,In_416,In_375);
nor U160 (N_160,In_348,In_309);
nand U161 (N_161,In_128,In_147);
and U162 (N_162,In_264,In_98);
and U163 (N_163,In_249,In_211);
xor U164 (N_164,In_395,In_110);
and U165 (N_165,In_189,In_173);
nor U166 (N_166,In_366,In_448);
or U167 (N_167,In_446,In_113);
or U168 (N_168,In_62,In_300);
and U169 (N_169,In_130,In_438);
or U170 (N_170,In_442,In_486);
nor U171 (N_171,In_291,In_139);
nand U172 (N_172,In_104,In_265);
nor U173 (N_173,In_259,In_496);
nor U174 (N_174,In_80,In_1);
or U175 (N_175,In_400,In_334);
or U176 (N_176,In_360,In_161);
nor U177 (N_177,In_79,In_299);
nor U178 (N_178,In_485,In_455);
and U179 (N_179,In_355,In_12);
or U180 (N_180,In_213,In_21);
and U181 (N_181,In_491,In_29);
nor U182 (N_182,In_156,In_162);
xor U183 (N_183,In_362,In_374);
or U184 (N_184,In_331,In_31);
or U185 (N_185,In_123,In_340);
nand U186 (N_186,In_71,In_472);
or U187 (N_187,In_163,In_275);
nor U188 (N_188,In_473,In_140);
xor U189 (N_189,In_181,In_169);
nor U190 (N_190,In_255,In_132);
nand U191 (N_191,In_83,In_447);
nand U192 (N_192,In_7,In_238);
or U193 (N_193,In_115,In_354);
nand U194 (N_194,In_351,In_172);
nor U195 (N_195,In_418,In_167);
nor U196 (N_196,In_246,In_145);
nor U197 (N_197,In_450,In_481);
nor U198 (N_198,In_97,In_256);
or U199 (N_199,In_13,In_120);
nor U200 (N_200,In_22,In_184);
or U201 (N_201,In_36,In_168);
and U202 (N_202,In_313,In_68);
nand U203 (N_203,In_57,In_205);
nor U204 (N_204,In_349,In_310);
or U205 (N_205,In_378,In_320);
and U206 (N_206,In_253,In_326);
or U207 (N_207,In_280,In_285);
nor U208 (N_208,In_346,In_327);
nand U209 (N_209,In_95,In_152);
xnor U210 (N_210,In_387,In_356);
nor U211 (N_211,In_352,In_250);
and U212 (N_212,In_333,In_70);
or U213 (N_213,In_166,In_452);
or U214 (N_214,In_198,In_487);
or U215 (N_215,In_193,In_469);
and U216 (N_216,In_292,In_37);
or U217 (N_217,In_428,In_397);
nor U218 (N_218,In_376,In_347);
nand U219 (N_219,In_93,In_341);
and U220 (N_220,In_306,In_59);
or U221 (N_221,In_330,In_430);
and U222 (N_222,In_410,In_389);
or U223 (N_223,In_38,In_338);
nand U224 (N_224,In_65,In_258);
nor U225 (N_225,In_131,In_85);
or U226 (N_226,In_422,In_386);
xnor U227 (N_227,In_407,In_247);
nand U228 (N_228,In_49,In_174);
nor U229 (N_229,In_380,In_480);
nor U230 (N_230,In_228,In_179);
or U231 (N_231,In_183,In_403);
nand U232 (N_232,In_467,In_236);
nor U233 (N_233,In_199,In_295);
and U234 (N_234,In_138,In_361);
and U235 (N_235,In_468,In_177);
nor U236 (N_236,In_439,In_212);
nand U237 (N_237,In_119,In_234);
or U238 (N_238,In_100,In_251);
nand U239 (N_239,In_436,In_107);
or U240 (N_240,In_368,In_24);
nand U241 (N_241,In_274,In_219);
and U242 (N_242,In_63,In_227);
and U243 (N_243,In_414,In_461);
or U244 (N_244,In_272,In_482);
nand U245 (N_245,In_257,In_406);
or U246 (N_246,In_239,In_408);
or U247 (N_247,In_191,In_315);
nor U248 (N_248,In_432,In_103);
nand U249 (N_249,In_437,In_273);
nand U250 (N_250,In_246,In_289);
or U251 (N_251,In_32,In_164);
nor U252 (N_252,In_143,In_214);
nand U253 (N_253,In_233,In_162);
or U254 (N_254,In_239,In_399);
nand U255 (N_255,In_300,In_469);
or U256 (N_256,In_474,In_185);
nor U257 (N_257,In_415,In_243);
and U258 (N_258,In_180,In_414);
or U259 (N_259,In_495,In_481);
and U260 (N_260,In_59,In_278);
nand U261 (N_261,In_217,In_468);
or U262 (N_262,In_244,In_443);
or U263 (N_263,In_192,In_59);
or U264 (N_264,In_202,In_363);
nor U265 (N_265,In_160,In_240);
nor U266 (N_266,In_359,In_75);
nor U267 (N_267,In_12,In_275);
and U268 (N_268,In_79,In_360);
nand U269 (N_269,In_434,In_77);
and U270 (N_270,In_388,In_132);
nand U271 (N_271,In_155,In_234);
and U272 (N_272,In_249,In_316);
and U273 (N_273,In_374,In_314);
nand U274 (N_274,In_243,In_86);
and U275 (N_275,In_324,In_101);
nor U276 (N_276,In_199,In_2);
nand U277 (N_277,In_454,In_451);
nor U278 (N_278,In_256,In_368);
nor U279 (N_279,In_201,In_485);
nor U280 (N_280,In_332,In_427);
nor U281 (N_281,In_34,In_350);
nand U282 (N_282,In_118,In_222);
xor U283 (N_283,In_424,In_333);
and U284 (N_284,In_228,In_240);
and U285 (N_285,In_185,In_331);
or U286 (N_286,In_286,In_8);
and U287 (N_287,In_174,In_372);
nand U288 (N_288,In_73,In_193);
and U289 (N_289,In_194,In_2);
and U290 (N_290,In_4,In_407);
nor U291 (N_291,In_475,In_403);
or U292 (N_292,In_87,In_452);
or U293 (N_293,In_385,In_13);
nor U294 (N_294,In_73,In_131);
nor U295 (N_295,In_98,In_448);
nor U296 (N_296,In_459,In_175);
nand U297 (N_297,In_268,In_449);
nor U298 (N_298,In_338,In_218);
nor U299 (N_299,In_192,In_483);
xnor U300 (N_300,In_288,In_409);
nor U301 (N_301,In_0,In_390);
and U302 (N_302,In_415,In_178);
or U303 (N_303,In_170,In_243);
or U304 (N_304,In_232,In_237);
and U305 (N_305,In_136,In_192);
or U306 (N_306,In_482,In_154);
and U307 (N_307,In_72,In_464);
and U308 (N_308,In_144,In_16);
or U309 (N_309,In_45,In_464);
and U310 (N_310,In_5,In_375);
nand U311 (N_311,In_405,In_214);
or U312 (N_312,In_250,In_21);
nor U313 (N_313,In_479,In_367);
nor U314 (N_314,In_360,In_175);
nor U315 (N_315,In_62,In_132);
nand U316 (N_316,In_102,In_149);
or U317 (N_317,In_435,In_101);
nand U318 (N_318,In_358,In_222);
or U319 (N_319,In_447,In_313);
nor U320 (N_320,In_15,In_370);
or U321 (N_321,In_328,In_415);
nand U322 (N_322,In_152,In_330);
nor U323 (N_323,In_321,In_174);
nand U324 (N_324,In_296,In_45);
or U325 (N_325,In_414,In_241);
and U326 (N_326,In_306,In_167);
and U327 (N_327,In_400,In_89);
or U328 (N_328,In_148,In_274);
and U329 (N_329,In_198,In_326);
and U330 (N_330,In_138,In_419);
nor U331 (N_331,In_420,In_341);
nor U332 (N_332,In_419,In_188);
or U333 (N_333,In_64,In_124);
nand U334 (N_334,In_184,In_471);
nor U335 (N_335,In_390,In_421);
nor U336 (N_336,In_174,In_77);
nand U337 (N_337,In_378,In_406);
nand U338 (N_338,In_40,In_50);
nor U339 (N_339,In_201,In_434);
or U340 (N_340,In_399,In_447);
nand U341 (N_341,In_430,In_209);
or U342 (N_342,In_270,In_465);
or U343 (N_343,In_195,In_481);
and U344 (N_344,In_438,In_290);
or U345 (N_345,In_183,In_307);
xnor U346 (N_346,In_179,In_74);
nor U347 (N_347,In_432,In_19);
nand U348 (N_348,In_232,In_112);
or U349 (N_349,In_221,In_235);
or U350 (N_350,In_343,In_68);
nor U351 (N_351,In_237,In_343);
or U352 (N_352,In_140,In_279);
and U353 (N_353,In_32,In_241);
or U354 (N_354,In_494,In_457);
or U355 (N_355,In_430,In_236);
nand U356 (N_356,In_287,In_127);
nor U357 (N_357,In_53,In_267);
nor U358 (N_358,In_276,In_284);
nand U359 (N_359,In_170,In_307);
or U360 (N_360,In_42,In_462);
or U361 (N_361,In_209,In_177);
nand U362 (N_362,In_403,In_63);
and U363 (N_363,In_27,In_248);
or U364 (N_364,In_212,In_344);
nor U365 (N_365,In_346,In_76);
or U366 (N_366,In_130,In_108);
and U367 (N_367,In_11,In_269);
nand U368 (N_368,In_190,In_117);
nor U369 (N_369,In_293,In_379);
or U370 (N_370,In_172,In_310);
or U371 (N_371,In_334,In_339);
nand U372 (N_372,In_9,In_466);
xor U373 (N_373,In_352,In_129);
and U374 (N_374,In_227,In_200);
or U375 (N_375,In_322,In_203);
nand U376 (N_376,In_156,In_227);
nand U377 (N_377,In_115,In_65);
or U378 (N_378,In_403,In_367);
and U379 (N_379,In_241,In_327);
nand U380 (N_380,In_304,In_294);
and U381 (N_381,In_483,In_208);
xnor U382 (N_382,In_440,In_418);
and U383 (N_383,In_26,In_357);
nand U384 (N_384,In_139,In_295);
nor U385 (N_385,In_425,In_386);
nand U386 (N_386,In_6,In_5);
nor U387 (N_387,In_140,In_402);
nor U388 (N_388,In_340,In_329);
nand U389 (N_389,In_200,In_194);
nand U390 (N_390,In_62,In_259);
nor U391 (N_391,In_390,In_8);
and U392 (N_392,In_17,In_439);
nor U393 (N_393,In_139,In_281);
nor U394 (N_394,In_45,In_330);
nand U395 (N_395,In_110,In_448);
nand U396 (N_396,In_444,In_287);
nand U397 (N_397,In_442,In_166);
and U398 (N_398,In_46,In_399);
nand U399 (N_399,In_260,In_407);
or U400 (N_400,In_331,In_306);
nand U401 (N_401,In_11,In_403);
and U402 (N_402,In_399,In_427);
or U403 (N_403,In_165,In_157);
nor U404 (N_404,In_351,In_400);
nand U405 (N_405,In_112,In_171);
or U406 (N_406,In_186,In_231);
nand U407 (N_407,In_476,In_210);
and U408 (N_408,In_42,In_179);
and U409 (N_409,In_162,In_1);
nand U410 (N_410,In_134,In_252);
xor U411 (N_411,In_55,In_418);
or U412 (N_412,In_264,In_256);
nor U413 (N_413,In_354,In_105);
and U414 (N_414,In_495,In_425);
or U415 (N_415,In_365,In_444);
and U416 (N_416,In_108,In_288);
nor U417 (N_417,In_79,In_232);
or U418 (N_418,In_144,In_455);
nand U419 (N_419,In_221,In_95);
and U420 (N_420,In_177,In_291);
and U421 (N_421,In_352,In_498);
nand U422 (N_422,In_105,In_495);
and U423 (N_423,In_88,In_376);
nand U424 (N_424,In_381,In_275);
and U425 (N_425,In_113,In_462);
nor U426 (N_426,In_64,In_483);
nand U427 (N_427,In_375,In_186);
or U428 (N_428,In_270,In_31);
or U429 (N_429,In_388,In_211);
or U430 (N_430,In_436,In_74);
and U431 (N_431,In_224,In_196);
or U432 (N_432,In_216,In_166);
or U433 (N_433,In_446,In_14);
nor U434 (N_434,In_422,In_134);
or U435 (N_435,In_362,In_496);
or U436 (N_436,In_206,In_456);
and U437 (N_437,In_55,In_21);
nand U438 (N_438,In_18,In_61);
nand U439 (N_439,In_315,In_480);
nor U440 (N_440,In_27,In_297);
nand U441 (N_441,In_18,In_81);
or U442 (N_442,In_228,In_352);
and U443 (N_443,In_113,In_201);
or U444 (N_444,In_94,In_176);
and U445 (N_445,In_318,In_300);
nor U446 (N_446,In_480,In_361);
nand U447 (N_447,In_59,In_85);
nand U448 (N_448,In_34,In_245);
or U449 (N_449,In_354,In_301);
nor U450 (N_450,In_296,In_92);
and U451 (N_451,In_354,In_203);
nand U452 (N_452,In_496,In_275);
or U453 (N_453,In_425,In_32);
and U454 (N_454,In_325,In_207);
and U455 (N_455,In_165,In_49);
nand U456 (N_456,In_54,In_363);
nor U457 (N_457,In_265,In_116);
or U458 (N_458,In_63,In_28);
and U459 (N_459,In_288,In_354);
nand U460 (N_460,In_418,In_261);
nor U461 (N_461,In_257,In_237);
or U462 (N_462,In_23,In_275);
nand U463 (N_463,In_314,In_288);
and U464 (N_464,In_297,In_294);
nor U465 (N_465,In_279,In_445);
and U466 (N_466,In_493,In_361);
or U467 (N_467,In_39,In_208);
or U468 (N_468,In_241,In_60);
and U469 (N_469,In_229,In_151);
nor U470 (N_470,In_480,In_270);
nor U471 (N_471,In_455,In_474);
nor U472 (N_472,In_479,In_355);
nand U473 (N_473,In_306,In_291);
and U474 (N_474,In_196,In_489);
nor U475 (N_475,In_113,In_251);
nand U476 (N_476,In_171,In_486);
and U477 (N_477,In_133,In_372);
or U478 (N_478,In_203,In_191);
or U479 (N_479,In_138,In_308);
nor U480 (N_480,In_431,In_150);
nand U481 (N_481,In_22,In_42);
nand U482 (N_482,In_445,In_305);
nor U483 (N_483,In_189,In_360);
nand U484 (N_484,In_388,In_380);
nand U485 (N_485,In_310,In_373);
and U486 (N_486,In_476,In_332);
nor U487 (N_487,In_217,In_125);
or U488 (N_488,In_363,In_259);
nand U489 (N_489,In_148,In_426);
nand U490 (N_490,In_352,In_213);
and U491 (N_491,In_254,In_465);
and U492 (N_492,In_226,In_301);
nor U493 (N_493,In_296,In_255);
nor U494 (N_494,In_24,In_14);
nand U495 (N_495,In_253,In_29);
or U496 (N_496,In_204,In_54);
or U497 (N_497,In_209,In_293);
nor U498 (N_498,In_348,In_251);
nor U499 (N_499,In_266,In_464);
nor U500 (N_500,In_352,In_478);
and U501 (N_501,In_262,In_156);
nand U502 (N_502,In_246,In_237);
nor U503 (N_503,In_24,In_354);
or U504 (N_504,In_180,In_48);
nor U505 (N_505,In_20,In_220);
nand U506 (N_506,In_460,In_309);
nand U507 (N_507,In_285,In_79);
nand U508 (N_508,In_25,In_143);
nand U509 (N_509,In_388,In_397);
nor U510 (N_510,In_330,In_269);
nor U511 (N_511,In_367,In_62);
nor U512 (N_512,In_357,In_224);
and U513 (N_513,In_365,In_203);
nand U514 (N_514,In_154,In_257);
or U515 (N_515,In_321,In_496);
and U516 (N_516,In_460,In_340);
nor U517 (N_517,In_208,In_232);
nand U518 (N_518,In_170,In_297);
or U519 (N_519,In_172,In_184);
and U520 (N_520,In_276,In_279);
and U521 (N_521,In_257,In_339);
or U522 (N_522,In_188,In_404);
and U523 (N_523,In_170,In_178);
nand U524 (N_524,In_396,In_164);
or U525 (N_525,In_91,In_330);
or U526 (N_526,In_356,In_108);
nand U527 (N_527,In_349,In_154);
or U528 (N_528,In_134,In_272);
nor U529 (N_529,In_160,In_389);
nor U530 (N_530,In_236,In_83);
nor U531 (N_531,In_22,In_155);
or U532 (N_532,In_243,In_117);
nand U533 (N_533,In_157,In_332);
and U534 (N_534,In_27,In_410);
nand U535 (N_535,In_72,In_56);
nand U536 (N_536,In_12,In_22);
nor U537 (N_537,In_220,In_458);
nor U538 (N_538,In_145,In_478);
or U539 (N_539,In_375,In_213);
nand U540 (N_540,In_310,In_288);
or U541 (N_541,In_403,In_277);
or U542 (N_542,In_432,In_383);
nand U543 (N_543,In_371,In_156);
nand U544 (N_544,In_320,In_262);
and U545 (N_545,In_281,In_37);
and U546 (N_546,In_259,In_261);
and U547 (N_547,In_143,In_47);
nand U548 (N_548,In_361,In_319);
nor U549 (N_549,In_106,In_89);
and U550 (N_550,In_191,In_290);
and U551 (N_551,In_377,In_294);
or U552 (N_552,In_254,In_455);
nor U553 (N_553,In_230,In_369);
nand U554 (N_554,In_239,In_311);
nand U555 (N_555,In_62,In_270);
and U556 (N_556,In_442,In_50);
nand U557 (N_557,In_369,In_170);
nand U558 (N_558,In_158,In_9);
nor U559 (N_559,In_18,In_432);
or U560 (N_560,In_29,In_131);
nand U561 (N_561,In_300,In_103);
nand U562 (N_562,In_202,In_386);
and U563 (N_563,In_414,In_79);
nor U564 (N_564,In_267,In_159);
and U565 (N_565,In_171,In_294);
nor U566 (N_566,In_199,In_48);
nand U567 (N_567,In_443,In_247);
or U568 (N_568,In_235,In_499);
and U569 (N_569,In_49,In_217);
nor U570 (N_570,In_410,In_406);
nor U571 (N_571,In_274,In_467);
nor U572 (N_572,In_369,In_439);
nor U573 (N_573,In_153,In_254);
or U574 (N_574,In_262,In_406);
nand U575 (N_575,In_238,In_370);
and U576 (N_576,In_415,In_214);
or U577 (N_577,In_370,In_333);
or U578 (N_578,In_284,In_247);
nand U579 (N_579,In_449,In_325);
nand U580 (N_580,In_127,In_183);
nand U581 (N_581,In_210,In_460);
or U582 (N_582,In_13,In_429);
or U583 (N_583,In_357,In_244);
xor U584 (N_584,In_121,In_388);
and U585 (N_585,In_401,In_267);
nand U586 (N_586,In_157,In_54);
nor U587 (N_587,In_432,In_425);
nand U588 (N_588,In_27,In_384);
nor U589 (N_589,In_279,In_110);
nor U590 (N_590,In_399,In_276);
and U591 (N_591,In_200,In_71);
nand U592 (N_592,In_453,In_170);
and U593 (N_593,In_121,In_202);
and U594 (N_594,In_139,In_156);
nand U595 (N_595,In_163,In_171);
nor U596 (N_596,In_235,In_466);
nor U597 (N_597,In_146,In_320);
nand U598 (N_598,In_11,In_392);
or U599 (N_599,In_224,In_232);
nor U600 (N_600,In_312,In_139);
nor U601 (N_601,In_254,In_464);
nand U602 (N_602,In_449,In_213);
and U603 (N_603,In_334,In_96);
nand U604 (N_604,In_370,In_462);
and U605 (N_605,In_161,In_398);
nand U606 (N_606,In_225,In_139);
nand U607 (N_607,In_99,In_320);
nor U608 (N_608,In_33,In_244);
xnor U609 (N_609,In_33,In_277);
and U610 (N_610,In_12,In_426);
nand U611 (N_611,In_90,In_130);
or U612 (N_612,In_405,In_170);
or U613 (N_613,In_306,In_416);
nor U614 (N_614,In_290,In_160);
xnor U615 (N_615,In_207,In_223);
nor U616 (N_616,In_221,In_322);
and U617 (N_617,In_472,In_165);
nand U618 (N_618,In_309,In_288);
or U619 (N_619,In_421,In_276);
and U620 (N_620,In_106,In_145);
and U621 (N_621,In_307,In_312);
or U622 (N_622,In_299,In_176);
nor U623 (N_623,In_283,In_272);
and U624 (N_624,In_450,In_485);
or U625 (N_625,In_439,In_183);
and U626 (N_626,In_262,In_337);
nor U627 (N_627,In_395,In_407);
or U628 (N_628,In_119,In_439);
nor U629 (N_629,In_364,In_398);
and U630 (N_630,In_335,In_27);
and U631 (N_631,In_291,In_171);
and U632 (N_632,In_251,In_487);
nand U633 (N_633,In_53,In_72);
or U634 (N_634,In_235,In_173);
or U635 (N_635,In_25,In_292);
nor U636 (N_636,In_224,In_197);
nand U637 (N_637,In_354,In_343);
nor U638 (N_638,In_39,In_42);
nand U639 (N_639,In_149,In_135);
and U640 (N_640,In_288,In_266);
nor U641 (N_641,In_42,In_313);
nor U642 (N_642,In_195,In_118);
nor U643 (N_643,In_347,In_37);
nand U644 (N_644,In_407,In_211);
nor U645 (N_645,In_3,In_66);
nor U646 (N_646,In_285,In_363);
xor U647 (N_647,In_58,In_207);
nand U648 (N_648,In_252,In_28);
or U649 (N_649,In_278,In_41);
nor U650 (N_650,In_297,In_51);
or U651 (N_651,In_152,In_99);
nand U652 (N_652,In_46,In_205);
and U653 (N_653,In_313,In_462);
nand U654 (N_654,In_50,In_109);
or U655 (N_655,In_120,In_287);
and U656 (N_656,In_144,In_67);
and U657 (N_657,In_153,In_73);
nor U658 (N_658,In_148,In_18);
and U659 (N_659,In_465,In_275);
nor U660 (N_660,In_455,In_440);
or U661 (N_661,In_293,In_156);
nor U662 (N_662,In_442,In_437);
nor U663 (N_663,In_364,In_54);
and U664 (N_664,In_40,In_308);
xor U665 (N_665,In_100,In_86);
nor U666 (N_666,In_403,In_323);
and U667 (N_667,In_493,In_442);
nor U668 (N_668,In_208,In_84);
nand U669 (N_669,In_459,In_403);
nor U670 (N_670,In_76,In_370);
nor U671 (N_671,In_57,In_293);
and U672 (N_672,In_211,In_125);
nand U673 (N_673,In_47,In_475);
or U674 (N_674,In_359,In_448);
and U675 (N_675,In_158,In_412);
or U676 (N_676,In_267,In_493);
nor U677 (N_677,In_223,In_424);
or U678 (N_678,In_395,In_376);
xnor U679 (N_679,In_473,In_378);
nor U680 (N_680,In_152,In_380);
nand U681 (N_681,In_360,In_84);
nor U682 (N_682,In_16,In_375);
nor U683 (N_683,In_115,In_218);
and U684 (N_684,In_493,In_457);
nor U685 (N_685,In_66,In_477);
or U686 (N_686,In_400,In_486);
nor U687 (N_687,In_482,In_144);
or U688 (N_688,In_395,In_31);
and U689 (N_689,In_340,In_235);
or U690 (N_690,In_330,In_102);
and U691 (N_691,In_343,In_311);
or U692 (N_692,In_17,In_336);
nand U693 (N_693,In_498,In_9);
nor U694 (N_694,In_280,In_241);
and U695 (N_695,In_7,In_381);
or U696 (N_696,In_64,In_443);
nor U697 (N_697,In_116,In_458);
nand U698 (N_698,In_198,In_482);
nand U699 (N_699,In_201,In_488);
nand U700 (N_700,In_221,In_280);
or U701 (N_701,In_250,In_88);
nand U702 (N_702,In_98,In_62);
and U703 (N_703,In_3,In_63);
nor U704 (N_704,In_326,In_160);
nor U705 (N_705,In_388,In_486);
nand U706 (N_706,In_195,In_235);
nor U707 (N_707,In_38,In_98);
and U708 (N_708,In_144,In_254);
and U709 (N_709,In_302,In_398);
or U710 (N_710,In_452,In_176);
or U711 (N_711,In_454,In_93);
or U712 (N_712,In_248,In_224);
and U713 (N_713,In_297,In_189);
nor U714 (N_714,In_60,In_149);
nor U715 (N_715,In_31,In_418);
or U716 (N_716,In_499,In_4);
or U717 (N_717,In_64,In_248);
nand U718 (N_718,In_279,In_306);
or U719 (N_719,In_402,In_420);
nand U720 (N_720,In_375,In_206);
nand U721 (N_721,In_282,In_312);
or U722 (N_722,In_174,In_186);
and U723 (N_723,In_40,In_269);
or U724 (N_724,In_121,In_381);
or U725 (N_725,In_66,In_244);
nand U726 (N_726,In_231,In_44);
or U727 (N_727,In_95,In_270);
and U728 (N_728,In_109,In_344);
or U729 (N_729,In_97,In_340);
and U730 (N_730,In_174,In_69);
nor U731 (N_731,In_157,In_254);
nor U732 (N_732,In_429,In_487);
nor U733 (N_733,In_32,In_53);
nand U734 (N_734,In_394,In_302);
nand U735 (N_735,In_252,In_330);
and U736 (N_736,In_267,In_413);
and U737 (N_737,In_205,In_119);
or U738 (N_738,In_349,In_254);
nor U739 (N_739,In_308,In_240);
nor U740 (N_740,In_3,In_411);
nor U741 (N_741,In_219,In_161);
nand U742 (N_742,In_441,In_314);
nand U743 (N_743,In_229,In_258);
nand U744 (N_744,In_241,In_300);
and U745 (N_745,In_467,In_175);
or U746 (N_746,In_91,In_257);
and U747 (N_747,In_240,In_68);
nand U748 (N_748,In_361,In_300);
and U749 (N_749,In_160,In_127);
and U750 (N_750,N_437,N_108);
or U751 (N_751,N_36,N_512);
nor U752 (N_752,N_454,N_481);
nand U753 (N_753,N_217,N_245);
and U754 (N_754,N_392,N_278);
nor U755 (N_755,N_148,N_327);
and U756 (N_756,N_55,N_310);
xnor U757 (N_757,N_445,N_339);
and U758 (N_758,N_220,N_233);
nand U759 (N_759,N_328,N_60);
and U760 (N_760,N_656,N_42);
xor U761 (N_761,N_8,N_336);
or U762 (N_762,N_645,N_133);
and U763 (N_763,N_492,N_222);
nor U764 (N_764,N_58,N_582);
and U765 (N_765,N_37,N_560);
or U766 (N_766,N_557,N_265);
or U767 (N_767,N_539,N_1);
or U768 (N_768,N_580,N_568);
or U769 (N_769,N_517,N_116);
nand U770 (N_770,N_349,N_446);
and U771 (N_771,N_204,N_367);
nor U772 (N_772,N_490,N_257);
xor U773 (N_773,N_718,N_246);
and U774 (N_774,N_375,N_681);
and U775 (N_775,N_166,N_597);
and U776 (N_776,N_225,N_387);
nand U777 (N_777,N_617,N_173);
nand U778 (N_778,N_659,N_156);
nor U779 (N_779,N_514,N_138);
nand U780 (N_780,N_348,N_22);
nand U781 (N_781,N_67,N_502);
and U782 (N_782,N_311,N_444);
nand U783 (N_783,N_425,N_559);
or U784 (N_784,N_322,N_356);
and U785 (N_785,N_149,N_118);
and U786 (N_786,N_408,N_88);
nor U787 (N_787,N_203,N_353);
or U788 (N_788,N_530,N_704);
and U789 (N_789,N_441,N_178);
nand U790 (N_790,N_23,N_41);
and U791 (N_791,N_355,N_135);
nand U792 (N_792,N_293,N_125);
and U793 (N_793,N_3,N_240);
and U794 (N_794,N_563,N_124);
nor U795 (N_795,N_43,N_50);
nand U796 (N_796,N_686,N_500);
nor U797 (N_797,N_341,N_301);
nand U798 (N_798,N_259,N_72);
or U799 (N_799,N_654,N_377);
nand U800 (N_800,N_325,N_176);
and U801 (N_801,N_611,N_529);
or U802 (N_802,N_522,N_131);
nand U803 (N_803,N_722,N_417);
or U804 (N_804,N_267,N_198);
xnor U805 (N_805,N_675,N_600);
nor U806 (N_806,N_456,N_360);
nor U807 (N_807,N_308,N_243);
or U808 (N_808,N_621,N_403);
and U809 (N_809,N_82,N_147);
and U810 (N_810,N_448,N_52);
and U811 (N_811,N_612,N_513);
and U812 (N_812,N_239,N_61);
and U813 (N_813,N_396,N_282);
and U814 (N_814,N_122,N_33);
and U815 (N_815,N_383,N_682);
xor U816 (N_816,N_496,N_478);
nand U817 (N_817,N_2,N_17);
nand U818 (N_818,N_343,N_13);
or U819 (N_819,N_29,N_488);
nor U820 (N_820,N_713,N_555);
and U821 (N_821,N_197,N_184);
nand U822 (N_822,N_56,N_30);
and U823 (N_823,N_525,N_276);
nor U824 (N_824,N_45,N_501);
and U825 (N_825,N_601,N_489);
and U826 (N_826,N_350,N_721);
and U827 (N_827,N_110,N_470);
nor U828 (N_828,N_191,N_273);
and U829 (N_829,N_141,N_683);
or U830 (N_830,N_119,N_380);
nor U831 (N_831,N_648,N_196);
or U832 (N_832,N_223,N_162);
nor U833 (N_833,N_723,N_26);
or U834 (N_834,N_104,N_661);
or U835 (N_835,N_81,N_363);
and U836 (N_836,N_618,N_77);
xor U837 (N_837,N_602,N_741);
xnor U838 (N_838,N_726,N_369);
or U839 (N_839,N_542,N_344);
and U840 (N_840,N_635,N_73);
and U841 (N_841,N_241,N_554);
xnor U842 (N_842,N_109,N_614);
nand U843 (N_843,N_66,N_113);
and U844 (N_844,N_609,N_290);
nor U845 (N_845,N_193,N_494);
nand U846 (N_846,N_691,N_743);
xnor U847 (N_847,N_631,N_440);
nor U848 (N_848,N_511,N_711);
nor U849 (N_849,N_676,N_351);
xor U850 (N_850,N_404,N_183);
and U851 (N_851,N_487,N_486);
or U852 (N_852,N_588,N_651);
nand U853 (N_853,N_309,N_587);
nor U854 (N_854,N_701,N_274);
or U855 (N_855,N_291,N_213);
nand U856 (N_856,N_376,N_594);
nor U857 (N_857,N_620,N_318);
and U858 (N_858,N_634,N_320);
and U859 (N_859,N_411,N_572);
or U860 (N_860,N_99,N_40);
or U861 (N_861,N_163,N_584);
nor U862 (N_862,N_698,N_644);
or U863 (N_863,N_628,N_570);
nand U864 (N_864,N_79,N_16);
nor U865 (N_865,N_10,N_117);
nor U866 (N_866,N_419,N_664);
and U867 (N_867,N_666,N_364);
and U868 (N_868,N_637,N_463);
and U869 (N_869,N_315,N_248);
or U870 (N_870,N_194,N_0);
nor U871 (N_871,N_564,N_158);
or U872 (N_872,N_665,N_192);
and U873 (N_873,N_283,N_548);
nor U874 (N_874,N_471,N_429);
nand U875 (N_875,N_253,N_385);
nor U876 (N_876,N_268,N_696);
and U877 (N_877,N_249,N_358);
nand U878 (N_878,N_716,N_205);
or U879 (N_879,N_107,N_256);
and U880 (N_880,N_640,N_672);
nor U881 (N_881,N_608,N_745);
and U882 (N_882,N_703,N_407);
or U883 (N_883,N_168,N_70);
nor U884 (N_884,N_468,N_98);
nor U885 (N_885,N_669,N_319);
nand U886 (N_886,N_679,N_323);
and U887 (N_887,N_516,N_483);
or U888 (N_888,N_78,N_238);
nand U889 (N_889,N_647,N_549);
nor U890 (N_890,N_366,N_532);
xor U891 (N_891,N_730,N_657);
and U892 (N_892,N_134,N_409);
and U893 (N_893,N_707,N_451);
nor U894 (N_894,N_174,N_93);
or U895 (N_895,N_544,N_578);
nand U896 (N_896,N_335,N_575);
or U897 (N_897,N_457,N_345);
and U898 (N_898,N_473,N_466);
nand U899 (N_899,N_458,N_215);
nand U900 (N_900,N_432,N_673);
nand U901 (N_901,N_386,N_632);
nand U902 (N_902,N_298,N_452);
nor U903 (N_903,N_434,N_221);
nor U904 (N_904,N_537,N_449);
or U905 (N_905,N_476,N_735);
nor U906 (N_906,N_284,N_209);
nand U907 (N_907,N_354,N_155);
nand U908 (N_908,N_330,N_394);
xor U909 (N_909,N_83,N_151);
nor U910 (N_910,N_433,N_201);
nor U911 (N_911,N_297,N_262);
nand U912 (N_912,N_97,N_625);
or U913 (N_913,N_210,N_615);
or U914 (N_914,N_80,N_269);
or U915 (N_915,N_674,N_84);
nand U916 (N_916,N_279,N_579);
or U917 (N_917,N_467,N_700);
nand U918 (N_918,N_391,N_303);
nand U919 (N_919,N_21,N_129);
or U920 (N_920,N_534,N_46);
nand U921 (N_921,N_300,N_485);
nor U922 (N_922,N_251,N_214);
nor U923 (N_923,N_27,N_410);
nor U924 (N_924,N_599,N_406);
or U925 (N_925,N_19,N_106);
or U926 (N_926,N_314,N_729);
nor U927 (N_927,N_736,N_447);
and U928 (N_928,N_480,N_724);
nor U929 (N_929,N_571,N_641);
nand U930 (N_930,N_38,N_188);
nand U931 (N_931,N_663,N_179);
and U932 (N_932,N_229,N_331);
and U933 (N_933,N_581,N_379);
nand U934 (N_934,N_312,N_164);
nand U935 (N_935,N_420,N_543);
or U936 (N_936,N_127,N_232);
and U937 (N_937,N_299,N_321);
nor U938 (N_938,N_551,N_405);
and U939 (N_939,N_727,N_623);
or U940 (N_940,N_275,N_206);
nand U941 (N_941,N_157,N_426);
and U942 (N_942,N_655,N_114);
or U943 (N_943,N_287,N_96);
or U944 (N_944,N_15,N_550);
nor U945 (N_945,N_535,N_677);
nor U946 (N_946,N_509,N_428);
nand U947 (N_947,N_748,N_424);
nand U948 (N_948,N_59,N_541);
or U949 (N_949,N_725,N_658);
nor U950 (N_950,N_585,N_622);
or U951 (N_951,N_636,N_576);
nor U952 (N_952,N_705,N_591);
nand U953 (N_953,N_398,N_167);
and U954 (N_954,N_740,N_236);
nand U955 (N_955,N_527,N_746);
and U956 (N_956,N_520,N_305);
and U957 (N_957,N_62,N_461);
nand U958 (N_958,N_140,N_553);
or U959 (N_959,N_31,N_90);
or U960 (N_960,N_402,N_639);
or U961 (N_961,N_68,N_606);
and U962 (N_962,N_695,N_684);
or U963 (N_963,N_296,N_261);
or U964 (N_964,N_629,N_250);
or U965 (N_965,N_733,N_277);
nand U966 (N_966,N_749,N_498);
and U967 (N_967,N_561,N_32);
xor U968 (N_968,N_732,N_258);
and U969 (N_969,N_49,N_190);
nor U970 (N_970,N_728,N_381);
nand U971 (N_971,N_373,N_14);
and U972 (N_972,N_263,N_720);
or U973 (N_973,N_175,N_742);
and U974 (N_974,N_415,N_4);
and U975 (N_975,N_393,N_226);
nand U976 (N_976,N_123,N_207);
or U977 (N_977,N_172,N_583);
nor U978 (N_978,N_247,N_706);
or U979 (N_979,N_289,N_271);
nand U980 (N_980,N_523,N_412);
and U981 (N_981,N_304,N_547);
or U982 (N_982,N_382,N_493);
nor U983 (N_983,N_649,N_101);
nor U984 (N_984,N_619,N_57);
nor U985 (N_985,N_159,N_285);
or U986 (N_986,N_567,N_738);
or U987 (N_987,N_89,N_211);
nand U988 (N_988,N_423,N_459);
nand U989 (N_989,N_421,N_199);
nand U990 (N_990,N_624,N_182);
nor U991 (N_991,N_528,N_145);
and U992 (N_992,N_177,N_688);
nor U993 (N_993,N_616,N_714);
and U994 (N_994,N_689,N_627);
or U995 (N_995,N_510,N_401);
and U996 (N_996,N_633,N_272);
and U997 (N_997,N_662,N_186);
or U998 (N_998,N_266,N_195);
or U999 (N_999,N_388,N_422);
and U1000 (N_1000,N_418,N_255);
and U1001 (N_1001,N_180,N_242);
or U1002 (N_1002,N_264,N_590);
nand U1003 (N_1003,N_592,N_613);
or U1004 (N_1004,N_34,N_717);
and U1005 (N_1005,N_48,N_39);
nand U1006 (N_1006,N_111,N_450);
xnor U1007 (N_1007,N_566,N_302);
nand U1008 (N_1008,N_260,N_455);
nand U1009 (N_1009,N_715,N_643);
nand U1010 (N_1010,N_413,N_552);
or U1011 (N_1011,N_333,N_646);
nand U1012 (N_1012,N_126,N_130);
nor U1013 (N_1013,N_737,N_593);
or U1014 (N_1014,N_165,N_115);
nand U1015 (N_1015,N_362,N_216);
nand U1016 (N_1016,N_538,N_218);
nand U1017 (N_1017,N_150,N_187);
nand U1018 (N_1018,N_153,N_63);
and U1019 (N_1019,N_252,N_105);
or U1020 (N_1020,N_292,N_556);
nor U1021 (N_1021,N_395,N_281);
or U1022 (N_1022,N_94,N_143);
nor U1023 (N_1023,N_306,N_650);
nand U1024 (N_1024,N_638,N_464);
nor U1025 (N_1025,N_462,N_6);
and U1026 (N_1026,N_660,N_694);
or U1027 (N_1027,N_202,N_161);
and U1028 (N_1028,N_230,N_25);
nand U1029 (N_1029,N_479,N_65);
nor U1030 (N_1030,N_497,N_365);
nor U1031 (N_1031,N_219,N_687);
and U1032 (N_1032,N_169,N_508);
xnor U1033 (N_1033,N_69,N_7);
or U1034 (N_1034,N_630,N_565);
nand U1035 (N_1035,N_372,N_137);
or U1036 (N_1036,N_712,N_121);
and U1037 (N_1037,N_670,N_35);
or U1038 (N_1038,N_697,N_189);
nor U1039 (N_1039,N_626,N_453);
or U1040 (N_1040,N_231,N_680);
nor U1041 (N_1041,N_295,N_503);
or U1042 (N_1042,N_54,N_739);
nand U1043 (N_1043,N_499,N_334);
nor U1044 (N_1044,N_469,N_504);
nor U1045 (N_1045,N_361,N_51);
or U1046 (N_1046,N_595,N_5);
or U1047 (N_1047,N_546,N_690);
and U1048 (N_1048,N_228,N_224);
nand U1049 (N_1049,N_235,N_416);
nor U1050 (N_1050,N_342,N_340);
or U1051 (N_1051,N_678,N_120);
and U1052 (N_1052,N_317,N_74);
nor U1053 (N_1053,N_536,N_146);
xor U1054 (N_1054,N_465,N_573);
nor U1055 (N_1055,N_671,N_438);
nand U1056 (N_1056,N_574,N_431);
and U1057 (N_1057,N_87,N_144);
or U1058 (N_1058,N_435,N_472);
and U1059 (N_1059,N_347,N_170);
or U1060 (N_1060,N_47,N_132);
and U1061 (N_1061,N_286,N_76);
nand U1062 (N_1062,N_185,N_491);
nor U1063 (N_1063,N_474,N_526);
and U1064 (N_1064,N_234,N_521);
nand U1065 (N_1065,N_324,N_316);
and U1066 (N_1066,N_92,N_100);
nor U1067 (N_1067,N_524,N_400);
nor U1068 (N_1068,N_598,N_288);
xnor U1069 (N_1069,N_731,N_53);
and U1070 (N_1070,N_569,N_142);
nor U1071 (N_1071,N_477,N_227);
or U1072 (N_1072,N_152,N_589);
nand U1073 (N_1073,N_495,N_280);
or U1074 (N_1074,N_352,N_443);
and U1075 (N_1075,N_603,N_531);
or U1076 (N_1076,N_747,N_371);
and U1077 (N_1077,N_519,N_693);
and U1078 (N_1078,N_160,N_653);
nand U1079 (N_1079,N_128,N_692);
nor U1080 (N_1080,N_610,N_702);
and U1081 (N_1081,N_540,N_294);
nor U1082 (N_1082,N_337,N_28);
or U1083 (N_1083,N_313,N_436);
and U1084 (N_1084,N_709,N_346);
nand U1085 (N_1085,N_154,N_667);
or U1086 (N_1086,N_484,N_719);
nand U1087 (N_1087,N_642,N_208);
and U1088 (N_1088,N_326,N_103);
or U1089 (N_1089,N_710,N_399);
nor U1090 (N_1090,N_475,N_439);
and U1091 (N_1091,N_482,N_545);
nand U1092 (N_1092,N_685,N_11);
xnor U1093 (N_1093,N_378,N_85);
and U1094 (N_1094,N_586,N_181);
nand U1095 (N_1095,N_577,N_427);
nand U1096 (N_1096,N_505,N_558);
and U1097 (N_1097,N_44,N_390);
or U1098 (N_1098,N_112,N_518);
nor U1099 (N_1099,N_734,N_368);
nor U1100 (N_1100,N_270,N_374);
xor U1101 (N_1101,N_430,N_384);
and U1102 (N_1102,N_102,N_200);
nor U1103 (N_1103,N_442,N_237);
nor U1104 (N_1104,N_64,N_332);
or U1105 (N_1105,N_389,N_708);
or U1106 (N_1106,N_71,N_95);
nand U1107 (N_1107,N_515,N_357);
or U1108 (N_1108,N_18,N_652);
and U1109 (N_1109,N_596,N_397);
or U1110 (N_1110,N_507,N_86);
or U1111 (N_1111,N_244,N_414);
nand U1112 (N_1112,N_171,N_254);
or U1113 (N_1113,N_307,N_24);
nor U1114 (N_1114,N_506,N_136);
nor U1115 (N_1115,N_562,N_91);
and U1116 (N_1116,N_75,N_699);
and U1117 (N_1117,N_533,N_9);
nand U1118 (N_1118,N_604,N_607);
nor U1119 (N_1119,N_744,N_359);
nand U1120 (N_1120,N_460,N_12);
nand U1121 (N_1121,N_329,N_370);
and U1122 (N_1122,N_668,N_139);
and U1123 (N_1123,N_338,N_20);
xor U1124 (N_1124,N_605,N_212);
nand U1125 (N_1125,N_570,N_413);
and U1126 (N_1126,N_438,N_398);
xnor U1127 (N_1127,N_288,N_540);
and U1128 (N_1128,N_745,N_155);
or U1129 (N_1129,N_652,N_721);
and U1130 (N_1130,N_56,N_676);
nor U1131 (N_1131,N_692,N_713);
nor U1132 (N_1132,N_668,N_556);
or U1133 (N_1133,N_433,N_690);
and U1134 (N_1134,N_409,N_402);
nor U1135 (N_1135,N_42,N_215);
nand U1136 (N_1136,N_625,N_222);
nor U1137 (N_1137,N_43,N_603);
nand U1138 (N_1138,N_157,N_177);
or U1139 (N_1139,N_12,N_650);
nor U1140 (N_1140,N_274,N_732);
and U1141 (N_1141,N_422,N_653);
or U1142 (N_1142,N_73,N_480);
or U1143 (N_1143,N_325,N_500);
or U1144 (N_1144,N_105,N_148);
nand U1145 (N_1145,N_680,N_335);
or U1146 (N_1146,N_56,N_719);
or U1147 (N_1147,N_479,N_378);
and U1148 (N_1148,N_344,N_70);
or U1149 (N_1149,N_438,N_49);
or U1150 (N_1150,N_105,N_185);
and U1151 (N_1151,N_109,N_683);
nand U1152 (N_1152,N_507,N_623);
and U1153 (N_1153,N_243,N_557);
nand U1154 (N_1154,N_160,N_186);
and U1155 (N_1155,N_93,N_168);
nand U1156 (N_1156,N_417,N_553);
and U1157 (N_1157,N_702,N_497);
and U1158 (N_1158,N_41,N_510);
and U1159 (N_1159,N_719,N_728);
and U1160 (N_1160,N_290,N_369);
or U1161 (N_1161,N_661,N_334);
and U1162 (N_1162,N_677,N_745);
or U1163 (N_1163,N_570,N_356);
nand U1164 (N_1164,N_599,N_505);
nand U1165 (N_1165,N_488,N_680);
and U1166 (N_1166,N_439,N_710);
or U1167 (N_1167,N_201,N_720);
or U1168 (N_1168,N_561,N_322);
and U1169 (N_1169,N_428,N_497);
nand U1170 (N_1170,N_426,N_178);
nand U1171 (N_1171,N_214,N_61);
or U1172 (N_1172,N_550,N_716);
and U1173 (N_1173,N_15,N_11);
nand U1174 (N_1174,N_297,N_439);
nand U1175 (N_1175,N_383,N_651);
nand U1176 (N_1176,N_79,N_250);
nand U1177 (N_1177,N_130,N_186);
or U1178 (N_1178,N_395,N_718);
nand U1179 (N_1179,N_232,N_692);
nor U1180 (N_1180,N_55,N_477);
nor U1181 (N_1181,N_657,N_38);
nand U1182 (N_1182,N_409,N_468);
or U1183 (N_1183,N_397,N_534);
or U1184 (N_1184,N_479,N_585);
or U1185 (N_1185,N_448,N_292);
nor U1186 (N_1186,N_23,N_167);
nor U1187 (N_1187,N_403,N_408);
nand U1188 (N_1188,N_465,N_334);
nor U1189 (N_1189,N_341,N_56);
and U1190 (N_1190,N_720,N_645);
nor U1191 (N_1191,N_664,N_162);
and U1192 (N_1192,N_378,N_496);
and U1193 (N_1193,N_276,N_337);
nand U1194 (N_1194,N_546,N_190);
nor U1195 (N_1195,N_505,N_708);
nand U1196 (N_1196,N_742,N_47);
nor U1197 (N_1197,N_245,N_433);
nand U1198 (N_1198,N_315,N_433);
nor U1199 (N_1199,N_336,N_622);
nor U1200 (N_1200,N_436,N_665);
or U1201 (N_1201,N_671,N_206);
nand U1202 (N_1202,N_80,N_135);
and U1203 (N_1203,N_239,N_291);
nand U1204 (N_1204,N_265,N_673);
or U1205 (N_1205,N_417,N_1);
or U1206 (N_1206,N_314,N_579);
nor U1207 (N_1207,N_687,N_680);
nor U1208 (N_1208,N_653,N_157);
and U1209 (N_1209,N_533,N_178);
and U1210 (N_1210,N_554,N_630);
nor U1211 (N_1211,N_334,N_464);
nand U1212 (N_1212,N_519,N_361);
or U1213 (N_1213,N_534,N_212);
nor U1214 (N_1214,N_470,N_259);
nor U1215 (N_1215,N_411,N_253);
nand U1216 (N_1216,N_243,N_203);
and U1217 (N_1217,N_245,N_165);
and U1218 (N_1218,N_586,N_407);
xor U1219 (N_1219,N_58,N_720);
and U1220 (N_1220,N_555,N_21);
nand U1221 (N_1221,N_541,N_575);
nand U1222 (N_1222,N_200,N_474);
nor U1223 (N_1223,N_707,N_543);
nor U1224 (N_1224,N_122,N_108);
nor U1225 (N_1225,N_490,N_728);
or U1226 (N_1226,N_172,N_66);
nand U1227 (N_1227,N_344,N_346);
nor U1228 (N_1228,N_267,N_626);
nand U1229 (N_1229,N_481,N_631);
nor U1230 (N_1230,N_572,N_595);
or U1231 (N_1231,N_143,N_188);
and U1232 (N_1232,N_659,N_192);
nor U1233 (N_1233,N_18,N_185);
or U1234 (N_1234,N_283,N_296);
nand U1235 (N_1235,N_262,N_228);
or U1236 (N_1236,N_409,N_488);
nand U1237 (N_1237,N_15,N_385);
or U1238 (N_1238,N_159,N_555);
nor U1239 (N_1239,N_144,N_666);
or U1240 (N_1240,N_399,N_656);
and U1241 (N_1241,N_585,N_146);
and U1242 (N_1242,N_661,N_275);
nand U1243 (N_1243,N_627,N_163);
or U1244 (N_1244,N_146,N_351);
nor U1245 (N_1245,N_405,N_197);
nor U1246 (N_1246,N_88,N_491);
and U1247 (N_1247,N_613,N_673);
nor U1248 (N_1248,N_282,N_337);
or U1249 (N_1249,N_667,N_663);
and U1250 (N_1250,N_215,N_144);
and U1251 (N_1251,N_507,N_251);
and U1252 (N_1252,N_262,N_496);
xor U1253 (N_1253,N_39,N_138);
nor U1254 (N_1254,N_513,N_730);
or U1255 (N_1255,N_321,N_364);
xnor U1256 (N_1256,N_608,N_71);
and U1257 (N_1257,N_102,N_517);
or U1258 (N_1258,N_411,N_479);
nand U1259 (N_1259,N_237,N_323);
nand U1260 (N_1260,N_452,N_118);
nor U1261 (N_1261,N_599,N_597);
or U1262 (N_1262,N_169,N_88);
nor U1263 (N_1263,N_101,N_520);
nor U1264 (N_1264,N_336,N_473);
or U1265 (N_1265,N_544,N_520);
and U1266 (N_1266,N_580,N_78);
or U1267 (N_1267,N_380,N_137);
or U1268 (N_1268,N_177,N_33);
and U1269 (N_1269,N_532,N_5);
and U1270 (N_1270,N_621,N_457);
nand U1271 (N_1271,N_47,N_566);
or U1272 (N_1272,N_415,N_201);
and U1273 (N_1273,N_353,N_595);
and U1274 (N_1274,N_328,N_386);
nor U1275 (N_1275,N_516,N_50);
nand U1276 (N_1276,N_559,N_256);
or U1277 (N_1277,N_574,N_280);
and U1278 (N_1278,N_496,N_610);
nor U1279 (N_1279,N_153,N_207);
or U1280 (N_1280,N_329,N_43);
nor U1281 (N_1281,N_54,N_614);
nand U1282 (N_1282,N_409,N_107);
and U1283 (N_1283,N_166,N_306);
nand U1284 (N_1284,N_162,N_259);
nor U1285 (N_1285,N_189,N_368);
nand U1286 (N_1286,N_484,N_240);
and U1287 (N_1287,N_216,N_608);
nor U1288 (N_1288,N_504,N_447);
xor U1289 (N_1289,N_99,N_670);
nand U1290 (N_1290,N_175,N_372);
and U1291 (N_1291,N_626,N_417);
or U1292 (N_1292,N_159,N_145);
and U1293 (N_1293,N_547,N_478);
xor U1294 (N_1294,N_240,N_424);
or U1295 (N_1295,N_693,N_649);
or U1296 (N_1296,N_723,N_360);
or U1297 (N_1297,N_456,N_40);
and U1298 (N_1298,N_706,N_156);
and U1299 (N_1299,N_5,N_738);
nand U1300 (N_1300,N_74,N_345);
and U1301 (N_1301,N_177,N_686);
nand U1302 (N_1302,N_336,N_94);
nand U1303 (N_1303,N_548,N_242);
nor U1304 (N_1304,N_666,N_606);
or U1305 (N_1305,N_145,N_746);
nor U1306 (N_1306,N_89,N_338);
nor U1307 (N_1307,N_59,N_676);
and U1308 (N_1308,N_377,N_743);
and U1309 (N_1309,N_160,N_374);
and U1310 (N_1310,N_182,N_170);
and U1311 (N_1311,N_655,N_55);
nand U1312 (N_1312,N_148,N_258);
or U1313 (N_1313,N_145,N_23);
xnor U1314 (N_1314,N_148,N_618);
or U1315 (N_1315,N_636,N_254);
and U1316 (N_1316,N_136,N_401);
and U1317 (N_1317,N_738,N_52);
or U1318 (N_1318,N_313,N_540);
nor U1319 (N_1319,N_485,N_16);
or U1320 (N_1320,N_372,N_418);
or U1321 (N_1321,N_134,N_47);
nand U1322 (N_1322,N_592,N_654);
nand U1323 (N_1323,N_580,N_73);
nand U1324 (N_1324,N_683,N_136);
and U1325 (N_1325,N_10,N_710);
nand U1326 (N_1326,N_397,N_86);
nand U1327 (N_1327,N_174,N_109);
and U1328 (N_1328,N_370,N_101);
and U1329 (N_1329,N_390,N_47);
nand U1330 (N_1330,N_519,N_442);
nand U1331 (N_1331,N_127,N_281);
or U1332 (N_1332,N_629,N_82);
nor U1333 (N_1333,N_589,N_567);
nor U1334 (N_1334,N_321,N_224);
or U1335 (N_1335,N_697,N_80);
nand U1336 (N_1336,N_438,N_65);
or U1337 (N_1337,N_81,N_270);
or U1338 (N_1338,N_378,N_603);
nand U1339 (N_1339,N_44,N_75);
nor U1340 (N_1340,N_72,N_682);
and U1341 (N_1341,N_481,N_413);
nand U1342 (N_1342,N_368,N_267);
and U1343 (N_1343,N_149,N_329);
nand U1344 (N_1344,N_535,N_232);
nand U1345 (N_1345,N_252,N_318);
or U1346 (N_1346,N_740,N_419);
nand U1347 (N_1347,N_592,N_438);
or U1348 (N_1348,N_390,N_587);
nand U1349 (N_1349,N_176,N_562);
or U1350 (N_1350,N_290,N_35);
and U1351 (N_1351,N_707,N_708);
xnor U1352 (N_1352,N_485,N_144);
and U1353 (N_1353,N_7,N_9);
or U1354 (N_1354,N_153,N_171);
nor U1355 (N_1355,N_35,N_569);
or U1356 (N_1356,N_724,N_46);
nand U1357 (N_1357,N_701,N_413);
xor U1358 (N_1358,N_154,N_646);
and U1359 (N_1359,N_228,N_687);
nor U1360 (N_1360,N_300,N_119);
xor U1361 (N_1361,N_625,N_425);
nor U1362 (N_1362,N_396,N_424);
and U1363 (N_1363,N_157,N_17);
or U1364 (N_1364,N_141,N_499);
and U1365 (N_1365,N_748,N_87);
or U1366 (N_1366,N_395,N_508);
nand U1367 (N_1367,N_411,N_337);
and U1368 (N_1368,N_32,N_541);
nand U1369 (N_1369,N_409,N_718);
and U1370 (N_1370,N_110,N_104);
and U1371 (N_1371,N_170,N_318);
nand U1372 (N_1372,N_39,N_111);
nand U1373 (N_1373,N_320,N_95);
nand U1374 (N_1374,N_196,N_154);
nor U1375 (N_1375,N_376,N_592);
or U1376 (N_1376,N_540,N_282);
nand U1377 (N_1377,N_29,N_105);
or U1378 (N_1378,N_33,N_532);
and U1379 (N_1379,N_471,N_250);
nand U1380 (N_1380,N_298,N_8);
nand U1381 (N_1381,N_577,N_723);
nand U1382 (N_1382,N_396,N_216);
nand U1383 (N_1383,N_724,N_643);
nand U1384 (N_1384,N_426,N_13);
nor U1385 (N_1385,N_460,N_643);
nor U1386 (N_1386,N_675,N_531);
nor U1387 (N_1387,N_365,N_587);
and U1388 (N_1388,N_294,N_363);
xnor U1389 (N_1389,N_20,N_598);
and U1390 (N_1390,N_336,N_7);
or U1391 (N_1391,N_226,N_508);
nand U1392 (N_1392,N_267,N_372);
nand U1393 (N_1393,N_214,N_596);
nor U1394 (N_1394,N_715,N_279);
nand U1395 (N_1395,N_695,N_439);
and U1396 (N_1396,N_685,N_340);
nand U1397 (N_1397,N_426,N_553);
nand U1398 (N_1398,N_115,N_240);
nand U1399 (N_1399,N_355,N_648);
or U1400 (N_1400,N_37,N_66);
nor U1401 (N_1401,N_639,N_563);
nand U1402 (N_1402,N_204,N_549);
and U1403 (N_1403,N_690,N_481);
nand U1404 (N_1404,N_28,N_687);
and U1405 (N_1405,N_283,N_37);
nor U1406 (N_1406,N_655,N_342);
nor U1407 (N_1407,N_333,N_210);
nor U1408 (N_1408,N_665,N_350);
nand U1409 (N_1409,N_276,N_538);
and U1410 (N_1410,N_252,N_312);
or U1411 (N_1411,N_2,N_549);
and U1412 (N_1412,N_256,N_306);
or U1413 (N_1413,N_106,N_358);
nand U1414 (N_1414,N_680,N_425);
nand U1415 (N_1415,N_10,N_580);
and U1416 (N_1416,N_459,N_702);
xnor U1417 (N_1417,N_148,N_584);
nor U1418 (N_1418,N_343,N_684);
nor U1419 (N_1419,N_719,N_668);
and U1420 (N_1420,N_111,N_470);
and U1421 (N_1421,N_131,N_237);
xor U1422 (N_1422,N_11,N_566);
nand U1423 (N_1423,N_237,N_61);
nor U1424 (N_1424,N_603,N_712);
or U1425 (N_1425,N_163,N_495);
or U1426 (N_1426,N_175,N_470);
and U1427 (N_1427,N_665,N_41);
nand U1428 (N_1428,N_253,N_179);
nand U1429 (N_1429,N_608,N_433);
and U1430 (N_1430,N_81,N_623);
or U1431 (N_1431,N_381,N_52);
and U1432 (N_1432,N_319,N_518);
nand U1433 (N_1433,N_380,N_13);
nor U1434 (N_1434,N_145,N_8);
nor U1435 (N_1435,N_27,N_205);
and U1436 (N_1436,N_704,N_225);
and U1437 (N_1437,N_177,N_552);
and U1438 (N_1438,N_241,N_244);
xor U1439 (N_1439,N_86,N_596);
nor U1440 (N_1440,N_321,N_260);
or U1441 (N_1441,N_114,N_68);
nand U1442 (N_1442,N_628,N_215);
nand U1443 (N_1443,N_732,N_553);
and U1444 (N_1444,N_219,N_213);
and U1445 (N_1445,N_48,N_383);
nor U1446 (N_1446,N_452,N_287);
nand U1447 (N_1447,N_554,N_93);
nor U1448 (N_1448,N_425,N_191);
nor U1449 (N_1449,N_572,N_277);
and U1450 (N_1450,N_647,N_590);
and U1451 (N_1451,N_285,N_521);
nor U1452 (N_1452,N_275,N_463);
nand U1453 (N_1453,N_571,N_643);
nand U1454 (N_1454,N_361,N_676);
and U1455 (N_1455,N_495,N_363);
or U1456 (N_1456,N_19,N_125);
and U1457 (N_1457,N_167,N_436);
nand U1458 (N_1458,N_283,N_309);
nor U1459 (N_1459,N_222,N_127);
nor U1460 (N_1460,N_237,N_196);
nor U1461 (N_1461,N_376,N_271);
nand U1462 (N_1462,N_531,N_629);
or U1463 (N_1463,N_155,N_3);
nor U1464 (N_1464,N_591,N_37);
nor U1465 (N_1465,N_363,N_455);
nand U1466 (N_1466,N_187,N_155);
or U1467 (N_1467,N_109,N_620);
nand U1468 (N_1468,N_580,N_65);
nand U1469 (N_1469,N_698,N_205);
nand U1470 (N_1470,N_1,N_707);
nor U1471 (N_1471,N_100,N_210);
nor U1472 (N_1472,N_613,N_181);
nor U1473 (N_1473,N_689,N_360);
or U1474 (N_1474,N_210,N_721);
nor U1475 (N_1475,N_331,N_61);
or U1476 (N_1476,N_546,N_225);
nand U1477 (N_1477,N_572,N_579);
xnor U1478 (N_1478,N_530,N_386);
or U1479 (N_1479,N_495,N_507);
nand U1480 (N_1480,N_626,N_173);
and U1481 (N_1481,N_507,N_65);
nor U1482 (N_1482,N_566,N_295);
nand U1483 (N_1483,N_99,N_209);
nor U1484 (N_1484,N_131,N_326);
nand U1485 (N_1485,N_479,N_684);
and U1486 (N_1486,N_393,N_301);
nor U1487 (N_1487,N_616,N_404);
nor U1488 (N_1488,N_261,N_464);
nand U1489 (N_1489,N_130,N_142);
or U1490 (N_1490,N_379,N_609);
and U1491 (N_1491,N_679,N_560);
nand U1492 (N_1492,N_579,N_68);
and U1493 (N_1493,N_737,N_139);
or U1494 (N_1494,N_719,N_154);
nand U1495 (N_1495,N_470,N_641);
nor U1496 (N_1496,N_572,N_121);
nor U1497 (N_1497,N_419,N_521);
or U1498 (N_1498,N_47,N_719);
nand U1499 (N_1499,N_480,N_341);
nand U1500 (N_1500,N_1477,N_943);
and U1501 (N_1501,N_1397,N_1199);
nand U1502 (N_1502,N_1354,N_845);
nand U1503 (N_1503,N_1083,N_844);
nand U1504 (N_1504,N_981,N_936);
nor U1505 (N_1505,N_1220,N_1028);
and U1506 (N_1506,N_1060,N_887);
and U1507 (N_1507,N_1058,N_1104);
or U1508 (N_1508,N_850,N_1044);
and U1509 (N_1509,N_1273,N_1209);
and U1510 (N_1510,N_1183,N_1421);
nand U1511 (N_1511,N_982,N_1266);
nor U1512 (N_1512,N_1188,N_757);
nor U1513 (N_1513,N_1186,N_1111);
and U1514 (N_1514,N_1461,N_1314);
nand U1515 (N_1515,N_860,N_1371);
nor U1516 (N_1516,N_1007,N_1338);
or U1517 (N_1517,N_1494,N_1377);
or U1518 (N_1518,N_1307,N_1232);
xnor U1519 (N_1519,N_1452,N_996);
nand U1520 (N_1520,N_900,N_1243);
or U1521 (N_1521,N_1348,N_920);
nand U1522 (N_1522,N_1327,N_788);
nor U1523 (N_1523,N_1445,N_1300);
and U1524 (N_1524,N_944,N_1481);
and U1525 (N_1525,N_924,N_762);
xor U1526 (N_1526,N_1207,N_1095);
xnor U1527 (N_1527,N_1178,N_1374);
or U1528 (N_1528,N_1379,N_1469);
or U1529 (N_1529,N_1238,N_1059);
nand U1530 (N_1530,N_822,N_1254);
nor U1531 (N_1531,N_902,N_1294);
or U1532 (N_1532,N_1335,N_1261);
nand U1533 (N_1533,N_1484,N_817);
nor U1534 (N_1534,N_997,N_759);
nor U1535 (N_1535,N_1226,N_1437);
and U1536 (N_1536,N_1200,N_1019);
or U1537 (N_1537,N_938,N_1233);
nor U1538 (N_1538,N_1342,N_808);
or U1539 (N_1539,N_935,N_1302);
nand U1540 (N_1540,N_1078,N_842);
and U1541 (N_1541,N_1463,N_1029);
xor U1542 (N_1542,N_959,N_960);
nand U1543 (N_1543,N_1466,N_1244);
nand U1544 (N_1544,N_1011,N_945);
or U1545 (N_1545,N_1073,N_1352);
or U1546 (N_1546,N_921,N_1239);
nor U1547 (N_1547,N_1031,N_1187);
nor U1548 (N_1548,N_1350,N_915);
nor U1549 (N_1549,N_1416,N_1107);
and U1550 (N_1550,N_1127,N_859);
and U1551 (N_1551,N_1419,N_894);
and U1552 (N_1552,N_1456,N_917);
and U1553 (N_1553,N_1412,N_846);
and U1554 (N_1554,N_1137,N_988);
and U1555 (N_1555,N_892,N_952);
nand U1556 (N_1556,N_1242,N_1424);
or U1557 (N_1557,N_1153,N_931);
and U1558 (N_1558,N_1084,N_1470);
and U1559 (N_1559,N_1049,N_918);
or U1560 (N_1560,N_1158,N_965);
nor U1561 (N_1561,N_1110,N_1376);
nand U1562 (N_1562,N_1334,N_893);
nor U1563 (N_1563,N_1215,N_912);
nor U1564 (N_1564,N_911,N_840);
nor U1565 (N_1565,N_1010,N_870);
or U1566 (N_1566,N_1042,N_1490);
and U1567 (N_1567,N_1034,N_1388);
nor U1568 (N_1568,N_1288,N_1202);
and U1569 (N_1569,N_1148,N_919);
or U1570 (N_1570,N_1402,N_1473);
and U1571 (N_1571,N_1015,N_1305);
nand U1572 (N_1572,N_841,N_1165);
nor U1573 (N_1573,N_1140,N_1144);
or U1574 (N_1574,N_856,N_929);
and U1575 (N_1575,N_1365,N_1033);
nor U1576 (N_1576,N_897,N_1077);
nor U1577 (N_1577,N_1050,N_1289);
or U1578 (N_1578,N_1337,N_1280);
or U1579 (N_1579,N_1359,N_1432);
nor U1580 (N_1580,N_883,N_1032);
nand U1581 (N_1581,N_833,N_1353);
or U1582 (N_1582,N_1414,N_984);
nor U1583 (N_1583,N_828,N_1169);
xor U1584 (N_1584,N_990,N_1035);
nand U1585 (N_1585,N_778,N_1223);
nor U1586 (N_1586,N_1038,N_946);
nand U1587 (N_1587,N_916,N_882);
nand U1588 (N_1588,N_1324,N_1047);
nor U1589 (N_1589,N_1429,N_1260);
nor U1590 (N_1590,N_980,N_1317);
or U1591 (N_1591,N_1340,N_1142);
nand U1592 (N_1592,N_1384,N_884);
and U1593 (N_1593,N_1003,N_1192);
nand U1594 (N_1594,N_881,N_1442);
and U1595 (N_1595,N_1120,N_1381);
nor U1596 (N_1596,N_750,N_906);
nor U1597 (N_1597,N_761,N_1193);
nand U1598 (N_1598,N_1292,N_871);
or U1599 (N_1599,N_1116,N_1052);
nand U1600 (N_1600,N_1449,N_1264);
and U1601 (N_1601,N_1085,N_1231);
and U1602 (N_1602,N_826,N_1299);
or U1603 (N_1603,N_1057,N_1407);
or U1604 (N_1604,N_1395,N_971);
or U1605 (N_1605,N_1166,N_1177);
and U1606 (N_1606,N_1203,N_795);
nor U1607 (N_1607,N_797,N_1304);
or U1608 (N_1608,N_1272,N_1139);
or U1609 (N_1609,N_1039,N_1357);
nand U1610 (N_1610,N_1228,N_1287);
and U1611 (N_1611,N_1064,N_798);
nand U1612 (N_1612,N_1176,N_1291);
nor U1613 (N_1613,N_1447,N_1441);
nand U1614 (N_1614,N_1126,N_1321);
nand U1615 (N_1615,N_839,N_809);
nor U1616 (N_1616,N_1418,N_1063);
or U1617 (N_1617,N_1322,N_854);
and U1618 (N_1618,N_1113,N_1005);
nor U1619 (N_1619,N_983,N_930);
nor U1620 (N_1620,N_1267,N_876);
nor U1621 (N_1621,N_1195,N_967);
nor U1622 (N_1622,N_868,N_825);
nand U1623 (N_1623,N_1062,N_1446);
nor U1624 (N_1624,N_977,N_1086);
nand U1625 (N_1625,N_942,N_1318);
and U1626 (N_1626,N_1349,N_1436);
nor U1627 (N_1627,N_888,N_1329);
and U1628 (N_1628,N_1043,N_1392);
nor U1629 (N_1629,N_1333,N_858);
and U1630 (N_1630,N_1236,N_1013);
or U1631 (N_1631,N_1184,N_1132);
nand U1632 (N_1632,N_1309,N_1467);
nor U1633 (N_1633,N_775,N_1450);
or U1634 (N_1634,N_1323,N_951);
and U1635 (N_1635,N_979,N_923);
nand U1636 (N_1636,N_1022,N_785);
and U1637 (N_1637,N_832,N_843);
or U1638 (N_1638,N_956,N_1235);
nor U1639 (N_1639,N_1451,N_1296);
xnor U1640 (N_1640,N_1024,N_1089);
or U1641 (N_1641,N_861,N_1016);
or U1642 (N_1642,N_973,N_1030);
nor U1643 (N_1643,N_818,N_1247);
nand U1644 (N_1644,N_899,N_986);
or U1645 (N_1645,N_1312,N_925);
nand U1646 (N_1646,N_816,N_1240);
and U1647 (N_1647,N_820,N_1316);
nand U1648 (N_1648,N_901,N_807);
nand U1649 (N_1649,N_1012,N_891);
and U1650 (N_1650,N_1366,N_954);
and U1651 (N_1651,N_1079,N_756);
and U1652 (N_1652,N_1141,N_1155);
nand U1653 (N_1653,N_1097,N_987);
nor U1654 (N_1654,N_1347,N_1303);
and U1655 (N_1655,N_1399,N_1105);
nand U1656 (N_1656,N_970,N_802);
or U1657 (N_1657,N_1219,N_1046);
and U1658 (N_1658,N_1315,N_1311);
nand U1659 (N_1659,N_964,N_1018);
and U1660 (N_1660,N_1131,N_1439);
nand U1661 (N_1661,N_1464,N_1382);
nor U1662 (N_1662,N_1213,N_769);
or U1663 (N_1663,N_1364,N_1306);
or U1664 (N_1664,N_1114,N_1076);
or U1665 (N_1665,N_875,N_771);
nand U1666 (N_1666,N_1409,N_1023);
nor U1667 (N_1667,N_1325,N_799);
or U1668 (N_1668,N_1008,N_1036);
nor U1669 (N_1669,N_1051,N_1135);
and U1670 (N_1670,N_910,N_1408);
nor U1671 (N_1671,N_1396,N_1265);
xor U1672 (N_1672,N_1027,N_1269);
and U1673 (N_1673,N_992,N_1164);
nand U1674 (N_1674,N_1246,N_1168);
and U1675 (N_1675,N_805,N_1401);
xor U1676 (N_1676,N_1259,N_1026);
or U1677 (N_1677,N_1128,N_1162);
and U1678 (N_1678,N_1257,N_889);
nor U1679 (N_1679,N_1152,N_914);
or U1680 (N_1680,N_1160,N_847);
or U1681 (N_1681,N_1041,N_790);
or U1682 (N_1682,N_776,N_1276);
nand U1683 (N_1683,N_1092,N_1413);
nor U1684 (N_1684,N_1072,N_1156);
and U1685 (N_1685,N_779,N_877);
nor U1686 (N_1686,N_1014,N_1275);
or U1687 (N_1687,N_1198,N_993);
and U1688 (N_1688,N_1251,N_1387);
and U1689 (N_1689,N_1189,N_1448);
xnor U1690 (N_1690,N_1194,N_878);
nor U1691 (N_1691,N_1081,N_1345);
nand U1692 (N_1692,N_1459,N_1151);
or U1693 (N_1693,N_772,N_950);
nor U1694 (N_1694,N_1403,N_994);
or U1695 (N_1695,N_789,N_1492);
nand U1696 (N_1696,N_1150,N_1344);
or U1697 (N_1697,N_1225,N_1270);
and U1698 (N_1698,N_1000,N_1175);
and U1699 (N_1699,N_1295,N_1098);
nand U1700 (N_1700,N_1230,N_1358);
and U1701 (N_1701,N_1117,N_1196);
and U1702 (N_1702,N_1025,N_1145);
or U1703 (N_1703,N_1278,N_922);
xor U1704 (N_1704,N_1282,N_1201);
and U1705 (N_1705,N_1115,N_1108);
or U1706 (N_1706,N_1373,N_1319);
nor U1707 (N_1707,N_815,N_1159);
xnor U1708 (N_1708,N_1332,N_1250);
nor U1709 (N_1709,N_796,N_794);
and U1710 (N_1710,N_1048,N_1245);
xnor U1711 (N_1711,N_1205,N_1167);
and U1712 (N_1712,N_1367,N_1037);
nor U1713 (N_1713,N_764,N_784);
nand U1714 (N_1714,N_1283,N_811);
nand U1715 (N_1715,N_1091,N_1458);
and U1716 (N_1716,N_1453,N_1454);
or U1717 (N_1717,N_985,N_958);
nor U1718 (N_1718,N_1431,N_1362);
or U1719 (N_1719,N_1191,N_1391);
nand U1720 (N_1720,N_1101,N_885);
and U1721 (N_1721,N_1020,N_904);
or U1722 (N_1722,N_913,N_969);
or U1723 (N_1723,N_1056,N_1130);
nor U1724 (N_1724,N_1301,N_926);
or U1725 (N_1725,N_873,N_1475);
nand U1726 (N_1726,N_1489,N_1171);
or U1727 (N_1727,N_1248,N_1222);
or U1728 (N_1728,N_1383,N_853);
and U1729 (N_1729,N_1087,N_1129);
or U1730 (N_1730,N_1380,N_780);
nor U1731 (N_1731,N_932,N_1368);
and U1732 (N_1732,N_783,N_961);
nand U1733 (N_1733,N_940,N_896);
nand U1734 (N_1734,N_1370,N_1218);
nand U1735 (N_1735,N_1069,N_1093);
nor U1736 (N_1736,N_862,N_1341);
nand U1737 (N_1737,N_1482,N_962);
and U1738 (N_1738,N_1343,N_1146);
nand U1739 (N_1739,N_1161,N_1217);
and U1740 (N_1740,N_806,N_903);
or U1741 (N_1741,N_879,N_869);
or U1742 (N_1742,N_1263,N_1181);
nand U1743 (N_1743,N_1001,N_1468);
and U1744 (N_1744,N_927,N_1009);
nor U1745 (N_1745,N_948,N_1285);
or U1746 (N_1746,N_1149,N_767);
and U1747 (N_1747,N_1179,N_1355);
or U1748 (N_1748,N_1124,N_1277);
nor U1749 (N_1749,N_836,N_1206);
or U1750 (N_1750,N_1075,N_1389);
or U1751 (N_1751,N_1157,N_1224);
nor U1752 (N_1752,N_1320,N_937);
xor U1753 (N_1753,N_1420,N_753);
nor U1754 (N_1754,N_1053,N_1180);
or U1755 (N_1755,N_786,N_1002);
nand U1756 (N_1756,N_1241,N_834);
or U1757 (N_1757,N_1268,N_804);
and U1758 (N_1758,N_1212,N_752);
nor U1759 (N_1759,N_1284,N_768);
nand U1760 (N_1760,N_895,N_1074);
and U1761 (N_1761,N_1274,N_1360);
nand U1762 (N_1762,N_1109,N_907);
and U1763 (N_1763,N_1483,N_765);
and U1764 (N_1764,N_1021,N_1182);
nor U1765 (N_1765,N_1185,N_1112);
nor U1766 (N_1766,N_1351,N_823);
nor U1767 (N_1767,N_1369,N_909);
or U1768 (N_1768,N_770,N_1485);
nor U1769 (N_1769,N_1390,N_1253);
nor U1770 (N_1770,N_872,N_934);
or U1771 (N_1771,N_1204,N_1136);
nand U1772 (N_1772,N_898,N_1460);
or U1773 (N_1773,N_972,N_821);
and U1774 (N_1774,N_995,N_947);
nor U1775 (N_1775,N_1099,N_1040);
nor U1776 (N_1776,N_1491,N_1465);
nor U1777 (N_1777,N_1308,N_1427);
nand U1778 (N_1778,N_1423,N_999);
or U1779 (N_1779,N_851,N_1444);
or U1780 (N_1780,N_1339,N_819);
and U1781 (N_1781,N_774,N_1174);
nand U1782 (N_1782,N_813,N_1071);
nand U1783 (N_1783,N_976,N_1495);
nor U1784 (N_1784,N_1102,N_1415);
and U1785 (N_1785,N_791,N_755);
nor U1786 (N_1786,N_827,N_837);
nand U1787 (N_1787,N_1411,N_1080);
nor U1788 (N_1788,N_1331,N_1106);
or U1789 (N_1789,N_1255,N_1123);
nand U1790 (N_1790,N_880,N_1271);
and U1791 (N_1791,N_1045,N_830);
nor U1792 (N_1792,N_1375,N_1118);
or U1793 (N_1793,N_803,N_1173);
or U1794 (N_1794,N_1190,N_1147);
nand U1795 (N_1795,N_1434,N_1090);
nor U1796 (N_1796,N_852,N_933);
nand U1797 (N_1797,N_1455,N_1088);
nor U1798 (N_1798,N_1234,N_835);
or U1799 (N_1799,N_1346,N_1386);
or U1800 (N_1800,N_787,N_1290);
nor U1801 (N_1801,N_792,N_978);
and U1802 (N_1802,N_855,N_864);
nor U1803 (N_1803,N_1258,N_1480);
nand U1804 (N_1804,N_1474,N_1252);
nand U1805 (N_1805,N_829,N_1493);
or U1806 (N_1806,N_1404,N_1067);
or U1807 (N_1807,N_1262,N_1486);
nand U1808 (N_1808,N_953,N_966);
nand U1809 (N_1809,N_1214,N_831);
nand U1810 (N_1810,N_1361,N_782);
nand U1811 (N_1811,N_1385,N_1488);
nor U1812 (N_1812,N_857,N_1497);
or U1813 (N_1813,N_863,N_1430);
and U1814 (N_1814,N_1279,N_1216);
or U1815 (N_1815,N_865,N_975);
nor U1816 (N_1816,N_1082,N_848);
and U1817 (N_1817,N_866,N_1208);
and U1818 (N_1818,N_1061,N_1433);
and U1819 (N_1819,N_838,N_949);
nor U1820 (N_1820,N_1096,N_1103);
and U1821 (N_1821,N_1457,N_1006);
or U1822 (N_1822,N_766,N_908);
nor U1823 (N_1823,N_1440,N_1065);
nand U1824 (N_1824,N_1487,N_801);
nand U1825 (N_1825,N_1336,N_1197);
xor U1826 (N_1826,N_989,N_1425);
and U1827 (N_1827,N_941,N_955);
and U1828 (N_1828,N_1400,N_974);
nand U1829 (N_1829,N_1394,N_1133);
nand U1830 (N_1830,N_1298,N_1054);
xor U1831 (N_1831,N_957,N_1293);
nand U1832 (N_1832,N_1055,N_1356);
nor U1833 (N_1833,N_1328,N_1017);
and U1834 (N_1834,N_939,N_1313);
nand U1835 (N_1835,N_1066,N_1472);
or U1836 (N_1836,N_773,N_814);
and U1837 (N_1837,N_1172,N_1438);
or U1838 (N_1838,N_1121,N_1211);
nand U1839 (N_1839,N_1256,N_1068);
and U1840 (N_1840,N_1372,N_751);
nor U1841 (N_1841,N_800,N_1143);
nor U1842 (N_1842,N_1227,N_777);
xnor U1843 (N_1843,N_1094,N_1237);
or U1844 (N_1844,N_1393,N_1443);
nor U1845 (N_1845,N_1499,N_810);
and U1846 (N_1846,N_1479,N_1435);
nor U1847 (N_1847,N_1221,N_1100);
nor U1848 (N_1848,N_998,N_1422);
or U1849 (N_1849,N_754,N_1426);
or U1850 (N_1850,N_1119,N_1210);
nor U1851 (N_1851,N_1163,N_890);
nand U1852 (N_1852,N_991,N_1428);
nand U1853 (N_1853,N_963,N_1310);
nand U1854 (N_1854,N_1297,N_1471);
nor U1855 (N_1855,N_1281,N_1417);
nand U1856 (N_1856,N_886,N_824);
and U1857 (N_1857,N_1122,N_874);
nand U1858 (N_1858,N_812,N_1406);
nand U1859 (N_1859,N_1398,N_1134);
nor U1860 (N_1860,N_1170,N_1154);
or U1861 (N_1861,N_1378,N_1286);
or U1862 (N_1862,N_968,N_1125);
nor U1863 (N_1863,N_928,N_905);
nand U1864 (N_1864,N_1138,N_1326);
and U1865 (N_1865,N_760,N_1229);
nor U1866 (N_1866,N_758,N_867);
and U1867 (N_1867,N_1410,N_781);
or U1868 (N_1868,N_1330,N_1476);
or U1869 (N_1869,N_1004,N_1498);
nor U1870 (N_1870,N_1462,N_1478);
or U1871 (N_1871,N_1496,N_1405);
nor U1872 (N_1872,N_763,N_849);
nand U1873 (N_1873,N_793,N_1249);
nand U1874 (N_1874,N_1363,N_1070);
or U1875 (N_1875,N_823,N_784);
or U1876 (N_1876,N_964,N_1492);
and U1877 (N_1877,N_971,N_1486);
and U1878 (N_1878,N_1225,N_1035);
or U1879 (N_1879,N_1308,N_968);
nor U1880 (N_1880,N_1431,N_1283);
nor U1881 (N_1881,N_825,N_757);
and U1882 (N_1882,N_1165,N_1328);
nor U1883 (N_1883,N_847,N_1161);
nand U1884 (N_1884,N_804,N_882);
and U1885 (N_1885,N_1011,N_1163);
or U1886 (N_1886,N_1131,N_795);
xor U1887 (N_1887,N_1471,N_789);
nand U1888 (N_1888,N_901,N_914);
or U1889 (N_1889,N_1478,N_1159);
nand U1890 (N_1890,N_1084,N_1341);
nor U1891 (N_1891,N_1445,N_1102);
nand U1892 (N_1892,N_1104,N_1015);
and U1893 (N_1893,N_965,N_944);
nor U1894 (N_1894,N_1080,N_1218);
nor U1895 (N_1895,N_1265,N_1020);
nand U1896 (N_1896,N_1382,N_756);
nor U1897 (N_1897,N_1091,N_892);
nor U1898 (N_1898,N_902,N_1069);
and U1899 (N_1899,N_862,N_1471);
or U1900 (N_1900,N_1123,N_1139);
and U1901 (N_1901,N_1460,N_1198);
and U1902 (N_1902,N_1421,N_1404);
and U1903 (N_1903,N_961,N_1219);
nand U1904 (N_1904,N_934,N_1079);
or U1905 (N_1905,N_1026,N_1104);
nand U1906 (N_1906,N_979,N_835);
and U1907 (N_1907,N_1001,N_1214);
nand U1908 (N_1908,N_770,N_1305);
nor U1909 (N_1909,N_957,N_825);
or U1910 (N_1910,N_1047,N_1106);
or U1911 (N_1911,N_1225,N_1255);
and U1912 (N_1912,N_1437,N_1433);
nor U1913 (N_1913,N_1311,N_960);
or U1914 (N_1914,N_940,N_1103);
or U1915 (N_1915,N_1071,N_1166);
nor U1916 (N_1916,N_931,N_1306);
nor U1917 (N_1917,N_786,N_1156);
nor U1918 (N_1918,N_1262,N_1214);
and U1919 (N_1919,N_1426,N_1462);
nand U1920 (N_1920,N_1161,N_1435);
or U1921 (N_1921,N_985,N_827);
or U1922 (N_1922,N_1456,N_924);
nand U1923 (N_1923,N_769,N_1178);
or U1924 (N_1924,N_1368,N_873);
nor U1925 (N_1925,N_877,N_1016);
nor U1926 (N_1926,N_934,N_818);
or U1927 (N_1927,N_956,N_1036);
and U1928 (N_1928,N_1061,N_1004);
nand U1929 (N_1929,N_1050,N_1363);
or U1930 (N_1930,N_1003,N_883);
nor U1931 (N_1931,N_1272,N_1487);
xor U1932 (N_1932,N_880,N_999);
nor U1933 (N_1933,N_914,N_1249);
nor U1934 (N_1934,N_1144,N_1184);
nor U1935 (N_1935,N_879,N_892);
and U1936 (N_1936,N_922,N_1340);
or U1937 (N_1937,N_992,N_1065);
nand U1938 (N_1938,N_937,N_1014);
xnor U1939 (N_1939,N_794,N_1060);
nor U1940 (N_1940,N_866,N_783);
and U1941 (N_1941,N_1356,N_804);
and U1942 (N_1942,N_1476,N_1052);
or U1943 (N_1943,N_1200,N_1493);
xnor U1944 (N_1944,N_1487,N_970);
and U1945 (N_1945,N_1050,N_932);
nand U1946 (N_1946,N_1084,N_1033);
nand U1947 (N_1947,N_1230,N_1200);
and U1948 (N_1948,N_1225,N_1229);
and U1949 (N_1949,N_1299,N_1067);
nor U1950 (N_1950,N_1330,N_1192);
or U1951 (N_1951,N_1029,N_1449);
nand U1952 (N_1952,N_1079,N_1327);
nand U1953 (N_1953,N_976,N_1364);
nand U1954 (N_1954,N_1350,N_1420);
nor U1955 (N_1955,N_1209,N_1067);
and U1956 (N_1956,N_1222,N_1095);
or U1957 (N_1957,N_1164,N_1008);
nand U1958 (N_1958,N_777,N_984);
and U1959 (N_1959,N_794,N_1180);
or U1960 (N_1960,N_1216,N_945);
or U1961 (N_1961,N_1178,N_904);
and U1962 (N_1962,N_1303,N_795);
nor U1963 (N_1963,N_1234,N_1076);
nand U1964 (N_1964,N_1004,N_894);
and U1965 (N_1965,N_1409,N_799);
nor U1966 (N_1966,N_750,N_968);
xor U1967 (N_1967,N_1214,N_1394);
nor U1968 (N_1968,N_1421,N_1417);
or U1969 (N_1969,N_1069,N_909);
or U1970 (N_1970,N_1296,N_1491);
nand U1971 (N_1971,N_1065,N_905);
nor U1972 (N_1972,N_859,N_1304);
and U1973 (N_1973,N_1100,N_1050);
nand U1974 (N_1974,N_1411,N_921);
nand U1975 (N_1975,N_973,N_1077);
xor U1976 (N_1976,N_1074,N_792);
nor U1977 (N_1977,N_968,N_1324);
nor U1978 (N_1978,N_972,N_1259);
or U1979 (N_1979,N_1311,N_1309);
and U1980 (N_1980,N_1057,N_1128);
nor U1981 (N_1981,N_869,N_1466);
or U1982 (N_1982,N_794,N_867);
or U1983 (N_1983,N_1017,N_837);
nand U1984 (N_1984,N_946,N_1077);
nand U1985 (N_1985,N_1013,N_869);
nor U1986 (N_1986,N_951,N_1168);
and U1987 (N_1987,N_1426,N_1329);
and U1988 (N_1988,N_1410,N_1130);
nor U1989 (N_1989,N_1462,N_1402);
or U1990 (N_1990,N_1180,N_1346);
nor U1991 (N_1991,N_1240,N_1423);
and U1992 (N_1992,N_1398,N_995);
nor U1993 (N_1993,N_855,N_1345);
and U1994 (N_1994,N_971,N_1021);
nor U1995 (N_1995,N_1260,N_1402);
and U1996 (N_1996,N_1014,N_1142);
nand U1997 (N_1997,N_965,N_1483);
or U1998 (N_1998,N_1386,N_968);
nor U1999 (N_1999,N_1333,N_1442);
or U2000 (N_2000,N_1423,N_1421);
or U2001 (N_2001,N_900,N_1470);
and U2002 (N_2002,N_1236,N_1119);
or U2003 (N_2003,N_1114,N_1008);
and U2004 (N_2004,N_1299,N_1017);
nor U2005 (N_2005,N_1178,N_1339);
nand U2006 (N_2006,N_1007,N_1436);
nor U2007 (N_2007,N_1182,N_1312);
nand U2008 (N_2008,N_998,N_971);
and U2009 (N_2009,N_900,N_1337);
nand U2010 (N_2010,N_1451,N_1108);
nor U2011 (N_2011,N_1491,N_1356);
and U2012 (N_2012,N_1474,N_1211);
and U2013 (N_2013,N_1167,N_1279);
nand U2014 (N_2014,N_1335,N_1166);
or U2015 (N_2015,N_1340,N_789);
nor U2016 (N_2016,N_902,N_834);
nor U2017 (N_2017,N_1335,N_870);
nand U2018 (N_2018,N_857,N_752);
and U2019 (N_2019,N_860,N_856);
or U2020 (N_2020,N_925,N_1156);
nand U2021 (N_2021,N_1111,N_1032);
or U2022 (N_2022,N_910,N_840);
nand U2023 (N_2023,N_1100,N_958);
nand U2024 (N_2024,N_825,N_1435);
nor U2025 (N_2025,N_836,N_1220);
nor U2026 (N_2026,N_1032,N_1053);
nor U2027 (N_2027,N_1294,N_752);
nand U2028 (N_2028,N_1284,N_1143);
or U2029 (N_2029,N_1163,N_955);
or U2030 (N_2030,N_1003,N_1417);
xor U2031 (N_2031,N_929,N_841);
or U2032 (N_2032,N_924,N_1348);
nor U2033 (N_2033,N_957,N_767);
nor U2034 (N_2034,N_1011,N_875);
and U2035 (N_2035,N_1444,N_907);
and U2036 (N_2036,N_792,N_958);
nor U2037 (N_2037,N_770,N_1184);
nand U2038 (N_2038,N_1421,N_957);
nand U2039 (N_2039,N_884,N_981);
nand U2040 (N_2040,N_824,N_1122);
nor U2041 (N_2041,N_1380,N_1486);
and U2042 (N_2042,N_1029,N_1476);
or U2043 (N_2043,N_1465,N_1116);
or U2044 (N_2044,N_1351,N_1122);
or U2045 (N_2045,N_767,N_769);
nand U2046 (N_2046,N_832,N_1462);
or U2047 (N_2047,N_1053,N_858);
nor U2048 (N_2048,N_1186,N_900);
nand U2049 (N_2049,N_835,N_1204);
nand U2050 (N_2050,N_1280,N_1224);
or U2051 (N_2051,N_999,N_988);
or U2052 (N_2052,N_1380,N_1338);
or U2053 (N_2053,N_1207,N_1254);
and U2054 (N_2054,N_840,N_1342);
and U2055 (N_2055,N_1128,N_1161);
and U2056 (N_2056,N_875,N_1040);
and U2057 (N_2057,N_1124,N_1056);
nor U2058 (N_2058,N_1389,N_780);
nor U2059 (N_2059,N_1125,N_992);
nor U2060 (N_2060,N_900,N_1455);
nor U2061 (N_2061,N_1159,N_761);
nor U2062 (N_2062,N_1284,N_1247);
and U2063 (N_2063,N_1239,N_1039);
xor U2064 (N_2064,N_1116,N_784);
and U2065 (N_2065,N_1437,N_971);
or U2066 (N_2066,N_942,N_1360);
and U2067 (N_2067,N_1126,N_936);
and U2068 (N_2068,N_764,N_940);
nor U2069 (N_2069,N_1318,N_825);
nor U2070 (N_2070,N_1226,N_982);
and U2071 (N_2071,N_984,N_1341);
and U2072 (N_2072,N_1015,N_881);
and U2073 (N_2073,N_778,N_1156);
and U2074 (N_2074,N_1251,N_1097);
nor U2075 (N_2075,N_899,N_963);
nand U2076 (N_2076,N_938,N_1487);
or U2077 (N_2077,N_961,N_1489);
and U2078 (N_2078,N_1016,N_894);
and U2079 (N_2079,N_1322,N_1084);
or U2080 (N_2080,N_1236,N_1345);
or U2081 (N_2081,N_1370,N_1057);
and U2082 (N_2082,N_1184,N_1454);
xnor U2083 (N_2083,N_1325,N_1047);
or U2084 (N_2084,N_1262,N_853);
and U2085 (N_2085,N_1277,N_1396);
nand U2086 (N_2086,N_1497,N_795);
nand U2087 (N_2087,N_1415,N_1140);
nor U2088 (N_2088,N_911,N_1289);
and U2089 (N_2089,N_1050,N_1149);
nor U2090 (N_2090,N_860,N_1423);
or U2091 (N_2091,N_1376,N_1010);
nand U2092 (N_2092,N_1067,N_1126);
nand U2093 (N_2093,N_1105,N_1096);
or U2094 (N_2094,N_1075,N_832);
nand U2095 (N_2095,N_1488,N_1087);
nor U2096 (N_2096,N_931,N_1232);
nand U2097 (N_2097,N_1222,N_1402);
or U2098 (N_2098,N_958,N_1126);
nor U2099 (N_2099,N_1298,N_994);
and U2100 (N_2100,N_1493,N_1126);
and U2101 (N_2101,N_1405,N_1371);
or U2102 (N_2102,N_963,N_1039);
nor U2103 (N_2103,N_1266,N_1028);
nand U2104 (N_2104,N_1013,N_944);
nand U2105 (N_2105,N_1052,N_1482);
and U2106 (N_2106,N_1259,N_833);
and U2107 (N_2107,N_1413,N_1245);
or U2108 (N_2108,N_1215,N_1237);
nor U2109 (N_2109,N_1121,N_1473);
nor U2110 (N_2110,N_904,N_777);
xnor U2111 (N_2111,N_854,N_1378);
or U2112 (N_2112,N_848,N_1282);
and U2113 (N_2113,N_1302,N_1249);
nand U2114 (N_2114,N_1137,N_1475);
and U2115 (N_2115,N_766,N_845);
xor U2116 (N_2116,N_960,N_976);
nand U2117 (N_2117,N_862,N_1462);
and U2118 (N_2118,N_1025,N_1289);
and U2119 (N_2119,N_1265,N_994);
xnor U2120 (N_2120,N_1341,N_955);
xor U2121 (N_2121,N_1238,N_1137);
and U2122 (N_2122,N_794,N_1343);
nor U2123 (N_2123,N_795,N_836);
nand U2124 (N_2124,N_793,N_916);
or U2125 (N_2125,N_1277,N_1223);
or U2126 (N_2126,N_1405,N_1042);
or U2127 (N_2127,N_1068,N_1350);
nand U2128 (N_2128,N_893,N_1002);
xnor U2129 (N_2129,N_1067,N_1253);
nor U2130 (N_2130,N_1085,N_1134);
nor U2131 (N_2131,N_886,N_1397);
nand U2132 (N_2132,N_1375,N_1427);
xnor U2133 (N_2133,N_1496,N_945);
nor U2134 (N_2134,N_976,N_795);
xnor U2135 (N_2135,N_1083,N_1495);
nand U2136 (N_2136,N_1366,N_1241);
nand U2137 (N_2137,N_982,N_1061);
and U2138 (N_2138,N_841,N_913);
nand U2139 (N_2139,N_1365,N_920);
nand U2140 (N_2140,N_1380,N_1278);
nand U2141 (N_2141,N_953,N_1327);
nor U2142 (N_2142,N_1239,N_1214);
nor U2143 (N_2143,N_938,N_1397);
nor U2144 (N_2144,N_1155,N_808);
and U2145 (N_2145,N_1146,N_1016);
nor U2146 (N_2146,N_1472,N_1491);
or U2147 (N_2147,N_1259,N_1495);
and U2148 (N_2148,N_989,N_1392);
and U2149 (N_2149,N_982,N_1264);
and U2150 (N_2150,N_952,N_1316);
nand U2151 (N_2151,N_933,N_1211);
or U2152 (N_2152,N_1349,N_925);
and U2153 (N_2153,N_1155,N_1376);
nand U2154 (N_2154,N_919,N_1305);
nand U2155 (N_2155,N_1349,N_964);
nor U2156 (N_2156,N_1250,N_1201);
nor U2157 (N_2157,N_1378,N_816);
nor U2158 (N_2158,N_860,N_1266);
or U2159 (N_2159,N_907,N_1092);
or U2160 (N_2160,N_998,N_1208);
nand U2161 (N_2161,N_956,N_777);
nand U2162 (N_2162,N_1391,N_955);
nor U2163 (N_2163,N_1210,N_972);
nor U2164 (N_2164,N_1034,N_1442);
or U2165 (N_2165,N_776,N_1054);
nor U2166 (N_2166,N_828,N_1477);
nor U2167 (N_2167,N_1277,N_912);
nor U2168 (N_2168,N_1274,N_764);
nor U2169 (N_2169,N_1368,N_1487);
nor U2170 (N_2170,N_1343,N_1144);
nand U2171 (N_2171,N_812,N_1331);
nor U2172 (N_2172,N_946,N_1493);
or U2173 (N_2173,N_1061,N_1417);
or U2174 (N_2174,N_1215,N_1081);
and U2175 (N_2175,N_1408,N_1497);
nor U2176 (N_2176,N_1069,N_1004);
and U2177 (N_2177,N_793,N_811);
and U2178 (N_2178,N_1144,N_1087);
and U2179 (N_2179,N_915,N_1434);
or U2180 (N_2180,N_1169,N_884);
or U2181 (N_2181,N_1440,N_1061);
and U2182 (N_2182,N_1350,N_815);
or U2183 (N_2183,N_1029,N_942);
nor U2184 (N_2184,N_1440,N_1232);
nor U2185 (N_2185,N_1099,N_1080);
nand U2186 (N_2186,N_1393,N_1002);
nor U2187 (N_2187,N_1183,N_1131);
or U2188 (N_2188,N_1319,N_909);
and U2189 (N_2189,N_1002,N_1323);
and U2190 (N_2190,N_818,N_1251);
or U2191 (N_2191,N_1271,N_1185);
or U2192 (N_2192,N_1024,N_904);
or U2193 (N_2193,N_1239,N_953);
and U2194 (N_2194,N_1011,N_1024);
and U2195 (N_2195,N_1088,N_1302);
or U2196 (N_2196,N_823,N_1132);
and U2197 (N_2197,N_1221,N_1011);
nor U2198 (N_2198,N_1450,N_1235);
xor U2199 (N_2199,N_1364,N_1003);
nor U2200 (N_2200,N_1098,N_1460);
and U2201 (N_2201,N_769,N_1334);
nor U2202 (N_2202,N_1196,N_800);
nand U2203 (N_2203,N_1148,N_1482);
or U2204 (N_2204,N_1161,N_877);
or U2205 (N_2205,N_815,N_833);
and U2206 (N_2206,N_942,N_964);
and U2207 (N_2207,N_1034,N_799);
nor U2208 (N_2208,N_1292,N_1037);
and U2209 (N_2209,N_1027,N_1421);
and U2210 (N_2210,N_1414,N_1489);
nor U2211 (N_2211,N_1004,N_1330);
and U2212 (N_2212,N_1182,N_1059);
nor U2213 (N_2213,N_1272,N_1145);
or U2214 (N_2214,N_854,N_1407);
nand U2215 (N_2215,N_1205,N_1156);
nand U2216 (N_2216,N_1341,N_1430);
nand U2217 (N_2217,N_1093,N_1451);
nor U2218 (N_2218,N_993,N_1194);
nand U2219 (N_2219,N_1139,N_935);
nand U2220 (N_2220,N_981,N_847);
or U2221 (N_2221,N_1088,N_1045);
and U2222 (N_2222,N_1373,N_827);
nand U2223 (N_2223,N_1112,N_1198);
and U2224 (N_2224,N_1165,N_997);
or U2225 (N_2225,N_1260,N_1485);
and U2226 (N_2226,N_1102,N_882);
or U2227 (N_2227,N_1151,N_755);
nor U2228 (N_2228,N_1320,N_1259);
or U2229 (N_2229,N_1244,N_930);
nand U2230 (N_2230,N_1346,N_1442);
nor U2231 (N_2231,N_1473,N_867);
nand U2232 (N_2232,N_998,N_1403);
xnor U2233 (N_2233,N_942,N_1468);
nand U2234 (N_2234,N_1463,N_979);
or U2235 (N_2235,N_961,N_916);
and U2236 (N_2236,N_878,N_1301);
nand U2237 (N_2237,N_906,N_850);
nor U2238 (N_2238,N_1149,N_1312);
and U2239 (N_2239,N_1152,N_1089);
nand U2240 (N_2240,N_1037,N_1023);
or U2241 (N_2241,N_1032,N_1334);
nand U2242 (N_2242,N_902,N_1185);
and U2243 (N_2243,N_1053,N_888);
and U2244 (N_2244,N_756,N_1002);
or U2245 (N_2245,N_1169,N_1352);
nand U2246 (N_2246,N_1074,N_1282);
nand U2247 (N_2247,N_857,N_1075);
nor U2248 (N_2248,N_1460,N_1428);
or U2249 (N_2249,N_840,N_1320);
nand U2250 (N_2250,N_1831,N_1529);
or U2251 (N_2251,N_1542,N_2227);
or U2252 (N_2252,N_2091,N_1829);
nand U2253 (N_2253,N_1580,N_1973);
nand U2254 (N_2254,N_1646,N_2169);
nor U2255 (N_2255,N_1846,N_2176);
and U2256 (N_2256,N_2014,N_1725);
or U2257 (N_2257,N_2185,N_1871);
nand U2258 (N_2258,N_1766,N_1563);
or U2259 (N_2259,N_1562,N_2055);
and U2260 (N_2260,N_1511,N_2145);
nor U2261 (N_2261,N_2222,N_2036);
or U2262 (N_2262,N_1988,N_2020);
xnor U2263 (N_2263,N_1697,N_1615);
and U2264 (N_2264,N_1716,N_1787);
nand U2265 (N_2265,N_2106,N_2130);
and U2266 (N_2266,N_2002,N_1554);
and U2267 (N_2267,N_1525,N_2080);
nand U2268 (N_2268,N_2008,N_1971);
and U2269 (N_2269,N_1944,N_2111);
nand U2270 (N_2270,N_1566,N_1813);
and U2271 (N_2271,N_2060,N_1791);
nor U2272 (N_2272,N_1966,N_1658);
or U2273 (N_2273,N_1885,N_2128);
and U2274 (N_2274,N_2153,N_1572);
or U2275 (N_2275,N_1873,N_2096);
and U2276 (N_2276,N_1962,N_2129);
nor U2277 (N_2277,N_2160,N_1760);
or U2278 (N_2278,N_2170,N_1628);
and U2279 (N_2279,N_2168,N_1901);
and U2280 (N_2280,N_1645,N_2074);
and U2281 (N_2281,N_1710,N_2174);
and U2282 (N_2282,N_1812,N_1505);
nand U2283 (N_2283,N_1926,N_1798);
and U2284 (N_2284,N_1826,N_1834);
or U2285 (N_2285,N_1877,N_1776);
or U2286 (N_2286,N_1661,N_2127);
nand U2287 (N_2287,N_1659,N_1643);
or U2288 (N_2288,N_1581,N_1539);
or U2289 (N_2289,N_1848,N_1941);
nand U2290 (N_2290,N_2249,N_2134);
nor U2291 (N_2291,N_1998,N_2173);
and U2292 (N_2292,N_1837,N_1928);
and U2293 (N_2293,N_1672,N_1815);
nand U2294 (N_2294,N_1788,N_2090);
nand U2295 (N_2295,N_2162,N_1553);
nand U2296 (N_2296,N_1743,N_1586);
or U2297 (N_2297,N_1949,N_1548);
or U2298 (N_2298,N_1981,N_1683);
nand U2299 (N_2299,N_2165,N_1573);
and U2300 (N_2300,N_2196,N_1509);
nor U2301 (N_2301,N_1731,N_1689);
or U2302 (N_2302,N_1965,N_1800);
or U2303 (N_2303,N_2052,N_2208);
or U2304 (N_2304,N_1501,N_2120);
nor U2305 (N_2305,N_1934,N_1518);
or U2306 (N_2306,N_1946,N_1708);
and U2307 (N_2307,N_1614,N_1742);
and U2308 (N_2308,N_1520,N_1709);
nor U2309 (N_2309,N_2105,N_1920);
nor U2310 (N_2310,N_1681,N_2190);
or U2311 (N_2311,N_1942,N_1889);
or U2312 (N_2312,N_2157,N_1842);
and U2313 (N_2313,N_1881,N_1841);
and U2314 (N_2314,N_1602,N_2107);
nor U2315 (N_2315,N_1648,N_2137);
nand U2316 (N_2316,N_1574,N_1622);
or U2317 (N_2317,N_1951,N_2067);
and U2318 (N_2318,N_1647,N_2035);
and U2319 (N_2319,N_2199,N_1961);
nor U2320 (N_2320,N_2118,N_1968);
or U2321 (N_2321,N_1953,N_1705);
nand U2322 (N_2322,N_1891,N_2141);
or U2323 (N_2323,N_1764,N_1932);
nand U2324 (N_2324,N_2124,N_1820);
or U2325 (N_2325,N_1744,N_1758);
or U2326 (N_2326,N_2212,N_1950);
or U2327 (N_2327,N_1666,N_2018);
nand U2328 (N_2328,N_2146,N_1836);
or U2329 (N_2329,N_1624,N_2037);
nand U2330 (N_2330,N_2030,N_1991);
nor U2331 (N_2331,N_1610,N_1723);
and U2332 (N_2332,N_2063,N_2187);
or U2333 (N_2333,N_1801,N_1783);
nand U2334 (N_2334,N_2047,N_1835);
and U2335 (N_2335,N_1995,N_2163);
or U2336 (N_2336,N_1908,N_1590);
nor U2337 (N_2337,N_1986,N_1588);
nand U2338 (N_2338,N_2087,N_2045);
nor U2339 (N_2339,N_1872,N_2103);
or U2340 (N_2340,N_2242,N_1858);
nand U2341 (N_2341,N_1746,N_1630);
and U2342 (N_2342,N_1990,N_1851);
nand U2343 (N_2343,N_1523,N_1938);
or U2344 (N_2344,N_1840,N_2081);
nor U2345 (N_2345,N_1636,N_1538);
or U2346 (N_2346,N_1900,N_2028);
or U2347 (N_2347,N_1568,N_1954);
xor U2348 (N_2348,N_2101,N_1671);
and U2349 (N_2349,N_1866,N_1641);
and U2350 (N_2350,N_1832,N_1748);
nand U2351 (N_2351,N_1603,N_1514);
or U2352 (N_2352,N_1605,N_1904);
nor U2353 (N_2353,N_1878,N_1741);
and U2354 (N_2354,N_1902,N_1660);
nor U2355 (N_2355,N_2201,N_2184);
and U2356 (N_2356,N_1888,N_1528);
or U2357 (N_2357,N_1515,N_2179);
nor U2358 (N_2358,N_2144,N_1668);
nand U2359 (N_2359,N_1897,N_1957);
and U2360 (N_2360,N_1856,N_2139);
nand U2361 (N_2361,N_1692,N_1870);
and U2362 (N_2362,N_1854,N_1594);
nor U2363 (N_2363,N_1596,N_1730);
nand U2364 (N_2364,N_1597,N_2076);
or U2365 (N_2365,N_1584,N_1571);
nor U2366 (N_2366,N_1770,N_1909);
or U2367 (N_2367,N_2217,N_1805);
and U2368 (N_2368,N_1508,N_1535);
nor U2369 (N_2369,N_2248,N_2099);
and U2370 (N_2370,N_1565,N_2016);
and U2371 (N_2371,N_1859,N_1694);
or U2372 (N_2372,N_1868,N_2131);
nor U2373 (N_2373,N_1773,N_2204);
nand U2374 (N_2374,N_2050,N_1550);
nor U2375 (N_2375,N_2155,N_2138);
and U2376 (N_2376,N_2188,N_1775);
and U2377 (N_2377,N_1952,N_1632);
nand U2378 (N_2378,N_2125,N_1917);
nor U2379 (N_2379,N_2186,N_1931);
nand U2380 (N_2380,N_2246,N_2164);
and U2381 (N_2381,N_2244,N_2051);
nor U2382 (N_2382,N_1778,N_1862);
and U2383 (N_2383,N_1827,N_1654);
or U2384 (N_2384,N_1886,N_1863);
nor U2385 (N_2385,N_2075,N_2082);
nor U2386 (N_2386,N_2073,N_1676);
or U2387 (N_2387,N_1793,N_1611);
and U2388 (N_2388,N_1945,N_1567);
nand U2389 (N_2389,N_2049,N_1806);
and U2390 (N_2390,N_1703,N_1513);
and U2391 (N_2391,N_1751,N_2236);
or U2392 (N_2392,N_1557,N_1790);
nor U2393 (N_2393,N_1559,N_1960);
nor U2394 (N_2394,N_1983,N_2033);
xnor U2395 (N_2395,N_2114,N_2159);
nor U2396 (N_2396,N_1750,N_2215);
and U2397 (N_2397,N_1560,N_1652);
nand U2398 (N_2398,N_2226,N_2247);
nor U2399 (N_2399,N_2024,N_1925);
or U2400 (N_2400,N_2143,N_1845);
and U2401 (N_2401,N_1556,N_2245);
nand U2402 (N_2402,N_1644,N_1534);
nand U2403 (N_2403,N_1687,N_1651);
nand U2404 (N_2404,N_1822,N_1795);
and U2405 (N_2405,N_1507,N_1627);
or U2406 (N_2406,N_1579,N_1818);
or U2407 (N_2407,N_1601,N_1718);
and U2408 (N_2408,N_2202,N_2189);
nor U2409 (N_2409,N_2092,N_2019);
nand U2410 (N_2410,N_1914,N_1617);
and U2411 (N_2411,N_1887,N_2011);
and U2412 (N_2412,N_1823,N_1635);
and U2413 (N_2413,N_2180,N_1591);
or U2414 (N_2414,N_1616,N_2191);
or U2415 (N_2415,N_1655,N_2219);
nor U2416 (N_2416,N_1940,N_1974);
or U2417 (N_2417,N_1752,N_2149);
nor U2418 (N_2418,N_2025,N_1698);
or U2419 (N_2419,N_1734,N_1702);
nor U2420 (N_2420,N_1719,N_2006);
or U2421 (N_2421,N_2150,N_1921);
and U2422 (N_2422,N_1516,N_1912);
and U2423 (N_2423,N_1879,N_1738);
nor U2424 (N_2424,N_1555,N_1656);
or U2425 (N_2425,N_1977,N_1970);
nand U2426 (N_2426,N_1850,N_2000);
nand U2427 (N_2427,N_1500,N_1869);
and U2428 (N_2428,N_2098,N_2009);
and U2429 (N_2429,N_1896,N_2234);
nand U2430 (N_2430,N_1558,N_1882);
nor U2431 (N_2431,N_2243,N_1670);
and U2432 (N_2432,N_2056,N_1544);
or U2433 (N_2433,N_2123,N_1789);
nand U2434 (N_2434,N_1722,N_2239);
nand U2435 (N_2435,N_1657,N_2086);
or U2436 (N_2436,N_1607,N_1996);
and U2437 (N_2437,N_2216,N_1989);
nand U2438 (N_2438,N_2083,N_1675);
xor U2439 (N_2439,N_1592,N_2210);
nor U2440 (N_2440,N_1502,N_1913);
nand U2441 (N_2441,N_1922,N_1807);
nand U2442 (N_2442,N_1701,N_1852);
or U2443 (N_2443,N_1633,N_1849);
or U2444 (N_2444,N_1691,N_1906);
nor U2445 (N_2445,N_1662,N_2079);
nand U2446 (N_2446,N_1857,N_1665);
nand U2447 (N_2447,N_1963,N_1915);
and U2448 (N_2448,N_1637,N_2094);
and U2449 (N_2449,N_2154,N_2078);
nor U2450 (N_2450,N_1564,N_2034);
and U2451 (N_2451,N_2031,N_1740);
or U2452 (N_2452,N_2233,N_1893);
nand U2453 (N_2453,N_1865,N_2178);
or U2454 (N_2454,N_1819,N_1677);
and U2455 (N_2455,N_2003,N_1690);
or U2456 (N_2456,N_2061,N_1583);
or U2457 (N_2457,N_1549,N_1679);
nand U2458 (N_2458,N_1796,N_1811);
nand U2459 (N_2459,N_1804,N_2228);
nor U2460 (N_2460,N_2133,N_1855);
or U2461 (N_2461,N_1833,N_2237);
or U2462 (N_2462,N_1861,N_1506);
nand U2463 (N_2463,N_1994,N_1980);
or U2464 (N_2464,N_1794,N_1761);
xnor U2465 (N_2465,N_1907,N_2238);
or U2466 (N_2466,N_2007,N_1682);
xor U2467 (N_2467,N_1510,N_1726);
and U2468 (N_2468,N_1784,N_2057);
nor U2469 (N_2469,N_1930,N_2070);
nor U2470 (N_2470,N_1967,N_1875);
nor U2471 (N_2471,N_2213,N_1598);
and U2472 (N_2472,N_2182,N_1543);
or U2473 (N_2473,N_1623,N_1969);
or U2474 (N_2474,N_1620,N_1604);
and U2475 (N_2475,N_1987,N_1985);
nor U2476 (N_2476,N_1678,N_1638);
or U2477 (N_2477,N_2241,N_2093);
or U2478 (N_2478,N_2206,N_1979);
xor U2479 (N_2479,N_1929,N_1927);
or U2480 (N_2480,N_2004,N_1541);
and U2481 (N_2481,N_2230,N_1608);
or U2482 (N_2482,N_2100,N_1768);
or U2483 (N_2483,N_2203,N_2108);
nor U2484 (N_2484,N_2117,N_1771);
nor U2485 (N_2485,N_2088,N_2113);
nor U2486 (N_2486,N_1814,N_1700);
or U2487 (N_2487,N_1905,N_2043);
nor U2488 (N_2488,N_1552,N_1755);
nor U2489 (N_2489,N_1809,N_1577);
nand U2490 (N_2490,N_2235,N_2112);
and U2491 (N_2491,N_1747,N_1729);
and U2492 (N_2492,N_2110,N_2231);
nand U2493 (N_2493,N_2209,N_1984);
or U2494 (N_2494,N_2029,N_1839);
nor U2495 (N_2495,N_1828,N_1728);
or U2496 (N_2496,N_2054,N_1792);
and U2497 (N_2497,N_1959,N_1774);
nor U2498 (N_2498,N_2224,N_2013);
xor U2499 (N_2499,N_1844,N_2071);
and U2500 (N_2500,N_1649,N_1585);
or U2501 (N_2501,N_1517,N_2042);
nor U2502 (N_2502,N_1883,N_1587);
nand U2503 (N_2503,N_2194,N_1777);
nand U2504 (N_2504,N_1578,N_2122);
nor U2505 (N_2505,N_2089,N_1561);
and U2506 (N_2506,N_1757,N_1547);
nand U2507 (N_2507,N_2147,N_1880);
and U2508 (N_2508,N_2175,N_1802);
nor U2509 (N_2509,N_1993,N_1720);
nand U2510 (N_2510,N_1634,N_1551);
nor U2511 (N_2511,N_1972,N_2161);
and U2512 (N_2512,N_2022,N_1680);
nand U2513 (N_2513,N_1684,N_2005);
or U2514 (N_2514,N_2062,N_1874);
nor U2515 (N_2515,N_1899,N_1753);
nor U2516 (N_2516,N_2229,N_2017);
and U2517 (N_2517,N_1919,N_2027);
nor U2518 (N_2518,N_1612,N_2132);
nand U2519 (N_2519,N_2152,N_1895);
nand U2520 (N_2520,N_1817,N_2142);
nor U2521 (N_2521,N_1745,N_2097);
nor U2522 (N_2522,N_2015,N_1733);
or U2523 (N_2523,N_1799,N_1727);
nand U2524 (N_2524,N_2148,N_2064);
and U2525 (N_2525,N_2046,N_2012);
nand U2526 (N_2526,N_1704,N_1504);
nand U2527 (N_2527,N_1876,N_1898);
and U2528 (N_2528,N_1699,N_1524);
nor U2529 (N_2529,N_1540,N_2223);
nand U2530 (N_2530,N_2225,N_2040);
and U2531 (N_2531,N_1736,N_1923);
and U2532 (N_2532,N_1955,N_1582);
and U2533 (N_2533,N_1939,N_1976);
nor U2534 (N_2534,N_1531,N_1824);
and U2535 (N_2535,N_1911,N_2023);
nor U2536 (N_2536,N_2084,N_1735);
and U2537 (N_2537,N_1759,N_1711);
and U2538 (N_2538,N_2021,N_1521);
and U2539 (N_2539,N_1707,N_1803);
nor U2540 (N_2540,N_1937,N_2032);
nor U2541 (N_2541,N_1712,N_2058);
and U2542 (N_2542,N_2072,N_2121);
nand U2543 (N_2543,N_2053,N_2192);
nor U2544 (N_2544,N_1780,N_2026);
nand U2545 (N_2545,N_1522,N_1715);
nand U2546 (N_2546,N_2193,N_1884);
nor U2547 (N_2547,N_2220,N_2177);
or U2548 (N_2548,N_1629,N_2200);
or U2549 (N_2549,N_1650,N_2240);
or U2550 (N_2550,N_2140,N_1958);
xor U2551 (N_2551,N_2104,N_1695);
and U2552 (N_2552,N_2172,N_1639);
nor U2553 (N_2553,N_1589,N_1956);
nand U2554 (N_2554,N_1943,N_2044);
nor U2555 (N_2555,N_2039,N_2195);
or U2556 (N_2556,N_1642,N_1892);
nor U2557 (N_2557,N_1536,N_2126);
and U2558 (N_2558,N_1935,N_1527);
nand U2559 (N_2559,N_1621,N_1537);
or U2560 (N_2560,N_2136,N_1686);
and U2561 (N_2561,N_2119,N_1864);
and U2562 (N_2562,N_1546,N_1673);
and U2563 (N_2563,N_1674,N_1890);
and U2564 (N_2564,N_1570,N_1714);
nor U2565 (N_2565,N_2102,N_1626);
nand U2566 (N_2566,N_1903,N_1847);
nor U2567 (N_2567,N_1948,N_1860);
nand U2568 (N_2568,N_1545,N_1664);
or U2569 (N_2569,N_1756,N_1693);
or U2570 (N_2570,N_1982,N_1772);
or U2571 (N_2571,N_1825,N_1816);
or U2572 (N_2572,N_1625,N_2068);
and U2573 (N_2573,N_1997,N_1838);
and U2574 (N_2574,N_2183,N_1754);
nand U2575 (N_2575,N_2198,N_1503);
nor U2576 (N_2576,N_2207,N_2001);
nand U2577 (N_2577,N_2151,N_1526);
nand U2578 (N_2578,N_1706,N_1779);
nor U2579 (N_2579,N_1867,N_2069);
nor U2580 (N_2580,N_1762,N_1782);
or U2581 (N_2581,N_1724,N_1749);
nand U2582 (N_2582,N_1618,N_1609);
or U2583 (N_2583,N_1853,N_1640);
nor U2584 (N_2584,N_1519,N_1786);
nor U2585 (N_2585,N_2221,N_2010);
and U2586 (N_2586,N_1685,N_2109);
and U2587 (N_2587,N_1575,N_1916);
and U2588 (N_2588,N_1732,N_2116);
and U2589 (N_2589,N_2059,N_1595);
nor U2590 (N_2590,N_2166,N_2077);
nor U2591 (N_2591,N_1781,N_1894);
or U2592 (N_2592,N_1924,N_1600);
nor U2593 (N_2593,N_2167,N_1739);
nor U2594 (N_2594,N_2065,N_2218);
and U2595 (N_2595,N_1593,N_1688);
or U2596 (N_2596,N_1696,N_1975);
xnor U2597 (N_2597,N_1978,N_1653);
and U2598 (N_2598,N_1721,N_1613);
nor U2599 (N_2599,N_2158,N_1830);
and U2600 (N_2600,N_1843,N_1999);
nor U2601 (N_2601,N_1933,N_1606);
xnor U2602 (N_2602,N_2115,N_1936);
or U2603 (N_2603,N_2041,N_1512);
nand U2604 (N_2604,N_2095,N_2197);
nand U2605 (N_2605,N_2205,N_2232);
and U2606 (N_2606,N_1785,N_1964);
or U2607 (N_2607,N_1599,N_1713);
or U2608 (N_2608,N_1918,N_1797);
nand U2609 (N_2609,N_2085,N_1737);
or U2610 (N_2610,N_2171,N_1992);
nand U2611 (N_2611,N_1569,N_2214);
and U2612 (N_2612,N_1947,N_1669);
nor U2613 (N_2613,N_1530,N_1821);
and U2614 (N_2614,N_1667,N_2048);
nand U2615 (N_2615,N_2156,N_1767);
and U2616 (N_2616,N_2066,N_1619);
and U2617 (N_2617,N_1910,N_1765);
nand U2618 (N_2618,N_2038,N_1810);
or U2619 (N_2619,N_2135,N_2181);
or U2620 (N_2620,N_2211,N_1663);
or U2621 (N_2621,N_1808,N_1769);
nand U2622 (N_2622,N_1533,N_1532);
nor U2623 (N_2623,N_1763,N_1631);
or U2624 (N_2624,N_1717,N_1576);
nor U2625 (N_2625,N_1996,N_2138);
nand U2626 (N_2626,N_1622,N_1978);
nor U2627 (N_2627,N_1868,N_2161);
and U2628 (N_2628,N_1563,N_1525);
and U2629 (N_2629,N_2053,N_1858);
or U2630 (N_2630,N_2211,N_1934);
and U2631 (N_2631,N_2144,N_1838);
xnor U2632 (N_2632,N_1932,N_2042);
nand U2633 (N_2633,N_1784,N_2060);
or U2634 (N_2634,N_1826,N_1538);
nor U2635 (N_2635,N_1508,N_2216);
nand U2636 (N_2636,N_1704,N_1891);
nor U2637 (N_2637,N_2209,N_1781);
nand U2638 (N_2638,N_1824,N_1918);
and U2639 (N_2639,N_1867,N_1662);
or U2640 (N_2640,N_2227,N_1764);
nor U2641 (N_2641,N_2193,N_2226);
nand U2642 (N_2642,N_2043,N_1799);
nand U2643 (N_2643,N_2192,N_1566);
nor U2644 (N_2644,N_1932,N_2123);
nand U2645 (N_2645,N_2122,N_2092);
nor U2646 (N_2646,N_1817,N_2240);
or U2647 (N_2647,N_2110,N_2046);
or U2648 (N_2648,N_1660,N_1571);
xor U2649 (N_2649,N_2210,N_1799);
nor U2650 (N_2650,N_2242,N_1894);
nor U2651 (N_2651,N_2008,N_1830);
nor U2652 (N_2652,N_2016,N_2140);
nand U2653 (N_2653,N_1720,N_2212);
or U2654 (N_2654,N_2057,N_1684);
and U2655 (N_2655,N_2018,N_2142);
and U2656 (N_2656,N_1714,N_1900);
nor U2657 (N_2657,N_1591,N_2098);
nand U2658 (N_2658,N_1641,N_2008);
or U2659 (N_2659,N_1826,N_1512);
and U2660 (N_2660,N_1838,N_1764);
nand U2661 (N_2661,N_2035,N_1995);
and U2662 (N_2662,N_2057,N_1826);
or U2663 (N_2663,N_1986,N_1643);
or U2664 (N_2664,N_2191,N_2118);
or U2665 (N_2665,N_2051,N_1985);
nor U2666 (N_2666,N_1967,N_2238);
and U2667 (N_2667,N_1858,N_2057);
and U2668 (N_2668,N_1832,N_1958);
or U2669 (N_2669,N_2210,N_1536);
nor U2670 (N_2670,N_1612,N_2133);
or U2671 (N_2671,N_1641,N_1541);
or U2672 (N_2672,N_1595,N_2028);
or U2673 (N_2673,N_1799,N_2221);
or U2674 (N_2674,N_2026,N_1615);
nor U2675 (N_2675,N_2233,N_2023);
nor U2676 (N_2676,N_2048,N_1953);
or U2677 (N_2677,N_1666,N_1520);
or U2678 (N_2678,N_2045,N_1777);
nand U2679 (N_2679,N_2105,N_2127);
nor U2680 (N_2680,N_1992,N_2210);
or U2681 (N_2681,N_1834,N_1773);
or U2682 (N_2682,N_1560,N_1721);
and U2683 (N_2683,N_2048,N_1974);
nand U2684 (N_2684,N_1558,N_1819);
nor U2685 (N_2685,N_2095,N_1902);
nand U2686 (N_2686,N_1986,N_1654);
nor U2687 (N_2687,N_2116,N_1740);
nand U2688 (N_2688,N_1899,N_1804);
xnor U2689 (N_2689,N_2001,N_1941);
nor U2690 (N_2690,N_2069,N_1698);
nor U2691 (N_2691,N_1920,N_1595);
and U2692 (N_2692,N_1850,N_1926);
and U2693 (N_2693,N_1864,N_2197);
nor U2694 (N_2694,N_1765,N_1661);
nand U2695 (N_2695,N_1594,N_1892);
and U2696 (N_2696,N_2202,N_1502);
or U2697 (N_2697,N_1646,N_1707);
nand U2698 (N_2698,N_1518,N_1689);
nor U2699 (N_2699,N_2033,N_2151);
nor U2700 (N_2700,N_1839,N_2192);
and U2701 (N_2701,N_1926,N_1948);
nand U2702 (N_2702,N_1611,N_2091);
or U2703 (N_2703,N_1735,N_2168);
or U2704 (N_2704,N_1541,N_2038);
and U2705 (N_2705,N_1696,N_2173);
and U2706 (N_2706,N_1749,N_2239);
nor U2707 (N_2707,N_1678,N_1964);
and U2708 (N_2708,N_2066,N_1804);
or U2709 (N_2709,N_1976,N_2101);
nor U2710 (N_2710,N_1960,N_1920);
or U2711 (N_2711,N_1738,N_1972);
nor U2712 (N_2712,N_2051,N_1927);
nor U2713 (N_2713,N_1907,N_2130);
nand U2714 (N_2714,N_1897,N_1563);
xnor U2715 (N_2715,N_1680,N_1656);
and U2716 (N_2716,N_1805,N_2055);
nor U2717 (N_2717,N_2132,N_2209);
nand U2718 (N_2718,N_1673,N_2216);
nor U2719 (N_2719,N_1678,N_2117);
or U2720 (N_2720,N_1676,N_1773);
nand U2721 (N_2721,N_2185,N_1872);
and U2722 (N_2722,N_1921,N_1608);
nor U2723 (N_2723,N_1517,N_1777);
nor U2724 (N_2724,N_1692,N_2087);
xor U2725 (N_2725,N_1664,N_1873);
or U2726 (N_2726,N_2212,N_1912);
and U2727 (N_2727,N_1546,N_2233);
or U2728 (N_2728,N_1879,N_2127);
nor U2729 (N_2729,N_2240,N_2164);
or U2730 (N_2730,N_2210,N_1588);
nor U2731 (N_2731,N_2205,N_1568);
nand U2732 (N_2732,N_1893,N_1815);
nand U2733 (N_2733,N_1624,N_1511);
or U2734 (N_2734,N_2185,N_1635);
or U2735 (N_2735,N_1685,N_1557);
or U2736 (N_2736,N_1849,N_1610);
nand U2737 (N_2737,N_2118,N_1901);
or U2738 (N_2738,N_2006,N_1952);
or U2739 (N_2739,N_1904,N_1912);
or U2740 (N_2740,N_2091,N_2030);
and U2741 (N_2741,N_2245,N_1824);
and U2742 (N_2742,N_1861,N_2000);
or U2743 (N_2743,N_2123,N_1733);
or U2744 (N_2744,N_1695,N_1525);
nand U2745 (N_2745,N_2073,N_2169);
and U2746 (N_2746,N_1729,N_2080);
and U2747 (N_2747,N_2216,N_1526);
xor U2748 (N_2748,N_2092,N_1623);
nand U2749 (N_2749,N_1567,N_2240);
nor U2750 (N_2750,N_1996,N_2180);
and U2751 (N_2751,N_1589,N_1869);
nor U2752 (N_2752,N_2236,N_1914);
nand U2753 (N_2753,N_1809,N_1773);
nand U2754 (N_2754,N_2119,N_2191);
or U2755 (N_2755,N_1867,N_1830);
nand U2756 (N_2756,N_2069,N_1515);
nor U2757 (N_2757,N_1965,N_1638);
nand U2758 (N_2758,N_2139,N_2043);
nor U2759 (N_2759,N_1635,N_1709);
and U2760 (N_2760,N_1941,N_1815);
nand U2761 (N_2761,N_1727,N_2116);
and U2762 (N_2762,N_2219,N_1762);
and U2763 (N_2763,N_2121,N_1952);
or U2764 (N_2764,N_1743,N_1950);
and U2765 (N_2765,N_1740,N_2193);
nor U2766 (N_2766,N_1842,N_1526);
nor U2767 (N_2767,N_2247,N_1675);
and U2768 (N_2768,N_2101,N_1783);
nor U2769 (N_2769,N_1739,N_1515);
or U2770 (N_2770,N_1974,N_1692);
or U2771 (N_2771,N_2046,N_2140);
and U2772 (N_2772,N_1528,N_1691);
nand U2773 (N_2773,N_2024,N_1579);
or U2774 (N_2774,N_2225,N_2049);
and U2775 (N_2775,N_1940,N_1673);
or U2776 (N_2776,N_1753,N_2215);
and U2777 (N_2777,N_1699,N_2042);
and U2778 (N_2778,N_1754,N_1745);
and U2779 (N_2779,N_1667,N_2031);
and U2780 (N_2780,N_1996,N_1902);
xor U2781 (N_2781,N_2094,N_2118);
and U2782 (N_2782,N_2052,N_1872);
or U2783 (N_2783,N_2179,N_1605);
nor U2784 (N_2784,N_1589,N_1773);
nand U2785 (N_2785,N_1791,N_1629);
nor U2786 (N_2786,N_2155,N_1820);
nor U2787 (N_2787,N_1593,N_1847);
and U2788 (N_2788,N_2176,N_2083);
and U2789 (N_2789,N_1787,N_1665);
nor U2790 (N_2790,N_2228,N_2213);
or U2791 (N_2791,N_1780,N_1520);
nor U2792 (N_2792,N_1531,N_2125);
or U2793 (N_2793,N_2010,N_2006);
or U2794 (N_2794,N_2146,N_1893);
and U2795 (N_2795,N_1958,N_1739);
and U2796 (N_2796,N_1567,N_2222);
nand U2797 (N_2797,N_1691,N_2028);
or U2798 (N_2798,N_2151,N_1868);
nand U2799 (N_2799,N_1940,N_1874);
nor U2800 (N_2800,N_1736,N_1572);
nor U2801 (N_2801,N_2100,N_1669);
and U2802 (N_2802,N_1709,N_2090);
and U2803 (N_2803,N_2236,N_2169);
xnor U2804 (N_2804,N_1974,N_1543);
or U2805 (N_2805,N_2046,N_1505);
or U2806 (N_2806,N_1524,N_1914);
nand U2807 (N_2807,N_1775,N_2119);
or U2808 (N_2808,N_1992,N_1554);
and U2809 (N_2809,N_1957,N_1605);
nor U2810 (N_2810,N_1788,N_1750);
or U2811 (N_2811,N_1860,N_1687);
and U2812 (N_2812,N_1733,N_1619);
nor U2813 (N_2813,N_2160,N_2242);
nor U2814 (N_2814,N_1742,N_2021);
nand U2815 (N_2815,N_1764,N_1520);
nand U2816 (N_2816,N_1905,N_2162);
nor U2817 (N_2817,N_1705,N_1751);
or U2818 (N_2818,N_2245,N_1859);
or U2819 (N_2819,N_2108,N_2042);
nor U2820 (N_2820,N_1866,N_1906);
nor U2821 (N_2821,N_1551,N_1730);
nand U2822 (N_2822,N_1858,N_1861);
and U2823 (N_2823,N_2112,N_1504);
nand U2824 (N_2824,N_1763,N_2007);
and U2825 (N_2825,N_2247,N_1527);
nor U2826 (N_2826,N_1591,N_2221);
nor U2827 (N_2827,N_2204,N_2022);
nor U2828 (N_2828,N_1722,N_2074);
or U2829 (N_2829,N_1569,N_1524);
nand U2830 (N_2830,N_1809,N_1882);
and U2831 (N_2831,N_1608,N_1721);
and U2832 (N_2832,N_1730,N_1746);
nand U2833 (N_2833,N_1797,N_2102);
and U2834 (N_2834,N_1580,N_2214);
or U2835 (N_2835,N_1594,N_2012);
and U2836 (N_2836,N_2034,N_1810);
or U2837 (N_2837,N_2143,N_1625);
nand U2838 (N_2838,N_1669,N_1598);
xnor U2839 (N_2839,N_2154,N_2115);
or U2840 (N_2840,N_2031,N_2038);
nand U2841 (N_2841,N_2009,N_1550);
and U2842 (N_2842,N_1884,N_2061);
and U2843 (N_2843,N_1973,N_1754);
and U2844 (N_2844,N_1904,N_1535);
and U2845 (N_2845,N_1542,N_1814);
nand U2846 (N_2846,N_1646,N_1854);
and U2847 (N_2847,N_2141,N_1537);
or U2848 (N_2848,N_2232,N_1873);
nor U2849 (N_2849,N_1542,N_1519);
and U2850 (N_2850,N_1586,N_1573);
and U2851 (N_2851,N_1992,N_1908);
nand U2852 (N_2852,N_2102,N_1586);
or U2853 (N_2853,N_1807,N_2076);
or U2854 (N_2854,N_2121,N_1582);
and U2855 (N_2855,N_1695,N_2201);
nand U2856 (N_2856,N_1904,N_1981);
and U2857 (N_2857,N_1803,N_1960);
or U2858 (N_2858,N_1780,N_2083);
nand U2859 (N_2859,N_1845,N_1651);
nand U2860 (N_2860,N_1661,N_2145);
xnor U2861 (N_2861,N_1636,N_2200);
and U2862 (N_2862,N_1558,N_1996);
nor U2863 (N_2863,N_1942,N_1805);
and U2864 (N_2864,N_1880,N_2152);
nand U2865 (N_2865,N_1963,N_1512);
nand U2866 (N_2866,N_1842,N_2139);
and U2867 (N_2867,N_2148,N_1666);
and U2868 (N_2868,N_1786,N_1659);
nand U2869 (N_2869,N_1716,N_1623);
or U2870 (N_2870,N_1957,N_1632);
nor U2871 (N_2871,N_1929,N_1611);
nor U2872 (N_2872,N_1893,N_1789);
or U2873 (N_2873,N_1659,N_2144);
nor U2874 (N_2874,N_1556,N_2058);
and U2875 (N_2875,N_2070,N_2015);
nand U2876 (N_2876,N_2159,N_1853);
or U2877 (N_2877,N_1869,N_2233);
or U2878 (N_2878,N_1557,N_1933);
and U2879 (N_2879,N_2243,N_2039);
or U2880 (N_2880,N_2027,N_2065);
nand U2881 (N_2881,N_1699,N_2111);
nor U2882 (N_2882,N_2209,N_1506);
or U2883 (N_2883,N_1903,N_2231);
and U2884 (N_2884,N_1702,N_1520);
nor U2885 (N_2885,N_1523,N_2039);
and U2886 (N_2886,N_1983,N_2041);
nand U2887 (N_2887,N_1877,N_2168);
or U2888 (N_2888,N_1847,N_2148);
nand U2889 (N_2889,N_1717,N_2154);
nor U2890 (N_2890,N_1769,N_2091);
nor U2891 (N_2891,N_2224,N_2056);
or U2892 (N_2892,N_1589,N_1818);
nand U2893 (N_2893,N_1583,N_2135);
or U2894 (N_2894,N_1578,N_2003);
nand U2895 (N_2895,N_2209,N_2076);
nand U2896 (N_2896,N_1749,N_1802);
nor U2897 (N_2897,N_1659,N_2028);
or U2898 (N_2898,N_1992,N_2167);
or U2899 (N_2899,N_2024,N_1859);
nand U2900 (N_2900,N_1739,N_1744);
and U2901 (N_2901,N_1814,N_2088);
nor U2902 (N_2902,N_2233,N_1824);
or U2903 (N_2903,N_1562,N_2075);
nor U2904 (N_2904,N_1883,N_1613);
or U2905 (N_2905,N_1835,N_2182);
nor U2906 (N_2906,N_2064,N_1634);
nand U2907 (N_2907,N_1828,N_1808);
xnor U2908 (N_2908,N_2207,N_1826);
or U2909 (N_2909,N_1728,N_2164);
nand U2910 (N_2910,N_1517,N_1970);
nand U2911 (N_2911,N_1510,N_1698);
or U2912 (N_2912,N_1581,N_1738);
nor U2913 (N_2913,N_1722,N_1945);
or U2914 (N_2914,N_1886,N_1610);
nor U2915 (N_2915,N_1736,N_2164);
nand U2916 (N_2916,N_1731,N_1860);
xnor U2917 (N_2917,N_1754,N_1822);
nor U2918 (N_2918,N_1859,N_1879);
and U2919 (N_2919,N_1967,N_1927);
nand U2920 (N_2920,N_1854,N_1519);
and U2921 (N_2921,N_2223,N_2071);
nor U2922 (N_2922,N_1629,N_1607);
and U2923 (N_2923,N_1743,N_1670);
nor U2924 (N_2924,N_2051,N_1838);
nor U2925 (N_2925,N_1886,N_1668);
and U2926 (N_2926,N_1760,N_1913);
and U2927 (N_2927,N_1581,N_2185);
nand U2928 (N_2928,N_2215,N_1557);
or U2929 (N_2929,N_1593,N_1807);
or U2930 (N_2930,N_1926,N_1879);
or U2931 (N_2931,N_1727,N_1724);
nand U2932 (N_2932,N_2107,N_1856);
and U2933 (N_2933,N_1881,N_1743);
nor U2934 (N_2934,N_1885,N_1986);
nand U2935 (N_2935,N_1643,N_2216);
and U2936 (N_2936,N_2034,N_1715);
nand U2937 (N_2937,N_1766,N_2246);
nand U2938 (N_2938,N_1683,N_1729);
nor U2939 (N_2939,N_1543,N_2231);
and U2940 (N_2940,N_2047,N_2226);
nand U2941 (N_2941,N_1676,N_1595);
or U2942 (N_2942,N_1840,N_1862);
nor U2943 (N_2943,N_2030,N_1758);
and U2944 (N_2944,N_2059,N_1544);
or U2945 (N_2945,N_1544,N_1683);
nand U2946 (N_2946,N_1588,N_1528);
and U2947 (N_2947,N_1908,N_2215);
nor U2948 (N_2948,N_1665,N_2147);
nand U2949 (N_2949,N_2247,N_1960);
nand U2950 (N_2950,N_1920,N_1509);
or U2951 (N_2951,N_2097,N_1614);
nor U2952 (N_2952,N_1523,N_2104);
nor U2953 (N_2953,N_2082,N_1853);
or U2954 (N_2954,N_1743,N_1879);
or U2955 (N_2955,N_1822,N_1688);
or U2956 (N_2956,N_1727,N_2005);
and U2957 (N_2957,N_1562,N_1521);
and U2958 (N_2958,N_1874,N_2167);
nand U2959 (N_2959,N_2133,N_2082);
nor U2960 (N_2960,N_2094,N_2056);
and U2961 (N_2961,N_1666,N_2135);
nand U2962 (N_2962,N_1613,N_1508);
nand U2963 (N_2963,N_2071,N_1686);
and U2964 (N_2964,N_2004,N_1638);
and U2965 (N_2965,N_1866,N_2211);
nand U2966 (N_2966,N_1587,N_1580);
nor U2967 (N_2967,N_1604,N_1550);
nor U2968 (N_2968,N_2144,N_1876);
nand U2969 (N_2969,N_2233,N_1620);
nand U2970 (N_2970,N_1960,N_2231);
or U2971 (N_2971,N_1994,N_1699);
xor U2972 (N_2972,N_1701,N_1747);
and U2973 (N_2973,N_1999,N_1698);
and U2974 (N_2974,N_1529,N_1548);
and U2975 (N_2975,N_1520,N_1931);
nor U2976 (N_2976,N_2154,N_1955);
nand U2977 (N_2977,N_1686,N_1706);
nor U2978 (N_2978,N_1562,N_1673);
and U2979 (N_2979,N_1939,N_1808);
nand U2980 (N_2980,N_2155,N_2143);
nor U2981 (N_2981,N_1702,N_1679);
and U2982 (N_2982,N_1986,N_2196);
nor U2983 (N_2983,N_2247,N_1947);
nand U2984 (N_2984,N_1654,N_1871);
or U2985 (N_2985,N_1669,N_1924);
nand U2986 (N_2986,N_1653,N_1654);
nand U2987 (N_2987,N_1856,N_1563);
and U2988 (N_2988,N_1627,N_1993);
or U2989 (N_2989,N_1679,N_1789);
or U2990 (N_2990,N_2161,N_1959);
nor U2991 (N_2991,N_2177,N_1802);
or U2992 (N_2992,N_1763,N_2225);
nand U2993 (N_2993,N_1765,N_1599);
or U2994 (N_2994,N_1740,N_2076);
and U2995 (N_2995,N_2147,N_1796);
nor U2996 (N_2996,N_2186,N_1703);
nor U2997 (N_2997,N_2081,N_1829);
nand U2998 (N_2998,N_1634,N_2138);
nand U2999 (N_2999,N_1749,N_1639);
nand UO_0 (O_0,N_2489,N_2958);
or UO_1 (O_1,N_2721,N_2401);
nand UO_2 (O_2,N_2473,N_2698);
or UO_3 (O_3,N_2281,N_2765);
nand UO_4 (O_4,N_2703,N_2335);
nor UO_5 (O_5,N_2614,N_2324);
or UO_6 (O_6,N_2944,N_2325);
and UO_7 (O_7,N_2546,N_2708);
and UO_8 (O_8,N_2596,N_2718);
or UO_9 (O_9,N_2522,N_2342);
xnor UO_10 (O_10,N_2599,N_2410);
nand UO_11 (O_11,N_2628,N_2555);
and UO_12 (O_12,N_2658,N_2274);
nor UO_13 (O_13,N_2682,N_2880);
or UO_14 (O_14,N_2809,N_2982);
or UO_15 (O_15,N_2971,N_2746);
or UO_16 (O_16,N_2615,N_2589);
or UO_17 (O_17,N_2283,N_2304);
and UO_18 (O_18,N_2623,N_2362);
nor UO_19 (O_19,N_2271,N_2756);
or UO_20 (O_20,N_2414,N_2578);
and UO_21 (O_21,N_2521,N_2326);
nor UO_22 (O_22,N_2752,N_2920);
nor UO_23 (O_23,N_2977,N_2520);
nand UO_24 (O_24,N_2277,N_2357);
or UO_25 (O_25,N_2939,N_2498);
or UO_26 (O_26,N_2418,N_2445);
nor UO_27 (O_27,N_2833,N_2874);
or UO_28 (O_28,N_2691,N_2426);
nor UO_29 (O_29,N_2406,N_2978);
nand UO_30 (O_30,N_2784,N_2303);
or UO_31 (O_31,N_2593,N_2581);
and UO_32 (O_32,N_2812,N_2926);
nor UO_33 (O_33,N_2517,N_2655);
and UO_34 (O_34,N_2495,N_2567);
xor UO_35 (O_35,N_2803,N_2781);
or UO_36 (O_36,N_2536,N_2435);
nor UO_37 (O_37,N_2523,N_2815);
or UO_38 (O_38,N_2910,N_2339);
and UO_39 (O_39,N_2308,N_2545);
or UO_40 (O_40,N_2286,N_2363);
and UO_41 (O_41,N_2798,N_2398);
nor UO_42 (O_42,N_2644,N_2710);
nor UO_43 (O_43,N_2707,N_2772);
nand UO_44 (O_44,N_2918,N_2715);
and UO_45 (O_45,N_2687,N_2816);
nand UO_46 (O_46,N_2998,N_2341);
and UO_47 (O_47,N_2646,N_2360);
nand UO_48 (O_48,N_2464,N_2935);
nand UO_49 (O_49,N_2257,N_2267);
nand UO_50 (O_50,N_2817,N_2359);
nand UO_51 (O_51,N_2588,N_2417);
nor UO_52 (O_52,N_2288,N_2709);
nand UO_53 (O_53,N_2885,N_2361);
nand UO_54 (O_54,N_2314,N_2569);
nor UO_55 (O_55,N_2748,N_2676);
nor UO_56 (O_56,N_2683,N_2871);
or UO_57 (O_57,N_2662,N_2867);
nand UO_58 (O_58,N_2862,N_2321);
nand UO_59 (O_59,N_2591,N_2810);
nor UO_60 (O_60,N_2639,N_2922);
nand UO_61 (O_61,N_2641,N_2976);
and UO_62 (O_62,N_2776,N_2847);
or UO_63 (O_63,N_2912,N_2309);
and UO_64 (O_64,N_2462,N_2433);
or UO_65 (O_65,N_2537,N_2270);
nor UO_66 (O_66,N_2497,N_2959);
and UO_67 (O_67,N_2893,N_2582);
nand UO_68 (O_68,N_2453,N_2346);
or UO_69 (O_69,N_2843,N_2684);
and UO_70 (O_70,N_2487,N_2524);
nand UO_71 (O_71,N_2492,N_2800);
nand UO_72 (O_72,N_2837,N_2826);
nor UO_73 (O_73,N_2732,N_2506);
nand UO_74 (O_74,N_2407,N_2962);
nor UO_75 (O_75,N_2383,N_2375);
nor UO_76 (O_76,N_2319,N_2884);
nand UO_77 (O_77,N_2377,N_2302);
or UO_78 (O_78,N_2534,N_2671);
or UO_79 (O_79,N_2737,N_2674);
or UO_80 (O_80,N_2617,N_2919);
or UO_81 (O_81,N_2866,N_2702);
nand UO_82 (O_82,N_2825,N_2597);
nand UO_83 (O_83,N_2380,N_2744);
and UO_84 (O_84,N_2908,N_2791);
nor UO_85 (O_85,N_2940,N_2528);
xnor UO_86 (O_86,N_2872,N_2430);
nand UO_87 (O_87,N_2423,N_2350);
nor UO_88 (O_88,N_2475,N_2562);
nor UO_89 (O_89,N_2481,N_2681);
or UO_90 (O_90,N_2619,N_2413);
and UO_91 (O_91,N_2992,N_2356);
nand UO_92 (O_92,N_2425,N_2519);
nor UO_93 (O_93,N_2811,N_2565);
nor UO_94 (O_94,N_2873,N_2889);
and UO_95 (O_95,N_2343,N_2332);
nand UO_96 (O_96,N_2392,N_2879);
and UO_97 (O_97,N_2738,N_2643);
nand UO_98 (O_98,N_2913,N_2938);
and UO_99 (O_99,N_2751,N_2364);
or UO_100 (O_100,N_2848,N_2952);
or UO_101 (O_101,N_2947,N_2807);
nor UO_102 (O_102,N_2793,N_2657);
nor UO_103 (O_103,N_2700,N_2263);
nor UO_104 (O_104,N_2921,N_2906);
or UO_105 (O_105,N_2768,N_2560);
or UO_106 (O_106,N_2750,N_2849);
or UO_107 (O_107,N_2653,N_2486);
or UO_108 (O_108,N_2675,N_2620);
nor UO_109 (O_109,N_2583,N_2666);
and UO_110 (O_110,N_2855,N_2600);
nand UO_111 (O_111,N_2911,N_2526);
nand UO_112 (O_112,N_2282,N_2261);
or UO_113 (O_113,N_2780,N_2693);
nor UO_114 (O_114,N_2496,N_2372);
nor UO_115 (O_115,N_2334,N_2504);
nor UO_116 (O_116,N_2818,N_2386);
nor UO_117 (O_117,N_2931,N_2408);
nor UO_118 (O_118,N_2891,N_2822);
nor UO_119 (O_119,N_2668,N_2654);
nand UO_120 (O_120,N_2353,N_2387);
nor UO_121 (O_121,N_2928,N_2769);
and UO_122 (O_122,N_2877,N_2777);
or UO_123 (O_123,N_2544,N_2859);
nand UO_124 (O_124,N_2667,N_2484);
nand UO_125 (O_125,N_2541,N_2965);
nand UO_126 (O_126,N_2340,N_2695);
and UO_127 (O_127,N_2986,N_2543);
nor UO_128 (O_128,N_2530,N_2411);
nand UO_129 (O_129,N_2923,N_2767);
and UO_130 (O_130,N_2846,N_2835);
nor UO_131 (O_131,N_2568,N_2967);
and UO_132 (O_132,N_2830,N_2990);
and UO_133 (O_133,N_2602,N_2421);
or UO_134 (O_134,N_2858,N_2685);
and UO_135 (O_135,N_2494,N_2905);
nand UO_136 (O_136,N_2397,N_2836);
and UO_137 (O_137,N_2594,N_2951);
or UO_138 (O_138,N_2892,N_2677);
or UO_139 (O_139,N_2839,N_2268);
nand UO_140 (O_140,N_2298,N_2451);
nand UO_141 (O_141,N_2660,N_2604);
and UO_142 (O_142,N_2650,N_2466);
or UO_143 (O_143,N_2757,N_2610);
or UO_144 (O_144,N_2382,N_2250);
nor UO_145 (O_145,N_2525,N_2786);
and UO_146 (O_146,N_2516,N_2424);
or UO_147 (O_147,N_2300,N_2799);
nand UO_148 (O_148,N_2575,N_2801);
nor UO_149 (O_149,N_2554,N_2564);
nor UO_150 (O_150,N_2539,N_2704);
or UO_151 (O_151,N_2624,N_2868);
nor UO_152 (O_152,N_2794,N_2946);
and UO_153 (O_153,N_2642,N_2476);
nand UO_154 (O_154,N_2754,N_2579);
or UO_155 (O_155,N_2284,N_2621);
xor UO_156 (O_156,N_2468,N_2507);
and UO_157 (O_157,N_2860,N_2988);
nor UO_158 (O_158,N_2755,N_2323);
nand UO_159 (O_159,N_2333,N_2804);
nand UO_160 (O_160,N_2348,N_2395);
xnor UO_161 (O_161,N_2483,N_2983);
or UO_162 (O_162,N_2994,N_2774);
or UO_163 (O_163,N_2500,N_2953);
nand UO_164 (O_164,N_2485,N_2638);
xor UO_165 (O_165,N_2742,N_2384);
nand UO_166 (O_166,N_2645,N_2369);
or UO_167 (O_167,N_2311,N_2924);
or UO_168 (O_168,N_2842,N_2743);
nand UO_169 (O_169,N_2491,N_2690);
nor UO_170 (O_170,N_2929,N_2694);
nand UO_171 (O_171,N_2907,N_2779);
nand UO_172 (O_172,N_2457,N_2449);
or UO_173 (O_173,N_2898,N_2775);
nor UO_174 (O_174,N_2735,N_2969);
nor UO_175 (O_175,N_2531,N_2570);
nand UO_176 (O_176,N_2741,N_2312);
nor UO_177 (O_177,N_2618,N_2727);
nor UO_178 (O_178,N_2405,N_2584);
xnor UO_179 (O_179,N_2995,N_2731);
nor UO_180 (O_180,N_2819,N_2396);
nand UO_181 (O_181,N_2699,N_2762);
or UO_182 (O_182,N_2553,N_2854);
nand UO_183 (O_183,N_2882,N_2264);
or UO_184 (O_184,N_2927,N_2814);
nand UO_185 (O_185,N_2412,N_2365);
or UO_186 (O_186,N_2381,N_2328);
nor UO_187 (O_187,N_2393,N_2566);
nor UO_188 (O_188,N_2251,N_2606);
nor UO_189 (O_189,N_2586,N_2488);
nor UO_190 (O_190,N_2469,N_2745);
or UO_191 (O_191,N_2447,N_2881);
or UO_192 (O_192,N_2279,N_2294);
nand UO_193 (O_193,N_2419,N_2499);
or UO_194 (O_194,N_2287,N_2649);
nor UO_195 (O_195,N_2502,N_2438);
and UO_196 (O_196,N_2930,N_2664);
nand UO_197 (O_197,N_2446,N_2612);
nand UO_198 (O_198,N_2637,N_2514);
and UO_199 (O_199,N_2463,N_2672);
nand UO_200 (O_200,N_2552,N_2291);
nand UO_201 (O_201,N_2840,N_2330);
and UO_202 (O_202,N_2626,N_2265);
and UO_203 (O_203,N_2831,N_2749);
and UO_204 (O_204,N_2821,N_2729);
or UO_205 (O_205,N_2436,N_2857);
nand UO_206 (O_206,N_2611,N_2997);
and UO_207 (O_207,N_2422,N_2452);
nand UO_208 (O_208,N_2511,N_2652);
or UO_209 (O_209,N_2409,N_2896);
nor UO_210 (O_210,N_2587,N_2595);
nand UO_211 (O_211,N_2439,N_2787);
and UO_212 (O_212,N_2991,N_2307);
nand UO_213 (O_213,N_2876,N_2764);
nor UO_214 (O_214,N_2945,N_2548);
nand UO_215 (O_215,N_2870,N_2974);
or UO_216 (O_216,N_2431,N_2996);
nand UO_217 (O_217,N_2673,N_2345);
nor UO_218 (O_218,N_2705,N_2761);
nand UO_219 (O_219,N_2442,N_2740);
nor UO_220 (O_220,N_2665,N_2782);
nor UO_221 (O_221,N_2972,N_2573);
nand UO_222 (O_222,N_2925,N_2434);
or UO_223 (O_223,N_2716,N_2585);
xor UO_224 (O_224,N_2322,N_2310);
and UO_225 (O_225,N_2461,N_2909);
nand UO_226 (O_226,N_2355,N_2805);
and UO_227 (O_227,N_2458,N_2917);
nand UO_228 (O_228,N_2973,N_2337);
or UO_229 (O_229,N_2460,N_2459);
or UO_230 (O_230,N_2366,N_2574);
and UO_231 (O_231,N_2295,N_2540);
nand UO_232 (O_232,N_2670,N_2255);
nor UO_233 (O_233,N_2900,N_2465);
nor UO_234 (O_234,N_2932,N_2558);
or UO_235 (O_235,N_2771,N_2622);
or UO_236 (O_236,N_2532,N_2806);
nor UO_237 (O_237,N_2285,N_2914);
nor UO_238 (O_238,N_2580,N_2915);
and UO_239 (O_239,N_2327,N_2313);
and UO_240 (O_240,N_2864,N_2474);
or UO_241 (O_241,N_2747,N_2299);
or UO_242 (O_242,N_2253,N_2680);
nand UO_243 (O_243,N_2933,N_2981);
and UO_244 (O_244,N_2301,N_2420);
or UO_245 (O_245,N_2987,N_2980);
nand UO_246 (O_246,N_2455,N_2989);
or UO_247 (O_247,N_2829,N_2320);
nand UO_248 (O_248,N_2450,N_2934);
nand UO_249 (O_249,N_2367,N_2789);
and UO_250 (O_250,N_2352,N_2961);
nand UO_251 (O_251,N_2571,N_2482);
xor UO_252 (O_252,N_2518,N_2713);
and UO_253 (O_253,N_2427,N_2609);
or UO_254 (O_254,N_2254,N_2441);
or UO_255 (O_255,N_2370,N_2289);
nand UO_256 (O_256,N_2607,N_2902);
nor UO_257 (O_257,N_2975,N_2454);
xor UO_258 (O_258,N_2493,N_2899);
nor UO_259 (O_259,N_2633,N_2338);
and UO_260 (O_260,N_2788,N_2358);
nor UO_261 (O_261,N_2853,N_2968);
and UO_262 (O_262,N_2505,N_2318);
or UO_263 (O_263,N_2634,N_2630);
nand UO_264 (O_264,N_2850,N_2942);
and UO_265 (O_265,N_2440,N_2883);
nor UO_266 (O_266,N_2416,N_2315);
and UO_267 (O_267,N_2717,N_2706);
and UO_268 (O_268,N_2719,N_2785);
nor UO_269 (O_269,N_2904,N_2797);
and UO_270 (O_270,N_2371,N_2444);
or UO_271 (O_271,N_2936,N_2557);
and UO_272 (O_272,N_2470,N_2515);
and UO_273 (O_273,N_2963,N_2888);
xnor UO_274 (O_274,N_2720,N_2613);
and UO_275 (O_275,N_2759,N_2479);
or UO_276 (O_276,N_2865,N_2603);
nand UO_277 (O_277,N_2916,N_2549);
and UO_278 (O_278,N_2559,N_2697);
and UO_279 (O_279,N_2722,N_2273);
or UO_280 (O_280,N_2527,N_2949);
or UO_281 (O_281,N_2394,N_2561);
nand UO_282 (O_282,N_2820,N_2692);
and UO_283 (O_283,N_2467,N_2349);
or UO_284 (O_284,N_2903,N_2448);
and UO_285 (O_285,N_2556,N_2937);
nor UO_286 (O_286,N_2533,N_2472);
xnor UO_287 (O_287,N_2766,N_2725);
nand UO_288 (O_288,N_2875,N_2813);
or UO_289 (O_289,N_2736,N_2950);
nand UO_290 (O_290,N_2262,N_2724);
or UO_291 (O_291,N_2429,N_2258);
and UO_292 (O_292,N_2790,N_2838);
or UO_293 (O_293,N_2266,N_2763);
or UO_294 (O_294,N_2778,N_2391);
xnor UO_295 (O_295,N_2689,N_2783);
nor UO_296 (O_296,N_2688,N_2389);
and UO_297 (O_297,N_2278,N_2714);
nand UO_298 (O_298,N_2632,N_2317);
nand UO_299 (O_299,N_2316,N_2276);
nand UO_300 (O_300,N_2792,N_2869);
or UO_301 (O_301,N_2796,N_2354);
nor UO_302 (O_302,N_2941,N_2576);
or UO_303 (O_303,N_2292,N_2844);
and UO_304 (O_304,N_2999,N_2629);
and UO_305 (O_305,N_2415,N_2828);
xnor UO_306 (O_306,N_2723,N_2378);
nor UO_307 (O_307,N_2547,N_2897);
nor UO_308 (O_308,N_2598,N_2669);
nand UO_309 (O_309,N_2402,N_2385);
nor UO_310 (O_310,N_2739,N_2651);
nor UO_311 (O_311,N_2404,N_2538);
or UO_312 (O_312,N_2960,N_2648);
nand UO_313 (O_313,N_2605,N_2635);
nand UO_314 (O_314,N_2252,N_2726);
and UO_315 (O_315,N_2970,N_2368);
nand UO_316 (O_316,N_2512,N_2728);
or UO_317 (O_317,N_2390,N_2376);
nor UO_318 (O_318,N_2509,N_2955);
and UO_319 (O_319,N_2964,N_2845);
and UO_320 (O_320,N_2647,N_2373);
and UO_321 (O_321,N_2656,N_2590);
nor UO_322 (O_322,N_2535,N_2403);
nor UO_323 (O_323,N_2686,N_2616);
nand UO_324 (O_324,N_2878,N_2513);
and UO_325 (O_325,N_2551,N_2795);
and UO_326 (O_326,N_2259,N_2661);
and UO_327 (O_327,N_2957,N_2437);
nor UO_328 (O_328,N_2269,N_2773);
nand UO_329 (O_329,N_2351,N_2374);
xnor UO_330 (O_330,N_2503,N_2956);
nor UO_331 (O_331,N_2490,N_2344);
and UO_332 (O_332,N_2501,N_2636);
nand UO_333 (O_333,N_2802,N_2592);
and UO_334 (O_334,N_2601,N_2443);
or UO_335 (O_335,N_2734,N_2379);
or UO_336 (O_336,N_2471,N_2834);
and UO_337 (O_337,N_2305,N_2823);
nand UO_338 (O_338,N_2895,N_2293);
or UO_339 (O_339,N_2280,N_2400);
nor UO_340 (O_340,N_2510,N_2542);
xnor UO_341 (O_341,N_2272,N_2640);
nor UO_342 (O_342,N_2659,N_2856);
nand UO_343 (O_343,N_2256,N_2678);
nand UO_344 (O_344,N_2890,N_2901);
and UO_345 (O_345,N_2753,N_2478);
nor UO_346 (O_346,N_2943,N_2984);
or UO_347 (O_347,N_2508,N_2477);
xnor UO_348 (O_348,N_2577,N_2712);
or UO_349 (O_349,N_2608,N_2388);
nand UO_350 (O_350,N_2887,N_2832);
or UO_351 (O_351,N_2863,N_2966);
or UO_352 (O_352,N_2572,N_2275);
and UO_353 (O_353,N_2948,N_2824);
or UO_354 (O_354,N_2529,N_2627);
or UO_355 (O_355,N_2730,N_2663);
or UO_356 (O_356,N_2456,N_2758);
or UO_357 (O_357,N_2290,N_2696);
and UO_358 (O_358,N_2399,N_2827);
xor UO_359 (O_359,N_2336,N_2297);
and UO_360 (O_360,N_2886,N_2631);
nor UO_361 (O_361,N_2701,N_2954);
and UO_362 (O_362,N_2331,N_2979);
nor UO_363 (O_363,N_2760,N_2993);
and UO_364 (O_364,N_2480,N_2625);
or UO_365 (O_365,N_2711,N_2841);
or UO_366 (O_366,N_2563,N_2861);
and UO_367 (O_367,N_2985,N_2852);
nor UO_368 (O_368,N_2679,N_2733);
xnor UO_369 (O_369,N_2808,N_2428);
nor UO_370 (O_370,N_2260,N_2347);
and UO_371 (O_371,N_2770,N_2329);
and UO_372 (O_372,N_2894,N_2550);
or UO_373 (O_373,N_2296,N_2432);
and UO_374 (O_374,N_2851,N_2306);
nor UO_375 (O_375,N_2295,N_2890);
nor UO_376 (O_376,N_2460,N_2693);
or UO_377 (O_377,N_2662,N_2331);
nor UO_378 (O_378,N_2900,N_2955);
and UO_379 (O_379,N_2820,N_2578);
and UO_380 (O_380,N_2879,N_2383);
and UO_381 (O_381,N_2301,N_2448);
and UO_382 (O_382,N_2616,N_2715);
nand UO_383 (O_383,N_2925,N_2762);
nor UO_384 (O_384,N_2660,N_2653);
nand UO_385 (O_385,N_2390,N_2375);
nand UO_386 (O_386,N_2528,N_2295);
nand UO_387 (O_387,N_2605,N_2984);
xnor UO_388 (O_388,N_2770,N_2829);
or UO_389 (O_389,N_2882,N_2389);
nor UO_390 (O_390,N_2535,N_2279);
nor UO_391 (O_391,N_2877,N_2562);
or UO_392 (O_392,N_2867,N_2949);
and UO_393 (O_393,N_2745,N_2630);
and UO_394 (O_394,N_2615,N_2261);
nor UO_395 (O_395,N_2391,N_2330);
or UO_396 (O_396,N_2791,N_2742);
and UO_397 (O_397,N_2600,N_2555);
and UO_398 (O_398,N_2479,N_2933);
nand UO_399 (O_399,N_2656,N_2425);
and UO_400 (O_400,N_2922,N_2790);
and UO_401 (O_401,N_2735,N_2272);
and UO_402 (O_402,N_2348,N_2837);
and UO_403 (O_403,N_2514,N_2859);
and UO_404 (O_404,N_2288,N_2815);
nand UO_405 (O_405,N_2962,N_2405);
nor UO_406 (O_406,N_2740,N_2942);
nor UO_407 (O_407,N_2609,N_2915);
nand UO_408 (O_408,N_2991,N_2293);
and UO_409 (O_409,N_2610,N_2839);
and UO_410 (O_410,N_2856,N_2465);
or UO_411 (O_411,N_2778,N_2742);
nor UO_412 (O_412,N_2558,N_2409);
or UO_413 (O_413,N_2706,N_2584);
xnor UO_414 (O_414,N_2400,N_2875);
and UO_415 (O_415,N_2789,N_2312);
nand UO_416 (O_416,N_2766,N_2598);
and UO_417 (O_417,N_2664,N_2561);
or UO_418 (O_418,N_2586,N_2477);
nand UO_419 (O_419,N_2950,N_2323);
nand UO_420 (O_420,N_2805,N_2506);
and UO_421 (O_421,N_2425,N_2579);
nor UO_422 (O_422,N_2376,N_2413);
and UO_423 (O_423,N_2807,N_2579);
nand UO_424 (O_424,N_2920,N_2615);
nor UO_425 (O_425,N_2536,N_2924);
nand UO_426 (O_426,N_2578,N_2705);
nand UO_427 (O_427,N_2440,N_2339);
nor UO_428 (O_428,N_2458,N_2407);
nand UO_429 (O_429,N_2965,N_2696);
or UO_430 (O_430,N_2406,N_2268);
nand UO_431 (O_431,N_2815,N_2484);
and UO_432 (O_432,N_2513,N_2259);
or UO_433 (O_433,N_2669,N_2948);
nand UO_434 (O_434,N_2618,N_2915);
nand UO_435 (O_435,N_2626,N_2996);
nand UO_436 (O_436,N_2556,N_2806);
and UO_437 (O_437,N_2616,N_2376);
and UO_438 (O_438,N_2719,N_2789);
and UO_439 (O_439,N_2748,N_2577);
or UO_440 (O_440,N_2682,N_2667);
nor UO_441 (O_441,N_2649,N_2816);
nor UO_442 (O_442,N_2911,N_2848);
nor UO_443 (O_443,N_2796,N_2770);
nand UO_444 (O_444,N_2782,N_2868);
and UO_445 (O_445,N_2337,N_2571);
nor UO_446 (O_446,N_2403,N_2676);
or UO_447 (O_447,N_2516,N_2647);
and UO_448 (O_448,N_2599,N_2564);
and UO_449 (O_449,N_2622,N_2424);
nor UO_450 (O_450,N_2965,N_2373);
nand UO_451 (O_451,N_2927,N_2953);
or UO_452 (O_452,N_2698,N_2541);
or UO_453 (O_453,N_2425,N_2838);
nand UO_454 (O_454,N_2674,N_2876);
nand UO_455 (O_455,N_2362,N_2581);
or UO_456 (O_456,N_2858,N_2810);
xor UO_457 (O_457,N_2801,N_2309);
or UO_458 (O_458,N_2624,N_2440);
xor UO_459 (O_459,N_2641,N_2712);
or UO_460 (O_460,N_2709,N_2655);
or UO_461 (O_461,N_2312,N_2370);
or UO_462 (O_462,N_2960,N_2598);
or UO_463 (O_463,N_2705,N_2349);
nor UO_464 (O_464,N_2439,N_2742);
nand UO_465 (O_465,N_2776,N_2496);
nor UO_466 (O_466,N_2813,N_2648);
and UO_467 (O_467,N_2469,N_2706);
nand UO_468 (O_468,N_2594,N_2957);
nand UO_469 (O_469,N_2875,N_2976);
nor UO_470 (O_470,N_2456,N_2707);
nor UO_471 (O_471,N_2820,N_2300);
nand UO_472 (O_472,N_2602,N_2374);
or UO_473 (O_473,N_2282,N_2318);
or UO_474 (O_474,N_2909,N_2282);
nand UO_475 (O_475,N_2838,N_2326);
nor UO_476 (O_476,N_2363,N_2537);
or UO_477 (O_477,N_2944,N_2914);
and UO_478 (O_478,N_2275,N_2254);
nand UO_479 (O_479,N_2700,N_2314);
and UO_480 (O_480,N_2970,N_2502);
nand UO_481 (O_481,N_2893,N_2515);
and UO_482 (O_482,N_2638,N_2458);
and UO_483 (O_483,N_2611,N_2987);
and UO_484 (O_484,N_2625,N_2519);
xnor UO_485 (O_485,N_2582,N_2379);
and UO_486 (O_486,N_2408,N_2676);
and UO_487 (O_487,N_2337,N_2286);
or UO_488 (O_488,N_2356,N_2458);
or UO_489 (O_489,N_2874,N_2306);
nand UO_490 (O_490,N_2380,N_2474);
or UO_491 (O_491,N_2837,N_2911);
and UO_492 (O_492,N_2639,N_2293);
or UO_493 (O_493,N_2490,N_2503);
or UO_494 (O_494,N_2768,N_2821);
nand UO_495 (O_495,N_2700,N_2376);
nor UO_496 (O_496,N_2282,N_2323);
nor UO_497 (O_497,N_2636,N_2520);
and UO_498 (O_498,N_2811,N_2749);
or UO_499 (O_499,N_2455,N_2502);
endmodule