module basic_500_3000_500_5_levels_2xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_439,In_358);
nor U1 (N_1,In_264,In_82);
or U2 (N_2,In_157,In_146);
nor U3 (N_3,In_5,In_407);
and U4 (N_4,In_245,In_239);
nand U5 (N_5,In_479,In_491);
nand U6 (N_6,In_111,In_107);
and U7 (N_7,In_202,In_267);
nor U8 (N_8,In_343,In_213);
nand U9 (N_9,In_97,In_122);
or U10 (N_10,In_277,In_387);
nor U11 (N_11,In_65,In_52);
nor U12 (N_12,In_105,In_353);
nand U13 (N_13,In_257,In_70);
nand U14 (N_14,In_204,In_216);
nand U15 (N_15,In_117,In_238);
nand U16 (N_16,In_258,In_31);
nand U17 (N_17,In_294,In_241);
and U18 (N_18,In_20,In_76);
nor U19 (N_19,In_135,In_64);
nand U20 (N_20,In_271,In_73);
and U21 (N_21,In_465,In_498);
nor U22 (N_22,In_136,In_433);
nor U23 (N_23,In_276,In_410);
nand U24 (N_24,In_392,In_50);
nor U25 (N_25,In_172,In_487);
nor U26 (N_26,In_337,In_299);
nand U27 (N_27,In_349,In_366);
or U28 (N_28,In_452,In_481);
nor U29 (N_29,In_362,In_103);
or U30 (N_30,In_368,In_468);
and U31 (N_31,In_333,In_104);
or U32 (N_32,In_119,In_340);
and U33 (N_33,In_28,In_6);
xnor U34 (N_34,In_401,In_39);
nand U35 (N_35,In_134,In_373);
nand U36 (N_36,In_77,In_272);
nand U37 (N_37,In_228,In_15);
nor U38 (N_38,In_389,In_398);
nand U39 (N_39,In_280,In_57);
and U40 (N_40,In_23,In_339);
and U41 (N_41,In_139,In_397);
nand U42 (N_42,In_209,In_173);
and U43 (N_43,In_35,In_447);
nand U44 (N_44,In_208,In_260);
nor U45 (N_45,In_315,In_462);
and U46 (N_46,In_273,In_59);
nand U47 (N_47,In_244,In_129);
and U48 (N_48,In_307,In_250);
and U49 (N_49,In_155,In_409);
or U50 (N_50,In_482,In_331);
nor U51 (N_51,In_302,In_259);
nand U52 (N_52,In_484,In_475);
nor U53 (N_53,In_150,In_198);
or U54 (N_54,In_360,In_25);
nand U55 (N_55,In_201,In_89);
nor U56 (N_56,In_143,In_14);
nand U57 (N_57,In_435,In_472);
and U58 (N_58,In_378,In_247);
or U59 (N_59,In_224,In_171);
nand U60 (N_60,In_66,In_131);
nand U61 (N_61,In_464,In_287);
and U62 (N_62,In_499,In_170);
xnor U63 (N_63,In_188,In_372);
nor U64 (N_64,In_110,In_399);
and U65 (N_65,In_185,In_81);
nor U66 (N_66,In_376,In_120);
nand U67 (N_67,In_69,In_470);
xnor U68 (N_68,In_268,In_488);
and U69 (N_69,In_453,In_182);
or U70 (N_70,In_256,In_304);
nand U71 (N_71,In_497,In_434);
nand U72 (N_72,In_218,In_12);
and U73 (N_73,In_412,In_48);
nor U74 (N_74,In_288,In_438);
nor U75 (N_75,In_379,In_269);
or U76 (N_76,In_251,In_400);
or U77 (N_77,In_467,In_477);
or U78 (N_78,In_441,In_444);
nand U79 (N_79,In_180,In_92);
or U80 (N_80,In_335,In_310);
nand U81 (N_81,In_386,In_419);
nand U82 (N_82,In_289,In_231);
nor U83 (N_83,In_496,In_169);
or U84 (N_84,In_388,In_174);
nand U85 (N_85,In_83,In_390);
and U86 (N_86,In_297,In_320);
or U87 (N_87,In_214,In_430);
or U88 (N_88,In_316,In_300);
and U89 (N_89,In_324,In_79);
and U90 (N_90,In_164,In_363);
nand U91 (N_91,In_413,In_232);
nand U92 (N_92,In_383,In_474);
or U93 (N_93,In_88,In_437);
and U94 (N_94,In_246,In_355);
nor U95 (N_95,In_163,In_417);
nand U96 (N_96,In_184,In_217);
nor U97 (N_97,In_203,In_255);
or U98 (N_98,In_91,In_40);
or U99 (N_99,In_42,In_114);
or U100 (N_100,In_27,In_22);
or U101 (N_101,In_321,In_431);
nand U102 (N_102,In_425,In_330);
nor U103 (N_103,In_151,In_305);
or U104 (N_104,In_235,In_221);
nor U105 (N_105,In_243,In_408);
and U106 (N_106,In_4,In_93);
or U107 (N_107,In_313,In_406);
and U108 (N_108,In_286,In_443);
or U109 (N_109,In_440,In_147);
nor U110 (N_110,In_87,In_108);
or U111 (N_111,In_225,In_402);
nor U112 (N_112,In_58,In_274);
nand U113 (N_113,In_153,In_265);
nor U114 (N_114,In_176,In_261);
nand U115 (N_115,In_455,In_160);
xor U116 (N_116,In_123,In_415);
or U117 (N_117,In_148,In_370);
and U118 (N_118,In_486,In_240);
and U119 (N_119,In_140,In_292);
or U120 (N_120,In_98,In_47);
or U121 (N_121,In_351,In_219);
nor U122 (N_122,In_442,In_347);
and U123 (N_123,In_327,In_112);
nand U124 (N_124,In_37,In_154);
or U125 (N_125,In_223,In_54);
or U126 (N_126,In_466,In_254);
nor U127 (N_127,In_190,In_473);
nand U128 (N_128,In_449,In_86);
nor U129 (N_129,In_211,In_63);
nor U130 (N_130,In_451,In_385);
nand U131 (N_131,In_314,In_226);
nand U132 (N_132,In_428,In_359);
or U133 (N_133,In_281,In_55);
nand U134 (N_134,In_301,In_306);
and U135 (N_135,In_44,In_90);
and U136 (N_136,In_200,In_236);
or U137 (N_137,In_233,In_16);
nor U138 (N_138,In_51,In_168);
nor U139 (N_139,In_361,In_195);
nand U140 (N_140,In_283,In_458);
nand U141 (N_141,In_7,In_354);
and U142 (N_142,In_404,In_423);
nand U143 (N_143,In_18,In_291);
or U144 (N_144,In_38,In_253);
or U145 (N_145,In_74,In_448);
and U146 (N_146,In_95,In_471);
nor U147 (N_147,In_152,In_341);
or U148 (N_148,In_290,In_285);
and U149 (N_149,In_100,In_414);
or U150 (N_150,In_179,In_344);
or U151 (N_151,In_326,In_445);
nand U152 (N_152,In_374,In_49);
or U153 (N_153,In_84,In_45);
nor U154 (N_154,In_421,In_193);
and U155 (N_155,In_207,In_365);
nor U156 (N_156,In_395,In_94);
nor U157 (N_157,In_127,In_29);
and U158 (N_158,In_113,In_75);
nand U159 (N_159,In_132,In_19);
nor U160 (N_160,In_189,In_270);
or U161 (N_161,In_165,In_336);
nand U162 (N_162,In_295,In_312);
and U163 (N_163,In_234,In_405);
nand U164 (N_164,In_426,In_192);
nand U165 (N_165,In_311,In_394);
or U166 (N_166,In_275,In_191);
nand U167 (N_167,In_391,In_137);
nor U168 (N_168,In_121,In_62);
or U169 (N_169,In_215,In_242);
nand U170 (N_170,In_125,In_375);
nand U171 (N_171,In_115,In_10);
or U172 (N_172,In_266,In_317);
and U173 (N_173,In_205,In_41);
nand U174 (N_174,In_116,In_357);
or U175 (N_175,In_175,In_124);
and U176 (N_176,In_356,In_308);
nand U177 (N_177,In_494,In_328);
nand U178 (N_178,In_377,In_43);
and U179 (N_179,In_478,In_24);
or U180 (N_180,In_282,In_446);
and U181 (N_181,In_485,In_342);
and U182 (N_182,In_323,In_220);
nand U183 (N_183,In_495,In_322);
xnor U184 (N_184,In_106,In_346);
and U185 (N_185,In_476,In_126);
nor U186 (N_186,In_483,In_457);
and U187 (N_187,In_145,In_30);
nor U188 (N_188,In_68,In_167);
and U189 (N_189,In_460,In_162);
nor U190 (N_190,In_133,In_101);
or U191 (N_191,In_102,In_416);
nand U192 (N_192,In_138,In_206);
and U193 (N_193,In_293,In_364);
or U194 (N_194,In_11,In_210);
nor U195 (N_195,In_469,In_325);
nand U196 (N_196,In_178,In_329);
nand U197 (N_197,In_450,In_85);
xor U198 (N_198,In_384,In_393);
nand U199 (N_199,In_380,In_298);
nand U200 (N_200,In_262,In_53);
nor U201 (N_201,In_493,In_263);
nor U202 (N_202,In_338,In_348);
nor U203 (N_203,In_489,In_17);
or U204 (N_204,In_9,In_0);
or U205 (N_205,In_99,In_199);
xor U206 (N_206,In_166,In_403);
nor U207 (N_207,In_454,In_352);
nor U208 (N_208,In_429,In_80);
and U209 (N_209,In_420,In_427);
nor U210 (N_210,In_141,In_480);
xnor U211 (N_211,In_248,In_72);
or U212 (N_212,In_303,In_418);
and U213 (N_213,In_144,In_332);
or U214 (N_214,In_33,In_46);
nand U215 (N_215,In_34,In_186);
and U216 (N_216,In_26,In_60);
nand U217 (N_217,In_230,In_284);
nor U218 (N_218,In_350,In_296);
nor U219 (N_219,In_411,In_396);
nand U220 (N_220,In_183,In_227);
xnor U221 (N_221,In_156,In_56);
or U222 (N_222,In_158,In_422);
nor U223 (N_223,In_130,In_278);
nor U224 (N_224,In_71,In_279);
nor U225 (N_225,In_367,In_432);
and U226 (N_226,In_61,In_369);
nor U227 (N_227,In_249,In_461);
nor U228 (N_228,In_2,In_318);
and U229 (N_229,In_3,In_381);
or U230 (N_230,In_212,In_109);
nand U231 (N_231,In_118,In_345);
and U232 (N_232,In_78,In_319);
and U233 (N_233,In_334,In_187);
and U234 (N_234,In_229,In_456);
and U235 (N_235,In_222,In_459);
nand U236 (N_236,In_436,In_194);
or U237 (N_237,In_196,In_36);
and U238 (N_238,In_177,In_309);
nor U239 (N_239,In_159,In_96);
or U240 (N_240,In_197,In_8);
nand U241 (N_241,In_490,In_128);
nor U242 (N_242,In_181,In_142);
nand U243 (N_243,In_1,In_252);
nand U244 (N_244,In_21,In_371);
and U245 (N_245,In_463,In_13);
and U246 (N_246,In_237,In_149);
or U247 (N_247,In_161,In_32);
or U248 (N_248,In_424,In_67);
and U249 (N_249,In_492,In_382);
and U250 (N_250,In_45,In_43);
xnor U251 (N_251,In_293,In_350);
or U252 (N_252,In_483,In_397);
or U253 (N_253,In_124,In_95);
and U254 (N_254,In_396,In_162);
nand U255 (N_255,In_138,In_238);
nand U256 (N_256,In_177,In_308);
nand U257 (N_257,In_67,In_299);
nand U258 (N_258,In_53,In_496);
and U259 (N_259,In_391,In_261);
or U260 (N_260,In_69,In_119);
nand U261 (N_261,In_387,In_369);
or U262 (N_262,In_117,In_396);
nor U263 (N_263,In_407,In_38);
or U264 (N_264,In_248,In_488);
or U265 (N_265,In_162,In_133);
and U266 (N_266,In_313,In_413);
and U267 (N_267,In_90,In_195);
nor U268 (N_268,In_204,In_438);
and U269 (N_269,In_457,In_312);
nand U270 (N_270,In_14,In_273);
nand U271 (N_271,In_389,In_104);
or U272 (N_272,In_149,In_83);
nor U273 (N_273,In_49,In_337);
or U274 (N_274,In_286,In_118);
or U275 (N_275,In_337,In_379);
and U276 (N_276,In_214,In_240);
nor U277 (N_277,In_470,In_292);
or U278 (N_278,In_231,In_122);
nor U279 (N_279,In_360,In_480);
nand U280 (N_280,In_175,In_443);
nor U281 (N_281,In_193,In_393);
or U282 (N_282,In_392,In_300);
and U283 (N_283,In_423,In_372);
or U284 (N_284,In_372,In_324);
and U285 (N_285,In_191,In_236);
and U286 (N_286,In_469,In_372);
nand U287 (N_287,In_287,In_373);
xnor U288 (N_288,In_488,In_270);
nor U289 (N_289,In_114,In_254);
nor U290 (N_290,In_369,In_408);
nand U291 (N_291,In_133,In_11);
nor U292 (N_292,In_79,In_357);
nor U293 (N_293,In_483,In_208);
nor U294 (N_294,In_385,In_152);
and U295 (N_295,In_18,In_307);
nand U296 (N_296,In_57,In_31);
and U297 (N_297,In_345,In_141);
or U298 (N_298,In_477,In_384);
nor U299 (N_299,In_64,In_384);
nand U300 (N_300,In_102,In_9);
or U301 (N_301,In_177,In_361);
or U302 (N_302,In_120,In_115);
nor U303 (N_303,In_353,In_22);
nand U304 (N_304,In_50,In_448);
and U305 (N_305,In_63,In_302);
nor U306 (N_306,In_98,In_498);
and U307 (N_307,In_221,In_491);
nor U308 (N_308,In_344,In_230);
nor U309 (N_309,In_437,In_476);
or U310 (N_310,In_148,In_28);
nor U311 (N_311,In_100,In_143);
and U312 (N_312,In_344,In_177);
and U313 (N_313,In_16,In_186);
nor U314 (N_314,In_150,In_25);
nand U315 (N_315,In_262,In_77);
nor U316 (N_316,In_83,In_433);
and U317 (N_317,In_470,In_171);
or U318 (N_318,In_292,In_485);
nor U319 (N_319,In_12,In_154);
nand U320 (N_320,In_471,In_363);
nand U321 (N_321,In_264,In_456);
nor U322 (N_322,In_460,In_340);
nor U323 (N_323,In_72,In_348);
and U324 (N_324,In_86,In_215);
nand U325 (N_325,In_435,In_457);
and U326 (N_326,In_226,In_18);
and U327 (N_327,In_307,In_30);
nand U328 (N_328,In_23,In_336);
or U329 (N_329,In_392,In_170);
or U330 (N_330,In_98,In_108);
nor U331 (N_331,In_442,In_127);
and U332 (N_332,In_399,In_266);
nor U333 (N_333,In_416,In_192);
and U334 (N_334,In_423,In_448);
or U335 (N_335,In_413,In_295);
nand U336 (N_336,In_198,In_39);
and U337 (N_337,In_272,In_389);
and U338 (N_338,In_343,In_107);
nand U339 (N_339,In_110,In_451);
nand U340 (N_340,In_156,In_230);
and U341 (N_341,In_294,In_96);
nand U342 (N_342,In_304,In_23);
nor U343 (N_343,In_227,In_140);
or U344 (N_344,In_459,In_342);
and U345 (N_345,In_131,In_173);
nand U346 (N_346,In_15,In_282);
nand U347 (N_347,In_1,In_65);
and U348 (N_348,In_303,In_221);
or U349 (N_349,In_476,In_155);
nor U350 (N_350,In_27,In_412);
nand U351 (N_351,In_448,In_455);
or U352 (N_352,In_395,In_70);
or U353 (N_353,In_440,In_373);
and U354 (N_354,In_275,In_224);
or U355 (N_355,In_217,In_174);
and U356 (N_356,In_16,In_187);
nand U357 (N_357,In_339,In_5);
nor U358 (N_358,In_187,In_244);
nand U359 (N_359,In_476,In_221);
nor U360 (N_360,In_257,In_90);
xnor U361 (N_361,In_248,In_430);
nand U362 (N_362,In_301,In_464);
or U363 (N_363,In_230,In_38);
or U364 (N_364,In_215,In_266);
nor U365 (N_365,In_466,In_467);
nor U366 (N_366,In_327,In_20);
and U367 (N_367,In_262,In_320);
and U368 (N_368,In_136,In_439);
and U369 (N_369,In_285,In_405);
nand U370 (N_370,In_300,In_294);
nor U371 (N_371,In_419,In_152);
nor U372 (N_372,In_83,In_247);
or U373 (N_373,In_122,In_317);
nor U374 (N_374,In_85,In_87);
nor U375 (N_375,In_375,In_58);
and U376 (N_376,In_492,In_295);
or U377 (N_377,In_246,In_88);
or U378 (N_378,In_244,In_156);
nor U379 (N_379,In_359,In_403);
nand U380 (N_380,In_450,In_223);
nand U381 (N_381,In_51,In_490);
nand U382 (N_382,In_363,In_62);
and U383 (N_383,In_245,In_165);
nor U384 (N_384,In_21,In_334);
nand U385 (N_385,In_20,In_245);
nor U386 (N_386,In_191,In_145);
nor U387 (N_387,In_216,In_489);
nand U388 (N_388,In_352,In_156);
or U389 (N_389,In_217,In_1);
or U390 (N_390,In_449,In_198);
nor U391 (N_391,In_372,In_489);
nand U392 (N_392,In_459,In_228);
and U393 (N_393,In_469,In_50);
nor U394 (N_394,In_115,In_489);
and U395 (N_395,In_51,In_375);
nand U396 (N_396,In_206,In_279);
nand U397 (N_397,In_468,In_262);
nand U398 (N_398,In_495,In_198);
or U399 (N_399,In_463,In_245);
and U400 (N_400,In_158,In_434);
nor U401 (N_401,In_396,In_202);
and U402 (N_402,In_489,In_424);
nor U403 (N_403,In_20,In_381);
nor U404 (N_404,In_485,In_311);
and U405 (N_405,In_188,In_368);
nor U406 (N_406,In_145,In_483);
nand U407 (N_407,In_364,In_110);
nand U408 (N_408,In_457,In_308);
and U409 (N_409,In_222,In_225);
xnor U410 (N_410,In_251,In_278);
or U411 (N_411,In_369,In_56);
or U412 (N_412,In_113,In_81);
nand U413 (N_413,In_384,In_337);
or U414 (N_414,In_372,In_211);
or U415 (N_415,In_494,In_429);
nand U416 (N_416,In_425,In_470);
and U417 (N_417,In_308,In_400);
nor U418 (N_418,In_284,In_79);
nor U419 (N_419,In_39,In_104);
nand U420 (N_420,In_430,In_484);
or U421 (N_421,In_381,In_433);
or U422 (N_422,In_102,In_255);
nor U423 (N_423,In_62,In_236);
and U424 (N_424,In_332,In_384);
nand U425 (N_425,In_373,In_69);
or U426 (N_426,In_190,In_160);
nand U427 (N_427,In_53,In_21);
nor U428 (N_428,In_380,In_299);
or U429 (N_429,In_116,In_133);
and U430 (N_430,In_15,In_206);
nand U431 (N_431,In_432,In_471);
nand U432 (N_432,In_294,In_414);
or U433 (N_433,In_60,In_478);
nand U434 (N_434,In_267,In_439);
nor U435 (N_435,In_305,In_274);
and U436 (N_436,In_56,In_364);
nor U437 (N_437,In_373,In_90);
nand U438 (N_438,In_188,In_41);
and U439 (N_439,In_364,In_92);
or U440 (N_440,In_296,In_226);
or U441 (N_441,In_75,In_356);
or U442 (N_442,In_186,In_115);
or U443 (N_443,In_499,In_172);
nand U444 (N_444,In_70,In_254);
and U445 (N_445,In_86,In_95);
or U446 (N_446,In_8,In_157);
or U447 (N_447,In_225,In_308);
and U448 (N_448,In_138,In_181);
nand U449 (N_449,In_395,In_98);
or U450 (N_450,In_484,In_22);
nand U451 (N_451,In_7,In_270);
nor U452 (N_452,In_282,In_131);
nor U453 (N_453,In_325,In_370);
nor U454 (N_454,In_129,In_495);
and U455 (N_455,In_451,In_292);
or U456 (N_456,In_99,In_329);
or U457 (N_457,In_68,In_381);
or U458 (N_458,In_16,In_324);
nor U459 (N_459,In_248,In_329);
and U460 (N_460,In_291,In_85);
and U461 (N_461,In_198,In_342);
or U462 (N_462,In_202,In_181);
nor U463 (N_463,In_128,In_344);
and U464 (N_464,In_42,In_453);
nand U465 (N_465,In_45,In_363);
and U466 (N_466,In_79,In_214);
nand U467 (N_467,In_52,In_157);
or U468 (N_468,In_169,In_457);
nor U469 (N_469,In_418,In_49);
and U470 (N_470,In_280,In_101);
or U471 (N_471,In_439,In_220);
and U472 (N_472,In_17,In_285);
nand U473 (N_473,In_195,In_237);
nand U474 (N_474,In_13,In_41);
or U475 (N_475,In_255,In_185);
and U476 (N_476,In_374,In_12);
and U477 (N_477,In_266,In_263);
and U478 (N_478,In_433,In_305);
and U479 (N_479,In_44,In_37);
and U480 (N_480,In_68,In_146);
and U481 (N_481,In_284,In_150);
or U482 (N_482,In_150,In_481);
nor U483 (N_483,In_195,In_95);
xor U484 (N_484,In_321,In_355);
nor U485 (N_485,In_69,In_420);
nor U486 (N_486,In_391,In_237);
xnor U487 (N_487,In_228,In_440);
nor U488 (N_488,In_332,In_245);
and U489 (N_489,In_468,In_444);
or U490 (N_490,In_406,In_133);
xnor U491 (N_491,In_177,In_171);
nor U492 (N_492,In_247,In_494);
nor U493 (N_493,In_240,In_12);
nand U494 (N_494,In_113,In_388);
nand U495 (N_495,In_113,In_427);
nor U496 (N_496,In_172,In_275);
nand U497 (N_497,In_288,In_39);
nor U498 (N_498,In_488,In_244);
nand U499 (N_499,In_217,In_233);
or U500 (N_500,In_271,In_9);
and U501 (N_501,In_309,In_23);
nor U502 (N_502,In_285,In_488);
or U503 (N_503,In_223,In_309);
nor U504 (N_504,In_223,In_478);
nor U505 (N_505,In_371,In_252);
nand U506 (N_506,In_439,In_324);
or U507 (N_507,In_414,In_149);
and U508 (N_508,In_1,In_277);
xor U509 (N_509,In_165,In_122);
nand U510 (N_510,In_249,In_163);
xor U511 (N_511,In_316,In_101);
nand U512 (N_512,In_194,In_485);
nor U513 (N_513,In_71,In_114);
or U514 (N_514,In_450,In_412);
or U515 (N_515,In_156,In_499);
and U516 (N_516,In_80,In_335);
or U517 (N_517,In_206,In_57);
or U518 (N_518,In_198,In_2);
and U519 (N_519,In_464,In_40);
nand U520 (N_520,In_429,In_364);
xor U521 (N_521,In_263,In_343);
and U522 (N_522,In_127,In_23);
nor U523 (N_523,In_354,In_341);
or U524 (N_524,In_301,In_99);
or U525 (N_525,In_252,In_56);
and U526 (N_526,In_382,In_417);
and U527 (N_527,In_331,In_243);
or U528 (N_528,In_204,In_295);
nand U529 (N_529,In_467,In_453);
or U530 (N_530,In_253,In_174);
nor U531 (N_531,In_3,In_472);
and U532 (N_532,In_18,In_46);
nand U533 (N_533,In_347,In_354);
nand U534 (N_534,In_212,In_282);
nor U535 (N_535,In_215,In_411);
or U536 (N_536,In_451,In_83);
nor U537 (N_537,In_263,In_355);
nor U538 (N_538,In_309,In_13);
or U539 (N_539,In_361,In_153);
and U540 (N_540,In_322,In_87);
nand U541 (N_541,In_111,In_265);
nor U542 (N_542,In_8,In_249);
and U543 (N_543,In_486,In_349);
nor U544 (N_544,In_490,In_267);
and U545 (N_545,In_314,In_309);
nor U546 (N_546,In_224,In_276);
nor U547 (N_547,In_106,In_25);
or U548 (N_548,In_200,In_355);
nand U549 (N_549,In_292,In_369);
and U550 (N_550,In_127,In_465);
nor U551 (N_551,In_122,In_57);
and U552 (N_552,In_317,In_117);
nor U553 (N_553,In_306,In_181);
or U554 (N_554,In_235,In_83);
nor U555 (N_555,In_256,In_338);
or U556 (N_556,In_83,In_283);
or U557 (N_557,In_492,In_404);
nand U558 (N_558,In_422,In_234);
and U559 (N_559,In_370,In_200);
or U560 (N_560,In_301,In_59);
nor U561 (N_561,In_46,In_14);
or U562 (N_562,In_384,In_78);
or U563 (N_563,In_210,In_289);
or U564 (N_564,In_80,In_445);
xnor U565 (N_565,In_397,In_180);
nand U566 (N_566,In_399,In_75);
and U567 (N_567,In_110,In_402);
or U568 (N_568,In_432,In_90);
or U569 (N_569,In_81,In_312);
nor U570 (N_570,In_197,In_252);
or U571 (N_571,In_365,In_47);
nand U572 (N_572,In_479,In_478);
nand U573 (N_573,In_194,In_33);
nand U574 (N_574,In_396,In_122);
nand U575 (N_575,In_489,In_458);
nand U576 (N_576,In_6,In_495);
nor U577 (N_577,In_214,In_481);
nor U578 (N_578,In_2,In_272);
or U579 (N_579,In_164,In_419);
nor U580 (N_580,In_133,In_50);
and U581 (N_581,In_86,In_92);
and U582 (N_582,In_397,In_316);
nor U583 (N_583,In_414,In_19);
nand U584 (N_584,In_36,In_141);
or U585 (N_585,In_321,In_499);
nand U586 (N_586,In_31,In_488);
nand U587 (N_587,In_409,In_458);
or U588 (N_588,In_122,In_309);
and U589 (N_589,In_498,In_316);
or U590 (N_590,In_421,In_288);
or U591 (N_591,In_76,In_361);
nand U592 (N_592,In_470,In_323);
or U593 (N_593,In_361,In_128);
nand U594 (N_594,In_137,In_187);
nor U595 (N_595,In_108,In_46);
nor U596 (N_596,In_197,In_362);
or U597 (N_597,In_21,In_332);
nand U598 (N_598,In_4,In_19);
nand U599 (N_599,In_278,In_168);
nand U600 (N_600,N_235,N_481);
or U601 (N_601,N_139,N_156);
nor U602 (N_602,N_464,N_459);
nand U603 (N_603,N_405,N_133);
and U604 (N_604,N_421,N_579);
or U605 (N_605,N_445,N_348);
and U606 (N_606,N_287,N_595);
and U607 (N_607,N_490,N_24);
nand U608 (N_608,N_57,N_442);
or U609 (N_609,N_425,N_402);
nand U610 (N_610,N_565,N_246);
xor U611 (N_611,N_503,N_341);
nand U612 (N_612,N_477,N_154);
and U613 (N_613,N_377,N_232);
xnor U614 (N_614,N_489,N_31);
and U615 (N_615,N_573,N_280);
or U616 (N_616,N_22,N_126);
nor U617 (N_617,N_479,N_282);
nand U618 (N_618,N_275,N_568);
and U619 (N_619,N_279,N_572);
nor U620 (N_620,N_149,N_314);
nor U621 (N_621,N_333,N_100);
and U622 (N_622,N_85,N_376);
or U623 (N_623,N_83,N_276);
or U624 (N_624,N_73,N_457);
nor U625 (N_625,N_122,N_75);
and U626 (N_626,N_550,N_35);
nor U627 (N_627,N_244,N_438);
and U628 (N_628,N_182,N_391);
nor U629 (N_629,N_554,N_32);
and U630 (N_630,N_549,N_253);
and U631 (N_631,N_51,N_309);
or U632 (N_632,N_157,N_559);
or U633 (N_633,N_423,N_251);
or U634 (N_634,N_177,N_527);
nand U635 (N_635,N_44,N_195);
nor U636 (N_636,N_353,N_240);
and U637 (N_637,N_140,N_321);
nand U638 (N_638,N_8,N_62);
nor U639 (N_639,N_270,N_265);
xnor U640 (N_640,N_381,N_170);
xor U641 (N_641,N_365,N_238);
or U642 (N_642,N_34,N_216);
nor U643 (N_643,N_493,N_249);
nor U644 (N_644,N_214,N_255);
nor U645 (N_645,N_10,N_413);
or U646 (N_646,N_553,N_98);
and U647 (N_647,N_103,N_460);
or U648 (N_648,N_4,N_307);
and U649 (N_649,N_9,N_525);
nor U650 (N_650,N_99,N_404);
and U651 (N_651,N_124,N_582);
nand U652 (N_652,N_310,N_332);
and U653 (N_653,N_323,N_450);
nor U654 (N_654,N_541,N_84);
and U655 (N_655,N_470,N_248);
nor U656 (N_656,N_151,N_507);
nor U657 (N_657,N_347,N_19);
nor U658 (N_658,N_218,N_302);
nand U659 (N_659,N_271,N_476);
nand U660 (N_660,N_107,N_74);
nand U661 (N_661,N_528,N_315);
nor U662 (N_662,N_494,N_184);
and U663 (N_663,N_327,N_574);
nand U664 (N_664,N_548,N_322);
nand U665 (N_665,N_570,N_48);
or U666 (N_666,N_96,N_209);
or U667 (N_667,N_432,N_12);
and U668 (N_668,N_500,N_65);
nand U669 (N_669,N_546,N_436);
nand U670 (N_670,N_552,N_43);
or U671 (N_671,N_33,N_147);
and U672 (N_672,N_378,N_13);
and U673 (N_673,N_516,N_152);
nand U674 (N_674,N_417,N_364);
or U675 (N_675,N_564,N_418);
nand U676 (N_676,N_491,N_303);
nand U677 (N_677,N_69,N_369);
or U678 (N_678,N_317,N_426);
or U679 (N_679,N_155,N_208);
and U680 (N_680,N_104,N_135);
nand U681 (N_681,N_112,N_586);
nor U682 (N_682,N_430,N_211);
and U683 (N_683,N_173,N_258);
and U684 (N_684,N_351,N_558);
nand U685 (N_685,N_326,N_411);
or U686 (N_686,N_120,N_106);
and U687 (N_687,N_439,N_367);
or U688 (N_688,N_560,N_121);
or U689 (N_689,N_360,N_409);
nand U690 (N_690,N_544,N_210);
nor U691 (N_691,N_483,N_264);
nand U692 (N_692,N_141,N_88);
and U693 (N_693,N_357,N_562);
and U694 (N_694,N_401,N_160);
nor U695 (N_695,N_190,N_262);
nor U696 (N_696,N_215,N_273);
nor U697 (N_697,N_437,N_578);
nor U698 (N_698,N_305,N_537);
and U699 (N_699,N_575,N_66);
nand U700 (N_700,N_545,N_236);
nor U701 (N_701,N_68,N_328);
nand U702 (N_702,N_338,N_174);
nor U703 (N_703,N_520,N_185);
xnor U704 (N_704,N_142,N_523);
nand U705 (N_705,N_186,N_343);
nand U706 (N_706,N_269,N_6);
or U707 (N_707,N_181,N_40);
or U708 (N_708,N_291,N_294);
or U709 (N_709,N_366,N_359);
and U710 (N_710,N_162,N_188);
and U711 (N_711,N_256,N_435);
nor U712 (N_712,N_410,N_311);
nor U713 (N_713,N_101,N_498);
or U714 (N_714,N_342,N_254);
or U715 (N_715,N_385,N_252);
and U716 (N_716,N_592,N_455);
nor U717 (N_717,N_581,N_340);
nand U718 (N_718,N_518,N_580);
nor U719 (N_719,N_495,N_227);
nand U720 (N_720,N_416,N_194);
or U721 (N_721,N_115,N_179);
nand U722 (N_722,N_241,N_199);
or U723 (N_723,N_488,N_233);
nor U724 (N_724,N_150,N_354);
nor U725 (N_725,N_221,N_557);
nor U726 (N_726,N_427,N_250);
or U727 (N_727,N_415,N_433);
and U728 (N_728,N_597,N_260);
or U729 (N_729,N_345,N_148);
or U730 (N_730,N_134,N_136);
and U731 (N_731,N_511,N_596);
nor U732 (N_732,N_113,N_517);
nand U733 (N_733,N_458,N_396);
and U734 (N_734,N_172,N_398);
nand U735 (N_735,N_5,N_577);
nor U736 (N_736,N_226,N_266);
and U737 (N_737,N_29,N_82);
nand U738 (N_738,N_487,N_95);
and U739 (N_739,N_299,N_325);
nand U740 (N_740,N_229,N_526);
or U741 (N_741,N_384,N_506);
or U742 (N_742,N_301,N_144);
xor U743 (N_743,N_16,N_118);
nor U744 (N_744,N_422,N_585);
nand U745 (N_745,N_499,N_175);
nand U746 (N_746,N_129,N_465);
nor U747 (N_747,N_213,N_1);
nor U748 (N_748,N_145,N_349);
nor U749 (N_749,N_382,N_510);
or U750 (N_750,N_454,N_428);
and U751 (N_751,N_368,N_36);
nor U752 (N_752,N_389,N_87);
and U753 (N_753,N_283,N_168);
nor U754 (N_754,N_219,N_370);
xor U755 (N_755,N_539,N_78);
nor U756 (N_756,N_164,N_289);
nor U757 (N_757,N_590,N_335);
or U758 (N_758,N_3,N_566);
nand U759 (N_759,N_452,N_485);
nor U760 (N_760,N_295,N_583);
or U761 (N_761,N_277,N_532);
nand U762 (N_762,N_390,N_166);
or U763 (N_763,N_358,N_480);
and U764 (N_764,N_64,N_478);
nand U765 (N_765,N_50,N_15);
and U766 (N_766,N_203,N_589);
nor U767 (N_767,N_412,N_443);
nor U768 (N_768,N_180,N_361);
and U769 (N_769,N_56,N_80);
nand U770 (N_770,N_469,N_515);
nand U771 (N_771,N_128,N_116);
nand U772 (N_772,N_59,N_290);
and U773 (N_773,N_334,N_37);
and U774 (N_774,N_30,N_400);
or U775 (N_775,N_392,N_547);
nor U776 (N_776,N_593,N_163);
and U777 (N_777,N_191,N_300);
nand U778 (N_778,N_60,N_234);
nor U779 (N_779,N_420,N_153);
nor U780 (N_780,N_339,N_521);
nand U781 (N_781,N_388,N_344);
and U782 (N_782,N_308,N_448);
nand U783 (N_783,N_383,N_200);
or U784 (N_784,N_239,N_441);
or U785 (N_785,N_513,N_535);
nor U786 (N_786,N_569,N_408);
or U787 (N_787,N_293,N_313);
or U788 (N_788,N_542,N_591);
nor U789 (N_789,N_414,N_159);
nor U790 (N_790,N_588,N_486);
or U791 (N_791,N_538,N_571);
or U792 (N_792,N_261,N_286);
nand U793 (N_793,N_449,N_397);
nor U794 (N_794,N_285,N_453);
nand U795 (N_795,N_55,N_504);
or U796 (N_796,N_54,N_529);
and U797 (N_797,N_551,N_161);
nor U798 (N_798,N_108,N_587);
nor U799 (N_799,N_67,N_268);
or U800 (N_800,N_471,N_374);
nand U801 (N_801,N_350,N_519);
nor U802 (N_802,N_501,N_114);
or U803 (N_803,N_187,N_594);
nor U804 (N_804,N_49,N_394);
and U805 (N_805,N_109,N_2);
nor U806 (N_806,N_20,N_380);
or U807 (N_807,N_356,N_93);
or U808 (N_808,N_70,N_89);
nor U809 (N_809,N_482,N_90);
or U810 (N_810,N_23,N_18);
nand U811 (N_811,N_63,N_496);
nor U812 (N_812,N_373,N_131);
and U813 (N_813,N_531,N_77);
nand U814 (N_814,N_312,N_263);
nor U815 (N_815,N_143,N_514);
or U816 (N_816,N_204,N_79);
or U817 (N_817,N_27,N_167);
or U818 (N_818,N_14,N_46);
or U819 (N_819,N_284,N_110);
nor U820 (N_820,N_524,N_138);
nor U821 (N_821,N_201,N_207);
and U822 (N_822,N_505,N_224);
or U823 (N_823,N_297,N_92);
nor U824 (N_824,N_444,N_395);
or U825 (N_825,N_509,N_292);
or U826 (N_826,N_363,N_462);
or U827 (N_827,N_272,N_205);
nor U828 (N_828,N_7,N_28);
nor U829 (N_829,N_362,N_387);
nand U830 (N_830,N_534,N_393);
nand U831 (N_831,N_91,N_336);
or U832 (N_832,N_561,N_26);
or U833 (N_833,N_379,N_97);
or U834 (N_834,N_0,N_267);
nor U835 (N_835,N_352,N_197);
nand U836 (N_836,N_225,N_288);
nor U837 (N_837,N_237,N_212);
nand U838 (N_838,N_223,N_176);
xor U839 (N_839,N_473,N_598);
nand U840 (N_840,N_502,N_316);
xor U841 (N_841,N_466,N_39);
nand U842 (N_842,N_247,N_72);
or U843 (N_843,N_324,N_447);
nor U844 (N_844,N_555,N_512);
or U845 (N_845,N_119,N_47);
and U846 (N_846,N_165,N_576);
and U847 (N_847,N_25,N_375);
and U848 (N_848,N_440,N_543);
and U849 (N_849,N_281,N_472);
and U850 (N_850,N_536,N_61);
and U851 (N_851,N_123,N_178);
or U852 (N_852,N_533,N_403);
nor U853 (N_853,N_296,N_306);
nor U854 (N_854,N_419,N_508);
xnor U855 (N_855,N_446,N_158);
nand U856 (N_856,N_319,N_274);
or U857 (N_857,N_242,N_217);
nor U858 (N_858,N_304,N_130);
nor U859 (N_859,N_228,N_346);
nor U860 (N_860,N_497,N_259);
or U861 (N_861,N_456,N_41);
nand U862 (N_862,N_463,N_222);
or U863 (N_863,N_146,N_53);
and U864 (N_864,N_424,N_245);
nor U865 (N_865,N_243,N_102);
nor U866 (N_866,N_125,N_220);
nand U867 (N_867,N_42,N_105);
or U868 (N_868,N_21,N_337);
or U869 (N_869,N_298,N_434);
or U870 (N_870,N_38,N_198);
and U871 (N_871,N_372,N_257);
and U872 (N_872,N_111,N_371);
nand U873 (N_873,N_386,N_399);
or U874 (N_874,N_17,N_522);
and U875 (N_875,N_563,N_406);
xor U876 (N_876,N_318,N_331);
nand U877 (N_877,N_484,N_206);
or U878 (N_878,N_193,N_599);
or U879 (N_879,N_86,N_183);
and U880 (N_880,N_45,N_530);
or U881 (N_881,N_474,N_71);
and U882 (N_882,N_451,N_584);
nand U883 (N_883,N_330,N_461);
nand U884 (N_884,N_355,N_468);
and U885 (N_885,N_189,N_556);
nand U886 (N_886,N_540,N_202);
nor U887 (N_887,N_429,N_81);
nand U888 (N_888,N_52,N_192);
or U889 (N_889,N_171,N_230);
nand U890 (N_890,N_117,N_137);
and U891 (N_891,N_132,N_567);
nand U892 (N_892,N_407,N_169);
and U893 (N_893,N_231,N_58);
or U894 (N_894,N_467,N_329);
or U895 (N_895,N_431,N_196);
nor U896 (N_896,N_475,N_11);
or U897 (N_897,N_278,N_94);
and U898 (N_898,N_320,N_127);
nand U899 (N_899,N_76,N_492);
nand U900 (N_900,N_154,N_523);
and U901 (N_901,N_253,N_114);
xnor U902 (N_902,N_78,N_58);
nor U903 (N_903,N_230,N_505);
and U904 (N_904,N_250,N_367);
nor U905 (N_905,N_235,N_198);
or U906 (N_906,N_293,N_453);
and U907 (N_907,N_535,N_36);
or U908 (N_908,N_164,N_557);
and U909 (N_909,N_186,N_525);
nand U910 (N_910,N_237,N_146);
nor U911 (N_911,N_521,N_489);
or U912 (N_912,N_530,N_220);
and U913 (N_913,N_426,N_60);
nor U914 (N_914,N_586,N_271);
or U915 (N_915,N_140,N_483);
and U916 (N_916,N_562,N_46);
and U917 (N_917,N_458,N_78);
or U918 (N_918,N_311,N_488);
or U919 (N_919,N_77,N_517);
or U920 (N_920,N_266,N_509);
nor U921 (N_921,N_466,N_90);
nor U922 (N_922,N_38,N_124);
nand U923 (N_923,N_232,N_130);
and U924 (N_924,N_379,N_429);
or U925 (N_925,N_505,N_249);
and U926 (N_926,N_331,N_557);
nand U927 (N_927,N_378,N_112);
nand U928 (N_928,N_246,N_394);
and U929 (N_929,N_310,N_377);
or U930 (N_930,N_558,N_247);
nor U931 (N_931,N_36,N_260);
nand U932 (N_932,N_592,N_429);
and U933 (N_933,N_499,N_39);
nand U934 (N_934,N_237,N_221);
and U935 (N_935,N_532,N_467);
nor U936 (N_936,N_555,N_437);
and U937 (N_937,N_282,N_116);
nand U938 (N_938,N_45,N_128);
nor U939 (N_939,N_106,N_357);
or U940 (N_940,N_27,N_356);
and U941 (N_941,N_145,N_443);
or U942 (N_942,N_168,N_578);
nor U943 (N_943,N_366,N_361);
nor U944 (N_944,N_80,N_575);
and U945 (N_945,N_463,N_311);
and U946 (N_946,N_455,N_131);
or U947 (N_947,N_271,N_450);
nand U948 (N_948,N_396,N_590);
or U949 (N_949,N_483,N_3);
nand U950 (N_950,N_268,N_97);
or U951 (N_951,N_23,N_101);
and U952 (N_952,N_570,N_172);
and U953 (N_953,N_115,N_233);
nand U954 (N_954,N_354,N_343);
nand U955 (N_955,N_96,N_67);
and U956 (N_956,N_67,N_306);
nand U957 (N_957,N_199,N_207);
nor U958 (N_958,N_237,N_550);
and U959 (N_959,N_42,N_256);
nor U960 (N_960,N_319,N_275);
and U961 (N_961,N_142,N_520);
and U962 (N_962,N_195,N_307);
or U963 (N_963,N_593,N_361);
xor U964 (N_964,N_468,N_231);
and U965 (N_965,N_199,N_134);
and U966 (N_966,N_8,N_459);
and U967 (N_967,N_537,N_39);
and U968 (N_968,N_352,N_239);
or U969 (N_969,N_589,N_115);
or U970 (N_970,N_487,N_106);
nand U971 (N_971,N_244,N_502);
or U972 (N_972,N_37,N_487);
nor U973 (N_973,N_103,N_44);
or U974 (N_974,N_349,N_460);
nor U975 (N_975,N_11,N_219);
and U976 (N_976,N_503,N_280);
nor U977 (N_977,N_403,N_392);
nand U978 (N_978,N_473,N_560);
nand U979 (N_979,N_598,N_234);
nand U980 (N_980,N_582,N_305);
or U981 (N_981,N_0,N_399);
or U982 (N_982,N_591,N_140);
nand U983 (N_983,N_554,N_79);
nor U984 (N_984,N_257,N_45);
nand U985 (N_985,N_496,N_225);
or U986 (N_986,N_514,N_14);
nor U987 (N_987,N_286,N_311);
or U988 (N_988,N_81,N_125);
nand U989 (N_989,N_86,N_522);
and U990 (N_990,N_491,N_585);
nand U991 (N_991,N_397,N_143);
and U992 (N_992,N_501,N_150);
and U993 (N_993,N_40,N_528);
nor U994 (N_994,N_416,N_259);
nor U995 (N_995,N_152,N_487);
and U996 (N_996,N_85,N_470);
nand U997 (N_997,N_327,N_357);
or U998 (N_998,N_454,N_193);
nand U999 (N_999,N_268,N_81);
and U1000 (N_1000,N_575,N_422);
and U1001 (N_1001,N_197,N_131);
nand U1002 (N_1002,N_371,N_370);
or U1003 (N_1003,N_257,N_567);
nand U1004 (N_1004,N_319,N_302);
nor U1005 (N_1005,N_483,N_427);
and U1006 (N_1006,N_598,N_179);
xnor U1007 (N_1007,N_137,N_345);
nor U1008 (N_1008,N_115,N_253);
and U1009 (N_1009,N_68,N_373);
and U1010 (N_1010,N_407,N_142);
nor U1011 (N_1011,N_548,N_178);
and U1012 (N_1012,N_479,N_277);
nand U1013 (N_1013,N_27,N_236);
nand U1014 (N_1014,N_208,N_106);
or U1015 (N_1015,N_28,N_458);
or U1016 (N_1016,N_325,N_393);
nand U1017 (N_1017,N_174,N_214);
or U1018 (N_1018,N_485,N_471);
and U1019 (N_1019,N_131,N_474);
nor U1020 (N_1020,N_473,N_176);
and U1021 (N_1021,N_395,N_467);
and U1022 (N_1022,N_333,N_544);
nor U1023 (N_1023,N_115,N_228);
or U1024 (N_1024,N_560,N_567);
nor U1025 (N_1025,N_581,N_210);
or U1026 (N_1026,N_129,N_222);
and U1027 (N_1027,N_414,N_186);
or U1028 (N_1028,N_249,N_241);
nand U1029 (N_1029,N_353,N_146);
nor U1030 (N_1030,N_554,N_99);
nor U1031 (N_1031,N_229,N_17);
or U1032 (N_1032,N_576,N_20);
and U1033 (N_1033,N_236,N_269);
nand U1034 (N_1034,N_21,N_228);
and U1035 (N_1035,N_462,N_82);
nor U1036 (N_1036,N_459,N_343);
nand U1037 (N_1037,N_599,N_468);
or U1038 (N_1038,N_429,N_499);
nor U1039 (N_1039,N_294,N_74);
nand U1040 (N_1040,N_97,N_411);
and U1041 (N_1041,N_122,N_542);
and U1042 (N_1042,N_443,N_402);
and U1043 (N_1043,N_529,N_355);
or U1044 (N_1044,N_344,N_535);
nand U1045 (N_1045,N_540,N_259);
and U1046 (N_1046,N_491,N_221);
or U1047 (N_1047,N_97,N_274);
or U1048 (N_1048,N_583,N_256);
and U1049 (N_1049,N_64,N_10);
nand U1050 (N_1050,N_578,N_371);
or U1051 (N_1051,N_428,N_332);
nor U1052 (N_1052,N_203,N_382);
nor U1053 (N_1053,N_512,N_398);
or U1054 (N_1054,N_283,N_209);
nor U1055 (N_1055,N_330,N_153);
nor U1056 (N_1056,N_550,N_436);
nor U1057 (N_1057,N_6,N_441);
nor U1058 (N_1058,N_365,N_492);
and U1059 (N_1059,N_209,N_117);
and U1060 (N_1060,N_341,N_157);
nand U1061 (N_1061,N_462,N_182);
nor U1062 (N_1062,N_481,N_296);
or U1063 (N_1063,N_558,N_88);
nand U1064 (N_1064,N_152,N_517);
nor U1065 (N_1065,N_338,N_109);
nor U1066 (N_1066,N_578,N_264);
or U1067 (N_1067,N_141,N_212);
and U1068 (N_1068,N_91,N_15);
nand U1069 (N_1069,N_575,N_518);
or U1070 (N_1070,N_558,N_329);
and U1071 (N_1071,N_37,N_503);
and U1072 (N_1072,N_295,N_396);
or U1073 (N_1073,N_245,N_130);
nor U1074 (N_1074,N_40,N_535);
nand U1075 (N_1075,N_125,N_357);
or U1076 (N_1076,N_158,N_430);
nor U1077 (N_1077,N_475,N_526);
and U1078 (N_1078,N_105,N_125);
nand U1079 (N_1079,N_121,N_546);
nor U1080 (N_1080,N_523,N_503);
or U1081 (N_1081,N_280,N_384);
nor U1082 (N_1082,N_563,N_569);
nand U1083 (N_1083,N_7,N_518);
and U1084 (N_1084,N_40,N_390);
nand U1085 (N_1085,N_262,N_406);
nor U1086 (N_1086,N_487,N_170);
nand U1087 (N_1087,N_441,N_62);
xnor U1088 (N_1088,N_262,N_551);
nand U1089 (N_1089,N_411,N_128);
nor U1090 (N_1090,N_282,N_10);
nand U1091 (N_1091,N_129,N_277);
and U1092 (N_1092,N_431,N_566);
and U1093 (N_1093,N_348,N_507);
nand U1094 (N_1094,N_577,N_576);
nor U1095 (N_1095,N_413,N_155);
and U1096 (N_1096,N_542,N_515);
nand U1097 (N_1097,N_406,N_174);
or U1098 (N_1098,N_17,N_254);
xor U1099 (N_1099,N_51,N_217);
or U1100 (N_1100,N_567,N_487);
nand U1101 (N_1101,N_316,N_574);
or U1102 (N_1102,N_544,N_451);
nor U1103 (N_1103,N_596,N_280);
nor U1104 (N_1104,N_382,N_158);
nand U1105 (N_1105,N_58,N_307);
and U1106 (N_1106,N_186,N_167);
nor U1107 (N_1107,N_202,N_421);
or U1108 (N_1108,N_163,N_452);
nand U1109 (N_1109,N_173,N_120);
xor U1110 (N_1110,N_209,N_63);
or U1111 (N_1111,N_444,N_271);
and U1112 (N_1112,N_40,N_220);
nor U1113 (N_1113,N_173,N_136);
and U1114 (N_1114,N_477,N_474);
or U1115 (N_1115,N_393,N_592);
nor U1116 (N_1116,N_140,N_563);
nor U1117 (N_1117,N_454,N_313);
nand U1118 (N_1118,N_347,N_335);
nand U1119 (N_1119,N_447,N_93);
nor U1120 (N_1120,N_253,N_494);
or U1121 (N_1121,N_105,N_349);
nor U1122 (N_1122,N_78,N_206);
nand U1123 (N_1123,N_162,N_440);
nand U1124 (N_1124,N_91,N_182);
nor U1125 (N_1125,N_567,N_8);
nor U1126 (N_1126,N_256,N_348);
and U1127 (N_1127,N_346,N_161);
nand U1128 (N_1128,N_226,N_46);
or U1129 (N_1129,N_169,N_214);
nand U1130 (N_1130,N_297,N_31);
nand U1131 (N_1131,N_512,N_287);
or U1132 (N_1132,N_365,N_189);
and U1133 (N_1133,N_291,N_206);
or U1134 (N_1134,N_16,N_295);
and U1135 (N_1135,N_387,N_460);
and U1136 (N_1136,N_96,N_434);
and U1137 (N_1137,N_554,N_205);
and U1138 (N_1138,N_15,N_549);
nand U1139 (N_1139,N_310,N_458);
or U1140 (N_1140,N_243,N_81);
nor U1141 (N_1141,N_550,N_141);
nor U1142 (N_1142,N_521,N_81);
nand U1143 (N_1143,N_161,N_479);
nor U1144 (N_1144,N_67,N_505);
or U1145 (N_1145,N_279,N_20);
xor U1146 (N_1146,N_113,N_417);
nor U1147 (N_1147,N_250,N_333);
nand U1148 (N_1148,N_35,N_276);
nor U1149 (N_1149,N_536,N_82);
nor U1150 (N_1150,N_386,N_518);
and U1151 (N_1151,N_161,N_268);
nor U1152 (N_1152,N_421,N_462);
nor U1153 (N_1153,N_231,N_478);
or U1154 (N_1154,N_308,N_235);
nor U1155 (N_1155,N_107,N_427);
and U1156 (N_1156,N_567,N_34);
or U1157 (N_1157,N_109,N_393);
nor U1158 (N_1158,N_579,N_439);
nor U1159 (N_1159,N_182,N_397);
nor U1160 (N_1160,N_297,N_149);
or U1161 (N_1161,N_129,N_33);
or U1162 (N_1162,N_205,N_452);
nor U1163 (N_1163,N_416,N_271);
nand U1164 (N_1164,N_83,N_252);
or U1165 (N_1165,N_6,N_393);
or U1166 (N_1166,N_143,N_105);
and U1167 (N_1167,N_484,N_283);
and U1168 (N_1168,N_389,N_42);
nor U1169 (N_1169,N_586,N_453);
nand U1170 (N_1170,N_338,N_166);
nor U1171 (N_1171,N_328,N_457);
nand U1172 (N_1172,N_575,N_284);
nor U1173 (N_1173,N_547,N_533);
or U1174 (N_1174,N_47,N_266);
nor U1175 (N_1175,N_387,N_524);
or U1176 (N_1176,N_348,N_500);
nor U1177 (N_1177,N_125,N_199);
nor U1178 (N_1178,N_582,N_261);
xnor U1179 (N_1179,N_575,N_330);
nand U1180 (N_1180,N_456,N_47);
xnor U1181 (N_1181,N_593,N_281);
or U1182 (N_1182,N_599,N_356);
or U1183 (N_1183,N_233,N_366);
or U1184 (N_1184,N_520,N_286);
nor U1185 (N_1185,N_229,N_445);
and U1186 (N_1186,N_75,N_155);
nand U1187 (N_1187,N_214,N_80);
nand U1188 (N_1188,N_281,N_231);
nand U1189 (N_1189,N_255,N_14);
or U1190 (N_1190,N_94,N_335);
nand U1191 (N_1191,N_69,N_190);
nor U1192 (N_1192,N_421,N_574);
nor U1193 (N_1193,N_492,N_177);
and U1194 (N_1194,N_373,N_515);
or U1195 (N_1195,N_109,N_500);
nand U1196 (N_1196,N_314,N_154);
and U1197 (N_1197,N_91,N_13);
nand U1198 (N_1198,N_248,N_142);
or U1199 (N_1199,N_122,N_242);
nor U1200 (N_1200,N_1178,N_664);
or U1201 (N_1201,N_917,N_704);
nand U1202 (N_1202,N_625,N_901);
or U1203 (N_1203,N_930,N_868);
and U1204 (N_1204,N_845,N_894);
nand U1205 (N_1205,N_1179,N_950);
and U1206 (N_1206,N_899,N_788);
nor U1207 (N_1207,N_759,N_748);
nand U1208 (N_1208,N_916,N_689);
nor U1209 (N_1209,N_1049,N_810);
or U1210 (N_1210,N_1104,N_896);
nor U1211 (N_1211,N_763,N_885);
nand U1212 (N_1212,N_1097,N_1060);
nor U1213 (N_1213,N_940,N_823);
or U1214 (N_1214,N_1164,N_1105);
nand U1215 (N_1215,N_730,N_1006);
or U1216 (N_1216,N_1038,N_1143);
and U1217 (N_1217,N_1007,N_1128);
nor U1218 (N_1218,N_771,N_884);
or U1219 (N_1219,N_862,N_696);
and U1220 (N_1220,N_942,N_692);
xnor U1221 (N_1221,N_765,N_774);
nor U1222 (N_1222,N_968,N_707);
or U1223 (N_1223,N_835,N_1051);
nand U1224 (N_1224,N_1155,N_630);
nor U1225 (N_1225,N_934,N_870);
and U1226 (N_1226,N_668,N_863);
xor U1227 (N_1227,N_1062,N_670);
and U1228 (N_1228,N_1187,N_860);
and U1229 (N_1229,N_826,N_632);
and U1230 (N_1230,N_912,N_639);
and U1231 (N_1231,N_1198,N_841);
and U1232 (N_1232,N_914,N_1027);
or U1233 (N_1233,N_705,N_1041);
nor U1234 (N_1234,N_1154,N_1093);
nor U1235 (N_1235,N_1050,N_606);
or U1236 (N_1236,N_687,N_770);
xnor U1237 (N_1237,N_1044,N_619);
nand U1238 (N_1238,N_666,N_722);
and U1239 (N_1239,N_731,N_654);
or U1240 (N_1240,N_641,N_711);
and U1241 (N_1241,N_811,N_1018);
or U1242 (N_1242,N_965,N_786);
and U1243 (N_1243,N_627,N_859);
xor U1244 (N_1244,N_1089,N_991);
or U1245 (N_1245,N_721,N_1034);
and U1246 (N_1246,N_1079,N_1037);
nor U1247 (N_1247,N_609,N_757);
or U1248 (N_1248,N_1111,N_970);
nor U1249 (N_1249,N_686,N_910);
and U1250 (N_1250,N_739,N_809);
or U1251 (N_1251,N_622,N_935);
xor U1252 (N_1252,N_645,N_742);
nor U1253 (N_1253,N_836,N_933);
nor U1254 (N_1254,N_720,N_915);
nor U1255 (N_1255,N_665,N_854);
nor U1256 (N_1256,N_685,N_655);
nor U1257 (N_1257,N_954,N_1152);
nand U1258 (N_1258,N_1072,N_1080);
nand U1259 (N_1259,N_659,N_701);
nand U1260 (N_1260,N_700,N_1162);
or U1261 (N_1261,N_679,N_853);
or U1262 (N_1262,N_657,N_649);
nor U1263 (N_1263,N_980,N_1009);
nand U1264 (N_1264,N_1077,N_618);
and U1265 (N_1265,N_617,N_732);
nand U1266 (N_1266,N_1107,N_989);
nand U1267 (N_1267,N_911,N_1197);
nor U1268 (N_1268,N_1048,N_1159);
and U1269 (N_1269,N_981,N_818);
nand U1270 (N_1270,N_620,N_1185);
xor U1271 (N_1271,N_672,N_1029);
or U1272 (N_1272,N_1015,N_1123);
nand U1273 (N_1273,N_1013,N_702);
and U1274 (N_1274,N_822,N_1098);
or U1275 (N_1275,N_1177,N_678);
and U1276 (N_1276,N_745,N_946);
and U1277 (N_1277,N_821,N_903);
and U1278 (N_1278,N_796,N_1022);
or U1279 (N_1279,N_1190,N_1075);
xnor U1280 (N_1280,N_847,N_754);
nand U1281 (N_1281,N_778,N_817);
nand U1282 (N_1282,N_755,N_1192);
nand U1283 (N_1283,N_1036,N_966);
and U1284 (N_1284,N_1199,N_1090);
nor U1285 (N_1285,N_1019,N_624);
or U1286 (N_1286,N_988,N_673);
or U1287 (N_1287,N_1172,N_1086);
and U1288 (N_1288,N_963,N_939);
nor U1289 (N_1289,N_974,N_1071);
nor U1290 (N_1290,N_651,N_1008);
xnor U1291 (N_1291,N_612,N_793);
nor U1292 (N_1292,N_777,N_864);
or U1293 (N_1293,N_886,N_958);
and U1294 (N_1294,N_772,N_955);
nand U1295 (N_1295,N_871,N_925);
or U1296 (N_1296,N_734,N_1134);
nand U1297 (N_1297,N_1180,N_1127);
nor U1298 (N_1298,N_648,N_636);
or U1299 (N_1299,N_1150,N_1167);
nand U1300 (N_1300,N_848,N_957);
nand U1301 (N_1301,N_795,N_1052);
nor U1302 (N_1302,N_891,N_1113);
nor U1303 (N_1303,N_1188,N_825);
nor U1304 (N_1304,N_824,N_1109);
nand U1305 (N_1305,N_808,N_1078);
or U1306 (N_1306,N_814,N_1042);
nand U1307 (N_1307,N_1108,N_1065);
nand U1308 (N_1308,N_1138,N_1116);
nor U1309 (N_1309,N_1045,N_984);
or U1310 (N_1310,N_855,N_875);
nor U1311 (N_1311,N_1012,N_913);
or U1312 (N_1312,N_756,N_768);
and U1313 (N_1313,N_837,N_1161);
nor U1314 (N_1314,N_923,N_1133);
or U1315 (N_1315,N_629,N_983);
and U1316 (N_1316,N_674,N_717);
nand U1317 (N_1317,N_943,N_727);
and U1318 (N_1318,N_713,N_775);
and U1319 (N_1319,N_872,N_741);
nand U1320 (N_1320,N_688,N_1103);
or U1321 (N_1321,N_782,N_849);
and U1322 (N_1322,N_779,N_1040);
and U1323 (N_1323,N_861,N_789);
and U1324 (N_1324,N_602,N_846);
and U1325 (N_1325,N_1100,N_610);
or U1326 (N_1326,N_724,N_681);
nand U1327 (N_1327,N_1053,N_1023);
and U1328 (N_1328,N_897,N_883);
nor U1329 (N_1329,N_764,N_1083);
or U1330 (N_1330,N_614,N_799);
or U1331 (N_1331,N_890,N_1119);
and U1332 (N_1332,N_706,N_921);
and U1333 (N_1333,N_656,N_747);
and U1334 (N_1334,N_1094,N_1136);
nand U1335 (N_1335,N_1194,N_878);
nor U1336 (N_1336,N_753,N_1130);
or U1337 (N_1337,N_893,N_1024);
and U1338 (N_1338,N_962,N_1026);
or U1339 (N_1339,N_807,N_882);
and U1340 (N_1340,N_1191,N_1066);
nand U1341 (N_1341,N_1073,N_1014);
nand U1342 (N_1342,N_1175,N_634);
or U1343 (N_1343,N_1149,N_876);
or U1344 (N_1344,N_1074,N_737);
and U1345 (N_1345,N_658,N_937);
and U1346 (N_1346,N_760,N_997);
or U1347 (N_1347,N_1033,N_813);
nand U1348 (N_1348,N_829,N_1035);
and U1349 (N_1349,N_1166,N_879);
or U1350 (N_1350,N_959,N_931);
or U1351 (N_1351,N_953,N_1115);
or U1352 (N_1352,N_738,N_839);
nor U1353 (N_1353,N_880,N_801);
nand U1354 (N_1354,N_712,N_1028);
nand U1355 (N_1355,N_675,N_716);
nor U1356 (N_1356,N_1055,N_708);
nand U1357 (N_1357,N_888,N_1156);
nand U1358 (N_1358,N_873,N_949);
nor U1359 (N_1359,N_792,N_797);
or U1360 (N_1360,N_964,N_1059);
and U1361 (N_1361,N_746,N_718);
nand U1362 (N_1362,N_918,N_1146);
and U1363 (N_1363,N_1032,N_909);
xnor U1364 (N_1364,N_740,N_699);
nand U1365 (N_1365,N_647,N_1047);
nor U1366 (N_1366,N_857,N_972);
or U1367 (N_1367,N_1176,N_1110);
and U1368 (N_1368,N_902,N_1114);
or U1369 (N_1369,N_604,N_616);
and U1370 (N_1370,N_867,N_979);
nor U1371 (N_1371,N_729,N_1112);
or U1372 (N_1372,N_723,N_1160);
nor U1373 (N_1373,N_733,N_1069);
or U1374 (N_1374,N_892,N_693);
nor U1375 (N_1375,N_626,N_714);
or U1376 (N_1376,N_928,N_631);
nand U1377 (N_1377,N_1144,N_1021);
nor U1378 (N_1378,N_802,N_736);
or U1379 (N_1379,N_956,N_850);
nand U1380 (N_1380,N_843,N_1000);
and U1381 (N_1381,N_1118,N_615);
and U1382 (N_1382,N_1129,N_1092);
nor U1383 (N_1383,N_804,N_780);
nand U1384 (N_1384,N_936,N_944);
nand U1385 (N_1385,N_1002,N_834);
nand U1386 (N_1386,N_652,N_697);
and U1387 (N_1387,N_1141,N_684);
and U1388 (N_1388,N_1170,N_787);
and U1389 (N_1389,N_851,N_613);
or U1390 (N_1390,N_1122,N_680);
or U1391 (N_1391,N_663,N_762);
or U1392 (N_1392,N_812,N_646);
and U1393 (N_1393,N_948,N_996);
and U1394 (N_1394,N_638,N_1039);
nand U1395 (N_1395,N_978,N_1082);
or U1396 (N_1396,N_1132,N_941);
nor U1397 (N_1397,N_869,N_600);
and U1398 (N_1398,N_858,N_1031);
nand U1399 (N_1399,N_1046,N_1151);
nand U1400 (N_1400,N_831,N_1001);
nor U1401 (N_1401,N_667,N_653);
nor U1402 (N_1402,N_920,N_1121);
and U1403 (N_1403,N_815,N_1184);
nor U1404 (N_1404,N_1157,N_1140);
nand U1405 (N_1405,N_1081,N_1124);
or U1406 (N_1406,N_660,N_1070);
nand U1407 (N_1407,N_895,N_904);
or U1408 (N_1408,N_994,N_1010);
and U1409 (N_1409,N_919,N_900);
nor U1410 (N_1410,N_1067,N_783);
and U1411 (N_1411,N_973,N_816);
and U1412 (N_1412,N_838,N_1125);
or U1413 (N_1413,N_924,N_866);
nor U1414 (N_1414,N_710,N_781);
or U1415 (N_1415,N_803,N_677);
or U1416 (N_1416,N_1163,N_932);
and U1417 (N_1417,N_800,N_785);
or U1418 (N_1418,N_889,N_1043);
and U1419 (N_1419,N_683,N_767);
and U1420 (N_1420,N_929,N_938);
nor U1421 (N_1421,N_1057,N_999);
and U1422 (N_1422,N_691,N_877);
or U1423 (N_1423,N_798,N_761);
or U1424 (N_1424,N_671,N_840);
nand U1425 (N_1425,N_990,N_976);
nand U1426 (N_1426,N_842,N_735);
and U1427 (N_1427,N_856,N_952);
or U1428 (N_1428,N_844,N_1131);
nand U1429 (N_1429,N_819,N_975);
and U1430 (N_1430,N_640,N_1117);
or U1431 (N_1431,N_881,N_947);
nand U1432 (N_1432,N_906,N_682);
nor U1433 (N_1433,N_828,N_1174);
and U1434 (N_1434,N_643,N_695);
and U1435 (N_1435,N_623,N_642);
nor U1436 (N_1436,N_1084,N_662);
nand U1437 (N_1437,N_715,N_1153);
nor U1438 (N_1438,N_1063,N_637);
nand U1439 (N_1439,N_1147,N_1095);
or U1440 (N_1440,N_1183,N_1145);
nor U1441 (N_1441,N_698,N_1142);
xnor U1442 (N_1442,N_971,N_1096);
nand U1443 (N_1443,N_773,N_749);
or U1444 (N_1444,N_1004,N_1158);
or U1445 (N_1445,N_926,N_1088);
or U1446 (N_1446,N_982,N_633);
and U1447 (N_1447,N_1005,N_1196);
and U1448 (N_1448,N_661,N_922);
and U1449 (N_1449,N_805,N_1181);
or U1450 (N_1450,N_1085,N_605);
and U1451 (N_1451,N_766,N_728);
nor U1452 (N_1452,N_719,N_874);
nand U1453 (N_1453,N_945,N_1061);
or U1454 (N_1454,N_628,N_743);
nand U1455 (N_1455,N_1173,N_1106);
and U1456 (N_1456,N_967,N_907);
nor U1457 (N_1457,N_603,N_690);
xnor U1458 (N_1458,N_905,N_1189);
and U1459 (N_1459,N_827,N_709);
and U1460 (N_1460,N_1139,N_1165);
nor U1461 (N_1461,N_977,N_601);
xor U1462 (N_1462,N_1169,N_611);
nor U1463 (N_1463,N_865,N_908);
and U1464 (N_1464,N_898,N_1056);
nand U1465 (N_1465,N_998,N_992);
nand U1466 (N_1466,N_769,N_794);
nand U1467 (N_1467,N_993,N_927);
nand U1468 (N_1468,N_1168,N_969);
or U1469 (N_1469,N_1020,N_621);
or U1470 (N_1470,N_1193,N_1016);
nand U1471 (N_1471,N_1126,N_985);
and U1472 (N_1472,N_1011,N_776);
nor U1473 (N_1473,N_1003,N_790);
nor U1474 (N_1474,N_887,N_703);
nand U1475 (N_1475,N_751,N_1087);
or U1476 (N_1476,N_986,N_694);
nor U1477 (N_1477,N_635,N_820);
nand U1478 (N_1478,N_960,N_1068);
nand U1479 (N_1479,N_987,N_725);
or U1480 (N_1480,N_607,N_806);
and U1481 (N_1481,N_1137,N_1091);
or U1482 (N_1482,N_1099,N_1025);
nor U1483 (N_1483,N_758,N_995);
nor U1484 (N_1484,N_852,N_1064);
or U1485 (N_1485,N_1030,N_1058);
and U1486 (N_1486,N_832,N_750);
or U1487 (N_1487,N_1054,N_644);
nand U1488 (N_1488,N_608,N_791);
and U1489 (N_1489,N_784,N_833);
nor U1490 (N_1490,N_726,N_1102);
or U1491 (N_1491,N_1171,N_1186);
or U1492 (N_1492,N_1120,N_1135);
and U1493 (N_1493,N_676,N_650);
and U1494 (N_1494,N_951,N_1017);
and U1495 (N_1495,N_1076,N_1101);
nand U1496 (N_1496,N_1148,N_1182);
and U1497 (N_1497,N_752,N_961);
nand U1498 (N_1498,N_744,N_830);
nand U1499 (N_1499,N_669,N_1195);
nand U1500 (N_1500,N_690,N_1083);
nand U1501 (N_1501,N_816,N_894);
and U1502 (N_1502,N_677,N_1058);
nor U1503 (N_1503,N_741,N_938);
or U1504 (N_1504,N_726,N_1184);
and U1505 (N_1505,N_992,N_1040);
xnor U1506 (N_1506,N_769,N_855);
nor U1507 (N_1507,N_773,N_921);
nor U1508 (N_1508,N_1123,N_941);
and U1509 (N_1509,N_804,N_784);
and U1510 (N_1510,N_982,N_677);
and U1511 (N_1511,N_658,N_623);
nor U1512 (N_1512,N_756,N_1159);
nor U1513 (N_1513,N_1173,N_1164);
nor U1514 (N_1514,N_757,N_972);
nor U1515 (N_1515,N_755,N_1001);
nor U1516 (N_1516,N_1128,N_897);
nand U1517 (N_1517,N_1065,N_1030);
nor U1518 (N_1518,N_791,N_631);
or U1519 (N_1519,N_996,N_644);
or U1520 (N_1520,N_843,N_815);
nand U1521 (N_1521,N_985,N_1165);
and U1522 (N_1522,N_1138,N_673);
and U1523 (N_1523,N_948,N_677);
nand U1524 (N_1524,N_1046,N_808);
nand U1525 (N_1525,N_731,N_1020);
nand U1526 (N_1526,N_749,N_838);
or U1527 (N_1527,N_683,N_1044);
or U1528 (N_1528,N_1033,N_774);
and U1529 (N_1529,N_869,N_826);
nor U1530 (N_1530,N_603,N_1161);
nor U1531 (N_1531,N_975,N_1089);
nor U1532 (N_1532,N_871,N_1056);
nand U1533 (N_1533,N_998,N_1025);
and U1534 (N_1534,N_722,N_1188);
and U1535 (N_1535,N_1039,N_862);
nand U1536 (N_1536,N_712,N_851);
nor U1537 (N_1537,N_875,N_1161);
and U1538 (N_1538,N_765,N_967);
and U1539 (N_1539,N_1042,N_716);
and U1540 (N_1540,N_621,N_882);
nor U1541 (N_1541,N_760,N_1047);
and U1542 (N_1542,N_971,N_1112);
nand U1543 (N_1543,N_1062,N_937);
nand U1544 (N_1544,N_642,N_951);
and U1545 (N_1545,N_966,N_825);
nand U1546 (N_1546,N_1186,N_747);
or U1547 (N_1547,N_759,N_776);
nand U1548 (N_1548,N_905,N_1049);
and U1549 (N_1549,N_751,N_1154);
or U1550 (N_1550,N_686,N_1116);
nor U1551 (N_1551,N_849,N_1191);
nand U1552 (N_1552,N_901,N_676);
nor U1553 (N_1553,N_1160,N_659);
or U1554 (N_1554,N_793,N_903);
nor U1555 (N_1555,N_854,N_690);
xor U1556 (N_1556,N_709,N_1191);
nand U1557 (N_1557,N_925,N_807);
and U1558 (N_1558,N_1075,N_712);
and U1559 (N_1559,N_656,N_932);
nor U1560 (N_1560,N_763,N_1120);
or U1561 (N_1561,N_1033,N_719);
nand U1562 (N_1562,N_952,N_1059);
or U1563 (N_1563,N_920,N_1046);
nor U1564 (N_1564,N_998,N_909);
xnor U1565 (N_1565,N_961,N_638);
nand U1566 (N_1566,N_977,N_1197);
and U1567 (N_1567,N_768,N_972);
and U1568 (N_1568,N_1104,N_1195);
xnor U1569 (N_1569,N_1014,N_1154);
and U1570 (N_1570,N_909,N_1036);
and U1571 (N_1571,N_1142,N_1173);
nor U1572 (N_1572,N_1098,N_1030);
or U1573 (N_1573,N_906,N_1008);
and U1574 (N_1574,N_1011,N_990);
nand U1575 (N_1575,N_905,N_956);
and U1576 (N_1576,N_959,N_676);
nand U1577 (N_1577,N_864,N_617);
nor U1578 (N_1578,N_983,N_972);
or U1579 (N_1579,N_1160,N_728);
nand U1580 (N_1580,N_744,N_953);
or U1581 (N_1581,N_1141,N_1095);
or U1582 (N_1582,N_981,N_881);
and U1583 (N_1583,N_632,N_961);
nand U1584 (N_1584,N_1076,N_1036);
or U1585 (N_1585,N_703,N_870);
and U1586 (N_1586,N_1172,N_653);
nor U1587 (N_1587,N_622,N_648);
and U1588 (N_1588,N_632,N_936);
nand U1589 (N_1589,N_780,N_600);
or U1590 (N_1590,N_892,N_926);
or U1591 (N_1591,N_1126,N_917);
nand U1592 (N_1592,N_1117,N_885);
nand U1593 (N_1593,N_749,N_846);
or U1594 (N_1594,N_1159,N_770);
xor U1595 (N_1595,N_854,N_916);
or U1596 (N_1596,N_971,N_703);
and U1597 (N_1597,N_783,N_930);
and U1598 (N_1598,N_870,N_1040);
or U1599 (N_1599,N_1086,N_1006);
nor U1600 (N_1600,N_707,N_760);
nor U1601 (N_1601,N_1165,N_734);
nor U1602 (N_1602,N_603,N_881);
or U1603 (N_1603,N_938,N_926);
nand U1604 (N_1604,N_688,N_806);
and U1605 (N_1605,N_965,N_742);
and U1606 (N_1606,N_672,N_890);
and U1607 (N_1607,N_1044,N_701);
nand U1608 (N_1608,N_1000,N_1140);
nor U1609 (N_1609,N_949,N_741);
or U1610 (N_1610,N_683,N_906);
nor U1611 (N_1611,N_1115,N_963);
or U1612 (N_1612,N_1023,N_1055);
xnor U1613 (N_1613,N_992,N_601);
nor U1614 (N_1614,N_735,N_618);
or U1615 (N_1615,N_893,N_1120);
nand U1616 (N_1616,N_1069,N_902);
nor U1617 (N_1617,N_1022,N_906);
or U1618 (N_1618,N_770,N_944);
or U1619 (N_1619,N_1171,N_964);
or U1620 (N_1620,N_831,N_734);
or U1621 (N_1621,N_872,N_757);
nand U1622 (N_1622,N_944,N_821);
nand U1623 (N_1623,N_902,N_1173);
nand U1624 (N_1624,N_816,N_718);
or U1625 (N_1625,N_783,N_1195);
nand U1626 (N_1626,N_1045,N_969);
nor U1627 (N_1627,N_850,N_1123);
nor U1628 (N_1628,N_1179,N_921);
nor U1629 (N_1629,N_733,N_899);
or U1630 (N_1630,N_781,N_625);
and U1631 (N_1631,N_876,N_720);
nor U1632 (N_1632,N_904,N_745);
nand U1633 (N_1633,N_1095,N_1124);
nor U1634 (N_1634,N_638,N_950);
nand U1635 (N_1635,N_1080,N_967);
or U1636 (N_1636,N_813,N_1149);
nor U1637 (N_1637,N_925,N_656);
xor U1638 (N_1638,N_1164,N_957);
xor U1639 (N_1639,N_1014,N_837);
nor U1640 (N_1640,N_1014,N_687);
xor U1641 (N_1641,N_731,N_1027);
and U1642 (N_1642,N_1050,N_846);
nand U1643 (N_1643,N_736,N_885);
or U1644 (N_1644,N_993,N_959);
or U1645 (N_1645,N_1009,N_653);
or U1646 (N_1646,N_757,N_1018);
or U1647 (N_1647,N_657,N_849);
or U1648 (N_1648,N_721,N_811);
nand U1649 (N_1649,N_684,N_759);
nand U1650 (N_1650,N_1060,N_1083);
xnor U1651 (N_1651,N_1063,N_1132);
or U1652 (N_1652,N_812,N_1117);
nand U1653 (N_1653,N_956,N_659);
and U1654 (N_1654,N_1020,N_759);
nand U1655 (N_1655,N_809,N_1010);
xor U1656 (N_1656,N_733,N_792);
nand U1657 (N_1657,N_779,N_951);
or U1658 (N_1658,N_791,N_1184);
nand U1659 (N_1659,N_604,N_915);
nor U1660 (N_1660,N_805,N_770);
nand U1661 (N_1661,N_994,N_805);
nor U1662 (N_1662,N_811,N_920);
and U1663 (N_1663,N_925,N_789);
or U1664 (N_1664,N_833,N_646);
nand U1665 (N_1665,N_785,N_790);
and U1666 (N_1666,N_631,N_927);
or U1667 (N_1667,N_1119,N_1026);
nor U1668 (N_1668,N_614,N_648);
nor U1669 (N_1669,N_965,N_998);
nand U1670 (N_1670,N_1072,N_980);
nand U1671 (N_1671,N_673,N_1187);
or U1672 (N_1672,N_1034,N_839);
nand U1673 (N_1673,N_869,N_1081);
or U1674 (N_1674,N_1067,N_1119);
or U1675 (N_1675,N_833,N_895);
and U1676 (N_1676,N_809,N_1021);
nand U1677 (N_1677,N_688,N_922);
xor U1678 (N_1678,N_1001,N_1047);
or U1679 (N_1679,N_943,N_667);
nand U1680 (N_1680,N_755,N_643);
and U1681 (N_1681,N_681,N_645);
or U1682 (N_1682,N_764,N_691);
nand U1683 (N_1683,N_986,N_653);
nor U1684 (N_1684,N_739,N_998);
nor U1685 (N_1685,N_893,N_936);
or U1686 (N_1686,N_680,N_819);
and U1687 (N_1687,N_900,N_676);
nand U1688 (N_1688,N_957,N_715);
and U1689 (N_1689,N_635,N_962);
and U1690 (N_1690,N_1139,N_1159);
and U1691 (N_1691,N_903,N_1075);
nand U1692 (N_1692,N_903,N_674);
nand U1693 (N_1693,N_1101,N_1169);
or U1694 (N_1694,N_690,N_684);
or U1695 (N_1695,N_918,N_941);
or U1696 (N_1696,N_668,N_1115);
xor U1697 (N_1697,N_1084,N_1061);
and U1698 (N_1698,N_819,N_1130);
and U1699 (N_1699,N_786,N_770);
and U1700 (N_1700,N_1144,N_1111);
nor U1701 (N_1701,N_1147,N_1020);
and U1702 (N_1702,N_1185,N_888);
or U1703 (N_1703,N_1144,N_1194);
nor U1704 (N_1704,N_1124,N_998);
or U1705 (N_1705,N_1149,N_928);
or U1706 (N_1706,N_710,N_815);
xnor U1707 (N_1707,N_713,N_1195);
nor U1708 (N_1708,N_797,N_925);
and U1709 (N_1709,N_1013,N_845);
nand U1710 (N_1710,N_845,N_1113);
nor U1711 (N_1711,N_1098,N_890);
and U1712 (N_1712,N_1139,N_1055);
nand U1713 (N_1713,N_1150,N_1096);
nor U1714 (N_1714,N_982,N_1056);
nand U1715 (N_1715,N_680,N_755);
or U1716 (N_1716,N_616,N_949);
nand U1717 (N_1717,N_1151,N_603);
or U1718 (N_1718,N_1126,N_1195);
or U1719 (N_1719,N_813,N_892);
or U1720 (N_1720,N_956,N_901);
nand U1721 (N_1721,N_827,N_936);
nand U1722 (N_1722,N_688,N_1089);
or U1723 (N_1723,N_1123,N_809);
and U1724 (N_1724,N_987,N_652);
and U1725 (N_1725,N_714,N_868);
nand U1726 (N_1726,N_673,N_786);
and U1727 (N_1727,N_660,N_710);
nor U1728 (N_1728,N_1082,N_1031);
nand U1729 (N_1729,N_997,N_991);
nand U1730 (N_1730,N_754,N_985);
and U1731 (N_1731,N_713,N_629);
nor U1732 (N_1732,N_635,N_861);
and U1733 (N_1733,N_919,N_842);
nor U1734 (N_1734,N_634,N_1099);
and U1735 (N_1735,N_1114,N_976);
nor U1736 (N_1736,N_1015,N_917);
nand U1737 (N_1737,N_643,N_1098);
nand U1738 (N_1738,N_734,N_935);
nor U1739 (N_1739,N_997,N_1178);
and U1740 (N_1740,N_814,N_661);
and U1741 (N_1741,N_1049,N_983);
or U1742 (N_1742,N_1032,N_1176);
or U1743 (N_1743,N_749,N_1085);
or U1744 (N_1744,N_967,N_863);
nand U1745 (N_1745,N_674,N_1084);
nand U1746 (N_1746,N_896,N_934);
nor U1747 (N_1747,N_676,N_1016);
and U1748 (N_1748,N_1024,N_954);
and U1749 (N_1749,N_1062,N_715);
xor U1750 (N_1750,N_1100,N_1198);
nand U1751 (N_1751,N_665,N_737);
or U1752 (N_1752,N_1178,N_922);
and U1753 (N_1753,N_975,N_904);
and U1754 (N_1754,N_1152,N_875);
xor U1755 (N_1755,N_1086,N_607);
xnor U1756 (N_1756,N_666,N_930);
nor U1757 (N_1757,N_1104,N_686);
or U1758 (N_1758,N_716,N_1104);
or U1759 (N_1759,N_617,N_904);
or U1760 (N_1760,N_747,N_1104);
nor U1761 (N_1761,N_745,N_817);
and U1762 (N_1762,N_608,N_831);
nor U1763 (N_1763,N_915,N_1007);
or U1764 (N_1764,N_952,N_1083);
nor U1765 (N_1765,N_1077,N_884);
nand U1766 (N_1766,N_1023,N_1003);
and U1767 (N_1767,N_719,N_735);
nor U1768 (N_1768,N_829,N_850);
nor U1769 (N_1769,N_1133,N_905);
or U1770 (N_1770,N_777,N_1008);
nand U1771 (N_1771,N_946,N_623);
and U1772 (N_1772,N_766,N_1109);
and U1773 (N_1773,N_999,N_782);
or U1774 (N_1774,N_814,N_669);
and U1775 (N_1775,N_999,N_678);
nand U1776 (N_1776,N_1061,N_1114);
xnor U1777 (N_1777,N_1067,N_833);
or U1778 (N_1778,N_850,N_723);
nand U1779 (N_1779,N_912,N_1174);
and U1780 (N_1780,N_700,N_704);
nor U1781 (N_1781,N_1040,N_1077);
nand U1782 (N_1782,N_1196,N_972);
and U1783 (N_1783,N_1095,N_950);
nand U1784 (N_1784,N_1083,N_912);
and U1785 (N_1785,N_879,N_956);
nor U1786 (N_1786,N_1045,N_828);
nand U1787 (N_1787,N_846,N_1190);
nor U1788 (N_1788,N_1031,N_1002);
nor U1789 (N_1789,N_1131,N_1025);
nand U1790 (N_1790,N_960,N_867);
nor U1791 (N_1791,N_807,N_1191);
nor U1792 (N_1792,N_710,N_618);
or U1793 (N_1793,N_781,N_1121);
nor U1794 (N_1794,N_760,N_932);
or U1795 (N_1795,N_725,N_833);
nand U1796 (N_1796,N_877,N_819);
nand U1797 (N_1797,N_604,N_886);
nor U1798 (N_1798,N_627,N_794);
xor U1799 (N_1799,N_1080,N_758);
nor U1800 (N_1800,N_1348,N_1547);
or U1801 (N_1801,N_1609,N_1437);
or U1802 (N_1802,N_1585,N_1444);
nand U1803 (N_1803,N_1646,N_1700);
nand U1804 (N_1804,N_1616,N_1783);
nor U1805 (N_1805,N_1400,N_1294);
and U1806 (N_1806,N_1758,N_1684);
or U1807 (N_1807,N_1429,N_1375);
nor U1808 (N_1808,N_1649,N_1426);
or U1809 (N_1809,N_1702,N_1371);
nand U1810 (N_1810,N_1680,N_1351);
or U1811 (N_1811,N_1264,N_1447);
nand U1812 (N_1812,N_1404,N_1655);
nor U1813 (N_1813,N_1201,N_1498);
and U1814 (N_1814,N_1712,N_1335);
nand U1815 (N_1815,N_1787,N_1548);
or U1816 (N_1816,N_1657,N_1673);
nor U1817 (N_1817,N_1604,N_1499);
or U1818 (N_1818,N_1295,N_1454);
nand U1819 (N_1819,N_1588,N_1645);
nand U1820 (N_1820,N_1734,N_1267);
and U1821 (N_1821,N_1664,N_1519);
nor U1822 (N_1822,N_1443,N_1324);
or U1823 (N_1823,N_1601,N_1225);
and U1824 (N_1824,N_1428,N_1279);
or U1825 (N_1825,N_1471,N_1597);
and U1826 (N_1826,N_1570,N_1651);
and U1827 (N_1827,N_1252,N_1514);
nor U1828 (N_1828,N_1674,N_1656);
nor U1829 (N_1829,N_1671,N_1448);
nand U1830 (N_1830,N_1511,N_1359);
nor U1831 (N_1831,N_1303,N_1515);
or U1832 (N_1832,N_1796,N_1211);
and U1833 (N_1833,N_1708,N_1624);
nor U1834 (N_1834,N_1338,N_1269);
or U1835 (N_1835,N_1383,N_1529);
nand U1836 (N_1836,N_1410,N_1579);
or U1837 (N_1837,N_1212,N_1685);
or U1838 (N_1838,N_1696,N_1461);
nor U1839 (N_1839,N_1272,N_1229);
and U1840 (N_1840,N_1524,N_1364);
or U1841 (N_1841,N_1350,N_1453);
or U1842 (N_1842,N_1670,N_1772);
nor U1843 (N_1843,N_1701,N_1724);
and U1844 (N_1844,N_1270,N_1779);
or U1845 (N_1845,N_1476,N_1532);
and U1846 (N_1846,N_1481,N_1276);
or U1847 (N_1847,N_1633,N_1480);
and U1848 (N_1848,N_1274,N_1574);
nor U1849 (N_1849,N_1500,N_1384);
or U1850 (N_1850,N_1320,N_1522);
or U1851 (N_1851,N_1330,N_1691);
nand U1852 (N_1852,N_1669,N_1341);
nand U1853 (N_1853,N_1305,N_1402);
or U1854 (N_1854,N_1623,N_1798);
nor U1855 (N_1855,N_1339,N_1366);
and U1856 (N_1856,N_1663,N_1730);
or U1857 (N_1857,N_1263,N_1788);
and U1858 (N_1858,N_1705,N_1586);
nor U1859 (N_1859,N_1243,N_1228);
nand U1860 (N_1860,N_1716,N_1729);
nor U1861 (N_1861,N_1769,N_1445);
or U1862 (N_1862,N_1304,N_1752);
nor U1863 (N_1863,N_1581,N_1695);
and U1864 (N_1864,N_1709,N_1761);
nand U1865 (N_1865,N_1284,N_1414);
nand U1866 (N_1866,N_1288,N_1707);
or U1867 (N_1867,N_1541,N_1205);
or U1868 (N_1868,N_1418,N_1227);
or U1869 (N_1869,N_1727,N_1732);
and U1870 (N_1870,N_1407,N_1391);
or U1871 (N_1871,N_1565,N_1714);
nand U1872 (N_1872,N_1754,N_1387);
nor U1873 (N_1873,N_1658,N_1667);
or U1874 (N_1874,N_1564,N_1449);
nor U1875 (N_1875,N_1254,N_1309);
or U1876 (N_1876,N_1283,N_1533);
or U1877 (N_1877,N_1567,N_1306);
or U1878 (N_1878,N_1736,N_1217);
and U1879 (N_1879,N_1537,N_1210);
nor U1880 (N_1880,N_1494,N_1509);
nor U1881 (N_1881,N_1568,N_1325);
or U1882 (N_1882,N_1462,N_1777);
and U1883 (N_1883,N_1208,N_1689);
nor U1884 (N_1884,N_1631,N_1472);
or U1885 (N_1885,N_1256,N_1662);
or U1886 (N_1886,N_1661,N_1213);
or U1887 (N_1887,N_1576,N_1654);
nor U1888 (N_1888,N_1452,N_1474);
nor U1889 (N_1889,N_1460,N_1742);
and U1890 (N_1890,N_1760,N_1678);
or U1891 (N_1891,N_1555,N_1679);
and U1892 (N_1892,N_1259,N_1411);
and U1893 (N_1893,N_1442,N_1334);
nor U1894 (N_1894,N_1572,N_1419);
nand U1895 (N_1895,N_1762,N_1245);
and U1896 (N_1896,N_1560,N_1326);
nand U1897 (N_1897,N_1451,N_1753);
nor U1898 (N_1898,N_1795,N_1425);
nand U1899 (N_1899,N_1374,N_1508);
nor U1900 (N_1900,N_1219,N_1526);
nand U1901 (N_1901,N_1506,N_1312);
or U1902 (N_1902,N_1469,N_1782);
nor U1903 (N_1903,N_1550,N_1482);
and U1904 (N_1904,N_1607,N_1751);
nor U1905 (N_1905,N_1590,N_1643);
nand U1906 (N_1906,N_1473,N_1580);
or U1907 (N_1907,N_1257,N_1323);
and U1908 (N_1908,N_1458,N_1492);
nor U1909 (N_1909,N_1440,N_1457);
nor U1910 (N_1910,N_1468,N_1766);
or U1911 (N_1911,N_1315,N_1546);
nor U1912 (N_1912,N_1553,N_1699);
nor U1913 (N_1913,N_1479,N_1289);
and U1914 (N_1914,N_1698,N_1441);
or U1915 (N_1915,N_1595,N_1393);
nand U1916 (N_1916,N_1220,N_1412);
and U1917 (N_1917,N_1518,N_1347);
nand U1918 (N_1918,N_1261,N_1693);
nand U1919 (N_1919,N_1557,N_1281);
nor U1920 (N_1920,N_1310,N_1436);
and U1921 (N_1921,N_1427,N_1744);
or U1922 (N_1922,N_1589,N_1369);
nor U1923 (N_1923,N_1490,N_1459);
xor U1924 (N_1924,N_1539,N_1573);
and U1925 (N_1925,N_1238,N_1642);
and U1926 (N_1926,N_1767,N_1439);
and U1927 (N_1927,N_1501,N_1596);
and U1928 (N_1928,N_1614,N_1781);
or U1929 (N_1929,N_1697,N_1349);
nand U1930 (N_1930,N_1307,N_1578);
and U1931 (N_1931,N_1389,N_1434);
and U1932 (N_1932,N_1582,N_1260);
nand U1933 (N_1933,N_1665,N_1619);
or U1934 (N_1934,N_1713,N_1398);
nand U1935 (N_1935,N_1620,N_1521);
nand U1936 (N_1936,N_1435,N_1241);
nand U1937 (N_1937,N_1372,N_1677);
or U1938 (N_1938,N_1632,N_1690);
or U1939 (N_1939,N_1226,N_1659);
or U1940 (N_1940,N_1799,N_1239);
or U1941 (N_1941,N_1485,N_1549);
or U1942 (N_1942,N_1255,N_1622);
or U1943 (N_1943,N_1466,N_1721);
nand U1944 (N_1944,N_1493,N_1647);
and U1945 (N_1945,N_1342,N_1528);
nand U1946 (N_1946,N_1456,N_1356);
nand U1947 (N_1947,N_1648,N_1629);
and U1948 (N_1948,N_1463,N_1794);
or U1949 (N_1949,N_1584,N_1785);
nand U1950 (N_1950,N_1681,N_1363);
or U1951 (N_1951,N_1365,N_1280);
or U1952 (N_1952,N_1401,N_1653);
nor U1953 (N_1953,N_1626,N_1298);
nand U1954 (N_1954,N_1333,N_1465);
nor U1955 (N_1955,N_1408,N_1415);
nor U1956 (N_1956,N_1242,N_1797);
nand U1957 (N_1957,N_1248,N_1599);
nand U1958 (N_1958,N_1244,N_1237);
and U1959 (N_1959,N_1683,N_1637);
and U1960 (N_1960,N_1543,N_1703);
and U1961 (N_1961,N_1396,N_1392);
or U1962 (N_1962,N_1345,N_1293);
or U1963 (N_1963,N_1748,N_1344);
and U1964 (N_1964,N_1329,N_1715);
nor U1965 (N_1965,N_1545,N_1223);
and U1966 (N_1966,N_1566,N_1406);
and U1967 (N_1967,N_1786,N_1755);
or U1968 (N_1968,N_1591,N_1497);
xnor U1969 (N_1969,N_1507,N_1577);
nand U1970 (N_1970,N_1611,N_1775);
and U1971 (N_1971,N_1368,N_1784);
nand U1972 (N_1972,N_1385,N_1353);
xor U1973 (N_1973,N_1793,N_1346);
and U1974 (N_1974,N_1361,N_1668);
nor U1975 (N_1975,N_1395,N_1525);
and U1976 (N_1976,N_1285,N_1612);
nor U1977 (N_1977,N_1692,N_1378);
and U1978 (N_1978,N_1236,N_1711);
or U1979 (N_1979,N_1706,N_1510);
nor U1980 (N_1980,N_1286,N_1438);
and U1981 (N_1981,N_1790,N_1571);
and U1982 (N_1982,N_1464,N_1486);
nor U1983 (N_1983,N_1757,N_1302);
or U1984 (N_1984,N_1749,N_1367);
and U1985 (N_1985,N_1308,N_1502);
and U1986 (N_1986,N_1328,N_1424);
and U1987 (N_1987,N_1535,N_1613);
and U1988 (N_1988,N_1605,N_1731);
nor U1989 (N_1989,N_1209,N_1523);
and U1990 (N_1990,N_1530,N_1446);
or U1991 (N_1991,N_1204,N_1373);
nor U1992 (N_1992,N_1296,N_1634);
nand U1993 (N_1993,N_1635,N_1215);
or U1994 (N_1994,N_1520,N_1627);
or U1995 (N_1995,N_1641,N_1247);
and U1996 (N_1996,N_1340,N_1603);
and U1997 (N_1997,N_1314,N_1686);
nand U1998 (N_1998,N_1625,N_1575);
and U1999 (N_1999,N_1455,N_1390);
and U2000 (N_2000,N_1773,N_1740);
nand U2001 (N_2001,N_1222,N_1399);
nand U2002 (N_2002,N_1231,N_1672);
and U2003 (N_2003,N_1676,N_1517);
and U2004 (N_2004,N_1376,N_1540);
nand U2005 (N_2005,N_1487,N_1527);
nand U2006 (N_2006,N_1475,N_1640);
nand U2007 (N_2007,N_1253,N_1216);
nand U2008 (N_2008,N_1600,N_1417);
and U2009 (N_2009,N_1606,N_1403);
nor U2010 (N_2010,N_1538,N_1770);
nand U2011 (N_2011,N_1470,N_1536);
and U2012 (N_2012,N_1483,N_1725);
and U2013 (N_2013,N_1618,N_1552);
xor U2014 (N_2014,N_1233,N_1316);
nor U2015 (N_2015,N_1594,N_1739);
and U2016 (N_2016,N_1206,N_1561);
or U2017 (N_2017,N_1512,N_1207);
and U2018 (N_2018,N_1318,N_1282);
or U2019 (N_2019,N_1652,N_1397);
nor U2020 (N_2020,N_1478,N_1450);
nand U2021 (N_2021,N_1221,N_1422);
nand U2022 (N_2022,N_1421,N_1583);
or U2023 (N_2023,N_1719,N_1299);
nor U2024 (N_2024,N_1733,N_1277);
xor U2025 (N_2025,N_1413,N_1592);
nor U2026 (N_2026,N_1666,N_1311);
and U2027 (N_2027,N_1224,N_1275);
or U2028 (N_2028,N_1743,N_1258);
or U2029 (N_2029,N_1551,N_1554);
or U2030 (N_2030,N_1746,N_1756);
nor U2031 (N_2031,N_1250,N_1776);
nand U2032 (N_2032,N_1763,N_1202);
nand U2033 (N_2033,N_1313,N_1336);
or U2034 (N_2034,N_1615,N_1630);
nand U2035 (N_2035,N_1682,N_1636);
or U2036 (N_2036,N_1544,N_1503);
and U2037 (N_2037,N_1513,N_1531);
or U2038 (N_2038,N_1496,N_1317);
and U2039 (N_2039,N_1268,N_1639);
nand U2040 (N_2040,N_1273,N_1660);
and U2041 (N_2041,N_1405,N_1278);
nor U2042 (N_2042,N_1562,N_1738);
nor U2043 (N_2043,N_1722,N_1377);
nand U2044 (N_2044,N_1694,N_1747);
nand U2045 (N_2045,N_1360,N_1778);
or U2046 (N_2046,N_1505,N_1416);
nand U2047 (N_2047,N_1558,N_1321);
and U2048 (N_2048,N_1780,N_1610);
nor U2049 (N_2049,N_1388,N_1290);
nor U2050 (N_2050,N_1266,N_1489);
nand U2051 (N_2051,N_1704,N_1382);
nor U2052 (N_2052,N_1297,N_1495);
or U2053 (N_2053,N_1559,N_1774);
or U2054 (N_2054,N_1218,N_1271);
nand U2055 (N_2055,N_1240,N_1357);
nand U2056 (N_2056,N_1792,N_1741);
or U2057 (N_2057,N_1381,N_1765);
nor U2058 (N_2058,N_1265,N_1431);
nor U2059 (N_2059,N_1687,N_1563);
xor U2060 (N_2060,N_1675,N_1602);
nand U2061 (N_2061,N_1644,N_1301);
and U2062 (N_2062,N_1735,N_1287);
and U2063 (N_2063,N_1332,N_1617);
and U2064 (N_2064,N_1467,N_1203);
nand U2065 (N_2065,N_1352,N_1331);
and U2066 (N_2066,N_1745,N_1737);
and U2067 (N_2067,N_1488,N_1717);
nand U2068 (N_2068,N_1292,N_1491);
and U2069 (N_2069,N_1587,N_1791);
nor U2070 (N_2070,N_1394,N_1726);
or U2071 (N_2071,N_1710,N_1354);
nand U2072 (N_2072,N_1628,N_1232);
nor U2073 (N_2073,N_1386,N_1516);
or U2074 (N_2074,N_1771,N_1319);
nand U2075 (N_2075,N_1504,N_1249);
nor U2076 (N_2076,N_1262,N_1593);
nor U2077 (N_2077,N_1477,N_1432);
and U2078 (N_2078,N_1423,N_1230);
and U2079 (N_2079,N_1246,N_1214);
nand U2080 (N_2080,N_1358,N_1235);
or U2081 (N_2081,N_1337,N_1598);
and U2082 (N_2082,N_1322,N_1300);
or U2083 (N_2083,N_1569,N_1251);
or U2084 (N_2084,N_1380,N_1720);
nand U2085 (N_2085,N_1718,N_1638);
nand U2086 (N_2086,N_1362,N_1355);
or U2087 (N_2087,N_1768,N_1723);
and U2088 (N_2088,N_1728,N_1650);
and U2089 (N_2089,N_1420,N_1608);
and U2090 (N_2090,N_1534,N_1484);
nor U2091 (N_2091,N_1433,N_1234);
and U2092 (N_2092,N_1750,N_1688);
or U2093 (N_2093,N_1542,N_1789);
nor U2094 (N_2094,N_1430,N_1759);
or U2095 (N_2095,N_1379,N_1200);
nand U2096 (N_2096,N_1764,N_1409);
nor U2097 (N_2097,N_1621,N_1343);
or U2098 (N_2098,N_1370,N_1291);
nand U2099 (N_2099,N_1556,N_1327);
nand U2100 (N_2100,N_1483,N_1319);
nand U2101 (N_2101,N_1781,N_1604);
nor U2102 (N_2102,N_1436,N_1646);
nand U2103 (N_2103,N_1236,N_1791);
and U2104 (N_2104,N_1231,N_1435);
and U2105 (N_2105,N_1666,N_1774);
and U2106 (N_2106,N_1249,N_1525);
nor U2107 (N_2107,N_1735,N_1564);
or U2108 (N_2108,N_1421,N_1784);
nor U2109 (N_2109,N_1775,N_1241);
nand U2110 (N_2110,N_1705,N_1347);
xnor U2111 (N_2111,N_1615,N_1283);
and U2112 (N_2112,N_1364,N_1473);
and U2113 (N_2113,N_1427,N_1789);
or U2114 (N_2114,N_1549,N_1661);
nor U2115 (N_2115,N_1289,N_1645);
or U2116 (N_2116,N_1752,N_1312);
and U2117 (N_2117,N_1673,N_1487);
or U2118 (N_2118,N_1367,N_1714);
nor U2119 (N_2119,N_1376,N_1563);
nand U2120 (N_2120,N_1349,N_1219);
nand U2121 (N_2121,N_1399,N_1459);
nand U2122 (N_2122,N_1559,N_1703);
nand U2123 (N_2123,N_1217,N_1692);
nor U2124 (N_2124,N_1714,N_1497);
nand U2125 (N_2125,N_1200,N_1561);
nand U2126 (N_2126,N_1693,N_1278);
and U2127 (N_2127,N_1234,N_1284);
or U2128 (N_2128,N_1342,N_1419);
nor U2129 (N_2129,N_1523,N_1411);
or U2130 (N_2130,N_1717,N_1537);
nand U2131 (N_2131,N_1554,N_1317);
nand U2132 (N_2132,N_1451,N_1771);
nor U2133 (N_2133,N_1458,N_1274);
nand U2134 (N_2134,N_1269,N_1378);
and U2135 (N_2135,N_1502,N_1298);
nand U2136 (N_2136,N_1570,N_1345);
nand U2137 (N_2137,N_1329,N_1687);
and U2138 (N_2138,N_1670,N_1287);
nor U2139 (N_2139,N_1559,N_1664);
nor U2140 (N_2140,N_1570,N_1402);
or U2141 (N_2141,N_1568,N_1669);
and U2142 (N_2142,N_1495,N_1742);
and U2143 (N_2143,N_1548,N_1513);
or U2144 (N_2144,N_1415,N_1393);
nand U2145 (N_2145,N_1622,N_1278);
nand U2146 (N_2146,N_1460,N_1333);
nand U2147 (N_2147,N_1725,N_1730);
nor U2148 (N_2148,N_1418,N_1484);
and U2149 (N_2149,N_1457,N_1730);
nand U2150 (N_2150,N_1273,N_1510);
and U2151 (N_2151,N_1447,N_1563);
xnor U2152 (N_2152,N_1351,N_1219);
nand U2153 (N_2153,N_1246,N_1234);
nor U2154 (N_2154,N_1654,N_1219);
or U2155 (N_2155,N_1242,N_1328);
or U2156 (N_2156,N_1580,N_1284);
and U2157 (N_2157,N_1233,N_1444);
nand U2158 (N_2158,N_1510,N_1723);
nor U2159 (N_2159,N_1529,N_1393);
and U2160 (N_2160,N_1248,N_1220);
nand U2161 (N_2161,N_1764,N_1217);
nor U2162 (N_2162,N_1692,N_1714);
or U2163 (N_2163,N_1244,N_1473);
nand U2164 (N_2164,N_1517,N_1777);
nand U2165 (N_2165,N_1403,N_1625);
nand U2166 (N_2166,N_1589,N_1256);
or U2167 (N_2167,N_1227,N_1453);
or U2168 (N_2168,N_1201,N_1557);
nand U2169 (N_2169,N_1610,N_1251);
or U2170 (N_2170,N_1371,N_1658);
xnor U2171 (N_2171,N_1516,N_1613);
nor U2172 (N_2172,N_1652,N_1760);
and U2173 (N_2173,N_1595,N_1714);
nand U2174 (N_2174,N_1722,N_1546);
or U2175 (N_2175,N_1294,N_1394);
nor U2176 (N_2176,N_1775,N_1353);
and U2177 (N_2177,N_1742,N_1380);
or U2178 (N_2178,N_1764,N_1613);
and U2179 (N_2179,N_1714,N_1233);
or U2180 (N_2180,N_1478,N_1243);
or U2181 (N_2181,N_1204,N_1587);
nor U2182 (N_2182,N_1410,N_1388);
nand U2183 (N_2183,N_1762,N_1350);
nand U2184 (N_2184,N_1273,N_1661);
or U2185 (N_2185,N_1314,N_1665);
or U2186 (N_2186,N_1410,N_1516);
and U2187 (N_2187,N_1513,N_1314);
or U2188 (N_2188,N_1359,N_1536);
nor U2189 (N_2189,N_1578,N_1763);
nor U2190 (N_2190,N_1656,N_1733);
xor U2191 (N_2191,N_1475,N_1490);
nand U2192 (N_2192,N_1600,N_1534);
and U2193 (N_2193,N_1761,N_1505);
or U2194 (N_2194,N_1651,N_1787);
and U2195 (N_2195,N_1502,N_1690);
nand U2196 (N_2196,N_1647,N_1562);
or U2197 (N_2197,N_1374,N_1283);
nand U2198 (N_2198,N_1498,N_1516);
nand U2199 (N_2199,N_1211,N_1382);
nand U2200 (N_2200,N_1754,N_1314);
and U2201 (N_2201,N_1213,N_1216);
or U2202 (N_2202,N_1740,N_1523);
or U2203 (N_2203,N_1560,N_1271);
nand U2204 (N_2204,N_1206,N_1443);
or U2205 (N_2205,N_1392,N_1686);
nand U2206 (N_2206,N_1734,N_1633);
nor U2207 (N_2207,N_1685,N_1692);
and U2208 (N_2208,N_1379,N_1588);
or U2209 (N_2209,N_1272,N_1226);
or U2210 (N_2210,N_1595,N_1664);
and U2211 (N_2211,N_1297,N_1520);
and U2212 (N_2212,N_1247,N_1470);
or U2213 (N_2213,N_1210,N_1423);
nand U2214 (N_2214,N_1758,N_1330);
or U2215 (N_2215,N_1610,N_1781);
nor U2216 (N_2216,N_1252,N_1341);
nor U2217 (N_2217,N_1392,N_1226);
nor U2218 (N_2218,N_1641,N_1273);
nand U2219 (N_2219,N_1681,N_1722);
or U2220 (N_2220,N_1278,N_1785);
nand U2221 (N_2221,N_1705,N_1321);
and U2222 (N_2222,N_1409,N_1239);
nand U2223 (N_2223,N_1344,N_1625);
nand U2224 (N_2224,N_1611,N_1568);
or U2225 (N_2225,N_1482,N_1724);
and U2226 (N_2226,N_1255,N_1645);
and U2227 (N_2227,N_1556,N_1639);
nand U2228 (N_2228,N_1237,N_1468);
or U2229 (N_2229,N_1736,N_1659);
and U2230 (N_2230,N_1235,N_1317);
nor U2231 (N_2231,N_1701,N_1748);
and U2232 (N_2232,N_1577,N_1414);
nand U2233 (N_2233,N_1492,N_1544);
nand U2234 (N_2234,N_1645,N_1441);
and U2235 (N_2235,N_1621,N_1214);
and U2236 (N_2236,N_1279,N_1645);
nand U2237 (N_2237,N_1268,N_1421);
nand U2238 (N_2238,N_1650,N_1544);
or U2239 (N_2239,N_1278,N_1269);
nand U2240 (N_2240,N_1607,N_1224);
nor U2241 (N_2241,N_1446,N_1473);
nand U2242 (N_2242,N_1594,N_1292);
nor U2243 (N_2243,N_1717,N_1262);
nand U2244 (N_2244,N_1597,N_1302);
nand U2245 (N_2245,N_1308,N_1411);
and U2246 (N_2246,N_1372,N_1427);
nand U2247 (N_2247,N_1773,N_1575);
nand U2248 (N_2248,N_1788,N_1376);
and U2249 (N_2249,N_1631,N_1618);
nor U2250 (N_2250,N_1515,N_1452);
or U2251 (N_2251,N_1212,N_1517);
nand U2252 (N_2252,N_1674,N_1689);
nor U2253 (N_2253,N_1440,N_1449);
nor U2254 (N_2254,N_1773,N_1359);
nand U2255 (N_2255,N_1761,N_1568);
or U2256 (N_2256,N_1552,N_1787);
nor U2257 (N_2257,N_1650,N_1513);
nand U2258 (N_2258,N_1604,N_1203);
nand U2259 (N_2259,N_1604,N_1750);
and U2260 (N_2260,N_1274,N_1495);
nor U2261 (N_2261,N_1313,N_1782);
nor U2262 (N_2262,N_1310,N_1499);
nor U2263 (N_2263,N_1482,N_1423);
and U2264 (N_2264,N_1270,N_1544);
nor U2265 (N_2265,N_1448,N_1677);
and U2266 (N_2266,N_1410,N_1219);
nand U2267 (N_2267,N_1337,N_1649);
nor U2268 (N_2268,N_1610,N_1554);
nand U2269 (N_2269,N_1331,N_1639);
nor U2270 (N_2270,N_1574,N_1617);
and U2271 (N_2271,N_1790,N_1664);
and U2272 (N_2272,N_1714,N_1377);
nor U2273 (N_2273,N_1640,N_1558);
nand U2274 (N_2274,N_1760,N_1268);
and U2275 (N_2275,N_1236,N_1761);
and U2276 (N_2276,N_1582,N_1225);
and U2277 (N_2277,N_1278,N_1410);
and U2278 (N_2278,N_1372,N_1513);
or U2279 (N_2279,N_1761,N_1339);
nor U2280 (N_2280,N_1438,N_1363);
nand U2281 (N_2281,N_1425,N_1613);
nor U2282 (N_2282,N_1393,N_1761);
nor U2283 (N_2283,N_1549,N_1228);
or U2284 (N_2284,N_1706,N_1783);
nor U2285 (N_2285,N_1336,N_1375);
nor U2286 (N_2286,N_1616,N_1438);
nor U2287 (N_2287,N_1274,N_1288);
nand U2288 (N_2288,N_1752,N_1570);
or U2289 (N_2289,N_1574,N_1758);
nand U2290 (N_2290,N_1380,N_1469);
or U2291 (N_2291,N_1549,N_1730);
nand U2292 (N_2292,N_1717,N_1628);
nor U2293 (N_2293,N_1328,N_1653);
and U2294 (N_2294,N_1490,N_1764);
nor U2295 (N_2295,N_1359,N_1381);
and U2296 (N_2296,N_1742,N_1357);
and U2297 (N_2297,N_1221,N_1402);
nor U2298 (N_2298,N_1595,N_1617);
nand U2299 (N_2299,N_1235,N_1302);
nand U2300 (N_2300,N_1698,N_1206);
xor U2301 (N_2301,N_1572,N_1751);
nand U2302 (N_2302,N_1757,N_1455);
nand U2303 (N_2303,N_1389,N_1219);
nor U2304 (N_2304,N_1365,N_1450);
and U2305 (N_2305,N_1222,N_1652);
xnor U2306 (N_2306,N_1237,N_1783);
and U2307 (N_2307,N_1347,N_1537);
and U2308 (N_2308,N_1597,N_1792);
xnor U2309 (N_2309,N_1516,N_1361);
or U2310 (N_2310,N_1470,N_1258);
and U2311 (N_2311,N_1285,N_1327);
nor U2312 (N_2312,N_1385,N_1568);
and U2313 (N_2313,N_1202,N_1787);
or U2314 (N_2314,N_1663,N_1435);
or U2315 (N_2315,N_1389,N_1490);
or U2316 (N_2316,N_1720,N_1721);
or U2317 (N_2317,N_1475,N_1295);
or U2318 (N_2318,N_1372,N_1485);
nand U2319 (N_2319,N_1257,N_1729);
nor U2320 (N_2320,N_1451,N_1227);
or U2321 (N_2321,N_1774,N_1459);
or U2322 (N_2322,N_1625,N_1463);
nand U2323 (N_2323,N_1419,N_1393);
nor U2324 (N_2324,N_1209,N_1747);
nand U2325 (N_2325,N_1627,N_1397);
nor U2326 (N_2326,N_1695,N_1330);
and U2327 (N_2327,N_1265,N_1329);
nand U2328 (N_2328,N_1608,N_1414);
nor U2329 (N_2329,N_1503,N_1478);
nor U2330 (N_2330,N_1756,N_1552);
nor U2331 (N_2331,N_1405,N_1660);
and U2332 (N_2332,N_1554,N_1791);
nand U2333 (N_2333,N_1680,N_1445);
nand U2334 (N_2334,N_1267,N_1760);
or U2335 (N_2335,N_1521,N_1362);
or U2336 (N_2336,N_1317,N_1428);
and U2337 (N_2337,N_1670,N_1515);
nand U2338 (N_2338,N_1347,N_1513);
nor U2339 (N_2339,N_1677,N_1512);
or U2340 (N_2340,N_1656,N_1316);
or U2341 (N_2341,N_1437,N_1266);
nor U2342 (N_2342,N_1454,N_1219);
nand U2343 (N_2343,N_1329,N_1608);
nor U2344 (N_2344,N_1400,N_1271);
nor U2345 (N_2345,N_1502,N_1390);
nor U2346 (N_2346,N_1552,N_1398);
and U2347 (N_2347,N_1668,N_1412);
or U2348 (N_2348,N_1694,N_1468);
and U2349 (N_2349,N_1404,N_1427);
nor U2350 (N_2350,N_1332,N_1588);
or U2351 (N_2351,N_1494,N_1417);
nand U2352 (N_2352,N_1275,N_1394);
and U2353 (N_2353,N_1470,N_1571);
and U2354 (N_2354,N_1514,N_1560);
and U2355 (N_2355,N_1313,N_1511);
nor U2356 (N_2356,N_1631,N_1375);
nand U2357 (N_2357,N_1764,N_1415);
or U2358 (N_2358,N_1783,N_1740);
nand U2359 (N_2359,N_1290,N_1457);
nor U2360 (N_2360,N_1600,N_1627);
nor U2361 (N_2361,N_1741,N_1798);
nand U2362 (N_2362,N_1503,N_1527);
nor U2363 (N_2363,N_1417,N_1794);
nor U2364 (N_2364,N_1302,N_1303);
and U2365 (N_2365,N_1649,N_1630);
nand U2366 (N_2366,N_1516,N_1539);
nand U2367 (N_2367,N_1492,N_1503);
or U2368 (N_2368,N_1649,N_1790);
xnor U2369 (N_2369,N_1781,N_1659);
and U2370 (N_2370,N_1294,N_1473);
nor U2371 (N_2371,N_1466,N_1381);
and U2372 (N_2372,N_1553,N_1510);
and U2373 (N_2373,N_1739,N_1511);
nand U2374 (N_2374,N_1326,N_1321);
nor U2375 (N_2375,N_1578,N_1430);
or U2376 (N_2376,N_1269,N_1523);
or U2377 (N_2377,N_1658,N_1569);
or U2378 (N_2378,N_1527,N_1299);
or U2379 (N_2379,N_1313,N_1636);
or U2380 (N_2380,N_1239,N_1785);
nand U2381 (N_2381,N_1348,N_1681);
or U2382 (N_2382,N_1374,N_1767);
or U2383 (N_2383,N_1611,N_1363);
nand U2384 (N_2384,N_1547,N_1767);
nor U2385 (N_2385,N_1269,N_1797);
nor U2386 (N_2386,N_1318,N_1692);
nand U2387 (N_2387,N_1769,N_1751);
and U2388 (N_2388,N_1209,N_1454);
and U2389 (N_2389,N_1501,N_1704);
nor U2390 (N_2390,N_1308,N_1529);
and U2391 (N_2391,N_1683,N_1417);
and U2392 (N_2392,N_1486,N_1387);
nand U2393 (N_2393,N_1473,N_1309);
and U2394 (N_2394,N_1555,N_1335);
or U2395 (N_2395,N_1595,N_1651);
xor U2396 (N_2396,N_1623,N_1425);
and U2397 (N_2397,N_1606,N_1332);
nor U2398 (N_2398,N_1201,N_1712);
or U2399 (N_2399,N_1276,N_1631);
or U2400 (N_2400,N_2222,N_1935);
and U2401 (N_2401,N_1821,N_2199);
or U2402 (N_2402,N_2015,N_2078);
nor U2403 (N_2403,N_2122,N_2289);
nor U2404 (N_2404,N_2027,N_2206);
or U2405 (N_2405,N_1995,N_2159);
or U2406 (N_2406,N_2371,N_1964);
nand U2407 (N_2407,N_2165,N_2195);
and U2408 (N_2408,N_1979,N_1846);
nor U2409 (N_2409,N_2064,N_1997);
and U2410 (N_2410,N_2103,N_1887);
and U2411 (N_2411,N_1963,N_2197);
or U2412 (N_2412,N_1880,N_2291);
or U2413 (N_2413,N_2353,N_2076);
or U2414 (N_2414,N_2178,N_2233);
nand U2415 (N_2415,N_2226,N_2342);
and U2416 (N_2416,N_1833,N_2272);
nor U2417 (N_2417,N_2120,N_2336);
nor U2418 (N_2418,N_2287,N_2067);
or U2419 (N_2419,N_1952,N_1975);
and U2420 (N_2420,N_1911,N_1940);
or U2421 (N_2421,N_2166,N_1917);
nor U2422 (N_2422,N_1897,N_2304);
or U2423 (N_2423,N_2100,N_1898);
or U2424 (N_2424,N_2230,N_1934);
or U2425 (N_2425,N_2388,N_2218);
nor U2426 (N_2426,N_2024,N_2071);
xor U2427 (N_2427,N_2126,N_2098);
nor U2428 (N_2428,N_2363,N_2247);
xnor U2429 (N_2429,N_2217,N_2032);
nand U2430 (N_2430,N_1852,N_2297);
nand U2431 (N_2431,N_2338,N_2393);
or U2432 (N_2432,N_1959,N_2150);
nor U2433 (N_2433,N_2055,N_2250);
nor U2434 (N_2434,N_2174,N_2106);
nand U2435 (N_2435,N_2257,N_2021);
or U2436 (N_2436,N_1892,N_2048);
nor U2437 (N_2437,N_2321,N_2181);
or U2438 (N_2438,N_2210,N_2031);
nor U2439 (N_2439,N_2141,N_2331);
and U2440 (N_2440,N_2223,N_2278);
xor U2441 (N_2441,N_2244,N_2175);
or U2442 (N_2442,N_2158,N_1907);
nor U2443 (N_2443,N_1908,N_2253);
and U2444 (N_2444,N_2144,N_1973);
nand U2445 (N_2445,N_2288,N_2377);
and U2446 (N_2446,N_2299,N_1832);
nor U2447 (N_2447,N_2203,N_1903);
nand U2448 (N_2448,N_1800,N_2315);
and U2449 (N_2449,N_2344,N_2038);
nor U2450 (N_2450,N_2266,N_1841);
nor U2451 (N_2451,N_2354,N_2105);
or U2452 (N_2452,N_2273,N_2161);
or U2453 (N_2453,N_2219,N_2232);
and U2454 (N_2454,N_2317,N_2379);
nor U2455 (N_2455,N_2039,N_1877);
or U2456 (N_2456,N_2019,N_1885);
or U2457 (N_2457,N_1828,N_2059);
nand U2458 (N_2458,N_1976,N_2115);
nand U2459 (N_2459,N_2153,N_1894);
nor U2460 (N_2460,N_2119,N_2137);
nand U2461 (N_2461,N_2383,N_2325);
and U2462 (N_2462,N_1998,N_1807);
or U2463 (N_2463,N_2054,N_1891);
nor U2464 (N_2464,N_2104,N_2111);
nor U2465 (N_2465,N_1947,N_2014);
and U2466 (N_2466,N_2235,N_2157);
nor U2467 (N_2467,N_2337,N_2227);
and U2468 (N_2468,N_2028,N_2171);
nand U2469 (N_2469,N_1856,N_2349);
and U2470 (N_2470,N_2183,N_1834);
and U2471 (N_2471,N_2148,N_1817);
nor U2472 (N_2472,N_1915,N_2134);
nor U2473 (N_2473,N_1905,N_1912);
nand U2474 (N_2474,N_1888,N_2369);
and U2475 (N_2475,N_1968,N_2225);
nor U2476 (N_2476,N_2351,N_1837);
and U2477 (N_2477,N_2163,N_2138);
and U2478 (N_2478,N_2298,N_2083);
nor U2479 (N_2479,N_2370,N_2186);
nor U2480 (N_2480,N_2133,N_2339);
nand U2481 (N_2481,N_2282,N_1902);
nor U2482 (N_2482,N_2312,N_2259);
or U2483 (N_2483,N_2075,N_1803);
nor U2484 (N_2484,N_2389,N_1873);
and U2485 (N_2485,N_2112,N_2207);
or U2486 (N_2486,N_2302,N_2306);
and U2487 (N_2487,N_1802,N_2065);
nand U2488 (N_2488,N_2080,N_1849);
and U2489 (N_2489,N_2135,N_2283);
nand U2490 (N_2490,N_2069,N_2290);
nor U2491 (N_2491,N_2011,N_2292);
or U2492 (N_2492,N_1906,N_1881);
or U2493 (N_2493,N_1999,N_2238);
or U2494 (N_2494,N_2193,N_2058);
nor U2495 (N_2495,N_1941,N_2117);
nor U2496 (N_2496,N_1960,N_2356);
nor U2497 (N_2497,N_2018,N_1890);
nand U2498 (N_2498,N_2375,N_2001);
nand U2499 (N_2499,N_2180,N_1962);
and U2500 (N_2500,N_2177,N_2258);
nand U2501 (N_2501,N_2160,N_1814);
and U2502 (N_2502,N_2307,N_2086);
and U2503 (N_2503,N_2154,N_2102);
or U2504 (N_2504,N_1801,N_2284);
nand U2505 (N_2505,N_2124,N_2364);
or U2506 (N_2506,N_2114,N_2190);
xnor U2507 (N_2507,N_2256,N_2125);
or U2508 (N_2508,N_2305,N_2034);
nand U2509 (N_2509,N_1991,N_2323);
nand U2510 (N_2510,N_1830,N_2335);
or U2511 (N_2511,N_2037,N_1904);
and U2512 (N_2512,N_2345,N_2254);
nand U2513 (N_2513,N_2139,N_2322);
nand U2514 (N_2514,N_2151,N_2188);
nor U2515 (N_2515,N_1989,N_1818);
nand U2516 (N_2516,N_2116,N_2172);
nand U2517 (N_2517,N_2264,N_1992);
nor U2518 (N_2518,N_1919,N_1838);
nor U2519 (N_2519,N_1861,N_2044);
nand U2520 (N_2520,N_1859,N_2189);
nand U2521 (N_2521,N_2090,N_2185);
nor U2522 (N_2522,N_2033,N_1813);
nand U2523 (N_2523,N_2212,N_2234);
nor U2524 (N_2524,N_2187,N_2070);
nor U2525 (N_2525,N_2316,N_2168);
and U2526 (N_2526,N_1874,N_2211);
and U2527 (N_2527,N_2201,N_2358);
and U2528 (N_2528,N_1878,N_2300);
or U2529 (N_2529,N_2333,N_2382);
nor U2530 (N_2530,N_2062,N_2167);
or U2531 (N_2531,N_2346,N_2350);
nand U2532 (N_2532,N_2255,N_1932);
or U2533 (N_2533,N_1825,N_1965);
nand U2534 (N_2534,N_1848,N_2368);
nand U2535 (N_2535,N_1827,N_2143);
or U2536 (N_2536,N_1842,N_1931);
nand U2537 (N_2537,N_2216,N_1980);
nor U2538 (N_2538,N_2051,N_1951);
nand U2539 (N_2539,N_2087,N_1829);
or U2540 (N_2540,N_2152,N_2142);
nand U2541 (N_2541,N_1996,N_1922);
nand U2542 (N_2542,N_1820,N_2136);
and U2543 (N_2543,N_2009,N_1847);
nor U2544 (N_2544,N_2396,N_1809);
nor U2545 (N_2545,N_2023,N_1851);
xnor U2546 (N_2546,N_2194,N_1805);
or U2547 (N_2547,N_2251,N_1966);
or U2548 (N_2548,N_2052,N_2224);
and U2549 (N_2549,N_2229,N_2343);
or U2550 (N_2550,N_2249,N_1916);
or U2551 (N_2551,N_2156,N_1871);
nor U2552 (N_2552,N_2005,N_2274);
and U2553 (N_2553,N_2096,N_1839);
and U2554 (N_2554,N_1853,N_2332);
nand U2555 (N_2555,N_2314,N_1987);
and U2556 (N_2556,N_1985,N_2089);
and U2557 (N_2557,N_2221,N_1938);
nand U2558 (N_2558,N_2360,N_1921);
nand U2559 (N_2559,N_1854,N_2241);
xnor U2560 (N_2560,N_1860,N_1896);
nand U2561 (N_2561,N_1981,N_2286);
and U2562 (N_2562,N_1812,N_2097);
and U2563 (N_2563,N_1901,N_2170);
nand U2564 (N_2564,N_1886,N_1819);
nor U2565 (N_2565,N_1993,N_2365);
nand U2566 (N_2566,N_1977,N_2285);
nor U2567 (N_2567,N_2085,N_2169);
nand U2568 (N_2568,N_2155,N_2303);
nand U2569 (N_2569,N_1953,N_2237);
or U2570 (N_2570,N_1969,N_1930);
and U2571 (N_2571,N_1806,N_2262);
nand U2572 (N_2572,N_1864,N_2056);
and U2573 (N_2573,N_2081,N_2109);
nor U2574 (N_2574,N_1900,N_2099);
or U2575 (N_2575,N_2327,N_1899);
nand U2576 (N_2576,N_2318,N_2091);
or U2577 (N_2577,N_2367,N_2003);
or U2578 (N_2578,N_2328,N_1811);
nor U2579 (N_2579,N_2362,N_2029);
nor U2580 (N_2580,N_2072,N_2392);
nor U2581 (N_2581,N_2025,N_2094);
nor U2582 (N_2582,N_2295,N_2118);
and U2583 (N_2583,N_1937,N_2095);
nor U2584 (N_2584,N_2068,N_2129);
and U2585 (N_2585,N_2004,N_1868);
nor U2586 (N_2586,N_2036,N_1843);
nor U2587 (N_2587,N_2202,N_2228);
nor U2588 (N_2588,N_2215,N_2010);
or U2589 (N_2589,N_1855,N_2042);
nand U2590 (N_2590,N_1914,N_1928);
or U2591 (N_2591,N_1869,N_2397);
nand U2592 (N_2592,N_1982,N_2270);
nor U2593 (N_2593,N_2173,N_1990);
nor U2594 (N_2594,N_2366,N_2309);
and U2595 (N_2595,N_1946,N_2191);
or U2596 (N_2596,N_2121,N_2016);
nand U2597 (N_2597,N_2209,N_2061);
or U2598 (N_2598,N_2008,N_2130);
nand U2599 (N_2599,N_2340,N_1920);
or U2600 (N_2600,N_1927,N_1956);
nand U2601 (N_2601,N_2162,N_2146);
or U2602 (N_2602,N_2088,N_1824);
nor U2603 (N_2603,N_2386,N_2341);
nor U2604 (N_2604,N_2108,N_2113);
nor U2605 (N_2605,N_2239,N_2220);
and U2606 (N_2606,N_2192,N_1823);
xor U2607 (N_2607,N_1961,N_2236);
nand U2608 (N_2608,N_2063,N_2140);
and U2609 (N_2609,N_2208,N_1836);
and U2610 (N_2610,N_1986,N_2301);
and U2611 (N_2611,N_1988,N_2231);
or U2612 (N_2612,N_2084,N_2006);
nand U2613 (N_2613,N_2296,N_2394);
nand U2614 (N_2614,N_2352,N_2281);
nand U2615 (N_2615,N_2007,N_2271);
and U2616 (N_2616,N_1967,N_1955);
or U2617 (N_2617,N_1876,N_1948);
nor U2618 (N_2618,N_1895,N_1943);
xnor U2619 (N_2619,N_1865,N_2050);
or U2620 (N_2620,N_2204,N_2280);
nor U2621 (N_2621,N_1850,N_2313);
and U2622 (N_2622,N_2261,N_2387);
or U2623 (N_2623,N_2391,N_2012);
nor U2624 (N_2624,N_2355,N_2373);
nand U2625 (N_2625,N_2110,N_1984);
nor U2626 (N_2626,N_1808,N_1972);
or U2627 (N_2627,N_2045,N_2214);
or U2628 (N_2628,N_2378,N_2348);
nand U2629 (N_2629,N_1858,N_2049);
and U2630 (N_2630,N_2310,N_1862);
nand U2631 (N_2631,N_1867,N_2380);
and U2632 (N_2632,N_2361,N_2182);
or U2633 (N_2633,N_2205,N_1857);
nor U2634 (N_2634,N_2057,N_1910);
or U2635 (N_2635,N_2093,N_1816);
nor U2636 (N_2636,N_2176,N_1870);
nor U2637 (N_2637,N_1913,N_1944);
nand U2638 (N_2638,N_2147,N_1909);
and U2639 (N_2639,N_1844,N_2243);
nor U2640 (N_2640,N_2041,N_2268);
or U2641 (N_2641,N_2079,N_2082);
or U2642 (N_2642,N_2017,N_2060);
nor U2643 (N_2643,N_2242,N_1840);
and U2644 (N_2644,N_2040,N_2320);
nor U2645 (N_2645,N_1923,N_2252);
nor U2646 (N_2646,N_1974,N_2043);
and U2647 (N_2647,N_1866,N_2213);
and U2648 (N_2648,N_1936,N_1958);
nand U2649 (N_2649,N_2319,N_1942);
xnor U2650 (N_2650,N_2184,N_2030);
nand U2651 (N_2651,N_1957,N_2077);
and U2652 (N_2652,N_1845,N_1971);
nand U2653 (N_2653,N_1822,N_2246);
nor U2654 (N_2654,N_1926,N_1978);
nand U2655 (N_2655,N_2020,N_2390);
nand U2656 (N_2656,N_1882,N_1918);
nand U2657 (N_2657,N_2053,N_1893);
nand U2658 (N_2658,N_2293,N_2276);
nor U2659 (N_2659,N_2046,N_2013);
and U2660 (N_2660,N_2308,N_1970);
and U2661 (N_2661,N_2198,N_2399);
nor U2662 (N_2662,N_1815,N_1835);
and U2663 (N_2663,N_2260,N_2334);
and U2664 (N_2664,N_2145,N_1884);
and U2665 (N_2665,N_2132,N_2240);
and U2666 (N_2666,N_2372,N_2330);
and U2667 (N_2667,N_2279,N_2179);
or U2668 (N_2668,N_2269,N_2398);
or U2669 (N_2669,N_2164,N_2376);
nand U2670 (N_2670,N_1883,N_2277);
nand U2671 (N_2671,N_2275,N_2128);
nor U2672 (N_2672,N_2347,N_1810);
nand U2673 (N_2673,N_2357,N_2395);
or U2674 (N_2674,N_2245,N_1804);
or U2675 (N_2675,N_2294,N_1954);
nand U2676 (N_2676,N_1831,N_1826);
or U2677 (N_2677,N_2374,N_1950);
nand U2678 (N_2678,N_2196,N_1929);
nand U2679 (N_2679,N_2359,N_2101);
and U2680 (N_2680,N_2248,N_2000);
xnor U2681 (N_2681,N_2047,N_2263);
and U2682 (N_2682,N_2107,N_1945);
nand U2683 (N_2683,N_1983,N_2022);
or U2684 (N_2684,N_1879,N_1994);
nor U2685 (N_2685,N_2073,N_2267);
or U2686 (N_2686,N_2384,N_2127);
nand U2687 (N_2687,N_2002,N_2324);
and U2688 (N_2688,N_2035,N_1875);
and U2689 (N_2689,N_2026,N_1949);
nor U2690 (N_2690,N_1872,N_2074);
or U2691 (N_2691,N_2131,N_1889);
xnor U2692 (N_2692,N_2385,N_2092);
nor U2693 (N_2693,N_2326,N_2066);
nor U2694 (N_2694,N_2149,N_2200);
nor U2695 (N_2695,N_2123,N_2329);
xnor U2696 (N_2696,N_1933,N_1939);
and U2697 (N_2697,N_2265,N_1863);
nand U2698 (N_2698,N_2381,N_1924);
or U2699 (N_2699,N_1925,N_2311);
and U2700 (N_2700,N_1836,N_2191);
nand U2701 (N_2701,N_1948,N_1986);
or U2702 (N_2702,N_2059,N_1959);
nor U2703 (N_2703,N_2145,N_2245);
nand U2704 (N_2704,N_2322,N_2182);
nand U2705 (N_2705,N_2030,N_2198);
nor U2706 (N_2706,N_2352,N_2136);
or U2707 (N_2707,N_1836,N_1824);
nor U2708 (N_2708,N_1989,N_1926);
nor U2709 (N_2709,N_1948,N_2358);
nor U2710 (N_2710,N_2117,N_2100);
nor U2711 (N_2711,N_1948,N_2184);
nand U2712 (N_2712,N_1902,N_2015);
or U2713 (N_2713,N_2297,N_1916);
nor U2714 (N_2714,N_2172,N_1941);
or U2715 (N_2715,N_2384,N_2099);
nor U2716 (N_2716,N_1845,N_1933);
and U2717 (N_2717,N_2271,N_2335);
nand U2718 (N_2718,N_2052,N_2393);
and U2719 (N_2719,N_2330,N_2257);
and U2720 (N_2720,N_1994,N_2140);
and U2721 (N_2721,N_1933,N_1912);
or U2722 (N_2722,N_1879,N_1866);
nand U2723 (N_2723,N_2203,N_2383);
nor U2724 (N_2724,N_2366,N_1891);
xor U2725 (N_2725,N_2083,N_2220);
or U2726 (N_2726,N_2283,N_1939);
or U2727 (N_2727,N_2269,N_2116);
nand U2728 (N_2728,N_1928,N_1926);
and U2729 (N_2729,N_2278,N_2344);
and U2730 (N_2730,N_2010,N_2378);
and U2731 (N_2731,N_2185,N_1810);
nand U2732 (N_2732,N_1976,N_1964);
nor U2733 (N_2733,N_2076,N_2272);
nor U2734 (N_2734,N_2355,N_2296);
nor U2735 (N_2735,N_2146,N_2273);
nor U2736 (N_2736,N_2253,N_2089);
and U2737 (N_2737,N_2226,N_1906);
nand U2738 (N_2738,N_2162,N_2180);
and U2739 (N_2739,N_1807,N_2144);
and U2740 (N_2740,N_2346,N_2244);
nand U2741 (N_2741,N_2036,N_2181);
nor U2742 (N_2742,N_2066,N_1819);
nand U2743 (N_2743,N_1820,N_1858);
nor U2744 (N_2744,N_2216,N_2117);
or U2745 (N_2745,N_1904,N_1963);
nand U2746 (N_2746,N_2059,N_2258);
or U2747 (N_2747,N_1923,N_2069);
nand U2748 (N_2748,N_2175,N_2209);
nor U2749 (N_2749,N_1844,N_2372);
and U2750 (N_2750,N_2003,N_1831);
or U2751 (N_2751,N_1928,N_1808);
nor U2752 (N_2752,N_2293,N_1870);
xor U2753 (N_2753,N_2027,N_2151);
or U2754 (N_2754,N_2382,N_1860);
nor U2755 (N_2755,N_2375,N_1855);
nand U2756 (N_2756,N_2080,N_1867);
nand U2757 (N_2757,N_2100,N_1957);
nand U2758 (N_2758,N_1963,N_1818);
and U2759 (N_2759,N_1984,N_2108);
nor U2760 (N_2760,N_2139,N_2173);
and U2761 (N_2761,N_2246,N_1877);
xor U2762 (N_2762,N_2359,N_1801);
nand U2763 (N_2763,N_2275,N_2022);
nand U2764 (N_2764,N_2239,N_1963);
xnor U2765 (N_2765,N_2181,N_1917);
nor U2766 (N_2766,N_2137,N_1919);
and U2767 (N_2767,N_2161,N_1997);
nor U2768 (N_2768,N_1881,N_1930);
nand U2769 (N_2769,N_2221,N_1841);
or U2770 (N_2770,N_2330,N_2198);
or U2771 (N_2771,N_2034,N_2129);
nand U2772 (N_2772,N_1906,N_2166);
nor U2773 (N_2773,N_1863,N_1956);
or U2774 (N_2774,N_2090,N_1978);
nor U2775 (N_2775,N_1865,N_2358);
and U2776 (N_2776,N_1979,N_2301);
or U2777 (N_2777,N_2052,N_2213);
nand U2778 (N_2778,N_2006,N_2115);
nand U2779 (N_2779,N_2041,N_2126);
and U2780 (N_2780,N_2287,N_2205);
or U2781 (N_2781,N_2347,N_1898);
xor U2782 (N_2782,N_2008,N_1861);
nand U2783 (N_2783,N_1801,N_2076);
or U2784 (N_2784,N_2160,N_2096);
or U2785 (N_2785,N_2087,N_1901);
nor U2786 (N_2786,N_1841,N_1942);
and U2787 (N_2787,N_2221,N_2042);
nand U2788 (N_2788,N_2230,N_2256);
nand U2789 (N_2789,N_2333,N_2176);
or U2790 (N_2790,N_1909,N_2027);
nand U2791 (N_2791,N_2068,N_2057);
nor U2792 (N_2792,N_2214,N_2244);
nor U2793 (N_2793,N_2057,N_2356);
and U2794 (N_2794,N_2284,N_2029);
nand U2795 (N_2795,N_2365,N_1954);
and U2796 (N_2796,N_2230,N_1901);
and U2797 (N_2797,N_2062,N_2182);
nand U2798 (N_2798,N_1949,N_2277);
or U2799 (N_2799,N_2285,N_1948);
and U2800 (N_2800,N_2195,N_2013);
or U2801 (N_2801,N_1845,N_2235);
xnor U2802 (N_2802,N_1914,N_2292);
and U2803 (N_2803,N_2099,N_2212);
and U2804 (N_2804,N_2086,N_1971);
nand U2805 (N_2805,N_2232,N_2039);
nand U2806 (N_2806,N_2300,N_1830);
or U2807 (N_2807,N_2239,N_2040);
and U2808 (N_2808,N_1808,N_1945);
nor U2809 (N_2809,N_2379,N_2391);
nor U2810 (N_2810,N_2347,N_2112);
nand U2811 (N_2811,N_2093,N_2030);
nand U2812 (N_2812,N_2153,N_1980);
nand U2813 (N_2813,N_2244,N_2267);
and U2814 (N_2814,N_2390,N_2120);
or U2815 (N_2815,N_2362,N_1857);
or U2816 (N_2816,N_2165,N_1931);
nand U2817 (N_2817,N_2280,N_2178);
and U2818 (N_2818,N_2225,N_2268);
nor U2819 (N_2819,N_2311,N_1833);
nand U2820 (N_2820,N_2285,N_1854);
or U2821 (N_2821,N_2074,N_1929);
nor U2822 (N_2822,N_2321,N_1904);
or U2823 (N_2823,N_1866,N_1979);
nand U2824 (N_2824,N_1986,N_1882);
or U2825 (N_2825,N_2387,N_2253);
and U2826 (N_2826,N_2170,N_2238);
and U2827 (N_2827,N_2278,N_2256);
and U2828 (N_2828,N_2048,N_2325);
nor U2829 (N_2829,N_2001,N_2077);
and U2830 (N_2830,N_1801,N_1917);
nor U2831 (N_2831,N_2160,N_1854);
or U2832 (N_2832,N_1808,N_2263);
nor U2833 (N_2833,N_2291,N_2271);
nand U2834 (N_2834,N_2346,N_1901);
nand U2835 (N_2835,N_2054,N_2068);
xnor U2836 (N_2836,N_2299,N_1896);
nor U2837 (N_2837,N_2371,N_1898);
nand U2838 (N_2838,N_1882,N_2213);
or U2839 (N_2839,N_2148,N_1833);
nor U2840 (N_2840,N_2013,N_2059);
nand U2841 (N_2841,N_2314,N_2080);
and U2842 (N_2842,N_2114,N_2374);
and U2843 (N_2843,N_2245,N_1886);
nand U2844 (N_2844,N_2165,N_2325);
nor U2845 (N_2845,N_2287,N_2076);
or U2846 (N_2846,N_2299,N_2052);
and U2847 (N_2847,N_2128,N_2127);
or U2848 (N_2848,N_2153,N_2325);
nand U2849 (N_2849,N_2379,N_1833);
nand U2850 (N_2850,N_2282,N_1984);
or U2851 (N_2851,N_2087,N_2134);
or U2852 (N_2852,N_2013,N_1879);
nand U2853 (N_2853,N_2135,N_2012);
nor U2854 (N_2854,N_2300,N_2190);
nand U2855 (N_2855,N_2143,N_1877);
and U2856 (N_2856,N_2380,N_1923);
or U2857 (N_2857,N_2082,N_1845);
and U2858 (N_2858,N_1963,N_2334);
or U2859 (N_2859,N_2016,N_1819);
nor U2860 (N_2860,N_2152,N_2226);
nand U2861 (N_2861,N_2083,N_2053);
or U2862 (N_2862,N_2372,N_1872);
or U2863 (N_2863,N_2141,N_2205);
and U2864 (N_2864,N_2273,N_2193);
nor U2865 (N_2865,N_1854,N_2375);
nand U2866 (N_2866,N_2369,N_2063);
nor U2867 (N_2867,N_1985,N_1997);
nand U2868 (N_2868,N_2381,N_1999);
and U2869 (N_2869,N_2303,N_1981);
nor U2870 (N_2870,N_1861,N_1900);
and U2871 (N_2871,N_1838,N_2334);
and U2872 (N_2872,N_1825,N_2052);
nand U2873 (N_2873,N_2113,N_1837);
nor U2874 (N_2874,N_2012,N_1956);
and U2875 (N_2875,N_1810,N_1949);
nand U2876 (N_2876,N_2311,N_2172);
or U2877 (N_2877,N_1800,N_2022);
or U2878 (N_2878,N_2334,N_1801);
nand U2879 (N_2879,N_1888,N_2376);
xnor U2880 (N_2880,N_1951,N_2367);
nand U2881 (N_2881,N_1825,N_2208);
nand U2882 (N_2882,N_1970,N_1997);
or U2883 (N_2883,N_1808,N_2358);
nand U2884 (N_2884,N_1954,N_1847);
nand U2885 (N_2885,N_2253,N_1813);
xor U2886 (N_2886,N_2025,N_2204);
or U2887 (N_2887,N_1869,N_2323);
nor U2888 (N_2888,N_1997,N_1829);
nand U2889 (N_2889,N_2148,N_2262);
nor U2890 (N_2890,N_1822,N_2148);
or U2891 (N_2891,N_1896,N_1871);
and U2892 (N_2892,N_1907,N_2033);
nand U2893 (N_2893,N_1837,N_2188);
and U2894 (N_2894,N_2282,N_2161);
and U2895 (N_2895,N_1801,N_2221);
and U2896 (N_2896,N_2025,N_1935);
nor U2897 (N_2897,N_2251,N_1871);
nor U2898 (N_2898,N_2249,N_1999);
nor U2899 (N_2899,N_2368,N_2266);
and U2900 (N_2900,N_2115,N_1955);
and U2901 (N_2901,N_2231,N_1897);
nand U2902 (N_2902,N_1835,N_2007);
nor U2903 (N_2903,N_1806,N_2391);
nand U2904 (N_2904,N_2348,N_2297);
and U2905 (N_2905,N_2022,N_2194);
nor U2906 (N_2906,N_1976,N_1841);
nand U2907 (N_2907,N_2175,N_2277);
nand U2908 (N_2908,N_1921,N_2115);
nand U2909 (N_2909,N_2114,N_1822);
and U2910 (N_2910,N_1947,N_2165);
or U2911 (N_2911,N_2045,N_2205);
and U2912 (N_2912,N_1916,N_1812);
and U2913 (N_2913,N_1867,N_2143);
nand U2914 (N_2914,N_1845,N_2002);
nand U2915 (N_2915,N_1860,N_1948);
nor U2916 (N_2916,N_1987,N_1899);
nor U2917 (N_2917,N_2081,N_1836);
nand U2918 (N_2918,N_2142,N_2351);
and U2919 (N_2919,N_2242,N_1806);
nor U2920 (N_2920,N_2290,N_1801);
nand U2921 (N_2921,N_2152,N_2077);
or U2922 (N_2922,N_2231,N_2180);
nor U2923 (N_2923,N_1830,N_1966);
nor U2924 (N_2924,N_2265,N_2161);
and U2925 (N_2925,N_2126,N_2181);
nor U2926 (N_2926,N_1873,N_2120);
or U2927 (N_2927,N_2237,N_2140);
or U2928 (N_2928,N_1907,N_2364);
nand U2929 (N_2929,N_1953,N_2170);
and U2930 (N_2930,N_2376,N_2385);
nor U2931 (N_2931,N_2123,N_2322);
or U2932 (N_2932,N_2247,N_2091);
nor U2933 (N_2933,N_2373,N_1930);
and U2934 (N_2934,N_1856,N_1859);
or U2935 (N_2935,N_2061,N_1999);
nand U2936 (N_2936,N_2122,N_2108);
nand U2937 (N_2937,N_2315,N_2372);
and U2938 (N_2938,N_2382,N_1814);
nand U2939 (N_2939,N_2308,N_2090);
and U2940 (N_2940,N_2022,N_2174);
nand U2941 (N_2941,N_2394,N_2000);
nor U2942 (N_2942,N_2125,N_1951);
and U2943 (N_2943,N_2133,N_2340);
nor U2944 (N_2944,N_2002,N_2367);
nand U2945 (N_2945,N_2038,N_2137);
or U2946 (N_2946,N_1986,N_1912);
nor U2947 (N_2947,N_1941,N_2165);
nand U2948 (N_2948,N_2306,N_2344);
and U2949 (N_2949,N_1965,N_2000);
nor U2950 (N_2950,N_1992,N_2135);
nand U2951 (N_2951,N_2113,N_1845);
nand U2952 (N_2952,N_2135,N_1976);
or U2953 (N_2953,N_2154,N_2132);
or U2954 (N_2954,N_1827,N_2390);
or U2955 (N_2955,N_2285,N_2102);
nand U2956 (N_2956,N_2052,N_2084);
and U2957 (N_2957,N_2210,N_2184);
nor U2958 (N_2958,N_2074,N_2326);
nor U2959 (N_2959,N_2354,N_1827);
and U2960 (N_2960,N_2283,N_2036);
and U2961 (N_2961,N_2044,N_2336);
or U2962 (N_2962,N_2266,N_1905);
nand U2963 (N_2963,N_1938,N_2367);
or U2964 (N_2964,N_2305,N_2369);
nor U2965 (N_2965,N_2272,N_1810);
nand U2966 (N_2966,N_2065,N_2324);
nor U2967 (N_2967,N_2384,N_2026);
nor U2968 (N_2968,N_2062,N_1951);
nor U2969 (N_2969,N_2270,N_2173);
nand U2970 (N_2970,N_2250,N_1937);
or U2971 (N_2971,N_2274,N_1938);
and U2972 (N_2972,N_2262,N_2088);
and U2973 (N_2973,N_1877,N_1908);
and U2974 (N_2974,N_2206,N_2340);
nand U2975 (N_2975,N_2391,N_2323);
or U2976 (N_2976,N_2038,N_2035);
and U2977 (N_2977,N_2187,N_2163);
or U2978 (N_2978,N_2294,N_2318);
nor U2979 (N_2979,N_1984,N_1852);
and U2980 (N_2980,N_1956,N_1984);
nand U2981 (N_2981,N_2106,N_2072);
and U2982 (N_2982,N_2155,N_2277);
nor U2983 (N_2983,N_1810,N_2315);
nand U2984 (N_2984,N_1800,N_2028);
nor U2985 (N_2985,N_2260,N_2010);
xor U2986 (N_2986,N_1833,N_2208);
and U2987 (N_2987,N_2031,N_2128);
nor U2988 (N_2988,N_1870,N_1815);
nand U2989 (N_2989,N_2148,N_2009);
nor U2990 (N_2990,N_1863,N_2379);
and U2991 (N_2991,N_1809,N_2189);
or U2992 (N_2992,N_2051,N_1955);
or U2993 (N_2993,N_1860,N_2301);
nand U2994 (N_2994,N_1977,N_1884);
and U2995 (N_2995,N_2356,N_2123);
nand U2996 (N_2996,N_1950,N_2213);
nor U2997 (N_2997,N_2091,N_2209);
or U2998 (N_2998,N_1921,N_2339);
and U2999 (N_2999,N_1806,N_2009);
nor UO_0 (O_0,N_2850,N_2993);
and UO_1 (O_1,N_2747,N_2615);
nand UO_2 (O_2,N_2537,N_2544);
nor UO_3 (O_3,N_2614,N_2547);
nor UO_4 (O_4,N_2569,N_2916);
and UO_5 (O_5,N_2434,N_2409);
or UO_6 (O_6,N_2908,N_2542);
or UO_7 (O_7,N_2701,N_2568);
or UO_8 (O_8,N_2667,N_2821);
or UO_9 (O_9,N_2834,N_2731);
nand UO_10 (O_10,N_2951,N_2982);
nor UO_11 (O_11,N_2684,N_2805);
and UO_12 (O_12,N_2425,N_2647);
nor UO_13 (O_13,N_2437,N_2489);
and UO_14 (O_14,N_2661,N_2632);
nand UO_15 (O_15,N_2702,N_2515);
nand UO_16 (O_16,N_2683,N_2750);
nand UO_17 (O_17,N_2773,N_2932);
or UO_18 (O_18,N_2506,N_2595);
and UO_19 (O_19,N_2630,N_2872);
nor UO_20 (O_20,N_2571,N_2934);
or UO_21 (O_21,N_2891,N_2740);
and UO_22 (O_22,N_2937,N_2407);
xor UO_23 (O_23,N_2966,N_2554);
nor UO_24 (O_24,N_2578,N_2924);
xor UO_25 (O_25,N_2759,N_2948);
or UO_26 (O_26,N_2593,N_2718);
nor UO_27 (O_27,N_2655,N_2816);
or UO_28 (O_28,N_2751,N_2873);
and UO_29 (O_29,N_2958,N_2915);
or UO_30 (O_30,N_2929,N_2758);
and UO_31 (O_31,N_2968,N_2820);
nand UO_32 (O_32,N_2481,N_2914);
or UO_33 (O_33,N_2854,N_2460);
nand UO_34 (O_34,N_2613,N_2516);
nor UO_35 (O_35,N_2763,N_2556);
or UO_36 (O_36,N_2996,N_2550);
and UO_37 (O_37,N_2653,N_2811);
nor UO_38 (O_38,N_2662,N_2863);
nand UO_39 (O_39,N_2959,N_2668);
nand UO_40 (O_40,N_2652,N_2415);
nand UO_41 (O_41,N_2988,N_2681);
and UO_42 (O_42,N_2831,N_2642);
or UO_43 (O_43,N_2723,N_2912);
nand UO_44 (O_44,N_2727,N_2498);
and UO_45 (O_45,N_2800,N_2899);
nor UO_46 (O_46,N_2448,N_2401);
nor UO_47 (O_47,N_2840,N_2509);
nand UO_48 (O_48,N_2422,N_2756);
nor UO_49 (O_49,N_2440,N_2430);
or UO_50 (O_50,N_2644,N_2960);
and UO_51 (O_51,N_2771,N_2815);
nor UO_52 (O_52,N_2480,N_2669);
nor UO_53 (O_53,N_2402,N_2772);
nor UO_54 (O_54,N_2824,N_2535);
and UO_55 (O_55,N_2781,N_2742);
nor UO_56 (O_56,N_2582,N_2566);
nor UO_57 (O_57,N_2736,N_2991);
nor UO_58 (O_58,N_2546,N_2706);
or UO_59 (O_59,N_2943,N_2628);
nand UO_60 (O_60,N_2689,N_2973);
nand UO_61 (O_61,N_2843,N_2787);
nand UO_62 (O_62,N_2984,N_2601);
and UO_63 (O_63,N_2594,N_2656);
nor UO_64 (O_64,N_2888,N_2471);
and UO_65 (O_65,N_2746,N_2637);
nand UO_66 (O_66,N_2472,N_2453);
nand UO_67 (O_67,N_2622,N_2627);
or UO_68 (O_68,N_2496,N_2592);
nand UO_69 (O_69,N_2676,N_2999);
nor UO_70 (O_70,N_2953,N_2579);
and UO_71 (O_71,N_2466,N_2427);
nand UO_72 (O_72,N_2512,N_2528);
or UO_73 (O_73,N_2874,N_2618);
or UO_74 (O_74,N_2995,N_2455);
nor UO_75 (O_75,N_2737,N_2513);
nor UO_76 (O_76,N_2970,N_2555);
nand UO_77 (O_77,N_2725,N_2467);
nor UO_78 (O_78,N_2621,N_2974);
nor UO_79 (O_79,N_2478,N_2581);
or UO_80 (O_80,N_2904,N_2584);
or UO_81 (O_81,N_2715,N_2711);
nand UO_82 (O_82,N_2954,N_2986);
and UO_83 (O_83,N_2531,N_2575);
or UO_84 (O_84,N_2545,N_2882);
nand UO_85 (O_85,N_2774,N_2673);
or UO_86 (O_86,N_2896,N_2983);
or UO_87 (O_87,N_2926,N_2499);
nand UO_88 (O_88,N_2977,N_2590);
or UO_89 (O_89,N_2950,N_2775);
or UO_90 (O_90,N_2892,N_2827);
or UO_91 (O_91,N_2610,N_2410);
nand UO_92 (O_92,N_2698,N_2998);
xnor UO_93 (O_93,N_2803,N_2769);
nor UO_94 (O_94,N_2732,N_2832);
nand UO_95 (O_95,N_2798,N_2743);
nand UO_96 (O_96,N_2606,N_2797);
nor UO_97 (O_97,N_2431,N_2757);
xor UO_98 (O_98,N_2646,N_2826);
or UO_99 (O_99,N_2664,N_2928);
or UO_100 (O_100,N_2487,N_2938);
nand UO_101 (O_101,N_2461,N_2458);
nor UO_102 (O_102,N_2690,N_2946);
or UO_103 (O_103,N_2792,N_2403);
and UO_104 (O_104,N_2865,N_2491);
or UO_105 (O_105,N_2710,N_2965);
or UO_106 (O_106,N_2573,N_2439);
nor UO_107 (O_107,N_2436,N_2881);
nor UO_108 (O_108,N_2859,N_2791);
nand UO_109 (O_109,N_2726,N_2910);
or UO_110 (O_110,N_2700,N_2432);
nand UO_111 (O_111,N_2452,N_2957);
and UO_112 (O_112,N_2780,N_2864);
nor UO_113 (O_113,N_2435,N_2519);
or UO_114 (O_114,N_2438,N_2482);
nor UO_115 (O_115,N_2521,N_2955);
nor UO_116 (O_116,N_2650,N_2465);
nor UO_117 (O_117,N_2479,N_2709);
or UO_118 (O_118,N_2877,N_2895);
and UO_119 (O_119,N_2503,N_2890);
or UO_120 (O_120,N_2539,N_2851);
nor UO_121 (O_121,N_2704,N_2806);
nor UO_122 (O_122,N_2623,N_2421);
nand UO_123 (O_123,N_2878,N_2540);
or UO_124 (O_124,N_2645,N_2901);
nor UO_125 (O_125,N_2449,N_2962);
nand UO_126 (O_126,N_2883,N_2484);
and UO_127 (O_127,N_2429,N_2490);
nor UO_128 (O_128,N_2524,N_2795);
nand UO_129 (O_129,N_2587,N_2909);
nor UO_130 (O_130,N_2752,N_2492);
nor UO_131 (O_131,N_2641,N_2994);
xnor UO_132 (O_132,N_2541,N_2852);
nand UO_133 (O_133,N_2720,N_2534);
nand UO_134 (O_134,N_2526,N_2708);
and UO_135 (O_135,N_2624,N_2860);
nor UO_136 (O_136,N_2703,N_2822);
or UO_137 (O_137,N_2707,N_2724);
and UO_138 (O_138,N_2404,N_2413);
nor UO_139 (O_139,N_2405,N_2975);
and UO_140 (O_140,N_2939,N_2788);
nand UO_141 (O_141,N_2952,N_2651);
xor UO_142 (O_142,N_2588,N_2730);
or UO_143 (O_143,N_2699,N_2412);
or UO_144 (O_144,N_2445,N_2533);
xor UO_145 (O_145,N_2680,N_2721);
and UO_146 (O_146,N_2940,N_2643);
nor UO_147 (O_147,N_2985,N_2903);
nor UO_148 (O_148,N_2557,N_2906);
nor UO_149 (O_149,N_2713,N_2599);
or UO_150 (O_150,N_2814,N_2518);
nand UO_151 (O_151,N_2495,N_2483);
nor UO_152 (O_152,N_2514,N_2799);
and UO_153 (O_153,N_2585,N_2944);
nor UO_154 (O_154,N_2898,N_2424);
or UO_155 (O_155,N_2817,N_2551);
nand UO_156 (O_156,N_2474,N_2619);
nor UO_157 (O_157,N_2931,N_2511);
nand UO_158 (O_158,N_2473,N_2635);
nand UO_159 (O_159,N_2530,N_2416);
nor UO_160 (O_160,N_2604,N_2576);
nand UO_161 (O_161,N_2971,N_2945);
or UO_162 (O_162,N_2470,N_2728);
nand UO_163 (O_163,N_2485,N_2688);
nand UO_164 (O_164,N_2505,N_2801);
nor UO_165 (O_165,N_2745,N_2666);
xor UO_166 (O_166,N_2504,N_2616);
or UO_167 (O_167,N_2612,N_2687);
nand UO_168 (O_168,N_2829,N_2523);
nor UO_169 (O_169,N_2411,N_2987);
or UO_170 (O_170,N_2672,N_2574);
and UO_171 (O_171,N_2639,N_2900);
or UO_172 (O_172,N_2770,N_2777);
nor UO_173 (O_173,N_2990,N_2572);
or UO_174 (O_174,N_2633,N_2497);
and UO_175 (O_175,N_2762,N_2560);
nand UO_176 (O_176,N_2935,N_2580);
and UO_177 (O_177,N_2459,N_2749);
and UO_178 (O_178,N_2714,N_2640);
and UO_179 (O_179,N_2845,N_2552);
nor UO_180 (O_180,N_2626,N_2857);
nand UO_181 (O_181,N_2789,N_2813);
nor UO_182 (O_182,N_2598,N_2441);
nand UO_183 (O_183,N_2921,N_2867);
or UO_184 (O_184,N_2920,N_2997);
and UO_185 (O_185,N_2469,N_2500);
nor UO_186 (O_186,N_2502,N_2716);
nand UO_187 (O_187,N_2693,N_2833);
nand UO_188 (O_188,N_2565,N_2722);
or UO_189 (O_189,N_2685,N_2744);
nand UO_190 (O_190,N_2433,N_2597);
nor UO_191 (O_191,N_2767,N_2885);
or UO_192 (O_192,N_2733,N_2527);
or UO_193 (O_193,N_2897,N_2942);
or UO_194 (O_194,N_2591,N_2947);
or UO_195 (O_195,N_2949,N_2790);
and UO_196 (O_196,N_2956,N_2869);
nor UO_197 (O_197,N_2918,N_2674);
or UO_198 (O_198,N_2712,N_2605);
or UO_199 (O_199,N_2548,N_2665);
and UO_200 (O_200,N_2629,N_2907);
and UO_201 (O_201,N_2917,N_2760);
nand UO_202 (O_202,N_2783,N_2420);
nand UO_203 (O_203,N_2784,N_2636);
nand UO_204 (O_204,N_2812,N_2922);
or UO_205 (O_205,N_2893,N_2563);
or UO_206 (O_206,N_2486,N_2675);
or UO_207 (O_207,N_2695,N_2753);
xor UO_208 (O_208,N_2611,N_2989);
or UO_209 (O_209,N_2444,N_2782);
or UO_210 (O_210,N_2553,N_2902);
or UO_211 (O_211,N_2558,N_2451);
nand UO_212 (O_212,N_2735,N_2858);
or UO_213 (O_213,N_2884,N_2961);
nor UO_214 (O_214,N_2638,N_2741);
nand UO_215 (O_215,N_2804,N_2980);
nand UO_216 (O_216,N_2905,N_2941);
nor UO_217 (O_217,N_2561,N_2889);
nor UO_218 (O_218,N_2870,N_2734);
or UO_219 (O_219,N_2810,N_2450);
nand UO_220 (O_220,N_2964,N_2856);
nand UO_221 (O_221,N_2835,N_2596);
and UO_222 (O_222,N_2525,N_2875);
nand UO_223 (O_223,N_2475,N_2844);
and UO_224 (O_224,N_2522,N_2508);
nand UO_225 (O_225,N_2507,N_2793);
or UO_226 (O_226,N_2755,N_2838);
and UO_227 (O_227,N_2494,N_2538);
or UO_228 (O_228,N_2764,N_2930);
nand UO_229 (O_229,N_2631,N_2696);
xor UO_230 (O_230,N_2738,N_2808);
and UO_231 (O_231,N_2697,N_2677);
nand UO_232 (O_232,N_2818,N_2686);
and UO_233 (O_233,N_2670,N_2691);
nor UO_234 (O_234,N_2570,N_2510);
or UO_235 (O_235,N_2879,N_2981);
nand UO_236 (O_236,N_2823,N_2678);
nand UO_237 (O_237,N_2849,N_2443);
nand UO_238 (O_238,N_2919,N_2933);
or UO_239 (O_239,N_2426,N_2887);
or UO_240 (O_240,N_2682,N_2786);
or UO_241 (O_241,N_2748,N_2419);
nor UO_242 (O_242,N_2754,N_2847);
or UO_243 (O_243,N_2841,N_2936);
or UO_244 (O_244,N_2853,N_2719);
and UO_245 (O_245,N_2520,N_2659);
and UO_246 (O_246,N_2848,N_2408);
or UO_247 (O_247,N_2583,N_2447);
nand UO_248 (O_248,N_2794,N_2717);
nand UO_249 (O_249,N_2969,N_2785);
and UO_250 (O_250,N_2559,N_2649);
and UO_251 (O_251,N_2603,N_2414);
or UO_252 (O_252,N_2428,N_2493);
or UO_253 (O_253,N_2457,N_2658);
nor UO_254 (O_254,N_2830,N_2979);
or UO_255 (O_255,N_2925,N_2468);
or UO_256 (O_256,N_2729,N_2976);
and UO_257 (O_257,N_2880,N_2654);
and UO_258 (O_258,N_2517,N_2765);
and UO_259 (O_259,N_2671,N_2417);
nand UO_260 (O_260,N_2807,N_2705);
nor UO_261 (O_261,N_2819,N_2549);
or UO_262 (O_262,N_2739,N_2602);
and UO_263 (O_263,N_2607,N_2400);
nand UO_264 (O_264,N_2634,N_2842);
or UO_265 (O_265,N_2657,N_2761);
or UO_266 (O_266,N_2600,N_2927);
nor UO_267 (O_267,N_2543,N_2779);
and UO_268 (O_268,N_2679,N_2442);
and UO_269 (O_269,N_2476,N_2406);
or UO_270 (O_270,N_2839,N_2648);
nand UO_271 (O_271,N_2894,N_2456);
nand UO_272 (O_272,N_2886,N_2868);
nand UO_273 (O_273,N_2463,N_2855);
and UO_274 (O_274,N_2992,N_2768);
and UO_275 (O_275,N_2871,N_2846);
and UO_276 (O_276,N_2418,N_2564);
nor UO_277 (O_277,N_2911,N_2862);
nand UO_278 (O_278,N_2609,N_2577);
nor UO_279 (O_279,N_2586,N_2825);
or UO_280 (O_280,N_2423,N_2608);
nand UO_281 (O_281,N_2625,N_2828);
nor UO_282 (O_282,N_2776,N_2978);
xor UO_283 (O_283,N_2796,N_2837);
nor UO_284 (O_284,N_2562,N_2967);
and UO_285 (O_285,N_2766,N_2532);
and UO_286 (O_286,N_2617,N_2620);
nand UO_287 (O_287,N_2536,N_2972);
nand UO_288 (O_288,N_2836,N_2660);
or UO_289 (O_289,N_2464,N_2809);
nor UO_290 (O_290,N_2963,N_2446);
or UO_291 (O_291,N_2802,N_2589);
and UO_292 (O_292,N_2876,N_2454);
nor UO_293 (O_293,N_2692,N_2866);
nand UO_294 (O_294,N_2663,N_2501);
nand UO_295 (O_295,N_2694,N_2462);
xnor UO_296 (O_296,N_2861,N_2923);
nand UO_297 (O_297,N_2913,N_2778);
nand UO_298 (O_298,N_2477,N_2488);
and UO_299 (O_299,N_2529,N_2567);
or UO_300 (O_300,N_2801,N_2459);
xor UO_301 (O_301,N_2917,N_2736);
or UO_302 (O_302,N_2649,N_2921);
nor UO_303 (O_303,N_2709,N_2894);
and UO_304 (O_304,N_2400,N_2677);
nor UO_305 (O_305,N_2959,N_2652);
and UO_306 (O_306,N_2878,N_2643);
and UO_307 (O_307,N_2792,N_2710);
and UO_308 (O_308,N_2703,N_2839);
or UO_309 (O_309,N_2701,N_2828);
or UO_310 (O_310,N_2487,N_2971);
or UO_311 (O_311,N_2627,N_2575);
nor UO_312 (O_312,N_2455,N_2911);
nor UO_313 (O_313,N_2983,N_2585);
nor UO_314 (O_314,N_2828,N_2988);
nor UO_315 (O_315,N_2733,N_2784);
and UO_316 (O_316,N_2406,N_2402);
nand UO_317 (O_317,N_2899,N_2607);
or UO_318 (O_318,N_2853,N_2666);
nor UO_319 (O_319,N_2725,N_2850);
and UO_320 (O_320,N_2675,N_2992);
nand UO_321 (O_321,N_2883,N_2881);
or UO_322 (O_322,N_2924,N_2875);
nand UO_323 (O_323,N_2691,N_2789);
nand UO_324 (O_324,N_2460,N_2839);
nand UO_325 (O_325,N_2595,N_2974);
and UO_326 (O_326,N_2701,N_2891);
nand UO_327 (O_327,N_2637,N_2842);
and UO_328 (O_328,N_2836,N_2544);
and UO_329 (O_329,N_2876,N_2498);
nor UO_330 (O_330,N_2450,N_2479);
nand UO_331 (O_331,N_2463,N_2779);
and UO_332 (O_332,N_2482,N_2989);
nor UO_333 (O_333,N_2612,N_2409);
nand UO_334 (O_334,N_2569,N_2811);
nand UO_335 (O_335,N_2618,N_2520);
and UO_336 (O_336,N_2551,N_2425);
nor UO_337 (O_337,N_2571,N_2488);
and UO_338 (O_338,N_2718,N_2707);
and UO_339 (O_339,N_2801,N_2660);
nor UO_340 (O_340,N_2655,N_2871);
or UO_341 (O_341,N_2938,N_2959);
nor UO_342 (O_342,N_2942,N_2917);
nor UO_343 (O_343,N_2779,N_2600);
or UO_344 (O_344,N_2490,N_2770);
nor UO_345 (O_345,N_2852,N_2870);
or UO_346 (O_346,N_2684,N_2678);
nand UO_347 (O_347,N_2800,N_2781);
and UO_348 (O_348,N_2895,N_2794);
nor UO_349 (O_349,N_2416,N_2879);
nor UO_350 (O_350,N_2503,N_2866);
nor UO_351 (O_351,N_2425,N_2803);
or UO_352 (O_352,N_2570,N_2624);
nor UO_353 (O_353,N_2886,N_2592);
and UO_354 (O_354,N_2627,N_2894);
or UO_355 (O_355,N_2642,N_2455);
or UO_356 (O_356,N_2979,N_2965);
nor UO_357 (O_357,N_2762,N_2813);
or UO_358 (O_358,N_2985,N_2521);
nand UO_359 (O_359,N_2515,N_2991);
nand UO_360 (O_360,N_2629,N_2981);
and UO_361 (O_361,N_2447,N_2994);
or UO_362 (O_362,N_2789,N_2595);
nand UO_363 (O_363,N_2906,N_2800);
nor UO_364 (O_364,N_2776,N_2436);
nor UO_365 (O_365,N_2676,N_2852);
and UO_366 (O_366,N_2560,N_2686);
and UO_367 (O_367,N_2848,N_2532);
nand UO_368 (O_368,N_2449,N_2658);
nand UO_369 (O_369,N_2931,N_2485);
xor UO_370 (O_370,N_2477,N_2687);
xnor UO_371 (O_371,N_2624,N_2641);
nor UO_372 (O_372,N_2835,N_2681);
nand UO_373 (O_373,N_2969,N_2549);
nand UO_374 (O_374,N_2444,N_2916);
nand UO_375 (O_375,N_2665,N_2893);
or UO_376 (O_376,N_2878,N_2464);
nor UO_377 (O_377,N_2459,N_2648);
nand UO_378 (O_378,N_2654,N_2818);
nand UO_379 (O_379,N_2556,N_2543);
nand UO_380 (O_380,N_2769,N_2535);
nand UO_381 (O_381,N_2810,N_2664);
or UO_382 (O_382,N_2629,N_2858);
and UO_383 (O_383,N_2661,N_2930);
nor UO_384 (O_384,N_2705,N_2841);
nand UO_385 (O_385,N_2489,N_2793);
nand UO_386 (O_386,N_2804,N_2592);
nand UO_387 (O_387,N_2632,N_2715);
nor UO_388 (O_388,N_2771,N_2481);
nor UO_389 (O_389,N_2508,N_2477);
and UO_390 (O_390,N_2665,N_2573);
nor UO_391 (O_391,N_2512,N_2831);
or UO_392 (O_392,N_2844,N_2899);
or UO_393 (O_393,N_2858,N_2882);
nand UO_394 (O_394,N_2537,N_2457);
and UO_395 (O_395,N_2427,N_2744);
or UO_396 (O_396,N_2571,N_2914);
and UO_397 (O_397,N_2829,N_2962);
or UO_398 (O_398,N_2682,N_2686);
nand UO_399 (O_399,N_2968,N_2594);
xnor UO_400 (O_400,N_2826,N_2573);
or UO_401 (O_401,N_2848,N_2830);
and UO_402 (O_402,N_2582,N_2926);
and UO_403 (O_403,N_2947,N_2611);
nand UO_404 (O_404,N_2713,N_2566);
or UO_405 (O_405,N_2933,N_2938);
nor UO_406 (O_406,N_2656,N_2514);
nand UO_407 (O_407,N_2497,N_2663);
and UO_408 (O_408,N_2456,N_2758);
and UO_409 (O_409,N_2823,N_2807);
xor UO_410 (O_410,N_2780,N_2443);
and UO_411 (O_411,N_2670,N_2528);
or UO_412 (O_412,N_2751,N_2742);
and UO_413 (O_413,N_2945,N_2434);
nor UO_414 (O_414,N_2813,N_2603);
and UO_415 (O_415,N_2729,N_2983);
nand UO_416 (O_416,N_2964,N_2902);
and UO_417 (O_417,N_2686,N_2400);
nor UO_418 (O_418,N_2499,N_2993);
nand UO_419 (O_419,N_2899,N_2493);
xor UO_420 (O_420,N_2522,N_2675);
and UO_421 (O_421,N_2805,N_2936);
or UO_422 (O_422,N_2490,N_2873);
or UO_423 (O_423,N_2407,N_2575);
nor UO_424 (O_424,N_2522,N_2949);
and UO_425 (O_425,N_2450,N_2715);
and UO_426 (O_426,N_2940,N_2519);
and UO_427 (O_427,N_2929,N_2427);
nand UO_428 (O_428,N_2590,N_2774);
or UO_429 (O_429,N_2439,N_2719);
or UO_430 (O_430,N_2437,N_2787);
xnor UO_431 (O_431,N_2639,N_2440);
or UO_432 (O_432,N_2515,N_2707);
nand UO_433 (O_433,N_2418,N_2850);
or UO_434 (O_434,N_2953,N_2499);
xnor UO_435 (O_435,N_2949,N_2612);
and UO_436 (O_436,N_2902,N_2481);
and UO_437 (O_437,N_2944,N_2407);
and UO_438 (O_438,N_2643,N_2586);
and UO_439 (O_439,N_2621,N_2922);
or UO_440 (O_440,N_2587,N_2654);
or UO_441 (O_441,N_2604,N_2818);
nand UO_442 (O_442,N_2567,N_2412);
xnor UO_443 (O_443,N_2852,N_2899);
and UO_444 (O_444,N_2709,N_2469);
and UO_445 (O_445,N_2813,N_2824);
nand UO_446 (O_446,N_2741,N_2950);
and UO_447 (O_447,N_2931,N_2827);
nor UO_448 (O_448,N_2485,N_2590);
or UO_449 (O_449,N_2827,N_2403);
and UO_450 (O_450,N_2553,N_2493);
or UO_451 (O_451,N_2804,N_2896);
and UO_452 (O_452,N_2924,N_2831);
nand UO_453 (O_453,N_2882,N_2861);
nand UO_454 (O_454,N_2668,N_2917);
and UO_455 (O_455,N_2701,N_2560);
xnor UO_456 (O_456,N_2593,N_2830);
or UO_457 (O_457,N_2548,N_2656);
and UO_458 (O_458,N_2822,N_2971);
and UO_459 (O_459,N_2528,N_2763);
nor UO_460 (O_460,N_2549,N_2731);
and UO_461 (O_461,N_2785,N_2939);
and UO_462 (O_462,N_2844,N_2596);
and UO_463 (O_463,N_2452,N_2597);
nand UO_464 (O_464,N_2789,N_2784);
nor UO_465 (O_465,N_2945,N_2548);
nor UO_466 (O_466,N_2811,N_2433);
or UO_467 (O_467,N_2419,N_2704);
and UO_468 (O_468,N_2782,N_2522);
nor UO_469 (O_469,N_2446,N_2412);
nor UO_470 (O_470,N_2612,N_2822);
nand UO_471 (O_471,N_2627,N_2493);
or UO_472 (O_472,N_2633,N_2945);
nand UO_473 (O_473,N_2991,N_2583);
and UO_474 (O_474,N_2760,N_2515);
nand UO_475 (O_475,N_2503,N_2887);
nand UO_476 (O_476,N_2586,N_2991);
and UO_477 (O_477,N_2585,N_2524);
and UO_478 (O_478,N_2637,N_2821);
and UO_479 (O_479,N_2427,N_2776);
nand UO_480 (O_480,N_2501,N_2824);
nor UO_481 (O_481,N_2983,N_2908);
nor UO_482 (O_482,N_2929,N_2523);
nor UO_483 (O_483,N_2407,N_2544);
and UO_484 (O_484,N_2717,N_2951);
or UO_485 (O_485,N_2601,N_2605);
or UO_486 (O_486,N_2447,N_2921);
nand UO_487 (O_487,N_2978,N_2440);
nor UO_488 (O_488,N_2891,N_2797);
and UO_489 (O_489,N_2735,N_2601);
or UO_490 (O_490,N_2800,N_2950);
nand UO_491 (O_491,N_2910,N_2931);
or UO_492 (O_492,N_2977,N_2772);
nand UO_493 (O_493,N_2461,N_2516);
or UO_494 (O_494,N_2932,N_2649);
and UO_495 (O_495,N_2695,N_2735);
nor UO_496 (O_496,N_2817,N_2954);
nor UO_497 (O_497,N_2462,N_2879);
and UO_498 (O_498,N_2569,N_2744);
xnor UO_499 (O_499,N_2996,N_2430);
endmodule