module basic_3000_30000_3500_20_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
or U0 (N_0,In_1240,In_1556);
and U1 (N_1,In_2597,In_1095);
nand U2 (N_2,In_2717,In_2613);
nor U3 (N_3,In_2590,In_2012);
nor U4 (N_4,In_276,In_1144);
and U5 (N_5,In_1883,In_1600);
xor U6 (N_6,In_2336,In_738);
nor U7 (N_7,In_506,In_2442);
nor U8 (N_8,In_842,In_2310);
or U9 (N_9,In_1957,In_1963);
nand U10 (N_10,In_562,In_986);
nor U11 (N_11,In_269,In_601);
nand U12 (N_12,In_2115,In_2788);
nor U13 (N_13,In_733,In_2672);
or U14 (N_14,In_649,In_1879);
nor U15 (N_15,In_2298,In_2969);
nor U16 (N_16,In_2749,In_1921);
xor U17 (N_17,In_716,In_1329);
nand U18 (N_18,In_284,In_1553);
xor U19 (N_19,In_850,In_2588);
and U20 (N_20,In_686,In_548);
nor U21 (N_21,In_982,In_1827);
nand U22 (N_22,In_1544,In_1984);
nand U23 (N_23,In_2091,In_2865);
nand U24 (N_24,In_1014,In_366);
and U25 (N_25,In_820,In_2350);
nand U26 (N_26,In_371,In_2827);
xnor U27 (N_27,In_66,In_1300);
nand U28 (N_28,In_1130,In_1295);
or U29 (N_29,In_2695,In_1842);
and U30 (N_30,In_1245,In_1395);
nand U31 (N_31,In_1381,In_248);
or U32 (N_32,In_1188,In_2516);
and U33 (N_33,In_1998,In_2947);
and U34 (N_34,In_1980,In_454);
nor U35 (N_35,In_2327,In_714);
nand U36 (N_36,In_2252,In_2525);
xnor U37 (N_37,In_2108,In_2368);
xnor U38 (N_38,In_2820,In_2742);
nor U39 (N_39,In_258,In_2348);
or U40 (N_40,In_134,In_2266);
nor U41 (N_41,In_1226,In_459);
xor U42 (N_42,In_1453,In_663);
nor U43 (N_43,In_473,In_2438);
or U44 (N_44,In_1511,In_1754);
xor U45 (N_45,In_2834,In_313);
nand U46 (N_46,In_1074,In_202);
nand U47 (N_47,In_1434,In_1782);
or U48 (N_48,In_1663,In_2522);
xnor U49 (N_49,In_179,In_634);
or U50 (N_50,In_2066,In_2104);
xnor U51 (N_51,In_1697,In_2250);
or U52 (N_52,In_104,In_2398);
nand U53 (N_53,In_1,In_130);
xor U54 (N_54,In_2406,In_1474);
nor U55 (N_55,In_144,In_1997);
nand U56 (N_56,In_1472,In_2445);
and U57 (N_57,In_885,In_1923);
nand U58 (N_58,In_1652,In_1868);
nor U59 (N_59,In_2378,In_2906);
or U60 (N_60,In_2913,In_679);
and U61 (N_61,In_346,In_871);
nand U62 (N_62,In_2692,In_542);
and U63 (N_63,In_1196,In_1840);
nand U64 (N_64,In_2410,In_1151);
and U65 (N_65,In_2386,In_2514);
nand U66 (N_66,In_1205,In_2685);
xnor U67 (N_67,In_1785,In_496);
nand U68 (N_68,In_1593,In_2646);
xor U69 (N_69,In_770,In_813);
xor U70 (N_70,In_1862,In_230);
xnor U71 (N_71,In_2923,In_183);
or U72 (N_72,In_1618,In_420);
nand U73 (N_73,In_537,In_2200);
xor U74 (N_74,In_290,In_1486);
nor U75 (N_75,In_1097,In_817);
nand U76 (N_76,In_941,In_2289);
nand U77 (N_77,In_2859,In_190);
xor U78 (N_78,In_1508,In_37);
or U79 (N_79,In_1276,In_1292);
nand U80 (N_80,In_538,In_2976);
or U81 (N_81,In_1443,In_1136);
xnor U82 (N_82,In_1212,In_1811);
and U83 (N_83,In_324,In_254);
or U84 (N_84,In_660,In_818);
nand U85 (N_85,In_809,In_1162);
and U86 (N_86,In_1447,In_1433);
nand U87 (N_87,In_2498,In_2482);
or U88 (N_88,In_484,In_2701);
nor U89 (N_89,In_2309,In_825);
and U90 (N_90,In_1849,In_1799);
xnor U91 (N_91,In_1523,In_341);
or U92 (N_92,In_235,In_376);
nor U93 (N_93,In_287,In_2562);
and U94 (N_94,In_2286,In_607);
or U95 (N_95,In_1002,In_596);
nand U96 (N_96,In_2433,In_852);
xnor U97 (N_97,In_1731,In_2822);
or U98 (N_98,In_2428,In_1279);
nand U99 (N_99,In_608,In_2813);
nand U100 (N_100,In_1435,In_2193);
nor U101 (N_101,In_1890,In_2006);
or U102 (N_102,In_1770,In_830);
and U103 (N_103,In_766,In_1837);
xnor U104 (N_104,In_905,In_4);
xnor U105 (N_105,In_2372,In_408);
nor U106 (N_106,In_2735,In_1104);
and U107 (N_107,In_1255,In_752);
xor U108 (N_108,In_2771,In_298);
xnor U109 (N_109,In_2149,In_1515);
and U110 (N_110,In_2322,In_2211);
and U111 (N_111,In_792,In_41);
nand U112 (N_112,In_288,In_2558);
and U113 (N_113,In_1666,In_1516);
nor U114 (N_114,In_461,In_502);
nand U115 (N_115,In_1535,In_2342);
nand U116 (N_116,In_526,In_1214);
or U117 (N_117,In_563,In_81);
nand U118 (N_118,In_923,In_693);
and U119 (N_119,In_838,In_297);
and U120 (N_120,In_1044,In_2244);
xnor U121 (N_121,In_2574,In_912);
xor U122 (N_122,In_1482,In_1971);
nor U123 (N_123,In_1901,In_406);
or U124 (N_124,In_1117,In_1277);
or U125 (N_125,In_477,In_2708);
xnor U126 (N_126,In_217,In_1354);
or U127 (N_127,In_1720,In_727);
nand U128 (N_128,In_724,In_673);
xnor U129 (N_129,In_200,In_1638);
nor U130 (N_130,In_631,In_2828);
or U131 (N_131,In_1684,In_2534);
nand U132 (N_132,In_334,In_1422);
xnor U133 (N_133,In_2796,In_2608);
nand U134 (N_134,In_1777,In_2996);
nand U135 (N_135,In_2292,In_1530);
and U136 (N_136,In_1886,In_2405);
and U137 (N_137,In_1787,In_2893);
xnor U138 (N_138,In_427,In_1824);
xor U139 (N_139,In_1471,In_469);
and U140 (N_140,In_403,In_2150);
nor U141 (N_141,In_2146,In_2112);
or U142 (N_142,In_633,In_1071);
or U143 (N_143,In_2468,In_1978);
and U144 (N_144,In_2496,In_2724);
or U145 (N_145,In_265,In_2073);
nor U146 (N_146,In_106,In_1333);
and U147 (N_147,In_1863,In_1759);
or U148 (N_148,In_1677,In_2639);
or U149 (N_149,In_1022,In_1539);
nor U150 (N_150,In_699,In_1178);
nand U151 (N_151,In_1410,In_1709);
nor U152 (N_152,In_1907,In_1451);
or U153 (N_153,In_2759,In_191);
nand U154 (N_154,In_1307,In_638);
nand U155 (N_155,In_1650,In_1909);
or U156 (N_156,In_533,In_89);
and U157 (N_157,In_1919,In_101);
nor U158 (N_158,In_811,In_1249);
nor U159 (N_159,In_2663,In_2751);
or U160 (N_160,In_2024,In_1867);
xor U161 (N_161,In_1937,In_2321);
xor U162 (N_162,In_2811,In_2352);
xnor U163 (N_163,In_128,In_2985);
xor U164 (N_164,In_2917,In_1804);
xnor U165 (N_165,In_1475,In_40);
or U166 (N_166,In_1135,In_1165);
nor U167 (N_167,In_2617,In_197);
and U168 (N_168,In_2915,In_2578);
nor U169 (N_169,In_2444,In_1414);
or U170 (N_170,In_886,In_2951);
or U171 (N_171,In_2557,In_1753);
and U172 (N_172,In_650,In_2623);
nand U173 (N_173,In_1749,In_2768);
and U174 (N_174,In_1316,In_675);
and U175 (N_175,In_1653,In_2414);
or U176 (N_176,In_1616,In_107);
xor U177 (N_177,In_2159,In_2866);
and U178 (N_178,In_2703,In_2688);
or U179 (N_179,In_1889,In_2598);
and U180 (N_180,In_1665,In_470);
nor U181 (N_181,In_536,In_2486);
or U182 (N_182,In_1432,In_1953);
nand U183 (N_183,In_2991,In_1066);
or U184 (N_184,In_246,In_2715);
and U185 (N_185,In_389,In_1747);
or U186 (N_186,In_2280,In_2532);
or U187 (N_187,In_2520,In_1239);
xnor U188 (N_188,In_262,In_1941);
and U189 (N_189,In_925,In_2824);
nand U190 (N_190,In_920,In_2876);
or U191 (N_191,In_1762,In_1915);
or U192 (N_192,In_1087,In_2090);
nand U193 (N_193,In_1325,In_1856);
and U194 (N_194,In_893,In_2704);
xnor U195 (N_195,In_29,In_209);
nor U196 (N_196,In_579,In_1826);
nand U197 (N_197,In_2587,In_2081);
nand U198 (N_198,In_917,In_954);
xor U199 (N_199,In_980,In_736);
nand U200 (N_200,In_1365,In_1994);
nor U201 (N_201,In_2973,In_708);
or U202 (N_202,In_2400,In_127);
nand U203 (N_203,In_1498,In_1960);
xnor U204 (N_204,In_1254,In_2860);
and U205 (N_205,In_869,In_315);
and U206 (N_206,In_1012,In_2698);
nor U207 (N_207,In_643,In_2541);
nor U208 (N_208,In_1568,In_2265);
or U209 (N_209,In_2925,In_2014);
or U210 (N_210,In_1814,In_2273);
or U211 (N_211,In_2157,In_2652);
xnor U212 (N_212,In_1949,In_985);
nand U213 (N_213,In_2584,In_602);
xor U214 (N_214,In_1779,In_2807);
or U215 (N_215,In_847,In_816);
xnor U216 (N_216,In_1194,In_1386);
xor U217 (N_217,In_2517,In_1331);
and U218 (N_218,In_2756,In_1200);
nor U219 (N_219,In_944,In_46);
xor U220 (N_220,In_256,In_2183);
and U221 (N_221,In_1263,In_336);
nor U222 (N_222,In_1791,In_1501);
or U223 (N_223,In_1664,In_1076);
nand U224 (N_224,In_1730,In_141);
nor U225 (N_225,In_1063,In_368);
xnor U226 (N_226,In_1131,In_27);
and U227 (N_227,In_1851,In_2540);
or U228 (N_228,In_1911,In_132);
and U229 (N_229,In_2366,In_424);
xnor U230 (N_230,In_822,In_908);
nor U231 (N_231,In_142,In_926);
and U232 (N_232,In_2840,In_1574);
xor U233 (N_233,In_2766,In_467);
or U234 (N_234,In_277,In_2376);
nor U235 (N_235,In_1109,In_2539);
nor U236 (N_236,In_2757,In_946);
nor U237 (N_237,In_1565,In_1428);
or U238 (N_238,In_2382,In_1606);
xnor U239 (N_239,In_2883,In_1213);
and U240 (N_240,In_181,In_1982);
xnor U241 (N_241,In_1764,In_2778);
xor U242 (N_242,In_97,In_1349);
xor U243 (N_243,In_2306,In_2094);
or U244 (N_244,In_2307,In_407);
xor U245 (N_245,In_1794,In_1658);
or U246 (N_246,In_2994,In_1636);
or U247 (N_247,In_1671,In_481);
or U248 (N_248,In_1455,In_2744);
nand U249 (N_249,In_1829,In_2293);
xor U250 (N_250,In_2015,In_1719);
nand U251 (N_251,In_965,In_966);
nor U252 (N_252,In_1098,In_2332);
and U253 (N_253,In_1152,In_300);
or U254 (N_254,In_1721,In_1114);
nor U255 (N_255,In_991,In_2997);
nand U256 (N_256,In_777,In_1489);
xnor U257 (N_257,In_1473,In_513);
xor U258 (N_258,In_2007,In_719);
or U259 (N_259,In_1018,In_165);
xnor U260 (N_260,In_2379,In_411);
xnor U261 (N_261,In_1776,In_689);
and U262 (N_262,In_466,In_1227);
or U263 (N_263,In_2419,In_1286);
nor U264 (N_264,In_2942,In_1154);
nand U265 (N_265,In_2555,In_2360);
and U266 (N_266,In_2396,In_1908);
nand U267 (N_267,In_1797,In_860);
and U268 (N_268,In_554,In_99);
and U269 (N_269,In_1113,In_74);
nor U270 (N_270,In_1020,In_1560);
nor U271 (N_271,In_2363,In_2047);
nor U272 (N_272,In_347,In_2491);
nor U273 (N_273,In_205,In_1297);
nand U274 (N_274,In_2791,In_52);
xor U275 (N_275,In_2592,In_995);
xnor U276 (N_276,In_2357,In_2920);
xnor U277 (N_277,In_2641,In_474);
nand U278 (N_278,In_1000,In_1605);
nand U279 (N_279,In_1241,In_531);
nand U280 (N_280,In_1427,In_31);
and U281 (N_281,In_2831,In_1407);
or U282 (N_282,In_2237,In_1185);
or U283 (N_283,In_176,In_2019);
nor U284 (N_284,In_2518,In_2814);
or U285 (N_285,In_2027,In_1742);
and U286 (N_286,In_159,In_422);
and U287 (N_287,In_806,In_1847);
and U288 (N_288,In_1094,In_1393);
nor U289 (N_289,In_2902,In_59);
xnor U290 (N_290,In_2215,In_942);
nor U291 (N_291,In_2671,In_943);
xnor U292 (N_292,In_2191,In_1882);
nor U293 (N_293,In_529,In_1064);
xor U294 (N_294,In_1929,In_1243);
xor U295 (N_295,In_2473,In_2537);
nor U296 (N_296,In_874,In_2053);
nor U297 (N_297,In_88,In_857);
xnor U298 (N_298,In_1256,In_1966);
nor U299 (N_299,In_453,In_2576);
nand U300 (N_300,In_1976,In_665);
nor U301 (N_301,In_2453,In_630);
nor U302 (N_302,In_1528,In_1841);
nand U303 (N_303,In_432,In_1751);
nor U304 (N_304,In_2201,In_1115);
nand U305 (N_305,In_1877,In_94);
xor U306 (N_306,In_567,In_1046);
xor U307 (N_307,In_2269,In_1502);
or U308 (N_308,In_8,In_624);
xor U309 (N_309,In_1716,In_69);
nor U310 (N_310,In_2088,In_763);
or U311 (N_311,In_2160,In_2817);
or U312 (N_312,In_2643,In_1924);
nand U313 (N_313,In_75,In_1081);
and U314 (N_314,In_2620,In_2448);
or U315 (N_315,In_273,In_2455);
and U316 (N_316,In_2572,In_1027);
nand U317 (N_317,In_1521,In_1536);
and U318 (N_318,In_1025,In_2471);
and U319 (N_319,In_1558,In_2675);
nor U320 (N_320,In_2806,In_1184);
and U321 (N_321,In_771,In_2536);
and U322 (N_322,In_556,In_2660);
or U323 (N_323,In_437,In_2511);
nand U324 (N_324,In_747,In_2039);
nor U325 (N_325,In_1445,In_87);
nor U326 (N_326,In_2916,In_1301);
or U327 (N_327,In_878,In_2107);
nor U328 (N_328,In_788,In_1004);
and U329 (N_329,In_677,In_2533);
nor U330 (N_330,In_2810,In_1830);
nand U331 (N_331,In_2062,In_417);
or U332 (N_332,In_683,In_2892);
or U333 (N_333,In_396,In_723);
or U334 (N_334,In_1543,In_2186);
nor U335 (N_335,In_354,In_1567);
xnor U336 (N_336,In_2037,In_47);
nor U337 (N_337,In_1400,In_530);
or U338 (N_338,In_220,In_267);
and U339 (N_339,In_261,In_867);
nor U340 (N_340,In_2154,In_85);
nor U341 (N_341,In_2839,In_1458);
or U342 (N_342,In_194,In_2317);
nor U343 (N_343,In_1028,In_2949);
nor U344 (N_344,In_2544,In_1487);
and U345 (N_345,In_1234,In_1030);
and U346 (N_346,In_2667,In_712);
and U347 (N_347,In_172,In_1357);
or U348 (N_348,In_2605,In_574);
nor U349 (N_349,In_930,In_519);
xnor U350 (N_350,In_2961,In_651);
nand U351 (N_351,In_2926,In_2980);
or U352 (N_352,In_974,In_2855);
xnor U353 (N_353,In_1013,In_1036);
or U354 (N_354,In_2478,In_522);
and U355 (N_355,In_1050,In_672);
and U356 (N_356,In_2456,In_421);
xnor U357 (N_357,In_1836,In_1037);
xor U358 (N_358,In_1617,In_1420);
nor U359 (N_359,In_711,In_802);
nand U360 (N_360,In_2978,In_222);
and U361 (N_361,In_2760,In_1660);
or U362 (N_362,In_1796,In_311);
and U363 (N_363,In_2480,In_2120);
and U364 (N_364,In_2678,In_185);
nor U365 (N_365,In_961,In_1099);
nand U366 (N_366,In_1436,In_2967);
xnor U367 (N_367,In_2458,In_591);
xor U368 (N_368,In_627,In_173);
and U369 (N_369,In_359,In_1913);
nand U370 (N_370,In_1808,In_2095);
nor U371 (N_371,In_2629,In_414);
xnor U372 (N_372,In_2083,In_786);
nand U373 (N_373,In_659,In_1372);
nor U374 (N_374,In_1049,In_600);
nand U375 (N_375,In_1399,In_1101);
and U376 (N_376,In_2064,In_1557);
or U377 (N_377,In_1326,In_2773);
and U378 (N_378,In_2426,In_1294);
nand U379 (N_379,In_388,In_737);
xnor U380 (N_380,In_2599,In_1225);
nor U381 (N_381,In_547,In_1067);
xnor U382 (N_382,In_726,In_2202);
nor U383 (N_383,In_2884,In_1158);
or U384 (N_384,In_2068,In_344);
or U385 (N_385,In_1467,In_2655);
and U386 (N_386,In_1148,In_709);
and U387 (N_387,In_772,In_2706);
xnor U388 (N_388,In_356,In_117);
or U389 (N_389,In_1051,In_2449);
nor U390 (N_390,In_1981,In_2836);
and U391 (N_391,In_2953,In_2738);
or U392 (N_392,In_1646,In_2278);
and U393 (N_393,In_1728,In_2649);
and U394 (N_394,In_1940,In_935);
and U395 (N_395,In_2508,In_2850);
nand U396 (N_396,In_1846,In_2938);
nand U397 (N_397,In_1138,In_757);
xor U398 (N_398,In_2575,In_2690);
nand U399 (N_399,In_2450,In_1571);
and U400 (N_400,In_1150,In_1033);
nor U401 (N_401,In_2345,In_2681);
and U402 (N_402,In_60,In_990);
nor U403 (N_403,In_2577,In_1576);
xnor U404 (N_404,In_2867,In_167);
and U405 (N_405,In_17,In_1793);
and U406 (N_406,In_2260,In_794);
xnor U407 (N_407,In_1705,In_762);
nand U408 (N_408,In_1038,In_2581);
xnor U409 (N_409,In_685,In_373);
or U410 (N_410,In_2846,In_2512);
and U411 (N_411,In_739,In_2754);
nand U412 (N_412,In_2647,In_2941);
nor U413 (N_413,In_2114,In_2238);
or U414 (N_414,In_833,In_1160);
nor U415 (N_415,In_2794,In_138);
nor U416 (N_416,In_2954,In_199);
and U417 (N_417,In_1387,In_2337);
nor U418 (N_418,In_1744,In_78);
nor U419 (N_419,In_2001,In_2972);
xor U420 (N_420,In_856,In_1272);
nand U421 (N_421,In_116,In_594);
and U422 (N_422,In_2950,In_2928);
or U423 (N_423,In_2294,In_446);
and U424 (N_424,In_1592,In_641);
nand U425 (N_425,In_465,In_2045);
xnor U426 (N_426,In_625,In_464);
or U427 (N_427,In_2711,In_2463);
and U428 (N_428,In_2870,In_1947);
and U429 (N_429,In_1577,In_1651);
nand U430 (N_430,In_1116,In_2714);
nand U431 (N_431,In_2586,In_545);
nor U432 (N_432,In_1362,In_773);
or U433 (N_433,In_2816,In_2462);
nand U434 (N_434,In_622,In_2563);
nand U435 (N_435,In_2825,In_916);
nand U436 (N_436,In_2644,In_2303);
and U437 (N_437,In_1710,In_2912);
and U438 (N_438,In_2819,In_1235);
nand U439 (N_439,In_1089,In_152);
nor U440 (N_440,In_330,In_2964);
nor U441 (N_441,In_2384,In_1555);
xnor U442 (N_442,In_20,In_1086);
nor U443 (N_443,In_2061,In_378);
nor U444 (N_444,In_968,In_653);
nor U445 (N_445,In_566,In_2944);
xor U446 (N_446,In_2199,In_2765);
and U447 (N_447,In_1419,In_2591);
xnor U448 (N_448,In_2287,In_2931);
and U449 (N_449,In_1681,In_1190);
nor U450 (N_450,In_1959,In_1268);
or U451 (N_451,In_399,In_1371);
and U452 (N_452,In_575,In_840);
nand U453 (N_453,In_2905,In_1201);
and U454 (N_454,In_2147,In_1090);
xor U455 (N_455,In_1992,In_1058);
nor U456 (N_456,In_2323,In_1654);
or U457 (N_457,In_2339,In_1338);
nor U458 (N_458,In_2922,In_807);
or U459 (N_459,In_1100,In_171);
nand U460 (N_460,In_541,In_2830);
and U461 (N_461,In_589,In_2399);
nor U462 (N_462,In_188,In_593);
or U463 (N_463,In_93,In_780);
or U464 (N_464,In_1513,In_428);
nand U465 (N_465,In_1674,In_2421);
nor U466 (N_466,In_1986,In_1634);
nor U467 (N_467,In_2325,In_2772);
or U468 (N_468,In_1792,In_789);
nand U469 (N_469,In_2175,In_2723);
and U470 (N_470,In_1054,In_1446);
and U471 (N_471,In_2677,In_448);
nor U472 (N_472,In_2390,In_439);
or U473 (N_473,In_2626,In_1526);
nor U474 (N_474,In_2111,In_2898);
xor U475 (N_475,In_225,In_866);
and U476 (N_476,In_100,In_2135);
or U477 (N_477,In_1912,In_2986);
nand U478 (N_478,In_2253,In_1355);
nand U479 (N_479,In_333,In_2437);
or U480 (N_480,In_1970,In_241);
and U481 (N_481,In_1962,In_76);
nand U482 (N_482,In_1163,In_884);
nand U483 (N_483,In_987,In_666);
and U484 (N_484,In_1549,In_215);
and U485 (N_485,In_992,In_1083);
nor U486 (N_486,In_933,In_1485);
nor U487 (N_487,In_2169,In_1891);
nor U488 (N_488,In_512,In_309);
nand U489 (N_489,In_102,In_1374);
or U490 (N_490,In_1659,In_1429);
nand U491 (N_491,In_1359,In_400);
or U492 (N_492,In_2279,In_1772);
xor U493 (N_493,In_1469,In_1449);
or U494 (N_494,In_2254,In_1496);
xor U495 (N_495,In_213,In_2609);
or U496 (N_496,In_725,In_2843);
xnor U497 (N_497,In_1897,In_1858);
nand U498 (N_498,In_2740,In_2194);
nor U499 (N_499,In_155,In_357);
nor U500 (N_500,In_2299,In_767);
or U501 (N_501,In_861,In_1554);
nand U502 (N_502,In_2495,In_2869);
xor U503 (N_503,In_201,In_2564);
xor U504 (N_504,In_490,In_1180);
nand U505 (N_505,In_887,In_903);
nor U506 (N_506,In_2113,In_1423);
and U507 (N_507,In_2624,In_2093);
or U508 (N_508,In_549,In_734);
or U509 (N_509,In_2259,In_883);
nor U510 (N_510,In_1503,In_815);
nand U511 (N_511,In_1611,In_1312);
or U512 (N_512,In_1084,In_555);
xnor U513 (N_513,In_1402,In_1639);
and U514 (N_514,In_2829,In_50);
xor U515 (N_515,In_1024,In_196);
and U516 (N_516,In_1609,In_2527);
nor U517 (N_517,In_463,In_303);
nand U518 (N_518,In_214,In_293);
nand U519 (N_519,In_449,In_1191);
nand U520 (N_520,In_2832,In_2367);
nor U521 (N_521,In_919,In_910);
and U522 (N_522,In_1106,In_1855);
xnor U523 (N_523,In_924,In_841);
or U524 (N_524,In_976,In_1869);
nor U525 (N_525,In_2638,In_2601);
nand U526 (N_526,In_999,In_2232);
nor U527 (N_527,In_970,In_2049);
xnor U528 (N_528,In_2021,In_169);
xor U529 (N_529,In_1497,In_2331);
or U530 (N_530,In_1735,In_2429);
nand U531 (N_531,In_80,In_1488);
xor U532 (N_532,In_2603,In_1586);
nor U533 (N_533,In_2957,In_1198);
or U534 (N_534,In_1872,In_1635);
nand U535 (N_535,In_2886,In_2727);
and U536 (N_536,In_1588,In_292);
xnor U537 (N_537,In_221,In_775);
xor U538 (N_538,In_2411,In_873);
and U539 (N_539,In_973,In_509);
xor U540 (N_540,In_621,In_617);
xnor U541 (N_541,In_2507,In_296);
xnor U542 (N_542,In_701,In_640);
and U543 (N_543,In_72,In_365);
and U544 (N_544,In_1053,In_1172);
xor U545 (N_545,In_978,In_342);
xor U546 (N_546,In_2805,In_655);
xor U547 (N_547,In_1859,In_2370);
or U548 (N_548,In_1061,In_375);
nor U549 (N_549,In_1688,In_1533);
and U550 (N_550,In_1578,In_2404);
or U551 (N_551,In_2580,In_206);
nand U552 (N_552,In_955,In_610);
or U553 (N_553,In_855,In_1337);
xnor U554 (N_554,In_12,In_2446);
xor U555 (N_555,In_2203,In_751);
nand U556 (N_556,In_1748,In_1368);
xor U557 (N_557,In_1975,In_2730);
or U558 (N_558,In_707,In_1266);
xnor U559 (N_559,In_2089,In_2901);
or U560 (N_560,In_581,In_1282);
nor U561 (N_561,In_741,In_695);
nand U562 (N_562,In_2600,In_2725);
and U563 (N_563,In_731,In_1507);
and U564 (N_564,In_1599,In_808);
and U565 (N_565,In_1480,In_1865);
or U566 (N_566,In_749,In_2402);
xnor U567 (N_567,In_688,In_1247);
xnor U568 (N_568,In_1902,In_2190);
and U569 (N_569,In_662,In_2070);
and U570 (N_570,In_1700,In_831);
nor U571 (N_571,In_1680,In_939);
nand U572 (N_572,In_1669,In_2621);
or U573 (N_573,In_750,In_2441);
nand U574 (N_574,In_2786,In_2128);
nor U575 (N_575,In_2180,In_765);
xnor U576 (N_576,In_2251,In_139);
and U577 (N_577,In_2427,In_2340);
and U578 (N_578,In_320,In_312);
xnor U579 (N_579,In_2758,In_36);
nand U580 (N_580,In_1179,In_2010);
xnor U581 (N_581,In_363,In_1060);
nor U582 (N_582,In_1009,In_480);
or U583 (N_583,In_544,In_1699);
nand U584 (N_584,In_1631,In_1570);
and U585 (N_585,In_1820,In_523);
nand U586 (N_586,In_255,In_73);
and U587 (N_587,In_501,In_722);
or U588 (N_588,In_285,In_1813);
xor U589 (N_589,In_232,In_2752);
nand U590 (N_590,In_402,In_2737);
nor U591 (N_591,In_1032,In_552);
xnor U592 (N_592,In_216,In_525);
xnor U593 (N_593,In_1857,In_2862);
and U594 (N_594,In_2878,In_1958);
and U595 (N_595,In_231,In_1819);
nor U596 (N_596,In_372,In_975);
and U597 (N_597,In_1714,In_45);
nand U598 (N_598,In_1270,In_355);
nor U599 (N_599,In_2492,In_2570);
or U600 (N_600,In_2891,In_800);
nor U601 (N_601,In_2267,In_2693);
or U602 (N_602,In_2418,In_1105);
nand U603 (N_603,In_1023,In_251);
and U604 (N_604,In_151,In_597);
xor U605 (N_605,In_1832,In_1134);
or U606 (N_606,In_472,In_48);
nor U607 (N_607,In_1126,In_543);
and U608 (N_608,In_2130,In_1287);
or U609 (N_609,In_2932,In_1085);
nand U610 (N_610,In_450,In_1645);
nand U611 (N_611,In_1623,In_1550);
or U612 (N_612,In_1717,In_2371);
nand U613 (N_613,In_2126,In_2223);
nor U614 (N_614,In_642,In_2679);
xor U615 (N_615,In_754,In_236);
nor U616 (N_616,In_1218,In_1630);
or U617 (N_617,In_2500,In_1026);
xnor U618 (N_618,In_1756,In_1661);
nor U619 (N_619,In_1195,In_2145);
nand U620 (N_620,In_2078,In_1798);
or U621 (N_621,In_2231,In_252);
xnor U622 (N_622,In_2447,In_2217);
xnor U623 (N_623,In_2395,In_2851);
nor U624 (N_624,In_948,In_1370);
and U625 (N_625,In_478,In_2314);
nor U626 (N_626,In_1088,In_3);
and U627 (N_627,In_1864,In_1142);
nor U628 (N_628,In_1120,In_1739);
nor U629 (N_629,In_805,In_2032);
or U630 (N_630,In_2753,In_1839);
and U631 (N_631,In_270,In_1649);
or U632 (N_632,In_598,In_1080);
nand U633 (N_633,In_1602,In_499);
xnor U634 (N_634,In_858,In_2995);
xor U635 (N_635,In_2783,In_1790);
xnor U636 (N_636,In_735,In_1233);
nor U637 (N_637,In_793,In_1206);
and U638 (N_638,In_2210,In_2241);
nor U639 (N_639,In_1708,In_1392);
xnor U640 (N_640,In_195,In_742);
or U641 (N_641,In_1942,In_86);
nor U642 (N_642,In_321,In_2640);
nand U643 (N_643,In_110,In_2416);
xnor U644 (N_644,In_1352,In_1173);
and U645 (N_645,In_361,In_1935);
or U646 (N_646,In_2140,In_799);
and U647 (N_647,In_535,In_2589);
nand U648 (N_648,In_2549,In_1668);
xnor U649 (N_649,In_2002,In_1604);
or U650 (N_650,In_118,In_515);
or U651 (N_651,In_35,In_380);
nor U652 (N_652,In_2595,In_1885);
xor U653 (N_653,In_1656,In_2712);
nor U654 (N_654,In_957,In_264);
nand U655 (N_655,In_1537,In_1375);
nor U656 (N_656,In_791,In_61);
nand U657 (N_657,In_233,In_2119);
and U658 (N_658,In_2543,In_1481);
nor U659 (N_659,In_1871,In_1512);
and U660 (N_660,In_1006,In_2628);
xnor U661 (N_661,In_2530,In_1632);
and U662 (N_662,In_964,In_801);
nor U663 (N_663,In_1424,In_2393);
and U664 (N_664,In_998,In_1219);
nand U665 (N_665,In_1361,In_2999);
and U666 (N_666,In_2682,In_1637);
nand U667 (N_667,In_1843,In_534);
nand U668 (N_668,In_184,In_326);
nor U669 (N_669,In_2689,In_550);
nor U670 (N_670,In_837,In_2556);
or U671 (N_671,In_1123,In_349);
nand U672 (N_672,In_1146,In_2245);
nor U673 (N_673,In_2664,In_2106);
nand U674 (N_674,In_797,In_2167);
or U675 (N_675,In_1275,In_674);
nand U676 (N_676,In_678,In_1450);
nand U677 (N_677,In_584,In_2579);
xnor U678 (N_678,In_419,In_1128);
xor U679 (N_679,In_83,In_839);
nor U680 (N_680,In_425,In_977);
and U681 (N_681,In_2110,In_2397);
nor U682 (N_682,In_569,In_2799);
or U683 (N_683,In_2283,In_2793);
nor U684 (N_684,In_2812,In_49);
and U685 (N_685,In_2782,In_1769);
and U686 (N_686,In_22,In_120);
xor U687 (N_687,In_1317,In_1015);
nand U688 (N_688,In_2435,In_950);
nor U689 (N_689,In_1224,In_2770);
xnor U690 (N_690,In_1591,In_1693);
or U691 (N_691,In_2247,In_2526);
nor U692 (N_692,In_1378,In_2940);
nor U693 (N_693,In_783,In_1622);
xor U694 (N_694,In_2687,In_646);
nand U695 (N_695,In_1517,In_637);
and U696 (N_696,In_395,In_2459);
nor U697 (N_697,In_1320,In_1293);
xnor U698 (N_698,In_1977,In_1587);
nor U699 (N_699,In_500,In_2505);
and U700 (N_700,In_2501,In_125);
xnor U701 (N_701,In_1801,In_2004);
and U702 (N_702,In_1621,In_1344);
xnor U703 (N_703,In_451,In_2041);
nand U704 (N_704,In_1768,In_2680);
and U705 (N_705,In_325,In_755);
nor U706 (N_706,In_2249,In_1290);
or U707 (N_707,In_2631,In_1367);
and U708 (N_708,In_362,In_2857);
nand U709 (N_709,In_2636,In_2596);
or U710 (N_710,In_1678,In_2958);
and U711 (N_711,In_728,In_644);
nor U712 (N_712,In_2550,In_1271);
nor U713 (N_713,In_1676,In_1875);
nor U714 (N_714,In_175,In_1928);
and U715 (N_715,In_2747,In_918);
and U716 (N_716,In_2207,In_2826);
nor U717 (N_717,In_2815,In_2476);
xor U718 (N_718,In_1703,In_2173);
or U719 (N_719,In_1389,In_2243);
and U720 (N_720,In_1418,In_826);
nor U721 (N_721,In_137,In_824);
and U722 (N_722,In_1724,In_1373);
xnor U723 (N_723,In_1725,In_1807);
and U724 (N_724,In_1581,In_2282);
xnor U725 (N_725,In_218,In_2567);
and U726 (N_726,In_1629,In_1822);
and U727 (N_727,In_1499,In_364);
xnor U728 (N_728,In_784,In_1221);
nor U729 (N_729,In_684,In_2308);
and U730 (N_730,In_24,In_9);
nor U731 (N_731,In_1974,In_19);
or U732 (N_732,In_1926,In_1267);
nand U733 (N_733,In_2979,In_1757);
nor U734 (N_734,In_2454,In_1314);
xor U735 (N_735,In_1057,In_1141);
and U736 (N_736,In_2178,In_1376);
nand U737 (N_737,In_1425,In_1147);
xor U738 (N_738,In_2082,In_2239);
nand U739 (N_739,In_2875,In_1823);
and U740 (N_740,In_1454,In_2984);
nor U741 (N_741,In_2022,In_1625);
and U742 (N_742,In_1563,In_63);
or U743 (N_743,In_828,In_2008);
nand U744 (N_744,In_163,In_460);
or U745 (N_745,In_2125,In_700);
or U746 (N_746,In_1189,In_2571);
and U747 (N_747,In_1421,In_648);
xnor U748 (N_748,In_33,In_2606);
or U749 (N_749,In_2559,In_1288);
nor U750 (N_750,In_2343,In_1127);
nand U751 (N_751,In_302,In_245);
nand U752 (N_752,In_2504,In_2143);
nor U753 (N_753,In_2256,In_2377);
and U754 (N_754,In_2166,In_1385);
nand U755 (N_755,In_1833,In_1334);
nand U756 (N_756,In_2277,In_415);
and U757 (N_757,In_2122,In_13);
nand U758 (N_758,In_2566,In_2457);
and U759 (N_759,In_2028,In_1806);
xnor U760 (N_760,In_2224,In_578);
and U761 (N_761,In_1197,In_1722);
nand U762 (N_762,In_226,In_1129);
nor U763 (N_763,In_1952,In_1401);
or U764 (N_764,In_1278,In_1948);
or U765 (N_765,In_1430,In_122);
xor U766 (N_766,In_224,In_1509);
and U767 (N_767,In_2197,In_2349);
nor U768 (N_768,In_53,In_620);
and U769 (N_769,In_2818,In_1895);
or U770 (N_770,In_1281,In_1667);
xnor U771 (N_771,In_1461,In_263);
nand U772 (N_772,In_1017,In_2510);
nor U773 (N_773,In_2187,In_2383);
xnor U774 (N_774,In_676,In_796);
and U775 (N_775,In_1615,In_518);
or U776 (N_776,In_1396,In_2248);
or U777 (N_777,In_1870,In_2117);
nor U778 (N_778,In_166,In_1273);
nand U779 (N_779,In_383,In_135);
or U780 (N_780,In_57,In_2852);
nand U781 (N_781,In_703,In_798);
nor U782 (N_782,In_259,In_2554);
nor U783 (N_783,In_2670,In_2084);
and U784 (N_784,In_2063,In_553);
and U785 (N_785,In_937,In_108);
nor U786 (N_786,In_894,In_2993);
xor U787 (N_787,In_2988,In_2461);
and U788 (N_788,In_2787,In_1069);
and U789 (N_789,In_1831,In_2802);
xor U790 (N_790,In_2914,In_2338);
nor U791 (N_791,In_862,In_2702);
xnor U792 (N_792,In_2489,In_743);
xnor U793 (N_793,In_1259,In_713);
nor U794 (N_794,In_1005,In_590);
xor U795 (N_795,In_2034,In_768);
or U796 (N_796,In_2403,In_5);
or U797 (N_797,In_1073,In_1746);
nand U798 (N_798,In_2479,In_2);
nand U799 (N_799,In_2910,In_1210);
nor U800 (N_800,In_68,In_129);
or U801 (N_801,In_2465,In_517);
xor U802 (N_802,In_2098,In_2475);
nor U803 (N_803,In_1884,In_1483);
and U804 (N_804,In_1111,In_1983);
xnor U805 (N_805,In_2023,In_2424);
and U806 (N_806,In_776,In_532);
or U807 (N_807,In_2761,In_299);
nand U808 (N_808,In_1476,In_993);
or U809 (N_809,In_2355,In_1236);
and U810 (N_810,In_1572,In_2423);
nor U811 (N_811,In_2177,In_940);
or U812 (N_812,In_2209,In_853);
nand U813 (N_813,In_1463,In_2152);
nor U814 (N_814,In_2198,In_632);
nand U815 (N_815,In_2043,In_1011);
nor U816 (N_816,In_1682,In_2375);
or U817 (N_817,In_2460,In_2176);
xor U818 (N_818,In_1763,In_2523);
and U819 (N_819,In_1156,In_350);
nor U820 (N_820,In_953,In_310);
nand U821 (N_821,In_1322,In_1967);
or U822 (N_822,In_1866,In_2669);
nand U823 (N_823,In_744,In_2102);
and U824 (N_824,In_2909,In_1741);
nor U825 (N_825,In_65,In_1457);
or U826 (N_826,In_385,In_1585);
and U827 (N_827,In_1532,In_331);
nand U828 (N_828,In_2746,In_2208);
or U829 (N_829,In_2301,In_2769);
and U830 (N_830,In_471,In_436);
and U831 (N_831,In_174,In_546);
xor U832 (N_832,In_2952,In_282);
nor U833 (N_833,In_2344,In_1335);
xor U834 (N_834,In_2962,In_1906);
nor U835 (N_835,In_718,In_1382);
nand U836 (N_836,In_2074,In_2612);
and U837 (N_837,In_2604,In_1304);
nor U838 (N_838,In_2674,In_1904);
nor U839 (N_839,In_698,In_2736);
xor U840 (N_840,In_803,In_1504);
nor U841 (N_841,In_1157,In_1031);
nor U842 (N_842,In_1415,In_2228);
or U843 (N_843,In_2904,In_1569);
xnor U844 (N_844,In_1738,In_2417);
and U845 (N_845,In_1444,In_1082);
nor U846 (N_846,In_2956,In_2075);
nor U847 (N_847,In_1118,In_2432);
and U848 (N_848,In_1723,In_337);
xor U849 (N_849,In_476,In_2362);
nand U850 (N_850,In_540,In_1726);
or U851 (N_851,In_2975,In_1518);
xor U852 (N_852,In_95,In_2132);
xor U853 (N_853,In_2118,In_1750);
nor U854 (N_854,In_1812,In_2431);
nand U855 (N_855,In_2519,In_691);
or U856 (N_856,In_1360,In_2161);
or U857 (N_857,In_680,In_2351);
or U858 (N_858,In_140,In_1743);
and U859 (N_859,In_2413,In_2837);
nor U860 (N_860,In_819,In_305);
and U861 (N_861,In_133,In_1112);
and U862 (N_862,In_2409,In_404);
nand U863 (N_863,In_34,In_187);
xnor U864 (N_864,In_2101,In_475);
xor U865 (N_865,In_397,In_343);
xnor U866 (N_866,In_322,In_2835);
and U867 (N_867,In_431,In_2035);
nand U868 (N_868,In_781,In_1285);
and U869 (N_869,In_623,In_1298);
or U870 (N_870,In_2436,In_2982);
and U871 (N_871,In_2439,In_2868);
nand U872 (N_872,In_2220,In_2650);
nor U873 (N_873,In_1564,In_576);
nor U874 (N_874,In_2937,In_1464);
or U875 (N_875,In_223,In_889);
nor U876 (N_876,In_2720,In_2930);
nand U877 (N_877,In_2493,In_182);
nand U878 (N_878,In_606,In_1850);
or U879 (N_879,In_2615,In_1965);
nand U880 (N_880,In_2296,In_2235);
or U881 (N_881,In_863,In_2585);
xnor U882 (N_882,In_1505,In_345);
nand U883 (N_883,In_1016,In_429);
nand U884 (N_884,In_1920,In_570);
and U885 (N_885,In_92,In_2633);
nor U886 (N_886,In_1413,In_1778);
and U887 (N_887,In_945,In_162);
nor U888 (N_888,In_1773,In_609);
nand U889 (N_889,In_1187,In_829);
xor U890 (N_890,In_921,In_960);
or U891 (N_891,In_2653,In_2743);
nor U892 (N_892,In_2718,In_661);
nor U893 (N_893,In_2033,In_1216);
or U894 (N_894,In_1280,In_2295);
and U895 (N_895,In_1110,In_119);
xnor U896 (N_896,In_178,In_1733);
and U897 (N_897,In_1478,In_2219);
xor U898 (N_898,In_2619,In_304);
or U899 (N_899,In_2316,In_1008);
nor U900 (N_900,In_2466,In_2469);
xnor U901 (N_901,In_2929,In_2899);
xnor U902 (N_902,In_2474,In_2728);
or U903 (N_903,In_2144,In_1493);
or U904 (N_904,In_168,In_443);
nand U905 (N_905,In_1608,In_1973);
and U906 (N_906,In_1169,In_1391);
xnor U907 (N_907,In_710,In_1752);
or U908 (N_908,In_1248,In_2470);
and U909 (N_909,In_2561,In_1815);
xnor U910 (N_910,In_1193,In_1186);
and U911 (N_911,In_1894,In_2359);
nor U912 (N_912,In_2472,In_1848);
nor U913 (N_913,In_1551,In_1404);
and U914 (N_914,In_1548,In_10);
xor U915 (N_915,In_1306,In_253);
nor U916 (N_916,In_382,In_2781);
or U917 (N_917,In_2987,In_932);
nor U918 (N_918,In_2524,In_870);
nor U919 (N_919,In_2464,In_746);
and U920 (N_920,In_2719,In_1330);
and U921 (N_921,In_785,In_2255);
and U922 (N_922,In_844,In_1995);
xnor U923 (N_923,In_67,In_1170);
nor U924 (N_924,In_1348,In_1047);
and U925 (N_925,In_2274,In_2528);
xor U926 (N_926,In_493,In_667);
nor U927 (N_927,In_891,In_979);
xnor U928 (N_928,In_121,In_2394);
or U929 (N_929,In_495,In_511);
nor U930 (N_930,In_203,In_988);
or U931 (N_931,In_307,In_2270);
nand U932 (N_932,In_2790,In_1264);
or U933 (N_933,In_1766,In_1495);
and U934 (N_934,In_2485,In_572);
or U935 (N_935,In_1524,In_1149);
xor U936 (N_936,In_2100,In_170);
or U937 (N_937,In_1573,In_565);
nand U938 (N_938,In_1706,In_2513);
or U939 (N_939,In_2484,In_2924);
or U940 (N_940,In_487,In_1122);
xnor U941 (N_941,In_1319,In_1091);
xnor U942 (N_942,In_2139,In_1861);
nand U943 (N_943,In_2092,In_2919);
xor U944 (N_944,In_875,In_2656);
nor U945 (N_945,In_2502,In_1800);
xor U946 (N_946,In_1470,In_1411);
or U947 (N_947,In_1010,In_1828);
nor U948 (N_948,In_1704,In_2127);
and U949 (N_949,In_2281,In_1070);
nor U950 (N_950,In_2369,In_962);
xnor U951 (N_951,In_670,In_2733);
nor U952 (N_952,In_668,In_2387);
and U953 (N_953,In_340,In_897);
and U954 (N_954,In_2809,In_1459);
xor U955 (N_955,In_497,In_394);
nand U956 (N_956,In_2434,In_1626);
nand U957 (N_957,In_193,In_1019);
xor U958 (N_958,In_1538,In_573);
or U959 (N_959,In_626,In_56);
or U960 (N_960,In_1075,In_2545);
and U961 (N_961,In_2654,In_1844);
or U962 (N_962,In_2583,In_1943);
nand U963 (N_963,In_1810,In_275);
nor U964 (N_964,In_1183,In_2731);
and U965 (N_965,In_39,In_2365);
xor U966 (N_966,In_412,In_913);
nor U967 (N_967,In_1405,In_645);
nor U968 (N_968,In_1531,In_2312);
nor U969 (N_969,In_1153,In_1440);
or U970 (N_970,In_2921,In_1021);
and U971 (N_971,In_1803,In_391);
or U972 (N_972,In_1985,In_1369);
nor U973 (N_973,In_2358,In_1439);
nand U974 (N_974,In_1584,In_1525);
nor U975 (N_975,In_1204,In_1874);
and U976 (N_976,In_2673,In_1552);
nand U977 (N_977,In_51,In_2767);
nor U978 (N_978,In_881,In_2755);
and U979 (N_979,In_1818,In_1506);
or U980 (N_980,In_1736,In_764);
nor U981 (N_981,In_1675,In_2780);
nand U982 (N_982,In_1363,In_1048);
nor U983 (N_983,In_1346,In_2845);
or U984 (N_984,In_257,In_317);
xor U985 (N_985,In_629,In_1683);
and U986 (N_986,In_2221,In_592);
or U987 (N_987,In_2181,In_2257);
and U988 (N_988,In_2529,In_2927);
xnor U989 (N_989,In_430,In_1289);
nand U990 (N_990,In_2745,In_585);
xor U991 (N_991,In_25,In_1887);
nor U992 (N_992,In_2762,In_969);
xor U993 (N_993,In_1466,In_1339);
or U994 (N_994,In_823,In_1880);
nor U995 (N_995,In_2123,In_2789);
xnor U996 (N_996,In_286,In_1696);
and U997 (N_997,In_704,In_1283);
and U998 (N_998,In_1460,In_105);
and U999 (N_999,In_458,In_507);
nor U1000 (N_1000,In_1690,In_2189);
or U1001 (N_1001,In_1644,In_1342);
nand U1002 (N_1002,In_2971,In_2025);
xor U1003 (N_1003,In_2206,In_11);
nand U1004 (N_1004,In_1917,In_1217);
or U1005 (N_1005,In_2748,In_2848);
or U1006 (N_1006,In_1903,In_503);
nor U1007 (N_1007,In_43,In_1269);
nand U1008 (N_1008,In_888,In_2630);
nand U1009 (N_1009,In_1612,In_1781);
nand U1010 (N_1010,In_124,In_1252);
and U1011 (N_1011,In_390,In_318);
nor U1012 (N_1012,In_2535,In_306);
or U1013 (N_1013,In_2713,In_2156);
xor U1014 (N_1014,In_1242,In_2691);
nand U1015 (N_1015,In_2380,In_2933);
xor U1016 (N_1016,In_413,In_314);
nand U1017 (N_1017,In_1296,In_2792);
nand U1018 (N_1018,In_656,In_2934);
nand U1019 (N_1019,In_103,In_2858);
or U1020 (N_1020,In_489,In_1207);
xor U1021 (N_1021,In_377,In_2392);
xor U1022 (N_1022,In_1366,In_2808);
nand U1023 (N_1023,In_2272,In_520);
xor U1024 (N_1024,In_452,In_687);
nand U1025 (N_1025,In_994,In_2204);
nor U1026 (N_1026,In_1946,In_1309);
xor U1027 (N_1027,In_244,In_1996);
and U1028 (N_1028,In_1484,In_2087);
nor U1029 (N_1029,In_58,In_1042);
xnor U1030 (N_1030,In_1168,In_1740);
nor U1031 (N_1031,In_2716,In_2864);
and U1032 (N_1032,In_2803,In_2784);
nor U1033 (N_1033,In_1442,In_2288);
xnor U1034 (N_1034,In_492,In_2907);
and U1035 (N_1035,In_947,In_238);
and U1036 (N_1036,In_2911,In_1056);
nand U1037 (N_1037,In_1452,In_756);
xor U1038 (N_1038,In_281,In_1816);
nor U1039 (N_1039,In_1133,In_1328);
xor U1040 (N_1040,In_1529,In_153);
nor U1041 (N_1041,In_42,In_2779);
and U1042 (N_1042,In_2521,In_1712);
nand U1043 (N_1043,In_2776,In_1838);
and U1044 (N_1044,In_234,In_1257);
nor U1045 (N_1045,In_438,In_561);
or U1046 (N_1046,In_2515,In_1718);
xnor U1047 (N_1047,In_2634,In_1802);
nor U1048 (N_1048,In_2229,In_938);
xnor U1049 (N_1049,In_418,In_468);
nand U1050 (N_1050,In_1695,In_2085);
and U1051 (N_1051,In_586,In_2889);
nor U1052 (N_1052,In_865,In_1145);
and U1053 (N_1053,In_1627,In_2333);
nor U1054 (N_1054,In_1274,In_1852);
nand U1055 (N_1055,In_690,In_628);
nand U1056 (N_1056,In_582,In_2388);
xnor U1057 (N_1057,In_1209,In_2841);
or U1058 (N_1058,In_1303,In_1161);
or U1059 (N_1059,In_657,In_1760);
nand U1060 (N_1060,In_2666,In_1343);
nand U1061 (N_1061,In_2943,In_1350);
or U1062 (N_1062,In_2842,In_1383);
or U1063 (N_1063,In_1534,In_984);
nand U1064 (N_1064,In_1582,In_1692);
and U1065 (N_1065,In_1045,In_2490);
nor U1066 (N_1066,In_934,In_614);
xor U1067 (N_1067,In_62,In_2887);
nor U1068 (N_1068,In_949,In_2172);
and U1069 (N_1069,In_1315,In_1327);
xor U1070 (N_1070,In_441,In_488);
xor U1071 (N_1071,In_2151,In_564);
and U1072 (N_1072,In_291,In_2134);
nor U1073 (N_1073,In_2657,In_2263);
and U1074 (N_1074,In_1972,In_2854);
nand U1075 (N_1075,In_2593,In_1341);
or U1076 (N_1076,In_1417,In_2795);
nand U1077 (N_1077,In_1477,In_156);
and U1078 (N_1078,In_790,In_1783);
or U1079 (N_1079,In_876,In_1251);
or U1080 (N_1080,In_1673,In_2565);
xor U1081 (N_1081,In_848,In_1437);
nor U1082 (N_1082,In_836,In_959);
nor U1083 (N_1083,In_2722,In_2148);
xnor U1084 (N_1084,In_482,In_1336);
and U1085 (N_1085,In_1999,In_2983);
nor U1086 (N_1086,In_1873,In_1701);
nor U1087 (N_1087,In_2353,In_2797);
or U1088 (N_1088,In_2648,In_846);
or U1089 (N_1089,In_758,In_2451);
xor U1090 (N_1090,In_1284,In_2056);
or U1091 (N_1091,In_1689,In_1107);
nor U1092 (N_1092,In_907,In_352);
xor U1093 (N_1093,In_705,In_1093);
or U1094 (N_1094,In_1078,In_2551);
or U1095 (N_1095,In_2320,In_2185);
nand U1096 (N_1096,In_2918,In_2129);
or U1097 (N_1097,In_2849,In_2665);
nand U1098 (N_1098,In_44,In_571);
or U1099 (N_1099,In_524,In_1789);
xor U1100 (N_1100,In_84,In_1388);
and U1101 (N_1101,In_2276,In_384);
or U1102 (N_1102,In_2894,In_1223);
nor U1103 (N_1103,In_1854,In_2881);
nand U1104 (N_1104,In_2430,In_271);
and U1105 (N_1105,In_835,In_2051);
and U1106 (N_1106,In_927,In_851);
and U1107 (N_1107,In_1961,In_639);
xnor U1108 (N_1108,In_229,In_1077);
nand U1109 (N_1109,In_2974,In_1096);
nor U1110 (N_1110,In_1408,In_211);
nor U1111 (N_1111,In_295,In_2271);
xor U1112 (N_1112,In_2304,In_2026);
or U1113 (N_1113,In_2319,In_2284);
and U1114 (N_1114,In_782,In_2044);
or U1115 (N_1115,In_2538,In_332);
nand U1116 (N_1116,In_1774,In_898);
nand U1117 (N_1117,In_2408,In_1364);
nand U1118 (N_1118,In_2594,In_652);
nor U1119 (N_1119,In_301,In_1159);
or U1120 (N_1120,In_1121,In_2821);
nand U1121 (N_1121,In_370,In_911);
and U1122 (N_1122,In_769,In_1072);
nand U1123 (N_1123,In_1922,In_996);
or U1124 (N_1124,In_2800,In_2328);
xnor U1125 (N_1125,In_588,In_2060);
or U1126 (N_1126,In_2017,In_2329);
xnor U1127 (N_1127,In_1479,In_1398);
nand U1128 (N_1128,In_2262,In_669);
or U1129 (N_1129,In_2030,In_821);
or U1130 (N_1130,In_2977,In_90);
and U1131 (N_1131,In_2141,In_207);
nor U1132 (N_1132,In_1302,In_180);
nand U1133 (N_1133,In_787,In_2179);
nand U1134 (N_1134,In_154,In_2546);
and U1135 (N_1135,In_2013,In_2109);
and U1136 (N_1136,In_1648,In_2116);
and U1137 (N_1137,In_2990,In_748);
xor U1138 (N_1138,In_2861,In_1598);
nor U1139 (N_1139,In_260,In_1566);
or U1140 (N_1140,In_1853,In_814);
nor U1141 (N_1141,In_2879,In_328);
nor U1142 (N_1142,In_1062,In_1672);
or U1143 (N_1143,In_1250,In_2880);
and U1144 (N_1144,In_2483,In_266);
nand U1145 (N_1145,In_2170,In_2050);
and U1146 (N_1146,In_1265,In_32);
and U1147 (N_1147,In_111,In_2547);
xnor U1148 (N_1148,In_1119,In_1641);
and U1149 (N_1149,In_1140,In_278);
or U1150 (N_1150,In_516,In_1727);
nand U1151 (N_1151,In_6,In_279);
nand U1152 (N_1152,In_1492,In_2391);
and U1153 (N_1153,In_1899,In_2096);
and U1154 (N_1154,In_2133,In_931);
or U1155 (N_1155,In_2683,In_1613);
and U1156 (N_1156,In_1817,In_2955);
and U1157 (N_1157,In_1351,In_1732);
or U1158 (N_1158,In_1640,In_1930);
nor U1159 (N_1159,In_983,In_2020);
xor U1160 (N_1160,In_832,In_1231);
xnor U1161 (N_1161,In_1412,In_989);
nand U1162 (N_1162,In_294,In_316);
nand U1163 (N_1163,In_1945,In_2335);
nor U1164 (N_1164,In_1795,In_1124);
xnor U1165 (N_1165,In_2077,In_1182);
nand U1166 (N_1166,In_1596,In_77);
xor U1167 (N_1167,In_392,In_696);
or U1168 (N_1168,In_2268,In_740);
or U1169 (N_1169,In_1137,In_1253);
nor U1170 (N_1170,In_2863,In_2700);
nor U1171 (N_1171,In_1786,In_868);
nand U1172 (N_1172,In_1597,In_2531);
or U1173 (N_1173,In_1881,In_250);
nor U1174 (N_1174,In_1954,In_228);
and U1175 (N_1175,In_2242,In_237);
nor U1176 (N_1176,In_1220,In_1347);
or U1177 (N_1177,In_1589,In_915);
xnor U1178 (N_1178,In_2174,In_2275);
or U1179 (N_1179,In_401,In_1299);
or U1180 (N_1180,In_2823,In_1229);
or U1181 (N_1181,In_2162,In_2622);
nand U1182 (N_1182,In_161,In_720);
nor U1183 (N_1183,In_2016,In_1232);
nor U1184 (N_1184,In_240,In_145);
nor U1185 (N_1185,In_1788,In_2305);
nand U1186 (N_1186,In_2945,In_2346);
nor U1187 (N_1187,In_1490,In_2285);
nor U1188 (N_1188,In_1092,In_2381);
nor U1189 (N_1189,In_2965,In_456);
or U1190 (N_1190,In_1065,In_1409);
or U1191 (N_1191,In_1456,In_587);
nand U1192 (N_1192,In_1007,In_2258);
nor U1193 (N_1193,In_901,In_131);
nor U1194 (N_1194,In_845,In_2155);
or U1195 (N_1195,In_2218,In_1003);
nor U1196 (N_1196,In_1969,In_398);
nand U1197 (N_1197,In_54,In_1167);
xor U1198 (N_1198,In_1103,In_895);
xor U1199 (N_1199,In_1878,In_929);
xnor U1200 (N_1200,In_615,In_1655);
xnor U1201 (N_1201,In_810,In_1102);
xnor U1202 (N_1202,In_1562,In_1579);
nand U1203 (N_1203,In_1761,In_353);
xor U1204 (N_1204,In_527,In_198);
xnor U1205 (N_1205,In_1698,In_1514);
or U1206 (N_1206,In_1662,In_1993);
nor U1207 (N_1207,In_697,In_1670);
xor U1208 (N_1208,In_843,In_1397);
xor U1209 (N_1209,In_618,In_560);
or U1210 (N_1210,In_227,In_160);
or U1211 (N_1211,In_1029,In_558);
nand U1212 (N_1212,In_2236,In_880);
or U1213 (N_1213,In_2291,In_902);
nor U1214 (N_1214,In_2182,In_2196);
and U1215 (N_1215,In_423,In_1001);
or U1216 (N_1216,In_882,In_123);
and U1217 (N_1217,In_922,In_2069);
nand U1218 (N_1218,In_854,In_2877);
and U1219 (N_1219,In_1384,In_2216);
nor U1220 (N_1220,In_189,In_1805);
nand U1221 (N_1221,In_890,In_16);
and U1222 (N_1222,In_2297,In_2131);
and U1223 (N_1223,In_1175,In_1711);
xnor U1224 (N_1224,In_483,In_1345);
nor U1225 (N_1225,In_1575,In_2058);
and U1226 (N_1226,In_38,In_812);
and U1227 (N_1227,In_528,In_1520);
or U1228 (N_1228,In_1527,In_23);
nand U1229 (N_1229,In_2214,In_1238);
nand U1230 (N_1230,In_1707,In_1228);
or U1231 (N_1231,In_2226,In_972);
xnor U1232 (N_1232,In_2936,In_2315);
or U1233 (N_1233,In_899,In_1758);
xor U1234 (N_1234,In_1547,In_1358);
or U1235 (N_1235,In_1380,In_1939);
nor U1236 (N_1236,In_339,In_2871);
or U1237 (N_1237,In_2568,In_928);
nand U1238 (N_1238,In_2872,In_760);
nor U1239 (N_1239,In_2777,In_1657);
xor U1240 (N_1240,In_2079,In_715);
nor U1241 (N_1241,In_2487,In_30);
and U1242 (N_1242,In_613,In_1590);
nand U1243 (N_1243,In_2052,In_2168);
xnor U1244 (N_1244,In_510,In_2099);
nor U1245 (N_1245,In_2960,In_2844);
nor U1246 (N_1246,In_2552,In_1540);
nor U1247 (N_1247,In_1192,In_896);
xor U1248 (N_1248,In_409,In_2948);
xor U1249 (N_1249,In_274,In_872);
nand U1250 (N_1250,In_612,In_381);
nand U1251 (N_1251,In_568,In_498);
xnor U1252 (N_1252,In_2833,In_2774);
nor U1253 (N_1253,In_149,In_1318);
xnor U1254 (N_1254,In_904,In_2055);
nor U1255 (N_1255,In_859,In_1171);
or U1256 (N_1256,In_2989,In_1944);
or U1257 (N_1257,In_849,In_2137);
and U1258 (N_1258,In_2420,In_2326);
nor U1259 (N_1259,In_79,In_2637);
nand U1260 (N_1260,In_2354,In_1491);
and U1261 (N_1261,In_2205,In_1702);
nand U1262 (N_1262,In_1687,In_1734);
nor U1263 (N_1263,In_2853,In_2227);
xnor U1264 (N_1264,In_1938,In_1755);
or U1265 (N_1265,In_1765,In_2324);
and U1266 (N_1266,In_2908,In_1546);
xor U1267 (N_1267,In_635,In_2042);
nor U1268 (N_1268,In_2124,In_2057);
or U1269 (N_1269,In_580,In_455);
or U1270 (N_1270,In_2040,In_2230);
nand U1271 (N_1271,In_1055,In_2347);
nor U1272 (N_1272,In_1559,In_2290);
nor U1273 (N_1273,In_1580,In_732);
and U1274 (N_1274,In_1771,In_551);
xor U1275 (N_1275,In_1834,In_971);
or U1276 (N_1276,In_351,In_2499);
xor U1277 (N_1277,In_636,In_126);
xor U1278 (N_1278,In_2164,In_1313);
or U1279 (N_1279,In_2697,In_759);
nor U1280 (N_1280,In_26,In_774);
xnor U1281 (N_1281,In_611,In_186);
nor U1282 (N_1282,In_1686,In_1934);
and U1283 (N_1283,In_91,In_2163);
xor U1284 (N_1284,In_1936,In_1323);
nand U1285 (N_1285,In_157,In_1767);
or U1286 (N_1286,In_1143,In_1356);
nand U1287 (N_1287,In_1494,In_2750);
nor U1288 (N_1288,In_2246,In_2509);
nor U1289 (N_1289,In_827,In_2240);
nand U1290 (N_1290,In_2452,In_539);
xor U1291 (N_1291,In_2497,In_323);
and U1292 (N_1292,In_1426,In_440);
or U1293 (N_1293,In_997,In_2165);
xor U1294 (N_1294,In_2036,In_1898);
nor U1295 (N_1295,In_909,In_2038);
and U1296 (N_1296,In_2192,In_1176);
xnor U1297 (N_1297,In_1968,In_2389);
or U1298 (N_1298,In_1500,In_682);
and U1299 (N_1299,In_1324,In_1035);
xor U1300 (N_1300,In_18,In_779);
nand U1301 (N_1301,In_1964,In_1394);
xor U1302 (N_1302,In_1988,In_605);
xor U1303 (N_1303,In_379,In_1164);
nor U1304 (N_1304,In_2885,In_1607);
and U1305 (N_1305,In_804,In_1835);
nand U1306 (N_1306,In_2659,In_729);
or U1307 (N_1307,In_1340,In_479);
and U1308 (N_1308,In_864,In_338);
xnor U1309 (N_1309,In_1208,In_2635);
nand U1310 (N_1310,In_1956,In_1780);
xor U1311 (N_1311,In_879,In_2097);
nor U1312 (N_1312,In_367,In_2573);
nand U1313 (N_1313,In_2658,In_2888);
nor U1314 (N_1314,In_692,In_2895);
or U1315 (N_1315,In_113,In_1079);
xnor U1316 (N_1316,In_1619,In_2707);
xor U1317 (N_1317,In_28,In_2067);
and U1318 (N_1318,In_150,In_1545);
xor U1319 (N_1319,In_2046,In_2318);
or U1320 (N_1320,In_369,In_2076);
nand U1321 (N_1321,In_96,In_2213);
xor U1322 (N_1322,In_717,In_410);
or U1323 (N_1323,In_2261,In_219);
or U1324 (N_1324,In_2300,In_753);
nor U1325 (N_1325,In_2407,In_967);
and U1326 (N_1326,In_2676,In_434);
and U1327 (N_1327,In_1034,In_1624);
xnor U1328 (N_1328,In_1910,In_1888);
nand U1329 (N_1329,In_2031,In_2625);
xnor U1330 (N_1330,In_1041,In_2602);
and U1331 (N_1331,In_2488,In_1643);
xnor U1332 (N_1332,In_1039,In_2009);
and U1333 (N_1333,In_2195,In_2618);
nand U1334 (N_1334,In_1933,In_1260);
and U1335 (N_1335,In_212,In_1925);
xnor U1336 (N_1336,In_55,In_1775);
nor U1337 (N_1337,In_2610,In_2373);
or U1338 (N_1338,In_1595,In_2661);
and U1339 (N_1339,In_1321,In_1892);
nand U1340 (N_1340,In_2054,In_2696);
xnor U1341 (N_1341,In_2798,In_2059);
and U1342 (N_1342,In_1955,In_1522);
or U1343 (N_1343,In_386,In_706);
nor U1344 (N_1344,In_2425,In_2607);
nor U1345 (N_1345,In_2412,In_2086);
nand U1346 (N_1346,In_761,In_1989);
xnor U1347 (N_1347,In_2734,In_952);
nand U1348 (N_1348,In_1896,In_1311);
xor U1349 (N_1349,In_671,In_98);
nand U1350 (N_1350,In_1620,In_1900);
nand U1351 (N_1351,In_1379,In_1211);
nor U1352 (N_1352,In_721,In_2018);
or U1353 (N_1353,In_208,In_2627);
nand U1354 (N_1354,In_1647,In_877);
nand U1355 (N_1355,In_147,In_1809);
nand U1356 (N_1356,In_112,In_1390);
and U1357 (N_1357,In_1713,In_730);
and U1358 (N_1358,In_2992,In_1308);
nor U1359 (N_1359,In_2233,In_1845);
nand U1360 (N_1360,In_143,In_1215);
nand U1361 (N_1361,In_892,In_2003);
and U1362 (N_1362,In_115,In_158);
xnor U1363 (N_1363,In_2153,In_2966);
and U1364 (N_1364,In_249,In_247);
and U1365 (N_1365,In_2847,In_956);
and U1366 (N_1366,In_557,In_7);
nand U1367 (N_1367,In_2005,In_2763);
and U1368 (N_1368,In_2341,In_2136);
and U1369 (N_1369,In_2080,In_1694);
xor U1370 (N_1370,In_1825,In_654);
nand U1371 (N_1371,In_283,In_658);
and U1372 (N_1372,In_2897,In_2856);
nor U1373 (N_1373,In_2684,In_2477);
nand U1374 (N_1374,In_2998,In_1203);
xnor U1375 (N_1375,In_2645,In_2668);
xnor U1376 (N_1376,In_146,In_1737);
nor U1377 (N_1377,In_2959,In_2970);
xor U1378 (N_1378,In_1448,In_1155);
nor U1379 (N_1379,In_308,In_442);
nand U1380 (N_1380,In_508,In_1353);
or U1381 (N_1381,In_2741,In_505);
xnor U1382 (N_1382,In_2374,In_1199);
nand U1383 (N_1383,In_192,In_177);
and U1384 (N_1384,In_444,In_2981);
or U1385 (N_1385,In_2709,In_2142);
nor U1386 (N_1386,In_2334,In_958);
nand U1387 (N_1387,In_1174,In_1932);
nand U1388 (N_1388,In_1462,In_2330);
nor U1389 (N_1389,In_2440,In_2222);
xnor U1390 (N_1390,In_2401,In_2616);
or U1391 (N_1391,In_109,In_2726);
nand U1392 (N_1392,In_1914,In_1305);
xor U1393 (N_1393,In_435,In_1043);
or U1394 (N_1394,In_2903,In_1403);
xor U1395 (N_1395,In_393,In_2662);
xor U1396 (N_1396,In_2029,In_2011);
and U1397 (N_1397,In_2065,In_1860);
nand U1398 (N_1398,In_2212,In_1510);
and U1399 (N_1399,In_1951,In_2103);
nor U1400 (N_1400,In_204,In_1468);
xor U1401 (N_1401,In_2071,In_1068);
and U1402 (N_1402,In_2686,In_1745);
xor U1403 (N_1403,In_433,In_2311);
nand U1404 (N_1404,In_494,In_1108);
or U1405 (N_1405,In_374,In_559);
and U1406 (N_1406,In_239,In_2225);
or U1407 (N_1407,In_2611,In_2614);
nand U1408 (N_1408,In_521,In_1691);
and U1409 (N_1409,In_1916,In_1685);
xnor U1410 (N_1410,In_1610,In_1991);
and U1411 (N_1411,In_335,In_1931);
nand U1412 (N_1412,In_2582,In_2739);
xnor U1413 (N_1413,In_2764,In_1821);
nand U1414 (N_1414,In_1715,In_0);
xor U1415 (N_1415,In_951,In_2900);
nor U1416 (N_1416,In_2481,In_1291);
nor U1417 (N_1417,In_2642,In_1332);
and U1418 (N_1418,In_164,In_1542);
nor U1419 (N_1419,In_963,In_906);
or U1420 (N_1420,In_1441,In_14);
nor U1421 (N_1421,In_1377,In_2732);
nor U1422 (N_1422,In_21,In_136);
and U1423 (N_1423,In_2105,In_447);
xor U1424 (N_1424,In_1139,In_1202);
nand U1425 (N_1425,In_1729,In_2890);
nand U1426 (N_1426,In_2171,In_1310);
or U1427 (N_1427,In_1633,In_1166);
and U1428 (N_1428,In_2494,In_1594);
nand U1429 (N_1429,In_486,In_2935);
and U1430 (N_1430,In_268,In_2560);
and U1431 (N_1431,In_2873,In_2361);
xnor U1432 (N_1432,In_485,In_647);
nor U1433 (N_1433,In_616,In_2506);
and U1434 (N_1434,In_2234,In_2138);
and U1435 (N_1435,In_319,In_514);
and U1436 (N_1436,In_2313,In_619);
or U1437 (N_1437,In_1979,In_360);
nand U1438 (N_1438,In_2264,In_1614);
nor U1439 (N_1439,In_2963,In_1246);
and U1440 (N_1440,In_936,In_2882);
xnor U1441 (N_1441,In_2158,In_1601);
xnor U1442 (N_1442,In_2699,In_1784);
xnor U1443 (N_1443,In_1628,In_1905);
and U1444 (N_1444,In_491,In_2548);
and U1445 (N_1445,In_1603,In_462);
and U1446 (N_1446,In_2553,In_1950);
and U1447 (N_1447,In_2874,In_148);
nand U1448 (N_1448,In_1679,In_1052);
and U1449 (N_1449,In_2048,In_71);
nor U1450 (N_1450,In_702,In_900);
or U1451 (N_1451,In_577,In_358);
nor U1452 (N_1452,In_2939,In_2569);
nor U1453 (N_1453,In_2775,In_1431);
nor U1454 (N_1454,In_1222,In_210);
and U1455 (N_1455,In_2710,In_2729);
xor U1456 (N_1456,In_2946,In_2651);
nor U1457 (N_1457,In_2302,In_745);
or U1458 (N_1458,In_2968,In_1438);
and U1459 (N_1459,In_2694,In_2364);
or U1460 (N_1460,In_2356,In_1258);
or U1461 (N_1461,In_681,In_914);
nand U1462 (N_1462,In_1261,In_2785);
nand U1463 (N_1463,In_603,In_327);
nor U1464 (N_1464,In_1987,In_2422);
nor U1465 (N_1465,In_2721,In_426);
nor U1466 (N_1466,In_416,In_70);
xor U1467 (N_1467,In_694,In_2121);
or U1468 (N_1468,In_289,In_2184);
nand U1469 (N_1469,In_1927,In_445);
and U1470 (N_1470,In_1642,In_1876);
nand U1471 (N_1471,In_280,In_1918);
nand U1472 (N_1472,In_1230,In_2385);
nor U1473 (N_1473,In_64,In_242);
or U1474 (N_1474,In_1132,In_795);
and U1475 (N_1475,In_2503,In_457);
and U1476 (N_1476,In_2072,In_2415);
nand U1477 (N_1477,In_1561,In_15);
or U1478 (N_1478,In_114,In_405);
nor U1479 (N_1479,In_1541,In_504);
and U1480 (N_1480,In_1990,In_2000);
nor U1481 (N_1481,In_2632,In_1125);
nor U1482 (N_1482,In_604,In_272);
xnor U1483 (N_1483,In_1244,In_2467);
or U1484 (N_1484,In_1406,In_2801);
and U1485 (N_1485,In_1181,In_2838);
and U1486 (N_1486,In_2443,In_243);
nand U1487 (N_1487,In_1583,In_82);
nand U1488 (N_1488,In_1893,In_664);
nor U1489 (N_1489,In_1262,In_387);
nor U1490 (N_1490,In_1177,In_1059);
nor U1491 (N_1491,In_2896,In_329);
and U1492 (N_1492,In_583,In_2542);
nand U1493 (N_1493,In_1465,In_2804);
or U1494 (N_1494,In_1040,In_599);
or U1495 (N_1495,In_1519,In_2188);
nor U1496 (N_1496,In_778,In_834);
nand U1497 (N_1497,In_1416,In_2705);
xor U1498 (N_1498,In_1237,In_595);
xor U1499 (N_1499,In_981,In_348);
and U1500 (N_1500,N_472,N_1227);
xnor U1501 (N_1501,N_381,N_61);
and U1502 (N_1502,N_1256,N_853);
nor U1503 (N_1503,N_768,N_88);
nor U1504 (N_1504,N_1281,N_288);
or U1505 (N_1505,N_886,N_12);
nand U1506 (N_1506,N_0,N_835);
and U1507 (N_1507,N_213,N_1312);
nand U1508 (N_1508,N_1289,N_1440);
nor U1509 (N_1509,N_58,N_916);
or U1510 (N_1510,N_1078,N_589);
xnor U1511 (N_1511,N_1496,N_1213);
or U1512 (N_1512,N_855,N_709);
nor U1513 (N_1513,N_161,N_441);
and U1514 (N_1514,N_964,N_374);
xor U1515 (N_1515,N_929,N_798);
or U1516 (N_1516,N_268,N_726);
or U1517 (N_1517,N_255,N_1446);
nand U1518 (N_1518,N_1303,N_222);
nand U1519 (N_1519,N_1058,N_465);
xor U1520 (N_1520,N_733,N_257);
and U1521 (N_1521,N_670,N_1450);
nand U1522 (N_1522,N_639,N_48);
nor U1523 (N_1523,N_1184,N_1234);
nand U1524 (N_1524,N_1403,N_749);
or U1525 (N_1525,N_773,N_1108);
or U1526 (N_1526,N_298,N_1352);
or U1527 (N_1527,N_907,N_1275);
xor U1528 (N_1528,N_29,N_637);
nor U1529 (N_1529,N_795,N_592);
and U1530 (N_1530,N_20,N_1123);
xnor U1531 (N_1531,N_883,N_112);
or U1532 (N_1532,N_574,N_411);
or U1533 (N_1533,N_201,N_157);
xnor U1534 (N_1534,N_1050,N_1170);
and U1535 (N_1535,N_276,N_126);
nor U1536 (N_1536,N_1410,N_1330);
xnor U1537 (N_1537,N_241,N_813);
and U1538 (N_1538,N_444,N_1262);
and U1539 (N_1539,N_32,N_1494);
or U1540 (N_1540,N_1044,N_753);
nor U1541 (N_1541,N_987,N_1358);
nand U1542 (N_1542,N_811,N_870);
or U1543 (N_1543,N_507,N_47);
nor U1544 (N_1544,N_777,N_363);
or U1545 (N_1545,N_1140,N_1382);
nor U1546 (N_1546,N_1096,N_707);
or U1547 (N_1547,N_718,N_921);
nand U1548 (N_1548,N_1128,N_1322);
nand U1549 (N_1549,N_346,N_851);
xnor U1550 (N_1550,N_1257,N_1197);
nand U1551 (N_1551,N_922,N_600);
xor U1552 (N_1552,N_1002,N_185);
nor U1553 (N_1553,N_1190,N_909);
or U1554 (N_1554,N_700,N_284);
xnor U1555 (N_1555,N_225,N_602);
nor U1556 (N_1556,N_857,N_1293);
nand U1557 (N_1557,N_5,N_817);
or U1558 (N_1558,N_1248,N_1138);
nand U1559 (N_1559,N_208,N_84);
nor U1560 (N_1560,N_515,N_859);
or U1561 (N_1561,N_1391,N_702);
xor U1562 (N_1562,N_1353,N_556);
xnor U1563 (N_1563,N_174,N_884);
or U1564 (N_1564,N_764,N_1119);
or U1565 (N_1565,N_349,N_1150);
nor U1566 (N_1566,N_1491,N_842);
xnor U1567 (N_1567,N_1431,N_575);
xnor U1568 (N_1568,N_933,N_117);
and U1569 (N_1569,N_214,N_1079);
and U1570 (N_1570,N_783,N_377);
xor U1571 (N_1571,N_1463,N_118);
xnor U1572 (N_1572,N_289,N_826);
nand U1573 (N_1573,N_1266,N_633);
and U1574 (N_1574,N_530,N_244);
and U1575 (N_1575,N_1042,N_337);
or U1576 (N_1576,N_119,N_999);
nor U1577 (N_1577,N_1471,N_1021);
nor U1578 (N_1578,N_429,N_442);
or U1579 (N_1579,N_123,N_1259);
nand U1580 (N_1580,N_1342,N_1393);
and U1581 (N_1581,N_1046,N_745);
xor U1582 (N_1582,N_784,N_1076);
nor U1583 (N_1583,N_182,N_1461);
and U1584 (N_1584,N_243,N_1339);
or U1585 (N_1585,N_997,N_1006);
nor U1586 (N_1586,N_199,N_1099);
or U1587 (N_1587,N_659,N_854);
or U1588 (N_1588,N_1204,N_548);
and U1589 (N_1589,N_164,N_1049);
nand U1590 (N_1590,N_1163,N_96);
and U1591 (N_1591,N_220,N_75);
or U1592 (N_1592,N_1287,N_821);
xnor U1593 (N_1593,N_620,N_1127);
xor U1594 (N_1594,N_1253,N_1378);
nand U1595 (N_1595,N_1379,N_62);
xor U1596 (N_1596,N_953,N_10);
or U1597 (N_1597,N_98,N_650);
xnor U1598 (N_1598,N_918,N_532);
nor U1599 (N_1599,N_168,N_673);
xnor U1600 (N_1600,N_1241,N_539);
xor U1601 (N_1601,N_800,N_323);
nand U1602 (N_1602,N_1026,N_1361);
and U1603 (N_1603,N_963,N_303);
and U1604 (N_1604,N_1242,N_1445);
xor U1605 (N_1605,N_756,N_1349);
or U1606 (N_1606,N_1404,N_196);
xnor U1607 (N_1607,N_1109,N_190);
nor U1608 (N_1608,N_551,N_277);
nor U1609 (N_1609,N_1484,N_451);
and U1610 (N_1610,N_45,N_209);
xor U1611 (N_1611,N_972,N_1004);
nand U1612 (N_1612,N_722,N_426);
or U1613 (N_1613,N_145,N_998);
or U1614 (N_1614,N_147,N_1413);
nand U1615 (N_1615,N_1177,N_934);
and U1616 (N_1616,N_1094,N_327);
nor U1617 (N_1617,N_1452,N_877);
or U1618 (N_1618,N_621,N_312);
and U1619 (N_1619,N_1301,N_1451);
and U1620 (N_1620,N_652,N_585);
and U1621 (N_1621,N_1149,N_200);
nand U1622 (N_1622,N_1251,N_17);
xor U1623 (N_1623,N_1316,N_1375);
or U1624 (N_1624,N_915,N_996);
nand U1625 (N_1625,N_1101,N_699);
and U1626 (N_1626,N_780,N_306);
nor U1627 (N_1627,N_81,N_1089);
or U1628 (N_1628,N_121,N_1203);
xnor U1629 (N_1629,N_986,N_634);
xnor U1630 (N_1630,N_1318,N_371);
or U1631 (N_1631,N_68,N_926);
xor U1632 (N_1632,N_1380,N_1386);
and U1633 (N_1633,N_177,N_344);
nand U1634 (N_1634,N_696,N_1146);
nand U1635 (N_1635,N_1070,N_719);
xnor U1636 (N_1636,N_341,N_1244);
xor U1637 (N_1637,N_1017,N_1037);
xor U1638 (N_1638,N_500,N_885);
nand U1639 (N_1639,N_601,N_927);
nand U1640 (N_1640,N_466,N_1456);
or U1641 (N_1641,N_1493,N_252);
and U1642 (N_1642,N_1336,N_1300);
xnor U1643 (N_1643,N_37,N_965);
nor U1644 (N_1644,N_829,N_26);
or U1645 (N_1645,N_408,N_1185);
nor U1646 (N_1646,N_1156,N_1284);
xor U1647 (N_1647,N_643,N_85);
xnor U1648 (N_1648,N_310,N_1286);
or U1649 (N_1649,N_1439,N_258);
nor U1650 (N_1650,N_1355,N_1229);
or U1651 (N_1651,N_4,N_1082);
nand U1652 (N_1652,N_526,N_412);
nor U1653 (N_1653,N_1181,N_171);
xnor U1654 (N_1654,N_528,N_1186);
or U1655 (N_1655,N_1106,N_361);
nor U1656 (N_1656,N_1205,N_1148);
and U1657 (N_1657,N_493,N_159);
or U1658 (N_1658,N_1290,N_490);
nor U1659 (N_1659,N_215,N_195);
nor U1660 (N_1660,N_597,N_937);
xnor U1661 (N_1661,N_815,N_140);
and U1662 (N_1662,N_744,N_906);
or U1663 (N_1663,N_486,N_852);
or U1664 (N_1664,N_1198,N_13);
xnor U1665 (N_1665,N_141,N_130);
nand U1666 (N_1666,N_1100,N_737);
xnor U1667 (N_1667,N_1480,N_967);
or U1668 (N_1668,N_116,N_1084);
or U1669 (N_1669,N_410,N_541);
nand U1670 (N_1670,N_1029,N_165);
and U1671 (N_1671,N_425,N_847);
and U1672 (N_1672,N_460,N_1160);
and U1673 (N_1673,N_33,N_1230);
xor U1674 (N_1674,N_446,N_66);
and U1675 (N_1675,N_770,N_137);
and U1676 (N_1676,N_1065,N_392);
xor U1677 (N_1677,N_248,N_1254);
nor U1678 (N_1678,N_1085,N_35);
and U1679 (N_1679,N_1191,N_698);
or U1680 (N_1680,N_15,N_259);
nor U1681 (N_1681,N_736,N_427);
nor U1682 (N_1682,N_475,N_588);
nand U1683 (N_1683,N_566,N_342);
and U1684 (N_1684,N_774,N_668);
or U1685 (N_1685,N_1299,N_318);
nor U1686 (N_1686,N_594,N_677);
xnor U1687 (N_1687,N_511,N_1436);
nand U1688 (N_1688,N_391,N_655);
nor U1689 (N_1689,N_1302,N_1053);
and U1690 (N_1690,N_343,N_1214);
xor U1691 (N_1691,N_1478,N_1343);
and U1692 (N_1692,N_582,N_1155);
or U1693 (N_1693,N_724,N_790);
and U1694 (N_1694,N_685,N_527);
nand U1695 (N_1695,N_1219,N_357);
and U1696 (N_1696,N_1143,N_1000);
and U1697 (N_1697,N_503,N_387);
nand U1698 (N_1698,N_524,N_1294);
and U1699 (N_1699,N_630,N_452);
nand U1700 (N_1700,N_1419,N_216);
nand U1701 (N_1701,N_115,N_192);
or U1702 (N_1702,N_521,N_665);
or U1703 (N_1703,N_1372,N_1488);
nand U1704 (N_1704,N_629,N_1189);
or U1705 (N_1705,N_207,N_474);
nor U1706 (N_1706,N_1088,N_928);
xnor U1707 (N_1707,N_1298,N_304);
and U1708 (N_1708,N_455,N_114);
or U1709 (N_1709,N_904,N_133);
nor U1710 (N_1710,N_1071,N_543);
nor U1711 (N_1711,N_1137,N_400);
or U1712 (N_1712,N_850,N_861);
xor U1713 (N_1713,N_890,N_499);
nor U1714 (N_1714,N_65,N_202);
or U1715 (N_1715,N_765,N_586);
and U1716 (N_1716,N_720,N_362);
nor U1717 (N_1717,N_1086,N_439);
xor U1718 (N_1718,N_791,N_966);
xor U1719 (N_1719,N_1485,N_666);
xor U1720 (N_1720,N_1033,N_492);
xor U1721 (N_1721,N_917,N_1272);
nand U1722 (N_1722,N_910,N_1060);
xor U1723 (N_1723,N_867,N_721);
xnor U1724 (N_1724,N_825,N_831);
and U1725 (N_1725,N_1247,N_148);
and U1726 (N_1726,N_135,N_804);
xnor U1727 (N_1727,N_172,N_271);
nand U1728 (N_1728,N_983,N_1048);
xnor U1729 (N_1729,N_43,N_42);
nor U1730 (N_1730,N_72,N_525);
and U1731 (N_1731,N_502,N_49);
nor U1732 (N_1732,N_674,N_664);
or U1733 (N_1733,N_739,N_1453);
or U1734 (N_1734,N_1279,N_865);
and U1735 (N_1735,N_1059,N_873);
or U1736 (N_1736,N_1359,N_266);
and U1737 (N_1737,N_1009,N_695);
nor U1738 (N_1738,N_1381,N_293);
nand U1739 (N_1739,N_734,N_275);
nand U1740 (N_1740,N_390,N_534);
or U1741 (N_1741,N_1310,N_1271);
xnor U1742 (N_1742,N_672,N_78);
or U1743 (N_1743,N_431,N_752);
or U1744 (N_1744,N_40,N_483);
xor U1745 (N_1745,N_833,N_1321);
nor U1746 (N_1746,N_1061,N_332);
or U1747 (N_1747,N_1144,N_540);
and U1748 (N_1748,N_1319,N_849);
nor U1749 (N_1749,N_616,N_805);
or U1750 (N_1750,N_892,N_338);
or U1751 (N_1751,N_1462,N_1005);
or U1752 (N_1752,N_605,N_100);
nand U1753 (N_1753,N_1398,N_944);
and U1754 (N_1754,N_836,N_1105);
nand U1755 (N_1755,N_863,N_82);
and U1756 (N_1756,N_505,N_1309);
nand U1757 (N_1757,N_754,N_254);
nor U1758 (N_1758,N_2,N_416);
nand U1759 (N_1759,N_1083,N_212);
or U1760 (N_1760,N_90,N_264);
and U1761 (N_1761,N_1092,N_260);
nor U1762 (N_1762,N_162,N_187);
xor U1763 (N_1763,N_728,N_478);
nor U1764 (N_1764,N_224,N_420);
xnor U1765 (N_1765,N_1187,N_1052);
nand U1766 (N_1766,N_529,N_1476);
nand U1767 (N_1767,N_1329,N_378);
nor U1768 (N_1768,N_705,N_227);
or U1769 (N_1769,N_1447,N_7);
or U1770 (N_1770,N_1387,N_691);
nor U1771 (N_1771,N_787,N_1276);
xor U1772 (N_1772,N_1296,N_1468);
nor U1773 (N_1773,N_314,N_287);
and U1774 (N_1774,N_569,N_463);
and U1775 (N_1775,N_622,N_393);
nor U1776 (N_1776,N_450,N_985);
or U1777 (N_1777,N_570,N_239);
or U1778 (N_1778,N_358,N_869);
xnor U1779 (N_1779,N_912,N_479);
nor U1780 (N_1780,N_626,N_579);
nand U1781 (N_1781,N_635,N_608);
nand U1782 (N_1782,N_1228,N_991);
nor U1783 (N_1783,N_714,N_485);
or U1784 (N_1784,N_1077,N_263);
and U1785 (N_1785,N_418,N_488);
xor U1786 (N_1786,N_1414,N_1067);
xor U1787 (N_1787,N_127,N_233);
nand U1788 (N_1788,N_373,N_644);
nand U1789 (N_1789,N_1133,N_1243);
nand U1790 (N_1790,N_91,N_1045);
and U1791 (N_1791,N_273,N_1420);
nand U1792 (N_1792,N_353,N_545);
xor U1793 (N_1793,N_1124,N_299);
nand U1794 (N_1794,N_546,N_560);
xnor U1795 (N_1795,N_975,N_1231);
xor U1796 (N_1796,N_671,N_710);
and U1797 (N_1797,N_830,N_992);
and U1798 (N_1798,N_1102,N_122);
and U1799 (N_1799,N_14,N_683);
or U1800 (N_1800,N_1240,N_487);
xor U1801 (N_1801,N_1348,N_1457);
xnor U1802 (N_1802,N_1364,N_181);
and U1803 (N_1803,N_129,N_1417);
nor U1804 (N_1804,N_766,N_267);
nor U1805 (N_1805,N_1104,N_1117);
nand U1806 (N_1806,N_236,N_464);
nor U1807 (N_1807,N_272,N_974);
nor U1808 (N_1808,N_802,N_154);
xnor U1809 (N_1809,N_428,N_1411);
nand U1810 (N_1810,N_661,N_1255);
nor U1811 (N_1811,N_237,N_1035);
nor U1812 (N_1812,N_941,N_1315);
nor U1813 (N_1813,N_593,N_368);
or U1814 (N_1814,N_134,N_1115);
xnor U1815 (N_1815,N_1154,N_175);
nand U1816 (N_1816,N_198,N_104);
xor U1817 (N_1817,N_1430,N_1020);
xor U1818 (N_1818,N_1014,N_150);
nor U1819 (N_1819,N_1278,N_1039);
and U1820 (N_1820,N_1224,N_1237);
nor U1821 (N_1821,N_102,N_1074);
xor U1822 (N_1822,N_1121,N_1483);
or U1823 (N_1823,N_348,N_1449);
nand U1824 (N_1824,N_269,N_846);
and U1825 (N_1825,N_1268,N_193);
nand U1826 (N_1826,N_249,N_1422);
nor U1827 (N_1827,N_581,N_39);
nor U1828 (N_1828,N_1261,N_1258);
xor U1829 (N_1829,N_956,N_191);
and U1830 (N_1830,N_583,N_519);
or U1831 (N_1831,N_1390,N_309);
nor U1832 (N_1832,N_1090,N_1209);
nor U1833 (N_1833,N_176,N_881);
nand U1834 (N_1834,N_615,N_701);
nand U1835 (N_1835,N_990,N_841);
nor U1836 (N_1836,N_1142,N_993);
nor U1837 (N_1837,N_603,N_1182);
nand U1838 (N_1838,N_59,N_989);
nand U1839 (N_1839,N_238,N_962);
or U1840 (N_1840,N_101,N_669);
or U1841 (N_1841,N_1377,N_895);
nand U1842 (N_1842,N_1428,N_1015);
xor U1843 (N_1843,N_523,N_1103);
nor U1844 (N_1844,N_415,N_935);
or U1845 (N_1845,N_291,N_839);
nor U1846 (N_1846,N_568,N_1054);
nand U1847 (N_1847,N_106,N_1384);
and U1848 (N_1848,N_845,N_509);
and U1849 (N_1849,N_470,N_1376);
nand U1850 (N_1850,N_1246,N_767);
and U1851 (N_1851,N_1098,N_54);
and U1852 (N_1852,N_1335,N_1345);
xor U1853 (N_1853,N_632,N_1110);
or U1854 (N_1854,N_206,N_960);
and U1855 (N_1855,N_1210,N_936);
or U1856 (N_1856,N_1273,N_375);
or U1857 (N_1857,N_1034,N_437);
xor U1858 (N_1858,N_366,N_471);
nand U1859 (N_1859,N_1194,N_1441);
xnor U1860 (N_1860,N_1129,N_1407);
nand U1861 (N_1861,N_432,N_223);
nand U1862 (N_1862,N_382,N_952);
nand U1863 (N_1863,N_1337,N_103);
or U1864 (N_1864,N_968,N_614);
nor U1865 (N_1865,N_913,N_41);
or U1866 (N_1866,N_781,N_55);
and U1867 (N_1867,N_1373,N_1196);
nand U1868 (N_1868,N_782,N_407);
or U1869 (N_1869,N_278,N_1306);
nor U1870 (N_1870,N_1135,N_796);
and U1871 (N_1871,N_402,N_607);
nand U1872 (N_1872,N_1388,N_775);
xnor U1873 (N_1873,N_786,N_105);
or U1874 (N_1874,N_1212,N_1317);
nor U1875 (N_1875,N_872,N_1486);
and U1876 (N_1876,N_856,N_1399);
xnor U1877 (N_1877,N_217,N_930);
xor U1878 (N_1878,N_875,N_414);
nand U1879 (N_1879,N_334,N_1164);
nand U1880 (N_1880,N_979,N_351);
nand U1881 (N_1881,N_294,N_868);
xor U1882 (N_1882,N_372,N_562);
nor U1883 (N_1883,N_1357,N_1490);
or U1884 (N_1884,N_792,N_751);
xnor U1885 (N_1885,N_1073,N_36);
or U1886 (N_1886,N_496,N_210);
xor U1887 (N_1887,N_1062,N_675);
nor U1888 (N_1888,N_1232,N_1166);
or U1889 (N_1889,N_571,N_1351);
nor U1890 (N_1890,N_183,N_1459);
or U1891 (N_1891,N_769,N_716);
nor U1892 (N_1892,N_297,N_226);
nor U1893 (N_1893,N_1003,N_1395);
or U1894 (N_1894,N_949,N_495);
xnor U1895 (N_1895,N_642,N_978);
or U1896 (N_1896,N_624,N_1469);
nor U1897 (N_1897,N_656,N_837);
and U1898 (N_1898,N_1499,N_1424);
or U1899 (N_1899,N_270,N_73);
nand U1900 (N_1900,N_1188,N_812);
xor U1901 (N_1901,N_16,N_506);
or U1902 (N_1902,N_572,N_23);
or U1903 (N_1903,N_1423,N_1113);
and U1904 (N_1904,N_827,N_794);
and U1905 (N_1905,N_557,N_189);
or U1906 (N_1906,N_347,N_584);
or U1907 (N_1907,N_328,N_128);
and U1908 (N_1908,N_77,N_717);
or U1909 (N_1909,N_553,N_283);
nor U1910 (N_1910,N_1027,N_247);
or U1911 (N_1911,N_1416,N_250);
nor U1912 (N_1912,N_1472,N_1016);
nor U1913 (N_1913,N_453,N_1282);
xor U1914 (N_1914,N_1013,N_604);
xnor U1915 (N_1915,N_840,N_689);
xor U1916 (N_1916,N_1385,N_340);
and U1917 (N_1917,N_435,N_1097);
nor U1918 (N_1918,N_1131,N_1460);
and U1919 (N_1919,N_538,N_1443);
and U1920 (N_1920,N_971,N_1314);
and U1921 (N_1921,N_1122,N_891);
nand U1922 (N_1922,N_379,N_1);
nand U1923 (N_1923,N_723,N_1285);
nand U1924 (N_1924,N_436,N_667);
xor U1925 (N_1925,N_305,N_1032);
and U1926 (N_1926,N_1206,N_771);
and U1927 (N_1927,N_370,N_71);
nor U1928 (N_1928,N_888,N_686);
nand U1929 (N_1929,N_1354,N_384);
nor U1930 (N_1930,N_413,N_564);
or U1931 (N_1931,N_711,N_552);
nand U1932 (N_1932,N_8,N_1183);
and U1933 (N_1933,N_676,N_163);
or U1934 (N_1934,N_120,N_645);
nor U1935 (N_1935,N_99,N_897);
and U1936 (N_1936,N_1208,N_433);
xnor U1937 (N_1937,N_38,N_1239);
nand U1938 (N_1938,N_1332,N_555);
nor U1939 (N_1939,N_1489,N_308);
xnor U1940 (N_1940,N_518,N_321);
and U1941 (N_1941,N_1167,N_1368);
and U1942 (N_1942,N_424,N_981);
nor U1943 (N_1943,N_27,N_461);
xor U1944 (N_1944,N_477,N_565);
nand U1945 (N_1945,N_793,N_882);
or U1946 (N_1946,N_1023,N_1292);
nor U1947 (N_1947,N_704,N_256);
or U1948 (N_1948,N_1169,N_919);
xor U1949 (N_1949,N_46,N_1400);
and U1950 (N_1950,N_322,N_834);
or U1951 (N_1951,N_326,N_285);
nor U1952 (N_1952,N_931,N_533);
nand U1953 (N_1953,N_755,N_520);
nand U1954 (N_1954,N_240,N_152);
and U1955 (N_1955,N_640,N_302);
nand U1956 (N_1956,N_1465,N_219);
nor U1957 (N_1957,N_1394,N_386);
or U1958 (N_1958,N_94,N_317);
nor U1959 (N_1959,N_1331,N_803);
or U1960 (N_1960,N_139,N_1371);
or U1961 (N_1961,N_893,N_83);
nand U1962 (N_1962,N_517,N_1217);
xnor U1963 (N_1963,N_1426,N_789);
nor U1964 (N_1964,N_712,N_596);
or U1965 (N_1965,N_491,N_1226);
and U1966 (N_1966,N_899,N_1307);
nor U1967 (N_1967,N_1161,N_876);
and U1968 (N_1968,N_409,N_727);
or U1969 (N_1969,N_591,N_959);
xnor U1970 (N_1970,N_482,N_434);
nand U1971 (N_1971,N_51,N_1324);
nand U1972 (N_1972,N_131,N_708);
nand U1973 (N_1973,N_738,N_394);
and U1974 (N_1974,N_544,N_1132);
xnor U1975 (N_1975,N_1047,N_973);
nor U1976 (N_1976,N_549,N_228);
nand U1977 (N_1977,N_653,N_497);
nor U1978 (N_1978,N_858,N_1432);
or U1979 (N_1979,N_898,N_900);
and U1980 (N_1980,N_619,N_567);
nor U1981 (N_1981,N_1173,N_443);
xor U1982 (N_1982,N_1220,N_292);
and U1983 (N_1983,N_184,N_1479);
or U1984 (N_1984,N_945,N_1093);
xnor U1985 (N_1985,N_300,N_1233);
and U1986 (N_1986,N_1136,N_142);
xor U1987 (N_1987,N_1201,N_662);
and U1988 (N_1988,N_489,N_1370);
xor U1989 (N_1989,N_692,N_138);
nor U1990 (N_1990,N_1277,N_628);
nor U1991 (N_1991,N_86,N_819);
or U1992 (N_1992,N_1091,N_24);
xor U1993 (N_1993,N_1218,N_820);
xnor U1994 (N_1994,N_136,N_143);
xor U1995 (N_1995,N_369,N_1326);
nor U1996 (N_1996,N_359,N_395);
xor U1997 (N_1997,N_1055,N_242);
and U1998 (N_1998,N_397,N_1141);
and U1999 (N_1999,N_611,N_818);
or U2000 (N_2000,N_245,N_1362);
nor U2001 (N_2001,N_69,N_1356);
xor U2002 (N_2002,N_958,N_180);
nor U2003 (N_2003,N_1374,N_403);
and U2004 (N_2004,N_1249,N_253);
nor U2005 (N_2005,N_335,N_1200);
or U2006 (N_2006,N_388,N_1360);
xnor U2007 (N_2007,N_1344,N_421);
or U2008 (N_2008,N_823,N_1111);
nor U2009 (N_2009,N_801,N_132);
or U2010 (N_2010,N_1025,N_367);
xor U2011 (N_2011,N_871,N_1069);
xnor U2012 (N_2012,N_160,N_398);
xor U2013 (N_2013,N_1291,N_1295);
nor U2014 (N_2014,N_896,N_1195);
and U2015 (N_2015,N_762,N_788);
or U2016 (N_2016,N_612,N_108);
or U2017 (N_2017,N_951,N_558);
nand U2018 (N_2018,N_481,N_301);
nor U2019 (N_2019,N_1406,N_1174);
xor U2020 (N_2020,N_325,N_1435);
nand U2021 (N_2021,N_550,N_679);
nand U2022 (N_2022,N_417,N_1147);
xnor U2023 (N_2023,N_943,N_1448);
xnor U2024 (N_2024,N_1001,N_1438);
xor U2025 (N_2025,N_1334,N_476);
or U2026 (N_2026,N_1180,N_438);
nand U2027 (N_2027,N_205,N_1482);
nor U2028 (N_2028,N_1120,N_1072);
and U2029 (N_2029,N_155,N_563);
nand U2030 (N_2030,N_204,N_824);
xnor U2031 (N_2031,N_1159,N_681);
or U2032 (N_2032,N_30,N_144);
xnor U2033 (N_2033,N_730,N_406);
nand U2034 (N_2034,N_844,N_295);
or U2035 (N_2035,N_331,N_862);
nor U2036 (N_2036,N_807,N_311);
and U2037 (N_2037,N_1207,N_504);
or U2038 (N_2038,N_1095,N_60);
nand U2039 (N_2039,N_468,N_64);
xor U2040 (N_2040,N_1270,N_419);
nand U2041 (N_2041,N_28,N_352);
nor U2042 (N_2042,N_561,N_889);
or U2043 (N_2043,N_1328,N_658);
and U2044 (N_2044,N_1225,N_947);
xnor U2045 (N_2045,N_942,N_1126);
or U2046 (N_2046,N_232,N_399);
xor U2047 (N_2047,N_364,N_687);
and U2048 (N_2048,N_262,N_731);
and U2049 (N_2049,N_660,N_1007);
and U2050 (N_2050,N_1475,N_946);
or U2051 (N_2051,N_810,N_146);
xnor U2052 (N_2052,N_158,N_230);
nand U2053 (N_2053,N_280,N_1288);
nand U2054 (N_2054,N_1112,N_1238);
nor U2055 (N_2055,N_153,N_1433);
or U2056 (N_2056,N_1019,N_536);
and U2057 (N_2057,N_961,N_110);
or U2058 (N_2058,N_107,N_1215);
nor U2059 (N_2059,N_623,N_1178);
xor U2060 (N_2060,N_1265,N_423);
xor U2061 (N_2061,N_954,N_537);
and U2062 (N_2062,N_984,N_587);
or U2063 (N_2063,N_1429,N_580);
nand U2064 (N_2064,N_1216,N_360);
xor U2065 (N_2065,N_1481,N_554);
nand U2066 (N_2066,N_1311,N_1418);
or U2067 (N_2067,N_1222,N_578);
and U2068 (N_2068,N_1158,N_678);
nand U2069 (N_2069,N_1415,N_1080);
nand U2070 (N_2070,N_87,N_448);
and U2071 (N_2071,N_860,N_785);
xnor U2072 (N_2072,N_447,N_950);
xnor U2073 (N_2073,N_814,N_590);
nor U2074 (N_2074,N_1434,N_1455);
nand U2075 (N_2075,N_599,N_1498);
xnor U2076 (N_2076,N_467,N_1350);
and U2077 (N_2077,N_422,N_290);
or U2078 (N_2078,N_50,N_67);
or U2079 (N_2079,N_976,N_315);
nor U2080 (N_2080,N_948,N_89);
nor U2081 (N_2081,N_1467,N_221);
or U2082 (N_2082,N_1041,N_761);
xnor U2083 (N_2083,N_380,N_166);
nand U2084 (N_2084,N_1260,N_808);
and U2085 (N_2085,N_21,N_151);
nand U2086 (N_2086,N_281,N_336);
xor U2087 (N_2087,N_1347,N_1068);
and U2088 (N_2088,N_229,N_79);
nor U2089 (N_2089,N_1341,N_806);
and U2090 (N_2090,N_354,N_1199);
and U2091 (N_2091,N_750,N_649);
and U2092 (N_2092,N_1157,N_879);
nand U2093 (N_2093,N_251,N_149);
nor U2094 (N_2094,N_648,N_778);
and U2095 (N_2095,N_1252,N_576);
xnor U2096 (N_2096,N_355,N_641);
xor U2097 (N_2097,N_908,N_235);
or U2098 (N_2098,N_779,N_279);
xnor U2099 (N_2099,N_535,N_547);
or U2100 (N_2100,N_169,N_1145);
or U2101 (N_2101,N_647,N_657);
nor U2102 (N_2102,N_1466,N_1162);
or U2103 (N_2103,N_457,N_878);
nand U2104 (N_2104,N_715,N_95);
or U2105 (N_2105,N_57,N_832);
xor U2106 (N_2106,N_449,N_809);
xnor U2107 (N_2107,N_1028,N_63);
or U2108 (N_2108,N_92,N_459);
xor U2109 (N_2109,N_194,N_97);
or U2110 (N_2110,N_1153,N_741);
or U2111 (N_2111,N_1038,N_383);
nand U2112 (N_2112,N_1018,N_1236);
and U2113 (N_2113,N_1269,N_109);
and U2114 (N_2114,N_1040,N_1363);
xor U2115 (N_2115,N_6,N_18);
or U2116 (N_2116,N_759,N_1168);
nor U2117 (N_2117,N_1125,N_1444);
nand U2118 (N_2118,N_9,N_982);
xnor U2119 (N_2119,N_940,N_1010);
or U2120 (N_2120,N_261,N_473);
nor U2121 (N_2121,N_1365,N_1396);
xor U2122 (N_2122,N_80,N_313);
or U2123 (N_2123,N_173,N_531);
nor U2124 (N_2124,N_735,N_1056);
nor U2125 (N_2125,N_350,N_1008);
or U2126 (N_2126,N_11,N_385);
xor U2127 (N_2127,N_559,N_1051);
nand U2128 (N_2128,N_1308,N_188);
nor U2129 (N_2129,N_1264,N_646);
xor U2130 (N_2130,N_508,N_203);
nor U2131 (N_2131,N_617,N_1030);
or U2132 (N_2132,N_498,N_939);
nand U2133 (N_2133,N_197,N_1130);
or U2134 (N_2134,N_1412,N_799);
nor U2135 (N_2135,N_693,N_1325);
nand U2136 (N_2136,N_932,N_329);
or U2137 (N_2137,N_828,N_1442);
and U2138 (N_2138,N_610,N_740);
nand U2139 (N_2139,N_1263,N_1474);
nand U2140 (N_2140,N_631,N_1202);
nand U2141 (N_2141,N_743,N_1392);
nor U2142 (N_2142,N_957,N_211);
or U2143 (N_2143,N_1297,N_1323);
nand U2144 (N_2144,N_1165,N_914);
or U2145 (N_2145,N_776,N_703);
and U2146 (N_2146,N_1011,N_1367);
and U2147 (N_2147,N_902,N_1402);
or U2148 (N_2148,N_440,N_980);
and U2149 (N_2149,N_1409,N_1081);
xor U2150 (N_2150,N_613,N_324);
or U2151 (N_2151,N_401,N_1346);
nor U2152 (N_2152,N_494,N_1024);
xnor U2153 (N_2153,N_955,N_430);
nor U2154 (N_2154,N_1464,N_1280);
xor U2155 (N_2155,N_838,N_246);
nor U2156 (N_2156,N_44,N_458);
and U2157 (N_2157,N_1333,N_843);
nand U2158 (N_2158,N_651,N_1211);
and U2159 (N_2159,N_1313,N_1107);
nand U2160 (N_2160,N_920,N_1458);
and U2161 (N_2161,N_1427,N_618);
nand U2162 (N_2162,N_1193,N_1383);
and U2163 (N_2163,N_772,N_113);
and U2164 (N_2164,N_333,N_1320);
and U2165 (N_2165,N_454,N_1172);
and U2166 (N_2166,N_1116,N_1340);
nand U2167 (N_2167,N_1389,N_1175);
xor U2168 (N_2168,N_1267,N_1031);
nand U2169 (N_2169,N_638,N_713);
xor U2170 (N_2170,N_1397,N_994);
or U2171 (N_2171,N_70,N_265);
nand U2172 (N_2172,N_682,N_680);
nor U2173 (N_2173,N_1064,N_816);
xnor U2174 (N_2174,N_1425,N_880);
and U2175 (N_2175,N_577,N_469);
nand U2176 (N_2176,N_690,N_1473);
nand U2177 (N_2177,N_1043,N_748);
nand U2178 (N_2178,N_725,N_501);
nand U2179 (N_2179,N_864,N_404);
or U2180 (N_2180,N_1497,N_763);
xor U2181 (N_2181,N_307,N_1235);
xnor U2182 (N_2182,N_627,N_179);
xnor U2183 (N_2183,N_988,N_510);
xor U2184 (N_2184,N_513,N_760);
nand U2185 (N_2185,N_522,N_286);
or U2186 (N_2186,N_911,N_1477);
and U2187 (N_2187,N_1274,N_925);
nand U2188 (N_2188,N_34,N_156);
and U2189 (N_2189,N_1192,N_19);
xnor U2190 (N_2190,N_684,N_977);
xnor U2191 (N_2191,N_25,N_445);
and U2192 (N_2192,N_595,N_654);
or U2193 (N_2193,N_218,N_376);
xnor U2194 (N_2194,N_1401,N_732);
or U2195 (N_2195,N_573,N_598);
nand U2196 (N_2196,N_1075,N_822);
xnor U2197 (N_2197,N_231,N_1221);
nor U2198 (N_2198,N_396,N_609);
and U2199 (N_2199,N_484,N_887);
and U2200 (N_2200,N_901,N_1114);
nor U2201 (N_2201,N_742,N_170);
nand U2202 (N_2202,N_1495,N_1118);
nand U2203 (N_2203,N_282,N_31);
and U2204 (N_2204,N_1405,N_1437);
nand U2205 (N_2205,N_76,N_516);
nand U2206 (N_2206,N_1304,N_514);
and U2207 (N_2207,N_405,N_1151);
nor U2208 (N_2208,N_1250,N_1338);
xnor U2209 (N_2209,N_706,N_52);
nand U2210 (N_2210,N_1421,N_694);
nor U2211 (N_2211,N_924,N_480);
nand U2212 (N_2212,N_1057,N_1063);
nor U2213 (N_2213,N_905,N_178);
nor U2214 (N_2214,N_1176,N_1492);
xor U2215 (N_2215,N_894,N_866);
xnor U2216 (N_2216,N_1179,N_167);
or U2217 (N_2217,N_697,N_316);
xnor U2218 (N_2218,N_1487,N_1327);
nor U2219 (N_2219,N_320,N_456);
nor U2220 (N_2220,N_111,N_186);
nand U2221 (N_2221,N_747,N_1036);
xor U2222 (N_2222,N_125,N_688);
nand U2223 (N_2223,N_758,N_389);
xor U2224 (N_2224,N_625,N_74);
or U2225 (N_2225,N_56,N_296);
or U2226 (N_2226,N_1305,N_356);
xnor U2227 (N_2227,N_969,N_938);
or U2228 (N_2228,N_797,N_1022);
xnor U2229 (N_2229,N_22,N_234);
nor U2230 (N_2230,N_542,N_757);
xnor U2231 (N_2231,N_995,N_512);
or U2232 (N_2232,N_339,N_462);
and U2233 (N_2233,N_3,N_606);
or U2234 (N_2234,N_1087,N_1470);
xor U2235 (N_2235,N_319,N_636);
and U2236 (N_2236,N_1171,N_729);
and U2237 (N_2237,N_1245,N_746);
nor U2238 (N_2238,N_923,N_1366);
or U2239 (N_2239,N_1012,N_1139);
xor U2240 (N_2240,N_124,N_53);
and U2241 (N_2241,N_903,N_330);
xor U2242 (N_2242,N_970,N_874);
and U2243 (N_2243,N_1152,N_663);
and U2244 (N_2244,N_1134,N_1454);
or U2245 (N_2245,N_1369,N_345);
nand U2246 (N_2246,N_274,N_93);
or U2247 (N_2247,N_1408,N_1223);
xnor U2248 (N_2248,N_1283,N_848);
nor U2249 (N_2249,N_1066,N_365);
or U2250 (N_2250,N_1073,N_570);
nand U2251 (N_2251,N_329,N_1167);
and U2252 (N_2252,N_1068,N_1275);
nand U2253 (N_2253,N_1068,N_1178);
or U2254 (N_2254,N_771,N_542);
xor U2255 (N_2255,N_1021,N_1232);
and U2256 (N_2256,N_927,N_850);
nand U2257 (N_2257,N_337,N_866);
nor U2258 (N_2258,N_10,N_859);
nand U2259 (N_2259,N_1321,N_576);
xnor U2260 (N_2260,N_1019,N_838);
and U2261 (N_2261,N_1255,N_232);
or U2262 (N_2262,N_471,N_433);
xnor U2263 (N_2263,N_582,N_39);
or U2264 (N_2264,N_273,N_225);
or U2265 (N_2265,N_1243,N_472);
and U2266 (N_2266,N_307,N_336);
and U2267 (N_2267,N_288,N_33);
xor U2268 (N_2268,N_879,N_185);
and U2269 (N_2269,N_662,N_186);
and U2270 (N_2270,N_796,N_4);
or U2271 (N_2271,N_5,N_483);
nand U2272 (N_2272,N_1292,N_19);
nand U2273 (N_2273,N_296,N_368);
or U2274 (N_2274,N_1050,N_122);
xor U2275 (N_2275,N_710,N_98);
nand U2276 (N_2276,N_551,N_140);
and U2277 (N_2277,N_760,N_529);
nand U2278 (N_2278,N_1441,N_1170);
nor U2279 (N_2279,N_986,N_331);
nand U2280 (N_2280,N_790,N_437);
nand U2281 (N_2281,N_617,N_698);
xor U2282 (N_2282,N_1281,N_701);
xor U2283 (N_2283,N_1169,N_657);
nand U2284 (N_2284,N_1465,N_1350);
nand U2285 (N_2285,N_276,N_322);
and U2286 (N_2286,N_1489,N_571);
nand U2287 (N_2287,N_10,N_1356);
xor U2288 (N_2288,N_1474,N_1052);
nand U2289 (N_2289,N_325,N_9);
and U2290 (N_2290,N_1492,N_1093);
xor U2291 (N_2291,N_829,N_1491);
xnor U2292 (N_2292,N_1492,N_870);
nand U2293 (N_2293,N_126,N_113);
or U2294 (N_2294,N_397,N_1468);
xnor U2295 (N_2295,N_473,N_1134);
and U2296 (N_2296,N_1329,N_966);
nand U2297 (N_2297,N_153,N_935);
or U2298 (N_2298,N_329,N_132);
and U2299 (N_2299,N_1393,N_457);
or U2300 (N_2300,N_340,N_18);
nor U2301 (N_2301,N_363,N_1100);
xor U2302 (N_2302,N_139,N_1450);
nor U2303 (N_2303,N_481,N_8);
and U2304 (N_2304,N_1325,N_1243);
or U2305 (N_2305,N_1408,N_911);
or U2306 (N_2306,N_1029,N_1268);
nand U2307 (N_2307,N_1315,N_119);
or U2308 (N_2308,N_252,N_106);
or U2309 (N_2309,N_73,N_852);
xnor U2310 (N_2310,N_1197,N_1187);
xnor U2311 (N_2311,N_454,N_394);
nor U2312 (N_2312,N_796,N_1408);
xnor U2313 (N_2313,N_1000,N_36);
nor U2314 (N_2314,N_882,N_1089);
nand U2315 (N_2315,N_1075,N_192);
xnor U2316 (N_2316,N_139,N_1027);
or U2317 (N_2317,N_338,N_988);
xor U2318 (N_2318,N_1019,N_953);
nand U2319 (N_2319,N_897,N_609);
nand U2320 (N_2320,N_1329,N_774);
or U2321 (N_2321,N_875,N_1170);
and U2322 (N_2322,N_401,N_1114);
xnor U2323 (N_2323,N_1451,N_475);
nand U2324 (N_2324,N_1223,N_1493);
and U2325 (N_2325,N_45,N_104);
nand U2326 (N_2326,N_74,N_1160);
or U2327 (N_2327,N_93,N_1102);
or U2328 (N_2328,N_910,N_531);
or U2329 (N_2329,N_1132,N_1422);
nand U2330 (N_2330,N_1409,N_1118);
nor U2331 (N_2331,N_790,N_775);
nand U2332 (N_2332,N_1056,N_778);
nor U2333 (N_2333,N_1048,N_60);
and U2334 (N_2334,N_661,N_282);
and U2335 (N_2335,N_549,N_100);
nor U2336 (N_2336,N_484,N_463);
xnor U2337 (N_2337,N_1349,N_865);
and U2338 (N_2338,N_236,N_719);
or U2339 (N_2339,N_1055,N_3);
nand U2340 (N_2340,N_617,N_1380);
nand U2341 (N_2341,N_255,N_948);
nand U2342 (N_2342,N_1435,N_329);
nand U2343 (N_2343,N_1173,N_452);
or U2344 (N_2344,N_257,N_1167);
and U2345 (N_2345,N_0,N_887);
nor U2346 (N_2346,N_27,N_355);
and U2347 (N_2347,N_305,N_1024);
and U2348 (N_2348,N_1119,N_645);
nor U2349 (N_2349,N_778,N_403);
nand U2350 (N_2350,N_179,N_1401);
nor U2351 (N_2351,N_708,N_1120);
xnor U2352 (N_2352,N_319,N_43);
nand U2353 (N_2353,N_1181,N_541);
xor U2354 (N_2354,N_4,N_1016);
nor U2355 (N_2355,N_75,N_1162);
or U2356 (N_2356,N_447,N_551);
nor U2357 (N_2357,N_612,N_807);
and U2358 (N_2358,N_1366,N_509);
and U2359 (N_2359,N_879,N_465);
or U2360 (N_2360,N_176,N_647);
and U2361 (N_2361,N_181,N_348);
or U2362 (N_2362,N_406,N_1059);
xor U2363 (N_2363,N_1377,N_99);
nand U2364 (N_2364,N_1254,N_1491);
nor U2365 (N_2365,N_33,N_27);
and U2366 (N_2366,N_7,N_1192);
and U2367 (N_2367,N_413,N_504);
nor U2368 (N_2368,N_975,N_1417);
and U2369 (N_2369,N_873,N_835);
and U2370 (N_2370,N_74,N_168);
and U2371 (N_2371,N_596,N_1282);
nand U2372 (N_2372,N_471,N_108);
xor U2373 (N_2373,N_175,N_270);
nor U2374 (N_2374,N_1342,N_171);
or U2375 (N_2375,N_590,N_791);
nor U2376 (N_2376,N_106,N_1403);
and U2377 (N_2377,N_733,N_1377);
and U2378 (N_2378,N_186,N_433);
nand U2379 (N_2379,N_66,N_170);
and U2380 (N_2380,N_1071,N_385);
xor U2381 (N_2381,N_538,N_1282);
nand U2382 (N_2382,N_1128,N_1138);
or U2383 (N_2383,N_40,N_1271);
and U2384 (N_2384,N_394,N_251);
or U2385 (N_2385,N_544,N_941);
nor U2386 (N_2386,N_1003,N_733);
xor U2387 (N_2387,N_622,N_1438);
nor U2388 (N_2388,N_834,N_712);
or U2389 (N_2389,N_1393,N_887);
and U2390 (N_2390,N_152,N_355);
and U2391 (N_2391,N_686,N_1428);
nor U2392 (N_2392,N_1295,N_715);
and U2393 (N_2393,N_1452,N_1339);
and U2394 (N_2394,N_526,N_929);
and U2395 (N_2395,N_35,N_421);
xor U2396 (N_2396,N_197,N_302);
or U2397 (N_2397,N_1212,N_790);
nor U2398 (N_2398,N_857,N_508);
nor U2399 (N_2399,N_555,N_948);
and U2400 (N_2400,N_827,N_87);
or U2401 (N_2401,N_694,N_225);
xor U2402 (N_2402,N_574,N_967);
and U2403 (N_2403,N_955,N_624);
xnor U2404 (N_2404,N_534,N_1340);
xnor U2405 (N_2405,N_666,N_1368);
and U2406 (N_2406,N_538,N_546);
nor U2407 (N_2407,N_105,N_622);
nand U2408 (N_2408,N_1039,N_801);
and U2409 (N_2409,N_1196,N_831);
nor U2410 (N_2410,N_1390,N_425);
nor U2411 (N_2411,N_1295,N_969);
and U2412 (N_2412,N_1496,N_1015);
nor U2413 (N_2413,N_741,N_785);
and U2414 (N_2414,N_982,N_907);
nand U2415 (N_2415,N_307,N_1206);
and U2416 (N_2416,N_775,N_681);
or U2417 (N_2417,N_174,N_662);
nor U2418 (N_2418,N_275,N_1367);
nor U2419 (N_2419,N_305,N_1047);
nand U2420 (N_2420,N_182,N_763);
and U2421 (N_2421,N_1254,N_846);
and U2422 (N_2422,N_876,N_1362);
and U2423 (N_2423,N_1166,N_606);
or U2424 (N_2424,N_1325,N_489);
or U2425 (N_2425,N_594,N_615);
and U2426 (N_2426,N_1449,N_1147);
nor U2427 (N_2427,N_1267,N_624);
or U2428 (N_2428,N_1171,N_872);
or U2429 (N_2429,N_1046,N_1095);
or U2430 (N_2430,N_27,N_1413);
nor U2431 (N_2431,N_817,N_1400);
nand U2432 (N_2432,N_69,N_885);
nor U2433 (N_2433,N_1412,N_1246);
and U2434 (N_2434,N_1179,N_1320);
and U2435 (N_2435,N_1156,N_128);
or U2436 (N_2436,N_5,N_254);
nor U2437 (N_2437,N_1322,N_1290);
and U2438 (N_2438,N_1036,N_890);
or U2439 (N_2439,N_50,N_1454);
nand U2440 (N_2440,N_651,N_958);
nor U2441 (N_2441,N_1063,N_278);
xor U2442 (N_2442,N_1039,N_673);
and U2443 (N_2443,N_1120,N_155);
and U2444 (N_2444,N_1331,N_219);
xor U2445 (N_2445,N_1050,N_1279);
or U2446 (N_2446,N_618,N_112);
and U2447 (N_2447,N_539,N_1149);
or U2448 (N_2448,N_152,N_728);
nand U2449 (N_2449,N_1013,N_874);
and U2450 (N_2450,N_1354,N_1128);
nand U2451 (N_2451,N_339,N_1312);
nor U2452 (N_2452,N_1186,N_192);
and U2453 (N_2453,N_557,N_431);
or U2454 (N_2454,N_1031,N_1113);
xnor U2455 (N_2455,N_195,N_144);
or U2456 (N_2456,N_759,N_1102);
and U2457 (N_2457,N_205,N_1025);
nand U2458 (N_2458,N_774,N_459);
and U2459 (N_2459,N_606,N_1436);
and U2460 (N_2460,N_622,N_463);
and U2461 (N_2461,N_832,N_1306);
xor U2462 (N_2462,N_1058,N_1082);
xor U2463 (N_2463,N_1183,N_654);
xnor U2464 (N_2464,N_517,N_522);
nand U2465 (N_2465,N_409,N_35);
nor U2466 (N_2466,N_200,N_923);
and U2467 (N_2467,N_798,N_837);
and U2468 (N_2468,N_214,N_147);
nor U2469 (N_2469,N_438,N_1007);
nand U2470 (N_2470,N_367,N_1250);
nand U2471 (N_2471,N_982,N_959);
or U2472 (N_2472,N_1499,N_1019);
or U2473 (N_2473,N_1280,N_300);
xnor U2474 (N_2474,N_930,N_842);
or U2475 (N_2475,N_1134,N_1339);
nor U2476 (N_2476,N_83,N_1036);
nor U2477 (N_2477,N_160,N_310);
nand U2478 (N_2478,N_984,N_1377);
and U2479 (N_2479,N_1158,N_393);
or U2480 (N_2480,N_438,N_277);
nor U2481 (N_2481,N_1483,N_1031);
nor U2482 (N_2482,N_522,N_743);
or U2483 (N_2483,N_1332,N_1238);
xor U2484 (N_2484,N_494,N_673);
or U2485 (N_2485,N_622,N_935);
or U2486 (N_2486,N_855,N_1070);
nor U2487 (N_2487,N_545,N_519);
or U2488 (N_2488,N_1224,N_767);
xnor U2489 (N_2489,N_1363,N_891);
and U2490 (N_2490,N_495,N_911);
nand U2491 (N_2491,N_1323,N_420);
xor U2492 (N_2492,N_74,N_530);
and U2493 (N_2493,N_1071,N_665);
xnor U2494 (N_2494,N_407,N_278);
nor U2495 (N_2495,N_1282,N_744);
nand U2496 (N_2496,N_267,N_706);
or U2497 (N_2497,N_1473,N_251);
nand U2498 (N_2498,N_377,N_78);
nor U2499 (N_2499,N_985,N_342);
xnor U2500 (N_2500,N_495,N_738);
nor U2501 (N_2501,N_1486,N_485);
and U2502 (N_2502,N_616,N_542);
or U2503 (N_2503,N_362,N_1213);
nor U2504 (N_2504,N_610,N_1213);
xor U2505 (N_2505,N_952,N_37);
or U2506 (N_2506,N_1099,N_578);
nand U2507 (N_2507,N_1366,N_336);
or U2508 (N_2508,N_722,N_86);
or U2509 (N_2509,N_846,N_270);
or U2510 (N_2510,N_984,N_116);
nor U2511 (N_2511,N_737,N_1441);
nor U2512 (N_2512,N_832,N_717);
xnor U2513 (N_2513,N_535,N_948);
nand U2514 (N_2514,N_267,N_148);
xnor U2515 (N_2515,N_72,N_619);
and U2516 (N_2516,N_1493,N_397);
and U2517 (N_2517,N_176,N_264);
xnor U2518 (N_2518,N_863,N_564);
and U2519 (N_2519,N_1483,N_140);
and U2520 (N_2520,N_483,N_444);
and U2521 (N_2521,N_534,N_823);
nand U2522 (N_2522,N_1047,N_177);
or U2523 (N_2523,N_1487,N_1443);
xnor U2524 (N_2524,N_1162,N_1425);
xor U2525 (N_2525,N_1161,N_517);
nand U2526 (N_2526,N_210,N_464);
nor U2527 (N_2527,N_600,N_1198);
xnor U2528 (N_2528,N_1232,N_446);
nand U2529 (N_2529,N_864,N_375);
xor U2530 (N_2530,N_1497,N_208);
xor U2531 (N_2531,N_602,N_492);
and U2532 (N_2532,N_991,N_467);
or U2533 (N_2533,N_87,N_64);
and U2534 (N_2534,N_632,N_1023);
nor U2535 (N_2535,N_806,N_762);
nand U2536 (N_2536,N_517,N_793);
or U2537 (N_2537,N_181,N_80);
nor U2538 (N_2538,N_204,N_1251);
or U2539 (N_2539,N_47,N_938);
and U2540 (N_2540,N_857,N_705);
xor U2541 (N_2541,N_1161,N_1423);
or U2542 (N_2542,N_1389,N_749);
nor U2543 (N_2543,N_408,N_225);
nor U2544 (N_2544,N_1191,N_973);
nor U2545 (N_2545,N_899,N_732);
xor U2546 (N_2546,N_924,N_221);
or U2547 (N_2547,N_518,N_1278);
and U2548 (N_2548,N_558,N_1176);
nand U2549 (N_2549,N_1254,N_984);
and U2550 (N_2550,N_752,N_994);
and U2551 (N_2551,N_1443,N_1098);
or U2552 (N_2552,N_407,N_1129);
and U2553 (N_2553,N_797,N_1011);
nor U2554 (N_2554,N_871,N_1076);
nor U2555 (N_2555,N_1172,N_364);
nor U2556 (N_2556,N_546,N_1350);
nor U2557 (N_2557,N_1386,N_1431);
and U2558 (N_2558,N_1368,N_1444);
xnor U2559 (N_2559,N_838,N_1326);
nor U2560 (N_2560,N_647,N_627);
or U2561 (N_2561,N_807,N_168);
nor U2562 (N_2562,N_227,N_781);
xnor U2563 (N_2563,N_889,N_1337);
nor U2564 (N_2564,N_1140,N_579);
xnor U2565 (N_2565,N_630,N_1121);
or U2566 (N_2566,N_1069,N_949);
and U2567 (N_2567,N_376,N_517);
nor U2568 (N_2568,N_875,N_139);
nand U2569 (N_2569,N_1272,N_818);
and U2570 (N_2570,N_932,N_1387);
nor U2571 (N_2571,N_1380,N_983);
xnor U2572 (N_2572,N_26,N_903);
nor U2573 (N_2573,N_437,N_1095);
or U2574 (N_2574,N_91,N_719);
or U2575 (N_2575,N_1048,N_588);
xnor U2576 (N_2576,N_35,N_196);
nand U2577 (N_2577,N_1258,N_816);
nor U2578 (N_2578,N_880,N_522);
nor U2579 (N_2579,N_917,N_139);
and U2580 (N_2580,N_291,N_702);
and U2581 (N_2581,N_695,N_952);
and U2582 (N_2582,N_340,N_1055);
nand U2583 (N_2583,N_169,N_1447);
or U2584 (N_2584,N_1405,N_1327);
nor U2585 (N_2585,N_205,N_780);
nand U2586 (N_2586,N_1041,N_1476);
and U2587 (N_2587,N_640,N_974);
and U2588 (N_2588,N_217,N_1042);
nor U2589 (N_2589,N_572,N_521);
xor U2590 (N_2590,N_95,N_1170);
nand U2591 (N_2591,N_846,N_1167);
nor U2592 (N_2592,N_230,N_270);
nor U2593 (N_2593,N_1092,N_14);
nor U2594 (N_2594,N_763,N_293);
or U2595 (N_2595,N_1108,N_1174);
or U2596 (N_2596,N_229,N_709);
and U2597 (N_2597,N_1429,N_810);
nand U2598 (N_2598,N_37,N_212);
or U2599 (N_2599,N_1373,N_1448);
nor U2600 (N_2600,N_417,N_791);
nand U2601 (N_2601,N_982,N_1341);
nand U2602 (N_2602,N_1256,N_986);
xnor U2603 (N_2603,N_772,N_1169);
or U2604 (N_2604,N_955,N_495);
or U2605 (N_2605,N_414,N_963);
or U2606 (N_2606,N_915,N_315);
nand U2607 (N_2607,N_1428,N_590);
xnor U2608 (N_2608,N_1328,N_996);
nand U2609 (N_2609,N_435,N_877);
nor U2610 (N_2610,N_1079,N_1107);
nand U2611 (N_2611,N_96,N_1402);
and U2612 (N_2612,N_670,N_1479);
and U2613 (N_2613,N_587,N_292);
or U2614 (N_2614,N_986,N_1025);
nand U2615 (N_2615,N_98,N_124);
or U2616 (N_2616,N_1135,N_123);
nor U2617 (N_2617,N_1088,N_282);
or U2618 (N_2618,N_1210,N_641);
xor U2619 (N_2619,N_1048,N_646);
or U2620 (N_2620,N_1393,N_1042);
or U2621 (N_2621,N_296,N_477);
or U2622 (N_2622,N_538,N_1434);
and U2623 (N_2623,N_446,N_1331);
or U2624 (N_2624,N_31,N_715);
xnor U2625 (N_2625,N_905,N_1387);
nand U2626 (N_2626,N_446,N_819);
nand U2627 (N_2627,N_421,N_51);
nor U2628 (N_2628,N_1189,N_945);
nand U2629 (N_2629,N_201,N_212);
and U2630 (N_2630,N_152,N_869);
nand U2631 (N_2631,N_1443,N_759);
or U2632 (N_2632,N_992,N_317);
or U2633 (N_2633,N_659,N_1388);
xor U2634 (N_2634,N_632,N_1475);
xor U2635 (N_2635,N_487,N_701);
xnor U2636 (N_2636,N_1167,N_1443);
xor U2637 (N_2637,N_242,N_1365);
and U2638 (N_2638,N_1006,N_712);
nand U2639 (N_2639,N_256,N_629);
and U2640 (N_2640,N_367,N_882);
nor U2641 (N_2641,N_736,N_1491);
and U2642 (N_2642,N_996,N_215);
nand U2643 (N_2643,N_1418,N_651);
and U2644 (N_2644,N_148,N_1090);
nand U2645 (N_2645,N_532,N_1386);
nor U2646 (N_2646,N_1139,N_630);
or U2647 (N_2647,N_787,N_1221);
xor U2648 (N_2648,N_53,N_938);
or U2649 (N_2649,N_195,N_12);
xnor U2650 (N_2650,N_759,N_182);
nand U2651 (N_2651,N_213,N_936);
or U2652 (N_2652,N_933,N_986);
or U2653 (N_2653,N_1028,N_981);
and U2654 (N_2654,N_289,N_1238);
and U2655 (N_2655,N_330,N_329);
and U2656 (N_2656,N_184,N_1355);
and U2657 (N_2657,N_1148,N_744);
nand U2658 (N_2658,N_863,N_553);
nor U2659 (N_2659,N_1491,N_69);
and U2660 (N_2660,N_409,N_527);
nand U2661 (N_2661,N_132,N_1455);
nor U2662 (N_2662,N_334,N_199);
nor U2663 (N_2663,N_214,N_56);
or U2664 (N_2664,N_67,N_1019);
nor U2665 (N_2665,N_115,N_1281);
nand U2666 (N_2666,N_366,N_665);
xor U2667 (N_2667,N_685,N_1042);
or U2668 (N_2668,N_287,N_1064);
nor U2669 (N_2669,N_1329,N_714);
or U2670 (N_2670,N_359,N_194);
nand U2671 (N_2671,N_738,N_133);
nor U2672 (N_2672,N_471,N_342);
nor U2673 (N_2673,N_83,N_158);
and U2674 (N_2674,N_538,N_198);
and U2675 (N_2675,N_1404,N_554);
or U2676 (N_2676,N_315,N_1429);
and U2677 (N_2677,N_931,N_586);
and U2678 (N_2678,N_855,N_978);
nand U2679 (N_2679,N_951,N_27);
and U2680 (N_2680,N_524,N_1013);
nand U2681 (N_2681,N_750,N_455);
xor U2682 (N_2682,N_174,N_1250);
or U2683 (N_2683,N_520,N_1317);
nand U2684 (N_2684,N_1069,N_1255);
xnor U2685 (N_2685,N_1483,N_71);
or U2686 (N_2686,N_804,N_1191);
or U2687 (N_2687,N_160,N_1317);
xor U2688 (N_2688,N_836,N_782);
and U2689 (N_2689,N_1101,N_148);
nor U2690 (N_2690,N_1307,N_107);
nand U2691 (N_2691,N_1065,N_215);
and U2692 (N_2692,N_1357,N_705);
nand U2693 (N_2693,N_320,N_1323);
and U2694 (N_2694,N_966,N_977);
xor U2695 (N_2695,N_272,N_406);
and U2696 (N_2696,N_1350,N_1343);
or U2697 (N_2697,N_1392,N_31);
nand U2698 (N_2698,N_639,N_758);
nor U2699 (N_2699,N_606,N_1494);
or U2700 (N_2700,N_1325,N_245);
and U2701 (N_2701,N_123,N_623);
nand U2702 (N_2702,N_1200,N_554);
xor U2703 (N_2703,N_164,N_635);
and U2704 (N_2704,N_839,N_516);
xor U2705 (N_2705,N_747,N_359);
nand U2706 (N_2706,N_1364,N_1287);
or U2707 (N_2707,N_1113,N_976);
or U2708 (N_2708,N_118,N_709);
and U2709 (N_2709,N_241,N_483);
xnor U2710 (N_2710,N_54,N_1353);
xor U2711 (N_2711,N_104,N_771);
xor U2712 (N_2712,N_219,N_1264);
nor U2713 (N_2713,N_485,N_156);
nor U2714 (N_2714,N_284,N_12);
nand U2715 (N_2715,N_920,N_254);
nand U2716 (N_2716,N_693,N_18);
xor U2717 (N_2717,N_1221,N_139);
nor U2718 (N_2718,N_90,N_1284);
and U2719 (N_2719,N_345,N_246);
nor U2720 (N_2720,N_28,N_1254);
nor U2721 (N_2721,N_1372,N_709);
nand U2722 (N_2722,N_758,N_1457);
nand U2723 (N_2723,N_1179,N_1198);
xnor U2724 (N_2724,N_832,N_1461);
or U2725 (N_2725,N_1282,N_1172);
and U2726 (N_2726,N_63,N_546);
nand U2727 (N_2727,N_834,N_417);
and U2728 (N_2728,N_386,N_1257);
nor U2729 (N_2729,N_147,N_192);
or U2730 (N_2730,N_553,N_1480);
and U2731 (N_2731,N_540,N_991);
nand U2732 (N_2732,N_1357,N_1367);
xnor U2733 (N_2733,N_545,N_1247);
or U2734 (N_2734,N_768,N_1090);
or U2735 (N_2735,N_1310,N_868);
and U2736 (N_2736,N_705,N_262);
nand U2737 (N_2737,N_169,N_830);
nand U2738 (N_2738,N_1488,N_132);
xor U2739 (N_2739,N_1006,N_1080);
or U2740 (N_2740,N_1300,N_458);
and U2741 (N_2741,N_37,N_793);
nand U2742 (N_2742,N_539,N_1453);
nand U2743 (N_2743,N_108,N_211);
nor U2744 (N_2744,N_712,N_173);
or U2745 (N_2745,N_954,N_1395);
and U2746 (N_2746,N_283,N_1275);
nor U2747 (N_2747,N_23,N_92);
or U2748 (N_2748,N_1014,N_1016);
nand U2749 (N_2749,N_194,N_833);
or U2750 (N_2750,N_1206,N_387);
nand U2751 (N_2751,N_102,N_462);
nor U2752 (N_2752,N_714,N_1390);
nor U2753 (N_2753,N_337,N_500);
and U2754 (N_2754,N_130,N_768);
nand U2755 (N_2755,N_273,N_485);
xnor U2756 (N_2756,N_253,N_220);
xor U2757 (N_2757,N_636,N_385);
xnor U2758 (N_2758,N_662,N_830);
or U2759 (N_2759,N_824,N_561);
nand U2760 (N_2760,N_1318,N_508);
nor U2761 (N_2761,N_410,N_75);
and U2762 (N_2762,N_106,N_457);
or U2763 (N_2763,N_111,N_327);
nand U2764 (N_2764,N_554,N_1383);
nand U2765 (N_2765,N_1161,N_1084);
xnor U2766 (N_2766,N_273,N_756);
nor U2767 (N_2767,N_1195,N_358);
and U2768 (N_2768,N_621,N_114);
or U2769 (N_2769,N_967,N_255);
nor U2770 (N_2770,N_1116,N_133);
xnor U2771 (N_2771,N_1319,N_507);
or U2772 (N_2772,N_1072,N_1275);
nor U2773 (N_2773,N_557,N_464);
or U2774 (N_2774,N_1142,N_824);
xor U2775 (N_2775,N_1043,N_1125);
and U2776 (N_2776,N_249,N_179);
and U2777 (N_2777,N_1288,N_1140);
nand U2778 (N_2778,N_1070,N_539);
nand U2779 (N_2779,N_68,N_1425);
xnor U2780 (N_2780,N_171,N_658);
nand U2781 (N_2781,N_1285,N_1439);
nand U2782 (N_2782,N_1086,N_334);
or U2783 (N_2783,N_78,N_162);
nor U2784 (N_2784,N_579,N_433);
xnor U2785 (N_2785,N_550,N_913);
xor U2786 (N_2786,N_305,N_533);
or U2787 (N_2787,N_1486,N_255);
nand U2788 (N_2788,N_651,N_190);
nand U2789 (N_2789,N_731,N_883);
nor U2790 (N_2790,N_236,N_239);
xor U2791 (N_2791,N_1248,N_735);
xnor U2792 (N_2792,N_697,N_820);
and U2793 (N_2793,N_893,N_1010);
or U2794 (N_2794,N_1430,N_963);
nor U2795 (N_2795,N_460,N_972);
nor U2796 (N_2796,N_1040,N_1072);
and U2797 (N_2797,N_1359,N_365);
and U2798 (N_2798,N_909,N_841);
nor U2799 (N_2799,N_1391,N_1316);
xnor U2800 (N_2800,N_732,N_1417);
nand U2801 (N_2801,N_841,N_713);
nor U2802 (N_2802,N_689,N_698);
xnor U2803 (N_2803,N_970,N_991);
and U2804 (N_2804,N_171,N_374);
nand U2805 (N_2805,N_1105,N_396);
xnor U2806 (N_2806,N_1289,N_508);
nor U2807 (N_2807,N_654,N_68);
and U2808 (N_2808,N_1072,N_664);
xor U2809 (N_2809,N_1314,N_826);
xnor U2810 (N_2810,N_202,N_75);
nor U2811 (N_2811,N_462,N_1177);
nand U2812 (N_2812,N_1276,N_136);
nand U2813 (N_2813,N_1083,N_899);
and U2814 (N_2814,N_886,N_1324);
nor U2815 (N_2815,N_247,N_501);
or U2816 (N_2816,N_388,N_1331);
or U2817 (N_2817,N_638,N_212);
or U2818 (N_2818,N_1410,N_635);
xor U2819 (N_2819,N_22,N_652);
nand U2820 (N_2820,N_1008,N_491);
nand U2821 (N_2821,N_1311,N_822);
and U2822 (N_2822,N_1164,N_708);
or U2823 (N_2823,N_433,N_1472);
or U2824 (N_2824,N_957,N_868);
and U2825 (N_2825,N_1112,N_89);
nand U2826 (N_2826,N_942,N_358);
or U2827 (N_2827,N_1286,N_1131);
or U2828 (N_2828,N_354,N_148);
nor U2829 (N_2829,N_1362,N_493);
xor U2830 (N_2830,N_764,N_180);
xor U2831 (N_2831,N_50,N_840);
nand U2832 (N_2832,N_252,N_1128);
and U2833 (N_2833,N_767,N_951);
nor U2834 (N_2834,N_535,N_814);
or U2835 (N_2835,N_1309,N_1407);
nor U2836 (N_2836,N_1038,N_1113);
nand U2837 (N_2837,N_116,N_259);
xnor U2838 (N_2838,N_429,N_74);
and U2839 (N_2839,N_39,N_1314);
xnor U2840 (N_2840,N_648,N_1354);
xor U2841 (N_2841,N_110,N_291);
and U2842 (N_2842,N_1319,N_1290);
nand U2843 (N_2843,N_1115,N_1226);
xnor U2844 (N_2844,N_201,N_1434);
xnor U2845 (N_2845,N_165,N_1258);
nor U2846 (N_2846,N_1041,N_409);
or U2847 (N_2847,N_121,N_855);
or U2848 (N_2848,N_1415,N_392);
nor U2849 (N_2849,N_1142,N_553);
xor U2850 (N_2850,N_1454,N_581);
nand U2851 (N_2851,N_147,N_340);
nand U2852 (N_2852,N_887,N_1462);
nor U2853 (N_2853,N_146,N_6);
or U2854 (N_2854,N_271,N_659);
xnor U2855 (N_2855,N_590,N_169);
nand U2856 (N_2856,N_1487,N_123);
or U2857 (N_2857,N_844,N_139);
or U2858 (N_2858,N_860,N_302);
xnor U2859 (N_2859,N_37,N_1244);
and U2860 (N_2860,N_421,N_946);
or U2861 (N_2861,N_390,N_683);
xnor U2862 (N_2862,N_915,N_1370);
xor U2863 (N_2863,N_1108,N_732);
nor U2864 (N_2864,N_1142,N_653);
nand U2865 (N_2865,N_121,N_1434);
and U2866 (N_2866,N_118,N_1329);
or U2867 (N_2867,N_42,N_591);
xor U2868 (N_2868,N_756,N_325);
nand U2869 (N_2869,N_441,N_448);
or U2870 (N_2870,N_1213,N_1482);
and U2871 (N_2871,N_1499,N_1455);
and U2872 (N_2872,N_1329,N_1160);
nor U2873 (N_2873,N_742,N_932);
xnor U2874 (N_2874,N_1476,N_988);
nand U2875 (N_2875,N_1037,N_590);
and U2876 (N_2876,N_1312,N_938);
xnor U2877 (N_2877,N_1404,N_490);
xor U2878 (N_2878,N_775,N_624);
nor U2879 (N_2879,N_993,N_1081);
nor U2880 (N_2880,N_1155,N_1495);
xnor U2881 (N_2881,N_1454,N_856);
nor U2882 (N_2882,N_858,N_1070);
nand U2883 (N_2883,N_1133,N_168);
or U2884 (N_2884,N_30,N_288);
nor U2885 (N_2885,N_1189,N_1496);
xnor U2886 (N_2886,N_318,N_1116);
or U2887 (N_2887,N_602,N_416);
xor U2888 (N_2888,N_369,N_313);
and U2889 (N_2889,N_897,N_70);
nand U2890 (N_2890,N_1365,N_413);
xor U2891 (N_2891,N_194,N_355);
xor U2892 (N_2892,N_1348,N_569);
xor U2893 (N_2893,N_259,N_506);
or U2894 (N_2894,N_879,N_488);
nor U2895 (N_2895,N_636,N_1047);
xnor U2896 (N_2896,N_1323,N_1491);
and U2897 (N_2897,N_255,N_1106);
xor U2898 (N_2898,N_707,N_1447);
or U2899 (N_2899,N_1018,N_1161);
or U2900 (N_2900,N_217,N_82);
or U2901 (N_2901,N_1151,N_631);
nand U2902 (N_2902,N_1493,N_1366);
and U2903 (N_2903,N_1070,N_1458);
nand U2904 (N_2904,N_1319,N_341);
xnor U2905 (N_2905,N_431,N_782);
and U2906 (N_2906,N_1383,N_882);
and U2907 (N_2907,N_692,N_809);
xor U2908 (N_2908,N_1142,N_1016);
nor U2909 (N_2909,N_97,N_491);
nor U2910 (N_2910,N_1162,N_1033);
and U2911 (N_2911,N_223,N_902);
nor U2912 (N_2912,N_488,N_53);
and U2913 (N_2913,N_1339,N_582);
nor U2914 (N_2914,N_1437,N_1384);
xnor U2915 (N_2915,N_51,N_1165);
or U2916 (N_2916,N_1238,N_933);
nand U2917 (N_2917,N_793,N_384);
and U2918 (N_2918,N_1064,N_799);
nor U2919 (N_2919,N_1339,N_1328);
nand U2920 (N_2920,N_497,N_78);
or U2921 (N_2921,N_1455,N_20);
nand U2922 (N_2922,N_1133,N_1349);
and U2923 (N_2923,N_569,N_1144);
nand U2924 (N_2924,N_231,N_750);
nor U2925 (N_2925,N_1388,N_710);
and U2926 (N_2926,N_1491,N_2);
nand U2927 (N_2927,N_149,N_561);
xor U2928 (N_2928,N_152,N_1410);
xnor U2929 (N_2929,N_334,N_898);
xnor U2930 (N_2930,N_686,N_790);
nor U2931 (N_2931,N_67,N_1024);
nand U2932 (N_2932,N_949,N_906);
nor U2933 (N_2933,N_151,N_393);
xor U2934 (N_2934,N_1146,N_396);
xnor U2935 (N_2935,N_1122,N_1275);
nand U2936 (N_2936,N_333,N_190);
and U2937 (N_2937,N_56,N_791);
or U2938 (N_2938,N_68,N_300);
or U2939 (N_2939,N_1413,N_1223);
or U2940 (N_2940,N_680,N_144);
nand U2941 (N_2941,N_122,N_1365);
or U2942 (N_2942,N_657,N_471);
or U2943 (N_2943,N_1438,N_1321);
nand U2944 (N_2944,N_457,N_1085);
xnor U2945 (N_2945,N_174,N_141);
nor U2946 (N_2946,N_801,N_1026);
nand U2947 (N_2947,N_1484,N_373);
nor U2948 (N_2948,N_1170,N_851);
nand U2949 (N_2949,N_1131,N_156);
nor U2950 (N_2950,N_1313,N_1454);
or U2951 (N_2951,N_850,N_403);
and U2952 (N_2952,N_851,N_650);
nor U2953 (N_2953,N_652,N_1298);
or U2954 (N_2954,N_403,N_807);
and U2955 (N_2955,N_1422,N_762);
or U2956 (N_2956,N_1124,N_1071);
xnor U2957 (N_2957,N_165,N_1289);
and U2958 (N_2958,N_1197,N_606);
nand U2959 (N_2959,N_354,N_48);
nand U2960 (N_2960,N_693,N_957);
nor U2961 (N_2961,N_1395,N_128);
nand U2962 (N_2962,N_594,N_786);
nor U2963 (N_2963,N_1245,N_45);
nand U2964 (N_2964,N_758,N_1091);
nand U2965 (N_2965,N_1497,N_1412);
nand U2966 (N_2966,N_689,N_987);
nand U2967 (N_2967,N_1402,N_65);
nor U2968 (N_2968,N_167,N_592);
nor U2969 (N_2969,N_229,N_1403);
or U2970 (N_2970,N_221,N_1481);
and U2971 (N_2971,N_647,N_763);
xor U2972 (N_2972,N_624,N_424);
and U2973 (N_2973,N_231,N_1141);
or U2974 (N_2974,N_704,N_394);
nand U2975 (N_2975,N_687,N_1051);
or U2976 (N_2976,N_466,N_1388);
or U2977 (N_2977,N_600,N_1328);
and U2978 (N_2978,N_830,N_1130);
xor U2979 (N_2979,N_428,N_335);
and U2980 (N_2980,N_1052,N_935);
and U2981 (N_2981,N_717,N_305);
xnor U2982 (N_2982,N_366,N_809);
xnor U2983 (N_2983,N_1290,N_95);
nor U2984 (N_2984,N_1363,N_557);
and U2985 (N_2985,N_1266,N_841);
nand U2986 (N_2986,N_634,N_278);
and U2987 (N_2987,N_220,N_693);
nor U2988 (N_2988,N_863,N_1146);
nor U2989 (N_2989,N_599,N_68);
nor U2990 (N_2990,N_279,N_950);
or U2991 (N_2991,N_355,N_819);
nor U2992 (N_2992,N_1055,N_504);
or U2993 (N_2993,N_293,N_983);
nand U2994 (N_2994,N_831,N_644);
nand U2995 (N_2995,N_506,N_1274);
or U2996 (N_2996,N_606,N_1365);
and U2997 (N_2997,N_1432,N_1101);
and U2998 (N_2998,N_73,N_791);
nand U2999 (N_2999,N_913,N_328);
nand U3000 (N_3000,N_2845,N_2837);
nand U3001 (N_3001,N_1832,N_1900);
or U3002 (N_3002,N_2194,N_2528);
and U3003 (N_3003,N_1674,N_2412);
or U3004 (N_3004,N_2140,N_2147);
xnor U3005 (N_3005,N_1979,N_2497);
nor U3006 (N_3006,N_1861,N_1935);
and U3007 (N_3007,N_2509,N_2268);
or U3008 (N_3008,N_2264,N_2239);
and U3009 (N_3009,N_1856,N_1599);
and U3010 (N_3010,N_2296,N_1573);
or U3011 (N_3011,N_1623,N_2563);
and U3012 (N_3012,N_1793,N_2463);
or U3013 (N_3013,N_2173,N_2215);
and U3014 (N_3014,N_1764,N_2907);
nor U3015 (N_3015,N_2921,N_1989);
nor U3016 (N_3016,N_1513,N_1788);
nor U3017 (N_3017,N_2090,N_2277);
xor U3018 (N_3018,N_2698,N_1562);
and U3019 (N_3019,N_2311,N_2930);
xor U3020 (N_3020,N_1571,N_1695);
nand U3021 (N_3021,N_2891,N_2785);
nor U3022 (N_3022,N_1522,N_1626);
and U3023 (N_3023,N_1679,N_2163);
nor U3024 (N_3024,N_1719,N_1576);
nor U3025 (N_3025,N_2975,N_2417);
or U3026 (N_3026,N_1745,N_1633);
xor U3027 (N_3027,N_2680,N_1639);
nand U3028 (N_3028,N_2848,N_1858);
or U3029 (N_3029,N_1780,N_1532);
and U3030 (N_3030,N_2692,N_2263);
and U3031 (N_3031,N_2396,N_2386);
or U3032 (N_3032,N_1803,N_2787);
and U3033 (N_3033,N_2513,N_2797);
nor U3034 (N_3034,N_2148,N_2336);
or U3035 (N_3035,N_2130,N_1661);
and U3036 (N_3036,N_2211,N_1903);
and U3037 (N_3037,N_1826,N_2355);
nor U3038 (N_3038,N_2932,N_2131);
nor U3039 (N_3039,N_2568,N_2841);
nor U3040 (N_3040,N_1967,N_2626);
nor U3041 (N_3041,N_1866,N_2811);
nor U3042 (N_3042,N_2636,N_2260);
and U3043 (N_3043,N_2561,N_2892);
xor U3044 (N_3044,N_2885,N_1564);
nand U3045 (N_3045,N_1638,N_1931);
or U3046 (N_3046,N_2049,N_1756);
nor U3047 (N_3047,N_1889,N_1666);
or U3048 (N_3048,N_2609,N_1586);
nor U3049 (N_3049,N_2861,N_1662);
and U3050 (N_3050,N_2805,N_2216);
xor U3051 (N_3051,N_2204,N_1555);
and U3052 (N_3052,N_2040,N_2987);
xnor U3053 (N_3053,N_2661,N_2723);
nand U3054 (N_3054,N_1942,N_1747);
xor U3055 (N_3055,N_1624,N_2525);
xor U3056 (N_3056,N_2757,N_1902);
nor U3057 (N_3057,N_2519,N_1701);
and U3058 (N_3058,N_2257,N_2766);
or U3059 (N_3059,N_2222,N_2562);
and U3060 (N_3060,N_1766,N_2832);
and U3061 (N_3061,N_2390,N_2421);
or U3062 (N_3062,N_2593,N_1930);
xnor U3063 (N_3063,N_1683,N_2056);
or U3064 (N_3064,N_2315,N_2476);
or U3065 (N_3065,N_2653,N_2182);
nor U3066 (N_3066,N_2498,N_2080);
or U3067 (N_3067,N_2247,N_1687);
or U3068 (N_3068,N_2475,N_2142);
or U3069 (N_3069,N_2784,N_2874);
nor U3070 (N_3070,N_1534,N_1837);
xor U3071 (N_3071,N_2026,N_1936);
or U3072 (N_3072,N_2377,N_1539);
and U3073 (N_3073,N_1946,N_1632);
nand U3074 (N_3074,N_2295,N_2686);
and U3075 (N_3075,N_2384,N_1763);
nand U3076 (N_3076,N_2279,N_1897);
xor U3077 (N_3077,N_2155,N_2484);
or U3078 (N_3078,N_1878,N_1822);
nand U3079 (N_3079,N_1870,N_1817);
and U3080 (N_3080,N_2812,N_2774);
and U3081 (N_3081,N_1727,N_2962);
xnor U3082 (N_3082,N_2794,N_1579);
nand U3083 (N_3083,N_2743,N_2491);
xor U3084 (N_3084,N_2226,N_2411);
or U3085 (N_3085,N_1997,N_2245);
nand U3086 (N_3086,N_2214,N_1651);
xnor U3087 (N_3087,N_2183,N_1899);
nand U3088 (N_3088,N_2150,N_2188);
or U3089 (N_3089,N_1739,N_2307);
xnor U3090 (N_3090,N_1986,N_2083);
and U3091 (N_3091,N_2343,N_2869);
and U3092 (N_3092,N_2993,N_1561);
nor U3093 (N_3093,N_2842,N_1804);
xor U3094 (N_3094,N_2508,N_1892);
nand U3095 (N_3095,N_2919,N_1553);
xnor U3096 (N_3096,N_2552,N_2868);
or U3097 (N_3097,N_1637,N_2485);
xor U3098 (N_3098,N_2046,N_2015);
xnor U3099 (N_3099,N_2413,N_2172);
nand U3100 (N_3100,N_1885,N_2925);
nand U3101 (N_3101,N_2543,N_2435);
and U3102 (N_3102,N_2077,N_1653);
and U3103 (N_3103,N_2756,N_2791);
xnor U3104 (N_3104,N_1733,N_2021);
and U3105 (N_3105,N_2713,N_2574);
or U3106 (N_3106,N_1536,N_1521);
and U3107 (N_3107,N_1867,N_1775);
nor U3108 (N_3108,N_2715,N_2909);
nor U3109 (N_3109,N_2641,N_1830);
nand U3110 (N_3110,N_2321,N_1730);
or U3111 (N_3111,N_2658,N_1659);
or U3112 (N_3112,N_2361,N_2855);
xnor U3113 (N_3113,N_2720,N_1808);
xnor U3114 (N_3114,N_1709,N_1590);
nand U3115 (N_3115,N_1919,N_1574);
or U3116 (N_3116,N_1517,N_2379);
nand U3117 (N_3117,N_1992,N_1966);
or U3118 (N_3118,N_1791,N_2983);
nor U3119 (N_3119,N_2044,N_1958);
nor U3120 (N_3120,N_2350,N_2726);
nand U3121 (N_3121,N_1834,N_2125);
xor U3122 (N_3122,N_1568,N_2996);
nand U3123 (N_3123,N_1960,N_1589);
nand U3124 (N_3124,N_2977,N_1615);
nor U3125 (N_3125,N_2195,N_2870);
nand U3126 (N_3126,N_2029,N_2093);
or U3127 (N_3127,N_2106,N_1577);
and U3128 (N_3128,N_2821,N_2037);
nand U3129 (N_3129,N_2569,N_1542);
nor U3130 (N_3130,N_1849,N_2980);
nand U3131 (N_3131,N_1508,N_2445);
or U3132 (N_3132,N_1620,N_2269);
or U3133 (N_3133,N_2433,N_2351);
nand U3134 (N_3134,N_1732,N_2630);
and U3135 (N_3135,N_2309,N_1748);
nor U3136 (N_3136,N_1660,N_2053);
xor U3137 (N_3137,N_1757,N_1514);
nor U3138 (N_3138,N_2085,N_2619);
nand U3139 (N_3139,N_2341,N_2542);
nand U3140 (N_3140,N_2141,N_2603);
xnor U3141 (N_3141,N_1749,N_2023);
or U3142 (N_3142,N_2673,N_2978);
and U3143 (N_3143,N_1614,N_1667);
and U3144 (N_3144,N_2681,N_2843);
nand U3145 (N_3145,N_2804,N_2225);
nand U3146 (N_3146,N_1621,N_2059);
and U3147 (N_3147,N_1565,N_2376);
nor U3148 (N_3148,N_1921,N_2096);
nand U3149 (N_3149,N_2894,N_2139);
and U3150 (N_3150,N_2359,N_1920);
or U3151 (N_3151,N_2221,N_2536);
or U3152 (N_3152,N_2920,N_2004);
xor U3153 (N_3153,N_2110,N_1669);
and U3154 (N_3154,N_2319,N_1691);
xnor U3155 (N_3155,N_1898,N_2905);
nor U3156 (N_3156,N_2814,N_1781);
nand U3157 (N_3157,N_2937,N_2378);
nand U3158 (N_3158,N_2911,N_2382);
and U3159 (N_3159,N_2599,N_2432);
or U3160 (N_3160,N_1972,N_2762);
and U3161 (N_3161,N_2388,N_1779);
and U3162 (N_3162,N_2428,N_2352);
and U3163 (N_3163,N_1926,N_2072);
xor U3164 (N_3164,N_1864,N_1641);
nor U3165 (N_3165,N_1770,N_1915);
xnor U3166 (N_3166,N_2954,N_2707);
xor U3167 (N_3167,N_1906,N_1887);
xnor U3168 (N_3168,N_2606,N_2864);
nor U3169 (N_3169,N_1708,N_2455);
or U3170 (N_3170,N_1742,N_1863);
nand U3171 (N_3171,N_2544,N_2403);
nand U3172 (N_3172,N_2638,N_2880);
or U3173 (N_3173,N_1681,N_1509);
and U3174 (N_3174,N_2482,N_2088);
nor U3175 (N_3175,N_2637,N_2575);
nand U3176 (N_3176,N_2285,N_2700);
and U3177 (N_3177,N_1760,N_2738);
xnor U3178 (N_3178,N_1957,N_1604);
and U3179 (N_3179,N_2986,N_2387);
xnor U3180 (N_3180,N_2200,N_2464);
xnor U3181 (N_3181,N_1968,N_2668);
or U3182 (N_3182,N_1649,N_2231);
and U3183 (N_3183,N_1777,N_2219);
nand U3184 (N_3184,N_2136,N_2358);
and U3185 (N_3185,N_1981,N_1538);
nor U3186 (N_3186,N_2557,N_2976);
or U3187 (N_3187,N_2076,N_2527);
or U3188 (N_3188,N_2656,N_2878);
and U3189 (N_3189,N_2457,N_2236);
or U3190 (N_3190,N_1888,N_2852);
and U3191 (N_3191,N_2752,N_2601);
nor U3192 (N_3192,N_1635,N_2313);
or U3193 (N_3193,N_2181,N_2960);
nor U3194 (N_3194,N_2753,N_2748);
or U3195 (N_3195,N_2467,N_2763);
nor U3196 (N_3196,N_1618,N_2663);
and U3197 (N_3197,N_1506,N_2929);
nor U3198 (N_3198,N_1663,N_2158);
nand U3199 (N_3199,N_2454,N_1551);
or U3200 (N_3200,N_1596,N_2511);
nand U3201 (N_3201,N_2688,N_1904);
and U3202 (N_3202,N_1790,N_1569);
and U3203 (N_3203,N_2685,N_2531);
nor U3204 (N_3204,N_2833,N_2157);
or U3205 (N_3205,N_2281,N_2906);
and U3206 (N_3206,N_1833,N_2910);
or U3207 (N_3207,N_2572,N_1873);
or U3208 (N_3208,N_2324,N_1690);
and U3209 (N_3209,N_1907,N_2126);
nor U3210 (N_3210,N_2375,N_1726);
and U3211 (N_3211,N_2866,N_2846);
and U3212 (N_3212,N_1927,N_2128);
or U3213 (N_3213,N_2782,N_2209);
xnor U3214 (N_3214,N_2771,N_1504);
nor U3215 (N_3215,N_1598,N_2108);
xor U3216 (N_3216,N_2600,N_1840);
or U3217 (N_3217,N_2566,N_2516);
nor U3218 (N_3218,N_2939,N_2585);
xor U3219 (N_3219,N_1525,N_2770);
and U3220 (N_3220,N_2144,N_2614);
xnor U3221 (N_3221,N_2474,N_2967);
nand U3222 (N_3222,N_1540,N_2876);
nor U3223 (N_3223,N_2777,N_2233);
or U3224 (N_3224,N_2442,N_2789);
nand U3225 (N_3225,N_2399,N_1723);
or U3226 (N_3226,N_1950,N_1563);
nor U3227 (N_3227,N_2969,N_2137);
xor U3228 (N_3228,N_2329,N_2075);
and U3229 (N_3229,N_2063,N_1990);
nor U3230 (N_3230,N_1601,N_2208);
nand U3231 (N_3231,N_2571,N_2573);
nand U3232 (N_3232,N_1941,N_1850);
and U3233 (N_3233,N_2510,N_2089);
nor U3234 (N_3234,N_2768,N_1627);
or U3235 (N_3235,N_2299,N_2617);
nor U3236 (N_3236,N_1984,N_2325);
or U3237 (N_3237,N_2642,N_2441);
or U3238 (N_3238,N_2270,N_2167);
nand U3239 (N_3239,N_2953,N_2010);
xor U3240 (N_3240,N_2320,N_2345);
or U3241 (N_3241,N_1758,N_2813);
xor U3242 (N_3242,N_1807,N_1933);
and U3243 (N_3243,N_1824,N_1693);
and U3244 (N_3244,N_2154,N_2731);
and U3245 (N_3245,N_1751,N_1880);
xnor U3246 (N_3246,N_1597,N_2312);
and U3247 (N_3247,N_2631,N_2248);
and U3248 (N_3248,N_1500,N_2549);
nand U3249 (N_3249,N_1510,N_1603);
xnor U3250 (N_3250,N_2280,N_1595);
xor U3251 (N_3251,N_2853,N_2815);
and U3252 (N_3252,N_1705,N_2149);
nor U3253 (N_3253,N_2207,N_2452);
and U3254 (N_3254,N_2469,N_2372);
and U3255 (N_3255,N_1810,N_2898);
and U3256 (N_3256,N_2045,N_2220);
nor U3257 (N_3257,N_2005,N_2458);
nor U3258 (N_3258,N_2169,N_1698);
nor U3259 (N_3259,N_1677,N_1657);
xor U3260 (N_3260,N_2471,N_2778);
nor U3261 (N_3261,N_2440,N_2449);
nor U3262 (N_3262,N_2702,N_2486);
or U3263 (N_3263,N_2335,N_2028);
xor U3264 (N_3264,N_2669,N_2696);
and U3265 (N_3265,N_2206,N_2301);
nand U3266 (N_3266,N_2618,N_1575);
and U3267 (N_3267,N_1797,N_2747);
xnor U3268 (N_3268,N_2775,N_2918);
or U3269 (N_3269,N_2646,N_1725);
nor U3270 (N_3270,N_2326,N_1721);
nand U3271 (N_3271,N_1668,N_1759);
nor U3272 (N_3272,N_1755,N_2662);
nand U3273 (N_3273,N_1865,N_2607);
nand U3274 (N_3274,N_2958,N_2951);
nand U3275 (N_3275,N_2589,N_1815);
nand U3276 (N_3276,N_2714,N_1648);
or U3277 (N_3277,N_2802,N_2480);
xnor U3278 (N_3278,N_2406,N_2462);
xor U3279 (N_3279,N_2941,N_2547);
and U3280 (N_3280,N_2587,N_1692);
nor U3281 (N_3281,N_2620,N_2114);
xnor U3282 (N_3282,N_2709,N_1868);
nor U3283 (N_3283,N_2119,N_1530);
nand U3284 (N_3284,N_2613,N_2357);
nand U3285 (N_3285,N_2256,N_2025);
and U3286 (N_3286,N_2177,N_1642);
nor U3287 (N_3287,N_2666,N_2538);
nor U3288 (N_3288,N_1531,N_1678);
and U3289 (N_3289,N_1718,N_1580);
or U3290 (N_3290,N_2780,N_1744);
nand U3291 (N_3291,N_1829,N_2875);
nor U3292 (N_3292,N_1993,N_2397);
and U3293 (N_3293,N_2253,N_2287);
nor U3294 (N_3294,N_1836,N_2303);
nand U3295 (N_3295,N_2900,N_1955);
or U3296 (N_3296,N_1855,N_2203);
nor U3297 (N_3297,N_2451,N_2481);
nand U3298 (N_3298,N_2009,N_2839);
nor U3299 (N_3299,N_1857,N_2973);
xnor U3300 (N_3300,N_1606,N_1910);
nor U3301 (N_3301,N_2316,N_1609);
nand U3302 (N_3302,N_2091,N_1913);
or U3303 (N_3303,N_2758,N_1636);
nor U3304 (N_3304,N_2156,N_1922);
nor U3305 (N_3305,N_2588,N_1932);
xnor U3306 (N_3306,N_2000,N_2460);
xnor U3307 (N_3307,N_2422,N_1511);
xor U3308 (N_3308,N_2665,N_2795);
and U3309 (N_3309,N_2470,N_2964);
nand U3310 (N_3310,N_2064,N_1812);
nor U3311 (N_3311,N_2302,N_2728);
nor U3312 (N_3312,N_2683,N_1588);
nor U3313 (N_3313,N_2830,N_2899);
xor U3314 (N_3314,N_2567,N_2152);
or U3315 (N_3315,N_2430,N_2927);
nand U3316 (N_3316,N_1684,N_1959);
or U3317 (N_3317,N_2250,N_1848);
xor U3318 (N_3318,N_2779,N_2252);
nor U3319 (N_3319,N_2041,N_2946);
nand U3320 (N_3320,N_2706,N_1631);
xnor U3321 (N_3321,N_2772,N_1784);
and U3322 (N_3322,N_2346,N_1617);
or U3323 (N_3323,N_2514,N_1852);
nor U3324 (N_3324,N_2734,N_1825);
and U3325 (N_3325,N_2087,N_2217);
or U3326 (N_3326,N_2385,N_1996);
and U3327 (N_3327,N_1835,N_2831);
xor U3328 (N_3328,N_2579,N_1792);
or U3329 (N_3329,N_1557,N_1844);
nor U3330 (N_3330,N_2006,N_2068);
nor U3331 (N_3331,N_2235,N_2998);
xnor U3332 (N_3332,N_2934,N_2404);
nand U3333 (N_3333,N_1696,N_2755);
and U3334 (N_3334,N_2115,N_2229);
nand U3335 (N_3335,N_1973,N_1610);
nand U3336 (N_3336,N_2950,N_2273);
and U3337 (N_3337,N_2013,N_2447);
nor U3338 (N_3338,N_2410,N_1533);
nand U3339 (N_3339,N_2165,N_2740);
or U3340 (N_3340,N_1643,N_1754);
nand U3341 (N_3341,N_1740,N_2232);
nand U3342 (N_3342,N_2807,N_2180);
and U3343 (N_3343,N_1847,N_2835);
xnor U3344 (N_3344,N_1991,N_1505);
nor U3345 (N_3345,N_2278,N_2790);
nor U3346 (N_3346,N_1673,N_1676);
xor U3347 (N_3347,N_2436,N_2674);
and U3348 (N_3348,N_2682,N_2366);
nor U3349 (N_3349,N_1975,N_2690);
and U3350 (N_3350,N_2213,N_1736);
nor U3351 (N_3351,N_1890,N_2550);
or U3352 (N_3352,N_2011,N_1543);
or U3353 (N_3353,N_2122,N_2548);
xor U3354 (N_3354,N_2847,N_1675);
or U3355 (N_3355,N_2365,N_1971);
nand U3356 (N_3356,N_2851,N_1717);
xnor U3357 (N_3357,N_2118,N_1944);
and U3358 (N_3358,N_2859,N_2796);
nand U3359 (N_3359,N_1896,N_2621);
nor U3360 (N_3360,N_2627,N_1951);
and U3361 (N_3361,N_2935,N_2305);
xor U3362 (N_3362,N_2761,N_2584);
nor U3363 (N_3363,N_1753,N_1916);
and U3364 (N_3364,N_2196,N_1943);
or U3365 (N_3365,N_2035,N_2995);
and U3366 (N_3366,N_1592,N_2506);
or U3367 (N_3367,N_2104,N_2423);
nor U3368 (N_3368,N_2730,N_2955);
or U3369 (N_3369,N_2988,N_1622);
nand U3370 (N_3370,N_2660,N_2529);
nor U3371 (N_3371,N_2494,N_2800);
and U3372 (N_3372,N_2776,N_2959);
nor U3373 (N_3373,N_2979,N_2395);
nor U3374 (N_3374,N_2348,N_2117);
and U3375 (N_3375,N_1702,N_2591);
nand U3376 (N_3376,N_2007,N_1908);
and U3377 (N_3377,N_2520,N_2697);
or U3378 (N_3378,N_1982,N_1948);
and U3379 (N_3379,N_2308,N_1771);
or U3380 (N_3380,N_1665,N_1528);
nor U3381 (N_3381,N_2556,N_1567);
xor U3382 (N_3382,N_2061,N_2888);
or U3383 (N_3383,N_2913,N_2582);
or U3384 (N_3384,N_2230,N_2570);
or U3385 (N_3385,N_2801,N_1854);
nor U3386 (N_3386,N_1816,N_1629);
xnor U3387 (N_3387,N_1560,N_2704);
xnor U3388 (N_3388,N_1529,N_1545);
nand U3389 (N_3389,N_1728,N_1554);
and U3390 (N_3390,N_2933,N_1895);
nor U3391 (N_3391,N_2294,N_2541);
and U3392 (N_3392,N_1987,N_2438);
nand U3393 (N_3393,N_1634,N_1947);
and U3394 (N_3394,N_1671,N_1819);
nor U3395 (N_3395,N_2717,N_2461);
nand U3396 (N_3396,N_2162,N_1827);
and U3397 (N_3397,N_2490,N_2971);
nand U3398 (N_3398,N_1512,N_1862);
nor U3399 (N_3399,N_1846,N_2291);
nand U3400 (N_3400,N_2625,N_1704);
nor U3401 (N_3401,N_2038,N_2071);
and U3402 (N_3402,N_1828,N_1587);
or U3403 (N_3403,N_2197,N_2394);
nand U3404 (N_3404,N_1535,N_2936);
nand U3405 (N_3405,N_2901,N_2459);
and U3406 (N_3406,N_2409,N_2065);
and U3407 (N_3407,N_2555,N_2810);
nor U3408 (N_3408,N_2465,N_2624);
xor U3409 (N_3409,N_2725,N_2949);
nand U3410 (N_3410,N_2434,N_2928);
and U3411 (N_3411,N_2699,N_1918);
and U3412 (N_3412,N_2254,N_2735);
or U3413 (N_3413,N_2691,N_1658);
xor U3414 (N_3414,N_2389,N_2545);
xnor U3415 (N_3415,N_2450,N_2178);
nand U3416 (N_3416,N_1547,N_2716);
nor U3417 (N_3417,N_2073,N_2676);
xor U3418 (N_3418,N_2840,N_2597);
nor U3419 (N_3419,N_2783,N_1762);
and U3420 (N_3420,N_2507,N_1516);
nor U3421 (N_3421,N_1934,N_2271);
nor U3422 (N_3422,N_2415,N_2292);
xor U3423 (N_3423,N_2737,N_2659);
and U3424 (N_3424,N_2654,N_1556);
nand U3425 (N_3425,N_2970,N_1891);
and U3426 (N_3426,N_1613,N_2478);
and U3427 (N_3427,N_2401,N_2289);
or U3428 (N_3428,N_2179,N_2168);
xor U3429 (N_3429,N_1507,N_2331);
xor U3430 (N_3430,N_2340,N_2185);
and U3431 (N_3431,N_2703,N_2337);
or U3432 (N_3432,N_2829,N_1976);
and U3433 (N_3433,N_2132,N_2749);
and U3434 (N_3434,N_1831,N_2966);
nand U3435 (N_3435,N_1884,N_1591);
nand U3436 (N_3436,N_2546,N_2218);
xnor U3437 (N_3437,N_2611,N_2535);
and U3438 (N_3438,N_2948,N_1746);
nand U3439 (N_3439,N_2184,N_2592);
xnor U3440 (N_3440,N_1672,N_2518);
and U3441 (N_3441,N_2327,N_2058);
nor U3442 (N_3442,N_2499,N_2741);
or U3443 (N_3443,N_1845,N_2825);
nor U3444 (N_3444,N_1616,N_2640);
or U3445 (N_3445,N_1795,N_2120);
and U3446 (N_3446,N_2223,N_2719);
or U3447 (N_3447,N_2773,N_2564);
or U3448 (N_3448,N_1820,N_2530);
or U3449 (N_3449,N_2754,N_1550);
xnor U3450 (N_3450,N_1761,N_2398);
and U3451 (N_3451,N_2596,N_1654);
nand U3452 (N_3452,N_1894,N_2055);
and U3453 (N_3453,N_2760,N_1785);
nor U3454 (N_3454,N_2989,N_2952);
or U3455 (N_3455,N_2405,N_2051);
or U3456 (N_3456,N_2836,N_2972);
nand U3457 (N_3457,N_2001,N_2739);
and U3458 (N_3458,N_1619,N_1954);
nor U3459 (N_3459,N_2266,N_2174);
nand U3460 (N_3460,N_2145,N_1809);
nand U3461 (N_3461,N_2082,N_2175);
xor U3462 (N_3462,N_2887,N_2342);
nor U3463 (N_3463,N_2241,N_1798);
xor U3464 (N_3464,N_1503,N_2062);
nor U3465 (N_3465,N_2135,N_2940);
and U3466 (N_3466,N_2402,N_1911);
nor U3467 (N_3467,N_1956,N_2227);
nor U3468 (N_3468,N_1743,N_2275);
nand U3469 (N_3469,N_2895,N_2590);
xor U3470 (N_3470,N_2306,N_2456);
xor U3471 (N_3471,N_1774,N_1682);
xor U3472 (N_3472,N_1706,N_2098);
and U3473 (N_3473,N_1901,N_2675);
or U3474 (N_3474,N_2027,N_2863);
and U3475 (N_3475,N_2304,N_2371);
xor U3476 (N_3476,N_1585,N_2968);
nand U3477 (N_3477,N_2879,N_2198);
xor U3478 (N_3478,N_2884,N_2820);
nor U3479 (N_3479,N_2473,N_2286);
and U3480 (N_3480,N_2672,N_2105);
nand U3481 (N_3481,N_1656,N_2828);
and U3482 (N_3482,N_2496,N_2657);
xor U3483 (N_3483,N_2356,N_2647);
nor U3484 (N_3484,N_2944,N_2290);
or U3485 (N_3485,N_1860,N_2437);
and U3486 (N_3486,N_1859,N_2212);
nand U3487 (N_3487,N_2808,N_2078);
nand U3488 (N_3488,N_2146,N_1985);
and U3489 (N_3489,N_1801,N_2267);
nand U3490 (N_3490,N_2809,N_2124);
and U3491 (N_3491,N_2099,N_2643);
or U3492 (N_3492,N_2111,N_1965);
or U3493 (N_3493,N_2374,N_2943);
nand U3494 (N_3494,N_1628,N_2274);
or U3495 (N_3495,N_2917,N_1806);
and U3496 (N_3496,N_2623,N_2865);
and U3497 (N_3497,N_2992,N_2466);
xor U3498 (N_3498,N_1977,N_1694);
and U3499 (N_3499,N_2444,N_2867);
nor U3500 (N_3500,N_2100,N_2488);
nor U3501 (N_3501,N_2667,N_2877);
and U3502 (N_3502,N_1713,N_2016);
and U3503 (N_3503,N_2202,N_2512);
xnor U3504 (N_3504,N_2559,N_1877);
nor U3505 (N_3505,N_2489,N_2393);
and U3506 (N_3506,N_2166,N_1841);
nand U3507 (N_3507,N_2890,N_1581);
xnor U3508 (N_3508,N_1879,N_2453);
nand U3509 (N_3509,N_2628,N_2081);
nand U3510 (N_3510,N_1800,N_2710);
xnor U3511 (N_3511,N_1664,N_1699);
and U3512 (N_3512,N_1605,N_2317);
nor U3513 (N_3513,N_1523,N_2322);
xor U3514 (N_3514,N_2522,N_1737);
or U3515 (N_3515,N_1988,N_2521);
and U3516 (N_3516,N_2261,N_2407);
xor U3517 (N_3517,N_2364,N_1731);
or U3518 (N_3518,N_2363,N_1980);
nand U3519 (N_3519,N_1594,N_2246);
xor U3520 (N_3520,N_2323,N_2997);
or U3521 (N_3521,N_1963,N_1640);
and U3522 (N_3522,N_1881,N_2418);
nand U3523 (N_3523,N_2502,N_2580);
xor U3524 (N_3524,N_1821,N_1787);
or U3525 (N_3525,N_2205,N_1722);
and U3526 (N_3526,N_2745,N_2565);
nor U3527 (N_3527,N_1611,N_2191);
or U3528 (N_3528,N_2727,N_2416);
nor U3529 (N_3529,N_2649,N_2050);
xnor U3530 (N_3530,N_2759,N_1612);
nor U3531 (N_3531,N_2515,N_2354);
nor U3532 (N_3532,N_2446,N_2963);
and U3533 (N_3533,N_1544,N_1924);
nand U3534 (N_3534,N_2908,N_2164);
or U3535 (N_3535,N_1874,N_1872);
nor U3536 (N_3536,N_2424,N_2903);
and U3537 (N_3537,N_1937,N_2608);
nand U3538 (N_3538,N_2786,N_1949);
and U3539 (N_3539,N_1767,N_1600);
and U3540 (N_3540,N_2882,N_1776);
nor U3541 (N_3541,N_2886,N_1549);
or U3542 (N_3542,N_2495,N_2014);
nand U3543 (N_3543,N_1978,N_2648);
xnor U3544 (N_3544,N_2926,N_1773);
or U3545 (N_3545,N_2504,N_1970);
nor U3546 (N_3546,N_1940,N_1735);
nor U3547 (N_3547,N_2769,N_1714);
nor U3548 (N_3548,N_2159,N_2799);
xor U3549 (N_3549,N_1558,N_1814);
xnor U3550 (N_3550,N_2722,N_1945);
and U3551 (N_3551,N_2003,N_2161);
xnor U3552 (N_3552,N_2956,N_1961);
nand U3553 (N_3553,N_1607,N_2965);
xor U3554 (N_3554,N_2032,N_2276);
and U3555 (N_3555,N_2602,N_1703);
nand U3556 (N_3556,N_2186,N_1520);
xor U3557 (N_3557,N_2282,N_1952);
and U3558 (N_3558,N_2539,N_2793);
nand U3559 (N_3559,N_1578,N_2834);
or U3560 (N_3560,N_2134,N_2806);
or U3561 (N_3561,N_1537,N_2540);
xor U3562 (N_3562,N_1686,N_2052);
nand U3563 (N_3563,N_2262,N_1502);
nor U3564 (N_3564,N_2103,N_1541);
xnor U3565 (N_3565,N_1974,N_2849);
or U3566 (N_3566,N_2171,N_2854);
nand U3567 (N_3567,N_2170,N_1724);
nand U3568 (N_3568,N_1647,N_2622);
nand U3569 (N_3569,N_2501,N_2981);
and U3570 (N_3570,N_2577,N_2718);
nor U3571 (N_3571,N_2687,N_2826);
xor U3572 (N_3572,N_2018,N_2655);
nand U3573 (N_3573,N_1650,N_1688);
xor U3574 (N_3574,N_2850,N_1738);
nor U3575 (N_3575,N_2604,N_2595);
or U3576 (N_3576,N_1939,N_2369);
nand U3577 (N_3577,N_1964,N_1802);
xor U3578 (N_3578,N_2650,N_1914);
xor U3579 (N_3579,N_2503,N_2916);
xor U3580 (N_3580,N_1741,N_2633);
or U3581 (N_3581,N_2036,N_2931);
and U3582 (N_3582,N_2048,N_2985);
nand U3583 (N_3583,N_2113,N_2468);
nand U3584 (N_3584,N_2610,N_1843);
nor U3585 (N_3585,N_2347,N_1608);
nand U3586 (N_3586,N_2199,N_2483);
or U3587 (N_3587,N_1519,N_2553);
and U3588 (N_3588,N_2915,N_2500);
xor U3589 (N_3589,N_2645,N_1584);
nand U3590 (N_3590,N_1734,N_1886);
nand U3591 (N_3591,N_2532,N_2999);
xnor U3592 (N_3592,N_2086,N_1711);
or U3593 (N_3593,N_2189,N_2733);
xnor U3594 (N_3594,N_2344,N_2057);
and U3595 (N_3595,N_1998,N_2712);
xor U3596 (N_3596,N_1799,N_2819);
nand U3597 (N_3597,N_1995,N_2781);
and U3598 (N_3598,N_2838,N_2938);
and U3599 (N_3599,N_2237,N_2678);
xnor U3600 (N_3600,N_2858,N_2238);
nand U3601 (N_3601,N_2912,N_1559);
xnor U3602 (N_3602,N_2079,N_2392);
nor U3603 (N_3603,N_2923,N_2581);
nor U3604 (N_3604,N_1796,N_1883);
and U3605 (N_3605,N_1707,N_2031);
or U3606 (N_3606,N_2067,N_2112);
nor U3607 (N_3607,N_2605,N_1851);
nor U3608 (N_3608,N_2872,N_2670);
nand U3609 (N_3609,N_2537,N_2896);
or U3610 (N_3610,N_1768,N_2897);
nand U3611 (N_3611,N_2914,N_1999);
xnor U3612 (N_3612,N_1700,N_2349);
or U3613 (N_3613,N_1909,N_1853);
nor U3614 (N_3614,N_1778,N_1783);
xor U3615 (N_3615,N_1752,N_1524);
nand U3616 (N_3616,N_2318,N_2060);
and U3617 (N_3617,N_1515,N_2695);
and U3618 (N_3618,N_2991,N_1527);
or U3619 (N_3619,N_2873,N_2517);
xnor U3620 (N_3620,N_2426,N_1923);
or U3621 (N_3621,N_2893,N_2639);
nand U3622 (N_3622,N_2750,N_2066);
nor U3623 (N_3623,N_2242,N_1566);
xor U3624 (N_3624,N_1813,N_2560);
xnor U3625 (N_3625,N_1750,N_2823);
nor U3626 (N_3626,N_2300,N_2822);
nor U3627 (N_3627,N_1917,N_2586);
and U3628 (N_3628,N_2109,N_2765);
or U3629 (N_3629,N_2258,N_2860);
or U3630 (N_3630,N_2904,N_1805);
and U3631 (N_3631,N_2024,N_1782);
nor U3632 (N_3632,N_1994,N_2526);
or U3633 (N_3633,N_2945,N_2074);
nand U3634 (N_3634,N_2803,N_1765);
or U3635 (N_3635,N_2283,N_2116);
nor U3636 (N_3636,N_2034,N_2127);
nand U3637 (N_3637,N_2133,N_2947);
nor U3638 (N_3638,N_2425,N_2333);
nand U3639 (N_3639,N_2736,N_1546);
or U3640 (N_3640,N_2862,N_2288);
nor U3641 (N_3641,N_2612,N_2693);
xor U3642 (N_3642,N_2551,N_2360);
or U3643 (N_3643,N_2974,N_1582);
nand U3644 (N_3644,N_2576,N_2054);
xnor U3645 (N_3645,N_2439,N_2187);
or U3646 (N_3646,N_2210,N_2234);
xnor U3647 (N_3647,N_2922,N_1712);
or U3648 (N_3648,N_2443,N_1838);
and U3649 (N_3649,N_2684,N_2240);
xor U3650 (N_3650,N_2729,N_2558);
nor U3651 (N_3651,N_2583,N_2990);
and U3652 (N_3652,N_2042,N_2265);
and U3653 (N_3653,N_2701,N_1729);
or U3654 (N_3654,N_2259,N_1680);
xnor U3655 (N_3655,N_2400,N_1842);
xor U3656 (N_3656,N_2689,N_2942);
and U3657 (N_3657,N_2721,N_2764);
and U3658 (N_3658,N_2431,N_2578);
nor U3659 (N_3659,N_1644,N_2871);
or U3660 (N_3660,N_2353,N_2994);
nand U3661 (N_3661,N_1501,N_1928);
or U3662 (N_3662,N_2651,N_2924);
nor U3663 (N_3663,N_2192,N_2448);
and U3664 (N_3664,N_2151,N_2744);
xnor U3665 (N_3665,N_1875,N_2671);
nand U3666 (N_3666,N_2984,N_2002);
nor U3667 (N_3667,N_1786,N_2043);
or U3668 (N_3668,N_1869,N_1583);
xnor U3669 (N_3669,N_1983,N_2523);
xor U3670 (N_3670,N_2534,N_2857);
and U3671 (N_3671,N_1716,N_2251);
and U3672 (N_3672,N_2957,N_2033);
nand U3673 (N_3673,N_2982,N_2160);
and U3674 (N_3674,N_2487,N_1593);
xor U3675 (N_3675,N_1882,N_2664);
nand U3676 (N_3676,N_1710,N_1929);
or U3677 (N_3677,N_2243,N_1969);
or U3678 (N_3678,N_2020,N_2533);
nor U3679 (N_3679,N_2107,N_1905);
nand U3680 (N_3680,N_2284,N_2047);
nand U3681 (N_3681,N_2370,N_2792);
and U3682 (N_3682,N_2094,N_2017);
and U3683 (N_3683,N_2095,N_2092);
or U3684 (N_3684,N_2070,N_2827);
xor U3685 (N_3685,N_2824,N_1570);
nand U3686 (N_3686,N_2429,N_1953);
or U3687 (N_3687,N_2201,N_1630);
xor U3688 (N_3688,N_1772,N_2694);
and U3689 (N_3689,N_2883,N_2635);
nand U3690 (N_3690,N_2368,N_1685);
and U3691 (N_3691,N_2334,N_1720);
xnor U3692 (N_3692,N_1876,N_1823);
and U3693 (N_3693,N_2746,N_2616);
nand U3694 (N_3694,N_1572,N_2615);
or U3695 (N_3695,N_1794,N_2069);
nor U3696 (N_3696,N_2554,N_2594);
xor U3697 (N_3697,N_2902,N_2030);
or U3698 (N_3698,N_2818,N_2310);
nor U3699 (N_3699,N_1652,N_2314);
xor U3700 (N_3700,N_1938,N_2419);
xnor U3701 (N_3701,N_2477,N_2751);
xor U3702 (N_3702,N_1646,N_2767);
nor U3703 (N_3703,N_2679,N_2084);
nor U3704 (N_3704,N_2677,N_2362);
nand U3705 (N_3705,N_2228,N_2881);
nor U3706 (N_3706,N_2598,N_2297);
or U3707 (N_3707,N_1655,N_1670);
nor U3708 (N_3708,N_2634,N_2138);
nor U3709 (N_3709,N_1625,N_2414);
nor U3710 (N_3710,N_1925,N_1548);
xnor U3711 (N_3711,N_2742,N_2224);
or U3712 (N_3712,N_2524,N_2479);
xor U3713 (N_3713,N_2391,N_2293);
xnor U3714 (N_3714,N_2798,N_1811);
and U3715 (N_3715,N_2121,N_2732);
xnor U3716 (N_3716,N_2249,N_1912);
nor U3717 (N_3717,N_2632,N_2383);
or U3718 (N_3718,N_2816,N_2008);
nand U3719 (N_3719,N_2330,N_2332);
or U3720 (N_3720,N_2708,N_2373);
nand U3721 (N_3721,N_2493,N_2255);
and U3722 (N_3722,N_2652,N_1839);
nand U3723 (N_3723,N_2420,N_1769);
nand U3724 (N_3724,N_1697,N_2123);
or U3725 (N_3725,N_1962,N_2039);
or U3726 (N_3726,N_2328,N_2817);
nand U3727 (N_3727,N_1602,N_1552);
and U3728 (N_3728,N_2505,N_2101);
nor U3729 (N_3729,N_2272,N_2472);
and U3730 (N_3730,N_1518,N_2190);
and U3731 (N_3731,N_1871,N_2176);
nor U3732 (N_3732,N_1526,N_1789);
or U3733 (N_3733,N_2102,N_1818);
or U3734 (N_3734,N_2961,N_2380);
or U3735 (N_3735,N_2724,N_2367);
and U3736 (N_3736,N_2097,N_2129);
xor U3737 (N_3737,N_2193,N_2705);
nand U3738 (N_3738,N_1689,N_2339);
and U3739 (N_3739,N_1715,N_2711);
nand U3740 (N_3740,N_2844,N_2153);
nor U3741 (N_3741,N_2889,N_2644);
nand U3742 (N_3742,N_2019,N_2856);
nand U3743 (N_3743,N_2492,N_2012);
and U3744 (N_3744,N_2298,N_2408);
nor U3745 (N_3745,N_2427,N_1645);
or U3746 (N_3746,N_2244,N_2338);
and U3747 (N_3747,N_2143,N_2788);
and U3748 (N_3748,N_2381,N_2629);
and U3749 (N_3749,N_2022,N_1893);
nor U3750 (N_3750,N_1626,N_1595);
and U3751 (N_3751,N_2631,N_2374);
or U3752 (N_3752,N_2540,N_2096);
xnor U3753 (N_3753,N_2131,N_2288);
xnor U3754 (N_3754,N_2553,N_2977);
nor U3755 (N_3755,N_2575,N_1631);
and U3756 (N_3756,N_2407,N_2966);
or U3757 (N_3757,N_2827,N_1653);
nor U3758 (N_3758,N_1723,N_1713);
or U3759 (N_3759,N_2975,N_2186);
nor U3760 (N_3760,N_1925,N_2504);
or U3761 (N_3761,N_2343,N_1819);
and U3762 (N_3762,N_2694,N_2353);
nand U3763 (N_3763,N_2619,N_2853);
xor U3764 (N_3764,N_1697,N_1772);
and U3765 (N_3765,N_2507,N_2495);
and U3766 (N_3766,N_2645,N_2197);
xnor U3767 (N_3767,N_2058,N_1983);
and U3768 (N_3768,N_1990,N_2003);
nand U3769 (N_3769,N_2791,N_2490);
xnor U3770 (N_3770,N_2693,N_2746);
nand U3771 (N_3771,N_1830,N_2793);
nor U3772 (N_3772,N_2519,N_2475);
or U3773 (N_3773,N_2691,N_1783);
nor U3774 (N_3774,N_2220,N_2645);
or U3775 (N_3775,N_2067,N_2386);
nor U3776 (N_3776,N_2261,N_2206);
or U3777 (N_3777,N_2867,N_2527);
or U3778 (N_3778,N_2377,N_2676);
or U3779 (N_3779,N_1876,N_2276);
nand U3780 (N_3780,N_2371,N_2750);
or U3781 (N_3781,N_2228,N_2638);
xor U3782 (N_3782,N_2427,N_1776);
and U3783 (N_3783,N_2717,N_2013);
nor U3784 (N_3784,N_2591,N_1508);
and U3785 (N_3785,N_2319,N_1844);
nor U3786 (N_3786,N_2589,N_2763);
nor U3787 (N_3787,N_2152,N_2912);
xnor U3788 (N_3788,N_2411,N_2381);
xnor U3789 (N_3789,N_1558,N_2348);
xor U3790 (N_3790,N_2380,N_1622);
nor U3791 (N_3791,N_2642,N_1866);
xnor U3792 (N_3792,N_2207,N_1695);
nor U3793 (N_3793,N_2175,N_1657);
nor U3794 (N_3794,N_2657,N_1897);
xor U3795 (N_3795,N_2219,N_2189);
xnor U3796 (N_3796,N_1648,N_2417);
xnor U3797 (N_3797,N_2956,N_2673);
and U3798 (N_3798,N_2975,N_2878);
xnor U3799 (N_3799,N_1851,N_2313);
and U3800 (N_3800,N_2433,N_1926);
or U3801 (N_3801,N_2849,N_2503);
nor U3802 (N_3802,N_1650,N_2086);
nor U3803 (N_3803,N_1840,N_2436);
xor U3804 (N_3804,N_2351,N_1583);
nand U3805 (N_3805,N_2281,N_1597);
or U3806 (N_3806,N_2527,N_1575);
nand U3807 (N_3807,N_1651,N_1613);
xnor U3808 (N_3808,N_2913,N_2305);
xor U3809 (N_3809,N_1673,N_2845);
xor U3810 (N_3810,N_2804,N_1511);
nand U3811 (N_3811,N_2832,N_2951);
nor U3812 (N_3812,N_2808,N_1583);
nor U3813 (N_3813,N_2992,N_2939);
and U3814 (N_3814,N_2851,N_2095);
and U3815 (N_3815,N_2705,N_1713);
xnor U3816 (N_3816,N_1717,N_2726);
xnor U3817 (N_3817,N_2792,N_1838);
nand U3818 (N_3818,N_2236,N_1871);
nand U3819 (N_3819,N_1839,N_2771);
xor U3820 (N_3820,N_2943,N_1533);
nand U3821 (N_3821,N_2285,N_2953);
nand U3822 (N_3822,N_1571,N_2935);
xnor U3823 (N_3823,N_2365,N_2805);
xor U3824 (N_3824,N_2194,N_2744);
or U3825 (N_3825,N_1845,N_2805);
xnor U3826 (N_3826,N_2003,N_1736);
xor U3827 (N_3827,N_1564,N_2207);
nand U3828 (N_3828,N_1523,N_2495);
xor U3829 (N_3829,N_1885,N_2023);
nor U3830 (N_3830,N_1814,N_1803);
and U3831 (N_3831,N_2659,N_1503);
nor U3832 (N_3832,N_1583,N_2683);
or U3833 (N_3833,N_2396,N_1716);
and U3834 (N_3834,N_2950,N_2499);
and U3835 (N_3835,N_2257,N_2252);
xnor U3836 (N_3836,N_2695,N_1558);
nand U3837 (N_3837,N_2399,N_2206);
or U3838 (N_3838,N_2353,N_2746);
xnor U3839 (N_3839,N_2364,N_2307);
or U3840 (N_3840,N_2962,N_2162);
xnor U3841 (N_3841,N_2244,N_2892);
nand U3842 (N_3842,N_1737,N_1571);
xor U3843 (N_3843,N_1866,N_2903);
and U3844 (N_3844,N_2393,N_1628);
and U3845 (N_3845,N_1733,N_2996);
xnor U3846 (N_3846,N_2919,N_2072);
or U3847 (N_3847,N_2786,N_2880);
nor U3848 (N_3848,N_2764,N_1915);
xor U3849 (N_3849,N_1848,N_2879);
nor U3850 (N_3850,N_1783,N_2019);
nor U3851 (N_3851,N_1672,N_2712);
and U3852 (N_3852,N_1717,N_2972);
nor U3853 (N_3853,N_1537,N_1882);
nor U3854 (N_3854,N_1851,N_2197);
and U3855 (N_3855,N_2101,N_2416);
or U3856 (N_3856,N_2222,N_2465);
nand U3857 (N_3857,N_1560,N_2661);
and U3858 (N_3858,N_2694,N_1968);
or U3859 (N_3859,N_2160,N_2069);
xnor U3860 (N_3860,N_2899,N_1671);
nor U3861 (N_3861,N_1928,N_1958);
and U3862 (N_3862,N_2231,N_1736);
and U3863 (N_3863,N_2950,N_2868);
and U3864 (N_3864,N_2702,N_1576);
or U3865 (N_3865,N_2081,N_2967);
and U3866 (N_3866,N_2673,N_2994);
nand U3867 (N_3867,N_2916,N_2970);
nor U3868 (N_3868,N_2143,N_2880);
and U3869 (N_3869,N_2554,N_2692);
nand U3870 (N_3870,N_1904,N_2412);
and U3871 (N_3871,N_2754,N_1813);
and U3872 (N_3872,N_2308,N_1721);
xnor U3873 (N_3873,N_2896,N_2351);
nor U3874 (N_3874,N_2249,N_2600);
nor U3875 (N_3875,N_1529,N_1921);
nor U3876 (N_3876,N_2945,N_2214);
and U3877 (N_3877,N_2677,N_2521);
and U3878 (N_3878,N_1890,N_2203);
and U3879 (N_3879,N_1699,N_1788);
nor U3880 (N_3880,N_2287,N_2771);
xnor U3881 (N_3881,N_1620,N_1750);
nor U3882 (N_3882,N_2762,N_1764);
nor U3883 (N_3883,N_2637,N_1881);
nor U3884 (N_3884,N_2368,N_1922);
or U3885 (N_3885,N_2601,N_2136);
nand U3886 (N_3886,N_2876,N_2835);
or U3887 (N_3887,N_1980,N_1694);
or U3888 (N_3888,N_1996,N_2408);
nor U3889 (N_3889,N_1657,N_1909);
nand U3890 (N_3890,N_2625,N_2531);
nand U3891 (N_3891,N_2924,N_2057);
and U3892 (N_3892,N_2559,N_1646);
xor U3893 (N_3893,N_2533,N_2314);
nor U3894 (N_3894,N_1695,N_2714);
and U3895 (N_3895,N_2757,N_2197);
or U3896 (N_3896,N_2453,N_2615);
and U3897 (N_3897,N_2256,N_2618);
or U3898 (N_3898,N_2166,N_2111);
and U3899 (N_3899,N_1840,N_2326);
and U3900 (N_3900,N_2711,N_1888);
nand U3901 (N_3901,N_1601,N_1980);
xnor U3902 (N_3902,N_2419,N_2642);
nor U3903 (N_3903,N_2455,N_2689);
xor U3904 (N_3904,N_1750,N_1833);
nor U3905 (N_3905,N_1987,N_1782);
xor U3906 (N_3906,N_2645,N_2372);
or U3907 (N_3907,N_2268,N_2145);
xnor U3908 (N_3908,N_2203,N_2567);
xor U3909 (N_3909,N_1608,N_1574);
nor U3910 (N_3910,N_2845,N_1823);
nand U3911 (N_3911,N_1713,N_2476);
or U3912 (N_3912,N_2691,N_1655);
or U3913 (N_3913,N_2532,N_2848);
or U3914 (N_3914,N_1989,N_2583);
or U3915 (N_3915,N_1550,N_1689);
nand U3916 (N_3916,N_1834,N_2023);
xnor U3917 (N_3917,N_1965,N_1848);
xnor U3918 (N_3918,N_2426,N_2318);
or U3919 (N_3919,N_1972,N_2456);
or U3920 (N_3920,N_2173,N_2355);
nor U3921 (N_3921,N_2074,N_1734);
and U3922 (N_3922,N_1792,N_2588);
or U3923 (N_3923,N_2521,N_2190);
and U3924 (N_3924,N_2777,N_2753);
or U3925 (N_3925,N_2654,N_2074);
or U3926 (N_3926,N_2771,N_1961);
xor U3927 (N_3927,N_2486,N_1558);
nand U3928 (N_3928,N_2285,N_1921);
nand U3929 (N_3929,N_2667,N_2561);
or U3930 (N_3930,N_2617,N_1923);
or U3931 (N_3931,N_1748,N_1967);
and U3932 (N_3932,N_2131,N_1620);
nor U3933 (N_3933,N_2725,N_2306);
xor U3934 (N_3934,N_1511,N_1689);
nor U3935 (N_3935,N_2521,N_2081);
nor U3936 (N_3936,N_2811,N_2443);
nor U3937 (N_3937,N_1967,N_2923);
nand U3938 (N_3938,N_1533,N_2203);
nor U3939 (N_3939,N_1502,N_2939);
nor U3940 (N_3940,N_2195,N_1795);
nand U3941 (N_3941,N_2307,N_2472);
nand U3942 (N_3942,N_2866,N_1998);
nand U3943 (N_3943,N_2202,N_1542);
and U3944 (N_3944,N_2460,N_2817);
and U3945 (N_3945,N_2567,N_2540);
nor U3946 (N_3946,N_2316,N_2855);
or U3947 (N_3947,N_1722,N_2809);
nor U3948 (N_3948,N_2033,N_1591);
xnor U3949 (N_3949,N_2921,N_2561);
nor U3950 (N_3950,N_2842,N_1968);
or U3951 (N_3951,N_2857,N_1956);
or U3952 (N_3952,N_2031,N_1864);
nand U3953 (N_3953,N_2772,N_2829);
nand U3954 (N_3954,N_1509,N_2103);
nor U3955 (N_3955,N_2670,N_2026);
nor U3956 (N_3956,N_2992,N_2674);
nand U3957 (N_3957,N_2701,N_2617);
nand U3958 (N_3958,N_2684,N_2283);
or U3959 (N_3959,N_2378,N_1995);
nand U3960 (N_3960,N_2837,N_2153);
or U3961 (N_3961,N_1770,N_2489);
or U3962 (N_3962,N_2375,N_1783);
nor U3963 (N_3963,N_2483,N_2702);
and U3964 (N_3964,N_2525,N_2222);
nor U3965 (N_3965,N_2955,N_1675);
xor U3966 (N_3966,N_2527,N_2560);
or U3967 (N_3967,N_2273,N_2775);
nand U3968 (N_3968,N_2725,N_2700);
and U3969 (N_3969,N_2956,N_1835);
and U3970 (N_3970,N_1819,N_2337);
nor U3971 (N_3971,N_2124,N_2858);
nor U3972 (N_3972,N_1867,N_1628);
and U3973 (N_3973,N_1528,N_1632);
nand U3974 (N_3974,N_1624,N_2204);
xnor U3975 (N_3975,N_1572,N_2527);
and U3976 (N_3976,N_2538,N_2391);
nand U3977 (N_3977,N_1890,N_2921);
nor U3978 (N_3978,N_2967,N_2530);
nor U3979 (N_3979,N_2300,N_2658);
xor U3980 (N_3980,N_2614,N_1736);
or U3981 (N_3981,N_2132,N_2014);
xor U3982 (N_3982,N_2870,N_1776);
xnor U3983 (N_3983,N_2886,N_2307);
and U3984 (N_3984,N_2915,N_1586);
or U3985 (N_3985,N_2546,N_1677);
and U3986 (N_3986,N_1659,N_1656);
and U3987 (N_3987,N_2893,N_1707);
xor U3988 (N_3988,N_2000,N_2185);
nand U3989 (N_3989,N_2501,N_2553);
nor U3990 (N_3990,N_2370,N_1547);
and U3991 (N_3991,N_2255,N_1536);
nor U3992 (N_3992,N_2616,N_2462);
or U3993 (N_3993,N_1543,N_2276);
or U3994 (N_3994,N_2770,N_2636);
or U3995 (N_3995,N_2482,N_2051);
nand U3996 (N_3996,N_2132,N_2745);
xnor U3997 (N_3997,N_1893,N_1877);
xor U3998 (N_3998,N_2028,N_2709);
and U3999 (N_3999,N_1678,N_1742);
nand U4000 (N_4000,N_2529,N_1975);
or U4001 (N_4001,N_2618,N_2479);
nor U4002 (N_4002,N_2577,N_2714);
xnor U4003 (N_4003,N_2630,N_2941);
nand U4004 (N_4004,N_1925,N_2764);
nand U4005 (N_4005,N_1750,N_1702);
nor U4006 (N_4006,N_2335,N_2398);
or U4007 (N_4007,N_2590,N_2761);
nor U4008 (N_4008,N_1905,N_1899);
xor U4009 (N_4009,N_2180,N_1613);
and U4010 (N_4010,N_2538,N_2368);
and U4011 (N_4011,N_1903,N_2103);
nor U4012 (N_4012,N_1694,N_1713);
xor U4013 (N_4013,N_2415,N_2502);
or U4014 (N_4014,N_2785,N_2194);
nor U4015 (N_4015,N_2994,N_2059);
xor U4016 (N_4016,N_2480,N_1500);
nand U4017 (N_4017,N_1683,N_2589);
and U4018 (N_4018,N_1567,N_2546);
or U4019 (N_4019,N_2658,N_1647);
nor U4020 (N_4020,N_2382,N_1718);
xnor U4021 (N_4021,N_2852,N_1587);
nor U4022 (N_4022,N_2848,N_2594);
nand U4023 (N_4023,N_1765,N_2138);
xnor U4024 (N_4024,N_2942,N_2286);
nand U4025 (N_4025,N_2456,N_2799);
nor U4026 (N_4026,N_2752,N_2629);
nand U4027 (N_4027,N_1747,N_2426);
or U4028 (N_4028,N_1519,N_1548);
and U4029 (N_4029,N_2566,N_2670);
and U4030 (N_4030,N_2245,N_2997);
nand U4031 (N_4031,N_2870,N_2285);
or U4032 (N_4032,N_1794,N_2373);
nand U4033 (N_4033,N_2172,N_1884);
and U4034 (N_4034,N_1657,N_2603);
or U4035 (N_4035,N_1938,N_2018);
xnor U4036 (N_4036,N_1835,N_2084);
and U4037 (N_4037,N_2985,N_1924);
or U4038 (N_4038,N_1868,N_2287);
nor U4039 (N_4039,N_2141,N_2466);
nor U4040 (N_4040,N_2147,N_2011);
xor U4041 (N_4041,N_1901,N_2707);
nor U4042 (N_4042,N_2457,N_2296);
xnor U4043 (N_4043,N_2754,N_2140);
xnor U4044 (N_4044,N_2694,N_2814);
nor U4045 (N_4045,N_1649,N_1995);
or U4046 (N_4046,N_2868,N_2489);
nor U4047 (N_4047,N_1579,N_1848);
or U4048 (N_4048,N_1619,N_2592);
nor U4049 (N_4049,N_2746,N_2352);
and U4050 (N_4050,N_2905,N_2353);
and U4051 (N_4051,N_1629,N_2009);
xor U4052 (N_4052,N_2862,N_2998);
nand U4053 (N_4053,N_2727,N_2704);
or U4054 (N_4054,N_2280,N_1676);
nor U4055 (N_4055,N_1641,N_2528);
xor U4056 (N_4056,N_1557,N_2096);
nand U4057 (N_4057,N_2282,N_2925);
nand U4058 (N_4058,N_2772,N_1664);
and U4059 (N_4059,N_2980,N_2695);
nand U4060 (N_4060,N_2331,N_2165);
and U4061 (N_4061,N_2366,N_1930);
and U4062 (N_4062,N_2121,N_2654);
nand U4063 (N_4063,N_1841,N_1515);
or U4064 (N_4064,N_2332,N_1722);
nand U4065 (N_4065,N_1827,N_2684);
and U4066 (N_4066,N_2740,N_2007);
nor U4067 (N_4067,N_2179,N_2808);
nand U4068 (N_4068,N_2720,N_2761);
nor U4069 (N_4069,N_1952,N_1979);
and U4070 (N_4070,N_2235,N_1956);
nand U4071 (N_4071,N_2216,N_2381);
nand U4072 (N_4072,N_1973,N_2602);
or U4073 (N_4073,N_2975,N_2949);
nor U4074 (N_4074,N_2517,N_2026);
nor U4075 (N_4075,N_2637,N_2861);
nand U4076 (N_4076,N_1562,N_2128);
nor U4077 (N_4077,N_2663,N_2088);
xnor U4078 (N_4078,N_1515,N_1937);
or U4079 (N_4079,N_2942,N_1911);
xor U4080 (N_4080,N_2177,N_1943);
and U4081 (N_4081,N_1872,N_1690);
and U4082 (N_4082,N_1692,N_1548);
nor U4083 (N_4083,N_2506,N_2130);
nor U4084 (N_4084,N_2620,N_2746);
and U4085 (N_4085,N_2746,N_2503);
and U4086 (N_4086,N_2018,N_2887);
or U4087 (N_4087,N_2189,N_2764);
nand U4088 (N_4088,N_2617,N_2271);
or U4089 (N_4089,N_1910,N_1967);
or U4090 (N_4090,N_2092,N_2736);
nor U4091 (N_4091,N_1706,N_2781);
or U4092 (N_4092,N_1973,N_2468);
or U4093 (N_4093,N_2636,N_2507);
or U4094 (N_4094,N_2830,N_2863);
or U4095 (N_4095,N_1954,N_1978);
or U4096 (N_4096,N_2377,N_2385);
nor U4097 (N_4097,N_2012,N_1530);
or U4098 (N_4098,N_2240,N_2233);
nor U4099 (N_4099,N_2522,N_1596);
and U4100 (N_4100,N_1819,N_1532);
nand U4101 (N_4101,N_1668,N_2495);
or U4102 (N_4102,N_2881,N_2646);
and U4103 (N_4103,N_2945,N_2211);
nand U4104 (N_4104,N_2085,N_2320);
nand U4105 (N_4105,N_2437,N_2648);
or U4106 (N_4106,N_2888,N_1792);
xnor U4107 (N_4107,N_2368,N_2165);
or U4108 (N_4108,N_2700,N_1745);
xnor U4109 (N_4109,N_2005,N_1980);
and U4110 (N_4110,N_2907,N_2656);
and U4111 (N_4111,N_2575,N_2344);
nand U4112 (N_4112,N_2452,N_1941);
or U4113 (N_4113,N_2376,N_2382);
and U4114 (N_4114,N_2714,N_1561);
or U4115 (N_4115,N_2150,N_1682);
nand U4116 (N_4116,N_2117,N_2292);
or U4117 (N_4117,N_1612,N_2641);
nor U4118 (N_4118,N_1509,N_1963);
nor U4119 (N_4119,N_2500,N_2242);
nor U4120 (N_4120,N_1828,N_2052);
xor U4121 (N_4121,N_2603,N_1799);
or U4122 (N_4122,N_2270,N_2125);
nor U4123 (N_4123,N_2845,N_2489);
xor U4124 (N_4124,N_1909,N_2261);
nand U4125 (N_4125,N_1721,N_1728);
xor U4126 (N_4126,N_1878,N_2494);
nor U4127 (N_4127,N_2263,N_2250);
and U4128 (N_4128,N_1692,N_1885);
xnor U4129 (N_4129,N_2442,N_2840);
and U4130 (N_4130,N_2844,N_2371);
xor U4131 (N_4131,N_2328,N_2359);
xnor U4132 (N_4132,N_2435,N_2469);
and U4133 (N_4133,N_2650,N_2619);
xor U4134 (N_4134,N_2854,N_2497);
nor U4135 (N_4135,N_2239,N_2450);
or U4136 (N_4136,N_1582,N_2817);
or U4137 (N_4137,N_1671,N_1535);
nor U4138 (N_4138,N_2167,N_1670);
or U4139 (N_4139,N_1952,N_1509);
nand U4140 (N_4140,N_2265,N_2951);
and U4141 (N_4141,N_2538,N_2895);
nor U4142 (N_4142,N_2095,N_2593);
nor U4143 (N_4143,N_2814,N_1769);
xor U4144 (N_4144,N_1610,N_1998);
and U4145 (N_4145,N_2026,N_1867);
nand U4146 (N_4146,N_2862,N_1893);
or U4147 (N_4147,N_2106,N_1579);
nand U4148 (N_4148,N_2777,N_2982);
xor U4149 (N_4149,N_2047,N_1528);
xor U4150 (N_4150,N_2846,N_2858);
and U4151 (N_4151,N_1871,N_2153);
nor U4152 (N_4152,N_1985,N_1704);
xnor U4153 (N_4153,N_1943,N_1760);
xor U4154 (N_4154,N_2918,N_2411);
or U4155 (N_4155,N_1579,N_2996);
nand U4156 (N_4156,N_2486,N_1639);
nor U4157 (N_4157,N_1828,N_2436);
nand U4158 (N_4158,N_2502,N_2711);
xor U4159 (N_4159,N_2599,N_2169);
nor U4160 (N_4160,N_1846,N_2416);
and U4161 (N_4161,N_2146,N_2360);
and U4162 (N_4162,N_1864,N_1690);
nand U4163 (N_4163,N_2452,N_1660);
nand U4164 (N_4164,N_1555,N_2055);
nand U4165 (N_4165,N_1760,N_1530);
xnor U4166 (N_4166,N_1806,N_1536);
xor U4167 (N_4167,N_2859,N_2648);
or U4168 (N_4168,N_1681,N_2347);
and U4169 (N_4169,N_1701,N_2369);
xor U4170 (N_4170,N_1904,N_1675);
or U4171 (N_4171,N_1677,N_2838);
or U4172 (N_4172,N_2291,N_2521);
xor U4173 (N_4173,N_2008,N_2498);
nor U4174 (N_4174,N_2620,N_1526);
or U4175 (N_4175,N_2963,N_2780);
xnor U4176 (N_4176,N_1637,N_2925);
nand U4177 (N_4177,N_2292,N_2058);
or U4178 (N_4178,N_1783,N_2846);
nand U4179 (N_4179,N_2513,N_1567);
xor U4180 (N_4180,N_2756,N_2855);
xor U4181 (N_4181,N_1868,N_2496);
and U4182 (N_4182,N_1732,N_2234);
nand U4183 (N_4183,N_1839,N_2272);
or U4184 (N_4184,N_2248,N_2563);
and U4185 (N_4185,N_2460,N_2594);
xnor U4186 (N_4186,N_1779,N_1643);
nor U4187 (N_4187,N_1782,N_2306);
nor U4188 (N_4188,N_2211,N_2255);
and U4189 (N_4189,N_2392,N_2834);
xnor U4190 (N_4190,N_1819,N_2916);
or U4191 (N_4191,N_2012,N_1541);
or U4192 (N_4192,N_1603,N_2321);
nand U4193 (N_4193,N_2457,N_2065);
or U4194 (N_4194,N_2843,N_1562);
xor U4195 (N_4195,N_2469,N_1582);
xnor U4196 (N_4196,N_1574,N_1686);
nor U4197 (N_4197,N_2801,N_1760);
or U4198 (N_4198,N_1952,N_2378);
or U4199 (N_4199,N_1527,N_1879);
nand U4200 (N_4200,N_2183,N_1961);
nor U4201 (N_4201,N_2775,N_2754);
xnor U4202 (N_4202,N_2742,N_2857);
nand U4203 (N_4203,N_1833,N_2823);
or U4204 (N_4204,N_1665,N_2979);
and U4205 (N_4205,N_2537,N_1527);
nor U4206 (N_4206,N_1598,N_2356);
nand U4207 (N_4207,N_2062,N_2904);
nor U4208 (N_4208,N_2224,N_2007);
nand U4209 (N_4209,N_2461,N_2785);
and U4210 (N_4210,N_2160,N_1768);
nor U4211 (N_4211,N_2455,N_1720);
and U4212 (N_4212,N_2507,N_2480);
and U4213 (N_4213,N_1718,N_1755);
nand U4214 (N_4214,N_2174,N_2533);
xnor U4215 (N_4215,N_2462,N_1516);
or U4216 (N_4216,N_2791,N_2556);
xor U4217 (N_4217,N_2915,N_2914);
xor U4218 (N_4218,N_2917,N_1605);
or U4219 (N_4219,N_2536,N_2663);
xnor U4220 (N_4220,N_2956,N_2486);
nor U4221 (N_4221,N_1919,N_2882);
nor U4222 (N_4222,N_2288,N_1705);
nor U4223 (N_4223,N_2302,N_2918);
or U4224 (N_4224,N_2468,N_2431);
xor U4225 (N_4225,N_1635,N_2002);
and U4226 (N_4226,N_2312,N_2766);
or U4227 (N_4227,N_2852,N_2874);
nand U4228 (N_4228,N_2948,N_2823);
and U4229 (N_4229,N_2857,N_2091);
or U4230 (N_4230,N_2732,N_2834);
nand U4231 (N_4231,N_2280,N_2929);
nand U4232 (N_4232,N_2745,N_2849);
nor U4233 (N_4233,N_1593,N_1970);
or U4234 (N_4234,N_2201,N_2154);
xnor U4235 (N_4235,N_2484,N_1692);
xnor U4236 (N_4236,N_2473,N_2953);
and U4237 (N_4237,N_1883,N_2372);
and U4238 (N_4238,N_2377,N_2711);
nor U4239 (N_4239,N_2911,N_1897);
xor U4240 (N_4240,N_2262,N_2420);
or U4241 (N_4241,N_2618,N_2842);
or U4242 (N_4242,N_2303,N_2509);
nand U4243 (N_4243,N_2459,N_1983);
or U4244 (N_4244,N_2751,N_2361);
xnor U4245 (N_4245,N_1744,N_2594);
and U4246 (N_4246,N_1721,N_2039);
or U4247 (N_4247,N_2180,N_1524);
nor U4248 (N_4248,N_1647,N_2917);
or U4249 (N_4249,N_2379,N_2070);
or U4250 (N_4250,N_2992,N_2410);
nand U4251 (N_4251,N_2086,N_2227);
or U4252 (N_4252,N_1866,N_2484);
nand U4253 (N_4253,N_1633,N_2033);
and U4254 (N_4254,N_1788,N_1997);
or U4255 (N_4255,N_2065,N_1744);
or U4256 (N_4256,N_1924,N_2716);
nor U4257 (N_4257,N_2600,N_1913);
or U4258 (N_4258,N_2075,N_1947);
nand U4259 (N_4259,N_2436,N_2621);
nor U4260 (N_4260,N_2874,N_2249);
or U4261 (N_4261,N_1836,N_1874);
nor U4262 (N_4262,N_2283,N_2195);
nor U4263 (N_4263,N_2695,N_2597);
xor U4264 (N_4264,N_2392,N_2869);
xor U4265 (N_4265,N_2582,N_1679);
or U4266 (N_4266,N_1661,N_2559);
or U4267 (N_4267,N_2818,N_1817);
or U4268 (N_4268,N_1521,N_2047);
and U4269 (N_4269,N_2922,N_2956);
and U4270 (N_4270,N_1571,N_2543);
or U4271 (N_4271,N_2700,N_2626);
or U4272 (N_4272,N_2177,N_2756);
and U4273 (N_4273,N_1787,N_1692);
nor U4274 (N_4274,N_1708,N_2430);
and U4275 (N_4275,N_2779,N_2921);
xor U4276 (N_4276,N_2824,N_2455);
nand U4277 (N_4277,N_2323,N_1894);
xnor U4278 (N_4278,N_2997,N_2823);
and U4279 (N_4279,N_2710,N_1919);
nand U4280 (N_4280,N_2645,N_2613);
xor U4281 (N_4281,N_2597,N_2853);
and U4282 (N_4282,N_2092,N_2081);
nand U4283 (N_4283,N_2049,N_2396);
xor U4284 (N_4284,N_2817,N_2736);
nand U4285 (N_4285,N_2780,N_2411);
xnor U4286 (N_4286,N_2559,N_1842);
or U4287 (N_4287,N_1826,N_1536);
nor U4288 (N_4288,N_1892,N_2989);
and U4289 (N_4289,N_2861,N_2651);
or U4290 (N_4290,N_2655,N_2150);
and U4291 (N_4291,N_1911,N_2550);
xnor U4292 (N_4292,N_2350,N_1765);
and U4293 (N_4293,N_2691,N_2015);
xor U4294 (N_4294,N_1913,N_2988);
nand U4295 (N_4295,N_2178,N_2738);
or U4296 (N_4296,N_1628,N_2022);
nor U4297 (N_4297,N_2439,N_2030);
nor U4298 (N_4298,N_2110,N_1793);
or U4299 (N_4299,N_1690,N_1543);
and U4300 (N_4300,N_1568,N_1885);
nand U4301 (N_4301,N_2365,N_2899);
xnor U4302 (N_4302,N_1730,N_2414);
nor U4303 (N_4303,N_2835,N_1878);
or U4304 (N_4304,N_2132,N_1721);
nand U4305 (N_4305,N_2995,N_2199);
nor U4306 (N_4306,N_2689,N_2697);
nand U4307 (N_4307,N_2309,N_2527);
nand U4308 (N_4308,N_1718,N_2451);
or U4309 (N_4309,N_1837,N_2575);
and U4310 (N_4310,N_2726,N_2517);
xor U4311 (N_4311,N_2220,N_2871);
nand U4312 (N_4312,N_1628,N_2417);
nand U4313 (N_4313,N_1975,N_2361);
nand U4314 (N_4314,N_1638,N_1976);
and U4315 (N_4315,N_2267,N_1988);
and U4316 (N_4316,N_1812,N_2209);
xnor U4317 (N_4317,N_1753,N_2029);
nor U4318 (N_4318,N_2436,N_2623);
or U4319 (N_4319,N_2625,N_1527);
xor U4320 (N_4320,N_2494,N_2088);
xor U4321 (N_4321,N_2914,N_2064);
and U4322 (N_4322,N_2259,N_1714);
and U4323 (N_4323,N_1721,N_1716);
nor U4324 (N_4324,N_2736,N_1995);
nor U4325 (N_4325,N_2555,N_2510);
nand U4326 (N_4326,N_2467,N_1775);
xnor U4327 (N_4327,N_2629,N_1890);
xor U4328 (N_4328,N_1686,N_2002);
and U4329 (N_4329,N_1558,N_2187);
xnor U4330 (N_4330,N_2147,N_1773);
and U4331 (N_4331,N_2025,N_2880);
or U4332 (N_4332,N_1750,N_1909);
and U4333 (N_4333,N_2196,N_2763);
nor U4334 (N_4334,N_2246,N_2241);
and U4335 (N_4335,N_2613,N_2267);
nand U4336 (N_4336,N_1909,N_2846);
nand U4337 (N_4337,N_2490,N_2767);
or U4338 (N_4338,N_2125,N_1554);
nand U4339 (N_4339,N_1891,N_1846);
xor U4340 (N_4340,N_2104,N_2036);
xor U4341 (N_4341,N_2554,N_2852);
nand U4342 (N_4342,N_2670,N_2359);
nor U4343 (N_4343,N_1647,N_2712);
nor U4344 (N_4344,N_1786,N_2683);
and U4345 (N_4345,N_2544,N_2426);
or U4346 (N_4346,N_1867,N_1632);
nand U4347 (N_4347,N_2622,N_2521);
or U4348 (N_4348,N_1914,N_1930);
and U4349 (N_4349,N_1987,N_2572);
or U4350 (N_4350,N_2575,N_2901);
nor U4351 (N_4351,N_2167,N_1744);
or U4352 (N_4352,N_1787,N_1960);
xnor U4353 (N_4353,N_2481,N_2468);
and U4354 (N_4354,N_2540,N_2270);
xnor U4355 (N_4355,N_2152,N_2190);
xnor U4356 (N_4356,N_1765,N_1824);
nand U4357 (N_4357,N_2439,N_1858);
nor U4358 (N_4358,N_1564,N_1625);
xor U4359 (N_4359,N_1794,N_2902);
or U4360 (N_4360,N_2785,N_2645);
and U4361 (N_4361,N_2774,N_2014);
nand U4362 (N_4362,N_2692,N_2863);
xnor U4363 (N_4363,N_2422,N_2216);
or U4364 (N_4364,N_1789,N_2587);
or U4365 (N_4365,N_1837,N_1985);
nand U4366 (N_4366,N_2171,N_2513);
or U4367 (N_4367,N_2054,N_2561);
nor U4368 (N_4368,N_2966,N_2372);
and U4369 (N_4369,N_1833,N_2030);
or U4370 (N_4370,N_2870,N_2265);
or U4371 (N_4371,N_2576,N_1832);
xnor U4372 (N_4372,N_1555,N_2047);
nor U4373 (N_4373,N_2978,N_2251);
or U4374 (N_4374,N_2377,N_1592);
nor U4375 (N_4375,N_2514,N_2875);
nor U4376 (N_4376,N_2571,N_2583);
nand U4377 (N_4377,N_2036,N_2397);
xor U4378 (N_4378,N_2502,N_2536);
xor U4379 (N_4379,N_1776,N_2402);
nor U4380 (N_4380,N_1806,N_1598);
xnor U4381 (N_4381,N_2191,N_2859);
and U4382 (N_4382,N_2015,N_2566);
xnor U4383 (N_4383,N_2759,N_2185);
nor U4384 (N_4384,N_1699,N_1826);
nor U4385 (N_4385,N_2362,N_2673);
nor U4386 (N_4386,N_1765,N_2876);
xnor U4387 (N_4387,N_2996,N_2402);
nor U4388 (N_4388,N_2087,N_1641);
and U4389 (N_4389,N_2796,N_2373);
or U4390 (N_4390,N_2667,N_2287);
nor U4391 (N_4391,N_1643,N_1670);
nor U4392 (N_4392,N_2476,N_1932);
nor U4393 (N_4393,N_1604,N_2539);
nor U4394 (N_4394,N_1742,N_1723);
nand U4395 (N_4395,N_1738,N_1779);
nand U4396 (N_4396,N_2111,N_2289);
or U4397 (N_4397,N_2148,N_1960);
or U4398 (N_4398,N_1958,N_2814);
or U4399 (N_4399,N_1632,N_2767);
and U4400 (N_4400,N_1551,N_2691);
nand U4401 (N_4401,N_1974,N_2359);
nor U4402 (N_4402,N_2348,N_1799);
nand U4403 (N_4403,N_2527,N_1601);
xnor U4404 (N_4404,N_2241,N_1717);
and U4405 (N_4405,N_2626,N_2573);
and U4406 (N_4406,N_2107,N_2815);
nor U4407 (N_4407,N_1626,N_2579);
nand U4408 (N_4408,N_2370,N_2116);
nand U4409 (N_4409,N_2075,N_2080);
xnor U4410 (N_4410,N_2925,N_2526);
or U4411 (N_4411,N_2280,N_2523);
nor U4412 (N_4412,N_1768,N_1653);
or U4413 (N_4413,N_2976,N_1698);
nor U4414 (N_4414,N_1533,N_1676);
xor U4415 (N_4415,N_2726,N_1790);
nand U4416 (N_4416,N_1879,N_2961);
and U4417 (N_4417,N_2592,N_2503);
and U4418 (N_4418,N_2677,N_1870);
or U4419 (N_4419,N_2409,N_1924);
and U4420 (N_4420,N_1952,N_2400);
nor U4421 (N_4421,N_2339,N_1730);
xnor U4422 (N_4422,N_2431,N_1868);
nand U4423 (N_4423,N_1675,N_2593);
or U4424 (N_4424,N_2430,N_2768);
and U4425 (N_4425,N_2049,N_1928);
and U4426 (N_4426,N_2454,N_1964);
or U4427 (N_4427,N_2379,N_1853);
or U4428 (N_4428,N_2816,N_1781);
nor U4429 (N_4429,N_2124,N_2884);
or U4430 (N_4430,N_2984,N_2867);
xnor U4431 (N_4431,N_1561,N_2833);
nor U4432 (N_4432,N_2609,N_2915);
nor U4433 (N_4433,N_2261,N_2213);
nor U4434 (N_4434,N_2483,N_2484);
nand U4435 (N_4435,N_1956,N_2591);
or U4436 (N_4436,N_2259,N_2481);
or U4437 (N_4437,N_2387,N_2358);
xnor U4438 (N_4438,N_1511,N_2242);
or U4439 (N_4439,N_1788,N_2543);
nand U4440 (N_4440,N_2952,N_1886);
xnor U4441 (N_4441,N_1844,N_1797);
and U4442 (N_4442,N_2669,N_2110);
nor U4443 (N_4443,N_2309,N_2894);
and U4444 (N_4444,N_2029,N_2852);
or U4445 (N_4445,N_2665,N_2137);
and U4446 (N_4446,N_2638,N_2361);
or U4447 (N_4447,N_2007,N_1786);
nand U4448 (N_4448,N_1570,N_2695);
nand U4449 (N_4449,N_2535,N_1903);
xnor U4450 (N_4450,N_2516,N_1777);
or U4451 (N_4451,N_2130,N_2454);
nor U4452 (N_4452,N_2617,N_1860);
and U4453 (N_4453,N_1607,N_2013);
nor U4454 (N_4454,N_2136,N_2415);
or U4455 (N_4455,N_2413,N_1568);
xor U4456 (N_4456,N_1507,N_2172);
or U4457 (N_4457,N_1853,N_2711);
nor U4458 (N_4458,N_2869,N_2650);
or U4459 (N_4459,N_2991,N_2477);
xnor U4460 (N_4460,N_2881,N_1789);
or U4461 (N_4461,N_2403,N_1854);
or U4462 (N_4462,N_1593,N_2379);
or U4463 (N_4463,N_2602,N_2202);
nand U4464 (N_4464,N_2381,N_2021);
or U4465 (N_4465,N_1698,N_1741);
xor U4466 (N_4466,N_2973,N_1658);
xnor U4467 (N_4467,N_2080,N_2857);
xor U4468 (N_4468,N_2981,N_1532);
nand U4469 (N_4469,N_2129,N_2265);
or U4470 (N_4470,N_1528,N_2327);
and U4471 (N_4471,N_2992,N_2362);
nand U4472 (N_4472,N_1886,N_1715);
nor U4473 (N_4473,N_2068,N_1635);
or U4474 (N_4474,N_2541,N_2647);
or U4475 (N_4475,N_2089,N_2202);
nor U4476 (N_4476,N_2652,N_2469);
or U4477 (N_4477,N_1599,N_1772);
nor U4478 (N_4478,N_2040,N_2390);
or U4479 (N_4479,N_1929,N_2028);
nand U4480 (N_4480,N_1592,N_1913);
and U4481 (N_4481,N_2892,N_1912);
nand U4482 (N_4482,N_1801,N_2700);
xnor U4483 (N_4483,N_2713,N_2931);
nand U4484 (N_4484,N_2221,N_2556);
and U4485 (N_4485,N_2905,N_1648);
nand U4486 (N_4486,N_2370,N_1691);
and U4487 (N_4487,N_1854,N_2407);
nor U4488 (N_4488,N_2147,N_2185);
and U4489 (N_4489,N_2767,N_1708);
and U4490 (N_4490,N_2311,N_2731);
and U4491 (N_4491,N_1851,N_2615);
and U4492 (N_4492,N_2868,N_2087);
and U4493 (N_4493,N_2933,N_1655);
or U4494 (N_4494,N_1836,N_1535);
nor U4495 (N_4495,N_2567,N_2321);
and U4496 (N_4496,N_1633,N_2051);
and U4497 (N_4497,N_1753,N_2291);
and U4498 (N_4498,N_1721,N_2725);
nor U4499 (N_4499,N_1690,N_1737);
nor U4500 (N_4500,N_3738,N_3389);
nand U4501 (N_4501,N_3044,N_3612);
nand U4502 (N_4502,N_3696,N_3261);
or U4503 (N_4503,N_3249,N_3663);
nand U4504 (N_4504,N_4104,N_3932);
and U4505 (N_4505,N_4206,N_4465);
and U4506 (N_4506,N_3807,N_3891);
nor U4507 (N_4507,N_3592,N_3434);
xnor U4508 (N_4508,N_3836,N_3223);
nand U4509 (N_4509,N_3340,N_4295);
nor U4510 (N_4510,N_4482,N_4382);
and U4511 (N_4511,N_3462,N_4256);
nand U4512 (N_4512,N_3130,N_3282);
nand U4513 (N_4513,N_3391,N_3294);
or U4514 (N_4514,N_3726,N_4394);
and U4515 (N_4515,N_3113,N_3021);
or U4516 (N_4516,N_3424,N_4257);
nor U4517 (N_4517,N_4378,N_3270);
nand U4518 (N_4518,N_3847,N_3892);
or U4519 (N_4519,N_3948,N_4049);
nand U4520 (N_4520,N_4313,N_3087);
or U4521 (N_4521,N_3715,N_3927);
xnor U4522 (N_4522,N_3097,N_4447);
and U4523 (N_4523,N_4199,N_3957);
nor U4524 (N_4524,N_3137,N_3503);
or U4525 (N_4525,N_3421,N_3330);
xor U4526 (N_4526,N_4287,N_3555);
nand U4527 (N_4527,N_3269,N_3737);
nand U4528 (N_4528,N_3474,N_3022);
xor U4529 (N_4529,N_4072,N_3094);
or U4530 (N_4530,N_3037,N_3714);
and U4531 (N_4531,N_4362,N_3406);
xnor U4532 (N_4532,N_4360,N_4121);
nor U4533 (N_4533,N_3817,N_3949);
xnor U4534 (N_4534,N_3786,N_3427);
xor U4535 (N_4535,N_3710,N_4216);
xnor U4536 (N_4536,N_4397,N_3335);
nor U4537 (N_4537,N_4289,N_3297);
or U4538 (N_4538,N_3851,N_3363);
and U4539 (N_4539,N_3060,N_4123);
nand U4540 (N_4540,N_4327,N_4107);
nand U4541 (N_4541,N_3532,N_4031);
nand U4542 (N_4542,N_4419,N_3005);
nor U4543 (N_4543,N_3629,N_3224);
xnor U4544 (N_4544,N_3546,N_3144);
nor U4545 (N_4545,N_4288,N_3965);
xnor U4546 (N_4546,N_3753,N_4304);
nand U4547 (N_4547,N_3093,N_4219);
nand U4548 (N_4548,N_4489,N_3562);
or U4549 (N_4549,N_3175,N_3861);
xor U4550 (N_4550,N_4042,N_3806);
or U4551 (N_4551,N_3325,N_3068);
xor U4552 (N_4552,N_3112,N_3464);
nor U4553 (N_4553,N_3413,N_3909);
xor U4554 (N_4554,N_3941,N_3057);
xnor U4555 (N_4555,N_3038,N_3517);
nor U4556 (N_4556,N_3179,N_3566);
nor U4557 (N_4557,N_3104,N_3796);
xor U4558 (N_4558,N_3230,N_4498);
nand U4559 (N_4559,N_4149,N_3280);
nand U4560 (N_4560,N_3305,N_3557);
nand U4561 (N_4561,N_4015,N_4366);
xor U4562 (N_4562,N_3442,N_3430);
nor U4563 (N_4563,N_4263,N_3400);
nor U4564 (N_4564,N_3604,N_3997);
nor U4565 (N_4565,N_4311,N_3480);
nand U4566 (N_4566,N_4211,N_3425);
nand U4567 (N_4567,N_3581,N_4208);
xnor U4568 (N_4568,N_3866,N_3132);
and U4569 (N_4569,N_4413,N_3928);
nor U4570 (N_4570,N_4356,N_3687);
nand U4571 (N_4571,N_3893,N_3667);
and U4572 (N_4572,N_3222,N_4492);
xor U4573 (N_4573,N_3247,N_3617);
nor U4574 (N_4574,N_3935,N_3439);
nor U4575 (N_4575,N_3128,N_3706);
nand U4576 (N_4576,N_3619,N_3189);
xnor U4577 (N_4577,N_4431,N_3039);
xnor U4578 (N_4578,N_3752,N_3637);
and U4579 (N_4579,N_3410,N_3301);
xnor U4580 (N_4580,N_4195,N_4071);
xnor U4581 (N_4581,N_3513,N_3934);
and U4582 (N_4582,N_3253,N_3493);
and U4583 (N_4583,N_4114,N_3390);
or U4584 (N_4584,N_3457,N_3521);
nor U4585 (N_4585,N_3600,N_3088);
nand U4586 (N_4586,N_3334,N_3947);
and U4587 (N_4587,N_3518,N_4461);
and U4588 (N_4588,N_3755,N_3489);
or U4589 (N_4589,N_3378,N_3570);
and U4590 (N_4590,N_4106,N_4325);
or U4591 (N_4591,N_3880,N_3913);
or U4592 (N_4592,N_4353,N_3638);
xnor U4593 (N_4593,N_3275,N_4004);
and U4594 (N_4594,N_3242,N_3746);
nand U4595 (N_4595,N_3551,N_3534);
xnor U4596 (N_4596,N_4487,N_3497);
or U4597 (N_4597,N_4010,N_4167);
and U4598 (N_4598,N_3114,N_4406);
xor U4599 (N_4599,N_4012,N_3279);
nor U4600 (N_4600,N_4109,N_3122);
xor U4601 (N_4601,N_3484,N_3429);
nor U4602 (N_4602,N_3111,N_3165);
or U4603 (N_4603,N_3998,N_3862);
or U4604 (N_4604,N_3795,N_3312);
and U4605 (N_4605,N_4145,N_3688);
and U4606 (N_4606,N_4280,N_3827);
and U4607 (N_4607,N_3085,N_3736);
nand U4608 (N_4608,N_3561,N_3857);
nand U4609 (N_4609,N_3138,N_3382);
xor U4610 (N_4610,N_3772,N_3356);
or U4611 (N_4611,N_3673,N_4125);
nor U4612 (N_4612,N_3315,N_3359);
nor U4613 (N_4613,N_4390,N_3770);
xnor U4614 (N_4614,N_3333,N_4239);
xnor U4615 (N_4615,N_3613,N_4450);
xor U4616 (N_4616,N_3593,N_3754);
xnor U4617 (N_4617,N_3731,N_3680);
xnor U4618 (N_4618,N_3336,N_4091);
xor U4619 (N_4619,N_3188,N_3103);
or U4620 (N_4620,N_3749,N_3956);
xor U4621 (N_4621,N_3937,N_3840);
xor U4622 (N_4622,N_3887,N_4395);
nor U4623 (N_4623,N_3106,N_3730);
and U4624 (N_4624,N_4210,N_4365);
nor U4625 (N_4625,N_3367,N_3711);
and U4626 (N_4626,N_3856,N_4359);
xnor U4627 (N_4627,N_3906,N_3785);
and U4628 (N_4628,N_3086,N_3853);
xnor U4629 (N_4629,N_4369,N_3951);
nor U4630 (N_4630,N_3355,N_3241);
nand U4631 (N_4631,N_3449,N_3184);
and U4632 (N_4632,N_3777,N_4396);
and U4633 (N_4633,N_3461,N_3441);
xor U4634 (N_4634,N_3623,N_3659);
or U4635 (N_4635,N_3601,N_3234);
or U4636 (N_4636,N_4120,N_4418);
nand U4637 (N_4637,N_3496,N_4126);
nor U4638 (N_4638,N_3860,N_4285);
nand U4639 (N_4639,N_3778,N_4033);
nor U4640 (N_4640,N_3990,N_4264);
nor U4641 (N_4641,N_3665,N_3588);
nor U4642 (N_4642,N_3351,N_3643);
and U4643 (N_4643,N_3048,N_3964);
xor U4644 (N_4644,N_3811,N_3712);
nor U4645 (N_4645,N_3759,N_3961);
nor U4646 (N_4646,N_3487,N_3657);
nand U4647 (N_4647,N_4217,N_3875);
and U4648 (N_4648,N_3285,N_4466);
or U4649 (N_4649,N_3215,N_3411);
or U4650 (N_4650,N_4041,N_3813);
nand U4651 (N_4651,N_4458,N_3842);
or U4652 (N_4652,N_3292,N_4053);
or U4653 (N_4653,N_3447,N_4028);
nand U4654 (N_4654,N_4163,N_4317);
nor U4655 (N_4655,N_3530,N_3058);
or U4656 (N_4656,N_3370,N_4349);
or U4657 (N_4657,N_3257,N_4342);
xor U4658 (N_4658,N_3975,N_3703);
or U4659 (N_4659,N_3376,N_4029);
nor U4660 (N_4660,N_3407,N_3290);
nand U4661 (N_4661,N_3387,N_3155);
nor U4662 (N_4662,N_3559,N_4261);
nand U4663 (N_4663,N_3074,N_4411);
and U4664 (N_4664,N_4456,N_3721);
nor U4665 (N_4665,N_3092,N_3879);
or U4666 (N_4666,N_3682,N_3101);
and U4667 (N_4667,N_3485,N_4192);
nand U4668 (N_4668,N_3606,N_3286);
or U4669 (N_4669,N_3140,N_3549);
nand U4670 (N_4670,N_3149,N_3541);
and U4671 (N_4671,N_4240,N_3126);
or U4672 (N_4672,N_3153,N_3668);
nand U4673 (N_4673,N_3124,N_3670);
or U4674 (N_4674,N_3550,N_4115);
xnor U4675 (N_4675,N_4426,N_4344);
or U4676 (N_4676,N_3248,N_4241);
nor U4677 (N_4677,N_3251,N_3078);
and U4678 (N_4678,N_3473,N_3708);
nand U4679 (N_4679,N_4139,N_3298);
or U4680 (N_4680,N_4337,N_3775);
or U4681 (N_4681,N_4333,N_4309);
or U4682 (N_4682,N_4372,N_3671);
nor U4683 (N_4683,N_3662,N_3147);
and U4684 (N_4684,N_4484,N_3574);
xor U4685 (N_4685,N_3723,N_3584);
and U4686 (N_4686,N_3924,N_4491);
and U4687 (N_4687,N_3416,N_3472);
or U4688 (N_4688,N_3573,N_3849);
or U4689 (N_4689,N_3564,N_3182);
nand U4690 (N_4690,N_4370,N_3426);
and U4691 (N_4691,N_3402,N_3572);
xor U4692 (N_4692,N_3996,N_3790);
nand U4693 (N_4693,N_4446,N_3967);
xor U4694 (N_4694,N_4059,N_4069);
xor U4695 (N_4695,N_3707,N_3156);
nor U4696 (N_4696,N_3963,N_3912);
or U4697 (N_4697,N_3739,N_3810);
or U4698 (N_4698,N_4250,N_3850);
nor U4699 (N_4699,N_4310,N_3004);
nor U4700 (N_4700,N_3970,N_4490);
and U4701 (N_4701,N_4300,N_4093);
nand U4702 (N_4702,N_4476,N_3198);
nand U4703 (N_4703,N_3586,N_3012);
and U4704 (N_4704,N_4019,N_4364);
or U4705 (N_4705,N_4132,N_3705);
and U4706 (N_4706,N_3616,N_3089);
or U4707 (N_4707,N_3864,N_3168);
nand U4708 (N_4708,N_4080,N_3405);
nand U4709 (N_4709,N_4144,N_4334);
and U4710 (N_4710,N_3832,N_3329);
xor U4711 (N_4711,N_4213,N_4345);
or U4712 (N_4712,N_4279,N_3268);
and U4713 (N_4713,N_3758,N_4226);
and U4714 (N_4714,N_3652,N_3505);
nand U4715 (N_4715,N_3898,N_3722);
or U4716 (N_4716,N_3981,N_3193);
xor U4717 (N_4717,N_3571,N_3107);
and U4718 (N_4718,N_3494,N_4453);
nor U4719 (N_4719,N_3046,N_3266);
or U4720 (N_4720,N_3980,N_3159);
and U4721 (N_4721,N_3150,N_3944);
and U4722 (N_4722,N_4255,N_4190);
xnor U4723 (N_4723,N_3302,N_3458);
xnor U4724 (N_4724,N_4194,N_3666);
or U4725 (N_4725,N_4005,N_3977);
xor U4726 (N_4726,N_3252,N_3782);
nand U4727 (N_4727,N_4245,N_3553);
xor U4728 (N_4728,N_3690,N_3255);
xnor U4729 (N_4729,N_4291,N_3139);
xnor U4730 (N_4730,N_3653,N_3136);
or U4731 (N_4731,N_4352,N_4314);
or U4732 (N_4732,N_4469,N_3774);
xnor U4733 (N_4733,N_3209,N_4141);
or U4734 (N_4734,N_3214,N_3904);
nor U4735 (N_4735,N_3431,N_4463);
nor U4736 (N_4736,N_4436,N_4297);
and U4737 (N_4737,N_3109,N_3542);
xnor U4738 (N_4738,N_3296,N_3056);
nand U4739 (N_4739,N_3190,N_4212);
and U4740 (N_4740,N_3191,N_4455);
and U4741 (N_4741,N_3900,N_4045);
nor U4742 (N_4742,N_3558,N_4388);
and U4743 (N_4743,N_4227,N_3834);
or U4744 (N_4744,N_3797,N_3733);
nor U4745 (N_4745,N_3920,N_3740);
or U4746 (N_4746,N_3554,N_3787);
nand U4747 (N_4747,N_3369,N_4242);
and U4748 (N_4748,N_4330,N_4203);
nand U4749 (N_4749,N_3066,N_3015);
nor U4750 (N_4750,N_3545,N_3640);
nor U4751 (N_4751,N_3658,N_3243);
xor U4752 (N_4752,N_4252,N_3865);
xor U4753 (N_4753,N_4236,N_4262);
or U4754 (N_4754,N_3470,N_3216);
nor U4755 (N_4755,N_3135,N_3311);
or U4756 (N_4756,N_3271,N_3764);
and U4757 (N_4757,N_3958,N_3256);
nand U4758 (N_4758,N_4368,N_4315);
or U4759 (N_4759,N_3694,N_4427);
and U4760 (N_4760,N_4068,N_4497);
xnor U4761 (N_4761,N_3664,N_3318);
or U4762 (N_4762,N_4493,N_3693);
and U4763 (N_4763,N_3615,N_4129);
and U4764 (N_4764,N_3281,N_3835);
and U4765 (N_4765,N_3988,N_4083);
nor U4766 (N_4766,N_3897,N_3506);
xor U4767 (N_4767,N_3531,N_4408);
or U4768 (N_4768,N_3767,N_3634);
or U4769 (N_4769,N_4283,N_4347);
or U4770 (N_4770,N_4034,N_3669);
nor U4771 (N_4771,N_3645,N_4063);
xnor U4772 (N_4772,N_3527,N_3784);
xnor U4773 (N_4773,N_3440,N_4156);
or U4774 (N_4774,N_4014,N_4001);
nor U4775 (N_4775,N_3729,N_4016);
nand U4776 (N_4776,N_3018,N_4169);
xnor U4777 (N_4777,N_3076,N_4064);
nor U4778 (N_4778,N_3308,N_4277);
nand U4779 (N_4779,N_4158,N_3742);
and U4780 (N_4780,N_4119,N_3220);
nand U4781 (N_4781,N_3953,N_3463);
xor U4782 (N_4782,N_3915,N_4374);
xor U4783 (N_4783,N_4073,N_3192);
or U4784 (N_4784,N_4273,N_4075);
or U4785 (N_4785,N_3607,N_4354);
xor U4786 (N_4786,N_3686,N_3969);
or U4787 (N_4787,N_3627,N_4112);
xor U4788 (N_4788,N_3199,N_4322);
or U4789 (N_4789,N_3419,N_3283);
or U4790 (N_4790,N_4017,N_4228);
nor U4791 (N_4791,N_4150,N_4441);
or U4792 (N_4792,N_3183,N_3435);
and U4793 (N_4793,N_3446,N_4442);
nand U4794 (N_4794,N_3264,N_3002);
nor U4795 (N_4795,N_3360,N_3852);
nand U4796 (N_4796,N_3186,N_4133);
xor U4797 (N_4797,N_4381,N_3217);
nor U4798 (N_4798,N_3259,N_3129);
and U4799 (N_4799,N_3701,N_3621);
nand U4800 (N_4800,N_3013,N_3535);
xnor U4801 (N_4801,N_3603,N_3397);
nand U4802 (N_4802,N_4409,N_3403);
nor U4803 (N_4803,N_4477,N_3418);
nor U4804 (N_4804,N_3151,N_3141);
or U4805 (N_4805,N_3077,N_3569);
or U4806 (N_4806,N_3067,N_3524);
nor U4807 (N_4807,N_3160,N_3986);
nor U4808 (N_4808,N_3143,N_4165);
and U4809 (N_4809,N_3587,N_4189);
and U4810 (N_4810,N_4043,N_3881);
xor U4811 (N_4811,N_3760,N_4100);
and U4812 (N_4812,N_3492,N_3218);
nand U4813 (N_4813,N_4421,N_4428);
nor U4814 (N_4814,N_3973,N_4435);
or U4815 (N_4815,N_3792,N_3033);
and U4816 (N_4816,N_4258,N_3029);
and U4817 (N_4817,N_3245,N_4022);
and U4818 (N_4818,N_4380,N_3519);
xnor U4819 (N_4819,N_3133,N_4479);
xnor U4820 (N_4820,N_4024,N_3971);
or U4821 (N_4821,N_3236,N_4050);
nor U4822 (N_4822,N_4485,N_3979);
nor U4823 (N_4823,N_3460,N_3848);
nand U4824 (N_4824,N_3206,N_3695);
nor U4825 (N_4825,N_4299,N_4478);
nor U4826 (N_4826,N_3233,N_3121);
xor U4827 (N_4827,N_3846,N_4102);
or U4828 (N_4828,N_3793,N_4302);
nand U4829 (N_4829,N_3942,N_3520);
xnor U4830 (N_4830,N_4124,N_4218);
nand U4831 (N_4831,N_3905,N_3577);
nor U4832 (N_4832,N_3801,N_3870);
and U4833 (N_4833,N_3594,N_3373);
or U4834 (N_4834,N_3872,N_3322);
xnor U4835 (N_4835,N_3580,N_4183);
and U4836 (N_4836,N_3277,N_3780);
or U4837 (N_4837,N_3874,N_3952);
xnor U4838 (N_4838,N_4018,N_3936);
nand U4839 (N_4839,N_3877,N_4009);
nand U4840 (N_4840,N_4496,N_4096);
and U4841 (N_4841,N_3211,N_4229);
nand U4842 (N_4842,N_3125,N_4243);
nor U4843 (N_4843,N_3345,N_3522);
nor U4844 (N_4844,N_4331,N_3099);
nor U4845 (N_4845,N_3450,N_3576);
and U4846 (N_4846,N_4099,N_4131);
xnor U4847 (N_4847,N_3393,N_3328);
nor U4848 (N_4848,N_3683,N_4305);
xnor U4849 (N_4849,N_4451,N_3946);
nor U4850 (N_4850,N_4276,N_3762);
xor U4851 (N_4851,N_4052,N_4320);
or U4852 (N_4852,N_3808,N_3278);
and U4853 (N_4853,N_4101,N_4298);
and U4854 (N_4854,N_3123,N_3000);
or U4855 (N_4855,N_4367,N_3228);
and U4856 (N_4856,N_3728,N_4201);
or U4857 (N_4857,N_4417,N_3174);
or U4858 (N_4858,N_4400,N_3339);
xnor U4859 (N_4859,N_3859,N_3999);
and U4860 (N_4860,N_3011,N_4020);
nand U4861 (N_4861,N_3704,N_3116);
nand U4862 (N_4862,N_3428,N_3317);
and U4863 (N_4863,N_3547,N_4248);
or U4864 (N_4864,N_3052,N_3326);
nor U4865 (N_4865,N_3933,N_3080);
and U4866 (N_4866,N_4346,N_4215);
xnor U4867 (N_4867,N_3105,N_3455);
xor U4868 (N_4868,N_3829,N_4225);
and U4869 (N_4869,N_4260,N_3609);
nand U4870 (N_4870,N_3036,N_3020);
nand U4871 (N_4871,N_3644,N_3605);
nand U4872 (N_4872,N_4172,N_3713);
or U4873 (N_4873,N_3632,N_3916);
xnor U4874 (N_4874,N_3984,N_4110);
nand U4875 (N_4875,N_3938,N_3639);
or U4876 (N_4876,N_3043,N_4232);
nand U4877 (N_4877,N_3741,N_3830);
xnor U4878 (N_4878,N_4200,N_3172);
or U4879 (N_4879,N_3955,N_3353);
or U4880 (N_4880,N_3922,N_3061);
or U4881 (N_4881,N_3161,N_3822);
nand U4882 (N_4882,N_3751,N_3047);
nor U4883 (N_4883,N_4293,N_4205);
and U4884 (N_4884,N_3420,N_3203);
nand U4885 (N_4885,N_3395,N_3091);
nor U4886 (N_4886,N_3945,N_3779);
nand U4887 (N_4887,N_3533,N_3661);
and U4888 (N_4888,N_4113,N_3173);
nor U4889 (N_4889,N_4452,N_3486);
xor U4890 (N_4890,N_4274,N_4142);
nand U4891 (N_4891,N_4323,N_3903);
or U4892 (N_4892,N_3219,N_3392);
nand U4893 (N_4893,N_3055,N_4003);
and U4894 (N_4894,N_4061,N_3119);
or U4895 (N_4895,N_3802,N_3293);
or U4896 (N_4896,N_4220,N_3364);
nand U4897 (N_4897,N_4209,N_4058);
nor U4898 (N_4898,N_4000,N_3525);
and U4899 (N_4899,N_4341,N_3647);
and U4900 (N_4900,N_4097,N_3347);
nand U4901 (N_4901,N_4433,N_3700);
or U4902 (N_4902,N_3982,N_4148);
or U4903 (N_4903,N_4173,N_4422);
or U4904 (N_4904,N_4281,N_3678);
and U4905 (N_4905,N_3498,N_3890);
nand U4906 (N_4906,N_3511,N_4087);
or U4907 (N_4907,N_3719,N_3110);
nand U4908 (N_4908,N_4384,N_3824);
or U4909 (N_4909,N_3943,N_4038);
nor U4910 (N_4910,N_4335,N_4412);
xnor U4911 (N_4911,N_3438,N_3907);
or U4912 (N_4912,N_3100,N_4157);
nand U4913 (N_4913,N_3783,N_4006);
xnor U4914 (N_4914,N_4207,N_4481);
and U4915 (N_4915,N_3869,N_3642);
nor U4916 (N_4916,N_3379,N_4191);
xor U4917 (N_4917,N_4269,N_3725);
and U4918 (N_4918,N_4238,N_3349);
xnor U4919 (N_4919,N_4271,N_3010);
and U4920 (N_4920,N_3622,N_4176);
and U4921 (N_4921,N_3478,N_3529);
xnor U4922 (N_4922,N_3962,N_3017);
nor U4923 (N_4923,N_4301,N_3095);
and U4924 (N_4924,N_4160,N_3655);
or U4925 (N_4925,N_4082,N_3540);
xor U4926 (N_4926,N_4094,N_3479);
xnor U4927 (N_4927,N_3398,N_3467);
nand U4928 (N_4928,N_3917,N_3205);
or U4929 (N_4929,N_4181,N_3225);
xor U4930 (N_4930,N_3567,N_3483);
xnor U4931 (N_4931,N_3888,N_3691);
nand U4932 (N_4932,N_3674,N_4127);
xnor U4933 (N_4933,N_3656,N_3276);
nand U4934 (N_4934,N_4424,N_3633);
xnor U4935 (N_4935,N_4079,N_3855);
and U4936 (N_4936,N_3361,N_4443);
nand U4937 (N_4937,N_3799,N_3102);
xor U4938 (N_4938,N_4403,N_3062);
nand U4939 (N_4939,N_4151,N_3028);
and U4940 (N_4940,N_3368,N_3819);
and U4941 (N_4941,N_3054,N_3254);
nand U4942 (N_4942,N_4355,N_4021);
nand U4943 (N_4943,N_4143,N_4055);
nor U4944 (N_4944,N_3303,N_3201);
nand U4945 (N_4945,N_3716,N_3162);
and U4946 (N_4946,N_3321,N_3884);
or U4947 (N_4947,N_4187,N_4338);
and U4948 (N_4948,N_4379,N_3596);
and U4949 (N_4949,N_4234,N_3024);
nor U4950 (N_4950,N_4222,N_4027);
or U4951 (N_4951,N_3288,N_3685);
and U4952 (N_4952,N_4040,N_4085);
or U4953 (N_4953,N_3063,N_3743);
or U4954 (N_4954,N_4472,N_3169);
xor U4955 (N_4955,N_4284,N_4383);
or U4956 (N_4956,N_4247,N_3001);
nor U4957 (N_4957,N_4468,N_3227);
xor U4958 (N_4958,N_4182,N_3776);
or U4959 (N_4959,N_3954,N_3757);
and U4960 (N_4960,N_3299,N_3514);
xor U4961 (N_4961,N_3471,N_4385);
xnor U4962 (N_4962,N_3994,N_3258);
nand U4963 (N_4963,N_3239,N_3631);
nor U4964 (N_4964,N_3763,N_3027);
nor U4965 (N_4965,N_4389,N_3930);
and U4966 (N_4966,N_3381,N_4170);
nor U4967 (N_4967,N_3375,N_3310);
nor U4968 (N_4968,N_3901,N_4321);
nand U4969 (N_4969,N_3374,N_4076);
nor U4970 (N_4970,N_3919,N_3309);
nor U4971 (N_4971,N_4373,N_3610);
xnor U4972 (N_4972,N_4230,N_3082);
xor U4973 (N_4973,N_3537,N_3090);
and U4974 (N_4974,N_4430,N_3451);
xnor U4975 (N_4975,N_3098,N_4398);
and U4976 (N_4976,N_3528,N_4056);
nand U4977 (N_4977,N_3350,N_3412);
nand U4978 (N_4978,N_4376,N_4259);
and U4979 (N_4979,N_4198,N_4117);
and U4980 (N_4980,N_3800,N_3641);
and U4981 (N_4981,N_3164,N_3443);
nand U4982 (N_4982,N_4499,N_3115);
and U4983 (N_4983,N_3651,N_3069);
xnor U4984 (N_4984,N_3826,N_3207);
and U4985 (N_4985,N_4386,N_3597);
nor U4986 (N_4986,N_3414,N_3702);
xor U4987 (N_4987,N_4319,N_3654);
nor U4988 (N_4988,N_4363,N_3724);
nor U4989 (N_4989,N_4032,N_4067);
nand U4990 (N_4990,N_3871,N_4474);
nor U4991 (N_4991,N_3346,N_3747);
nor U4992 (N_4992,N_4483,N_3974);
xor U4993 (N_4993,N_4159,N_3625);
nand U4994 (N_4994,N_3265,N_4030);
or U4995 (N_4995,N_4007,N_3157);
nand U4996 (N_4996,N_3194,N_3180);
or U4997 (N_4997,N_3096,N_3422);
or U4998 (N_4998,N_3007,N_3882);
and U4999 (N_4999,N_3291,N_3766);
nand U5000 (N_5000,N_3798,N_3185);
or U5001 (N_5001,N_4343,N_4088);
xor U5002 (N_5002,N_3026,N_3081);
xor U5003 (N_5003,N_3515,N_3885);
or U5004 (N_5004,N_4164,N_3003);
nand U5005 (N_5005,N_4204,N_4166);
nor U5006 (N_5006,N_4268,N_3926);
nor U5007 (N_5007,N_3635,N_3985);
or U5008 (N_5008,N_3548,N_4282);
xnor U5009 (N_5009,N_3598,N_3131);
nor U5010 (N_5010,N_3921,N_4171);
nor U5011 (N_5011,N_4196,N_4401);
nand U5012 (N_5012,N_3163,N_3423);
or U5013 (N_5013,N_3009,N_3568);
xnor U5014 (N_5014,N_3142,N_4078);
nor U5015 (N_5015,N_3262,N_3019);
xor U5016 (N_5016,N_4002,N_3432);
or U5017 (N_5017,N_3448,N_4066);
xnor U5018 (N_5018,N_4193,N_3868);
xor U5019 (N_5019,N_3481,N_4445);
nand U5020 (N_5020,N_3679,N_3684);
xnor U5021 (N_5021,N_3059,N_3459);
and U5022 (N_5022,N_3823,N_4074);
or U5023 (N_5023,N_3578,N_4065);
xnor U5024 (N_5024,N_3734,N_3501);
nand U5025 (N_5025,N_3371,N_3079);
xor U5026 (N_5026,N_3883,N_3748);
xnor U5027 (N_5027,N_3354,N_3959);
nand U5028 (N_5028,N_4415,N_3267);
or U5029 (N_5029,N_4202,N_4186);
and U5030 (N_5030,N_4306,N_4392);
or U5031 (N_5031,N_3341,N_4116);
or U5032 (N_5032,N_3244,N_3681);
xor U5033 (N_5033,N_4486,N_4168);
and U5034 (N_5034,N_3908,N_3231);
and U5035 (N_5035,N_3342,N_4275);
nor U5036 (N_5036,N_3120,N_3365);
xor U5037 (N_5037,N_3692,N_3611);
xnor U5038 (N_5038,N_3040,N_3358);
nor U5039 (N_5039,N_3025,N_3475);
nor U5040 (N_5040,N_3476,N_3675);
and U5041 (N_5041,N_3595,N_4475);
or U5042 (N_5042,N_3972,N_3697);
xor U5043 (N_5043,N_3127,N_3176);
nor U5044 (N_5044,N_3895,N_3499);
xnor U5045 (N_5045,N_3923,N_4251);
and U5046 (N_5046,N_3626,N_3344);
nor U5047 (N_5047,N_4439,N_4081);
or U5048 (N_5048,N_4197,N_4437);
and U5049 (N_5049,N_3436,N_4153);
and U5050 (N_5050,N_4423,N_3388);
or U5051 (N_5051,N_3745,N_3992);
xnor U5052 (N_5052,N_4253,N_4254);
or U5053 (N_5053,N_3821,N_3732);
or U5054 (N_5054,N_3065,N_4077);
xor U5055 (N_5055,N_3825,N_3968);
nand U5056 (N_5056,N_3383,N_4296);
nor U5057 (N_5057,N_3837,N_3590);
xnor U5058 (N_5058,N_3454,N_4135);
or U5059 (N_5059,N_3075,N_4023);
and U5060 (N_5060,N_3196,N_3589);
nor U5061 (N_5061,N_3357,N_3332);
and U5062 (N_5062,N_4457,N_4326);
xnor U5063 (N_5063,N_4350,N_4184);
nand U5064 (N_5064,N_4420,N_4152);
xor U5065 (N_5065,N_3544,N_3049);
or U5066 (N_5066,N_3030,N_3698);
and U5067 (N_5067,N_3976,N_4039);
or U5068 (N_5068,N_4438,N_3343);
nand U5069 (N_5069,N_4224,N_4324);
nor U5070 (N_5070,N_4312,N_3717);
nand U5071 (N_5071,N_3689,N_4128);
nand U5072 (N_5072,N_3507,N_4410);
nand U5073 (N_5073,N_3445,N_3274);
and U5074 (N_5074,N_3940,N_3289);
and U5075 (N_5075,N_3646,N_3051);
xor U5076 (N_5076,N_3841,N_3839);
xor U5077 (N_5077,N_3991,N_3415);
xor U5078 (N_5078,N_3319,N_4351);
xnor U5079 (N_5079,N_3628,N_3768);
or U5080 (N_5080,N_3240,N_4013);
nand U5081 (N_5081,N_4174,N_3295);
and U5082 (N_5082,N_4308,N_4294);
or U5083 (N_5083,N_4051,N_4233);
nor U5084 (N_5084,N_3744,N_3023);
and U5085 (N_5085,N_3272,N_4092);
and U5086 (N_5086,N_3773,N_3929);
or U5087 (N_5087,N_4473,N_4459);
xnor U5088 (N_5088,N_3208,N_4026);
or U5089 (N_5089,N_3504,N_3833);
or U5090 (N_5090,N_4084,N_3452);
nand U5091 (N_5091,N_3352,N_4432);
or U5092 (N_5092,N_4278,N_4361);
nor U5093 (N_5093,N_3650,N_3512);
nor U5094 (N_5094,N_3618,N_3204);
and U5095 (N_5095,N_3181,N_3386);
xnor U5096 (N_5096,N_4292,N_3016);
nand U5097 (N_5097,N_4155,N_4161);
and U5098 (N_5098,N_4391,N_4494);
or U5099 (N_5099,N_3565,N_3444);
nand U5100 (N_5100,N_3585,N_3950);
or U5101 (N_5101,N_3469,N_3781);
xnor U5102 (N_5102,N_4495,N_3314);
or U5103 (N_5103,N_3878,N_4290);
xnor U5104 (N_5104,N_3466,N_3636);
xor U5105 (N_5105,N_3989,N_3006);
or U5106 (N_5106,N_3399,N_3300);
and U5107 (N_5107,N_3794,N_3803);
nor U5108 (N_5108,N_3939,N_3408);
nor U5109 (N_5109,N_3212,N_4471);
nor U5110 (N_5110,N_3502,N_3608);
nand U5111 (N_5111,N_4025,N_3845);
or U5112 (N_5112,N_3815,N_4348);
xnor U5113 (N_5113,N_3134,N_3516);
xor U5114 (N_5114,N_4444,N_4223);
and U5115 (N_5115,N_3931,N_3649);
nor U5116 (N_5116,N_4098,N_3526);
nor U5117 (N_5117,N_4462,N_4328);
xnor U5118 (N_5118,N_3490,N_3306);
nor U5119 (N_5119,N_4070,N_3084);
or U5120 (N_5120,N_4048,N_3477);
and U5121 (N_5121,N_4449,N_4303);
nand U5122 (N_5122,N_4393,N_4235);
nor U5123 (N_5123,N_4405,N_4246);
nand U5124 (N_5124,N_3284,N_4086);
or U5125 (N_5125,N_3791,N_3672);
or U5126 (N_5126,N_4138,N_3324);
xnor U5127 (N_5127,N_4095,N_3575);
nand U5128 (N_5128,N_3894,N_3876);
and U5129 (N_5129,N_3831,N_3195);
nor U5130 (N_5130,N_3167,N_4387);
nor U5131 (N_5131,N_3050,N_3536);
xor U5132 (N_5132,N_4185,N_4062);
xor U5133 (N_5133,N_3083,N_3660);
and U5134 (N_5134,N_3867,N_4329);
xnor U5135 (N_5135,N_3108,N_3579);
xnor U5136 (N_5136,N_4464,N_3246);
nor U5137 (N_5137,N_4371,N_4488);
or U5138 (N_5138,N_4054,N_3031);
and U5139 (N_5139,N_3453,N_3273);
nor U5140 (N_5140,N_3210,N_3582);
nand U5141 (N_5141,N_4429,N_3032);
nor U5142 (N_5142,N_3323,N_3146);
or U5143 (N_5143,N_3820,N_3816);
and U5144 (N_5144,N_3404,N_3510);
nor U5145 (N_5145,N_3488,N_3396);
nor U5146 (N_5146,N_4060,N_4244);
or U5147 (N_5147,N_4035,N_3232);
nand U5148 (N_5148,N_3735,N_3699);
or U5149 (N_5149,N_3543,N_3720);
nor U5150 (N_5150,N_3509,N_3709);
nor U5151 (N_5151,N_3788,N_3539);
and U5152 (N_5152,N_3761,N_3171);
and U5153 (N_5153,N_3914,N_3508);
and U5154 (N_5154,N_3327,N_3394);
and U5155 (N_5155,N_3072,N_4270);
nand U5156 (N_5156,N_4177,N_4286);
nand U5157 (N_5157,N_3238,N_3035);
nand U5158 (N_5158,N_3899,N_4057);
nor U5159 (N_5159,N_4404,N_3338);
nor U5160 (N_5160,N_3482,N_4448);
or U5161 (N_5161,N_4358,N_4375);
and U5162 (N_5162,N_3117,N_3409);
and U5163 (N_5163,N_3911,N_3630);
xnor U5164 (N_5164,N_3987,N_3154);
and U5165 (N_5165,N_4154,N_4090);
or U5166 (N_5166,N_3818,N_4402);
and U5167 (N_5167,N_3313,N_3202);
nor U5168 (N_5168,N_3377,N_3602);
nand U5169 (N_5169,N_3614,N_3380);
or U5170 (N_5170,N_3118,N_4399);
nand U5171 (N_5171,N_3263,N_3805);
xor U5172 (N_5172,N_3307,N_3401);
and U5173 (N_5173,N_3648,N_3260);
nand U5174 (N_5174,N_4307,N_3008);
nand U5175 (N_5175,N_3563,N_4265);
nand U5176 (N_5176,N_3229,N_3372);
nand U5177 (N_5177,N_3560,N_3902);
and U5178 (N_5178,N_3993,N_3896);
and U5179 (N_5179,N_3362,N_3178);
nor U5180 (N_5180,N_4272,N_3070);
or U5181 (N_5181,N_3538,N_4231);
or U5182 (N_5182,N_4454,N_3769);
nand U5183 (N_5183,N_4460,N_3221);
or U5184 (N_5184,N_3620,N_3583);
nand U5185 (N_5185,N_4467,N_3765);
xnor U5186 (N_5186,N_3200,N_4044);
nor U5187 (N_5187,N_3491,N_4011);
or U5188 (N_5188,N_3437,N_3828);
nand U5189 (N_5189,N_3148,N_4180);
xnor U5190 (N_5190,N_3873,N_3287);
and U5191 (N_5191,N_3858,N_3995);
xnor U5192 (N_5192,N_3495,N_3152);
nand U5193 (N_5193,N_4111,N_4036);
and U5194 (N_5194,N_3417,N_3844);
xor U5195 (N_5195,N_3465,N_3348);
and U5196 (N_5196,N_3910,N_3456);
and U5197 (N_5197,N_3983,N_3804);
xnor U5198 (N_5198,N_4136,N_3814);
nor U5199 (N_5199,N_3771,N_3809);
or U5200 (N_5200,N_4008,N_3235);
and U5201 (N_5201,N_4249,N_4179);
or U5202 (N_5202,N_3523,N_3320);
nand U5203 (N_5203,N_4416,N_3366);
or U5204 (N_5204,N_4221,N_3843);
and U5205 (N_5205,N_3158,N_3756);
xnor U5206 (N_5206,N_4134,N_3960);
nand U5207 (N_5207,N_3966,N_4047);
xor U5208 (N_5208,N_3886,N_3925);
and U5209 (N_5209,N_3041,N_4037);
xor U5210 (N_5210,N_4140,N_4108);
nor U5211 (N_5211,N_3556,N_4137);
nor U5212 (N_5212,N_3250,N_4175);
nand U5213 (N_5213,N_4414,N_3599);
nand U5214 (N_5214,N_3034,N_3718);
xor U5215 (N_5215,N_4122,N_3789);
xnor U5216 (N_5216,N_3677,N_3624);
nand U5217 (N_5217,N_4188,N_4318);
nor U5218 (N_5218,N_4440,N_4377);
and U5219 (N_5219,N_3727,N_4178);
nand U5220 (N_5220,N_3838,N_3237);
nor U5221 (N_5221,N_3337,N_4214);
nand U5222 (N_5222,N_3064,N_4340);
nor U5223 (N_5223,N_3166,N_3854);
xnor U5224 (N_5224,N_3889,N_4237);
and U5225 (N_5225,N_4480,N_3591);
and U5226 (N_5226,N_4118,N_3213);
and U5227 (N_5227,N_4434,N_4105);
nand U5228 (N_5228,N_4316,N_3042);
xor U5229 (N_5229,N_3750,N_4339);
or U5230 (N_5230,N_3468,N_4089);
nor U5231 (N_5231,N_4332,N_4147);
xnor U5232 (N_5232,N_4046,N_3014);
xnor U5233 (N_5233,N_3384,N_3331);
or U5234 (N_5234,N_4336,N_3978);
xnor U5235 (N_5235,N_3177,N_4425);
nor U5236 (N_5236,N_4470,N_3316);
and U5237 (N_5237,N_4407,N_3433);
xor U5238 (N_5238,N_4266,N_3071);
nor U5239 (N_5239,N_3197,N_3676);
or U5240 (N_5240,N_3385,N_3073);
or U5241 (N_5241,N_3187,N_4130);
nand U5242 (N_5242,N_3170,N_3812);
or U5243 (N_5243,N_3500,N_3053);
nor U5244 (N_5244,N_3918,N_3226);
nand U5245 (N_5245,N_3045,N_3145);
xnor U5246 (N_5246,N_4357,N_3863);
nand U5247 (N_5247,N_4162,N_4146);
nor U5248 (N_5248,N_3304,N_3552);
nor U5249 (N_5249,N_4103,N_4267);
or U5250 (N_5250,N_3759,N_3849);
nand U5251 (N_5251,N_4126,N_3246);
nand U5252 (N_5252,N_3645,N_3642);
nand U5253 (N_5253,N_3764,N_3827);
xnor U5254 (N_5254,N_3165,N_4077);
and U5255 (N_5255,N_3624,N_4269);
xor U5256 (N_5256,N_4080,N_3644);
nand U5257 (N_5257,N_3270,N_3996);
or U5258 (N_5258,N_4201,N_3135);
and U5259 (N_5259,N_3035,N_3130);
or U5260 (N_5260,N_4142,N_3663);
and U5261 (N_5261,N_3666,N_3051);
xnor U5262 (N_5262,N_3923,N_3273);
nor U5263 (N_5263,N_3730,N_3388);
nand U5264 (N_5264,N_3889,N_3961);
nor U5265 (N_5265,N_3499,N_4341);
xor U5266 (N_5266,N_4496,N_4100);
and U5267 (N_5267,N_3167,N_3201);
and U5268 (N_5268,N_4014,N_4074);
or U5269 (N_5269,N_3093,N_4431);
nor U5270 (N_5270,N_3346,N_4316);
nand U5271 (N_5271,N_4148,N_3385);
and U5272 (N_5272,N_3173,N_3427);
nand U5273 (N_5273,N_4220,N_3892);
xor U5274 (N_5274,N_3699,N_3616);
nor U5275 (N_5275,N_4021,N_4198);
and U5276 (N_5276,N_3535,N_3805);
or U5277 (N_5277,N_3666,N_3431);
and U5278 (N_5278,N_4347,N_4339);
xnor U5279 (N_5279,N_3591,N_3813);
and U5280 (N_5280,N_3146,N_4114);
or U5281 (N_5281,N_3407,N_4461);
or U5282 (N_5282,N_3784,N_3810);
nor U5283 (N_5283,N_3327,N_3199);
nor U5284 (N_5284,N_3079,N_4142);
nor U5285 (N_5285,N_3489,N_3483);
nor U5286 (N_5286,N_4113,N_3514);
xor U5287 (N_5287,N_3463,N_3933);
nand U5288 (N_5288,N_3011,N_4167);
or U5289 (N_5289,N_3386,N_4448);
nand U5290 (N_5290,N_3519,N_3119);
nand U5291 (N_5291,N_3845,N_4285);
xnor U5292 (N_5292,N_3413,N_3928);
nand U5293 (N_5293,N_3159,N_3074);
nor U5294 (N_5294,N_4396,N_3679);
nand U5295 (N_5295,N_4439,N_3070);
and U5296 (N_5296,N_4123,N_3683);
and U5297 (N_5297,N_3451,N_4334);
or U5298 (N_5298,N_3085,N_3441);
nand U5299 (N_5299,N_3927,N_3764);
and U5300 (N_5300,N_4204,N_4104);
nand U5301 (N_5301,N_3391,N_3486);
and U5302 (N_5302,N_3735,N_4336);
and U5303 (N_5303,N_4323,N_4101);
nor U5304 (N_5304,N_3229,N_3224);
nand U5305 (N_5305,N_3937,N_3217);
nor U5306 (N_5306,N_3680,N_3118);
nand U5307 (N_5307,N_3394,N_3550);
nor U5308 (N_5308,N_3252,N_4436);
xnor U5309 (N_5309,N_3353,N_4064);
nor U5310 (N_5310,N_3040,N_4307);
nand U5311 (N_5311,N_4284,N_3351);
and U5312 (N_5312,N_3250,N_3334);
or U5313 (N_5313,N_3355,N_3302);
or U5314 (N_5314,N_3357,N_3921);
or U5315 (N_5315,N_3755,N_4173);
nor U5316 (N_5316,N_3559,N_3128);
and U5317 (N_5317,N_3626,N_3255);
nor U5318 (N_5318,N_3681,N_4342);
nor U5319 (N_5319,N_3736,N_3067);
nand U5320 (N_5320,N_3644,N_4070);
or U5321 (N_5321,N_3584,N_4078);
nand U5322 (N_5322,N_3106,N_4397);
nand U5323 (N_5323,N_3537,N_3405);
nand U5324 (N_5324,N_4108,N_4190);
nand U5325 (N_5325,N_4151,N_4394);
nand U5326 (N_5326,N_3877,N_3471);
nor U5327 (N_5327,N_3730,N_3621);
nand U5328 (N_5328,N_3876,N_3809);
xor U5329 (N_5329,N_3193,N_3860);
nor U5330 (N_5330,N_3004,N_3779);
xor U5331 (N_5331,N_4496,N_3776);
nand U5332 (N_5332,N_4471,N_3805);
or U5333 (N_5333,N_3840,N_4085);
nand U5334 (N_5334,N_3141,N_3267);
xor U5335 (N_5335,N_3362,N_3599);
or U5336 (N_5336,N_3216,N_4348);
nor U5337 (N_5337,N_3258,N_4404);
and U5338 (N_5338,N_3063,N_3068);
or U5339 (N_5339,N_3311,N_4181);
and U5340 (N_5340,N_4007,N_4152);
or U5341 (N_5341,N_3612,N_4016);
nand U5342 (N_5342,N_4174,N_3227);
nor U5343 (N_5343,N_3867,N_4392);
xor U5344 (N_5344,N_3399,N_4471);
nor U5345 (N_5345,N_4312,N_3481);
xor U5346 (N_5346,N_3722,N_4186);
or U5347 (N_5347,N_3216,N_3233);
nor U5348 (N_5348,N_4456,N_3515);
nor U5349 (N_5349,N_4118,N_3203);
xor U5350 (N_5350,N_3994,N_3693);
or U5351 (N_5351,N_3668,N_4270);
nand U5352 (N_5352,N_3457,N_3340);
and U5353 (N_5353,N_3608,N_3970);
nand U5354 (N_5354,N_3163,N_4039);
or U5355 (N_5355,N_4391,N_4272);
nand U5356 (N_5356,N_3428,N_3747);
nand U5357 (N_5357,N_3547,N_3507);
nand U5358 (N_5358,N_4011,N_4119);
xor U5359 (N_5359,N_3045,N_3252);
nor U5360 (N_5360,N_3716,N_3118);
nand U5361 (N_5361,N_3737,N_3117);
nor U5362 (N_5362,N_4134,N_4286);
nand U5363 (N_5363,N_4256,N_3887);
xnor U5364 (N_5364,N_3162,N_3047);
nor U5365 (N_5365,N_4124,N_3097);
nand U5366 (N_5366,N_4321,N_3462);
nor U5367 (N_5367,N_3352,N_4443);
nand U5368 (N_5368,N_3489,N_4325);
and U5369 (N_5369,N_3003,N_3801);
and U5370 (N_5370,N_4283,N_3030);
nor U5371 (N_5371,N_3802,N_4288);
xor U5372 (N_5372,N_4372,N_3007);
nor U5373 (N_5373,N_4270,N_3020);
and U5374 (N_5374,N_3584,N_3757);
and U5375 (N_5375,N_3312,N_4176);
xor U5376 (N_5376,N_4280,N_4358);
or U5377 (N_5377,N_3960,N_3732);
nor U5378 (N_5378,N_4409,N_4007);
xor U5379 (N_5379,N_3246,N_3649);
or U5380 (N_5380,N_3684,N_4299);
and U5381 (N_5381,N_4053,N_3718);
xor U5382 (N_5382,N_3072,N_4087);
and U5383 (N_5383,N_4082,N_3978);
nand U5384 (N_5384,N_3342,N_4089);
nor U5385 (N_5385,N_3680,N_3679);
or U5386 (N_5386,N_3035,N_4169);
nand U5387 (N_5387,N_3674,N_4325);
or U5388 (N_5388,N_3792,N_3700);
xnor U5389 (N_5389,N_3408,N_3536);
xor U5390 (N_5390,N_3506,N_3628);
and U5391 (N_5391,N_4289,N_3694);
or U5392 (N_5392,N_3977,N_3583);
xor U5393 (N_5393,N_4468,N_3113);
nor U5394 (N_5394,N_4095,N_3791);
and U5395 (N_5395,N_3552,N_3094);
nand U5396 (N_5396,N_4413,N_3549);
nand U5397 (N_5397,N_3274,N_3119);
or U5398 (N_5398,N_3495,N_3215);
nor U5399 (N_5399,N_3780,N_4436);
xnor U5400 (N_5400,N_3922,N_4419);
and U5401 (N_5401,N_3940,N_4290);
nand U5402 (N_5402,N_3864,N_4090);
and U5403 (N_5403,N_3174,N_4007);
and U5404 (N_5404,N_4128,N_3617);
nor U5405 (N_5405,N_3633,N_4493);
nand U5406 (N_5406,N_3321,N_3291);
nand U5407 (N_5407,N_3208,N_3390);
and U5408 (N_5408,N_4187,N_3869);
or U5409 (N_5409,N_4253,N_3569);
xor U5410 (N_5410,N_4193,N_3338);
xor U5411 (N_5411,N_4360,N_3634);
nand U5412 (N_5412,N_4371,N_3555);
nand U5413 (N_5413,N_3419,N_4230);
or U5414 (N_5414,N_3766,N_3474);
or U5415 (N_5415,N_3301,N_3082);
and U5416 (N_5416,N_3719,N_3126);
nand U5417 (N_5417,N_3549,N_4298);
and U5418 (N_5418,N_3025,N_3951);
xnor U5419 (N_5419,N_3064,N_4119);
nor U5420 (N_5420,N_3509,N_3851);
xnor U5421 (N_5421,N_3515,N_3112);
and U5422 (N_5422,N_3023,N_3891);
or U5423 (N_5423,N_3921,N_3865);
or U5424 (N_5424,N_3873,N_3116);
xor U5425 (N_5425,N_3331,N_4338);
nor U5426 (N_5426,N_3218,N_4401);
or U5427 (N_5427,N_4154,N_3218);
nor U5428 (N_5428,N_3844,N_4199);
nand U5429 (N_5429,N_3474,N_3880);
or U5430 (N_5430,N_4412,N_4072);
nor U5431 (N_5431,N_4242,N_4034);
and U5432 (N_5432,N_3170,N_3512);
nand U5433 (N_5433,N_3369,N_3844);
nand U5434 (N_5434,N_3101,N_4477);
xor U5435 (N_5435,N_3353,N_3613);
nand U5436 (N_5436,N_3793,N_4096);
xnor U5437 (N_5437,N_3799,N_3720);
or U5438 (N_5438,N_3690,N_3676);
nand U5439 (N_5439,N_4111,N_3383);
xnor U5440 (N_5440,N_3472,N_4068);
or U5441 (N_5441,N_3060,N_3490);
or U5442 (N_5442,N_3534,N_4247);
and U5443 (N_5443,N_4397,N_3053);
or U5444 (N_5444,N_4158,N_3812);
nand U5445 (N_5445,N_3367,N_3570);
nand U5446 (N_5446,N_3847,N_4315);
or U5447 (N_5447,N_4495,N_4281);
or U5448 (N_5448,N_3790,N_4443);
xnor U5449 (N_5449,N_3729,N_3222);
nand U5450 (N_5450,N_3387,N_4489);
nor U5451 (N_5451,N_3158,N_3265);
nand U5452 (N_5452,N_3849,N_4430);
nand U5453 (N_5453,N_3275,N_3989);
nand U5454 (N_5454,N_3906,N_3466);
and U5455 (N_5455,N_3519,N_3922);
xor U5456 (N_5456,N_4235,N_4119);
and U5457 (N_5457,N_4157,N_4109);
or U5458 (N_5458,N_3385,N_4228);
nand U5459 (N_5459,N_3336,N_3698);
xnor U5460 (N_5460,N_4344,N_4202);
nand U5461 (N_5461,N_3791,N_3418);
or U5462 (N_5462,N_3732,N_3375);
nor U5463 (N_5463,N_3884,N_4348);
or U5464 (N_5464,N_3280,N_3682);
nor U5465 (N_5465,N_4495,N_3263);
and U5466 (N_5466,N_3509,N_3485);
and U5467 (N_5467,N_4389,N_3511);
or U5468 (N_5468,N_3372,N_3516);
xor U5469 (N_5469,N_4421,N_3811);
nor U5470 (N_5470,N_3736,N_3284);
xnor U5471 (N_5471,N_3242,N_3988);
nand U5472 (N_5472,N_3201,N_3760);
nand U5473 (N_5473,N_3066,N_3325);
or U5474 (N_5474,N_3917,N_3345);
nand U5475 (N_5475,N_3255,N_4123);
xnor U5476 (N_5476,N_4261,N_3454);
nand U5477 (N_5477,N_3634,N_3147);
and U5478 (N_5478,N_4172,N_4070);
and U5479 (N_5479,N_3141,N_4087);
nor U5480 (N_5480,N_4099,N_3618);
or U5481 (N_5481,N_3625,N_3600);
or U5482 (N_5482,N_4430,N_3591);
and U5483 (N_5483,N_3474,N_3773);
nor U5484 (N_5484,N_3172,N_3013);
and U5485 (N_5485,N_3059,N_3554);
nor U5486 (N_5486,N_3795,N_4070);
nand U5487 (N_5487,N_3475,N_4207);
nor U5488 (N_5488,N_3776,N_4462);
and U5489 (N_5489,N_3101,N_4234);
or U5490 (N_5490,N_4343,N_4129);
or U5491 (N_5491,N_3492,N_4087);
nand U5492 (N_5492,N_3452,N_4270);
or U5493 (N_5493,N_3620,N_4448);
nand U5494 (N_5494,N_4417,N_3218);
nor U5495 (N_5495,N_3235,N_3688);
and U5496 (N_5496,N_4450,N_4045);
nand U5497 (N_5497,N_4134,N_3607);
nand U5498 (N_5498,N_4252,N_3904);
or U5499 (N_5499,N_3551,N_3023);
nor U5500 (N_5500,N_3514,N_3985);
nor U5501 (N_5501,N_3328,N_3727);
nor U5502 (N_5502,N_3945,N_4413);
nand U5503 (N_5503,N_3974,N_3765);
or U5504 (N_5504,N_3166,N_4359);
nand U5505 (N_5505,N_4175,N_3087);
nand U5506 (N_5506,N_3279,N_4312);
xor U5507 (N_5507,N_3092,N_3011);
nand U5508 (N_5508,N_3223,N_3803);
and U5509 (N_5509,N_3884,N_4258);
xnor U5510 (N_5510,N_4455,N_4006);
nand U5511 (N_5511,N_3678,N_3823);
xor U5512 (N_5512,N_3528,N_3343);
and U5513 (N_5513,N_4180,N_3144);
and U5514 (N_5514,N_3465,N_4403);
nor U5515 (N_5515,N_4138,N_3943);
xor U5516 (N_5516,N_3049,N_4331);
nor U5517 (N_5517,N_4477,N_4294);
xnor U5518 (N_5518,N_3892,N_3562);
nand U5519 (N_5519,N_3081,N_4200);
or U5520 (N_5520,N_3889,N_3096);
and U5521 (N_5521,N_4291,N_3706);
xor U5522 (N_5522,N_4241,N_3777);
nand U5523 (N_5523,N_4277,N_4228);
and U5524 (N_5524,N_3131,N_3792);
or U5525 (N_5525,N_3570,N_3196);
or U5526 (N_5526,N_4054,N_3929);
nor U5527 (N_5527,N_3804,N_3295);
and U5528 (N_5528,N_4176,N_4159);
and U5529 (N_5529,N_3951,N_3707);
nor U5530 (N_5530,N_3052,N_4044);
and U5531 (N_5531,N_3245,N_3107);
and U5532 (N_5532,N_4239,N_3445);
xor U5533 (N_5533,N_3830,N_3438);
xnor U5534 (N_5534,N_4144,N_3615);
or U5535 (N_5535,N_3714,N_3170);
nor U5536 (N_5536,N_3964,N_4351);
nor U5537 (N_5537,N_3368,N_3634);
nand U5538 (N_5538,N_3174,N_4178);
nor U5539 (N_5539,N_3689,N_3680);
nor U5540 (N_5540,N_3432,N_3354);
or U5541 (N_5541,N_3421,N_4032);
nor U5542 (N_5542,N_4199,N_4478);
and U5543 (N_5543,N_4022,N_3447);
or U5544 (N_5544,N_4188,N_3277);
nand U5545 (N_5545,N_3546,N_3786);
nor U5546 (N_5546,N_3344,N_3163);
xor U5547 (N_5547,N_3018,N_4312);
or U5548 (N_5548,N_3180,N_3868);
xnor U5549 (N_5549,N_4361,N_3357);
and U5550 (N_5550,N_3349,N_3622);
xnor U5551 (N_5551,N_3081,N_3804);
nor U5552 (N_5552,N_3457,N_3534);
or U5553 (N_5553,N_3709,N_4433);
nor U5554 (N_5554,N_4258,N_3374);
nand U5555 (N_5555,N_4452,N_3396);
and U5556 (N_5556,N_4234,N_4439);
or U5557 (N_5557,N_4189,N_4241);
xor U5558 (N_5558,N_3341,N_3542);
xnor U5559 (N_5559,N_4193,N_3167);
and U5560 (N_5560,N_4382,N_3287);
and U5561 (N_5561,N_4079,N_4246);
xnor U5562 (N_5562,N_3547,N_3294);
nand U5563 (N_5563,N_3657,N_4461);
nand U5564 (N_5564,N_3368,N_3728);
and U5565 (N_5565,N_4453,N_3978);
or U5566 (N_5566,N_3665,N_3404);
or U5567 (N_5567,N_3155,N_4475);
xnor U5568 (N_5568,N_3971,N_3974);
or U5569 (N_5569,N_3208,N_3542);
nand U5570 (N_5570,N_3459,N_4026);
and U5571 (N_5571,N_3407,N_4329);
or U5572 (N_5572,N_3587,N_4169);
and U5573 (N_5573,N_4415,N_4366);
and U5574 (N_5574,N_3242,N_3860);
or U5575 (N_5575,N_3894,N_3400);
nand U5576 (N_5576,N_3205,N_3703);
and U5577 (N_5577,N_4107,N_4146);
xor U5578 (N_5578,N_3662,N_3007);
or U5579 (N_5579,N_3191,N_3172);
xnor U5580 (N_5580,N_3981,N_4083);
nor U5581 (N_5581,N_4048,N_3925);
and U5582 (N_5582,N_3215,N_3249);
xor U5583 (N_5583,N_4311,N_3146);
and U5584 (N_5584,N_4061,N_3777);
xnor U5585 (N_5585,N_4189,N_3336);
nand U5586 (N_5586,N_4168,N_4318);
and U5587 (N_5587,N_3991,N_3172);
and U5588 (N_5588,N_3206,N_3350);
nor U5589 (N_5589,N_3655,N_3280);
or U5590 (N_5590,N_4409,N_4422);
nor U5591 (N_5591,N_3997,N_3690);
and U5592 (N_5592,N_3154,N_3767);
and U5593 (N_5593,N_3113,N_3407);
xor U5594 (N_5594,N_3195,N_4449);
nor U5595 (N_5595,N_3446,N_3909);
nand U5596 (N_5596,N_3681,N_3173);
or U5597 (N_5597,N_3866,N_3713);
and U5598 (N_5598,N_4363,N_4333);
xnor U5599 (N_5599,N_4336,N_4032);
nor U5600 (N_5600,N_3162,N_4033);
and U5601 (N_5601,N_4115,N_3279);
xnor U5602 (N_5602,N_3132,N_3809);
xnor U5603 (N_5603,N_4471,N_3373);
or U5604 (N_5604,N_3554,N_3781);
xnor U5605 (N_5605,N_4423,N_4019);
nand U5606 (N_5606,N_3069,N_4068);
and U5607 (N_5607,N_3503,N_3162);
xor U5608 (N_5608,N_4086,N_4297);
nor U5609 (N_5609,N_4310,N_3091);
nand U5610 (N_5610,N_4459,N_4155);
nor U5611 (N_5611,N_3256,N_3812);
nand U5612 (N_5612,N_3746,N_3581);
nand U5613 (N_5613,N_3307,N_4179);
or U5614 (N_5614,N_3703,N_4421);
nand U5615 (N_5615,N_3832,N_3801);
or U5616 (N_5616,N_3866,N_3799);
or U5617 (N_5617,N_3632,N_3691);
nor U5618 (N_5618,N_3017,N_4152);
or U5619 (N_5619,N_3005,N_4083);
xor U5620 (N_5620,N_3475,N_3155);
xnor U5621 (N_5621,N_3712,N_4395);
or U5622 (N_5622,N_3462,N_3602);
or U5623 (N_5623,N_4271,N_3668);
and U5624 (N_5624,N_3779,N_3241);
xnor U5625 (N_5625,N_4002,N_3650);
xnor U5626 (N_5626,N_3346,N_4461);
and U5627 (N_5627,N_3215,N_4411);
or U5628 (N_5628,N_3374,N_4084);
or U5629 (N_5629,N_3607,N_3219);
xnor U5630 (N_5630,N_4053,N_3668);
nand U5631 (N_5631,N_4335,N_3448);
and U5632 (N_5632,N_3364,N_3239);
nand U5633 (N_5633,N_3517,N_3795);
and U5634 (N_5634,N_4323,N_3660);
and U5635 (N_5635,N_3692,N_4079);
nor U5636 (N_5636,N_4057,N_3173);
xnor U5637 (N_5637,N_3995,N_3126);
xor U5638 (N_5638,N_4362,N_3693);
xnor U5639 (N_5639,N_3717,N_3850);
xnor U5640 (N_5640,N_4045,N_3329);
nor U5641 (N_5641,N_3522,N_3339);
xor U5642 (N_5642,N_3879,N_3261);
nand U5643 (N_5643,N_4306,N_3076);
xnor U5644 (N_5644,N_3581,N_3651);
nand U5645 (N_5645,N_4462,N_3398);
nor U5646 (N_5646,N_3031,N_3361);
nand U5647 (N_5647,N_4169,N_4037);
or U5648 (N_5648,N_4011,N_3378);
and U5649 (N_5649,N_4399,N_3058);
xor U5650 (N_5650,N_3346,N_3189);
xnor U5651 (N_5651,N_3463,N_3160);
nor U5652 (N_5652,N_3826,N_3383);
xnor U5653 (N_5653,N_4100,N_3413);
or U5654 (N_5654,N_3693,N_4001);
xor U5655 (N_5655,N_3012,N_4172);
nor U5656 (N_5656,N_3673,N_3179);
or U5657 (N_5657,N_4128,N_3790);
and U5658 (N_5658,N_4464,N_3466);
nor U5659 (N_5659,N_3810,N_4127);
xor U5660 (N_5660,N_4269,N_3412);
or U5661 (N_5661,N_3077,N_4469);
and U5662 (N_5662,N_4344,N_4482);
xor U5663 (N_5663,N_3467,N_4461);
and U5664 (N_5664,N_4087,N_4377);
nor U5665 (N_5665,N_4043,N_4285);
xor U5666 (N_5666,N_3079,N_4102);
and U5667 (N_5667,N_4415,N_4088);
and U5668 (N_5668,N_3933,N_4426);
or U5669 (N_5669,N_3043,N_4360);
or U5670 (N_5670,N_3233,N_3989);
nand U5671 (N_5671,N_4341,N_3304);
xor U5672 (N_5672,N_3115,N_3058);
or U5673 (N_5673,N_3282,N_4230);
nor U5674 (N_5674,N_3953,N_3192);
xor U5675 (N_5675,N_4487,N_4371);
and U5676 (N_5676,N_3680,N_3293);
and U5677 (N_5677,N_3279,N_4126);
nand U5678 (N_5678,N_4210,N_3290);
xnor U5679 (N_5679,N_3243,N_3692);
or U5680 (N_5680,N_4362,N_3034);
or U5681 (N_5681,N_3613,N_4438);
xnor U5682 (N_5682,N_3745,N_3846);
nor U5683 (N_5683,N_3270,N_3345);
xor U5684 (N_5684,N_3319,N_4392);
nand U5685 (N_5685,N_3937,N_4015);
or U5686 (N_5686,N_4376,N_4193);
nor U5687 (N_5687,N_3828,N_4331);
nand U5688 (N_5688,N_3783,N_3626);
and U5689 (N_5689,N_3580,N_4121);
nand U5690 (N_5690,N_3131,N_3886);
or U5691 (N_5691,N_3488,N_3649);
and U5692 (N_5692,N_3060,N_3524);
nand U5693 (N_5693,N_3644,N_3221);
xor U5694 (N_5694,N_3234,N_3985);
xor U5695 (N_5695,N_3726,N_3789);
or U5696 (N_5696,N_3518,N_4277);
nor U5697 (N_5697,N_3146,N_3529);
and U5698 (N_5698,N_3248,N_3856);
nand U5699 (N_5699,N_3308,N_4248);
nor U5700 (N_5700,N_3121,N_3677);
nand U5701 (N_5701,N_4152,N_3528);
nand U5702 (N_5702,N_3173,N_3622);
xor U5703 (N_5703,N_3276,N_3797);
nor U5704 (N_5704,N_3134,N_4023);
nand U5705 (N_5705,N_3497,N_3030);
xnor U5706 (N_5706,N_3485,N_3743);
or U5707 (N_5707,N_3176,N_4041);
nor U5708 (N_5708,N_4167,N_3251);
nand U5709 (N_5709,N_3150,N_3887);
nor U5710 (N_5710,N_3856,N_3397);
nor U5711 (N_5711,N_4192,N_3217);
nand U5712 (N_5712,N_4005,N_4135);
nor U5713 (N_5713,N_4256,N_4228);
nand U5714 (N_5714,N_3394,N_4332);
and U5715 (N_5715,N_3644,N_4467);
nor U5716 (N_5716,N_3601,N_4471);
or U5717 (N_5717,N_3135,N_3588);
or U5718 (N_5718,N_3448,N_3224);
and U5719 (N_5719,N_3227,N_3614);
xnor U5720 (N_5720,N_4226,N_4312);
and U5721 (N_5721,N_4038,N_3350);
xor U5722 (N_5722,N_3905,N_3501);
or U5723 (N_5723,N_3945,N_4287);
xor U5724 (N_5724,N_3301,N_4357);
and U5725 (N_5725,N_3338,N_4197);
and U5726 (N_5726,N_4215,N_3940);
and U5727 (N_5727,N_3298,N_4096);
nor U5728 (N_5728,N_3592,N_3258);
and U5729 (N_5729,N_4312,N_4164);
nor U5730 (N_5730,N_3766,N_3425);
or U5731 (N_5731,N_3049,N_3484);
and U5732 (N_5732,N_3246,N_4147);
nand U5733 (N_5733,N_4232,N_3948);
or U5734 (N_5734,N_4263,N_3609);
nor U5735 (N_5735,N_4288,N_3096);
xnor U5736 (N_5736,N_3560,N_4002);
and U5737 (N_5737,N_3189,N_3432);
nand U5738 (N_5738,N_3508,N_3421);
xnor U5739 (N_5739,N_4376,N_3896);
xor U5740 (N_5740,N_3543,N_4488);
or U5741 (N_5741,N_3972,N_3631);
nor U5742 (N_5742,N_3446,N_3224);
or U5743 (N_5743,N_3633,N_3925);
or U5744 (N_5744,N_4285,N_4044);
or U5745 (N_5745,N_4293,N_3340);
nor U5746 (N_5746,N_3327,N_3098);
nor U5747 (N_5747,N_4415,N_3287);
nor U5748 (N_5748,N_4483,N_3712);
xor U5749 (N_5749,N_3921,N_4028);
nand U5750 (N_5750,N_4303,N_3078);
nand U5751 (N_5751,N_3054,N_3972);
nor U5752 (N_5752,N_3589,N_3018);
nand U5753 (N_5753,N_4111,N_3447);
xor U5754 (N_5754,N_3865,N_3112);
nor U5755 (N_5755,N_4283,N_3993);
or U5756 (N_5756,N_3130,N_3216);
and U5757 (N_5757,N_3783,N_4036);
xor U5758 (N_5758,N_3500,N_4095);
xor U5759 (N_5759,N_3582,N_4120);
or U5760 (N_5760,N_3486,N_4153);
nor U5761 (N_5761,N_4458,N_3110);
xnor U5762 (N_5762,N_3176,N_4442);
and U5763 (N_5763,N_4489,N_3875);
and U5764 (N_5764,N_3367,N_3402);
and U5765 (N_5765,N_3485,N_3177);
or U5766 (N_5766,N_3437,N_3992);
and U5767 (N_5767,N_4336,N_3452);
xor U5768 (N_5768,N_4092,N_3315);
xor U5769 (N_5769,N_3029,N_3637);
and U5770 (N_5770,N_3872,N_4153);
nand U5771 (N_5771,N_3438,N_3746);
xor U5772 (N_5772,N_3170,N_4415);
nand U5773 (N_5773,N_3320,N_4443);
nor U5774 (N_5774,N_3477,N_3262);
nor U5775 (N_5775,N_3100,N_4081);
xor U5776 (N_5776,N_4228,N_3304);
nand U5777 (N_5777,N_3502,N_4366);
xor U5778 (N_5778,N_3959,N_3777);
xnor U5779 (N_5779,N_3598,N_3836);
xor U5780 (N_5780,N_3470,N_4114);
nand U5781 (N_5781,N_3016,N_3680);
or U5782 (N_5782,N_3046,N_4204);
nor U5783 (N_5783,N_3012,N_4190);
or U5784 (N_5784,N_3732,N_4398);
nand U5785 (N_5785,N_3787,N_4222);
xnor U5786 (N_5786,N_3022,N_3223);
or U5787 (N_5787,N_3325,N_4389);
xnor U5788 (N_5788,N_3930,N_3214);
nor U5789 (N_5789,N_4068,N_4129);
and U5790 (N_5790,N_4420,N_4296);
nor U5791 (N_5791,N_3180,N_3338);
and U5792 (N_5792,N_4240,N_4392);
and U5793 (N_5793,N_3356,N_3728);
nand U5794 (N_5794,N_3072,N_4350);
or U5795 (N_5795,N_3707,N_3469);
nand U5796 (N_5796,N_3535,N_3352);
nor U5797 (N_5797,N_4105,N_3478);
or U5798 (N_5798,N_4204,N_3477);
or U5799 (N_5799,N_3282,N_4334);
nand U5800 (N_5800,N_3015,N_3480);
nor U5801 (N_5801,N_4499,N_4467);
nand U5802 (N_5802,N_3722,N_3582);
or U5803 (N_5803,N_3550,N_3131);
nor U5804 (N_5804,N_3165,N_3670);
and U5805 (N_5805,N_4387,N_3200);
xor U5806 (N_5806,N_4457,N_4274);
xor U5807 (N_5807,N_3137,N_3088);
nand U5808 (N_5808,N_3475,N_3893);
xnor U5809 (N_5809,N_4330,N_3676);
xnor U5810 (N_5810,N_4249,N_3922);
and U5811 (N_5811,N_3173,N_3761);
nand U5812 (N_5812,N_3872,N_3803);
nand U5813 (N_5813,N_3539,N_4436);
or U5814 (N_5814,N_4425,N_4102);
nand U5815 (N_5815,N_3201,N_4450);
xnor U5816 (N_5816,N_4011,N_3504);
nor U5817 (N_5817,N_3516,N_3169);
nor U5818 (N_5818,N_4422,N_4433);
or U5819 (N_5819,N_3292,N_4046);
nor U5820 (N_5820,N_3258,N_3543);
and U5821 (N_5821,N_3569,N_4341);
xnor U5822 (N_5822,N_4161,N_4253);
nor U5823 (N_5823,N_3906,N_3185);
xor U5824 (N_5824,N_3596,N_3626);
or U5825 (N_5825,N_3882,N_3795);
or U5826 (N_5826,N_4271,N_4093);
and U5827 (N_5827,N_4380,N_3349);
nor U5828 (N_5828,N_3896,N_4143);
and U5829 (N_5829,N_4250,N_3238);
or U5830 (N_5830,N_3832,N_3776);
or U5831 (N_5831,N_3648,N_3834);
or U5832 (N_5832,N_3053,N_3998);
nand U5833 (N_5833,N_3940,N_3182);
or U5834 (N_5834,N_3380,N_4098);
xnor U5835 (N_5835,N_3471,N_4446);
nand U5836 (N_5836,N_4413,N_3268);
nand U5837 (N_5837,N_3728,N_3464);
and U5838 (N_5838,N_3203,N_3556);
and U5839 (N_5839,N_3899,N_3046);
nor U5840 (N_5840,N_3100,N_4295);
nand U5841 (N_5841,N_3508,N_4461);
and U5842 (N_5842,N_3020,N_4400);
nand U5843 (N_5843,N_4174,N_3501);
xnor U5844 (N_5844,N_3427,N_3250);
and U5845 (N_5845,N_3530,N_4283);
and U5846 (N_5846,N_4115,N_4272);
nor U5847 (N_5847,N_4270,N_3482);
nand U5848 (N_5848,N_3667,N_4182);
nand U5849 (N_5849,N_3203,N_3348);
nand U5850 (N_5850,N_3600,N_4282);
xor U5851 (N_5851,N_4211,N_4364);
nor U5852 (N_5852,N_3324,N_3414);
nor U5853 (N_5853,N_3325,N_3123);
nand U5854 (N_5854,N_3632,N_3192);
or U5855 (N_5855,N_3586,N_3802);
nand U5856 (N_5856,N_4257,N_3317);
nor U5857 (N_5857,N_3650,N_4342);
nand U5858 (N_5858,N_4328,N_4313);
or U5859 (N_5859,N_4278,N_3564);
nand U5860 (N_5860,N_3903,N_4311);
and U5861 (N_5861,N_4053,N_3251);
nor U5862 (N_5862,N_4489,N_3008);
or U5863 (N_5863,N_3259,N_3524);
xnor U5864 (N_5864,N_3430,N_3499);
nand U5865 (N_5865,N_4117,N_4138);
xor U5866 (N_5866,N_3577,N_4393);
and U5867 (N_5867,N_3790,N_3646);
nor U5868 (N_5868,N_3746,N_3214);
nand U5869 (N_5869,N_4346,N_3785);
nand U5870 (N_5870,N_3609,N_3238);
nand U5871 (N_5871,N_3545,N_3876);
and U5872 (N_5872,N_4474,N_4047);
or U5873 (N_5873,N_4404,N_3707);
nand U5874 (N_5874,N_3546,N_4341);
xnor U5875 (N_5875,N_3762,N_3456);
and U5876 (N_5876,N_3338,N_3353);
xnor U5877 (N_5877,N_3505,N_3607);
and U5878 (N_5878,N_3045,N_3948);
or U5879 (N_5879,N_3633,N_3026);
xor U5880 (N_5880,N_3750,N_3450);
nand U5881 (N_5881,N_3600,N_4391);
nor U5882 (N_5882,N_3795,N_3837);
nand U5883 (N_5883,N_3341,N_4484);
xnor U5884 (N_5884,N_3531,N_3346);
nor U5885 (N_5885,N_3581,N_3924);
nand U5886 (N_5886,N_3637,N_3300);
or U5887 (N_5887,N_3638,N_3908);
or U5888 (N_5888,N_3363,N_3407);
nand U5889 (N_5889,N_3176,N_3024);
nor U5890 (N_5890,N_4014,N_3413);
or U5891 (N_5891,N_3826,N_3962);
and U5892 (N_5892,N_3107,N_3760);
nand U5893 (N_5893,N_4480,N_3468);
nor U5894 (N_5894,N_4049,N_3310);
nor U5895 (N_5895,N_4338,N_4223);
and U5896 (N_5896,N_3903,N_4339);
nand U5897 (N_5897,N_3924,N_3162);
and U5898 (N_5898,N_4366,N_4075);
nor U5899 (N_5899,N_3236,N_3683);
nor U5900 (N_5900,N_3360,N_3137);
nor U5901 (N_5901,N_4326,N_3490);
xnor U5902 (N_5902,N_3710,N_4236);
or U5903 (N_5903,N_3604,N_3916);
nor U5904 (N_5904,N_3278,N_3661);
and U5905 (N_5905,N_3093,N_4002);
or U5906 (N_5906,N_3908,N_3409);
xor U5907 (N_5907,N_3309,N_3067);
nor U5908 (N_5908,N_3979,N_3092);
nor U5909 (N_5909,N_4216,N_4321);
nor U5910 (N_5910,N_3325,N_3278);
xor U5911 (N_5911,N_3824,N_4391);
nand U5912 (N_5912,N_3874,N_3036);
xor U5913 (N_5913,N_3821,N_4278);
xnor U5914 (N_5914,N_3220,N_4331);
xor U5915 (N_5915,N_3687,N_4483);
xor U5916 (N_5916,N_4130,N_3398);
nand U5917 (N_5917,N_4463,N_4043);
nand U5918 (N_5918,N_3709,N_3412);
nor U5919 (N_5919,N_3073,N_3453);
nor U5920 (N_5920,N_3653,N_3632);
and U5921 (N_5921,N_4192,N_3591);
xor U5922 (N_5922,N_3358,N_3194);
or U5923 (N_5923,N_3230,N_3776);
and U5924 (N_5924,N_3973,N_3096);
nor U5925 (N_5925,N_3538,N_4451);
or U5926 (N_5926,N_4109,N_4191);
nand U5927 (N_5927,N_3955,N_3099);
and U5928 (N_5928,N_3735,N_3719);
xnor U5929 (N_5929,N_3177,N_3840);
xnor U5930 (N_5930,N_4127,N_3189);
nand U5931 (N_5931,N_3367,N_3475);
nor U5932 (N_5932,N_3134,N_3635);
and U5933 (N_5933,N_4268,N_3779);
or U5934 (N_5934,N_4075,N_3466);
nor U5935 (N_5935,N_3038,N_3176);
nor U5936 (N_5936,N_4187,N_3760);
nand U5937 (N_5937,N_3848,N_3309);
xor U5938 (N_5938,N_3857,N_3304);
xnor U5939 (N_5939,N_3319,N_3934);
nand U5940 (N_5940,N_3080,N_4115);
nor U5941 (N_5941,N_3726,N_3752);
nor U5942 (N_5942,N_4067,N_3287);
nand U5943 (N_5943,N_3364,N_3541);
and U5944 (N_5944,N_3029,N_4296);
and U5945 (N_5945,N_3689,N_3258);
and U5946 (N_5946,N_4345,N_3440);
and U5947 (N_5947,N_3048,N_4268);
or U5948 (N_5948,N_3864,N_3737);
nor U5949 (N_5949,N_4183,N_3737);
and U5950 (N_5950,N_4129,N_3803);
xor U5951 (N_5951,N_4003,N_4388);
or U5952 (N_5952,N_4472,N_3263);
nand U5953 (N_5953,N_3751,N_3541);
or U5954 (N_5954,N_3479,N_4068);
nand U5955 (N_5955,N_3923,N_3371);
nor U5956 (N_5956,N_4453,N_3959);
nand U5957 (N_5957,N_3157,N_4230);
or U5958 (N_5958,N_3149,N_4323);
and U5959 (N_5959,N_3636,N_3007);
or U5960 (N_5960,N_4456,N_3537);
xnor U5961 (N_5961,N_3300,N_3439);
or U5962 (N_5962,N_3804,N_3888);
nor U5963 (N_5963,N_4450,N_4098);
nand U5964 (N_5964,N_3831,N_4065);
nor U5965 (N_5965,N_3460,N_3132);
or U5966 (N_5966,N_4327,N_3136);
and U5967 (N_5967,N_3914,N_3831);
or U5968 (N_5968,N_3582,N_3494);
xnor U5969 (N_5969,N_3410,N_3781);
nor U5970 (N_5970,N_4145,N_3741);
and U5971 (N_5971,N_4441,N_4114);
xnor U5972 (N_5972,N_3380,N_4251);
nand U5973 (N_5973,N_3515,N_3590);
and U5974 (N_5974,N_4117,N_3153);
nor U5975 (N_5975,N_4233,N_4440);
xnor U5976 (N_5976,N_4231,N_3961);
xor U5977 (N_5977,N_3752,N_4040);
nor U5978 (N_5978,N_3746,N_3250);
nand U5979 (N_5979,N_4069,N_4470);
nand U5980 (N_5980,N_3317,N_4374);
or U5981 (N_5981,N_4139,N_4068);
or U5982 (N_5982,N_3270,N_4034);
nand U5983 (N_5983,N_3398,N_4181);
nor U5984 (N_5984,N_3707,N_3545);
xor U5985 (N_5985,N_4441,N_3803);
nor U5986 (N_5986,N_4060,N_3431);
or U5987 (N_5987,N_3729,N_4397);
or U5988 (N_5988,N_3738,N_4255);
and U5989 (N_5989,N_3846,N_4458);
and U5990 (N_5990,N_4486,N_3306);
and U5991 (N_5991,N_4229,N_4185);
nor U5992 (N_5992,N_4302,N_3429);
or U5993 (N_5993,N_3420,N_3344);
nand U5994 (N_5994,N_3296,N_3402);
nor U5995 (N_5995,N_3537,N_3723);
or U5996 (N_5996,N_4158,N_3352);
xor U5997 (N_5997,N_3391,N_4248);
nor U5998 (N_5998,N_3670,N_3793);
nand U5999 (N_5999,N_3641,N_3627);
nand U6000 (N_6000,N_4773,N_5429);
xnor U6001 (N_6001,N_5334,N_5109);
nand U6002 (N_6002,N_5759,N_5187);
or U6003 (N_6003,N_4526,N_5596);
or U6004 (N_6004,N_5328,N_5948);
and U6005 (N_6005,N_5515,N_5487);
xor U6006 (N_6006,N_5704,N_4923);
nor U6007 (N_6007,N_5947,N_4638);
xnor U6008 (N_6008,N_5053,N_5922);
and U6009 (N_6009,N_5047,N_4739);
nor U6010 (N_6010,N_5503,N_5159);
or U6011 (N_6011,N_4574,N_4755);
nor U6012 (N_6012,N_5273,N_4600);
or U6013 (N_6013,N_5306,N_5703);
and U6014 (N_6014,N_4531,N_5702);
nand U6015 (N_6015,N_5483,N_5789);
nand U6016 (N_6016,N_4653,N_4919);
and U6017 (N_6017,N_5643,N_5447);
or U6018 (N_6018,N_5965,N_4680);
nand U6019 (N_6019,N_5903,N_5087);
and U6020 (N_6020,N_5930,N_4826);
xnor U6021 (N_6021,N_5344,N_5021);
or U6022 (N_6022,N_4718,N_5891);
and U6023 (N_6023,N_5630,N_4814);
and U6024 (N_6024,N_4895,N_5131);
nand U6025 (N_6025,N_5178,N_5627);
nand U6026 (N_6026,N_5175,N_4796);
nor U6027 (N_6027,N_5130,N_5761);
and U6028 (N_6028,N_4539,N_5656);
xor U6029 (N_6029,N_4803,N_5524);
and U6030 (N_6030,N_4972,N_4524);
nand U6031 (N_6031,N_5068,N_5368);
xor U6032 (N_6032,N_4947,N_4554);
nand U6033 (N_6033,N_5757,N_5488);
nand U6034 (N_6034,N_4980,N_4909);
or U6035 (N_6035,N_5267,N_5218);
xnor U6036 (N_6036,N_5354,N_5849);
xor U6037 (N_6037,N_4593,N_4964);
xnor U6038 (N_6038,N_5451,N_5241);
xor U6039 (N_6039,N_5244,N_4658);
nor U6040 (N_6040,N_5998,N_5291);
xnor U6041 (N_6041,N_5138,N_4590);
nand U6042 (N_6042,N_5339,N_5404);
nand U6043 (N_6043,N_5409,N_5917);
nand U6044 (N_6044,N_4904,N_4830);
xor U6045 (N_6045,N_5071,N_4829);
nor U6046 (N_6046,N_5696,N_5212);
or U6047 (N_6047,N_5500,N_5106);
nand U6048 (N_6048,N_4965,N_5502);
and U6049 (N_6049,N_5282,N_5747);
xor U6050 (N_6050,N_5126,N_5443);
or U6051 (N_6051,N_4963,N_4881);
or U6052 (N_6052,N_5372,N_4591);
nand U6053 (N_6053,N_5235,N_5842);
nor U6054 (N_6054,N_4940,N_4686);
xor U6055 (N_6055,N_5781,N_5464);
or U6056 (N_6056,N_5101,N_5380);
or U6057 (N_6057,N_4956,N_5915);
nand U6058 (N_6058,N_5543,N_5466);
nor U6059 (N_6059,N_5506,N_4903);
nor U6060 (N_6060,N_5225,N_5685);
nor U6061 (N_6061,N_4777,N_5712);
nor U6062 (N_6062,N_4995,N_5496);
and U6063 (N_6063,N_5582,N_5555);
and U6064 (N_6064,N_5918,N_5646);
or U6065 (N_6065,N_5631,N_5878);
or U6066 (N_6066,N_4540,N_5529);
nand U6067 (N_6067,N_5705,N_4737);
nor U6068 (N_6068,N_5504,N_4886);
and U6069 (N_6069,N_4618,N_5557);
nand U6070 (N_6070,N_4620,N_5804);
nor U6071 (N_6071,N_5371,N_5148);
or U6072 (N_6072,N_5462,N_5883);
nand U6073 (N_6073,N_5049,N_4669);
or U6074 (N_6074,N_4579,N_5870);
xnor U6075 (N_6075,N_4671,N_5052);
or U6076 (N_6076,N_5573,N_4977);
nor U6077 (N_6077,N_4610,N_5024);
nor U6078 (N_6078,N_5494,N_5223);
or U6079 (N_6079,N_4897,N_5424);
nand U6080 (N_6080,N_5015,N_4882);
or U6081 (N_6081,N_4894,N_5739);
nand U6082 (N_6082,N_5194,N_4797);
and U6083 (N_6083,N_5280,N_5365);
or U6084 (N_6084,N_4549,N_4901);
nor U6085 (N_6085,N_5511,N_5410);
or U6086 (N_6086,N_4898,N_5794);
or U6087 (N_6087,N_4890,N_5632);
xor U6088 (N_6088,N_5304,N_5420);
and U6089 (N_6089,N_4765,N_5377);
xor U6090 (N_6090,N_5875,N_5622);
and U6091 (N_6091,N_5871,N_5990);
xor U6092 (N_6092,N_5142,N_4966);
or U6093 (N_6093,N_5208,N_4553);
or U6094 (N_6094,N_5214,N_5825);
or U6095 (N_6095,N_5498,N_5690);
and U6096 (N_6096,N_5754,N_4837);
and U6097 (N_6097,N_5128,N_5394);
and U6098 (N_6098,N_5822,N_5821);
nor U6099 (N_6099,N_5248,N_4706);
xnor U6100 (N_6100,N_5165,N_4793);
nand U6101 (N_6101,N_5491,N_4850);
xnor U6102 (N_6102,N_5960,N_5499);
nor U6103 (N_6103,N_5415,N_5993);
nor U6104 (N_6104,N_4536,N_4592);
xor U6105 (N_6105,N_5872,N_5076);
and U6106 (N_6106,N_5974,N_5433);
nor U6107 (N_6107,N_5820,N_4975);
nand U6108 (N_6108,N_5356,N_5459);
nand U6109 (N_6109,N_5294,N_5327);
xnor U6110 (N_6110,N_5714,N_5120);
nor U6111 (N_6111,N_4869,N_4845);
xor U6112 (N_6112,N_5609,N_5036);
or U6113 (N_6113,N_5069,N_4884);
nand U6114 (N_6114,N_4585,N_5435);
nand U6115 (N_6115,N_5749,N_4629);
nand U6116 (N_6116,N_5580,N_4883);
nor U6117 (N_6117,N_5710,N_4717);
xnor U6118 (N_6118,N_5261,N_5363);
nor U6119 (N_6119,N_5230,N_5110);
and U6120 (N_6120,N_5341,N_5833);
or U6121 (N_6121,N_4969,N_4509);
nand U6122 (N_6122,N_5654,N_5669);
and U6123 (N_6123,N_4785,N_5364);
xor U6124 (N_6124,N_5533,N_5064);
nor U6125 (N_6125,N_5736,N_4985);
nand U6126 (N_6126,N_5399,N_5886);
nand U6127 (N_6127,N_4959,N_5001);
nor U6128 (N_6128,N_4728,N_5285);
or U6129 (N_6129,N_5122,N_5127);
or U6130 (N_6130,N_5684,N_4954);
or U6131 (N_6131,N_5207,N_5297);
xnor U6132 (N_6132,N_5318,N_4968);
nand U6133 (N_6133,N_5890,N_5492);
and U6134 (N_6134,N_4730,N_5783);
nand U6135 (N_6135,N_4819,N_5608);
or U6136 (N_6136,N_5835,N_5994);
or U6137 (N_6137,N_4582,N_5210);
and U6138 (N_6138,N_4707,N_4696);
nor U6139 (N_6139,N_5260,N_4668);
or U6140 (N_6140,N_4973,N_5062);
or U6141 (N_6141,N_4564,N_5427);
and U6142 (N_6142,N_4587,N_5626);
or U6143 (N_6143,N_5302,N_5834);
nor U6144 (N_6144,N_5139,N_5920);
nand U6145 (N_6145,N_5895,N_4609);
and U6146 (N_6146,N_4544,N_4512);
or U6147 (N_6147,N_5972,N_5751);
or U6148 (N_6148,N_5839,N_5495);
xor U6149 (N_6149,N_5253,N_5800);
or U6150 (N_6150,N_4948,N_5135);
and U6151 (N_6151,N_5486,N_5648);
or U6152 (N_6152,N_4580,N_4859);
and U6153 (N_6153,N_4682,N_4925);
or U6154 (N_6154,N_4659,N_5811);
nor U6155 (N_6155,N_5475,N_4762);
nor U6156 (N_6156,N_4831,N_4603);
nor U6157 (N_6157,N_5659,N_4503);
nand U6158 (N_6158,N_4839,N_5108);
or U6159 (N_6159,N_4945,N_5432);
nor U6160 (N_6160,N_5768,N_5683);
and U6161 (N_6161,N_5211,N_5750);
nor U6162 (N_6162,N_5061,N_5925);
or U6163 (N_6163,N_5691,N_5414);
nor U6164 (N_6164,N_4676,N_5317);
xnor U6165 (N_6165,N_5172,N_4962);
nor U6166 (N_6166,N_5828,N_5154);
and U6167 (N_6167,N_5619,N_4644);
and U6168 (N_6168,N_5634,N_5203);
and U6169 (N_6169,N_5545,N_4841);
nand U6170 (N_6170,N_5314,N_4936);
nor U6171 (N_6171,N_4781,N_4753);
and U6172 (N_6172,N_5168,N_5284);
nand U6173 (N_6173,N_5124,N_5269);
or U6174 (N_6174,N_5330,N_5186);
nor U6175 (N_6175,N_5863,N_5660);
or U6176 (N_6176,N_5664,N_4763);
xor U6177 (N_6177,N_5150,N_4997);
xor U6178 (N_6178,N_4601,N_5647);
and U6179 (N_6179,N_5801,N_4971);
xnor U6180 (N_6180,N_5033,N_5578);
nor U6181 (N_6181,N_4542,N_5549);
xnor U6182 (N_6182,N_5478,N_4703);
xnor U6183 (N_6183,N_4723,N_5403);
nand U6184 (N_6184,N_5125,N_5376);
and U6185 (N_6185,N_5778,N_4943);
xor U6186 (N_6186,N_5075,N_5985);
xor U6187 (N_6187,N_4566,N_5694);
xnor U6188 (N_6188,N_4999,N_5472);
xor U6189 (N_6189,N_4941,N_4705);
or U6190 (N_6190,N_5845,N_5787);
or U6191 (N_6191,N_5926,N_5590);
nor U6192 (N_6192,N_4749,N_5020);
xor U6193 (N_6193,N_4887,N_5982);
nand U6194 (N_6194,N_4533,N_5426);
nand U6195 (N_6195,N_5671,N_4993);
xnor U6196 (N_6196,N_5591,N_5098);
and U6197 (N_6197,N_4710,N_5239);
xor U6198 (N_6198,N_5322,N_5114);
and U6199 (N_6199,N_5968,N_5310);
or U6200 (N_6200,N_5229,N_5594);
or U6201 (N_6201,N_4761,N_5850);
or U6202 (N_6202,N_4513,N_5575);
nor U6203 (N_6203,N_5640,N_4545);
xor U6204 (N_6204,N_4873,N_5692);
xor U6205 (N_6205,N_5010,N_5962);
or U6206 (N_6206,N_4987,N_4794);
and U6207 (N_6207,N_5852,N_4674);
nor U6208 (N_6208,N_4608,N_4507);
xor U6209 (N_6209,N_5123,N_4506);
and U6210 (N_6210,N_4516,N_5234);
nand U6211 (N_6211,N_5205,N_5658);
or U6212 (N_6212,N_5966,N_5748);
or U6213 (N_6213,N_5044,N_5772);
and U6214 (N_6214,N_5180,N_5119);
nand U6215 (N_6215,N_5961,N_5535);
nor U6216 (N_6216,N_4976,N_5182);
xor U6217 (N_6217,N_5653,N_5516);
and U6218 (N_6218,N_5100,N_4858);
or U6219 (N_6219,N_4892,N_5538);
nor U6220 (N_6220,N_4934,N_5989);
or U6221 (N_6221,N_5268,N_5290);
nand U6222 (N_6222,N_4701,N_5406);
and U6223 (N_6223,N_5458,N_4991);
xnor U6224 (N_6224,N_4888,N_5308);
nor U6225 (N_6225,N_4571,N_4769);
or U6226 (N_6226,N_5559,N_4570);
or U6227 (N_6227,N_5348,N_5995);
or U6228 (N_6228,N_5721,N_5861);
nand U6229 (N_6229,N_4950,N_5367);
xnor U6230 (N_6230,N_5166,N_4700);
nor U6231 (N_6231,N_4688,N_5209);
or U6232 (N_6232,N_4970,N_5774);
xor U6233 (N_6233,N_5507,N_4863);
or U6234 (N_6234,N_5170,N_5666);
nand U6235 (N_6235,N_5058,N_4846);
xor U6236 (N_6236,N_5574,N_5140);
and U6237 (N_6237,N_5887,N_5089);
and U6238 (N_6238,N_5636,N_5732);
nand U6239 (N_6239,N_4684,N_4988);
xnor U6240 (N_6240,N_5323,N_4729);
and U6241 (N_6241,N_4791,N_5333);
or U6242 (N_6242,N_5407,N_4534);
nand U6243 (N_6243,N_5534,N_4655);
nor U6244 (N_6244,N_5465,N_4986);
or U6245 (N_6245,N_5688,N_4896);
nand U6246 (N_6246,N_5892,N_4984);
and U6247 (N_6247,N_5275,N_5734);
or U6248 (N_6248,N_4646,N_5481);
nor U6249 (N_6249,N_4535,N_4860);
nor U6250 (N_6250,N_4619,N_5790);
and U6251 (N_6251,N_5980,N_4625);
or U6252 (N_6252,N_4685,N_4810);
nand U6253 (N_6253,N_5798,N_5616);
xor U6254 (N_6254,N_4944,N_5191);
and U6255 (N_6255,N_5865,N_4690);
and U6256 (N_6256,N_5817,N_5246);
nor U6257 (N_6257,N_4842,N_5944);
and U6258 (N_6258,N_5085,N_4586);
xnor U6259 (N_6259,N_4771,N_5908);
and U6260 (N_6260,N_5793,N_5400);
or U6261 (N_6261,N_5661,N_5039);
xnor U6262 (N_6262,N_4935,N_4556);
nor U6263 (N_6263,N_5625,N_4721);
and U6264 (N_6264,N_4648,N_5358);
nor U6265 (N_6265,N_4900,N_5652);
or U6266 (N_6266,N_5452,N_5564);
xnor U6267 (N_6267,N_5397,N_4800);
and U6268 (N_6268,N_5855,N_4697);
nor U6269 (N_6269,N_5031,N_4760);
or U6270 (N_6270,N_5796,N_4645);
or U6271 (N_6271,N_5450,N_4661);
nor U6272 (N_6272,N_5996,N_4809);
nand U6273 (N_6273,N_4546,N_5907);
or U6274 (N_6274,N_5866,N_4640);
and U6275 (N_6275,N_5293,N_5336);
and U6276 (N_6276,N_5715,N_5467);
nor U6277 (N_6277,N_5206,N_5179);
or U6278 (N_6278,N_5086,N_5489);
nand U6279 (N_6279,N_5614,N_5418);
and U6280 (N_6280,N_5392,N_4994);
xor U6281 (N_6281,N_4930,N_5271);
nand U6282 (N_6282,N_4530,N_5473);
or U6283 (N_6283,N_5836,N_5526);
nor U6284 (N_6284,N_4905,N_5542);
and U6285 (N_6285,N_5411,N_5813);
nor U6286 (N_6286,N_5355,N_4504);
nor U6287 (N_6287,N_5588,N_5988);
and U6288 (N_6288,N_5357,N_5953);
and U6289 (N_6289,N_5065,N_5784);
nor U6290 (N_6290,N_4879,N_5074);
or U6291 (N_6291,N_5107,N_4612);
nor U6292 (N_6292,N_4912,N_5373);
nand U6293 (N_6293,N_5252,N_5583);
or U6294 (N_6294,N_5862,N_5025);
nor U6295 (N_6295,N_5532,N_4604);
nand U6296 (N_6296,N_5600,N_4522);
xor U6297 (N_6297,N_4689,N_5837);
nand U6298 (N_6298,N_5675,N_4584);
and U6299 (N_6299,N_5490,N_4572);
xnor U6300 (N_6300,N_5421,N_4937);
xor U6301 (N_6301,N_5188,N_5933);
and U6302 (N_6302,N_5519,N_5164);
xnor U6303 (N_6303,N_5547,N_4624);
nand U6304 (N_6304,N_4704,N_5117);
and U6305 (N_6305,N_5566,N_4577);
nand U6306 (N_6306,N_5799,N_5957);
nand U6307 (N_6307,N_5932,N_4820);
or U6308 (N_6308,N_5196,N_4754);
nand U6309 (N_6309,N_5349,N_5169);
nor U6310 (N_6310,N_5711,N_4508);
xnor U6311 (N_6311,N_4691,N_5938);
and U6312 (N_6312,N_4727,N_5958);
or U6313 (N_6313,N_5325,N_5343);
nand U6314 (N_6314,N_5305,N_5389);
or U6315 (N_6315,N_4982,N_5551);
or U6316 (N_6316,N_5073,N_5092);
and U6317 (N_6317,N_5359,N_4938);
and U6318 (N_6318,N_5552,N_5617);
or U6319 (N_6319,N_5638,N_5278);
nor U6320 (N_6320,N_5263,N_5904);
nand U6321 (N_6321,N_5642,N_4872);
nor U6322 (N_6322,N_5174,N_5782);
nand U6323 (N_6323,N_5022,N_5760);
nor U6324 (N_6324,N_5620,N_5541);
nor U6325 (N_6325,N_4630,N_5824);
nand U6326 (N_6326,N_4654,N_5222);
nor U6327 (N_6327,N_5550,N_5449);
nand U6328 (N_6328,N_4775,N_4731);
xnor U6329 (N_6329,N_5158,N_5160);
xor U6330 (N_6330,N_4565,N_5381);
nand U6331 (N_6331,N_5242,N_5934);
and U6332 (N_6332,N_5350,N_5385);
xnor U6333 (N_6333,N_4548,N_4924);
xnor U6334 (N_6334,N_4525,N_4695);
nand U6335 (N_6335,N_5697,N_5192);
or U6336 (N_6336,N_4650,N_4768);
xor U6337 (N_6337,N_5238,N_5665);
nor U6338 (N_6338,N_5416,N_5718);
xnor U6339 (N_6339,N_5561,N_5303);
nor U6340 (N_6340,N_5040,N_5581);
or U6341 (N_6341,N_5037,N_5687);
xnor U6342 (N_6342,N_5019,N_5362);
nor U6343 (N_6343,N_5914,N_5729);
xor U6344 (N_6344,N_4741,N_5240);
and U6345 (N_6345,N_5147,N_4817);
or U6346 (N_6346,N_5963,N_5227);
nand U6347 (N_6347,N_4505,N_4597);
and U6348 (N_6348,N_5606,N_5233);
or U6349 (N_6349,N_5510,N_5383);
nor U6350 (N_6350,N_5902,N_4569);
nand U6351 (N_6351,N_4926,N_4878);
or U6352 (N_6352,N_5973,N_5059);
and U6353 (N_6353,N_4917,N_5943);
nand U6354 (N_6354,N_5528,N_4871);
nand U6355 (N_6355,N_5807,N_5931);
xor U6356 (N_6356,N_5326,N_5346);
xor U6357 (N_6357,N_4665,N_4520);
or U6358 (N_6358,N_4621,N_5942);
xnor U6359 (N_6359,N_5482,N_5522);
xor U6360 (N_6360,N_5030,N_5497);
and U6361 (N_6361,N_4713,N_4805);
xor U6362 (N_6362,N_5558,N_4742);
and U6363 (N_6363,N_5078,N_4672);
or U6364 (N_6364,N_5217,N_5713);
or U6365 (N_6365,N_4679,N_5689);
or U6366 (N_6366,N_5032,N_5624);
nor U6367 (N_6367,N_5141,N_5144);
or U6368 (N_6368,N_5706,N_5313);
or U6369 (N_6369,N_5262,N_5909);
and U6370 (N_6370,N_5716,N_4617);
nor U6371 (N_6371,N_4596,N_5352);
nand U6372 (N_6372,N_5319,N_4631);
nand U6373 (N_6373,N_5765,N_5727);
and U6374 (N_6374,N_5929,N_5826);
nand U6375 (N_6375,N_4551,N_4594);
nor U6376 (N_6376,N_5779,N_5231);
xor U6377 (N_6377,N_5412,N_5093);
nand U6378 (N_6378,N_4996,N_5113);
and U6379 (N_6379,N_5738,N_5115);
nor U6380 (N_6380,N_5423,N_5539);
nor U6381 (N_6381,N_4989,N_5224);
or U6382 (N_6382,N_5129,N_4849);
xor U6383 (N_6383,N_5876,N_5655);
or U6384 (N_6384,N_5361,N_4720);
and U6385 (N_6385,N_5805,N_4714);
and U6386 (N_6386,N_5257,N_4974);
and U6387 (N_6387,N_5080,N_4613);
and U6388 (N_6388,N_5476,N_5593);
nor U6389 (N_6389,N_4847,N_4877);
nor U6390 (N_6390,N_5088,N_5770);
xnor U6391 (N_6391,N_5637,N_4795);
and U6392 (N_6392,N_5949,N_5753);
and U6393 (N_6393,N_5369,N_4666);
nand U6394 (N_6394,N_4560,N_4957);
xnor U6395 (N_6395,N_5288,N_4527);
nand U6396 (N_6396,N_4519,N_5151);
nor U6397 (N_6397,N_4615,N_5668);
nor U6398 (N_6398,N_5898,N_5514);
nand U6399 (N_6399,N_5347,N_5844);
nor U6400 (N_6400,N_5266,N_5457);
and U6401 (N_6401,N_5301,N_5201);
nand U6402 (N_6402,N_4914,N_4766);
nand U6403 (N_6403,N_4783,N_5220);
nand U6404 (N_6404,N_4614,N_5145);
nand U6405 (N_6405,N_5513,N_5621);
nor U6406 (N_6406,N_5084,N_5448);
nand U6407 (N_6407,N_4902,N_4911);
or U6408 (N_6408,N_4708,N_4824);
or U6409 (N_6409,N_5454,N_5795);
and U6410 (N_6410,N_5888,N_4855);
nand U6411 (N_6411,N_5924,N_5309);
xor U6412 (N_6412,N_5708,N_5936);
or U6413 (N_6413,N_4568,N_5353);
and U6414 (N_6414,N_5132,N_5298);
nor U6415 (N_6415,N_4838,N_5742);
and U6416 (N_6416,N_5598,N_5374);
nand U6417 (N_6417,N_5786,N_5912);
or U6418 (N_6418,N_5913,N_5873);
and U6419 (N_6419,N_4874,N_4663);
xor U6420 (N_6420,N_5480,N_4677);
xor U6421 (N_6421,N_5332,N_5366);
or U6422 (N_6422,N_4643,N_4960);
nand U6423 (N_6423,N_4853,N_4811);
nand U6424 (N_6424,N_5921,N_4748);
or U6425 (N_6425,N_5446,N_5463);
and U6426 (N_6426,N_5830,N_5281);
xor U6427 (N_6427,N_4514,N_4583);
nand U6428 (N_6428,N_4547,N_5417);
nor U6429 (N_6429,N_5901,N_5629);
or U6430 (N_6430,N_5011,N_5964);
nor U6431 (N_6431,N_5384,N_5556);
or U6432 (N_6432,N_4744,N_5846);
and U6433 (N_6433,N_4555,N_5342);
nand U6434 (N_6434,N_5885,N_4670);
and U6435 (N_6435,N_5816,N_4918);
xnor U6436 (N_6436,N_4511,N_5419);
xnor U6437 (N_6437,N_5893,N_4848);
nor U6438 (N_6438,N_5563,N_5243);
nand U6439 (N_6439,N_5752,N_4920);
nor U6440 (N_6440,N_4702,N_5329);
and U6441 (N_6441,N_4589,N_5766);
nor U6442 (N_6442,N_4861,N_4857);
and U6443 (N_6443,N_4864,N_5610);
xnor U6444 (N_6444,N_5916,N_5405);
and U6445 (N_6445,N_5681,N_5940);
nor U6446 (N_6446,N_5111,N_5858);
xor U6447 (N_6447,N_5340,N_5678);
nor U6448 (N_6448,N_5345,N_5613);
xor U6449 (N_6449,N_4953,N_4823);
or U6450 (N_6450,N_5853,N_5012);
nor U6451 (N_6451,N_5388,N_5969);
or U6452 (N_6452,N_4757,N_4808);
nor U6453 (N_6453,N_5202,N_5177);
and U6454 (N_6454,N_5009,N_4758);
or U6455 (N_6455,N_4538,N_4906);
nor U6456 (N_6456,N_5562,N_5152);
and U6457 (N_6457,N_5823,N_5283);
nor U6458 (N_6458,N_5264,N_5173);
or U6459 (N_6459,N_4868,N_5146);
and U6460 (N_6460,N_4818,N_4578);
and U6461 (N_6461,N_5584,N_5808);
nor U6462 (N_6462,N_4628,N_5398);
nand U6463 (N_6463,N_5693,N_4747);
nor U6464 (N_6464,N_5276,N_4598);
nor U6465 (N_6465,N_5193,N_4709);
or U6466 (N_6466,N_5512,N_5091);
xor U6467 (N_6467,N_5952,N_5444);
nor U6468 (N_6468,N_5181,N_5767);
nor U6469 (N_6469,N_5540,N_5521);
nor U6470 (N_6470,N_4699,N_5859);
nor U6471 (N_6471,N_5247,N_5546);
nor U6472 (N_6472,N_4929,N_4532);
or U6473 (N_6473,N_4932,N_4942);
xor U6474 (N_6474,N_4961,N_5587);
nand U6475 (N_6475,N_5937,N_4518);
nor U6476 (N_6476,N_5818,N_4812);
nor U6477 (N_6477,N_5396,N_4559);
nand U6478 (N_6478,N_5945,N_5992);
nand U6479 (N_6479,N_5469,N_5649);
nor U6480 (N_6480,N_4622,N_4635);
xor U6481 (N_6481,N_4876,N_5197);
nor U6482 (N_6482,N_5055,N_5440);
nand U6483 (N_6483,N_4541,N_5889);
or U6484 (N_6484,N_5956,N_4664);
nor U6485 (N_6485,N_5189,N_4743);
xor U6486 (N_6486,N_5723,N_5097);
nor U6487 (N_6487,N_4693,N_4740);
or U6488 (N_6488,N_5300,N_4832);
nor U6489 (N_6489,N_5679,N_4799);
xnor U6490 (N_6490,N_5571,N_4933);
xnor U6491 (N_6491,N_5221,N_5335);
xnor U6492 (N_6492,N_5390,N_5250);
nor U6493 (N_6493,N_5360,N_5215);
nand U6494 (N_6494,N_5395,N_4978);
or U6495 (N_6495,N_5579,N_5762);
nor U6496 (N_6496,N_4588,N_5485);
or U6497 (N_6497,N_4567,N_4833);
nand U6498 (N_6498,N_5635,N_4642);
and U6499 (N_6499,N_5810,N_4807);
and U6500 (N_6500,N_5112,N_5628);
or U6501 (N_6501,N_5195,N_4675);
nand U6502 (N_6502,N_4722,N_5868);
or U6503 (N_6503,N_4813,N_5641);
xor U6504 (N_6504,N_4637,N_5070);
nand U6505 (N_6505,N_5391,N_4623);
or U6506 (N_6506,N_5589,N_4836);
or U6507 (N_6507,N_5331,N_5975);
or U6508 (N_6508,N_5042,N_4652);
nand U6509 (N_6509,N_4899,N_5560);
nand U6510 (N_6510,N_4502,N_5028);
or U6511 (N_6511,N_4711,N_5981);
nand U6512 (N_6512,N_5296,N_4735);
and U6513 (N_6513,N_5536,N_5508);
and U6514 (N_6514,N_5874,N_5370);
xnor U6515 (N_6515,N_5900,N_5569);
nor U6516 (N_6516,N_5585,N_5682);
xnor U6517 (N_6517,N_5006,N_5814);
nand U6518 (N_6518,N_4607,N_4922);
xor U6519 (N_6519,N_4557,N_5163);
nor U6520 (N_6520,N_5910,N_5501);
and U6521 (N_6521,N_5623,N_4678);
nor U6522 (N_6522,N_5453,N_5434);
or U6523 (N_6523,N_4774,N_5894);
or U6524 (N_6524,N_5484,N_4804);
xnor U6525 (N_6525,N_5758,N_5717);
or U6526 (N_6526,N_5987,N_5984);
or U6527 (N_6527,N_4834,N_4752);
and U6528 (N_6528,N_5848,N_5976);
or U6529 (N_6529,N_5950,N_4854);
or U6530 (N_6530,N_5431,N_4719);
or U6531 (N_6531,N_4790,N_5577);
or U6532 (N_6532,N_4776,N_4802);
nor U6533 (N_6533,N_5773,N_5063);
or U6534 (N_6534,N_5763,N_5066);
nand U6535 (N_6535,N_5155,N_4780);
nand U6536 (N_6536,N_5645,N_4647);
and U6537 (N_6537,N_5438,N_5245);
nand U6538 (N_6538,N_5102,N_5456);
nor U6539 (N_6539,N_5258,N_4751);
nor U6540 (N_6540,N_5236,N_5134);
or U6541 (N_6541,N_4952,N_4716);
or U6542 (N_6542,N_5809,N_5707);
nor U6543 (N_6543,N_5072,N_5698);
xor U6544 (N_6544,N_5274,N_4537);
and U6545 (N_6545,N_5000,N_5157);
and U6546 (N_6546,N_5199,N_4715);
or U6547 (N_6547,N_4875,N_5518);
nand U6548 (N_6548,N_4928,N_5612);
and U6549 (N_6549,N_4784,N_5094);
nor U6550 (N_6550,N_5884,N_5460);
and U6551 (N_6551,N_5797,N_5272);
nor U6552 (N_6552,N_4563,N_4990);
nand U6553 (N_6553,N_5604,N_5057);
nand U6554 (N_6554,N_5054,N_5686);
and U6555 (N_6555,N_5847,N_4649);
and U6556 (N_6556,N_4725,N_4770);
nor U6557 (N_6557,N_5295,N_5838);
and U6558 (N_6558,N_4651,N_5307);
nand U6559 (N_6559,N_4889,N_5286);
nand U6560 (N_6560,N_5840,N_5375);
and U6561 (N_6561,N_5746,N_4660);
and U6562 (N_6562,N_5014,N_5544);
and U6563 (N_6563,N_4732,N_5699);
nor U6564 (N_6564,N_4673,N_5277);
nor U6565 (N_6565,N_5387,N_4616);
or U6566 (N_6566,N_5941,N_4927);
xnor U6567 (N_6567,N_5316,N_5724);
or U6568 (N_6568,N_4611,N_4633);
or U6569 (N_6569,N_5255,N_5676);
or U6570 (N_6570,N_4981,N_4543);
xnor U6571 (N_6571,N_5785,N_5565);
xor U6572 (N_6572,N_4552,N_4798);
nand U6573 (N_6573,N_5819,N_5149);
nor U6574 (N_6574,N_5437,N_5315);
nand U6575 (N_6575,N_5156,N_5928);
and U6576 (N_6576,N_5603,N_5035);
and U6577 (N_6577,N_4756,N_5897);
nor U6578 (N_6578,N_5899,N_5116);
nor U6579 (N_6579,N_5905,N_5553);
nor U6580 (N_6580,N_5531,N_4786);
and U6581 (N_6581,N_4891,N_4595);
and U6582 (N_6582,N_5095,N_5572);
xor U6583 (N_6583,N_5857,N_5190);
xnor U6584 (N_6584,N_5537,N_5121);
nand U6585 (N_6585,N_5324,N_5923);
and U6586 (N_6586,N_4801,N_5027);
nand U6587 (N_6587,N_5137,N_5935);
xnor U6588 (N_6588,N_5812,N_5788);
and U6589 (N_6589,N_4787,N_5425);
nand U6590 (N_6590,N_5198,N_5722);
nor U6591 (N_6591,N_5841,N_4867);
nor U6592 (N_6592,N_5077,N_4632);
nand U6593 (N_6593,N_5408,N_4626);
or U6594 (N_6594,N_5393,N_5979);
nand U6595 (N_6595,N_5046,N_5806);
and U6596 (N_6596,N_5016,N_5946);
nand U6597 (N_6597,N_5311,N_4844);
xnor U6598 (N_6598,N_5663,N_5312);
or U6599 (N_6599,N_5554,N_5136);
or U6600 (N_6600,N_5041,N_5096);
or U6601 (N_6601,N_5219,N_5445);
xnor U6602 (N_6602,N_4558,N_5843);
nand U6603 (N_6603,N_5607,N_5803);
and U6604 (N_6604,N_5200,N_4683);
xor U6605 (N_6605,N_5143,N_4528);
or U6606 (N_6606,N_5701,N_5680);
and U6607 (N_6607,N_5743,N_5771);
and U6608 (N_6608,N_5733,N_5650);
and U6609 (N_6609,N_4967,N_5470);
xor U6610 (N_6610,N_5213,N_4806);
nand U6611 (N_6611,N_5048,N_5045);
and U6612 (N_6612,N_5008,N_5954);
and U6613 (N_6613,N_5337,N_4792);
and U6614 (N_6614,N_5568,N_4517);
nand U6615 (N_6615,N_4908,N_5441);
and U6616 (N_6616,N_5105,N_5651);
and U6617 (N_6617,N_4951,N_4681);
nor U6618 (N_6618,N_4843,N_5527);
nand U6619 (N_6619,N_5442,N_5735);
nand U6620 (N_6620,N_5256,N_5270);
and U6621 (N_6621,N_5461,N_5530);
or U6622 (N_6622,N_5017,N_5378);
xnor U6623 (N_6623,N_4822,N_5402);
or U6624 (N_6624,N_5896,N_5869);
nand U6625 (N_6625,N_4521,N_4767);
nor U6626 (N_6626,N_5618,N_4733);
xnor U6627 (N_6627,N_4913,N_5662);
or U6628 (N_6628,N_5162,N_4827);
or U6629 (N_6629,N_5351,N_5730);
and U6630 (N_6630,N_5018,N_5971);
xnor U6631 (N_6631,N_4529,N_5104);
and U6632 (N_6632,N_5249,N_5237);
nor U6633 (N_6633,N_5599,N_5856);
nor U6634 (N_6634,N_4575,N_5780);
nand U6635 (N_6635,N_5977,N_5677);
or U6636 (N_6636,N_5428,N_5967);
nand U6637 (N_6637,N_4955,N_4816);
xnor U6638 (N_6638,N_5775,N_5386);
nor U6639 (N_6639,N_4515,N_5505);
xor U6640 (N_6640,N_4738,N_4726);
and U6641 (N_6641,N_4550,N_5764);
nand U6642 (N_6642,N_5864,N_5602);
or U6643 (N_6643,N_4852,N_5289);
and U6644 (N_6644,N_5455,N_5867);
and U6645 (N_6645,N_4764,N_5401);
and U6646 (N_6646,N_4500,N_5379);
and U6647 (N_6647,N_5576,N_4835);
or U6648 (N_6648,N_5051,N_5430);
and U6649 (N_6649,N_4983,N_5720);
nand U6650 (N_6650,N_4501,N_5951);
xnor U6651 (N_6651,N_4992,N_4627);
nand U6652 (N_6652,N_4687,N_5725);
or U6653 (N_6653,N_5999,N_4778);
and U6654 (N_6654,N_5023,N_5667);
or U6655 (N_6655,N_4510,N_5597);
or U6656 (N_6656,N_5183,N_5474);
and U6657 (N_6657,N_5851,N_5700);
or U6658 (N_6658,N_5005,N_4788);
nor U6659 (N_6659,N_4866,N_5287);
xnor U6660 (N_6660,N_5882,N_5939);
and U6661 (N_6661,N_5745,N_5744);
and U6662 (N_6662,N_5970,N_4907);
or U6663 (N_6663,N_4636,N_4639);
and U6664 (N_6664,N_5978,N_5525);
and U6665 (N_6665,N_4759,N_4602);
or U6666 (N_6666,N_5791,N_5060);
nor U6667 (N_6667,N_5517,N_5657);
xnor U6668 (N_6668,N_4880,N_5176);
or U6669 (N_6669,N_5633,N_5832);
nor U6670 (N_6670,N_5567,N_4931);
nand U6671 (N_6671,N_4851,N_4856);
or U6672 (N_6672,N_5983,N_4734);
nor U6673 (N_6673,N_4949,N_5226);
nor U6674 (N_6674,N_5672,N_5171);
and U6675 (N_6675,N_5731,N_5959);
nor U6676 (N_6676,N_5471,N_4745);
nor U6677 (N_6677,N_5879,N_5161);
and U6678 (N_6678,N_5003,N_5259);
nand U6679 (N_6679,N_4573,N_4576);
nand U6680 (N_6680,N_5719,N_4523);
and U6681 (N_6681,N_4915,N_4662);
nand U6682 (N_6682,N_5911,N_5413);
or U6683 (N_6683,N_5099,N_5509);
nor U6684 (N_6684,N_4667,N_4840);
nor U6685 (N_6685,N_5251,N_5728);
nor U6686 (N_6686,N_4581,N_5860);
nor U6687 (N_6687,N_5955,N_5185);
xor U6688 (N_6688,N_5493,N_4634);
xnor U6689 (N_6689,N_4870,N_4782);
nand U6690 (N_6690,N_5265,N_5067);
nor U6691 (N_6691,N_5740,N_5854);
nor U6692 (N_6692,N_5204,N_4825);
nand U6693 (N_6693,N_4746,N_5133);
or U6694 (N_6694,N_5615,N_4921);
and U6695 (N_6695,N_5382,N_4862);
xor U6696 (N_6696,N_4979,N_5338);
xor U6697 (N_6697,N_4736,N_5468);
nor U6698 (N_6698,N_5601,N_5043);
nor U6699 (N_6699,N_5320,N_4916);
and U6700 (N_6700,N_5997,N_4910);
nand U6701 (N_6701,N_4561,N_5299);
nand U6702 (N_6702,N_5991,N_4893);
xnor U6703 (N_6703,N_5079,N_5292);
and U6704 (N_6704,N_5709,N_5802);
xnor U6705 (N_6705,N_5232,N_5279);
nor U6706 (N_6706,N_5477,N_5674);
or U6707 (N_6707,N_5479,N_5007);
xor U6708 (N_6708,N_5034,N_4998);
or U6709 (N_6709,N_4694,N_4698);
nor U6710 (N_6710,N_5986,N_5611);
and U6711 (N_6711,N_4815,N_4712);
nor U6712 (N_6712,N_4958,N_4946);
xor U6713 (N_6713,N_5026,N_5831);
nor U6714 (N_6714,N_5906,N_5090);
or U6715 (N_6715,N_5737,N_4562);
or U6716 (N_6716,N_4885,N_5002);
nand U6717 (N_6717,N_5439,N_5777);
or U6718 (N_6718,N_4606,N_4599);
nor U6719 (N_6719,N_5321,N_5167);
and U6720 (N_6720,N_5927,N_5670);
nor U6721 (N_6721,N_4657,N_5881);
or U6722 (N_6722,N_5595,N_5029);
xnor U6723 (N_6723,N_5013,N_5755);
or U6724 (N_6724,N_5216,N_5038);
nand U6725 (N_6725,N_5880,N_4789);
xnor U6726 (N_6726,N_5254,N_5726);
xnor U6727 (N_6727,N_5639,N_4605);
nand U6728 (N_6728,N_5081,N_5082);
xor U6729 (N_6729,N_4779,N_5548);
nor U6730 (N_6730,N_5792,N_5673);
and U6731 (N_6731,N_5184,N_4821);
and U6732 (N_6732,N_5422,N_5829);
nor U6733 (N_6733,N_5004,N_4939);
and U6734 (N_6734,N_4656,N_5592);
nand U6735 (N_6735,N_5877,N_5153);
nor U6736 (N_6736,N_4865,N_4641);
and U6737 (N_6737,N_4692,N_4772);
nand U6738 (N_6738,N_5769,N_5436);
and U6739 (N_6739,N_5056,N_5228);
xnor U6740 (N_6740,N_5118,N_5520);
nor U6741 (N_6741,N_5644,N_5523);
nor U6742 (N_6742,N_5815,N_5586);
nand U6743 (N_6743,N_4724,N_4750);
nor U6744 (N_6744,N_5083,N_4828);
nor U6745 (N_6745,N_5695,N_5776);
nor U6746 (N_6746,N_5756,N_5103);
xnor U6747 (N_6747,N_5570,N_5605);
or U6748 (N_6748,N_5741,N_5827);
and U6749 (N_6749,N_5919,N_5050);
or U6750 (N_6750,N_5065,N_5372);
xor U6751 (N_6751,N_4942,N_5560);
nand U6752 (N_6752,N_5907,N_5318);
nor U6753 (N_6753,N_5087,N_5802);
nor U6754 (N_6754,N_5303,N_5540);
or U6755 (N_6755,N_4579,N_5524);
nand U6756 (N_6756,N_4526,N_5274);
nand U6757 (N_6757,N_4836,N_4922);
nand U6758 (N_6758,N_5382,N_5546);
and U6759 (N_6759,N_5023,N_5347);
nor U6760 (N_6760,N_5220,N_5414);
xnor U6761 (N_6761,N_5594,N_4975);
or U6762 (N_6762,N_4761,N_4913);
or U6763 (N_6763,N_5125,N_5646);
xnor U6764 (N_6764,N_4944,N_5292);
xnor U6765 (N_6765,N_5147,N_5773);
or U6766 (N_6766,N_5289,N_4863);
nand U6767 (N_6767,N_4617,N_4859);
nand U6768 (N_6768,N_5379,N_5307);
nand U6769 (N_6769,N_4836,N_5899);
and U6770 (N_6770,N_4733,N_5905);
nor U6771 (N_6771,N_5709,N_4827);
xor U6772 (N_6772,N_5726,N_5619);
and U6773 (N_6773,N_4594,N_5736);
nor U6774 (N_6774,N_5346,N_4668);
nor U6775 (N_6775,N_5625,N_5256);
and U6776 (N_6776,N_5457,N_5289);
nand U6777 (N_6777,N_4615,N_5939);
nand U6778 (N_6778,N_4537,N_5587);
nor U6779 (N_6779,N_5107,N_5757);
or U6780 (N_6780,N_4553,N_5615);
xor U6781 (N_6781,N_4960,N_5032);
xnor U6782 (N_6782,N_5765,N_4551);
nand U6783 (N_6783,N_4779,N_5061);
or U6784 (N_6784,N_5645,N_4705);
or U6785 (N_6785,N_5827,N_5889);
xor U6786 (N_6786,N_5118,N_5204);
and U6787 (N_6787,N_5738,N_5010);
nor U6788 (N_6788,N_4703,N_5415);
nor U6789 (N_6789,N_5700,N_5502);
xor U6790 (N_6790,N_5712,N_5993);
nor U6791 (N_6791,N_4837,N_5526);
and U6792 (N_6792,N_4630,N_5269);
xnor U6793 (N_6793,N_4659,N_5361);
nor U6794 (N_6794,N_5471,N_5517);
nand U6795 (N_6795,N_4707,N_5035);
or U6796 (N_6796,N_5068,N_4622);
nand U6797 (N_6797,N_5907,N_5728);
nand U6798 (N_6798,N_5677,N_5160);
or U6799 (N_6799,N_5063,N_4686);
or U6800 (N_6800,N_5899,N_5296);
xnor U6801 (N_6801,N_5235,N_4763);
xnor U6802 (N_6802,N_5372,N_5662);
nand U6803 (N_6803,N_5988,N_5739);
nor U6804 (N_6804,N_5652,N_5408);
xnor U6805 (N_6805,N_5003,N_5703);
or U6806 (N_6806,N_5751,N_5570);
and U6807 (N_6807,N_5270,N_5590);
nor U6808 (N_6808,N_5692,N_4633);
xnor U6809 (N_6809,N_4812,N_5975);
xnor U6810 (N_6810,N_5118,N_5514);
or U6811 (N_6811,N_4529,N_4635);
and U6812 (N_6812,N_5916,N_5673);
and U6813 (N_6813,N_5314,N_5611);
or U6814 (N_6814,N_5911,N_5455);
xor U6815 (N_6815,N_5811,N_5607);
and U6816 (N_6816,N_5121,N_5162);
xor U6817 (N_6817,N_5804,N_5420);
and U6818 (N_6818,N_5908,N_4651);
or U6819 (N_6819,N_5082,N_5037);
or U6820 (N_6820,N_5646,N_5932);
or U6821 (N_6821,N_4565,N_4961);
or U6822 (N_6822,N_5336,N_4555);
and U6823 (N_6823,N_5659,N_5898);
xor U6824 (N_6824,N_5347,N_5288);
or U6825 (N_6825,N_4805,N_4597);
xor U6826 (N_6826,N_5242,N_5941);
or U6827 (N_6827,N_4878,N_5247);
nor U6828 (N_6828,N_4931,N_5427);
nor U6829 (N_6829,N_5171,N_5541);
nor U6830 (N_6830,N_4807,N_5917);
and U6831 (N_6831,N_4656,N_5906);
nor U6832 (N_6832,N_5710,N_5711);
and U6833 (N_6833,N_5139,N_4727);
xor U6834 (N_6834,N_5181,N_5948);
nor U6835 (N_6835,N_4513,N_4633);
nor U6836 (N_6836,N_5664,N_5545);
xor U6837 (N_6837,N_5456,N_5176);
or U6838 (N_6838,N_5816,N_5556);
nand U6839 (N_6839,N_4773,N_4875);
nand U6840 (N_6840,N_4967,N_4544);
nor U6841 (N_6841,N_4539,N_5430);
nand U6842 (N_6842,N_5691,N_5107);
or U6843 (N_6843,N_5927,N_5112);
xor U6844 (N_6844,N_4863,N_5419);
xor U6845 (N_6845,N_4684,N_5665);
nand U6846 (N_6846,N_4628,N_4808);
nor U6847 (N_6847,N_5797,N_5604);
nor U6848 (N_6848,N_5421,N_5843);
or U6849 (N_6849,N_5710,N_5260);
xnor U6850 (N_6850,N_5007,N_5543);
nand U6851 (N_6851,N_4942,N_5900);
and U6852 (N_6852,N_5042,N_5184);
nand U6853 (N_6853,N_5588,N_4570);
and U6854 (N_6854,N_4655,N_5535);
nand U6855 (N_6855,N_5280,N_5635);
nor U6856 (N_6856,N_5427,N_4826);
xnor U6857 (N_6857,N_4685,N_5767);
nand U6858 (N_6858,N_5368,N_5015);
or U6859 (N_6859,N_5888,N_5360);
nor U6860 (N_6860,N_5975,N_4782);
and U6861 (N_6861,N_5472,N_4992);
nor U6862 (N_6862,N_5823,N_4544);
nand U6863 (N_6863,N_5092,N_4656);
or U6864 (N_6864,N_5722,N_5953);
or U6865 (N_6865,N_5098,N_5449);
xor U6866 (N_6866,N_5919,N_5929);
nand U6867 (N_6867,N_5099,N_5781);
xor U6868 (N_6868,N_5053,N_5923);
and U6869 (N_6869,N_5883,N_5593);
and U6870 (N_6870,N_5676,N_5113);
xor U6871 (N_6871,N_5848,N_5285);
nand U6872 (N_6872,N_5127,N_5588);
xor U6873 (N_6873,N_5875,N_5556);
and U6874 (N_6874,N_5671,N_5475);
nor U6875 (N_6875,N_5182,N_5007);
xor U6876 (N_6876,N_4937,N_4692);
xnor U6877 (N_6877,N_5956,N_5038);
nor U6878 (N_6878,N_5080,N_5939);
or U6879 (N_6879,N_5149,N_4794);
nand U6880 (N_6880,N_5845,N_5232);
and U6881 (N_6881,N_5410,N_5099);
or U6882 (N_6882,N_4819,N_5590);
nor U6883 (N_6883,N_4811,N_5529);
nand U6884 (N_6884,N_5449,N_4689);
xor U6885 (N_6885,N_5841,N_5872);
xnor U6886 (N_6886,N_5785,N_5079);
nand U6887 (N_6887,N_4538,N_4657);
nor U6888 (N_6888,N_5197,N_4549);
and U6889 (N_6889,N_5079,N_5598);
nor U6890 (N_6890,N_5912,N_5734);
xnor U6891 (N_6891,N_4942,N_5092);
nor U6892 (N_6892,N_4564,N_4902);
xor U6893 (N_6893,N_4622,N_5970);
and U6894 (N_6894,N_5517,N_4937);
or U6895 (N_6895,N_4758,N_4628);
nand U6896 (N_6896,N_4974,N_5088);
nand U6897 (N_6897,N_5556,N_5628);
nor U6898 (N_6898,N_5374,N_4647);
nor U6899 (N_6899,N_5683,N_5053);
nand U6900 (N_6900,N_5867,N_4893);
xnor U6901 (N_6901,N_5885,N_4544);
or U6902 (N_6902,N_4511,N_5518);
and U6903 (N_6903,N_5427,N_5747);
nor U6904 (N_6904,N_5424,N_5827);
or U6905 (N_6905,N_5175,N_5425);
xor U6906 (N_6906,N_5125,N_5739);
or U6907 (N_6907,N_5342,N_4843);
nand U6908 (N_6908,N_4666,N_4958);
and U6909 (N_6909,N_5614,N_4622);
or U6910 (N_6910,N_4662,N_5688);
nand U6911 (N_6911,N_5389,N_5941);
nor U6912 (N_6912,N_4790,N_5628);
xor U6913 (N_6913,N_4954,N_5892);
and U6914 (N_6914,N_5375,N_5151);
xnor U6915 (N_6915,N_5460,N_5280);
nor U6916 (N_6916,N_5390,N_4719);
and U6917 (N_6917,N_5713,N_5272);
nand U6918 (N_6918,N_5697,N_5166);
nand U6919 (N_6919,N_5370,N_5082);
xnor U6920 (N_6920,N_5282,N_4916);
or U6921 (N_6921,N_5656,N_5774);
or U6922 (N_6922,N_5843,N_5790);
or U6923 (N_6923,N_5898,N_4853);
or U6924 (N_6924,N_5221,N_4530);
or U6925 (N_6925,N_5014,N_5070);
xor U6926 (N_6926,N_4972,N_5585);
or U6927 (N_6927,N_5051,N_5878);
xor U6928 (N_6928,N_5191,N_5716);
xnor U6929 (N_6929,N_5241,N_5915);
xor U6930 (N_6930,N_4978,N_5436);
xor U6931 (N_6931,N_5821,N_5352);
nor U6932 (N_6932,N_4724,N_5975);
nand U6933 (N_6933,N_5476,N_5956);
and U6934 (N_6934,N_5561,N_5563);
or U6935 (N_6935,N_5890,N_4896);
nor U6936 (N_6936,N_4916,N_4933);
nor U6937 (N_6937,N_4704,N_5191);
nor U6938 (N_6938,N_5849,N_5405);
and U6939 (N_6939,N_4868,N_4738);
nand U6940 (N_6940,N_4967,N_5322);
xnor U6941 (N_6941,N_5034,N_4833);
xnor U6942 (N_6942,N_5072,N_5297);
or U6943 (N_6943,N_5599,N_5853);
or U6944 (N_6944,N_4913,N_5121);
nor U6945 (N_6945,N_5050,N_4743);
or U6946 (N_6946,N_4883,N_5018);
nand U6947 (N_6947,N_5038,N_5007);
and U6948 (N_6948,N_4917,N_4691);
and U6949 (N_6949,N_4923,N_5623);
nor U6950 (N_6950,N_5938,N_5242);
nand U6951 (N_6951,N_5701,N_5051);
nor U6952 (N_6952,N_5663,N_5788);
nor U6953 (N_6953,N_5667,N_4972);
nor U6954 (N_6954,N_5118,N_4938);
or U6955 (N_6955,N_5449,N_5747);
nand U6956 (N_6956,N_4514,N_4624);
xnor U6957 (N_6957,N_4814,N_4887);
nand U6958 (N_6958,N_4818,N_4532);
and U6959 (N_6959,N_5339,N_5671);
nor U6960 (N_6960,N_5369,N_5396);
and U6961 (N_6961,N_4506,N_4937);
nor U6962 (N_6962,N_5993,N_5830);
and U6963 (N_6963,N_5719,N_5275);
and U6964 (N_6964,N_5393,N_5598);
or U6965 (N_6965,N_5636,N_5734);
or U6966 (N_6966,N_5592,N_5173);
and U6967 (N_6967,N_5907,N_4551);
nand U6968 (N_6968,N_5003,N_5652);
xnor U6969 (N_6969,N_5056,N_5878);
or U6970 (N_6970,N_5786,N_5937);
xnor U6971 (N_6971,N_5766,N_5498);
or U6972 (N_6972,N_5704,N_5870);
or U6973 (N_6973,N_5292,N_5972);
nand U6974 (N_6974,N_5737,N_5348);
xor U6975 (N_6975,N_5139,N_4648);
nor U6976 (N_6976,N_5828,N_5316);
xnor U6977 (N_6977,N_5161,N_4811);
nand U6978 (N_6978,N_5949,N_4572);
xnor U6979 (N_6979,N_5019,N_5645);
xor U6980 (N_6980,N_5204,N_5526);
nand U6981 (N_6981,N_5580,N_4654);
nor U6982 (N_6982,N_5640,N_5865);
and U6983 (N_6983,N_4729,N_5470);
xnor U6984 (N_6984,N_4718,N_4775);
xor U6985 (N_6985,N_5875,N_5014);
nand U6986 (N_6986,N_5862,N_5088);
and U6987 (N_6987,N_4959,N_5870);
nor U6988 (N_6988,N_5065,N_5806);
and U6989 (N_6989,N_5965,N_4524);
and U6990 (N_6990,N_5637,N_4810);
and U6991 (N_6991,N_5456,N_5676);
xor U6992 (N_6992,N_5715,N_5437);
or U6993 (N_6993,N_5386,N_4973);
xor U6994 (N_6994,N_5499,N_5281);
nor U6995 (N_6995,N_5590,N_5148);
nand U6996 (N_6996,N_4611,N_5434);
nand U6997 (N_6997,N_5934,N_5977);
nand U6998 (N_6998,N_5042,N_5399);
nor U6999 (N_6999,N_5347,N_4986);
or U7000 (N_7000,N_5237,N_5013);
xor U7001 (N_7001,N_5822,N_5002);
xor U7002 (N_7002,N_5082,N_5640);
nand U7003 (N_7003,N_5328,N_5287);
and U7004 (N_7004,N_5316,N_5297);
or U7005 (N_7005,N_5607,N_4502);
xor U7006 (N_7006,N_4955,N_4990);
nor U7007 (N_7007,N_5692,N_4996);
xor U7008 (N_7008,N_5668,N_5828);
or U7009 (N_7009,N_4543,N_4525);
or U7010 (N_7010,N_5010,N_5793);
xnor U7011 (N_7011,N_5319,N_4679);
xor U7012 (N_7012,N_4525,N_5291);
or U7013 (N_7013,N_5154,N_4638);
nand U7014 (N_7014,N_4963,N_5573);
nor U7015 (N_7015,N_5250,N_4579);
nand U7016 (N_7016,N_4980,N_4514);
or U7017 (N_7017,N_4558,N_5785);
nor U7018 (N_7018,N_5928,N_5750);
xor U7019 (N_7019,N_4749,N_4831);
xor U7020 (N_7020,N_5045,N_4871);
nor U7021 (N_7021,N_5949,N_5633);
and U7022 (N_7022,N_5045,N_5904);
nand U7023 (N_7023,N_4824,N_5912);
or U7024 (N_7024,N_4676,N_5491);
nand U7025 (N_7025,N_4699,N_4542);
nand U7026 (N_7026,N_5435,N_4935);
nand U7027 (N_7027,N_5352,N_5049);
or U7028 (N_7028,N_5753,N_4602);
nand U7029 (N_7029,N_4607,N_4973);
nor U7030 (N_7030,N_5497,N_5610);
or U7031 (N_7031,N_4534,N_5505);
or U7032 (N_7032,N_5561,N_5150);
or U7033 (N_7033,N_5895,N_5579);
nor U7034 (N_7034,N_4868,N_5713);
xnor U7035 (N_7035,N_4555,N_5726);
nor U7036 (N_7036,N_4505,N_4626);
nor U7037 (N_7037,N_5234,N_5966);
or U7038 (N_7038,N_5238,N_4565);
and U7039 (N_7039,N_5546,N_4733);
or U7040 (N_7040,N_5486,N_4651);
nor U7041 (N_7041,N_5085,N_4746);
xnor U7042 (N_7042,N_5422,N_5849);
xnor U7043 (N_7043,N_5766,N_5753);
nor U7044 (N_7044,N_4923,N_4732);
nand U7045 (N_7045,N_5083,N_5932);
nor U7046 (N_7046,N_5477,N_4592);
nand U7047 (N_7047,N_5151,N_5419);
nor U7048 (N_7048,N_5363,N_4896);
or U7049 (N_7049,N_4934,N_5881);
nor U7050 (N_7050,N_5344,N_5529);
or U7051 (N_7051,N_5154,N_4871);
or U7052 (N_7052,N_4954,N_5937);
nand U7053 (N_7053,N_5573,N_5810);
nand U7054 (N_7054,N_4621,N_4616);
nor U7055 (N_7055,N_5539,N_5584);
or U7056 (N_7056,N_4578,N_5041);
or U7057 (N_7057,N_4643,N_5379);
nand U7058 (N_7058,N_5280,N_5312);
and U7059 (N_7059,N_5305,N_5083);
and U7060 (N_7060,N_4858,N_4721);
or U7061 (N_7061,N_5363,N_4790);
nor U7062 (N_7062,N_5948,N_5990);
or U7063 (N_7063,N_5406,N_5400);
xnor U7064 (N_7064,N_4840,N_5783);
and U7065 (N_7065,N_5892,N_4938);
and U7066 (N_7066,N_5052,N_5602);
and U7067 (N_7067,N_4539,N_5908);
or U7068 (N_7068,N_5931,N_5847);
nand U7069 (N_7069,N_5445,N_5423);
nor U7070 (N_7070,N_5029,N_5121);
and U7071 (N_7071,N_5441,N_4965);
xnor U7072 (N_7072,N_5925,N_5438);
or U7073 (N_7073,N_5914,N_4646);
nor U7074 (N_7074,N_4779,N_4679);
nor U7075 (N_7075,N_4841,N_5639);
and U7076 (N_7076,N_5805,N_4573);
xnor U7077 (N_7077,N_4639,N_4966);
xnor U7078 (N_7078,N_5292,N_4777);
xnor U7079 (N_7079,N_5319,N_5882);
or U7080 (N_7080,N_5930,N_5369);
or U7081 (N_7081,N_5345,N_5507);
or U7082 (N_7082,N_5754,N_5243);
and U7083 (N_7083,N_5274,N_5089);
xnor U7084 (N_7084,N_5403,N_5301);
and U7085 (N_7085,N_5824,N_4761);
xor U7086 (N_7086,N_4688,N_5482);
xor U7087 (N_7087,N_5812,N_4561);
nand U7088 (N_7088,N_4737,N_5418);
or U7089 (N_7089,N_4689,N_5468);
and U7090 (N_7090,N_5475,N_4895);
and U7091 (N_7091,N_5940,N_5865);
nor U7092 (N_7092,N_4775,N_4984);
nor U7093 (N_7093,N_4736,N_5186);
nor U7094 (N_7094,N_4825,N_5416);
or U7095 (N_7095,N_5132,N_5177);
and U7096 (N_7096,N_5579,N_5863);
nor U7097 (N_7097,N_4622,N_5698);
xor U7098 (N_7098,N_4791,N_5371);
xor U7099 (N_7099,N_4778,N_4672);
nand U7100 (N_7100,N_5944,N_5668);
nand U7101 (N_7101,N_4892,N_5339);
and U7102 (N_7102,N_5283,N_4955);
nor U7103 (N_7103,N_4787,N_5858);
and U7104 (N_7104,N_5619,N_5148);
nor U7105 (N_7105,N_5387,N_5016);
and U7106 (N_7106,N_5477,N_4933);
and U7107 (N_7107,N_4941,N_4830);
nor U7108 (N_7108,N_5222,N_4927);
xor U7109 (N_7109,N_5093,N_5130);
nand U7110 (N_7110,N_5862,N_4703);
and U7111 (N_7111,N_4554,N_5485);
xnor U7112 (N_7112,N_5138,N_4846);
nand U7113 (N_7113,N_5800,N_5753);
nor U7114 (N_7114,N_5493,N_5163);
xor U7115 (N_7115,N_4624,N_5589);
xor U7116 (N_7116,N_4587,N_5214);
and U7117 (N_7117,N_5387,N_4506);
xnor U7118 (N_7118,N_4520,N_4603);
nor U7119 (N_7119,N_4894,N_5064);
nand U7120 (N_7120,N_5268,N_5693);
and U7121 (N_7121,N_4920,N_5552);
and U7122 (N_7122,N_5579,N_5228);
nor U7123 (N_7123,N_5152,N_5783);
nor U7124 (N_7124,N_5870,N_4768);
and U7125 (N_7125,N_4623,N_4679);
and U7126 (N_7126,N_5920,N_5805);
nand U7127 (N_7127,N_4623,N_4738);
or U7128 (N_7128,N_5722,N_5428);
nor U7129 (N_7129,N_5478,N_5686);
nor U7130 (N_7130,N_5083,N_5486);
nand U7131 (N_7131,N_5904,N_5834);
and U7132 (N_7132,N_5266,N_4723);
nand U7133 (N_7133,N_5171,N_5034);
nor U7134 (N_7134,N_5565,N_5957);
or U7135 (N_7135,N_5891,N_4666);
and U7136 (N_7136,N_5028,N_5607);
xnor U7137 (N_7137,N_5875,N_5744);
nand U7138 (N_7138,N_5954,N_4562);
xnor U7139 (N_7139,N_5168,N_5207);
xor U7140 (N_7140,N_5097,N_5783);
or U7141 (N_7141,N_4592,N_5271);
nand U7142 (N_7142,N_5179,N_4535);
nor U7143 (N_7143,N_5656,N_5579);
xnor U7144 (N_7144,N_4750,N_5468);
nor U7145 (N_7145,N_5008,N_5158);
xnor U7146 (N_7146,N_5641,N_4920);
nor U7147 (N_7147,N_5034,N_4999);
or U7148 (N_7148,N_4518,N_5852);
xnor U7149 (N_7149,N_5127,N_5136);
nor U7150 (N_7150,N_5440,N_4827);
and U7151 (N_7151,N_5334,N_4563);
or U7152 (N_7152,N_5177,N_5877);
nor U7153 (N_7153,N_5907,N_4841);
or U7154 (N_7154,N_4952,N_4755);
nand U7155 (N_7155,N_5359,N_5361);
nand U7156 (N_7156,N_4925,N_5260);
xor U7157 (N_7157,N_4756,N_4782);
xor U7158 (N_7158,N_4778,N_4547);
xnor U7159 (N_7159,N_5968,N_5226);
xor U7160 (N_7160,N_4616,N_4904);
xor U7161 (N_7161,N_5279,N_4870);
xor U7162 (N_7162,N_5641,N_5742);
nand U7163 (N_7163,N_5153,N_5688);
xnor U7164 (N_7164,N_4616,N_4800);
xor U7165 (N_7165,N_5653,N_5645);
or U7166 (N_7166,N_5516,N_5463);
nand U7167 (N_7167,N_5639,N_4786);
nor U7168 (N_7168,N_5093,N_5090);
nor U7169 (N_7169,N_5718,N_5260);
nand U7170 (N_7170,N_5360,N_5761);
nor U7171 (N_7171,N_4706,N_4586);
and U7172 (N_7172,N_4824,N_4553);
and U7173 (N_7173,N_4536,N_5270);
nor U7174 (N_7174,N_5259,N_4658);
xor U7175 (N_7175,N_4682,N_5804);
nor U7176 (N_7176,N_5469,N_5199);
or U7177 (N_7177,N_4802,N_5963);
and U7178 (N_7178,N_5993,N_5217);
and U7179 (N_7179,N_5921,N_4871);
nor U7180 (N_7180,N_5980,N_5886);
or U7181 (N_7181,N_4732,N_4722);
nand U7182 (N_7182,N_4512,N_5612);
nand U7183 (N_7183,N_5259,N_4638);
or U7184 (N_7184,N_5748,N_4586);
and U7185 (N_7185,N_4699,N_4777);
nor U7186 (N_7186,N_5354,N_5759);
or U7187 (N_7187,N_5197,N_4695);
nand U7188 (N_7188,N_5985,N_4527);
and U7189 (N_7189,N_5528,N_5851);
xnor U7190 (N_7190,N_4831,N_5996);
and U7191 (N_7191,N_5295,N_4555);
or U7192 (N_7192,N_5663,N_4606);
nand U7193 (N_7193,N_4879,N_4563);
and U7194 (N_7194,N_4782,N_4511);
or U7195 (N_7195,N_5750,N_5539);
and U7196 (N_7196,N_5142,N_4955);
xor U7197 (N_7197,N_5004,N_5135);
or U7198 (N_7198,N_5817,N_4850);
xnor U7199 (N_7199,N_4628,N_5331);
nor U7200 (N_7200,N_5132,N_4690);
nand U7201 (N_7201,N_4528,N_5423);
or U7202 (N_7202,N_4602,N_5959);
nand U7203 (N_7203,N_5886,N_5128);
or U7204 (N_7204,N_4802,N_4775);
xnor U7205 (N_7205,N_4598,N_5406);
or U7206 (N_7206,N_5240,N_5040);
nor U7207 (N_7207,N_5224,N_5541);
or U7208 (N_7208,N_5652,N_4663);
xor U7209 (N_7209,N_4993,N_5958);
nand U7210 (N_7210,N_5478,N_5534);
or U7211 (N_7211,N_4540,N_4812);
nor U7212 (N_7212,N_4788,N_4977);
nand U7213 (N_7213,N_5987,N_4931);
nor U7214 (N_7214,N_5615,N_5544);
and U7215 (N_7215,N_5802,N_5322);
xnor U7216 (N_7216,N_5612,N_5167);
nor U7217 (N_7217,N_5124,N_5435);
nand U7218 (N_7218,N_5452,N_4964);
and U7219 (N_7219,N_4906,N_5797);
xor U7220 (N_7220,N_4624,N_5980);
and U7221 (N_7221,N_5231,N_5637);
nor U7222 (N_7222,N_5934,N_5292);
and U7223 (N_7223,N_5498,N_4570);
nor U7224 (N_7224,N_5891,N_5929);
nor U7225 (N_7225,N_5698,N_5527);
xnor U7226 (N_7226,N_5286,N_4989);
nor U7227 (N_7227,N_4887,N_5731);
or U7228 (N_7228,N_4767,N_5878);
and U7229 (N_7229,N_5540,N_4583);
nand U7230 (N_7230,N_5970,N_5761);
nor U7231 (N_7231,N_5193,N_4719);
nand U7232 (N_7232,N_5892,N_5004);
xnor U7233 (N_7233,N_4937,N_4908);
or U7234 (N_7234,N_5612,N_5778);
xnor U7235 (N_7235,N_5945,N_5889);
nor U7236 (N_7236,N_4926,N_5453);
xnor U7237 (N_7237,N_4597,N_5482);
xor U7238 (N_7238,N_5289,N_5118);
xnor U7239 (N_7239,N_5732,N_4864);
nor U7240 (N_7240,N_5819,N_5453);
nand U7241 (N_7241,N_5828,N_5945);
or U7242 (N_7242,N_5837,N_5689);
nor U7243 (N_7243,N_5285,N_4558);
nor U7244 (N_7244,N_5165,N_5609);
and U7245 (N_7245,N_4528,N_5891);
nor U7246 (N_7246,N_4564,N_5067);
nor U7247 (N_7247,N_5552,N_5626);
or U7248 (N_7248,N_4770,N_4609);
nor U7249 (N_7249,N_4661,N_5812);
nand U7250 (N_7250,N_5740,N_5342);
or U7251 (N_7251,N_5405,N_5155);
xor U7252 (N_7252,N_4856,N_5430);
or U7253 (N_7253,N_4997,N_5416);
nand U7254 (N_7254,N_5824,N_4560);
and U7255 (N_7255,N_4718,N_5652);
and U7256 (N_7256,N_4735,N_5202);
and U7257 (N_7257,N_5946,N_4525);
nand U7258 (N_7258,N_4587,N_4514);
and U7259 (N_7259,N_4852,N_5343);
nor U7260 (N_7260,N_4641,N_4967);
nand U7261 (N_7261,N_5016,N_5568);
nor U7262 (N_7262,N_5508,N_5172);
and U7263 (N_7263,N_4868,N_5587);
or U7264 (N_7264,N_5530,N_5211);
and U7265 (N_7265,N_5839,N_5763);
or U7266 (N_7266,N_5412,N_5886);
or U7267 (N_7267,N_4938,N_5008);
xor U7268 (N_7268,N_5499,N_5620);
or U7269 (N_7269,N_5421,N_5603);
xnor U7270 (N_7270,N_4562,N_4760);
nor U7271 (N_7271,N_5203,N_4948);
and U7272 (N_7272,N_5151,N_5029);
and U7273 (N_7273,N_4818,N_4910);
nand U7274 (N_7274,N_4920,N_5716);
or U7275 (N_7275,N_5616,N_4855);
and U7276 (N_7276,N_5698,N_4793);
nor U7277 (N_7277,N_5558,N_4687);
xnor U7278 (N_7278,N_4596,N_5032);
nand U7279 (N_7279,N_5859,N_5681);
and U7280 (N_7280,N_5813,N_5836);
xnor U7281 (N_7281,N_5398,N_5088);
nor U7282 (N_7282,N_4597,N_4743);
nor U7283 (N_7283,N_5013,N_4647);
and U7284 (N_7284,N_4744,N_5958);
nand U7285 (N_7285,N_4938,N_4606);
and U7286 (N_7286,N_4746,N_4873);
nand U7287 (N_7287,N_4694,N_5526);
xor U7288 (N_7288,N_5520,N_5060);
xnor U7289 (N_7289,N_4952,N_5629);
or U7290 (N_7290,N_5256,N_5859);
or U7291 (N_7291,N_4786,N_4764);
nor U7292 (N_7292,N_5896,N_5761);
or U7293 (N_7293,N_5012,N_5076);
and U7294 (N_7294,N_5067,N_5678);
xor U7295 (N_7295,N_5952,N_5932);
or U7296 (N_7296,N_4698,N_5805);
xnor U7297 (N_7297,N_5820,N_5346);
nor U7298 (N_7298,N_4708,N_5543);
xnor U7299 (N_7299,N_4855,N_5730);
xnor U7300 (N_7300,N_5607,N_4814);
or U7301 (N_7301,N_4783,N_4849);
or U7302 (N_7302,N_4505,N_5598);
nand U7303 (N_7303,N_5948,N_5256);
nor U7304 (N_7304,N_5787,N_5791);
and U7305 (N_7305,N_5564,N_4609);
nor U7306 (N_7306,N_5322,N_5724);
xnor U7307 (N_7307,N_5853,N_5534);
xnor U7308 (N_7308,N_5674,N_5406);
xor U7309 (N_7309,N_4884,N_5595);
nor U7310 (N_7310,N_5203,N_5536);
xor U7311 (N_7311,N_4827,N_5871);
and U7312 (N_7312,N_4797,N_5790);
nor U7313 (N_7313,N_4751,N_5696);
nand U7314 (N_7314,N_5300,N_5331);
and U7315 (N_7315,N_5502,N_5394);
or U7316 (N_7316,N_5912,N_5762);
nor U7317 (N_7317,N_5939,N_4992);
or U7318 (N_7318,N_4852,N_5083);
or U7319 (N_7319,N_5651,N_5991);
nor U7320 (N_7320,N_5647,N_5245);
xor U7321 (N_7321,N_4975,N_5481);
or U7322 (N_7322,N_5216,N_5379);
and U7323 (N_7323,N_5886,N_5967);
and U7324 (N_7324,N_5842,N_5488);
nor U7325 (N_7325,N_5085,N_5377);
nand U7326 (N_7326,N_5659,N_5696);
nor U7327 (N_7327,N_5326,N_4864);
nand U7328 (N_7328,N_5802,N_5234);
or U7329 (N_7329,N_4898,N_5455);
and U7330 (N_7330,N_4504,N_5528);
or U7331 (N_7331,N_5041,N_4954);
nand U7332 (N_7332,N_5098,N_4738);
xnor U7333 (N_7333,N_5807,N_5598);
and U7334 (N_7334,N_5818,N_5775);
or U7335 (N_7335,N_5035,N_5359);
nand U7336 (N_7336,N_5903,N_4565);
and U7337 (N_7337,N_5750,N_4532);
and U7338 (N_7338,N_5529,N_4747);
nand U7339 (N_7339,N_5821,N_4691);
xnor U7340 (N_7340,N_5544,N_4783);
nand U7341 (N_7341,N_4960,N_5062);
xor U7342 (N_7342,N_4514,N_4837);
nand U7343 (N_7343,N_5596,N_5464);
xor U7344 (N_7344,N_5949,N_4881);
xor U7345 (N_7345,N_5129,N_5549);
or U7346 (N_7346,N_4912,N_5736);
or U7347 (N_7347,N_5676,N_4648);
and U7348 (N_7348,N_4510,N_5133);
nor U7349 (N_7349,N_4998,N_4867);
and U7350 (N_7350,N_4875,N_5865);
or U7351 (N_7351,N_5402,N_5881);
and U7352 (N_7352,N_5472,N_4593);
xnor U7353 (N_7353,N_5712,N_5686);
xor U7354 (N_7354,N_5342,N_5300);
nand U7355 (N_7355,N_5197,N_5768);
and U7356 (N_7356,N_5647,N_4931);
or U7357 (N_7357,N_4921,N_5825);
nor U7358 (N_7358,N_5766,N_5920);
xor U7359 (N_7359,N_5127,N_5570);
nand U7360 (N_7360,N_5302,N_4716);
and U7361 (N_7361,N_4648,N_4608);
xnor U7362 (N_7362,N_4560,N_4834);
and U7363 (N_7363,N_4779,N_4933);
nor U7364 (N_7364,N_5166,N_5765);
nor U7365 (N_7365,N_5392,N_5913);
nand U7366 (N_7366,N_5181,N_4823);
nand U7367 (N_7367,N_5474,N_5081);
xor U7368 (N_7368,N_4960,N_5554);
or U7369 (N_7369,N_4905,N_5254);
nor U7370 (N_7370,N_5006,N_4891);
xor U7371 (N_7371,N_5689,N_5684);
nand U7372 (N_7372,N_4604,N_4782);
and U7373 (N_7373,N_5784,N_5571);
and U7374 (N_7374,N_5659,N_5891);
and U7375 (N_7375,N_4762,N_5131);
nand U7376 (N_7376,N_5579,N_5413);
or U7377 (N_7377,N_4888,N_5254);
nor U7378 (N_7378,N_4714,N_4698);
and U7379 (N_7379,N_4665,N_5473);
nor U7380 (N_7380,N_5445,N_4954);
or U7381 (N_7381,N_4996,N_5866);
or U7382 (N_7382,N_4729,N_5457);
nand U7383 (N_7383,N_4819,N_5933);
nor U7384 (N_7384,N_5914,N_4987);
nor U7385 (N_7385,N_5275,N_5155);
or U7386 (N_7386,N_5328,N_5698);
or U7387 (N_7387,N_5052,N_5085);
xnor U7388 (N_7388,N_5651,N_5086);
xor U7389 (N_7389,N_4623,N_5449);
or U7390 (N_7390,N_4939,N_5797);
nand U7391 (N_7391,N_5653,N_4771);
or U7392 (N_7392,N_5296,N_5403);
and U7393 (N_7393,N_5304,N_5940);
nor U7394 (N_7394,N_5791,N_5982);
and U7395 (N_7395,N_5020,N_5292);
nand U7396 (N_7396,N_5095,N_5026);
nand U7397 (N_7397,N_4791,N_5448);
nor U7398 (N_7398,N_5462,N_5833);
nand U7399 (N_7399,N_5779,N_4995);
nor U7400 (N_7400,N_4764,N_4959);
nor U7401 (N_7401,N_5336,N_5867);
or U7402 (N_7402,N_5655,N_4883);
and U7403 (N_7403,N_5705,N_5776);
xor U7404 (N_7404,N_4508,N_5494);
and U7405 (N_7405,N_5775,N_4559);
xnor U7406 (N_7406,N_5594,N_4912);
or U7407 (N_7407,N_5455,N_5215);
xnor U7408 (N_7408,N_4600,N_4915);
and U7409 (N_7409,N_5837,N_5705);
nor U7410 (N_7410,N_5413,N_5235);
nand U7411 (N_7411,N_4953,N_5380);
or U7412 (N_7412,N_5387,N_5713);
or U7413 (N_7413,N_5113,N_4896);
and U7414 (N_7414,N_5189,N_5442);
nor U7415 (N_7415,N_4891,N_5792);
or U7416 (N_7416,N_4682,N_5427);
nand U7417 (N_7417,N_5603,N_5797);
xnor U7418 (N_7418,N_5991,N_5989);
and U7419 (N_7419,N_4576,N_5638);
or U7420 (N_7420,N_5506,N_5161);
and U7421 (N_7421,N_4801,N_4772);
nand U7422 (N_7422,N_4611,N_5223);
xor U7423 (N_7423,N_5437,N_4620);
or U7424 (N_7424,N_5318,N_5972);
nor U7425 (N_7425,N_4588,N_5374);
nand U7426 (N_7426,N_5365,N_4657);
nand U7427 (N_7427,N_5946,N_4906);
nor U7428 (N_7428,N_5662,N_4692);
or U7429 (N_7429,N_5580,N_4913);
nand U7430 (N_7430,N_5764,N_4733);
nor U7431 (N_7431,N_5339,N_4913);
nand U7432 (N_7432,N_5590,N_5831);
nand U7433 (N_7433,N_5755,N_5425);
and U7434 (N_7434,N_4748,N_5502);
and U7435 (N_7435,N_4870,N_5056);
xor U7436 (N_7436,N_4662,N_4820);
or U7437 (N_7437,N_5707,N_4528);
or U7438 (N_7438,N_5403,N_5196);
nand U7439 (N_7439,N_4756,N_5981);
nor U7440 (N_7440,N_4576,N_5648);
xnor U7441 (N_7441,N_5419,N_5320);
nand U7442 (N_7442,N_4948,N_5273);
nand U7443 (N_7443,N_5162,N_5297);
or U7444 (N_7444,N_5293,N_5128);
or U7445 (N_7445,N_5492,N_5094);
xnor U7446 (N_7446,N_4880,N_5178);
and U7447 (N_7447,N_5786,N_5261);
and U7448 (N_7448,N_4901,N_4520);
xnor U7449 (N_7449,N_5730,N_5353);
xnor U7450 (N_7450,N_5844,N_4643);
or U7451 (N_7451,N_4501,N_5874);
nand U7452 (N_7452,N_5604,N_4601);
and U7453 (N_7453,N_5176,N_5081);
nand U7454 (N_7454,N_4759,N_5877);
xor U7455 (N_7455,N_5654,N_4760);
nand U7456 (N_7456,N_4636,N_5894);
nand U7457 (N_7457,N_5737,N_5774);
and U7458 (N_7458,N_5191,N_5437);
xor U7459 (N_7459,N_5009,N_5664);
nand U7460 (N_7460,N_5815,N_5973);
or U7461 (N_7461,N_5568,N_5360);
nor U7462 (N_7462,N_5767,N_5532);
or U7463 (N_7463,N_4974,N_5734);
or U7464 (N_7464,N_5542,N_4921);
or U7465 (N_7465,N_4887,N_5349);
xor U7466 (N_7466,N_5697,N_5711);
and U7467 (N_7467,N_4542,N_5448);
or U7468 (N_7468,N_4928,N_5159);
nand U7469 (N_7469,N_4699,N_5455);
nor U7470 (N_7470,N_4503,N_5978);
nand U7471 (N_7471,N_4873,N_5155);
nor U7472 (N_7472,N_5254,N_4896);
xor U7473 (N_7473,N_5712,N_5187);
nand U7474 (N_7474,N_5883,N_5233);
and U7475 (N_7475,N_5929,N_4898);
nand U7476 (N_7476,N_5135,N_4801);
nand U7477 (N_7477,N_4607,N_4993);
nand U7478 (N_7478,N_5553,N_5399);
or U7479 (N_7479,N_4778,N_5238);
nand U7480 (N_7480,N_5927,N_5429);
nor U7481 (N_7481,N_4690,N_4796);
and U7482 (N_7482,N_5083,N_4793);
xnor U7483 (N_7483,N_4920,N_5109);
and U7484 (N_7484,N_4544,N_5037);
xor U7485 (N_7485,N_4649,N_4840);
nand U7486 (N_7486,N_4904,N_4697);
nand U7487 (N_7487,N_4558,N_5559);
xnor U7488 (N_7488,N_5499,N_5702);
nand U7489 (N_7489,N_4615,N_4568);
or U7490 (N_7490,N_4833,N_5378);
and U7491 (N_7491,N_4972,N_5466);
and U7492 (N_7492,N_5839,N_5883);
xnor U7493 (N_7493,N_4927,N_4745);
nand U7494 (N_7494,N_4823,N_4794);
and U7495 (N_7495,N_4684,N_5462);
xnor U7496 (N_7496,N_5748,N_5638);
and U7497 (N_7497,N_5258,N_4749);
nor U7498 (N_7498,N_5902,N_5578);
and U7499 (N_7499,N_5575,N_5567);
nand U7500 (N_7500,N_6263,N_7305);
xnor U7501 (N_7501,N_6573,N_6184);
or U7502 (N_7502,N_6260,N_6160);
nand U7503 (N_7503,N_6781,N_7453);
nor U7504 (N_7504,N_7312,N_6509);
xnor U7505 (N_7505,N_7205,N_6652);
and U7506 (N_7506,N_6982,N_6090);
nor U7507 (N_7507,N_6758,N_7058);
or U7508 (N_7508,N_7252,N_6675);
or U7509 (N_7509,N_6516,N_6695);
or U7510 (N_7510,N_6454,N_6269);
xor U7511 (N_7511,N_6512,N_7237);
xnor U7512 (N_7512,N_6299,N_7286);
nand U7513 (N_7513,N_7056,N_6570);
nand U7514 (N_7514,N_6693,N_6863);
nand U7515 (N_7515,N_7002,N_7417);
and U7516 (N_7516,N_7333,N_7410);
nand U7517 (N_7517,N_6772,N_7052);
or U7518 (N_7518,N_6705,N_7262);
xor U7519 (N_7519,N_7368,N_6368);
xnor U7520 (N_7520,N_6644,N_6403);
nor U7521 (N_7521,N_6195,N_6285);
nor U7522 (N_7522,N_7078,N_6432);
nor U7523 (N_7523,N_6942,N_6922);
nand U7524 (N_7524,N_7126,N_6630);
xnor U7525 (N_7525,N_6120,N_6887);
nor U7526 (N_7526,N_6629,N_7362);
or U7527 (N_7527,N_6397,N_6335);
nand U7528 (N_7528,N_6989,N_6823);
nand U7529 (N_7529,N_7353,N_6882);
nor U7530 (N_7530,N_6796,N_7354);
nand U7531 (N_7531,N_6498,N_6464);
nor U7532 (N_7532,N_6200,N_6606);
xor U7533 (N_7533,N_6838,N_6615);
nor U7534 (N_7534,N_6961,N_7068);
nor U7535 (N_7535,N_6717,N_6788);
and U7536 (N_7536,N_6850,N_7287);
or U7537 (N_7537,N_6411,N_6480);
nor U7538 (N_7538,N_6847,N_6142);
xnor U7539 (N_7539,N_6429,N_6848);
or U7540 (N_7540,N_7090,N_7170);
xor U7541 (N_7541,N_6414,N_6499);
nor U7542 (N_7542,N_6144,N_6814);
xor U7543 (N_7543,N_6618,N_7399);
nand U7544 (N_7544,N_6953,N_6459);
nand U7545 (N_7545,N_6580,N_6568);
nand U7546 (N_7546,N_7080,N_6928);
and U7547 (N_7547,N_6486,N_6474);
and U7548 (N_7548,N_6558,N_7440);
or U7549 (N_7549,N_7036,N_6751);
nor U7550 (N_7550,N_6321,N_6510);
and U7551 (N_7551,N_6654,N_6956);
or U7552 (N_7552,N_6380,N_6344);
nor U7553 (N_7553,N_6419,N_6258);
nand U7554 (N_7554,N_6778,N_6291);
nor U7555 (N_7555,N_7495,N_7418);
xor U7556 (N_7556,N_7271,N_6867);
nand U7557 (N_7557,N_7427,N_7109);
xor U7558 (N_7558,N_7321,N_7269);
nand U7559 (N_7559,N_6387,N_6314);
and U7560 (N_7560,N_6378,N_6660);
and U7561 (N_7561,N_6213,N_6614);
xnor U7562 (N_7562,N_7493,N_7363);
and U7563 (N_7563,N_6275,N_6806);
nor U7564 (N_7564,N_6991,N_6050);
xor U7565 (N_7565,N_6721,N_6117);
or U7566 (N_7566,N_6186,N_7101);
xnor U7567 (N_7567,N_6697,N_6044);
and U7568 (N_7568,N_7055,N_6755);
nor U7569 (N_7569,N_6904,N_7226);
nor U7570 (N_7570,N_6469,N_7290);
or U7571 (N_7571,N_6312,N_6185);
xnor U7572 (N_7572,N_6390,N_6409);
or U7573 (N_7573,N_6552,N_6119);
nor U7574 (N_7574,N_7185,N_7326);
nand U7575 (N_7575,N_7412,N_6156);
nor U7576 (N_7576,N_6106,N_6007);
nor U7577 (N_7577,N_7172,N_6797);
nor U7578 (N_7578,N_7367,N_6651);
and U7579 (N_7579,N_7050,N_6364);
nand U7580 (N_7580,N_6140,N_7190);
xor U7581 (N_7581,N_6954,N_7065);
nand U7582 (N_7582,N_6886,N_6520);
nand U7583 (N_7583,N_6218,N_6040);
xnor U7584 (N_7584,N_6227,N_6794);
xnor U7585 (N_7585,N_7432,N_6866);
nand U7586 (N_7586,N_7365,N_6791);
and U7587 (N_7587,N_7415,N_6501);
and U7588 (N_7588,N_7298,N_6547);
and U7589 (N_7589,N_6889,N_7392);
nor U7590 (N_7590,N_7039,N_6496);
nor U7591 (N_7591,N_7144,N_7475);
nand U7592 (N_7592,N_6030,N_7494);
and U7593 (N_7593,N_6545,N_6827);
xnor U7594 (N_7594,N_6656,N_6821);
nor U7595 (N_7595,N_6530,N_6198);
xor U7596 (N_7596,N_7349,N_6853);
nor U7597 (N_7597,N_6650,N_6912);
nand U7598 (N_7598,N_6988,N_7281);
nor U7599 (N_7599,N_7132,N_6241);
and U7600 (N_7600,N_7469,N_7441);
xor U7601 (N_7601,N_6825,N_7238);
or U7602 (N_7602,N_6097,N_7089);
nor U7603 (N_7603,N_6233,N_7169);
and U7604 (N_7604,N_7084,N_6094);
nor U7605 (N_7605,N_6288,N_6899);
nor U7606 (N_7606,N_6465,N_6808);
or U7607 (N_7607,N_7146,N_7168);
nor U7608 (N_7608,N_7316,N_7092);
and U7609 (N_7609,N_6166,N_7087);
nor U7610 (N_7610,N_7425,N_6162);
or U7611 (N_7611,N_6408,N_6016);
nor U7612 (N_7612,N_7193,N_7402);
nand U7613 (N_7613,N_6301,N_6603);
nor U7614 (N_7614,N_7008,N_7389);
xnor U7615 (N_7615,N_6715,N_6575);
nor U7616 (N_7616,N_6209,N_7187);
and U7617 (N_7617,N_6271,N_7308);
xnor U7618 (N_7618,N_6990,N_7026);
or U7619 (N_7619,N_7470,N_7260);
nor U7620 (N_7620,N_6177,N_6785);
nand U7621 (N_7621,N_7229,N_6522);
xor U7622 (N_7622,N_7433,N_6243);
nand U7623 (N_7623,N_7214,N_7018);
nor U7624 (N_7624,N_7143,N_7306);
and U7625 (N_7625,N_6687,N_6639);
or U7626 (N_7626,N_7405,N_6001);
nor U7627 (N_7627,N_7436,N_7459);
nand U7628 (N_7628,N_7227,N_6828);
and U7629 (N_7629,N_6951,N_7319);
or U7630 (N_7630,N_6784,N_6153);
nor U7631 (N_7631,N_6457,N_6586);
nor U7632 (N_7632,N_6182,N_6556);
or U7633 (N_7633,N_6625,N_7067);
nor U7634 (N_7634,N_6888,N_7166);
nand U7635 (N_7635,N_6613,N_6935);
nand U7636 (N_7636,N_7485,N_7449);
and U7637 (N_7637,N_6192,N_7247);
or U7638 (N_7638,N_6400,N_7408);
nor U7639 (N_7639,N_6957,N_7279);
xor U7640 (N_7640,N_6984,N_6497);
nor U7641 (N_7641,N_6643,N_6730);
nor U7642 (N_7642,N_6421,N_7335);
nor U7643 (N_7643,N_7243,N_6324);
and U7644 (N_7644,N_7157,N_7372);
nand U7645 (N_7645,N_6423,N_7300);
and U7646 (N_7646,N_6684,N_6566);
nor U7647 (N_7647,N_6923,N_6031);
and U7648 (N_7648,N_6065,N_7009);
and U7649 (N_7649,N_6565,N_7409);
xor U7650 (N_7650,N_6392,N_6770);
nor U7651 (N_7651,N_6217,N_6122);
nand U7652 (N_7652,N_6399,N_6608);
or U7653 (N_7653,N_6318,N_6537);
nor U7654 (N_7654,N_6444,N_6960);
nor U7655 (N_7655,N_6698,N_6374);
nand U7656 (N_7656,N_6685,N_6450);
nor U7657 (N_7657,N_6436,N_6679);
and U7658 (N_7658,N_6041,N_6925);
nand U7659 (N_7659,N_6631,N_7322);
xnor U7660 (N_7660,N_6930,N_6800);
nand U7661 (N_7661,N_6809,N_7284);
and U7662 (N_7662,N_7122,N_6190);
nand U7663 (N_7663,N_6860,N_6962);
xor U7664 (N_7664,N_6975,N_6420);
xnor U7665 (N_7665,N_6527,N_6402);
and U7666 (N_7666,N_6668,N_6810);
xnor U7667 (N_7667,N_7048,N_6289);
or U7668 (N_7668,N_7047,N_6619);
or U7669 (N_7669,N_6861,N_6495);
xor U7670 (N_7670,N_7438,N_7446);
nand U7671 (N_7671,N_7134,N_6026);
xnor U7672 (N_7672,N_6385,N_6091);
nor U7673 (N_7673,N_6014,N_7334);
xor U7674 (N_7674,N_6865,N_6560);
nor U7675 (N_7675,N_6023,N_7096);
and U7676 (N_7676,N_6169,N_7153);
or U7677 (N_7677,N_6722,N_6105);
nand U7678 (N_7678,N_6987,N_6313);
nor U7679 (N_7679,N_6264,N_6396);
nor U7680 (N_7680,N_7406,N_6920);
and U7681 (N_7681,N_7159,N_6058);
nor U7682 (N_7682,N_6536,N_6820);
xor U7683 (N_7683,N_7378,N_7171);
nand U7684 (N_7684,N_6756,N_6354);
and U7685 (N_7685,N_6736,N_6242);
or U7686 (N_7686,N_6910,N_6789);
xor U7687 (N_7687,N_7401,N_6112);
nand U7688 (N_7688,N_6085,N_6482);
xor U7689 (N_7689,N_7232,N_7258);
nand U7690 (N_7690,N_7294,N_6895);
or U7691 (N_7691,N_7288,N_6471);
or U7692 (N_7692,N_7314,N_7194);
and U7693 (N_7693,N_6587,N_7278);
nand U7694 (N_7694,N_6333,N_7221);
or U7695 (N_7695,N_7366,N_7043);
nor U7696 (N_7696,N_6008,N_7060);
nand U7697 (N_7697,N_6894,N_6326);
and U7698 (N_7698,N_6753,N_6079);
or U7699 (N_7699,N_6035,N_7376);
nor U7700 (N_7700,N_6940,N_6890);
nand U7701 (N_7701,N_6662,N_6102);
nor U7702 (N_7702,N_6529,N_7100);
and U7703 (N_7703,N_6015,N_7184);
and U7704 (N_7704,N_7424,N_7492);
xnor U7705 (N_7705,N_6308,N_7352);
nand U7706 (N_7706,N_6274,N_7098);
nand U7707 (N_7707,N_7498,N_7200);
or U7708 (N_7708,N_6857,N_6924);
or U7709 (N_7709,N_6086,N_7397);
xor U7710 (N_7710,N_6624,N_6633);
nand U7711 (N_7711,N_6148,N_6569);
xor U7712 (N_7712,N_6362,N_7370);
and U7713 (N_7713,N_7374,N_7325);
and U7714 (N_7714,N_6858,N_6401);
nor U7715 (N_7715,N_6022,N_6768);
or U7716 (N_7716,N_6971,N_7158);
nand U7717 (N_7717,N_6416,N_7398);
nand U7718 (N_7718,N_7387,N_6357);
xnor U7719 (N_7719,N_6595,N_6795);
nor U7720 (N_7720,N_7155,N_6383);
xnor U7721 (N_7721,N_7219,N_7458);
nand U7722 (N_7722,N_6173,N_6761);
xnor U7723 (N_7723,N_6124,N_6053);
or U7724 (N_7724,N_7430,N_6798);
nand U7725 (N_7725,N_6234,N_7267);
nand U7726 (N_7726,N_6902,N_6508);
nand U7727 (N_7727,N_7042,N_7347);
nand U7728 (N_7728,N_7324,N_6579);
and U7729 (N_7729,N_7484,N_6430);
or U7730 (N_7730,N_6748,N_7491);
or U7731 (N_7731,N_6208,N_7212);
nor U7732 (N_7732,N_6492,N_7123);
xor U7733 (N_7733,N_6244,N_6270);
or U7734 (N_7734,N_7094,N_7105);
xor U7735 (N_7735,N_6188,N_6726);
and U7736 (N_7736,N_7361,N_6881);
xor U7737 (N_7737,N_7463,N_7173);
nand U7738 (N_7738,N_6535,N_6371);
nor U7739 (N_7739,N_6365,N_6011);
nor U7740 (N_7740,N_6716,N_6412);
and U7741 (N_7741,N_7106,N_6159);
and U7742 (N_7742,N_7077,N_7206);
or U7743 (N_7743,N_6127,N_6750);
nand U7744 (N_7744,N_6002,N_7150);
or U7745 (N_7745,N_6245,N_7407);
and U7746 (N_7746,N_6331,N_7054);
and U7747 (N_7747,N_6210,N_7473);
nand U7748 (N_7748,N_6557,N_7391);
nor U7749 (N_7749,N_6702,N_6384);
xnor U7750 (N_7750,N_6841,N_7195);
or U7751 (N_7751,N_6948,N_7477);
xnor U7752 (N_7752,N_6178,N_7444);
nor U7753 (N_7753,N_6534,N_6605);
or U7754 (N_7754,N_7442,N_6714);
or U7755 (N_7755,N_6347,N_6804);
and U7756 (N_7756,N_7455,N_6845);
and U7757 (N_7757,N_6332,N_6191);
nor U7758 (N_7758,N_6507,N_6329);
xnor U7759 (N_7759,N_6203,N_6708);
xor U7760 (N_7760,N_6012,N_7383);
nor U7761 (N_7761,N_7480,N_6147);
and U7762 (N_7762,N_6811,N_7293);
xnor U7763 (N_7763,N_6638,N_7456);
xnor U7764 (N_7764,N_6334,N_7251);
nor U7765 (N_7765,N_6039,N_6790);
or U7766 (N_7766,N_6712,N_6749);
or U7767 (N_7767,N_6746,N_6974);
or U7768 (N_7768,N_6862,N_6303);
nand U7769 (N_7769,N_6844,N_7088);
or U7770 (N_7770,N_6546,N_7236);
xor U7771 (N_7771,N_7131,N_7142);
nand U7772 (N_7772,N_6434,N_6010);
or U7773 (N_7773,N_7420,N_7472);
and U7774 (N_7774,N_6338,N_6181);
nor U7775 (N_7775,N_6438,N_7296);
xor U7776 (N_7776,N_7192,N_6455);
nand U7777 (N_7777,N_6729,N_6513);
nor U7778 (N_7778,N_6377,N_6095);
and U7779 (N_7779,N_6123,N_6594);
and U7780 (N_7780,N_6665,N_6248);
nor U7781 (N_7781,N_6045,N_6907);
or U7782 (N_7782,N_6348,N_6817);
nand U7783 (N_7783,N_6372,N_6027);
or U7784 (N_7784,N_6916,N_7327);
xnor U7785 (N_7785,N_7255,N_7450);
nor U7786 (N_7786,N_6057,N_6009);
and U7787 (N_7787,N_7220,N_6885);
nand U7788 (N_7788,N_7075,N_6601);
and U7789 (N_7789,N_7435,N_6251);
nor U7790 (N_7790,N_7309,N_7351);
or U7791 (N_7791,N_7264,N_7299);
nand U7792 (N_7792,N_7431,N_7259);
xor U7793 (N_7793,N_6305,N_7209);
xor U7794 (N_7794,N_7315,N_7328);
or U7795 (N_7795,N_7462,N_7041);
nand U7796 (N_7796,N_6448,N_7481);
or U7797 (N_7797,N_6109,N_6164);
and U7798 (N_7798,N_6076,N_6478);
nor U7799 (N_7799,N_6143,N_7426);
and U7800 (N_7800,N_6686,N_6366);
nor U7801 (N_7801,N_6336,N_6391);
nor U7802 (N_7802,N_6253,N_6946);
xnor U7803 (N_7803,N_6875,N_6118);
nand U7804 (N_7804,N_6997,N_7489);
xnor U7805 (N_7805,N_7307,N_6533);
or U7806 (N_7806,N_7360,N_6757);
nor U7807 (N_7807,N_6637,N_7265);
or U7808 (N_7808,N_6232,N_6514);
nor U7809 (N_7809,N_7428,N_6062);
xor U7810 (N_7810,N_6723,N_6874);
nor U7811 (N_7811,N_6226,N_7464);
nor U7812 (N_7812,N_6792,N_6503);
nand U7813 (N_7813,N_6175,N_7429);
and U7814 (N_7814,N_6493,N_6970);
nand U7815 (N_7815,N_6571,N_6256);
and U7816 (N_7816,N_6539,N_7053);
nand U7817 (N_7817,N_7160,N_6060);
or U7818 (N_7818,N_7413,N_7006);
and U7819 (N_7819,N_6903,N_7276);
xnor U7820 (N_7820,N_6963,N_6891);
or U7821 (N_7821,N_7266,N_6771);
or U7822 (N_7822,N_6939,N_7046);
nor U7823 (N_7823,N_7059,N_6612);
nor U7824 (N_7824,N_6413,N_7063);
nor U7825 (N_7825,N_6355,N_6727);
xor U7826 (N_7826,N_6292,N_6082);
or U7827 (N_7827,N_6080,N_6635);
or U7828 (N_7828,N_6165,N_6311);
nand U7829 (N_7829,N_7081,N_6295);
and U7830 (N_7830,N_6944,N_6674);
or U7831 (N_7831,N_7177,N_6719);
and U7832 (N_7832,N_6277,N_7051);
nand U7833 (N_7833,N_7454,N_7274);
nand U7834 (N_7834,N_6734,N_6739);
and U7835 (N_7835,N_7019,N_6302);
nor U7836 (N_7836,N_6363,N_6135);
and U7837 (N_7837,N_6659,N_6950);
and U7838 (N_7838,N_6740,N_7437);
nand U7839 (N_7839,N_7496,N_6056);
and U7840 (N_7840,N_6913,N_6621);
or U7841 (N_7841,N_7031,N_7341);
nor U7842 (N_7842,N_7049,N_6979);
or U7843 (N_7843,N_6350,N_6004);
nand U7844 (N_7844,N_6111,N_6880);
and U7845 (N_7845,N_6054,N_7490);
nand U7846 (N_7846,N_6231,N_7057);
or U7847 (N_7847,N_6265,N_6752);
nor U7848 (N_7848,N_6460,N_6688);
and U7849 (N_7849,N_6968,N_6511);
or U7850 (N_7850,N_6024,N_6774);
nor U7851 (N_7851,N_7014,N_7117);
xor U7852 (N_7852,N_6351,N_6765);
xor U7853 (N_7853,N_6937,N_6307);
or U7854 (N_7854,N_7215,N_6819);
nor U7855 (N_7855,N_6561,N_7275);
or U7856 (N_7856,N_6491,N_6067);
xnor U7857 (N_7857,N_6196,N_7186);
nor U7858 (N_7858,N_6610,N_7384);
nand U7859 (N_7859,N_6515,N_6786);
xnor U7860 (N_7860,N_6171,N_6049);
or U7861 (N_7861,N_6290,N_6517);
nand U7862 (N_7862,N_7145,N_6699);
or U7863 (N_7863,N_6607,N_6843);
nand U7864 (N_7864,N_6223,N_6589);
or U7865 (N_7865,N_7128,N_6425);
xnor U7866 (N_7866,N_7311,N_6958);
nand U7867 (N_7867,N_7213,N_7253);
xor U7868 (N_7868,N_6107,N_7329);
and U7869 (N_7869,N_6528,N_6868);
xor U7870 (N_7870,N_7071,N_6976);
and U7871 (N_7871,N_6315,N_6361);
nor U7872 (N_7872,N_6911,N_6849);
or U7873 (N_7873,N_7246,N_6622);
nand U7874 (N_7874,N_6706,N_6405);
nor U7875 (N_7875,N_6458,N_6276);
or U7876 (N_7876,N_7460,N_7204);
nor U7877 (N_7877,N_7216,N_6576);
and U7878 (N_7878,N_6407,N_7350);
nand U7879 (N_7879,N_6918,N_6319);
or U7880 (N_7880,N_6801,N_6394);
or U7881 (N_7881,N_6461,N_6896);
nor U7882 (N_7882,N_7097,N_6246);
and U7883 (N_7883,N_7140,N_7448);
nor U7884 (N_7884,N_6667,N_6055);
xnor U7885 (N_7885,N_7165,N_7467);
and U7886 (N_7886,N_7116,N_6428);
nand U7887 (N_7887,N_6360,N_7332);
and U7888 (N_7888,N_6980,N_6871);
xnor U7889 (N_7889,N_6846,N_6006);
nor U7890 (N_7890,N_6061,N_7261);
and U7891 (N_7891,N_6297,N_6367);
or U7892 (N_7892,N_6933,N_6489);
and U7893 (N_7893,N_7111,N_6051);
xnor U7894 (N_7894,N_7000,N_6092);
and U7895 (N_7895,N_6952,N_6833);
nand U7896 (N_7896,N_7024,N_7277);
xnor U7897 (N_7897,N_6393,N_7414);
nand U7898 (N_7898,N_6658,N_6404);
xnor U7899 (N_7899,N_6449,N_6905);
or U7900 (N_7900,N_6731,N_6257);
nand U7901 (N_7901,N_7248,N_7297);
nor U7902 (N_7902,N_6852,N_7202);
or U7903 (N_7903,N_6463,N_6657);
nor U7904 (N_7904,N_7379,N_6212);
and U7905 (N_7905,N_6475,N_6627);
or U7906 (N_7906,N_7044,N_6653);
or U7907 (N_7907,N_7156,N_7241);
nand U7908 (N_7908,N_6389,N_6851);
and U7909 (N_7909,N_7218,N_6998);
or U7910 (N_7910,N_6345,N_6353);
nand U7911 (N_7911,N_7005,N_7239);
and U7912 (N_7912,N_6059,N_6128);
nor U7913 (N_7913,N_6676,N_6700);
and U7914 (N_7914,N_6115,N_6168);
or U7915 (N_7915,N_6272,N_6479);
nand U7916 (N_7916,N_6646,N_7447);
nor U7917 (N_7917,N_6069,N_7465);
nand U7918 (N_7918,N_6893,N_6818);
nor U7919 (N_7919,N_7154,N_6042);
or U7920 (N_7920,N_6926,N_6661);
and U7921 (N_7921,N_6525,N_6611);
xnor U7922 (N_7922,N_7189,N_7345);
xor U7923 (N_7923,N_6735,N_7124);
and U7924 (N_7924,N_6532,N_6793);
xor U7925 (N_7925,N_7176,N_6945);
xnor U7926 (N_7926,N_7110,N_6578);
or U7927 (N_7927,N_7061,N_6609);
nand U7928 (N_7928,N_6077,N_7240);
or U7929 (N_7929,N_7004,N_6013);
or U7930 (N_7930,N_7183,N_6211);
nor U7931 (N_7931,N_6028,N_6375);
and U7932 (N_7932,N_6839,N_6000);
nor U7933 (N_7933,N_6284,N_6519);
and U7934 (N_7934,N_6278,N_7025);
and U7935 (N_7935,N_6626,N_6078);
nor U7936 (N_7936,N_6999,N_6268);
xnor U7937 (N_7937,N_6125,N_6266);
nand U7938 (N_7938,N_6996,N_7147);
nand U7939 (N_7939,N_6538,N_7196);
nor U7940 (N_7940,N_6029,N_6395);
xor U7941 (N_7941,N_6352,N_6098);
nand U7942 (N_7942,N_6725,N_6955);
nand U7943 (N_7943,N_7268,N_7223);
nor U7944 (N_7944,N_7163,N_7069);
nor U7945 (N_7945,N_6966,N_6897);
nor U7946 (N_7946,N_6046,N_7434);
and U7947 (N_7947,N_6762,N_6099);
or U7948 (N_7948,N_6179,N_7303);
and U7949 (N_7949,N_6835,N_6878);
nand U7950 (N_7950,N_6692,N_7330);
nand U7951 (N_7951,N_6487,N_6167);
xor U7952 (N_7952,N_7076,N_6710);
nor U7953 (N_7953,N_7461,N_6711);
xor U7954 (N_7954,N_6456,N_7010);
nand U7955 (N_7955,N_6864,N_7107);
xor U7956 (N_7956,N_6373,N_6550);
xor U7957 (N_7957,N_7201,N_6322);
xnor U7958 (N_7958,N_6296,N_7029);
nor U7959 (N_7959,N_6985,N_6340);
nand U7960 (N_7960,N_6669,N_6591);
nand U7961 (N_7961,N_6604,N_6590);
or U7962 (N_7962,N_6207,N_6929);
nor U7963 (N_7963,N_6317,N_6139);
nor U7964 (N_7964,N_7452,N_6398);
nor U7965 (N_7965,N_6254,N_6807);
or U7966 (N_7966,N_6193,N_6084);
xnor U7967 (N_7967,N_7375,N_6187);
or U7968 (N_7968,N_7443,N_6154);
or U7969 (N_7969,N_6995,N_6647);
and U7970 (N_7970,N_7017,N_6540);
xnor U7971 (N_7971,N_7358,N_6504);
or U7972 (N_7972,N_7211,N_6342);
nand U7973 (N_7973,N_6328,N_7093);
nand U7974 (N_7974,N_6743,N_7033);
nor U7975 (N_7975,N_6066,N_6671);
nor U7976 (N_7976,N_6883,N_6718);
and U7977 (N_7977,N_7445,N_6453);
nand U7978 (N_7978,N_7359,N_7273);
nand U7979 (N_7979,N_7250,N_7451);
xnor U7980 (N_7980,N_6488,N_6523);
xnor U7981 (N_7981,N_6225,N_6113);
nor U7982 (N_7982,N_7181,N_7355);
or U7983 (N_7983,N_6502,N_7289);
and U7984 (N_7984,N_7331,N_7103);
nand U7985 (N_7985,N_6306,N_6673);
or U7986 (N_7986,N_6349,N_7112);
and U7987 (N_7987,N_7182,N_6145);
or U7988 (N_7988,N_7035,N_6415);
nor U7989 (N_7989,N_7070,N_6634);
xnor U7990 (N_7990,N_6327,N_6931);
xnor U7991 (N_7991,N_6019,N_7479);
or U7992 (N_7992,N_6677,N_6442);
nand U7993 (N_7993,N_7283,N_6994);
and U7994 (N_7994,N_6047,N_6898);
or U7995 (N_7995,N_6494,N_6096);
and U7996 (N_7996,N_6856,N_6252);
xor U7997 (N_7997,N_7400,N_7476);
nor U7998 (N_7998,N_6678,N_7377);
or U7999 (N_7999,N_7272,N_7235);
or U8000 (N_8000,N_6737,N_6551);
and U8001 (N_8001,N_7021,N_6172);
or U8002 (N_8002,N_7313,N_6909);
nand U8003 (N_8003,N_6205,N_6577);
nand U8004 (N_8004,N_7217,N_7118);
xor U8005 (N_8005,N_6732,N_6034);
nor U8006 (N_8006,N_6199,N_6917);
nor U8007 (N_8007,N_6616,N_6541);
xor U8008 (N_8008,N_7073,N_7161);
and U8009 (N_8009,N_6183,N_6690);
and U8010 (N_8010,N_6766,N_7032);
nand U8011 (N_8011,N_6132,N_6215);
xor U8012 (N_8012,N_6572,N_6379);
nand U8013 (N_8013,N_6206,N_6703);
nor U8014 (N_8014,N_6287,N_6033);
or U8015 (N_8015,N_7136,N_6549);
nand U8016 (N_8016,N_6131,N_6236);
or U8017 (N_8017,N_7208,N_6418);
nand U8018 (N_8018,N_6914,N_6815);
and U8019 (N_8019,N_7007,N_6564);
nand U8020 (N_8020,N_7488,N_7468);
or U8021 (N_8021,N_6531,N_6842);
nor U8022 (N_8022,N_6467,N_6741);
xor U8023 (N_8023,N_7079,N_7318);
xor U8024 (N_8024,N_6149,N_7395);
and U8025 (N_8025,N_6070,N_7139);
or U8026 (N_8026,N_6481,N_6623);
xnor U8027 (N_8027,N_6689,N_6776);
xor U8028 (N_8028,N_6599,N_6081);
and U8029 (N_8029,N_6435,N_6691);
nand U8030 (N_8030,N_6443,N_6137);
or U8031 (N_8031,N_7346,N_7127);
and U8032 (N_8032,N_7040,N_7086);
nor U8033 (N_8033,N_6642,N_7027);
nand U8034 (N_8034,N_6358,N_7231);
nand U8035 (N_8035,N_6410,N_7233);
and U8036 (N_8036,N_6900,N_6562);
or U8037 (N_8037,N_6855,N_7317);
nor U8038 (N_8038,N_6073,N_7038);
nand U8039 (N_8039,N_6204,N_6584);
nand U8040 (N_8040,N_7234,N_6422);
nand U8041 (N_8041,N_6240,N_7104);
or U8042 (N_8042,N_6943,N_6554);
nand U8043 (N_8043,N_6176,N_6052);
or U8044 (N_8044,N_7419,N_7030);
and U8045 (N_8045,N_6043,N_6466);
or U8046 (N_8046,N_6967,N_7403);
or U8047 (N_8047,N_7371,N_6018);
nor U8048 (N_8048,N_6949,N_7125);
xnor U8049 (N_8049,N_6655,N_6230);
or U8050 (N_8050,N_6104,N_6600);
nor U8051 (N_8051,N_6921,N_6663);
nand U8052 (N_8052,N_7179,N_7091);
nand U8053 (N_8053,N_6598,N_7137);
and U8054 (N_8054,N_6760,N_6174);
nand U8055 (N_8055,N_7390,N_7295);
xnor U8056 (N_8056,N_7245,N_6947);
nand U8057 (N_8057,N_7285,N_6477);
nand U8058 (N_8058,N_6282,N_7224);
xnor U8059 (N_8059,N_6720,N_7373);
nor U8060 (N_8060,N_6777,N_6802);
nor U8061 (N_8061,N_6406,N_6170);
and U8062 (N_8062,N_7225,N_6259);
nand U8063 (N_8063,N_7364,N_7003);
or U8064 (N_8064,N_6701,N_6431);
nand U8065 (N_8065,N_7152,N_6381);
or U8066 (N_8066,N_7343,N_6025);
nand U8067 (N_8067,N_6682,N_7338);
or U8068 (N_8068,N_6830,N_6472);
nor U8069 (N_8069,N_6021,N_6239);
and U8070 (N_8070,N_7337,N_7422);
nor U8071 (N_8071,N_6280,N_6037);
or U8072 (N_8072,N_6068,N_6048);
and U8073 (N_8073,N_6884,N_6518);
nor U8074 (N_8074,N_7499,N_7487);
nand U8075 (N_8075,N_6320,N_7486);
nor U8076 (N_8076,N_6202,N_6640);
xnor U8077 (N_8077,N_6965,N_6433);
nor U8078 (N_8078,N_7012,N_6892);
xnor U8079 (N_8079,N_7222,N_6873);
nor U8080 (N_8080,N_7066,N_6670);
xor U8081 (N_8081,N_6707,N_6969);
nor U8082 (N_8082,N_6075,N_6574);
xor U8083 (N_8083,N_7404,N_6837);
xnor U8084 (N_8084,N_6840,N_6088);
nand U8085 (N_8085,N_6709,N_6369);
nor U8086 (N_8086,N_6216,N_6005);
or U8087 (N_8087,N_7028,N_6704);
xor U8088 (N_8088,N_6927,N_6138);
xor U8089 (N_8089,N_6993,N_6728);
xor U8090 (N_8090,N_7175,N_7045);
and U8091 (N_8091,N_6228,N_6158);
nand U8092 (N_8092,N_6286,N_6738);
and U8093 (N_8093,N_6273,N_6992);
nor U8094 (N_8094,N_6462,N_6683);
nand U8095 (N_8095,N_6483,N_7254);
nor U8096 (N_8096,N_6473,N_6386);
nand U8097 (N_8097,N_7034,N_7013);
and U8098 (N_8098,N_7257,N_6129);
nand U8099 (N_8099,N_6110,N_6316);
or U8100 (N_8100,N_7396,N_7180);
xnor U8101 (N_8101,N_6229,N_7411);
and U8102 (N_8102,N_6831,N_6447);
xor U8103 (N_8103,N_6816,N_6593);
nor U8104 (N_8104,N_7497,N_6304);
or U8105 (N_8105,N_6445,N_6267);
xnor U8106 (N_8106,N_6754,N_6832);
nor U8107 (N_8107,N_7416,N_7301);
xor U8108 (N_8108,N_6221,N_7323);
xnor U8109 (N_8109,N_7114,N_7388);
and U8110 (N_8110,N_6908,N_7135);
and U8111 (N_8111,N_7011,N_7138);
nor U8112 (N_8112,N_6346,N_7188);
or U8113 (N_8113,N_6238,N_6973);
or U8114 (N_8114,N_6972,N_6836);
xnor U8115 (N_8115,N_7113,N_6180);
nand U8116 (N_8116,N_7198,N_6281);
or U8117 (N_8117,N_6262,N_6964);
nor U8118 (N_8118,N_6812,N_6876);
nor U8119 (N_8119,N_6093,N_6803);
or U8120 (N_8120,N_6769,N_7381);
nor U8121 (N_8121,N_6544,N_7263);
nand U8122 (N_8122,N_6764,N_6103);
nand U8123 (N_8123,N_6424,N_6426);
nor U8124 (N_8124,N_7457,N_6775);
and U8125 (N_8125,N_7304,N_6649);
or U8126 (N_8126,N_6934,N_6744);
nand U8127 (N_8127,N_6805,N_6592);
and U8128 (N_8128,N_6915,N_6247);
nand U8129 (N_8129,N_6468,N_6141);
and U8130 (N_8130,N_7471,N_6323);
nor U8131 (N_8131,N_6133,N_6901);
xor U8132 (N_8132,N_6294,N_6506);
and U8133 (N_8133,N_6108,N_7382);
and U8134 (N_8134,N_7108,N_6521);
xor U8135 (N_8135,N_7120,N_6126);
and U8136 (N_8136,N_6003,N_6427);
or U8137 (N_8137,N_6869,N_6074);
and U8138 (N_8138,N_6745,N_6696);
or U8139 (N_8139,N_7199,N_6724);
xor U8140 (N_8140,N_6330,N_6063);
nor U8141 (N_8141,N_6672,N_6747);
or U8142 (N_8142,N_6214,N_6343);
or U8143 (N_8143,N_6936,N_6780);
or U8144 (N_8144,N_7421,N_6620);
or U8145 (N_8145,N_6870,N_7072);
xor U8146 (N_8146,N_6919,N_6524);
and U8147 (N_8147,N_6388,N_6567);
nand U8148 (N_8148,N_7394,N_7129);
and U8149 (N_8149,N_6293,N_6596);
nor U8150 (N_8150,N_6136,N_6356);
nand U8151 (N_8151,N_7244,N_6938);
nand U8152 (N_8152,N_7291,N_6249);
nand U8153 (N_8153,N_6219,N_7482);
or U8154 (N_8154,N_7151,N_7242);
xnor U8155 (N_8155,N_6201,N_6382);
and U8156 (N_8156,N_6879,N_6986);
xor U8157 (N_8157,N_7174,N_7385);
and U8158 (N_8158,N_6834,N_6645);
and U8159 (N_8159,N_6485,N_6981);
xnor U8160 (N_8160,N_6829,N_7102);
and U8161 (N_8161,N_7210,N_6100);
or U8162 (N_8162,N_7310,N_7203);
nor U8163 (N_8163,N_6439,N_6452);
nor U8164 (N_8164,N_6680,N_7466);
nand U8165 (N_8165,N_6799,N_6470);
or U8166 (N_8166,N_6555,N_6543);
nor U8167 (N_8167,N_7074,N_7228);
or U8168 (N_8168,N_6451,N_6150);
nor U8169 (N_8169,N_6681,N_6261);
xor U8170 (N_8170,N_7357,N_6636);
or U8171 (N_8171,N_7148,N_6114);
nand U8172 (N_8172,N_7478,N_7121);
xor U8173 (N_8173,N_6283,N_7167);
or U8174 (N_8174,N_6759,N_6255);
nand U8175 (N_8175,N_6032,N_7022);
nand U8176 (N_8176,N_6983,N_6309);
nor U8177 (N_8177,N_6742,N_6977);
xnor U8178 (N_8178,N_7099,N_7342);
xor U8179 (N_8179,N_7474,N_6146);
nor U8180 (N_8180,N_7082,N_6089);
nor U8181 (N_8181,N_6563,N_7119);
nand U8182 (N_8182,N_7340,N_6163);
xor U8183 (N_8183,N_6341,N_7023);
nor U8184 (N_8184,N_6664,N_6194);
nand U8185 (N_8185,N_6542,N_6582);
and U8186 (N_8186,N_7141,N_6130);
nand U8187 (N_8187,N_6222,N_7483);
xnor U8188 (N_8188,N_6476,N_6859);
nor U8189 (N_8189,N_6121,N_7083);
nor U8190 (N_8190,N_6713,N_6822);
nand U8191 (N_8191,N_6036,N_7302);
nor U8192 (N_8192,N_7339,N_6941);
xor U8193 (N_8193,N_7282,N_7149);
or U8194 (N_8194,N_6441,N_6484);
nor U8195 (N_8195,N_6197,N_6505);
xnor U8196 (N_8196,N_6083,N_7020);
nor U8197 (N_8197,N_6161,N_7178);
or U8198 (N_8198,N_6157,N_6339);
xor U8199 (N_8199,N_6824,N_6583);
nor U8200 (N_8200,N_6250,N_6906);
nor U8201 (N_8201,N_6101,N_7270);
nand U8202 (N_8202,N_6628,N_7369);
nor U8203 (N_8203,N_6490,N_6826);
and U8204 (N_8204,N_6155,N_7037);
or U8205 (N_8205,N_6134,N_6548);
nor U8206 (N_8206,N_6733,N_6151);
nor U8207 (N_8207,N_6632,N_6666);
xor U8208 (N_8208,N_6087,N_6526);
nor U8209 (N_8209,N_6779,N_7386);
nor U8210 (N_8210,N_6559,N_6189);
or U8211 (N_8211,N_7336,N_7095);
and U8212 (N_8212,N_6588,N_6782);
and U8213 (N_8213,N_6116,N_6767);
nand U8214 (N_8214,N_6813,N_7230);
nor U8215 (N_8215,N_6440,N_6298);
nand U8216 (N_8216,N_7292,N_6585);
nand U8217 (N_8217,N_7115,N_6932);
nor U8218 (N_8218,N_6978,N_6872);
nand U8219 (N_8219,N_6017,N_6959);
nor U8220 (N_8220,N_7164,N_6854);
nor U8221 (N_8221,N_6072,N_6300);
or U8222 (N_8222,N_6038,N_6641);
nand U8223 (N_8223,N_6763,N_6581);
xor U8224 (N_8224,N_7356,N_6617);
and U8225 (N_8225,N_7015,N_6224);
nor U8226 (N_8226,N_6220,N_7085);
xnor U8227 (N_8227,N_6648,N_6020);
xnor U8228 (N_8228,N_7320,N_6597);
nand U8229 (N_8229,N_6310,N_7423);
xnor U8230 (N_8230,N_6446,N_7348);
or U8231 (N_8231,N_6773,N_7393);
and U8232 (N_8232,N_6877,N_7380);
nand U8233 (N_8233,N_7062,N_6064);
and U8234 (N_8234,N_7280,N_6325);
and U8235 (N_8235,N_6553,N_6417);
nor U8236 (N_8236,N_6237,N_6370);
or U8237 (N_8237,N_6783,N_6152);
nand U8238 (N_8238,N_7001,N_6437);
and U8239 (N_8239,N_7256,N_6235);
nor U8240 (N_8240,N_7133,N_7191);
nand U8241 (N_8241,N_6359,N_6602);
nand U8242 (N_8242,N_7249,N_7064);
nor U8243 (N_8243,N_6337,N_6279);
and U8244 (N_8244,N_7016,N_7130);
nand U8245 (N_8245,N_7162,N_6376);
xnor U8246 (N_8246,N_6500,N_6694);
nor U8247 (N_8247,N_6787,N_7439);
xor U8248 (N_8248,N_7344,N_6071);
xor U8249 (N_8249,N_7207,N_7197);
or U8250 (N_8250,N_7428,N_6432);
or U8251 (N_8251,N_6725,N_6662);
nor U8252 (N_8252,N_6695,N_6002);
xnor U8253 (N_8253,N_6106,N_6687);
nor U8254 (N_8254,N_6945,N_6394);
nand U8255 (N_8255,N_7171,N_7462);
nand U8256 (N_8256,N_6125,N_6008);
or U8257 (N_8257,N_7442,N_6529);
xnor U8258 (N_8258,N_6922,N_6644);
nor U8259 (N_8259,N_7381,N_7489);
or U8260 (N_8260,N_7316,N_6276);
nor U8261 (N_8261,N_6788,N_7466);
nand U8262 (N_8262,N_6769,N_7003);
nand U8263 (N_8263,N_7393,N_6155);
nor U8264 (N_8264,N_7045,N_6500);
and U8265 (N_8265,N_7313,N_6678);
xor U8266 (N_8266,N_7429,N_7406);
xor U8267 (N_8267,N_7016,N_6093);
nor U8268 (N_8268,N_7429,N_6806);
xnor U8269 (N_8269,N_6357,N_7308);
xor U8270 (N_8270,N_7448,N_6242);
or U8271 (N_8271,N_6199,N_6373);
or U8272 (N_8272,N_6252,N_6775);
nor U8273 (N_8273,N_6921,N_6456);
nand U8274 (N_8274,N_6941,N_6268);
or U8275 (N_8275,N_6551,N_6553);
nand U8276 (N_8276,N_6738,N_7283);
nor U8277 (N_8277,N_6253,N_6920);
and U8278 (N_8278,N_6939,N_6608);
nand U8279 (N_8279,N_7344,N_7347);
nand U8280 (N_8280,N_6432,N_6699);
nor U8281 (N_8281,N_7026,N_6360);
nor U8282 (N_8282,N_6772,N_6599);
xor U8283 (N_8283,N_6819,N_6128);
or U8284 (N_8284,N_6528,N_6658);
xor U8285 (N_8285,N_7378,N_6398);
nand U8286 (N_8286,N_7249,N_6608);
and U8287 (N_8287,N_6743,N_7089);
and U8288 (N_8288,N_6555,N_6220);
and U8289 (N_8289,N_6285,N_6789);
nand U8290 (N_8290,N_6316,N_6852);
nand U8291 (N_8291,N_6041,N_6222);
nand U8292 (N_8292,N_6397,N_6180);
nor U8293 (N_8293,N_6073,N_7255);
nand U8294 (N_8294,N_6077,N_6370);
nor U8295 (N_8295,N_6349,N_6064);
xnor U8296 (N_8296,N_6309,N_6838);
nand U8297 (N_8297,N_7121,N_6094);
xnor U8298 (N_8298,N_6052,N_6852);
xor U8299 (N_8299,N_6738,N_6182);
or U8300 (N_8300,N_6633,N_7053);
nand U8301 (N_8301,N_6433,N_6394);
xor U8302 (N_8302,N_7485,N_6901);
or U8303 (N_8303,N_6329,N_6851);
nor U8304 (N_8304,N_7225,N_7469);
nand U8305 (N_8305,N_7481,N_7200);
xnor U8306 (N_8306,N_7492,N_6241);
or U8307 (N_8307,N_6267,N_6541);
xor U8308 (N_8308,N_6553,N_7151);
or U8309 (N_8309,N_6270,N_6825);
or U8310 (N_8310,N_7038,N_7207);
or U8311 (N_8311,N_7215,N_6741);
or U8312 (N_8312,N_6622,N_6742);
nand U8313 (N_8313,N_6595,N_6322);
nand U8314 (N_8314,N_6191,N_6371);
nor U8315 (N_8315,N_6959,N_6462);
nand U8316 (N_8316,N_6397,N_6538);
nor U8317 (N_8317,N_6269,N_7369);
nand U8318 (N_8318,N_6359,N_7172);
or U8319 (N_8319,N_6083,N_7480);
nor U8320 (N_8320,N_6715,N_7196);
nand U8321 (N_8321,N_6963,N_6407);
nor U8322 (N_8322,N_6274,N_6233);
nor U8323 (N_8323,N_7496,N_6816);
xnor U8324 (N_8324,N_7243,N_6893);
nand U8325 (N_8325,N_7362,N_7346);
and U8326 (N_8326,N_6756,N_6389);
and U8327 (N_8327,N_6745,N_6359);
nand U8328 (N_8328,N_6427,N_7244);
nand U8329 (N_8329,N_7473,N_7427);
xor U8330 (N_8330,N_6205,N_7030);
or U8331 (N_8331,N_6545,N_7153);
nand U8332 (N_8332,N_6026,N_7268);
xor U8333 (N_8333,N_6845,N_7324);
xnor U8334 (N_8334,N_7065,N_6173);
nor U8335 (N_8335,N_6977,N_6495);
xnor U8336 (N_8336,N_6755,N_6342);
nor U8337 (N_8337,N_7296,N_7083);
and U8338 (N_8338,N_6517,N_6371);
nand U8339 (N_8339,N_6538,N_7366);
xor U8340 (N_8340,N_6392,N_7107);
nor U8341 (N_8341,N_6348,N_7448);
and U8342 (N_8342,N_7158,N_6607);
or U8343 (N_8343,N_6139,N_6786);
nor U8344 (N_8344,N_7113,N_6601);
xor U8345 (N_8345,N_6095,N_7158);
or U8346 (N_8346,N_6865,N_6648);
and U8347 (N_8347,N_7078,N_6077);
nor U8348 (N_8348,N_7099,N_6161);
and U8349 (N_8349,N_7445,N_6282);
xnor U8350 (N_8350,N_6490,N_6773);
nand U8351 (N_8351,N_6098,N_6318);
or U8352 (N_8352,N_6149,N_7045);
and U8353 (N_8353,N_7317,N_6588);
nand U8354 (N_8354,N_6788,N_7080);
or U8355 (N_8355,N_6935,N_7318);
nand U8356 (N_8356,N_6565,N_6290);
xor U8357 (N_8357,N_6658,N_6023);
nand U8358 (N_8358,N_6988,N_6048);
nor U8359 (N_8359,N_6201,N_6747);
xor U8360 (N_8360,N_7009,N_6408);
and U8361 (N_8361,N_6243,N_6016);
xnor U8362 (N_8362,N_6999,N_6342);
nor U8363 (N_8363,N_6305,N_6582);
or U8364 (N_8364,N_6459,N_7108);
nor U8365 (N_8365,N_7387,N_7254);
nor U8366 (N_8366,N_6356,N_7171);
and U8367 (N_8367,N_7189,N_6524);
nand U8368 (N_8368,N_6401,N_6899);
nand U8369 (N_8369,N_7199,N_7039);
nand U8370 (N_8370,N_7036,N_6992);
nor U8371 (N_8371,N_6248,N_6046);
or U8372 (N_8372,N_6865,N_7317);
xor U8373 (N_8373,N_6436,N_6536);
and U8374 (N_8374,N_6229,N_6290);
xnor U8375 (N_8375,N_6419,N_7025);
and U8376 (N_8376,N_6541,N_7040);
or U8377 (N_8377,N_6054,N_7082);
xnor U8378 (N_8378,N_6427,N_7305);
and U8379 (N_8379,N_7071,N_6329);
xor U8380 (N_8380,N_7404,N_6433);
nand U8381 (N_8381,N_6441,N_7039);
or U8382 (N_8382,N_7086,N_7107);
xor U8383 (N_8383,N_6330,N_7117);
or U8384 (N_8384,N_6027,N_6045);
or U8385 (N_8385,N_6071,N_6070);
nand U8386 (N_8386,N_6651,N_6763);
nor U8387 (N_8387,N_7381,N_6547);
xor U8388 (N_8388,N_7215,N_6470);
xor U8389 (N_8389,N_7202,N_7300);
or U8390 (N_8390,N_6526,N_7370);
nand U8391 (N_8391,N_6191,N_6085);
nor U8392 (N_8392,N_6650,N_6644);
and U8393 (N_8393,N_6471,N_6541);
or U8394 (N_8394,N_7197,N_7292);
or U8395 (N_8395,N_7172,N_6081);
nor U8396 (N_8396,N_6050,N_6378);
nand U8397 (N_8397,N_7261,N_6370);
nand U8398 (N_8398,N_6229,N_6575);
nand U8399 (N_8399,N_6084,N_6393);
and U8400 (N_8400,N_7463,N_7334);
nand U8401 (N_8401,N_6551,N_6182);
nand U8402 (N_8402,N_6647,N_6520);
or U8403 (N_8403,N_7130,N_6235);
nand U8404 (N_8404,N_6251,N_7142);
nor U8405 (N_8405,N_7443,N_6738);
nor U8406 (N_8406,N_6964,N_7448);
or U8407 (N_8407,N_6313,N_6785);
nor U8408 (N_8408,N_6139,N_7492);
or U8409 (N_8409,N_7455,N_6956);
and U8410 (N_8410,N_6230,N_7095);
or U8411 (N_8411,N_6227,N_6065);
nor U8412 (N_8412,N_6485,N_7248);
or U8413 (N_8413,N_6284,N_6614);
nor U8414 (N_8414,N_6089,N_6191);
nand U8415 (N_8415,N_6932,N_6020);
xnor U8416 (N_8416,N_6444,N_6633);
and U8417 (N_8417,N_6861,N_7343);
nor U8418 (N_8418,N_6018,N_7093);
nand U8419 (N_8419,N_7016,N_7487);
and U8420 (N_8420,N_7423,N_6004);
nand U8421 (N_8421,N_7071,N_7422);
xnor U8422 (N_8422,N_6028,N_6448);
nand U8423 (N_8423,N_7032,N_7064);
nor U8424 (N_8424,N_7333,N_6412);
or U8425 (N_8425,N_7139,N_7452);
xnor U8426 (N_8426,N_6603,N_7174);
or U8427 (N_8427,N_6080,N_7375);
nor U8428 (N_8428,N_6808,N_7441);
nor U8429 (N_8429,N_6409,N_7128);
nand U8430 (N_8430,N_6178,N_7098);
nor U8431 (N_8431,N_7191,N_6017);
nand U8432 (N_8432,N_6634,N_6973);
xor U8433 (N_8433,N_6566,N_6944);
nand U8434 (N_8434,N_6592,N_6135);
nor U8435 (N_8435,N_6100,N_6306);
xor U8436 (N_8436,N_7484,N_6612);
nand U8437 (N_8437,N_6950,N_6279);
and U8438 (N_8438,N_6503,N_6084);
nor U8439 (N_8439,N_7303,N_7008);
or U8440 (N_8440,N_6944,N_6891);
nor U8441 (N_8441,N_6211,N_6459);
nand U8442 (N_8442,N_7415,N_6217);
and U8443 (N_8443,N_6575,N_7232);
or U8444 (N_8444,N_6283,N_6233);
xnor U8445 (N_8445,N_6943,N_7195);
nor U8446 (N_8446,N_6069,N_6930);
xor U8447 (N_8447,N_6289,N_7354);
nand U8448 (N_8448,N_6102,N_6131);
nor U8449 (N_8449,N_6665,N_6510);
nand U8450 (N_8450,N_6134,N_7413);
nor U8451 (N_8451,N_6770,N_6355);
or U8452 (N_8452,N_6202,N_7415);
xor U8453 (N_8453,N_6395,N_6377);
or U8454 (N_8454,N_7118,N_6548);
nand U8455 (N_8455,N_6992,N_6335);
xor U8456 (N_8456,N_7220,N_7152);
xor U8457 (N_8457,N_7182,N_7270);
or U8458 (N_8458,N_6342,N_6006);
xnor U8459 (N_8459,N_7147,N_7438);
or U8460 (N_8460,N_6802,N_6089);
or U8461 (N_8461,N_6157,N_6699);
nand U8462 (N_8462,N_6980,N_6839);
xnor U8463 (N_8463,N_6712,N_6099);
xnor U8464 (N_8464,N_7346,N_6733);
xnor U8465 (N_8465,N_6670,N_7052);
nand U8466 (N_8466,N_6546,N_7053);
nor U8467 (N_8467,N_6138,N_6115);
and U8468 (N_8468,N_6718,N_6954);
nand U8469 (N_8469,N_7381,N_6048);
or U8470 (N_8470,N_6851,N_6067);
nand U8471 (N_8471,N_6724,N_6883);
and U8472 (N_8472,N_6426,N_6165);
or U8473 (N_8473,N_6034,N_6024);
nor U8474 (N_8474,N_6497,N_6075);
or U8475 (N_8475,N_6907,N_6801);
nor U8476 (N_8476,N_7237,N_6766);
or U8477 (N_8477,N_6276,N_6784);
nand U8478 (N_8478,N_6906,N_6573);
nand U8479 (N_8479,N_6738,N_6264);
xor U8480 (N_8480,N_6745,N_7342);
nand U8481 (N_8481,N_7327,N_6821);
nor U8482 (N_8482,N_6201,N_6323);
or U8483 (N_8483,N_7276,N_6026);
and U8484 (N_8484,N_6170,N_7026);
xor U8485 (N_8485,N_7139,N_7106);
xnor U8486 (N_8486,N_6787,N_7249);
or U8487 (N_8487,N_6975,N_6526);
xor U8488 (N_8488,N_7061,N_6907);
nor U8489 (N_8489,N_6189,N_6164);
or U8490 (N_8490,N_7448,N_6907);
or U8491 (N_8491,N_6193,N_6536);
or U8492 (N_8492,N_6011,N_6359);
xor U8493 (N_8493,N_7183,N_6794);
nand U8494 (N_8494,N_6495,N_7373);
and U8495 (N_8495,N_6412,N_6212);
or U8496 (N_8496,N_6781,N_7359);
or U8497 (N_8497,N_6791,N_7462);
nor U8498 (N_8498,N_6783,N_6601);
nor U8499 (N_8499,N_6630,N_7235);
nor U8500 (N_8500,N_7315,N_6042);
and U8501 (N_8501,N_6209,N_6185);
xnor U8502 (N_8502,N_6489,N_6434);
and U8503 (N_8503,N_6514,N_6834);
and U8504 (N_8504,N_7311,N_6257);
nor U8505 (N_8505,N_6350,N_6982);
nor U8506 (N_8506,N_7219,N_6040);
or U8507 (N_8507,N_6027,N_6066);
and U8508 (N_8508,N_6875,N_6293);
nor U8509 (N_8509,N_7268,N_7104);
or U8510 (N_8510,N_7374,N_6533);
xor U8511 (N_8511,N_6006,N_7162);
nand U8512 (N_8512,N_6713,N_7157);
and U8513 (N_8513,N_7423,N_6474);
nor U8514 (N_8514,N_6450,N_6494);
or U8515 (N_8515,N_6682,N_6612);
xnor U8516 (N_8516,N_6106,N_7201);
or U8517 (N_8517,N_6819,N_7149);
or U8518 (N_8518,N_6564,N_6322);
or U8519 (N_8519,N_6614,N_6781);
and U8520 (N_8520,N_6445,N_6807);
or U8521 (N_8521,N_6185,N_6085);
xor U8522 (N_8522,N_7470,N_6750);
nor U8523 (N_8523,N_6514,N_7461);
or U8524 (N_8524,N_6105,N_7382);
nor U8525 (N_8525,N_7032,N_7179);
or U8526 (N_8526,N_6682,N_6485);
nand U8527 (N_8527,N_6764,N_7076);
nand U8528 (N_8528,N_7064,N_7086);
and U8529 (N_8529,N_6665,N_7115);
nand U8530 (N_8530,N_6311,N_7318);
or U8531 (N_8531,N_6019,N_6585);
nand U8532 (N_8532,N_6961,N_6053);
or U8533 (N_8533,N_6590,N_6110);
xnor U8534 (N_8534,N_7384,N_6695);
xnor U8535 (N_8535,N_7218,N_6908);
xor U8536 (N_8536,N_7108,N_7308);
xnor U8537 (N_8537,N_6875,N_6879);
nand U8538 (N_8538,N_6475,N_6031);
and U8539 (N_8539,N_6129,N_6739);
nor U8540 (N_8540,N_7007,N_7119);
and U8541 (N_8541,N_7162,N_7405);
or U8542 (N_8542,N_6730,N_7010);
and U8543 (N_8543,N_6264,N_6294);
and U8544 (N_8544,N_6103,N_6761);
or U8545 (N_8545,N_6198,N_6597);
and U8546 (N_8546,N_7383,N_6279);
nand U8547 (N_8547,N_6876,N_6280);
xor U8548 (N_8548,N_6974,N_7278);
nand U8549 (N_8549,N_6829,N_6987);
xor U8550 (N_8550,N_6954,N_6534);
xor U8551 (N_8551,N_7343,N_6047);
xor U8552 (N_8552,N_7028,N_6035);
and U8553 (N_8553,N_7498,N_6685);
nor U8554 (N_8554,N_6264,N_7296);
nor U8555 (N_8555,N_7292,N_6168);
and U8556 (N_8556,N_7471,N_6386);
and U8557 (N_8557,N_7274,N_6563);
nor U8558 (N_8558,N_7372,N_7304);
xnor U8559 (N_8559,N_7475,N_6300);
nor U8560 (N_8560,N_7425,N_6115);
or U8561 (N_8561,N_6556,N_6424);
nor U8562 (N_8562,N_7281,N_6044);
xnor U8563 (N_8563,N_6865,N_6104);
and U8564 (N_8564,N_6764,N_6613);
nand U8565 (N_8565,N_6204,N_6730);
or U8566 (N_8566,N_6873,N_7342);
and U8567 (N_8567,N_6499,N_6586);
nand U8568 (N_8568,N_6923,N_6808);
and U8569 (N_8569,N_7476,N_6101);
xor U8570 (N_8570,N_6341,N_7348);
nand U8571 (N_8571,N_6559,N_6930);
nand U8572 (N_8572,N_7328,N_6263);
nand U8573 (N_8573,N_7213,N_6761);
nand U8574 (N_8574,N_6295,N_6669);
and U8575 (N_8575,N_6516,N_6160);
or U8576 (N_8576,N_6961,N_6464);
nand U8577 (N_8577,N_6781,N_6881);
xor U8578 (N_8578,N_7184,N_6874);
nor U8579 (N_8579,N_6218,N_6473);
nor U8580 (N_8580,N_6547,N_6717);
and U8581 (N_8581,N_6162,N_6585);
or U8582 (N_8582,N_7077,N_6067);
nor U8583 (N_8583,N_6732,N_6462);
or U8584 (N_8584,N_6909,N_7435);
nor U8585 (N_8585,N_6708,N_6430);
xor U8586 (N_8586,N_6215,N_6377);
nor U8587 (N_8587,N_6260,N_7423);
and U8588 (N_8588,N_7225,N_6176);
nor U8589 (N_8589,N_6367,N_6690);
nand U8590 (N_8590,N_7434,N_6341);
and U8591 (N_8591,N_6603,N_7151);
and U8592 (N_8592,N_6152,N_6005);
xnor U8593 (N_8593,N_6835,N_7323);
and U8594 (N_8594,N_6814,N_6193);
or U8595 (N_8595,N_7282,N_7322);
nor U8596 (N_8596,N_6477,N_7080);
or U8597 (N_8597,N_6757,N_7131);
xor U8598 (N_8598,N_7021,N_6839);
nor U8599 (N_8599,N_6946,N_6093);
or U8600 (N_8600,N_6235,N_6081);
and U8601 (N_8601,N_6900,N_6341);
and U8602 (N_8602,N_7046,N_7428);
and U8603 (N_8603,N_6179,N_6529);
or U8604 (N_8604,N_6469,N_6731);
and U8605 (N_8605,N_7264,N_6851);
nand U8606 (N_8606,N_7130,N_6405);
or U8607 (N_8607,N_6785,N_6021);
nor U8608 (N_8608,N_6275,N_6870);
or U8609 (N_8609,N_7066,N_6333);
xnor U8610 (N_8610,N_7208,N_6836);
xnor U8611 (N_8611,N_7443,N_6458);
nand U8612 (N_8612,N_6089,N_6159);
nand U8613 (N_8613,N_7005,N_6861);
nor U8614 (N_8614,N_6298,N_6532);
and U8615 (N_8615,N_6527,N_7044);
xnor U8616 (N_8616,N_6642,N_7325);
xnor U8617 (N_8617,N_6993,N_6423);
or U8618 (N_8618,N_7467,N_7368);
xnor U8619 (N_8619,N_6588,N_6614);
nand U8620 (N_8620,N_6990,N_6476);
nand U8621 (N_8621,N_6921,N_7450);
xor U8622 (N_8622,N_6270,N_7197);
xor U8623 (N_8623,N_7275,N_6720);
nor U8624 (N_8624,N_7211,N_6623);
or U8625 (N_8625,N_7155,N_7458);
or U8626 (N_8626,N_6315,N_6311);
xor U8627 (N_8627,N_6106,N_6886);
and U8628 (N_8628,N_6040,N_6874);
or U8629 (N_8629,N_7379,N_6736);
and U8630 (N_8630,N_7214,N_6474);
nor U8631 (N_8631,N_6549,N_6189);
and U8632 (N_8632,N_6500,N_6107);
nor U8633 (N_8633,N_7391,N_6051);
nor U8634 (N_8634,N_7205,N_7239);
and U8635 (N_8635,N_7292,N_6574);
and U8636 (N_8636,N_6948,N_7189);
nand U8637 (N_8637,N_6485,N_6711);
or U8638 (N_8638,N_6462,N_6764);
or U8639 (N_8639,N_7230,N_6027);
or U8640 (N_8640,N_6801,N_6921);
and U8641 (N_8641,N_6292,N_6939);
and U8642 (N_8642,N_6122,N_6691);
xor U8643 (N_8643,N_7392,N_7391);
xnor U8644 (N_8644,N_6096,N_7069);
nor U8645 (N_8645,N_7249,N_6356);
nand U8646 (N_8646,N_6825,N_6747);
and U8647 (N_8647,N_6656,N_6764);
xnor U8648 (N_8648,N_6314,N_6028);
xnor U8649 (N_8649,N_6910,N_6739);
or U8650 (N_8650,N_6328,N_6407);
nor U8651 (N_8651,N_6376,N_6403);
and U8652 (N_8652,N_6797,N_7068);
xor U8653 (N_8653,N_6560,N_6427);
or U8654 (N_8654,N_7357,N_7184);
xor U8655 (N_8655,N_7389,N_7252);
nand U8656 (N_8656,N_6638,N_6699);
and U8657 (N_8657,N_7451,N_7258);
xor U8658 (N_8658,N_7491,N_6354);
or U8659 (N_8659,N_6160,N_6137);
xor U8660 (N_8660,N_6787,N_7453);
or U8661 (N_8661,N_6029,N_6942);
xor U8662 (N_8662,N_6216,N_6436);
xor U8663 (N_8663,N_6342,N_6969);
nor U8664 (N_8664,N_7463,N_7129);
xnor U8665 (N_8665,N_7105,N_6929);
and U8666 (N_8666,N_6191,N_6094);
or U8667 (N_8667,N_6229,N_6540);
xnor U8668 (N_8668,N_7199,N_6874);
nand U8669 (N_8669,N_6927,N_6866);
nor U8670 (N_8670,N_7138,N_6554);
or U8671 (N_8671,N_6776,N_7157);
nor U8672 (N_8672,N_7234,N_6593);
nor U8673 (N_8673,N_6668,N_6667);
and U8674 (N_8674,N_7047,N_6511);
xor U8675 (N_8675,N_7239,N_6436);
nand U8676 (N_8676,N_6739,N_7437);
nand U8677 (N_8677,N_6490,N_6880);
nand U8678 (N_8678,N_6853,N_6795);
and U8679 (N_8679,N_6809,N_6684);
xor U8680 (N_8680,N_6444,N_6814);
and U8681 (N_8681,N_6217,N_7418);
and U8682 (N_8682,N_6576,N_6963);
xor U8683 (N_8683,N_7076,N_6064);
and U8684 (N_8684,N_7243,N_6867);
nor U8685 (N_8685,N_6592,N_7331);
xor U8686 (N_8686,N_7246,N_6170);
and U8687 (N_8687,N_6179,N_7366);
nand U8688 (N_8688,N_6444,N_7275);
nor U8689 (N_8689,N_6703,N_7271);
or U8690 (N_8690,N_6312,N_7236);
or U8691 (N_8691,N_7058,N_7149);
nor U8692 (N_8692,N_6392,N_6123);
nor U8693 (N_8693,N_7368,N_6010);
nor U8694 (N_8694,N_6495,N_7483);
and U8695 (N_8695,N_6807,N_6198);
or U8696 (N_8696,N_6948,N_7022);
xnor U8697 (N_8697,N_7042,N_6652);
or U8698 (N_8698,N_6238,N_6157);
nor U8699 (N_8699,N_6102,N_6229);
and U8700 (N_8700,N_7418,N_6032);
nor U8701 (N_8701,N_6314,N_6288);
nand U8702 (N_8702,N_7092,N_7486);
or U8703 (N_8703,N_6168,N_6961);
nor U8704 (N_8704,N_7435,N_6930);
xnor U8705 (N_8705,N_6166,N_7477);
or U8706 (N_8706,N_6124,N_6545);
xnor U8707 (N_8707,N_7319,N_6288);
nor U8708 (N_8708,N_7339,N_7412);
nor U8709 (N_8709,N_7482,N_6275);
xor U8710 (N_8710,N_6390,N_6888);
nor U8711 (N_8711,N_7373,N_6726);
nand U8712 (N_8712,N_7415,N_7480);
nor U8713 (N_8713,N_7466,N_6724);
or U8714 (N_8714,N_6916,N_6678);
and U8715 (N_8715,N_7021,N_6493);
nand U8716 (N_8716,N_6503,N_7284);
nor U8717 (N_8717,N_6692,N_6834);
nand U8718 (N_8718,N_6483,N_6208);
or U8719 (N_8719,N_6514,N_6552);
nor U8720 (N_8720,N_6113,N_6855);
nor U8721 (N_8721,N_7086,N_6391);
nand U8722 (N_8722,N_6070,N_6380);
or U8723 (N_8723,N_7488,N_6417);
nand U8724 (N_8724,N_7077,N_6260);
xnor U8725 (N_8725,N_6088,N_6300);
nand U8726 (N_8726,N_6808,N_7143);
xnor U8727 (N_8727,N_6161,N_7014);
or U8728 (N_8728,N_7448,N_6675);
nand U8729 (N_8729,N_6471,N_7349);
or U8730 (N_8730,N_6343,N_7354);
or U8731 (N_8731,N_6850,N_7295);
nor U8732 (N_8732,N_7130,N_6920);
nor U8733 (N_8733,N_6816,N_6603);
nand U8734 (N_8734,N_6087,N_6086);
or U8735 (N_8735,N_6165,N_6811);
nor U8736 (N_8736,N_7115,N_6370);
or U8737 (N_8737,N_6460,N_7329);
and U8738 (N_8738,N_6913,N_6588);
xor U8739 (N_8739,N_6857,N_6469);
or U8740 (N_8740,N_7119,N_6142);
nand U8741 (N_8741,N_6113,N_6667);
nand U8742 (N_8742,N_6563,N_7102);
xor U8743 (N_8743,N_6929,N_6409);
and U8744 (N_8744,N_6495,N_6656);
nor U8745 (N_8745,N_7107,N_7390);
nor U8746 (N_8746,N_6012,N_7012);
nand U8747 (N_8747,N_7419,N_7411);
nand U8748 (N_8748,N_6662,N_6557);
nand U8749 (N_8749,N_6227,N_7466);
nand U8750 (N_8750,N_6276,N_6626);
or U8751 (N_8751,N_7066,N_6242);
nor U8752 (N_8752,N_7334,N_6858);
nor U8753 (N_8753,N_6144,N_6154);
and U8754 (N_8754,N_6474,N_6147);
or U8755 (N_8755,N_7350,N_7312);
nor U8756 (N_8756,N_6826,N_6594);
and U8757 (N_8757,N_6200,N_6138);
and U8758 (N_8758,N_7058,N_6079);
xnor U8759 (N_8759,N_7328,N_7329);
nand U8760 (N_8760,N_6501,N_7150);
nor U8761 (N_8761,N_6445,N_6745);
xor U8762 (N_8762,N_6699,N_7272);
xnor U8763 (N_8763,N_7300,N_6031);
and U8764 (N_8764,N_6084,N_6551);
or U8765 (N_8765,N_7437,N_6923);
nand U8766 (N_8766,N_6506,N_6642);
nor U8767 (N_8767,N_6299,N_6568);
nand U8768 (N_8768,N_7080,N_6187);
or U8769 (N_8769,N_6169,N_6149);
or U8770 (N_8770,N_6448,N_7463);
xnor U8771 (N_8771,N_6507,N_6901);
xor U8772 (N_8772,N_7116,N_7174);
or U8773 (N_8773,N_7253,N_6531);
nand U8774 (N_8774,N_7087,N_7273);
and U8775 (N_8775,N_7102,N_6217);
xor U8776 (N_8776,N_7012,N_7403);
xor U8777 (N_8777,N_7093,N_6345);
xor U8778 (N_8778,N_6076,N_6732);
and U8779 (N_8779,N_6688,N_6837);
nor U8780 (N_8780,N_6380,N_6055);
nor U8781 (N_8781,N_7188,N_6258);
nand U8782 (N_8782,N_6424,N_6764);
or U8783 (N_8783,N_6170,N_6261);
or U8784 (N_8784,N_6793,N_7218);
and U8785 (N_8785,N_6386,N_6479);
nor U8786 (N_8786,N_6311,N_6896);
and U8787 (N_8787,N_7323,N_7196);
or U8788 (N_8788,N_6308,N_6583);
or U8789 (N_8789,N_7212,N_7379);
nand U8790 (N_8790,N_6974,N_6614);
nor U8791 (N_8791,N_7210,N_7051);
and U8792 (N_8792,N_6806,N_7209);
nor U8793 (N_8793,N_7127,N_6139);
xnor U8794 (N_8794,N_6916,N_7175);
or U8795 (N_8795,N_6273,N_6106);
nand U8796 (N_8796,N_6995,N_6634);
or U8797 (N_8797,N_6571,N_6088);
xor U8798 (N_8798,N_7063,N_7113);
nand U8799 (N_8799,N_6068,N_6279);
nor U8800 (N_8800,N_6514,N_7216);
nand U8801 (N_8801,N_7111,N_6256);
xnor U8802 (N_8802,N_6896,N_7431);
nand U8803 (N_8803,N_6116,N_7062);
nand U8804 (N_8804,N_6494,N_7248);
and U8805 (N_8805,N_6300,N_7116);
xnor U8806 (N_8806,N_7153,N_6077);
and U8807 (N_8807,N_6387,N_7053);
xor U8808 (N_8808,N_7360,N_7157);
or U8809 (N_8809,N_6495,N_6823);
or U8810 (N_8810,N_6834,N_7120);
or U8811 (N_8811,N_7460,N_6221);
nor U8812 (N_8812,N_6139,N_6289);
xnor U8813 (N_8813,N_6388,N_7256);
and U8814 (N_8814,N_6178,N_6062);
or U8815 (N_8815,N_7428,N_6486);
nor U8816 (N_8816,N_7387,N_6125);
nand U8817 (N_8817,N_6685,N_7420);
nor U8818 (N_8818,N_6407,N_7166);
nand U8819 (N_8819,N_6743,N_7150);
nand U8820 (N_8820,N_6971,N_6766);
xnor U8821 (N_8821,N_6767,N_6486);
nand U8822 (N_8822,N_6938,N_6839);
nor U8823 (N_8823,N_6991,N_6942);
xnor U8824 (N_8824,N_7054,N_6419);
nor U8825 (N_8825,N_7134,N_7272);
nor U8826 (N_8826,N_6292,N_7197);
nand U8827 (N_8827,N_7134,N_6965);
xor U8828 (N_8828,N_6633,N_6295);
and U8829 (N_8829,N_6358,N_7155);
nand U8830 (N_8830,N_6595,N_6045);
nand U8831 (N_8831,N_6472,N_6476);
xnor U8832 (N_8832,N_6344,N_6107);
and U8833 (N_8833,N_7431,N_6915);
xor U8834 (N_8834,N_6720,N_6958);
nand U8835 (N_8835,N_7287,N_6882);
nor U8836 (N_8836,N_7130,N_6864);
or U8837 (N_8837,N_6193,N_7435);
nor U8838 (N_8838,N_6534,N_6985);
or U8839 (N_8839,N_6543,N_6311);
and U8840 (N_8840,N_7295,N_7006);
nor U8841 (N_8841,N_6442,N_6494);
or U8842 (N_8842,N_7028,N_6971);
xnor U8843 (N_8843,N_6743,N_6732);
nor U8844 (N_8844,N_6751,N_7329);
and U8845 (N_8845,N_6780,N_6053);
nor U8846 (N_8846,N_6125,N_6372);
xnor U8847 (N_8847,N_6501,N_6617);
or U8848 (N_8848,N_6990,N_6117);
nand U8849 (N_8849,N_6511,N_7237);
nor U8850 (N_8850,N_7207,N_7283);
nand U8851 (N_8851,N_7375,N_6567);
nor U8852 (N_8852,N_6925,N_6369);
or U8853 (N_8853,N_7111,N_7486);
or U8854 (N_8854,N_6017,N_7471);
or U8855 (N_8855,N_6096,N_6122);
nor U8856 (N_8856,N_6299,N_6670);
nand U8857 (N_8857,N_6284,N_6220);
and U8858 (N_8858,N_7265,N_6904);
and U8859 (N_8859,N_6188,N_6172);
nor U8860 (N_8860,N_6906,N_7069);
or U8861 (N_8861,N_6559,N_6166);
nor U8862 (N_8862,N_7155,N_6730);
xor U8863 (N_8863,N_7372,N_6313);
xnor U8864 (N_8864,N_6756,N_7185);
or U8865 (N_8865,N_7392,N_6987);
nor U8866 (N_8866,N_6441,N_6156);
and U8867 (N_8867,N_6437,N_6419);
xnor U8868 (N_8868,N_7305,N_7256);
or U8869 (N_8869,N_6903,N_7437);
or U8870 (N_8870,N_7289,N_6948);
and U8871 (N_8871,N_6325,N_7372);
and U8872 (N_8872,N_6366,N_6164);
xor U8873 (N_8873,N_6233,N_6934);
nand U8874 (N_8874,N_6497,N_6041);
and U8875 (N_8875,N_6059,N_6580);
xor U8876 (N_8876,N_7408,N_7172);
and U8877 (N_8877,N_6815,N_7150);
and U8878 (N_8878,N_6235,N_6991);
nor U8879 (N_8879,N_7316,N_6198);
nor U8880 (N_8880,N_7273,N_6730);
or U8881 (N_8881,N_7376,N_7239);
xnor U8882 (N_8882,N_6511,N_6717);
xnor U8883 (N_8883,N_6465,N_6387);
nor U8884 (N_8884,N_7063,N_6847);
xor U8885 (N_8885,N_6327,N_6743);
nor U8886 (N_8886,N_6317,N_6129);
nand U8887 (N_8887,N_7184,N_6572);
or U8888 (N_8888,N_6234,N_7256);
nand U8889 (N_8889,N_6528,N_7234);
xor U8890 (N_8890,N_7438,N_6733);
and U8891 (N_8891,N_6797,N_7047);
xor U8892 (N_8892,N_6975,N_7356);
or U8893 (N_8893,N_6155,N_6490);
or U8894 (N_8894,N_7097,N_6125);
nor U8895 (N_8895,N_6059,N_7121);
and U8896 (N_8896,N_6678,N_6133);
nor U8897 (N_8897,N_7446,N_6374);
nand U8898 (N_8898,N_7101,N_7057);
and U8899 (N_8899,N_6718,N_6454);
xor U8900 (N_8900,N_6647,N_7009);
nor U8901 (N_8901,N_6515,N_7389);
xor U8902 (N_8902,N_6561,N_7005);
and U8903 (N_8903,N_6358,N_6136);
or U8904 (N_8904,N_7207,N_6248);
nand U8905 (N_8905,N_6293,N_7344);
nand U8906 (N_8906,N_7470,N_6175);
or U8907 (N_8907,N_7228,N_6734);
nand U8908 (N_8908,N_7456,N_7383);
or U8909 (N_8909,N_6449,N_6181);
and U8910 (N_8910,N_6799,N_7015);
or U8911 (N_8911,N_6170,N_6504);
or U8912 (N_8912,N_7243,N_6412);
xor U8913 (N_8913,N_6119,N_6362);
nor U8914 (N_8914,N_7144,N_6005);
nor U8915 (N_8915,N_6480,N_6629);
xor U8916 (N_8916,N_6335,N_6404);
nor U8917 (N_8917,N_7486,N_6111);
or U8918 (N_8918,N_6876,N_6972);
nand U8919 (N_8919,N_7481,N_6214);
and U8920 (N_8920,N_6526,N_6530);
nor U8921 (N_8921,N_6844,N_6372);
nor U8922 (N_8922,N_6264,N_7421);
and U8923 (N_8923,N_6726,N_7235);
nand U8924 (N_8924,N_6355,N_6293);
xnor U8925 (N_8925,N_7248,N_7414);
xor U8926 (N_8926,N_7462,N_7194);
nand U8927 (N_8927,N_7206,N_6734);
or U8928 (N_8928,N_7351,N_6619);
and U8929 (N_8929,N_6848,N_7346);
nor U8930 (N_8930,N_6903,N_6559);
xnor U8931 (N_8931,N_6673,N_7495);
nor U8932 (N_8932,N_6250,N_6939);
nand U8933 (N_8933,N_6900,N_6904);
or U8934 (N_8934,N_6714,N_7320);
xnor U8935 (N_8935,N_7202,N_7458);
or U8936 (N_8936,N_6175,N_7168);
xor U8937 (N_8937,N_7286,N_6425);
and U8938 (N_8938,N_6427,N_6607);
nand U8939 (N_8939,N_7123,N_6311);
or U8940 (N_8940,N_6927,N_7056);
nand U8941 (N_8941,N_7359,N_6528);
or U8942 (N_8942,N_7453,N_7202);
xnor U8943 (N_8943,N_6437,N_6931);
nand U8944 (N_8944,N_7216,N_6560);
and U8945 (N_8945,N_6654,N_6200);
nand U8946 (N_8946,N_6748,N_6675);
nor U8947 (N_8947,N_7322,N_7372);
xor U8948 (N_8948,N_6787,N_6140);
xor U8949 (N_8949,N_6190,N_6222);
xnor U8950 (N_8950,N_6024,N_7196);
or U8951 (N_8951,N_6329,N_6280);
nand U8952 (N_8952,N_6132,N_6931);
or U8953 (N_8953,N_6399,N_6886);
nor U8954 (N_8954,N_6161,N_6456);
and U8955 (N_8955,N_7105,N_6370);
or U8956 (N_8956,N_6418,N_6187);
nand U8957 (N_8957,N_7030,N_6404);
xnor U8958 (N_8958,N_6876,N_6925);
or U8959 (N_8959,N_6110,N_6353);
nor U8960 (N_8960,N_6061,N_7046);
or U8961 (N_8961,N_6490,N_6526);
nand U8962 (N_8962,N_7126,N_7422);
nand U8963 (N_8963,N_6379,N_7467);
nor U8964 (N_8964,N_6542,N_7362);
nor U8965 (N_8965,N_6628,N_7248);
xor U8966 (N_8966,N_7462,N_6428);
nor U8967 (N_8967,N_7384,N_7399);
or U8968 (N_8968,N_7048,N_6480);
and U8969 (N_8969,N_7134,N_6039);
or U8970 (N_8970,N_6319,N_6486);
or U8971 (N_8971,N_7015,N_6742);
nand U8972 (N_8972,N_6628,N_6556);
and U8973 (N_8973,N_6885,N_6274);
xor U8974 (N_8974,N_7064,N_6374);
and U8975 (N_8975,N_6667,N_7351);
and U8976 (N_8976,N_6284,N_6465);
xnor U8977 (N_8977,N_6781,N_6132);
xnor U8978 (N_8978,N_6212,N_6167);
nor U8979 (N_8979,N_6503,N_7092);
nand U8980 (N_8980,N_7244,N_6142);
nand U8981 (N_8981,N_6386,N_7105);
and U8982 (N_8982,N_6339,N_6917);
and U8983 (N_8983,N_7207,N_6187);
xor U8984 (N_8984,N_6915,N_6224);
nor U8985 (N_8985,N_6535,N_6651);
xor U8986 (N_8986,N_6975,N_6293);
xor U8987 (N_8987,N_7497,N_7321);
nand U8988 (N_8988,N_6421,N_6910);
nor U8989 (N_8989,N_6829,N_6211);
and U8990 (N_8990,N_6976,N_6246);
and U8991 (N_8991,N_6411,N_7379);
and U8992 (N_8992,N_7432,N_6311);
and U8993 (N_8993,N_6800,N_6610);
nand U8994 (N_8994,N_6518,N_6968);
or U8995 (N_8995,N_7363,N_7179);
nand U8996 (N_8996,N_6137,N_6521);
or U8997 (N_8997,N_6467,N_6277);
xnor U8998 (N_8998,N_7277,N_7474);
nor U8999 (N_8999,N_6859,N_6208);
nand U9000 (N_9000,N_7891,N_8029);
xnor U9001 (N_9001,N_7860,N_8685);
xor U9002 (N_9002,N_8561,N_8400);
nand U9003 (N_9003,N_7838,N_7926);
nor U9004 (N_9004,N_8449,N_7754);
xnor U9005 (N_9005,N_8057,N_8578);
nand U9006 (N_9006,N_8089,N_8211);
or U9007 (N_9007,N_7656,N_8048);
and U9008 (N_9008,N_8562,N_8762);
xor U9009 (N_9009,N_8208,N_8337);
and U9010 (N_9010,N_7861,N_7547);
xor U9011 (N_9011,N_8277,N_7577);
nand U9012 (N_9012,N_8259,N_8042);
or U9013 (N_9013,N_8328,N_8765);
nand U9014 (N_9014,N_8172,N_7956);
nor U9015 (N_9015,N_8114,N_7884);
and U9016 (N_9016,N_7742,N_8973);
xnor U9017 (N_9017,N_7998,N_8223);
nor U9018 (N_9018,N_8791,N_8509);
nand U9019 (N_9019,N_8673,N_7999);
or U9020 (N_9020,N_8885,N_8501);
xor U9021 (N_9021,N_8555,N_8644);
and U9022 (N_9022,N_8248,N_8675);
or U9023 (N_9023,N_8435,N_8087);
and U9024 (N_9024,N_7526,N_8462);
or U9025 (N_9025,N_7714,N_7992);
xnor U9026 (N_9026,N_8035,N_7532);
xnor U9027 (N_9027,N_8932,N_8626);
xor U9028 (N_9028,N_7903,N_8394);
or U9029 (N_9029,N_8471,N_7734);
and U9030 (N_9030,N_8786,N_8537);
and U9031 (N_9031,N_8752,N_8000);
or U9032 (N_9032,N_8303,N_8881);
nand U9033 (N_9033,N_8202,N_7557);
and U9034 (N_9034,N_7990,N_8733);
nand U9035 (N_9035,N_7963,N_8031);
xnor U9036 (N_9036,N_8748,N_7661);
xor U9037 (N_9037,N_8794,N_7600);
or U9038 (N_9038,N_8479,N_8192);
or U9039 (N_9039,N_8205,N_7589);
or U9040 (N_9040,N_8126,N_8313);
nor U9041 (N_9041,N_8852,N_7737);
nor U9042 (N_9042,N_8286,N_7684);
nand U9043 (N_9043,N_8961,N_7668);
nand U9044 (N_9044,N_8164,N_8056);
and U9045 (N_9045,N_8331,N_7788);
or U9046 (N_9046,N_8174,N_8522);
or U9047 (N_9047,N_8798,N_7873);
xor U9048 (N_9048,N_8054,N_7604);
xor U9049 (N_9049,N_7858,N_7978);
nor U9050 (N_9050,N_8840,N_7627);
nor U9051 (N_9051,N_8540,N_8942);
or U9052 (N_9052,N_8153,N_8834);
and U9053 (N_9053,N_7753,N_7853);
nor U9054 (N_9054,N_8472,N_7987);
and U9055 (N_9055,N_8838,N_8173);
nor U9056 (N_9056,N_7962,N_8293);
xnor U9057 (N_9057,N_8399,N_8257);
and U9058 (N_9058,N_7545,N_7761);
nor U9059 (N_9059,N_8005,N_8861);
nand U9060 (N_9060,N_8769,N_7509);
and U9061 (N_9061,N_8037,N_8222);
and U9062 (N_9062,N_7541,N_7955);
or U9063 (N_9063,N_7824,N_8782);
nand U9064 (N_9064,N_8619,N_8758);
nor U9065 (N_9065,N_7881,N_7582);
nand U9066 (N_9066,N_7679,N_8046);
nand U9067 (N_9067,N_8159,N_7615);
and U9068 (N_9068,N_8781,N_7691);
nand U9069 (N_9069,N_8504,N_8948);
and U9070 (N_9070,N_7569,N_7747);
nand U9071 (N_9071,N_7562,N_8298);
nor U9072 (N_9072,N_8141,N_8997);
nand U9073 (N_9073,N_7603,N_8166);
and U9074 (N_9074,N_8712,N_7941);
and U9075 (N_9075,N_7806,N_8571);
or U9076 (N_9076,N_7576,N_8783);
xor U9077 (N_9077,N_8774,N_8220);
nor U9078 (N_9078,N_8474,N_8591);
xnor U9079 (N_9079,N_8886,N_7528);
and U9080 (N_9080,N_8241,N_8289);
or U9081 (N_9081,N_8610,N_8689);
or U9082 (N_9082,N_8221,N_8483);
and U9083 (N_9083,N_8801,N_8498);
xor U9084 (N_9084,N_8149,N_8217);
nor U9085 (N_9085,N_7800,N_8735);
nor U9086 (N_9086,N_7676,N_8928);
and U9087 (N_9087,N_8269,N_8442);
and U9088 (N_9088,N_8341,N_7588);
or U9089 (N_9089,N_7949,N_8891);
and U9090 (N_9090,N_7720,N_8841);
nand U9091 (N_9091,N_8092,N_8078);
xor U9092 (N_9092,N_8396,N_8660);
xnor U9093 (N_9093,N_8193,N_8875);
xnor U9094 (N_9094,N_8258,N_8249);
or U9095 (N_9095,N_7880,N_8470);
or U9096 (N_9096,N_7560,N_8291);
or U9097 (N_9097,N_8454,N_7531);
and U9098 (N_9098,N_8709,N_8937);
nand U9099 (N_9099,N_8326,N_7702);
xor U9100 (N_9100,N_8314,N_8920);
or U9101 (N_9101,N_8790,N_8379);
nand U9102 (N_9102,N_7601,N_8130);
nand U9103 (N_9103,N_8066,N_8960);
or U9104 (N_9104,N_7634,N_7748);
and U9105 (N_9105,N_8308,N_7515);
or U9106 (N_9106,N_7638,N_8635);
nor U9107 (N_9107,N_8332,N_8162);
or U9108 (N_9108,N_8287,N_8495);
and U9109 (N_9109,N_8953,N_7837);
or U9110 (N_9110,N_7697,N_7643);
xnor U9111 (N_9111,N_8980,N_8648);
and U9112 (N_9112,N_8378,N_7633);
and U9113 (N_9113,N_7721,N_7639);
and U9114 (N_9114,N_8702,N_7713);
nand U9115 (N_9115,N_8389,N_7566);
nand U9116 (N_9116,N_8867,N_7756);
nor U9117 (N_9117,N_8055,N_7820);
xor U9118 (N_9118,N_8465,N_8693);
nor U9119 (N_9119,N_8404,N_8184);
xor U9120 (N_9120,N_7695,N_8746);
or U9121 (N_9121,N_8910,N_8132);
nor U9122 (N_9122,N_8124,N_7674);
nor U9123 (N_9123,N_8323,N_8030);
xnor U9124 (N_9124,N_8219,N_8821);
or U9125 (N_9125,N_8139,N_8455);
or U9126 (N_9126,N_8760,N_8897);
or U9127 (N_9127,N_8008,N_8300);
and U9128 (N_9128,N_8866,N_7896);
and U9129 (N_9129,N_8939,N_7755);
nand U9130 (N_9130,N_8371,N_7723);
or U9131 (N_9131,N_7518,N_8788);
or U9132 (N_9132,N_8186,N_8520);
xor U9133 (N_9133,N_7868,N_7758);
xnor U9134 (N_9134,N_8240,N_8377);
or U9135 (N_9135,N_7645,N_8687);
nand U9136 (N_9136,N_8297,N_8707);
xor U9137 (N_9137,N_7696,N_8111);
and U9138 (N_9138,N_8083,N_7961);
or U9139 (N_9139,N_7670,N_7908);
and U9140 (N_9140,N_8517,N_8344);
nand U9141 (N_9141,N_8958,N_7527);
or U9142 (N_9142,N_8409,N_8535);
xor U9143 (N_9143,N_8959,N_8523);
or U9144 (N_9144,N_8573,N_8188);
xnor U9145 (N_9145,N_8178,N_8858);
nor U9146 (N_9146,N_8432,N_7530);
and U9147 (N_9147,N_8368,N_7997);
or U9148 (N_9148,N_8025,N_7623);
nand U9149 (N_9149,N_7834,N_7984);
xnor U9150 (N_9150,N_7664,N_8954);
or U9151 (N_9151,N_8271,N_8252);
xnor U9152 (N_9152,N_8775,N_7535);
nand U9153 (N_9153,N_8991,N_7829);
nand U9154 (N_9154,N_8697,N_8630);
and U9155 (N_9155,N_8677,N_8096);
or U9156 (N_9156,N_8397,N_8700);
or U9157 (N_9157,N_8235,N_8052);
xnor U9158 (N_9158,N_8737,N_7692);
nor U9159 (N_9159,N_7916,N_8988);
nand U9160 (N_9160,N_8779,N_7799);
and U9161 (N_9161,N_8104,N_8723);
nand U9162 (N_9162,N_8170,N_8246);
and U9163 (N_9163,N_7804,N_8533);
xor U9164 (N_9164,N_8012,N_8179);
and U9165 (N_9165,N_8545,N_7842);
nor U9166 (N_9166,N_8429,N_8094);
nand U9167 (N_9167,N_8759,N_8450);
nand U9168 (N_9168,N_8091,N_8811);
xnor U9169 (N_9169,N_7777,N_7845);
or U9170 (N_9170,N_8721,N_8070);
nor U9171 (N_9171,N_8730,N_7939);
xnor U9172 (N_9172,N_7621,N_7705);
and U9173 (N_9173,N_8224,N_8169);
nor U9174 (N_9174,N_8382,N_8815);
nand U9175 (N_9175,N_8419,N_7964);
and U9176 (N_9176,N_7631,N_8098);
or U9177 (N_9177,N_8418,N_8696);
nor U9178 (N_9178,N_8985,N_8206);
nand U9179 (N_9179,N_8044,N_8216);
xor U9180 (N_9180,N_8156,N_8907);
or U9181 (N_9181,N_7865,N_8107);
xor U9182 (N_9182,N_8952,N_7584);
xnor U9183 (N_9183,N_8975,N_8013);
or U9184 (N_9184,N_7520,N_8040);
and U9185 (N_9185,N_8503,N_7869);
or U9186 (N_9186,N_8965,N_8142);
or U9187 (N_9187,N_7878,N_8065);
nor U9188 (N_9188,N_8494,N_8380);
xnor U9189 (N_9189,N_7906,N_7875);
nand U9190 (N_9190,N_8238,N_7613);
or U9191 (N_9191,N_8936,N_7585);
and U9192 (N_9192,N_7924,N_8436);
nand U9193 (N_9193,N_8925,N_7813);
and U9194 (N_9194,N_8233,N_8416);
nor U9195 (N_9195,N_7625,N_8434);
nand U9196 (N_9196,N_7636,N_7708);
or U9197 (N_9197,N_8972,N_8940);
xor U9198 (N_9198,N_8295,N_8899);
nor U9199 (N_9199,N_8789,N_7701);
nor U9200 (N_9200,N_7759,N_7918);
nor U9201 (N_9201,N_8951,N_8684);
xor U9202 (N_9202,N_8294,N_8809);
nor U9203 (N_9203,N_8309,N_8989);
and U9204 (N_9204,N_7943,N_8366);
or U9205 (N_9205,N_8490,N_7938);
xnor U9206 (N_9206,N_7780,N_8706);
nand U9207 (N_9207,N_7840,N_8900);
nor U9208 (N_9208,N_8964,N_8278);
xor U9209 (N_9209,N_8019,N_7743);
nand U9210 (N_9210,N_8641,N_8225);
or U9211 (N_9211,N_7681,N_8129);
xor U9212 (N_9212,N_8829,N_8110);
nand U9213 (N_9213,N_8672,N_8489);
nor U9214 (N_9214,N_8370,N_8667);
nor U9215 (N_9215,N_7640,N_8011);
nand U9216 (N_9216,N_8830,N_8082);
and U9217 (N_9217,N_8236,N_8045);
nand U9218 (N_9218,N_7523,N_8227);
or U9219 (N_9219,N_8873,N_8812);
or U9220 (N_9220,N_8979,N_8800);
nand U9221 (N_9221,N_7719,N_7921);
or U9222 (N_9222,N_7744,N_7790);
nor U9223 (N_9223,N_7770,N_7879);
and U9224 (N_9224,N_7966,N_7682);
nand U9225 (N_9225,N_8357,N_8947);
or U9226 (N_9226,N_7774,N_8021);
nor U9227 (N_9227,N_7826,N_7792);
and U9228 (N_9228,N_7814,N_8376);
xor U9229 (N_9229,N_7712,N_8664);
nor U9230 (N_9230,N_8616,N_8460);
and U9231 (N_9231,N_8974,N_8995);
or U9232 (N_9232,N_7767,N_7765);
nand U9233 (N_9233,N_7630,N_7717);
nand U9234 (N_9234,N_8403,N_8656);
nand U9235 (N_9235,N_8254,N_8681);
or U9236 (N_9236,N_8967,N_8551);
nand U9237 (N_9237,N_8999,N_8074);
xnor U9238 (N_9238,N_7936,N_8133);
nand U9239 (N_9239,N_8405,N_8549);
nand U9240 (N_9240,N_8304,N_8844);
or U9241 (N_9241,N_8971,N_7874);
nand U9242 (N_9242,N_8556,N_8699);
or U9243 (N_9243,N_8546,N_8349);
and U9244 (N_9244,N_8905,N_7923);
nor U9245 (N_9245,N_8725,N_8365);
nand U9246 (N_9246,N_7766,N_8524);
nand U9247 (N_9247,N_8652,N_8682);
nand U9248 (N_9248,N_8207,N_8741);
or U9249 (N_9249,N_8039,N_8024);
and U9250 (N_9250,N_7822,N_8198);
nand U9251 (N_9251,N_8793,N_8753);
nor U9252 (N_9252,N_8547,N_8391);
xor U9253 (N_9253,N_8962,N_8468);
or U9254 (N_9254,N_8768,N_8077);
or U9255 (N_9255,N_8705,N_8569);
nor U9256 (N_9256,N_8525,N_8923);
nor U9257 (N_9257,N_8305,N_8736);
xor U9258 (N_9258,N_7781,N_7993);
nand U9259 (N_9259,N_8588,N_8724);
nand U9260 (N_9260,N_7660,N_7843);
xnor U9261 (N_9261,N_8580,N_8778);
or U9262 (N_9262,N_8375,N_8500);
and U9263 (N_9263,N_8451,N_7501);
or U9264 (N_9264,N_8009,N_7649);
or U9265 (N_9265,N_7779,N_8846);
xor U9266 (N_9266,N_8679,N_8154);
nand U9267 (N_9267,N_8015,N_8457);
and U9268 (N_9268,N_7534,N_8281);
or U9269 (N_9269,N_8069,N_7946);
or U9270 (N_9270,N_8329,N_8292);
nor U9271 (N_9271,N_8744,N_8134);
and U9272 (N_9272,N_8034,N_8890);
nand U9273 (N_9273,N_8876,N_8742);
nand U9274 (N_9274,N_8718,N_8464);
nor U9275 (N_9275,N_7666,N_8101);
nand U9276 (N_9276,N_8143,N_8387);
nand U9277 (N_9277,N_7740,N_8552);
xor U9278 (N_9278,N_7893,N_8417);
nand U9279 (N_9279,N_8084,N_8112);
nand U9280 (N_9280,N_8529,N_7854);
nand U9281 (N_9281,N_8734,N_8182);
xnor U9282 (N_9282,N_8051,N_8837);
nand U9283 (N_9283,N_8893,N_7716);
nor U9284 (N_9284,N_7763,N_7904);
xor U9285 (N_9285,N_8427,N_8691);
and U9286 (N_9286,N_8502,N_8898);
and U9287 (N_9287,N_8076,N_7828);
nand U9288 (N_9288,N_8270,N_7876);
xnor U9289 (N_9289,N_7972,N_7706);
xor U9290 (N_9290,N_8116,N_8311);
nand U9291 (N_9291,N_8301,N_8181);
nor U9292 (N_9292,N_8544,N_8606);
or U9293 (N_9293,N_8430,N_7995);
nor U9294 (N_9294,N_8804,N_7727);
nor U9295 (N_9295,N_7544,N_8532);
xnor U9296 (N_9296,N_8986,N_7887);
or U9297 (N_9297,N_7561,N_8582);
or U9298 (N_9298,N_7646,N_7699);
nand U9299 (N_9299,N_7506,N_8513);
or U9300 (N_9300,N_8296,N_8410);
nand U9301 (N_9301,N_8272,N_7986);
xnor U9302 (N_9302,N_8658,N_8835);
or U9303 (N_9303,N_8872,N_7787);
xnor U9304 (N_9304,N_8137,N_8594);
or U9305 (N_9305,N_8369,N_7839);
or U9306 (N_9306,N_8439,N_7605);
nand U9307 (N_9307,N_7968,N_8674);
and U9308 (N_9308,N_8497,N_8823);
or U9309 (N_9309,N_8516,N_8362);
nor U9310 (N_9310,N_8053,N_7795);
xor U9311 (N_9311,N_7500,N_8756);
nand U9312 (N_9312,N_8950,N_8888);
xor U9313 (N_9313,N_7953,N_8147);
or U9314 (N_9314,N_7899,N_8381);
nor U9315 (N_9315,N_8437,N_8374);
or U9316 (N_9316,N_8118,N_8026);
or U9317 (N_9317,N_8854,N_8845);
or U9318 (N_9318,N_8097,N_7622);
or U9319 (N_9319,N_8433,N_8102);
or U9320 (N_9320,N_8302,N_7760);
xor U9321 (N_9321,N_8061,N_7927);
or U9322 (N_9322,N_8336,N_8847);
nor U9323 (N_9323,N_8550,N_8659);
and U9324 (N_9324,N_8827,N_7565);
nand U9325 (N_9325,N_8175,N_7957);
xnor U9326 (N_9326,N_8728,N_8010);
nor U9327 (N_9327,N_8536,N_7819);
xnor U9328 (N_9328,N_8617,N_7581);
xnor U9329 (N_9329,N_7898,N_8319);
xor U9330 (N_9330,N_8507,N_7726);
nand U9331 (N_9331,N_8957,N_8956);
and U9332 (N_9332,N_7857,N_8796);
and U9333 (N_9333,N_8386,N_7889);
nand U9334 (N_9334,N_7967,N_8242);
nand U9335 (N_9335,N_8711,N_8438);
xor U9336 (N_9336,N_8828,N_8559);
xor U9337 (N_9337,N_7508,N_8354);
and U9338 (N_9338,N_8627,N_8968);
xnor U9339 (N_9339,N_8683,N_7546);
nor U9340 (N_9340,N_8817,N_8036);
or U9341 (N_9341,N_8637,N_8935);
nand U9342 (N_9342,N_8738,N_8231);
or U9343 (N_9343,N_8632,N_7920);
and U9344 (N_9344,N_7662,N_8339);
xnor U9345 (N_9345,N_8745,N_7606);
xor U9346 (N_9346,N_8719,N_8239);
and U9347 (N_9347,N_7933,N_8245);
nand U9348 (N_9348,N_8187,N_7832);
or U9349 (N_9349,N_8398,N_8895);
or U9350 (N_9350,N_8848,N_8856);
nand U9351 (N_9351,N_8813,N_8592);
or U9352 (N_9352,N_7882,N_7772);
nand U9353 (N_9353,N_8315,N_7988);
xor U9354 (N_9354,N_8058,N_8018);
nand U9355 (N_9355,N_8933,N_8415);
or U9356 (N_9356,N_7659,N_7808);
xor U9357 (N_9357,N_7590,N_8190);
or U9358 (N_9358,N_7607,N_8978);
or U9359 (N_9359,N_8447,N_7729);
xor U9360 (N_9360,N_8140,N_8203);
xor U9361 (N_9361,N_8818,N_8992);
and U9362 (N_9362,N_7652,N_8824);
nor U9363 (N_9363,N_7771,N_8108);
and U9364 (N_9364,N_8963,N_7746);
and U9365 (N_9365,N_7852,N_8138);
and U9366 (N_9366,N_8668,N_8717);
xor U9367 (N_9367,N_7786,N_8943);
nor U9368 (N_9368,N_8911,N_8176);
xnor U9369 (N_9369,N_7870,N_8966);
nor U9370 (N_9370,N_7610,N_8148);
xnor U9371 (N_9371,N_8625,N_7977);
xor U9372 (N_9372,N_7710,N_7574);
nor U9373 (N_9373,N_8327,N_8444);
or U9374 (N_9374,N_8612,N_7563);
and U9375 (N_9375,N_8448,N_8064);
and U9376 (N_9376,N_7959,N_7841);
or U9377 (N_9377,N_7930,N_8251);
xor U9378 (N_9378,N_8476,N_8320);
and U9379 (N_9379,N_7970,N_8440);
nand U9380 (N_9380,N_7653,N_7846);
nand U9381 (N_9381,N_8539,N_8004);
xnor U9382 (N_9382,N_8808,N_7592);
nand U9383 (N_9383,N_8067,N_7626);
or U9384 (N_9384,N_7942,N_7703);
nand U9385 (N_9385,N_7764,N_7807);
and U9386 (N_9386,N_8420,N_8931);
xnor U9387 (N_9387,N_8563,N_7883);
xor U9388 (N_9388,N_7715,N_8060);
xor U9389 (N_9389,N_8915,N_8708);
xnor U9390 (N_9390,N_8127,N_8456);
nand U9391 (N_9391,N_8250,N_8079);
and U9392 (N_9392,N_8215,N_7902);
xor U9393 (N_9393,N_8445,N_8859);
and U9394 (N_9394,N_7954,N_7752);
nor U9395 (N_9395,N_8145,N_8321);
nor U9396 (N_9396,N_8347,N_7655);
xnor U9397 (N_9397,N_8653,N_8651);
xor U9398 (N_9398,N_8570,N_7594);
nor U9399 (N_9399,N_8209,N_8784);
and U9400 (N_9400,N_8715,N_8038);
nor U9401 (N_9401,N_8600,N_7671);
or U9402 (N_9402,N_8863,N_8831);
xor U9403 (N_9403,N_7917,N_8896);
nand U9404 (N_9404,N_8361,N_8628);
xor U9405 (N_9405,N_7980,N_7648);
nand U9406 (N_9406,N_8643,N_8740);
nor U9407 (N_9407,N_8312,N_8528);
nand U9408 (N_9408,N_8214,N_8969);
nor U9409 (N_9409,N_8595,N_7644);
nand U9410 (N_9410,N_7973,N_8572);
or U9411 (N_9411,N_7886,N_7794);
or U9412 (N_9412,N_8299,N_8767);
or U9413 (N_9413,N_7549,N_8688);
xnor U9414 (N_9414,N_8634,N_8355);
nor U9415 (N_9415,N_8698,N_8534);
and U9416 (N_9416,N_7778,N_8695);
nand U9417 (N_9417,N_8623,N_7619);
nor U9418 (N_9418,N_8493,N_8340);
nand U9419 (N_9419,N_8820,N_8977);
and U9420 (N_9420,N_8482,N_7536);
or U9421 (N_9421,N_8904,N_8566);
xor U9422 (N_9422,N_8560,N_8877);
nand U9423 (N_9423,N_8189,N_8099);
xnor U9424 (N_9424,N_8716,N_7782);
or U9425 (N_9425,N_8324,N_8491);
xor U9426 (N_9426,N_7816,N_8605);
nor U9427 (N_9427,N_7683,N_7791);
and U9428 (N_9428,N_8666,N_8373);
or U9429 (N_9429,N_8194,N_8212);
xnor U9430 (N_9430,N_8351,N_8285);
and U9431 (N_9431,N_7969,N_8113);
nor U9432 (N_9432,N_8115,N_8307);
nand U9433 (N_9433,N_8185,N_8624);
xor U9434 (N_9434,N_7564,N_7618);
or U9435 (N_9435,N_7912,N_8622);
nor U9436 (N_9436,N_8732,N_8575);
nand U9437 (N_9437,N_8508,N_8201);
xnor U9438 (N_9438,N_8917,N_8047);
or U9439 (N_9439,N_7913,N_8511);
nor U9440 (N_9440,N_8929,N_8348);
nor U9441 (N_9441,N_8274,N_8343);
or U9442 (N_9442,N_8144,N_7556);
or U9443 (N_9443,N_8938,N_8392);
nor U9444 (N_9444,N_8894,N_8710);
or U9445 (N_9445,N_8049,N_8123);
and U9446 (N_9446,N_7950,N_7735);
nor U9447 (N_9447,N_8467,N_8325);
and U9448 (N_9448,N_8395,N_8776);
or U9449 (N_9449,N_8629,N_8244);
or U9450 (N_9450,N_8086,N_8168);
nand U9451 (N_9451,N_8983,N_7810);
nor U9452 (N_9452,N_8155,N_8955);
nand U9453 (N_9453,N_7543,N_8871);
nor U9454 (N_9454,N_7925,N_8330);
or U9455 (N_9455,N_8264,N_8880);
or U9456 (N_9456,N_8128,N_7855);
or U9457 (N_9457,N_8317,N_8263);
nand U9458 (N_9458,N_8136,N_8574);
xnor U9459 (N_9459,N_8267,N_7749);
xnor U9460 (N_9460,N_8506,N_7629);
xnor U9461 (N_9461,N_7504,N_8633);
nand U9462 (N_9462,N_7524,N_7687);
nand U9463 (N_9463,N_8346,N_7597);
nor U9464 (N_9464,N_7669,N_7700);
xor U9465 (N_9465,N_8833,N_8469);
and U9466 (N_9466,N_7709,N_7751);
or U9467 (N_9467,N_7718,N_8869);
nand U9468 (N_9468,N_8849,N_8860);
and U9469 (N_9469,N_8865,N_7690);
nor U9470 (N_9470,N_8825,N_8874);
and U9471 (N_9471,N_7572,N_8638);
xor U9472 (N_9472,N_8541,N_7647);
and U9473 (N_9473,N_8177,N_8596);
nor U9474 (N_9474,N_8996,N_8080);
nor U9475 (N_9475,N_8657,N_7975);
nor U9476 (N_9476,N_8577,N_8879);
and U9477 (N_9477,N_8771,N_8288);
or U9478 (N_9478,N_8165,N_8713);
or U9479 (N_9479,N_7981,N_8807);
xnor U9480 (N_9480,N_8268,N_7821);
nand U9481 (N_9481,N_7624,N_8538);
nand U9482 (N_9482,N_8926,N_8063);
or U9483 (N_9483,N_7910,N_8739);
and U9484 (N_9484,N_8477,N_8488);
xor U9485 (N_9485,N_8255,N_8558);
nor U9486 (N_9486,N_7673,N_7935);
nand U9487 (N_9487,N_8645,N_8350);
or U9488 (N_9488,N_7940,N_7632);
nor U9489 (N_9489,N_8729,N_7741);
xor U9490 (N_9490,N_8601,N_8003);
xor U9491 (N_9491,N_8527,N_7548);
nor U9492 (N_9492,N_8990,N_8543);
nand U9493 (N_9493,N_8090,N_8542);
and U9494 (N_9494,N_8665,N_7952);
or U9495 (N_9495,N_8088,N_7991);
or U9496 (N_9496,N_8704,N_8836);
or U9497 (N_9497,N_7937,N_8001);
or U9498 (N_9498,N_7551,N_7686);
nor U9499 (N_9499,N_7785,N_8889);
and U9500 (N_9500,N_8318,N_7725);
nand U9501 (N_9501,N_8806,N_8908);
nor U9502 (N_9502,N_8671,N_7586);
and U9503 (N_9503,N_8919,N_8383);
or U9504 (N_9504,N_8647,N_7689);
xnor U9505 (N_9505,N_7704,N_8649);
and U9506 (N_9506,N_7510,N_7784);
nand U9507 (N_9507,N_8982,N_8353);
xnor U9508 (N_9508,N_8810,N_7979);
xnor U9509 (N_9509,N_8218,N_7602);
xor U9510 (N_9510,N_8870,N_8797);
nand U9511 (N_9511,N_8480,N_7578);
or U9512 (N_9512,N_7836,N_8411);
nand U9513 (N_9513,N_7730,N_8703);
and U9514 (N_9514,N_7895,N_7680);
and U9515 (N_9515,N_8531,N_7919);
nor U9516 (N_9516,N_7722,N_8050);
nor U9517 (N_9517,N_8388,N_8458);
nand U9518 (N_9518,N_8661,N_7511);
nand U9519 (N_9519,N_8423,N_8984);
and U9520 (N_9520,N_7947,N_8196);
or U9521 (N_9521,N_8822,N_8994);
nor U9522 (N_9522,N_8016,N_7905);
nand U9523 (N_9523,N_8290,N_7614);
nor U9524 (N_9524,N_8020,N_8478);
and U9525 (N_9525,N_8342,N_8075);
and U9526 (N_9526,N_8443,N_8043);
xor U9527 (N_9527,N_8152,N_8213);
and U9528 (N_9528,N_8690,N_8505);
xnor U9529 (N_9529,N_8461,N_8930);
and U9530 (N_9530,N_7976,N_8199);
nor U9531 (N_9531,N_8441,N_8914);
and U9532 (N_9532,N_8568,N_8526);
xnor U9533 (N_9533,N_8777,N_7863);
xnor U9534 (N_9534,N_7555,N_7591);
nand U9535 (N_9535,N_7512,N_7573);
xor U9536 (N_9536,N_8655,N_8587);
nor U9537 (N_9537,N_8204,N_7522);
nand U9538 (N_9538,N_8260,N_7525);
nand U9539 (N_9539,N_7550,N_8662);
or U9540 (N_9540,N_7609,N_8028);
and U9541 (N_9541,N_7797,N_8059);
xnor U9542 (N_9542,N_8484,N_8322);
nor U9543 (N_9543,N_8243,N_8604);
and U9544 (N_9544,N_8426,N_8639);
or U9545 (N_9545,N_7616,N_7866);
or U9546 (N_9546,N_8642,N_7915);
nand U9547 (N_9547,N_8007,N_7803);
xor U9548 (N_9548,N_8275,N_8581);
nand U9549 (N_9549,N_7812,N_8934);
nand U9550 (N_9550,N_8200,N_7985);
nand U9551 (N_9551,N_7796,N_7934);
nand U9552 (N_9552,N_8473,N_8564);
nand U9553 (N_9553,N_7732,N_8903);
and U9554 (N_9554,N_8692,N_8614);
and U9555 (N_9555,N_8453,N_7983);
or U9556 (N_9556,N_8256,N_7678);
and U9557 (N_9557,N_7529,N_8412);
nand U9558 (N_9558,N_7989,N_8266);
xor U9559 (N_9559,N_7533,N_8770);
nand U9560 (N_9560,N_8431,N_7775);
nor U9561 (N_9561,N_7635,N_8843);
nand U9562 (N_9562,N_8901,N_7773);
nand U9563 (N_9563,N_8731,N_7974);
and U9564 (N_9564,N_8210,N_8613);
xor U9565 (N_9565,N_8576,N_8422);
or U9566 (N_9566,N_8819,N_7892);
nor U9567 (N_9567,N_8727,N_7818);
nor U9568 (N_9568,N_8095,N_8654);
nand U9569 (N_9569,N_7769,N_8921);
and U9570 (N_9570,N_8229,N_8615);
nor U9571 (N_9571,N_8916,N_8424);
nand U9572 (N_9572,N_8557,N_7517);
and U9573 (N_9573,N_8862,N_8125);
xor U9574 (N_9574,N_8747,N_8180);
or U9575 (N_9575,N_7587,N_7599);
and U9576 (N_9576,N_8071,N_7542);
nand U9577 (N_9577,N_8117,N_7877);
and U9578 (N_9578,N_8384,N_7608);
and U9579 (N_9579,N_7503,N_8763);
or U9580 (N_9580,N_8022,N_8912);
or U9581 (N_9581,N_8882,N_8232);
and U9582 (N_9582,N_7731,N_8226);
nor U9583 (N_9583,N_7844,N_8390);
nand U9584 (N_9584,N_8805,N_7568);
or U9585 (N_9585,N_7872,N_7583);
xnor U9586 (N_9586,N_7817,N_8585);
nor U9587 (N_9587,N_8496,N_8492);
xnor U9588 (N_9588,N_8487,N_8726);
xor U9589 (N_9589,N_8761,N_8103);
or U9590 (N_9590,N_7728,N_8584);
and U9591 (N_9591,N_7693,N_8230);
nor U9592 (N_9592,N_8987,N_8764);
or U9593 (N_9593,N_8565,N_8081);
nor U9594 (N_9594,N_8814,N_8032);
or U9595 (N_9595,N_8754,N_7783);
nor U9596 (N_9596,N_8393,N_8485);
nor U9597 (N_9597,N_8402,N_7929);
nand U9598 (N_9598,N_8262,N_7944);
nand U9599 (N_9599,N_8119,N_8428);
nand U9600 (N_9600,N_7554,N_8620);
nand U9601 (N_9601,N_8481,N_8135);
or U9602 (N_9602,N_8519,N_8832);
nor U9603 (N_9603,N_8799,N_7514);
nand U9604 (N_9604,N_8131,N_7971);
nor U9605 (N_9605,N_7823,N_8787);
or U9606 (N_9606,N_8085,N_8406);
or U9607 (N_9607,N_8105,N_7733);
or U9608 (N_9608,N_8772,N_8593);
nand U9609 (N_9609,N_8548,N_8282);
and U9610 (N_9610,N_7833,N_8073);
and U9611 (N_9611,N_7830,N_8106);
nor U9612 (N_9612,N_7711,N_8646);
xnor U9613 (N_9613,N_8868,N_8006);
and U9614 (N_9614,N_8253,N_8033);
and U9615 (N_9615,N_8163,N_7580);
xor U9616 (N_9616,N_8553,N_8607);
xor U9617 (N_9617,N_7798,N_7805);
nor U9618 (N_9618,N_7768,N_8598);
nor U9619 (N_9619,N_8466,N_7932);
nor U9620 (N_9620,N_7596,N_7888);
or U9621 (N_9621,N_8247,N_7856);
nor U9622 (N_9622,N_7505,N_8945);
nor U9623 (N_9623,N_8273,N_8195);
or U9624 (N_9624,N_8680,N_8167);
nand U9625 (N_9625,N_8228,N_8237);
or U9626 (N_9626,N_7724,N_8372);
xnor U9627 (N_9627,N_8803,N_8678);
nor U9628 (N_9628,N_8636,N_8883);
xor U9629 (N_9629,N_7847,N_7825);
or U9630 (N_9630,N_8486,N_8414);
nor U9631 (N_9631,N_7739,N_8676);
nand U9632 (N_9632,N_8352,N_8521);
nor U9633 (N_9633,N_7945,N_8234);
nand U9634 (N_9634,N_7651,N_8191);
or U9635 (N_9635,N_8949,N_8918);
or U9636 (N_9636,N_7922,N_7827);
xnor U9637 (N_9637,N_8062,N_7931);
and U9638 (N_9638,N_7848,N_7579);
nor U9639 (N_9639,N_7885,N_8276);
or U9640 (N_9640,N_8892,N_7907);
and U9641 (N_9641,N_8385,N_8590);
and U9642 (N_9642,N_8407,N_7502);
nand U9643 (N_9643,N_8618,N_8650);
nor U9644 (N_9644,N_7862,N_8686);
nor U9645 (N_9645,N_8452,N_8878);
xnor U9646 (N_9646,N_8068,N_8851);
or U9647 (N_9647,N_7567,N_8345);
xnor U9648 (N_9648,N_8023,N_8792);
nor U9649 (N_9649,N_7811,N_8408);
nand U9650 (N_9650,N_7871,N_8183);
or U9651 (N_9651,N_8766,N_8002);
or U9652 (N_9652,N_8816,N_8884);
nor U9653 (N_9653,N_8621,N_8902);
xnor U9654 (N_9654,N_8158,N_8359);
or U9655 (N_9655,N_7575,N_7552);
nor U9656 (N_9656,N_8640,N_7658);
or U9657 (N_9657,N_7571,N_7507);
xnor U9658 (N_9658,N_8981,N_8946);
and U9659 (N_9659,N_7698,N_8161);
xor U9660 (N_9660,N_7864,N_8367);
nand U9661 (N_9661,N_7815,N_8122);
and U9662 (N_9662,N_8993,N_8512);
or U9663 (N_9663,N_8280,N_8554);
nand U9664 (N_9664,N_8171,N_8714);
nor U9665 (N_9665,N_8589,N_7958);
and U9666 (N_9666,N_8017,N_8701);
nor U9667 (N_9667,N_8425,N_7558);
and U9668 (N_9668,N_8780,N_7802);
nor U9669 (N_9669,N_7672,N_7894);
or U9670 (N_9670,N_8014,N_7617);
nand U9671 (N_9671,N_8608,N_8157);
or U9672 (N_9672,N_7707,N_7835);
nand U9673 (N_9673,N_8755,N_8749);
xor U9674 (N_9674,N_8853,N_7637);
nand U9675 (N_9675,N_8510,N_7867);
and U9676 (N_9676,N_7789,N_7685);
and U9677 (N_9677,N_7628,N_8611);
or U9678 (N_9678,N_7996,N_8316);
nand U9679 (N_9679,N_8750,N_7901);
or U9680 (N_9680,N_8864,N_7521);
xnor U9681 (N_9681,N_7519,N_8121);
or U9682 (N_9682,N_8670,N_7793);
and U9683 (N_9683,N_8785,N_8499);
nand U9684 (N_9684,N_7745,N_8333);
xnor U9685 (N_9685,N_8924,N_8100);
nor U9686 (N_9686,N_8463,N_8941);
or U9687 (N_9687,N_8694,N_7620);
and U9688 (N_9688,N_7914,N_7537);
xnor U9689 (N_9689,N_7570,N_7757);
xor U9690 (N_9690,N_7801,N_7762);
xnor U9691 (N_9691,N_7611,N_8151);
xor U9692 (N_9692,N_7650,N_7897);
nand U9693 (N_9693,N_8356,N_8720);
xnor U9694 (N_9694,N_7928,N_8976);
xor U9695 (N_9695,N_8583,N_8631);
nand U9696 (N_9696,N_8970,N_8306);
nand U9697 (N_9697,N_8413,N_7951);
and U9698 (N_9698,N_8826,N_8146);
and U9699 (N_9699,N_8335,N_8515);
nand U9700 (N_9700,N_7694,N_8475);
and U9701 (N_9701,N_8150,N_7851);
and U9702 (N_9702,N_7593,N_7654);
nand U9703 (N_9703,N_8358,N_7994);
xnor U9704 (N_9704,N_8093,N_8743);
nand U9705 (N_9705,N_8567,N_7948);
nand U9706 (N_9706,N_8839,N_8109);
and U9707 (N_9707,N_8599,N_7675);
xor U9708 (N_9708,N_7850,N_8913);
xnor U9709 (N_9709,N_7960,N_7657);
nor U9710 (N_9710,N_8850,N_8609);
xor U9711 (N_9711,N_8459,N_7750);
nor U9712 (N_9712,N_8857,N_8751);
and U9713 (N_9713,N_7516,N_7553);
or U9714 (N_9714,N_8530,N_8279);
xnor U9715 (N_9715,N_8998,N_7900);
and U9716 (N_9716,N_8773,N_7665);
nor U9717 (N_9717,N_8663,N_8334);
nand U9718 (N_9718,N_8757,N_8602);
or U9719 (N_9719,N_7982,N_8603);
or U9720 (N_9720,N_7513,N_7641);
nor U9721 (N_9721,N_8842,N_7809);
nor U9722 (N_9722,N_8310,N_7890);
xor U9723 (N_9723,N_8927,N_8197);
and U9724 (N_9724,N_7831,N_8363);
and U9725 (N_9725,N_8284,N_8265);
nor U9726 (N_9726,N_7859,N_8261);
and U9727 (N_9727,N_8906,N_8364);
or U9728 (N_9728,N_7595,N_7559);
nand U9729 (N_9729,N_8579,N_8401);
nor U9730 (N_9730,N_7688,N_7677);
or U9731 (N_9731,N_8160,N_7849);
or U9732 (N_9732,N_8909,N_7540);
nand U9733 (N_9733,N_8944,N_7539);
xor U9734 (N_9734,N_8041,N_7776);
or U9735 (N_9735,N_7538,N_7911);
and U9736 (N_9736,N_8360,N_8922);
or U9737 (N_9737,N_7642,N_8072);
xnor U9738 (N_9738,N_7965,N_7736);
xnor U9739 (N_9739,N_8446,N_7663);
or U9740 (N_9740,N_8802,N_8027);
nand U9741 (N_9741,N_7612,N_8669);
xor U9742 (N_9742,N_7738,N_8120);
nand U9743 (N_9743,N_7598,N_7667);
and U9744 (N_9744,N_8518,N_8887);
nand U9745 (N_9745,N_7909,N_8597);
or U9746 (N_9746,N_8722,N_8421);
nor U9747 (N_9747,N_8586,N_8283);
nand U9748 (N_9748,N_8855,N_8514);
nor U9749 (N_9749,N_8795,N_8338);
or U9750 (N_9750,N_7867,N_8697);
nor U9751 (N_9751,N_8741,N_7744);
nor U9752 (N_9752,N_8840,N_8367);
nor U9753 (N_9753,N_8877,N_7722);
or U9754 (N_9754,N_8604,N_8099);
or U9755 (N_9755,N_7636,N_7686);
xnor U9756 (N_9756,N_7503,N_8839);
nand U9757 (N_9757,N_7771,N_8419);
xnor U9758 (N_9758,N_7699,N_8957);
xnor U9759 (N_9759,N_7790,N_8172);
and U9760 (N_9760,N_7790,N_7539);
nor U9761 (N_9761,N_8248,N_7691);
and U9762 (N_9762,N_7628,N_7714);
nand U9763 (N_9763,N_8026,N_8311);
nand U9764 (N_9764,N_8758,N_8963);
nor U9765 (N_9765,N_8684,N_8916);
nand U9766 (N_9766,N_7615,N_8494);
xnor U9767 (N_9767,N_8115,N_8084);
nand U9768 (N_9768,N_8262,N_7938);
xor U9769 (N_9769,N_8994,N_7579);
nand U9770 (N_9770,N_8982,N_8284);
or U9771 (N_9771,N_8484,N_7543);
nor U9772 (N_9772,N_7742,N_7571);
xor U9773 (N_9773,N_8365,N_7531);
or U9774 (N_9774,N_8245,N_7898);
nor U9775 (N_9775,N_7934,N_8074);
or U9776 (N_9776,N_7726,N_7869);
xnor U9777 (N_9777,N_8840,N_8736);
nor U9778 (N_9778,N_8841,N_7564);
xnor U9779 (N_9779,N_8000,N_8611);
nand U9780 (N_9780,N_8052,N_8453);
and U9781 (N_9781,N_8733,N_7961);
nand U9782 (N_9782,N_8089,N_7767);
nand U9783 (N_9783,N_8197,N_8886);
xor U9784 (N_9784,N_8420,N_8232);
xnor U9785 (N_9785,N_7883,N_8417);
xnor U9786 (N_9786,N_7775,N_8568);
nand U9787 (N_9787,N_7699,N_7703);
or U9788 (N_9788,N_8898,N_8617);
xnor U9789 (N_9789,N_8642,N_8570);
xnor U9790 (N_9790,N_7740,N_7941);
nor U9791 (N_9791,N_7914,N_7660);
nor U9792 (N_9792,N_8095,N_8870);
nor U9793 (N_9793,N_8755,N_8532);
nor U9794 (N_9794,N_8121,N_7897);
nand U9795 (N_9795,N_7654,N_8173);
xnor U9796 (N_9796,N_7905,N_7652);
and U9797 (N_9797,N_7736,N_8232);
nand U9798 (N_9798,N_7771,N_7576);
nand U9799 (N_9799,N_8031,N_7863);
and U9800 (N_9800,N_8533,N_7973);
and U9801 (N_9801,N_8550,N_8951);
or U9802 (N_9802,N_7810,N_8610);
xor U9803 (N_9803,N_7936,N_8279);
nand U9804 (N_9804,N_8791,N_7876);
xnor U9805 (N_9805,N_8757,N_7879);
xor U9806 (N_9806,N_8808,N_7584);
nand U9807 (N_9807,N_7525,N_8321);
or U9808 (N_9808,N_8874,N_7563);
nor U9809 (N_9809,N_8579,N_8181);
and U9810 (N_9810,N_8981,N_7634);
and U9811 (N_9811,N_8444,N_7670);
and U9812 (N_9812,N_7580,N_7545);
xnor U9813 (N_9813,N_8832,N_7878);
nand U9814 (N_9814,N_8849,N_8754);
nand U9815 (N_9815,N_7583,N_8908);
and U9816 (N_9816,N_8894,N_8242);
and U9817 (N_9817,N_8230,N_8784);
and U9818 (N_9818,N_8915,N_7712);
or U9819 (N_9819,N_7587,N_8528);
or U9820 (N_9820,N_8818,N_8186);
or U9821 (N_9821,N_8610,N_8087);
xor U9822 (N_9822,N_8399,N_8402);
xnor U9823 (N_9823,N_8264,N_8798);
xor U9824 (N_9824,N_7795,N_8510);
nor U9825 (N_9825,N_7692,N_8655);
xor U9826 (N_9826,N_7831,N_8761);
and U9827 (N_9827,N_8198,N_8970);
and U9828 (N_9828,N_8877,N_8974);
or U9829 (N_9829,N_8176,N_8196);
nor U9830 (N_9830,N_7581,N_8115);
nand U9831 (N_9831,N_7980,N_7921);
xor U9832 (N_9832,N_8287,N_8860);
and U9833 (N_9833,N_8119,N_8863);
or U9834 (N_9834,N_8846,N_7531);
nor U9835 (N_9835,N_8218,N_8801);
or U9836 (N_9836,N_8749,N_8255);
xor U9837 (N_9837,N_7968,N_8893);
and U9838 (N_9838,N_7702,N_8379);
xor U9839 (N_9839,N_8563,N_8132);
or U9840 (N_9840,N_8769,N_8572);
nand U9841 (N_9841,N_7812,N_8563);
nor U9842 (N_9842,N_7553,N_8328);
and U9843 (N_9843,N_8249,N_8064);
nand U9844 (N_9844,N_8738,N_7562);
and U9845 (N_9845,N_8826,N_8176);
xor U9846 (N_9846,N_8777,N_8518);
nand U9847 (N_9847,N_8005,N_8415);
nand U9848 (N_9848,N_8734,N_8886);
and U9849 (N_9849,N_8075,N_7778);
or U9850 (N_9850,N_8351,N_8768);
xnor U9851 (N_9851,N_8067,N_8779);
or U9852 (N_9852,N_7623,N_7895);
and U9853 (N_9853,N_8294,N_8125);
nand U9854 (N_9854,N_8997,N_8955);
nand U9855 (N_9855,N_7551,N_8700);
nand U9856 (N_9856,N_8226,N_8348);
and U9857 (N_9857,N_8434,N_8576);
or U9858 (N_9858,N_7791,N_8654);
or U9859 (N_9859,N_8363,N_8959);
nor U9860 (N_9860,N_8839,N_8779);
xnor U9861 (N_9861,N_8231,N_8421);
nand U9862 (N_9862,N_8603,N_8907);
and U9863 (N_9863,N_7985,N_7652);
nand U9864 (N_9864,N_8563,N_7958);
xor U9865 (N_9865,N_8885,N_8733);
xnor U9866 (N_9866,N_8044,N_7559);
nand U9867 (N_9867,N_8663,N_8216);
or U9868 (N_9868,N_8510,N_7593);
and U9869 (N_9869,N_7575,N_8449);
xor U9870 (N_9870,N_8275,N_8372);
xnor U9871 (N_9871,N_8454,N_8384);
xor U9872 (N_9872,N_8841,N_8689);
and U9873 (N_9873,N_8818,N_8822);
xor U9874 (N_9874,N_8464,N_7932);
xor U9875 (N_9875,N_8026,N_7800);
or U9876 (N_9876,N_8143,N_7811);
or U9877 (N_9877,N_7908,N_8518);
and U9878 (N_9878,N_8264,N_7985);
or U9879 (N_9879,N_8304,N_8213);
and U9880 (N_9880,N_8520,N_8740);
or U9881 (N_9881,N_7926,N_7698);
and U9882 (N_9882,N_7683,N_8144);
nor U9883 (N_9883,N_8940,N_8537);
xnor U9884 (N_9884,N_8823,N_8072);
or U9885 (N_9885,N_8475,N_8530);
xnor U9886 (N_9886,N_8233,N_8102);
and U9887 (N_9887,N_8936,N_8531);
or U9888 (N_9888,N_8214,N_8544);
or U9889 (N_9889,N_8068,N_8478);
xor U9890 (N_9890,N_7611,N_8680);
xor U9891 (N_9891,N_8684,N_8918);
nand U9892 (N_9892,N_7959,N_8512);
and U9893 (N_9893,N_8848,N_8701);
xnor U9894 (N_9894,N_8876,N_8048);
and U9895 (N_9895,N_7583,N_8320);
nor U9896 (N_9896,N_8257,N_8006);
or U9897 (N_9897,N_8907,N_8380);
nor U9898 (N_9898,N_8826,N_7512);
xor U9899 (N_9899,N_7664,N_8892);
xnor U9900 (N_9900,N_7898,N_8867);
xnor U9901 (N_9901,N_8740,N_8105);
xor U9902 (N_9902,N_8891,N_8421);
xnor U9903 (N_9903,N_8721,N_8502);
nor U9904 (N_9904,N_8345,N_7665);
xnor U9905 (N_9905,N_7567,N_8229);
nor U9906 (N_9906,N_8382,N_8330);
xnor U9907 (N_9907,N_7864,N_7675);
xnor U9908 (N_9908,N_7542,N_7980);
nor U9909 (N_9909,N_8597,N_8159);
and U9910 (N_9910,N_8722,N_8512);
nor U9911 (N_9911,N_7606,N_7551);
and U9912 (N_9912,N_8227,N_7689);
or U9913 (N_9913,N_8084,N_8620);
nand U9914 (N_9914,N_8378,N_7816);
xnor U9915 (N_9915,N_8855,N_8427);
xnor U9916 (N_9916,N_8657,N_7666);
nor U9917 (N_9917,N_8490,N_8030);
nand U9918 (N_9918,N_8016,N_7641);
and U9919 (N_9919,N_7636,N_8168);
or U9920 (N_9920,N_8116,N_7984);
nand U9921 (N_9921,N_7675,N_7577);
and U9922 (N_9922,N_8457,N_8296);
xnor U9923 (N_9923,N_7953,N_8361);
xnor U9924 (N_9924,N_8699,N_8946);
nor U9925 (N_9925,N_7774,N_8091);
or U9926 (N_9926,N_8759,N_7620);
and U9927 (N_9927,N_8459,N_7636);
nor U9928 (N_9928,N_8057,N_8451);
or U9929 (N_9929,N_7856,N_7613);
nand U9930 (N_9930,N_8471,N_8936);
nand U9931 (N_9931,N_7826,N_8497);
and U9932 (N_9932,N_8172,N_8727);
xnor U9933 (N_9933,N_8237,N_8832);
or U9934 (N_9934,N_8855,N_8363);
and U9935 (N_9935,N_7970,N_8863);
xor U9936 (N_9936,N_8095,N_7543);
nand U9937 (N_9937,N_7675,N_7986);
nor U9938 (N_9938,N_8410,N_8281);
nor U9939 (N_9939,N_7793,N_8075);
xor U9940 (N_9940,N_7798,N_7741);
and U9941 (N_9941,N_8977,N_8178);
or U9942 (N_9942,N_8868,N_7663);
or U9943 (N_9943,N_8525,N_7757);
nand U9944 (N_9944,N_8152,N_7790);
nand U9945 (N_9945,N_8563,N_8779);
xnor U9946 (N_9946,N_8035,N_8373);
or U9947 (N_9947,N_7928,N_8736);
xnor U9948 (N_9948,N_8905,N_7686);
nand U9949 (N_9949,N_8774,N_8746);
nor U9950 (N_9950,N_8115,N_8077);
and U9951 (N_9951,N_7686,N_8782);
nand U9952 (N_9952,N_8629,N_8610);
and U9953 (N_9953,N_7633,N_8486);
nor U9954 (N_9954,N_7812,N_7712);
nor U9955 (N_9955,N_7789,N_8798);
and U9956 (N_9956,N_7595,N_8402);
nand U9957 (N_9957,N_8658,N_7759);
and U9958 (N_9958,N_8925,N_8807);
and U9959 (N_9959,N_7980,N_8854);
and U9960 (N_9960,N_8076,N_7968);
nor U9961 (N_9961,N_7832,N_8311);
nor U9962 (N_9962,N_8500,N_8776);
xnor U9963 (N_9963,N_8255,N_8058);
nor U9964 (N_9964,N_7910,N_8213);
and U9965 (N_9965,N_7935,N_7800);
nand U9966 (N_9966,N_7732,N_8526);
or U9967 (N_9967,N_8790,N_8564);
nor U9968 (N_9968,N_8191,N_8536);
nor U9969 (N_9969,N_8915,N_8525);
or U9970 (N_9970,N_7664,N_7747);
or U9971 (N_9971,N_7727,N_8307);
or U9972 (N_9972,N_7817,N_7687);
nor U9973 (N_9973,N_8066,N_8668);
nor U9974 (N_9974,N_8933,N_7598);
nor U9975 (N_9975,N_8696,N_7671);
or U9976 (N_9976,N_8826,N_8668);
or U9977 (N_9977,N_7758,N_7958);
nand U9978 (N_9978,N_8527,N_8984);
nor U9979 (N_9979,N_8601,N_7894);
and U9980 (N_9980,N_8573,N_8396);
nand U9981 (N_9981,N_8280,N_7982);
nor U9982 (N_9982,N_7811,N_7783);
nand U9983 (N_9983,N_8139,N_8021);
nor U9984 (N_9984,N_8100,N_8527);
and U9985 (N_9985,N_8797,N_7967);
xnor U9986 (N_9986,N_8081,N_7744);
xor U9987 (N_9987,N_8082,N_8237);
xnor U9988 (N_9988,N_7779,N_8013);
xor U9989 (N_9989,N_8762,N_7567);
nor U9990 (N_9990,N_8896,N_8635);
nor U9991 (N_9991,N_8966,N_7512);
and U9992 (N_9992,N_8987,N_8113);
nand U9993 (N_9993,N_8682,N_8909);
nand U9994 (N_9994,N_8703,N_8353);
and U9995 (N_9995,N_7738,N_8333);
nor U9996 (N_9996,N_7651,N_7807);
and U9997 (N_9997,N_7671,N_8212);
nor U9998 (N_9998,N_7669,N_8871);
xor U9999 (N_9999,N_8799,N_8890);
nand U10000 (N_10000,N_8460,N_8252);
xnor U10001 (N_10001,N_8627,N_7946);
nor U10002 (N_10002,N_8972,N_8983);
xnor U10003 (N_10003,N_8401,N_7818);
and U10004 (N_10004,N_8233,N_8685);
or U10005 (N_10005,N_8613,N_7854);
nand U10006 (N_10006,N_7970,N_8772);
or U10007 (N_10007,N_8135,N_8058);
nand U10008 (N_10008,N_8149,N_7990);
and U10009 (N_10009,N_8017,N_7929);
nor U10010 (N_10010,N_7529,N_7570);
and U10011 (N_10011,N_8015,N_8111);
nor U10012 (N_10012,N_8901,N_7790);
nor U10013 (N_10013,N_8640,N_8129);
nand U10014 (N_10014,N_7706,N_8259);
or U10015 (N_10015,N_7541,N_7924);
and U10016 (N_10016,N_8280,N_8774);
xor U10017 (N_10017,N_8446,N_8030);
and U10018 (N_10018,N_8692,N_8809);
and U10019 (N_10019,N_8683,N_8691);
xor U10020 (N_10020,N_8155,N_8431);
nor U10021 (N_10021,N_8704,N_8411);
and U10022 (N_10022,N_8129,N_8741);
or U10023 (N_10023,N_8254,N_8063);
or U10024 (N_10024,N_7865,N_8434);
nand U10025 (N_10025,N_7877,N_7725);
or U10026 (N_10026,N_8511,N_8214);
or U10027 (N_10027,N_8354,N_7861);
nor U10028 (N_10028,N_8473,N_8258);
xor U10029 (N_10029,N_7780,N_8404);
nor U10030 (N_10030,N_7660,N_8669);
xnor U10031 (N_10031,N_8068,N_8881);
nor U10032 (N_10032,N_8338,N_8832);
nand U10033 (N_10033,N_8012,N_8151);
or U10034 (N_10034,N_8901,N_8160);
nor U10035 (N_10035,N_8621,N_8729);
and U10036 (N_10036,N_8507,N_8234);
and U10037 (N_10037,N_7504,N_8851);
nor U10038 (N_10038,N_8741,N_7776);
xor U10039 (N_10039,N_7879,N_7851);
xnor U10040 (N_10040,N_8582,N_8944);
and U10041 (N_10041,N_8961,N_8240);
nor U10042 (N_10042,N_8687,N_8228);
nor U10043 (N_10043,N_7594,N_7653);
or U10044 (N_10044,N_7799,N_8224);
nor U10045 (N_10045,N_7774,N_8858);
or U10046 (N_10046,N_8041,N_7701);
xor U10047 (N_10047,N_8430,N_8550);
and U10048 (N_10048,N_7966,N_8550);
or U10049 (N_10049,N_7655,N_8244);
and U10050 (N_10050,N_8140,N_7503);
nor U10051 (N_10051,N_7841,N_8370);
or U10052 (N_10052,N_7509,N_8600);
nand U10053 (N_10053,N_8288,N_8948);
or U10054 (N_10054,N_8543,N_8947);
nand U10055 (N_10055,N_7853,N_8731);
and U10056 (N_10056,N_7660,N_7587);
and U10057 (N_10057,N_8195,N_8191);
nor U10058 (N_10058,N_8155,N_8776);
xnor U10059 (N_10059,N_8085,N_7933);
or U10060 (N_10060,N_8532,N_8663);
or U10061 (N_10061,N_8559,N_8148);
and U10062 (N_10062,N_8878,N_8278);
and U10063 (N_10063,N_8406,N_7555);
xnor U10064 (N_10064,N_8707,N_8533);
and U10065 (N_10065,N_8453,N_7643);
or U10066 (N_10066,N_7787,N_8845);
xnor U10067 (N_10067,N_8245,N_8189);
and U10068 (N_10068,N_8343,N_8982);
and U10069 (N_10069,N_7949,N_8770);
xnor U10070 (N_10070,N_8379,N_8609);
and U10071 (N_10071,N_8408,N_8189);
xor U10072 (N_10072,N_8802,N_7998);
xor U10073 (N_10073,N_8914,N_8281);
or U10074 (N_10074,N_8683,N_8855);
nand U10075 (N_10075,N_8933,N_7674);
nand U10076 (N_10076,N_8551,N_8319);
nor U10077 (N_10077,N_8582,N_8845);
xnor U10078 (N_10078,N_7589,N_8263);
nor U10079 (N_10079,N_8104,N_8054);
nor U10080 (N_10080,N_7914,N_8376);
nand U10081 (N_10081,N_7729,N_8455);
or U10082 (N_10082,N_8107,N_8036);
and U10083 (N_10083,N_8603,N_8771);
nor U10084 (N_10084,N_8579,N_7948);
nand U10085 (N_10085,N_8748,N_8632);
nand U10086 (N_10086,N_8076,N_8738);
xor U10087 (N_10087,N_8415,N_8584);
or U10088 (N_10088,N_8186,N_8417);
nor U10089 (N_10089,N_8627,N_7727);
xnor U10090 (N_10090,N_7636,N_7646);
nand U10091 (N_10091,N_8683,N_8279);
xnor U10092 (N_10092,N_7846,N_7982);
or U10093 (N_10093,N_8557,N_8533);
or U10094 (N_10094,N_7774,N_8797);
nor U10095 (N_10095,N_7998,N_8107);
and U10096 (N_10096,N_7817,N_7804);
nor U10097 (N_10097,N_8907,N_8623);
or U10098 (N_10098,N_8115,N_8091);
xnor U10099 (N_10099,N_8904,N_7909);
and U10100 (N_10100,N_8049,N_8042);
nor U10101 (N_10101,N_8867,N_8569);
nor U10102 (N_10102,N_8279,N_8150);
nor U10103 (N_10103,N_8473,N_7729);
xor U10104 (N_10104,N_8655,N_8904);
or U10105 (N_10105,N_7518,N_8570);
or U10106 (N_10106,N_7694,N_8557);
nor U10107 (N_10107,N_8876,N_8366);
and U10108 (N_10108,N_8145,N_7683);
and U10109 (N_10109,N_7643,N_8086);
xor U10110 (N_10110,N_7511,N_8144);
nand U10111 (N_10111,N_8381,N_7841);
nor U10112 (N_10112,N_8676,N_8096);
nand U10113 (N_10113,N_7778,N_8050);
and U10114 (N_10114,N_8558,N_8129);
or U10115 (N_10115,N_7792,N_7894);
or U10116 (N_10116,N_7550,N_7603);
nand U10117 (N_10117,N_7832,N_8281);
nand U10118 (N_10118,N_8873,N_8595);
nand U10119 (N_10119,N_8641,N_8833);
and U10120 (N_10120,N_8344,N_8799);
nor U10121 (N_10121,N_7581,N_8997);
xnor U10122 (N_10122,N_8232,N_8304);
xor U10123 (N_10123,N_8290,N_8989);
xnor U10124 (N_10124,N_8028,N_8851);
or U10125 (N_10125,N_7568,N_7616);
xor U10126 (N_10126,N_8288,N_8656);
xnor U10127 (N_10127,N_7929,N_8069);
and U10128 (N_10128,N_8843,N_8609);
nor U10129 (N_10129,N_8716,N_8606);
nor U10130 (N_10130,N_7735,N_7919);
or U10131 (N_10131,N_7721,N_8000);
or U10132 (N_10132,N_8465,N_8791);
nand U10133 (N_10133,N_8315,N_7929);
nand U10134 (N_10134,N_8538,N_7816);
xor U10135 (N_10135,N_8381,N_7600);
or U10136 (N_10136,N_8443,N_8265);
or U10137 (N_10137,N_8867,N_7869);
or U10138 (N_10138,N_7831,N_8325);
and U10139 (N_10139,N_8906,N_7668);
nand U10140 (N_10140,N_8475,N_8294);
or U10141 (N_10141,N_8083,N_7982);
and U10142 (N_10142,N_8777,N_8941);
nor U10143 (N_10143,N_8851,N_8987);
xnor U10144 (N_10144,N_8076,N_7577);
or U10145 (N_10145,N_7507,N_8522);
xnor U10146 (N_10146,N_8846,N_8580);
xnor U10147 (N_10147,N_8824,N_7728);
xor U10148 (N_10148,N_7560,N_7614);
and U10149 (N_10149,N_8809,N_8014);
nand U10150 (N_10150,N_7952,N_8751);
and U10151 (N_10151,N_8220,N_7991);
or U10152 (N_10152,N_8322,N_7601);
or U10153 (N_10153,N_8846,N_8383);
nor U10154 (N_10154,N_7890,N_8182);
nor U10155 (N_10155,N_8540,N_8518);
nand U10156 (N_10156,N_7710,N_8572);
or U10157 (N_10157,N_7520,N_8350);
or U10158 (N_10158,N_8046,N_8124);
and U10159 (N_10159,N_7777,N_7957);
nor U10160 (N_10160,N_8259,N_8312);
xnor U10161 (N_10161,N_8466,N_7666);
nor U10162 (N_10162,N_7870,N_7512);
and U10163 (N_10163,N_8820,N_8148);
nor U10164 (N_10164,N_8989,N_8918);
and U10165 (N_10165,N_7618,N_8429);
nor U10166 (N_10166,N_8501,N_7882);
nand U10167 (N_10167,N_7790,N_8960);
xor U10168 (N_10168,N_7685,N_8096);
or U10169 (N_10169,N_8983,N_8744);
nand U10170 (N_10170,N_8389,N_7925);
nor U10171 (N_10171,N_8827,N_8731);
nor U10172 (N_10172,N_8628,N_8815);
nand U10173 (N_10173,N_8724,N_8429);
nor U10174 (N_10174,N_8567,N_8421);
or U10175 (N_10175,N_8958,N_8001);
nand U10176 (N_10176,N_8594,N_8059);
xnor U10177 (N_10177,N_8238,N_8605);
nor U10178 (N_10178,N_8168,N_7503);
nand U10179 (N_10179,N_7833,N_7686);
nor U10180 (N_10180,N_8998,N_8266);
nand U10181 (N_10181,N_8500,N_7840);
nor U10182 (N_10182,N_8546,N_8593);
or U10183 (N_10183,N_8763,N_8025);
or U10184 (N_10184,N_8249,N_8463);
xor U10185 (N_10185,N_8267,N_8956);
xnor U10186 (N_10186,N_8007,N_8561);
xnor U10187 (N_10187,N_8326,N_8455);
or U10188 (N_10188,N_8352,N_7769);
xor U10189 (N_10189,N_8703,N_8147);
nor U10190 (N_10190,N_7785,N_7597);
or U10191 (N_10191,N_8765,N_8246);
nor U10192 (N_10192,N_8902,N_8014);
or U10193 (N_10193,N_8914,N_8538);
and U10194 (N_10194,N_7632,N_7804);
nand U10195 (N_10195,N_8390,N_8949);
and U10196 (N_10196,N_8862,N_8528);
and U10197 (N_10197,N_7572,N_7660);
nor U10198 (N_10198,N_8007,N_7730);
and U10199 (N_10199,N_7693,N_8752);
nand U10200 (N_10200,N_8023,N_8754);
and U10201 (N_10201,N_8922,N_8662);
nor U10202 (N_10202,N_7885,N_7864);
nor U10203 (N_10203,N_7643,N_7692);
xor U10204 (N_10204,N_7770,N_8844);
nand U10205 (N_10205,N_7841,N_8066);
nand U10206 (N_10206,N_8772,N_8330);
or U10207 (N_10207,N_8879,N_8633);
nor U10208 (N_10208,N_7596,N_7917);
nand U10209 (N_10209,N_7894,N_8046);
and U10210 (N_10210,N_8289,N_7747);
nand U10211 (N_10211,N_8251,N_8929);
and U10212 (N_10212,N_7849,N_8715);
nand U10213 (N_10213,N_8298,N_8461);
nor U10214 (N_10214,N_8596,N_8367);
nor U10215 (N_10215,N_7592,N_8370);
nand U10216 (N_10216,N_8715,N_7638);
xnor U10217 (N_10217,N_8950,N_8297);
or U10218 (N_10218,N_8892,N_8596);
and U10219 (N_10219,N_8087,N_7651);
nor U10220 (N_10220,N_7833,N_8412);
and U10221 (N_10221,N_8024,N_8975);
xnor U10222 (N_10222,N_8405,N_8291);
nand U10223 (N_10223,N_8392,N_8393);
and U10224 (N_10224,N_8349,N_8075);
and U10225 (N_10225,N_8313,N_7719);
and U10226 (N_10226,N_8391,N_8627);
and U10227 (N_10227,N_7996,N_7995);
xnor U10228 (N_10228,N_8375,N_8605);
nand U10229 (N_10229,N_7719,N_8290);
xnor U10230 (N_10230,N_7700,N_7736);
and U10231 (N_10231,N_7836,N_7745);
and U10232 (N_10232,N_8745,N_7760);
or U10233 (N_10233,N_7708,N_8969);
nand U10234 (N_10234,N_7602,N_8758);
and U10235 (N_10235,N_7870,N_8442);
xor U10236 (N_10236,N_8450,N_8816);
nor U10237 (N_10237,N_8866,N_8030);
or U10238 (N_10238,N_8239,N_7806);
nand U10239 (N_10239,N_7557,N_8723);
and U10240 (N_10240,N_7937,N_7840);
and U10241 (N_10241,N_8886,N_8118);
xnor U10242 (N_10242,N_8707,N_7602);
nor U10243 (N_10243,N_8355,N_8309);
xor U10244 (N_10244,N_8576,N_8217);
or U10245 (N_10245,N_7707,N_7883);
nor U10246 (N_10246,N_8917,N_7633);
nand U10247 (N_10247,N_8901,N_8100);
nand U10248 (N_10248,N_8252,N_8939);
xnor U10249 (N_10249,N_7537,N_7551);
xnor U10250 (N_10250,N_7969,N_8621);
xnor U10251 (N_10251,N_8906,N_7602);
nand U10252 (N_10252,N_8551,N_8304);
and U10253 (N_10253,N_8034,N_8533);
nor U10254 (N_10254,N_8227,N_8904);
xor U10255 (N_10255,N_8704,N_8105);
xor U10256 (N_10256,N_7685,N_8558);
and U10257 (N_10257,N_8745,N_8821);
nor U10258 (N_10258,N_8423,N_7782);
nand U10259 (N_10259,N_8343,N_8947);
and U10260 (N_10260,N_8480,N_8357);
nand U10261 (N_10261,N_8208,N_7572);
nand U10262 (N_10262,N_8692,N_8828);
nand U10263 (N_10263,N_8513,N_8930);
nand U10264 (N_10264,N_7647,N_7618);
xor U10265 (N_10265,N_8128,N_7683);
nor U10266 (N_10266,N_8096,N_8945);
and U10267 (N_10267,N_8783,N_8942);
nand U10268 (N_10268,N_8197,N_8615);
xnor U10269 (N_10269,N_7649,N_8294);
nand U10270 (N_10270,N_8128,N_7619);
xor U10271 (N_10271,N_8265,N_8768);
xnor U10272 (N_10272,N_8131,N_8290);
and U10273 (N_10273,N_7724,N_8511);
nor U10274 (N_10274,N_8476,N_7869);
or U10275 (N_10275,N_7982,N_7768);
xor U10276 (N_10276,N_8161,N_8397);
and U10277 (N_10277,N_8147,N_7922);
and U10278 (N_10278,N_7670,N_8896);
or U10279 (N_10279,N_8477,N_8547);
and U10280 (N_10280,N_8638,N_7936);
xnor U10281 (N_10281,N_8817,N_8078);
nor U10282 (N_10282,N_7966,N_7607);
or U10283 (N_10283,N_8640,N_8189);
nor U10284 (N_10284,N_8484,N_8221);
nor U10285 (N_10285,N_8207,N_8843);
xor U10286 (N_10286,N_8770,N_7567);
nor U10287 (N_10287,N_8578,N_8912);
nor U10288 (N_10288,N_8643,N_8520);
or U10289 (N_10289,N_8126,N_8486);
and U10290 (N_10290,N_7715,N_7931);
xor U10291 (N_10291,N_8675,N_7501);
xnor U10292 (N_10292,N_8691,N_7656);
nor U10293 (N_10293,N_8556,N_7725);
nand U10294 (N_10294,N_8438,N_8510);
xnor U10295 (N_10295,N_8172,N_7518);
xor U10296 (N_10296,N_8151,N_8894);
nor U10297 (N_10297,N_8141,N_7659);
nand U10298 (N_10298,N_8189,N_7580);
nand U10299 (N_10299,N_8423,N_8861);
xnor U10300 (N_10300,N_8660,N_8709);
and U10301 (N_10301,N_8506,N_7507);
nor U10302 (N_10302,N_8665,N_7711);
and U10303 (N_10303,N_8412,N_7907);
and U10304 (N_10304,N_7876,N_8550);
and U10305 (N_10305,N_8787,N_7560);
nor U10306 (N_10306,N_7602,N_7595);
xnor U10307 (N_10307,N_8002,N_7600);
and U10308 (N_10308,N_7653,N_8884);
or U10309 (N_10309,N_8514,N_8661);
xor U10310 (N_10310,N_8426,N_8166);
and U10311 (N_10311,N_7585,N_8017);
xnor U10312 (N_10312,N_7748,N_7763);
nor U10313 (N_10313,N_8807,N_7869);
nor U10314 (N_10314,N_7743,N_7909);
xnor U10315 (N_10315,N_8839,N_8199);
and U10316 (N_10316,N_8022,N_8477);
nand U10317 (N_10317,N_8478,N_8454);
xor U10318 (N_10318,N_8762,N_8430);
or U10319 (N_10319,N_7697,N_7837);
or U10320 (N_10320,N_7594,N_8663);
and U10321 (N_10321,N_8292,N_8597);
xnor U10322 (N_10322,N_8319,N_8792);
nor U10323 (N_10323,N_8057,N_7918);
or U10324 (N_10324,N_8853,N_8205);
and U10325 (N_10325,N_8101,N_8414);
nor U10326 (N_10326,N_8739,N_7592);
or U10327 (N_10327,N_8640,N_7919);
or U10328 (N_10328,N_8882,N_7946);
xnor U10329 (N_10329,N_7613,N_7709);
nand U10330 (N_10330,N_7823,N_7691);
and U10331 (N_10331,N_8414,N_8889);
xnor U10332 (N_10332,N_8569,N_8800);
or U10333 (N_10333,N_7899,N_8928);
nand U10334 (N_10334,N_8663,N_7704);
or U10335 (N_10335,N_8433,N_8213);
nor U10336 (N_10336,N_7688,N_8379);
or U10337 (N_10337,N_7868,N_8949);
xnor U10338 (N_10338,N_8636,N_8697);
or U10339 (N_10339,N_7754,N_8136);
xnor U10340 (N_10340,N_8964,N_7678);
nor U10341 (N_10341,N_7701,N_7656);
xor U10342 (N_10342,N_8870,N_8239);
xnor U10343 (N_10343,N_8807,N_8482);
nor U10344 (N_10344,N_8419,N_7743);
and U10345 (N_10345,N_8415,N_8569);
or U10346 (N_10346,N_8288,N_8867);
nor U10347 (N_10347,N_7542,N_7671);
and U10348 (N_10348,N_7811,N_7593);
nor U10349 (N_10349,N_8228,N_8174);
or U10350 (N_10350,N_7833,N_8783);
nand U10351 (N_10351,N_7588,N_8652);
xor U10352 (N_10352,N_8977,N_7568);
or U10353 (N_10353,N_7632,N_8126);
nor U10354 (N_10354,N_8525,N_8232);
xnor U10355 (N_10355,N_7953,N_8413);
or U10356 (N_10356,N_7599,N_7869);
xnor U10357 (N_10357,N_8129,N_7758);
nand U10358 (N_10358,N_7789,N_8378);
nor U10359 (N_10359,N_7507,N_8988);
or U10360 (N_10360,N_8445,N_8952);
or U10361 (N_10361,N_8978,N_7566);
nand U10362 (N_10362,N_8918,N_8916);
xor U10363 (N_10363,N_7683,N_8888);
nor U10364 (N_10364,N_8076,N_8864);
xor U10365 (N_10365,N_8886,N_8536);
xor U10366 (N_10366,N_7949,N_7753);
or U10367 (N_10367,N_7818,N_7562);
xor U10368 (N_10368,N_8986,N_7714);
and U10369 (N_10369,N_8887,N_8743);
xnor U10370 (N_10370,N_8278,N_7986);
and U10371 (N_10371,N_8077,N_8367);
or U10372 (N_10372,N_8395,N_8256);
and U10373 (N_10373,N_8354,N_8794);
and U10374 (N_10374,N_8526,N_7849);
nor U10375 (N_10375,N_7879,N_8626);
or U10376 (N_10376,N_8310,N_8547);
or U10377 (N_10377,N_8849,N_7629);
nand U10378 (N_10378,N_8605,N_8794);
and U10379 (N_10379,N_8244,N_7892);
or U10380 (N_10380,N_8558,N_7509);
xor U10381 (N_10381,N_8956,N_7589);
xnor U10382 (N_10382,N_7838,N_8793);
nand U10383 (N_10383,N_8345,N_8043);
and U10384 (N_10384,N_8490,N_7508);
and U10385 (N_10385,N_7559,N_7942);
nand U10386 (N_10386,N_8486,N_8890);
nor U10387 (N_10387,N_7779,N_7943);
xor U10388 (N_10388,N_7815,N_8392);
and U10389 (N_10389,N_8436,N_8411);
and U10390 (N_10390,N_8485,N_8845);
or U10391 (N_10391,N_7545,N_7902);
xnor U10392 (N_10392,N_8234,N_8800);
nor U10393 (N_10393,N_7658,N_7881);
nand U10394 (N_10394,N_8386,N_8496);
or U10395 (N_10395,N_7923,N_8760);
or U10396 (N_10396,N_8331,N_8838);
and U10397 (N_10397,N_8515,N_8510);
nand U10398 (N_10398,N_8950,N_8885);
or U10399 (N_10399,N_7608,N_7511);
or U10400 (N_10400,N_8924,N_8179);
and U10401 (N_10401,N_7932,N_7969);
or U10402 (N_10402,N_7952,N_7817);
or U10403 (N_10403,N_7922,N_8578);
nand U10404 (N_10404,N_7844,N_8471);
and U10405 (N_10405,N_7581,N_7613);
nand U10406 (N_10406,N_8807,N_7984);
and U10407 (N_10407,N_8492,N_8373);
nor U10408 (N_10408,N_7699,N_7910);
nor U10409 (N_10409,N_8468,N_8218);
nor U10410 (N_10410,N_7603,N_7821);
or U10411 (N_10411,N_8482,N_7833);
xnor U10412 (N_10412,N_8119,N_8818);
nor U10413 (N_10413,N_8931,N_8470);
or U10414 (N_10414,N_7953,N_8286);
nand U10415 (N_10415,N_8048,N_7858);
or U10416 (N_10416,N_8917,N_8413);
xor U10417 (N_10417,N_8951,N_8415);
nor U10418 (N_10418,N_7590,N_8251);
or U10419 (N_10419,N_8537,N_8303);
nor U10420 (N_10420,N_7607,N_7949);
or U10421 (N_10421,N_8498,N_7846);
xor U10422 (N_10422,N_8993,N_8945);
nor U10423 (N_10423,N_8385,N_7594);
or U10424 (N_10424,N_8703,N_8522);
nor U10425 (N_10425,N_7624,N_8372);
or U10426 (N_10426,N_8381,N_8266);
nor U10427 (N_10427,N_7573,N_8392);
and U10428 (N_10428,N_8388,N_8027);
xnor U10429 (N_10429,N_8454,N_8169);
nand U10430 (N_10430,N_8324,N_7699);
xor U10431 (N_10431,N_8258,N_8282);
nand U10432 (N_10432,N_8362,N_8826);
xnor U10433 (N_10433,N_7768,N_8423);
xnor U10434 (N_10434,N_7980,N_7649);
nor U10435 (N_10435,N_7813,N_7713);
xor U10436 (N_10436,N_7785,N_7507);
and U10437 (N_10437,N_7928,N_8000);
nand U10438 (N_10438,N_8863,N_7613);
or U10439 (N_10439,N_7755,N_8687);
or U10440 (N_10440,N_8470,N_8223);
nor U10441 (N_10441,N_8519,N_8793);
nor U10442 (N_10442,N_8349,N_7963);
and U10443 (N_10443,N_8300,N_8387);
or U10444 (N_10444,N_8190,N_7874);
nor U10445 (N_10445,N_7852,N_7532);
or U10446 (N_10446,N_8266,N_8173);
or U10447 (N_10447,N_8049,N_8756);
nand U10448 (N_10448,N_7672,N_8334);
nor U10449 (N_10449,N_7760,N_8853);
nor U10450 (N_10450,N_7921,N_8481);
xor U10451 (N_10451,N_8590,N_8023);
and U10452 (N_10452,N_8118,N_8460);
xnor U10453 (N_10453,N_7985,N_8316);
nand U10454 (N_10454,N_8168,N_7773);
or U10455 (N_10455,N_8666,N_7853);
and U10456 (N_10456,N_8332,N_8852);
xor U10457 (N_10457,N_8468,N_8767);
and U10458 (N_10458,N_8548,N_7997);
xor U10459 (N_10459,N_8099,N_8004);
and U10460 (N_10460,N_8907,N_8415);
nand U10461 (N_10461,N_7533,N_7780);
nand U10462 (N_10462,N_8896,N_7517);
xnor U10463 (N_10463,N_7676,N_8579);
or U10464 (N_10464,N_7638,N_8352);
nor U10465 (N_10465,N_8297,N_8629);
nor U10466 (N_10466,N_7531,N_8019);
and U10467 (N_10467,N_8536,N_7615);
nor U10468 (N_10468,N_7741,N_7999);
nand U10469 (N_10469,N_8221,N_8433);
xor U10470 (N_10470,N_8173,N_8386);
xor U10471 (N_10471,N_8598,N_8529);
nand U10472 (N_10472,N_8069,N_8854);
or U10473 (N_10473,N_7817,N_8705);
nand U10474 (N_10474,N_8059,N_8944);
nand U10475 (N_10475,N_8183,N_8765);
xor U10476 (N_10476,N_7548,N_8355);
nor U10477 (N_10477,N_8140,N_8754);
and U10478 (N_10478,N_8116,N_7779);
and U10479 (N_10479,N_8050,N_8275);
nor U10480 (N_10480,N_8513,N_8413);
and U10481 (N_10481,N_8391,N_7598);
nand U10482 (N_10482,N_8329,N_8840);
xnor U10483 (N_10483,N_8025,N_8942);
xor U10484 (N_10484,N_7777,N_8452);
nor U10485 (N_10485,N_8233,N_8855);
or U10486 (N_10486,N_7839,N_8255);
nor U10487 (N_10487,N_8422,N_8467);
nand U10488 (N_10488,N_8515,N_8622);
or U10489 (N_10489,N_7763,N_8273);
and U10490 (N_10490,N_7538,N_7719);
or U10491 (N_10491,N_8962,N_8564);
nand U10492 (N_10492,N_8696,N_8435);
nand U10493 (N_10493,N_7883,N_7584);
nor U10494 (N_10494,N_8726,N_7799);
and U10495 (N_10495,N_8727,N_8678);
nor U10496 (N_10496,N_8314,N_7633);
or U10497 (N_10497,N_8239,N_8480);
and U10498 (N_10498,N_7508,N_8363);
nor U10499 (N_10499,N_8954,N_8664);
nand U10500 (N_10500,N_10292,N_9819);
nand U10501 (N_10501,N_9318,N_9433);
and U10502 (N_10502,N_9117,N_9578);
nand U10503 (N_10503,N_9376,N_10400);
and U10504 (N_10504,N_9983,N_9229);
nand U10505 (N_10505,N_9100,N_9539);
nor U10506 (N_10506,N_9803,N_9021);
xnor U10507 (N_10507,N_9381,N_9604);
nand U10508 (N_10508,N_10397,N_10326);
nand U10509 (N_10509,N_9617,N_10383);
xor U10510 (N_10510,N_9715,N_9032);
nor U10511 (N_10511,N_9847,N_9927);
xnor U10512 (N_10512,N_10165,N_9861);
or U10513 (N_10513,N_9203,N_9115);
or U10514 (N_10514,N_10078,N_10461);
and U10515 (N_10515,N_9120,N_9002);
or U10516 (N_10516,N_9190,N_9896);
xnor U10517 (N_10517,N_9828,N_10142);
or U10518 (N_10518,N_9742,N_9736);
and U10519 (N_10519,N_10258,N_9790);
and U10520 (N_10520,N_9471,N_10191);
or U10521 (N_10521,N_9659,N_9406);
nor U10522 (N_10522,N_9633,N_9294);
nand U10523 (N_10523,N_10216,N_9375);
and U10524 (N_10524,N_9152,N_9603);
and U10525 (N_10525,N_9958,N_10232);
or U10526 (N_10526,N_10371,N_10441);
xor U10527 (N_10527,N_9883,N_9220);
nor U10528 (N_10528,N_9254,N_9587);
nor U10529 (N_10529,N_10422,N_10040);
and U10530 (N_10530,N_10217,N_10331);
xnor U10531 (N_10531,N_9218,N_9372);
or U10532 (N_10532,N_10032,N_9174);
nand U10533 (N_10533,N_9399,N_10457);
or U10534 (N_10534,N_10474,N_9078);
nand U10535 (N_10535,N_9644,N_9760);
xnor U10536 (N_10536,N_9669,N_10025);
xnor U10537 (N_10537,N_9003,N_10027);
nand U10538 (N_10538,N_9223,N_9501);
and U10539 (N_10539,N_9682,N_9383);
and U10540 (N_10540,N_10442,N_9188);
or U10541 (N_10541,N_9343,N_10072);
xnor U10542 (N_10542,N_10269,N_9425);
or U10543 (N_10543,N_9873,N_9573);
nand U10544 (N_10544,N_9692,N_10486);
xor U10545 (N_10545,N_9072,N_10396);
nor U10546 (N_10546,N_9065,N_9206);
and U10547 (N_10547,N_10263,N_9080);
nor U10548 (N_10548,N_9811,N_10021);
and U10549 (N_10549,N_10398,N_9976);
and U10550 (N_10550,N_9909,N_9332);
and U10551 (N_10551,N_10446,N_9673);
nor U10552 (N_10552,N_9066,N_9582);
nand U10553 (N_10553,N_9487,N_9470);
nand U10554 (N_10554,N_10332,N_9815);
nor U10555 (N_10555,N_10384,N_9794);
nor U10556 (N_10556,N_9562,N_9747);
xor U10557 (N_10557,N_9805,N_10096);
nand U10558 (N_10558,N_10162,N_10494);
xnor U10559 (N_10559,N_10117,N_9738);
and U10560 (N_10560,N_9986,N_10133);
and U10561 (N_10561,N_9102,N_9314);
nor U10562 (N_10562,N_9391,N_10039);
nor U10563 (N_10563,N_10158,N_9639);
nand U10564 (N_10564,N_9018,N_9311);
and U10565 (N_10565,N_10024,N_10427);
xnor U10566 (N_10566,N_9952,N_10315);
and U10567 (N_10567,N_9169,N_9288);
or U10568 (N_10568,N_10282,N_9774);
nand U10569 (N_10569,N_9557,N_9723);
and U10570 (N_10570,N_10256,N_9729);
nor U10571 (N_10571,N_10083,N_9704);
nor U10572 (N_10572,N_10219,N_9705);
or U10573 (N_10573,N_10174,N_10353);
or U10574 (N_10574,N_9610,N_9154);
xor U10575 (N_10575,N_9429,N_9697);
nand U10576 (N_10576,N_10112,N_9473);
and U10577 (N_10577,N_9313,N_9533);
xor U10578 (N_10578,N_10048,N_10073);
or U10579 (N_10579,N_9276,N_9139);
xor U10580 (N_10580,N_9933,N_9205);
nor U10581 (N_10581,N_9296,N_10336);
nor U10582 (N_10582,N_9202,N_9567);
xnor U10583 (N_10583,N_9106,N_9667);
nor U10584 (N_10584,N_9676,N_9595);
and U10585 (N_10585,N_10028,N_9367);
nand U10586 (N_10586,N_10119,N_9784);
nor U10587 (N_10587,N_9321,N_9920);
xor U10588 (N_10588,N_9163,N_10321);
xor U10589 (N_10589,N_9849,N_9108);
nor U10590 (N_10590,N_9802,N_9387);
and U10591 (N_10591,N_10405,N_10118);
nor U10592 (N_10592,N_9962,N_9484);
and U10593 (N_10593,N_9428,N_9778);
and U10594 (N_10594,N_9486,N_9678);
nor U10595 (N_10595,N_10190,N_9044);
and U10596 (N_10596,N_10064,N_9488);
or U10597 (N_10597,N_10287,N_9431);
nor U10598 (N_10598,N_9224,N_9377);
nor U10599 (N_10599,N_9073,N_10199);
or U10600 (N_10600,N_9545,N_10387);
xor U10601 (N_10601,N_9326,N_10401);
xnor U10602 (N_10602,N_9445,N_10068);
xnor U10603 (N_10603,N_9892,N_9137);
nor U10604 (N_10604,N_9170,N_9565);
xor U10605 (N_10605,N_9750,N_9325);
nor U10606 (N_10606,N_9746,N_9996);
xnor U10607 (N_10607,N_9404,N_9788);
nand U10608 (N_10608,N_9273,N_9081);
nand U10609 (N_10609,N_10140,N_9505);
xor U10610 (N_10610,N_10276,N_10323);
nor U10611 (N_10611,N_9845,N_9623);
or U10612 (N_10612,N_9358,N_9319);
nor U10613 (N_10613,N_9987,N_10286);
nor U10614 (N_10614,N_9140,N_10128);
or U10615 (N_10615,N_9625,N_9439);
nand U10616 (N_10616,N_9159,N_9844);
xor U10617 (N_10617,N_9010,N_9193);
nor U10618 (N_10618,N_9379,N_9440);
or U10619 (N_10619,N_10380,N_9960);
and U10620 (N_10620,N_9878,N_10409);
xor U10621 (N_10621,N_10430,N_9568);
and U10622 (N_10622,N_10322,N_9123);
or U10623 (N_10623,N_10000,N_10364);
nand U10624 (N_10624,N_9558,N_10333);
nor U10625 (N_10625,N_10127,N_10469);
and U10626 (N_10626,N_9171,N_9918);
nand U10627 (N_10627,N_9212,N_9201);
xor U10628 (N_10628,N_9700,N_9852);
xnor U10629 (N_10629,N_10221,N_9300);
nand U10630 (N_10630,N_9219,N_9214);
and U10631 (N_10631,N_9025,N_9243);
nor U10632 (N_10632,N_9907,N_10490);
and U10633 (N_10633,N_10202,N_10359);
and U10634 (N_10634,N_9011,N_10186);
and U10635 (N_10635,N_9055,N_10463);
and U10636 (N_10636,N_9616,N_9506);
or U10637 (N_10637,N_9244,N_10204);
nor U10638 (N_10638,N_10223,N_9683);
xor U10639 (N_10639,N_10077,N_9238);
or U10640 (N_10640,N_10339,N_9248);
and U10641 (N_10641,N_9129,N_10376);
or U10642 (N_10642,N_9999,N_9782);
xnor U10643 (N_10643,N_10407,N_10374);
nor U10644 (N_10644,N_9196,N_9001);
xnor U10645 (N_10645,N_9030,N_9923);
nor U10646 (N_10646,N_9405,N_10420);
nor U10647 (N_10647,N_9540,N_9753);
and U10648 (N_10648,N_9773,N_9324);
and U10649 (N_10649,N_9088,N_9458);
nand U10650 (N_10650,N_9929,N_9452);
and U10651 (N_10651,N_9004,N_9037);
nor U10652 (N_10652,N_10355,N_9831);
or U10653 (N_10653,N_9624,N_9327);
nand U10654 (N_10654,N_10370,N_9389);
nand U10655 (N_10655,N_9530,N_9880);
nand U10656 (N_10656,N_9368,N_10379);
xor U10657 (N_10657,N_9531,N_9369);
or U10658 (N_10658,N_10498,N_9741);
and U10659 (N_10659,N_9752,N_9620);
and U10660 (N_10660,N_9413,N_9974);
or U10661 (N_10661,N_9510,N_9841);
and U10662 (N_10662,N_10145,N_9083);
nand U10663 (N_10663,N_9519,N_9813);
nor U10664 (N_10664,N_9945,N_10134);
nor U10665 (N_10665,N_9019,N_10449);
nor U10666 (N_10666,N_9550,N_9045);
nand U10667 (N_10667,N_10260,N_9434);
and U10668 (N_10668,N_9396,N_10382);
nor U10669 (N_10669,N_9270,N_9232);
nor U10670 (N_10670,N_10470,N_10104);
and U10671 (N_10671,N_10002,N_9971);
and U10672 (N_10672,N_9643,N_9581);
xor U10673 (N_10673,N_9076,N_9717);
nor U10674 (N_10674,N_10302,N_9577);
xor U10675 (N_10675,N_9937,N_9121);
nor U10676 (N_10676,N_10460,N_9951);
and U10677 (N_10677,N_10121,N_9257);
nand U10678 (N_10678,N_10168,N_10488);
nor U10679 (N_10679,N_9725,N_9442);
nor U10680 (N_10680,N_9580,N_10419);
and U10681 (N_10681,N_9388,N_9972);
nand U10682 (N_10682,N_10054,N_10154);
and U10683 (N_10683,N_9928,N_10088);
xor U10684 (N_10684,N_9652,N_9417);
nor U10685 (N_10685,N_9259,N_9598);
or U10686 (N_10686,N_9876,N_10106);
nor U10687 (N_10687,N_9733,N_10171);
nor U10688 (N_10688,N_10259,N_9146);
nor U10689 (N_10689,N_10307,N_9204);
nor U10690 (N_10690,N_10099,N_9251);
and U10691 (N_10691,N_9503,N_10246);
xnor U10692 (N_10692,N_10212,N_9973);
xor U10693 (N_10693,N_9386,N_9908);
or U10694 (N_10694,N_9284,N_9754);
nor U10695 (N_10695,N_9250,N_9593);
or U10696 (N_10696,N_9240,N_9661);
or U10697 (N_10697,N_10185,N_10319);
nor U10698 (N_10698,N_9082,N_10176);
nand U10699 (N_10699,N_10354,N_10362);
xor U10700 (N_10700,N_9013,N_9990);
xor U10701 (N_10701,N_9299,N_10139);
nor U10702 (N_10702,N_10147,N_10464);
xor U10703 (N_10703,N_9921,N_10055);
and U10704 (N_10704,N_9810,N_9077);
or U10705 (N_10705,N_10426,N_9268);
nand U10706 (N_10706,N_9217,N_10489);
nand U10707 (N_10707,N_10479,N_9925);
and U10708 (N_10708,N_9247,N_10350);
or U10709 (N_10709,N_10043,N_9427);
or U10710 (N_10710,N_9655,N_10241);
nand U10711 (N_10711,N_9838,N_9776);
nor U10712 (N_10712,N_9791,N_9910);
and U10713 (N_10713,N_9104,N_10492);
nor U10714 (N_10714,N_9511,N_9069);
xor U10715 (N_10715,N_9895,N_9561);
or U10716 (N_10716,N_10472,N_9096);
nand U10717 (N_10717,N_10141,N_9969);
nand U10718 (N_10718,N_10338,N_9239);
and U10719 (N_10719,N_9517,N_10455);
nand U10720 (N_10720,N_10136,N_9820);
and U10721 (N_10721,N_9571,N_9160);
nand U10722 (N_10722,N_9144,N_9767);
nand U10723 (N_10723,N_9543,N_10225);
and U10724 (N_10724,N_9830,N_9266);
or U10725 (N_10725,N_9267,N_9320);
xnor U10726 (N_10726,N_9789,N_10238);
nand U10727 (N_10727,N_9843,N_9832);
nor U10728 (N_10728,N_9063,N_10310);
nand U10729 (N_10729,N_9863,N_9640);
or U10730 (N_10730,N_9265,N_10063);
nor U10731 (N_10731,N_9353,N_9615);
and U10732 (N_10732,N_9521,N_9614);
and U10733 (N_10733,N_9913,N_9946);
nor U10734 (N_10734,N_9197,N_10095);
nand U10735 (N_10735,N_9411,N_10081);
nor U10736 (N_10736,N_10074,N_10208);
nor U10737 (N_10737,N_9961,N_9835);
nand U10738 (N_10738,N_10229,N_9891);
and U10739 (N_10739,N_9138,N_10318);
or U10740 (N_10740,N_9443,N_9457);
or U10741 (N_10741,N_10428,N_9061);
nand U10742 (N_10742,N_9674,N_9438);
nand U10743 (N_10743,N_9315,N_9497);
nand U10744 (N_10744,N_9017,N_9936);
xnor U10745 (N_10745,N_9529,N_9829);
and U10746 (N_10746,N_10448,N_10497);
nor U10747 (N_10747,N_9415,N_10007);
xor U10748 (N_10748,N_10248,N_9304);
xnor U10749 (N_10749,N_9708,N_9498);
or U10750 (N_10750,N_9934,N_10042);
or U10751 (N_10751,N_9119,N_10393);
nand U10752 (N_10752,N_9357,N_9028);
or U10753 (N_10753,N_9978,N_9074);
or U10754 (N_10754,N_9000,N_9619);
or U10755 (N_10755,N_10161,N_9341);
or U10756 (N_10756,N_10148,N_9477);
nor U10757 (N_10757,N_9950,N_9956);
or U10758 (N_10758,N_9173,N_10451);
or U10759 (N_10759,N_9134,N_9964);
and U10760 (N_10760,N_9221,N_9448);
xnor U10761 (N_10761,N_10423,N_10218);
nor U10762 (N_10762,N_9101,N_10080);
xor U10763 (N_10763,N_10102,N_10456);
and U10764 (N_10764,N_9185,N_9801);
xnor U10765 (N_10765,N_9600,N_9275);
nand U10766 (N_10766,N_9485,N_9271);
nand U10767 (N_10767,N_9014,N_9097);
xor U10768 (N_10768,N_10358,N_9762);
nand U10769 (N_10769,N_9260,N_9085);
nor U10770 (N_10770,N_9766,N_9869);
or U10771 (N_10771,N_9574,N_9730);
or U10772 (N_10772,N_10316,N_9351);
nand U10773 (N_10773,N_9131,N_9851);
and U10774 (N_10774,N_9435,N_10004);
xnor U10775 (N_10775,N_9594,N_9356);
nand U10776 (N_10776,N_9671,N_10014);
nand U10777 (N_10777,N_10485,N_9544);
xnor U10778 (N_10778,N_10361,N_10325);
nor U10779 (N_10779,N_9982,N_10299);
nand U10780 (N_10780,N_10335,N_9666);
and U10781 (N_10781,N_10312,N_10167);
xnor U10782 (N_10782,N_9105,N_9157);
nand U10783 (N_10783,N_9938,N_10372);
or U10784 (N_10784,N_10010,N_10352);
or U10785 (N_10785,N_9775,N_9126);
nand U10786 (N_10786,N_10105,N_9043);
and U10787 (N_10787,N_10107,N_9191);
xor U10788 (N_10788,N_10347,N_10421);
or U10789 (N_10789,N_9068,N_9451);
xor U10790 (N_10790,N_10130,N_9309);
and U10791 (N_10791,N_9226,N_9542);
nor U10792 (N_10792,N_9227,N_10293);
or U10793 (N_10793,N_10245,N_9513);
xor U10794 (N_10794,N_9493,N_9397);
nor U10795 (N_10795,N_10045,N_9153);
nand U10796 (N_10796,N_9524,N_9207);
nor U10797 (N_10797,N_9344,N_10329);
nand U10798 (N_10798,N_9359,N_10473);
nor U10799 (N_10799,N_9716,N_9461);
nor U10800 (N_10800,N_9366,N_9349);
xnor U10801 (N_10801,N_10151,N_9967);
or U10802 (N_10802,N_10035,N_10041);
or U10803 (N_10803,N_9904,N_9162);
nor U10804 (N_10804,N_9350,N_9328);
or U10805 (N_10805,N_10327,N_9648);
nor U10806 (N_10806,N_9899,N_9371);
nand U10807 (N_10807,N_10023,N_9049);
nand U10808 (N_10808,N_10179,N_9302);
and U10809 (N_10809,N_9935,N_9823);
and U10810 (N_10810,N_9208,N_9165);
xor U10811 (N_10811,N_10275,N_9817);
xnor U10812 (N_10812,N_9979,N_9145);
nand U10813 (N_10813,N_10252,N_9148);
and U10814 (N_10814,N_10018,N_9130);
nor U10815 (N_10815,N_9086,N_10163);
and U10816 (N_10816,N_10328,N_9155);
nand U10817 (N_10817,N_9618,N_10373);
nor U10818 (N_10818,N_10062,N_9739);
nor U10819 (N_10819,N_9881,N_10126);
nor U10820 (N_10820,N_9884,N_9732);
and U10821 (N_10821,N_10052,N_9491);
or U10822 (N_10822,N_9476,N_9256);
and U10823 (N_10823,N_9418,N_9720);
or U10824 (N_10824,N_9807,N_9702);
or U10825 (N_10825,N_9283,N_9382);
nor U10826 (N_10826,N_9797,N_9585);
nand U10827 (N_10827,N_9213,N_9981);
xor U10828 (N_10828,N_9871,N_10349);
nand U10829 (N_10829,N_10075,N_9589);
nand U10830 (N_10830,N_9826,N_9555);
or U10831 (N_10831,N_10173,N_10155);
nor U10832 (N_10832,N_9735,N_9612);
nand U10833 (N_10833,N_9424,N_10272);
nor U10834 (N_10834,N_9308,N_10187);
xnor U10835 (N_10835,N_9989,N_10069);
nor U10836 (N_10836,N_10006,N_9184);
and U10837 (N_10837,N_9111,N_9164);
nand U10838 (N_10838,N_9384,N_9740);
or U10839 (N_10839,N_10255,N_9809);
and U10840 (N_10840,N_10305,N_9690);
nand U10841 (N_10841,N_9274,N_10411);
and U10842 (N_10842,N_10109,N_9727);
nand U10843 (N_10843,N_10091,N_9930);
nand U10844 (N_10844,N_9701,N_9412);
xnor U10845 (N_10845,N_9850,N_10012);
xor U10846 (N_10846,N_9495,N_9575);
nor U10847 (N_10847,N_9877,N_10342);
and U10848 (N_10848,N_9804,N_9834);
nand U10849 (N_10849,N_10233,N_9158);
xnor U10850 (N_10850,N_9998,N_9919);
and U10851 (N_10851,N_9970,N_10029);
nand U10852 (N_10852,N_10424,N_9479);
and U10853 (N_10853,N_9020,N_9997);
xnor U10854 (N_10854,N_10297,N_9355);
and U10855 (N_10855,N_9765,N_10468);
nor U10856 (N_10856,N_9955,N_9722);
and U10857 (N_10857,N_9903,N_9363);
xor U10858 (N_10858,N_9005,N_9711);
nand U10859 (N_10859,N_10070,N_10476);
and U10860 (N_10860,N_10390,N_9535);
and U10861 (N_10861,N_10159,N_9514);
and U10862 (N_10862,N_10237,N_10434);
nand U10863 (N_10863,N_9024,N_9291);
nor U10864 (N_10864,N_9772,N_9954);
and U10865 (N_10865,N_9756,N_9520);
nor U10866 (N_10866,N_10435,N_9475);
nand U10867 (N_10867,N_9922,N_9052);
nor U10868 (N_10868,N_10235,N_9179);
nand U10869 (N_10869,N_9109,N_10129);
and U10870 (N_10870,N_9125,N_9712);
nand U10871 (N_10871,N_9337,N_10381);
nor U10872 (N_10872,N_10280,N_10125);
and U10873 (N_10873,N_9241,N_10164);
xor U10874 (N_10874,N_9912,N_10429);
xor U10875 (N_10875,N_9305,N_10357);
or U10876 (N_10876,N_9657,N_9348);
or U10877 (N_10877,N_9079,N_10298);
and U10878 (N_10878,N_10443,N_10416);
or U10879 (N_10879,N_9286,N_9637);
or U10880 (N_10880,N_9113,N_9761);
or U10881 (N_10881,N_9222,N_9649);
nand U10882 (N_10882,N_9679,N_9340);
nand U10883 (N_10883,N_9848,N_9507);
nor U10884 (N_10884,N_9691,N_10089);
nand U10885 (N_10885,N_9398,N_9818);
nand U10886 (N_10886,N_10182,N_9446);
nand U10887 (N_10887,N_9898,N_9882);
or U10888 (N_10888,N_10487,N_9792);
nand U10889 (N_10889,N_9062,N_9602);
xor U10890 (N_10890,N_10022,N_9093);
xor U10891 (N_10891,N_10399,N_9846);
xor U10892 (N_10892,N_9480,N_9576);
xor U10893 (N_10893,N_9658,N_9734);
or U10894 (N_10894,N_10412,N_9749);
nor U10895 (N_10895,N_9454,N_10076);
xnor U10896 (N_10896,N_10279,N_9075);
nand U10897 (N_10897,N_10092,N_9868);
xor U10898 (N_10898,N_10013,N_10211);
xnor U10899 (N_10899,N_9168,N_9855);
and U10900 (N_10900,N_9133,N_10153);
nor U10901 (N_10901,N_10183,N_9632);
xnor U10902 (N_10902,N_9149,N_9806);
or U10903 (N_10903,N_10239,N_9499);
and U10904 (N_10904,N_9569,N_9858);
xnor U10905 (N_10905,N_9686,N_9401);
xor U10906 (N_10906,N_9675,N_10224);
nand U10907 (N_10907,N_10348,N_10471);
nor U10908 (N_10908,N_9862,N_10122);
and U10909 (N_10909,N_9916,N_9837);
nor U10910 (N_10910,N_10200,N_9629);
nand U10911 (N_10911,N_10261,N_10184);
nand U10912 (N_10912,N_9795,N_9006);
and U10913 (N_10913,N_10392,N_9410);
and U10914 (N_10914,N_10213,N_10295);
and U10915 (N_10915,N_9246,N_9768);
xnor U10916 (N_10916,N_9465,N_9853);
xnor U10917 (N_10917,N_10031,N_10491);
xor U10918 (N_10918,N_9748,N_9022);
and U10919 (N_10919,N_9988,N_9474);
nand U10920 (N_10920,N_9255,N_9242);
nand U10921 (N_10921,N_9180,N_10444);
nand U10922 (N_10922,N_10100,N_10300);
and U10923 (N_10923,N_10047,N_9258);
nand U10924 (N_10924,N_10222,N_10466);
nor U10925 (N_10925,N_9127,N_9360);
xor U10926 (N_10926,N_9769,N_10138);
or U10927 (N_10927,N_9780,N_10116);
nor U10928 (N_10928,N_9745,N_9609);
nand U10929 (N_10929,N_9293,N_9685);
and U10930 (N_10930,N_10137,N_10493);
or U10931 (N_10931,N_9161,N_9995);
nand U10932 (N_10932,N_9588,N_10437);
nor U10933 (N_10933,N_9546,N_9426);
and U10934 (N_10934,N_10196,N_9630);
or U10935 (N_10935,N_9572,N_10389);
nor U10936 (N_10936,N_10236,N_9894);
or U10937 (N_10937,N_9634,N_9508);
nor U10938 (N_10938,N_9210,N_9622);
or U10939 (N_10939,N_9586,N_9627);
and U10940 (N_10940,N_9195,N_9905);
and U10941 (N_10941,N_10368,N_9347);
nand U10942 (N_10942,N_9089,N_9516);
nand U10943 (N_10943,N_9036,N_9867);
xor U10944 (N_10944,N_10367,N_9796);
xor U10945 (N_10945,N_10417,N_10090);
xnor U10946 (N_10946,N_9092,N_9352);
or U10947 (N_10947,N_9541,N_9468);
nand U10948 (N_10948,N_9114,N_10240);
nand U10949 (N_10949,N_10250,N_9591);
nor U10950 (N_10950,N_9714,N_10017);
or U10951 (N_10951,N_9570,N_9890);
nor U10952 (N_10952,N_10330,N_9538);
nor U10953 (N_10953,N_10378,N_9755);
or U10954 (N_10954,N_9249,N_10049);
nor U10955 (N_10955,N_9166,N_9500);
or U10956 (N_10956,N_9141,N_9663);
or U10957 (N_10957,N_9422,N_10169);
or U10958 (N_10958,N_9502,N_9306);
nor U10959 (N_10959,N_10231,N_9728);
and U10960 (N_10960,N_9118,N_10290);
nor U10961 (N_10961,N_9211,N_9023);
xor U10962 (N_10962,N_10103,N_9719);
xor U10963 (N_10963,N_10085,N_10243);
xor U10964 (N_10964,N_9653,N_9966);
nand U10965 (N_10965,N_10046,N_10150);
and U10966 (N_10966,N_10135,N_9940);
xnor U10967 (N_10967,N_9393,N_9509);
or U10968 (N_10968,N_9525,N_9628);
xnor U10969 (N_10969,N_10281,N_9112);
and U10970 (N_10970,N_9447,N_9482);
nor U10971 (N_10971,N_9060,N_9449);
nand U10972 (N_10972,N_9551,N_9994);
xnor U10973 (N_10973,N_9726,N_9307);
nor U10974 (N_10974,N_9459,N_9186);
and U10975 (N_10975,N_10160,N_9414);
or U10976 (N_10976,N_9054,N_9606);
nand U10977 (N_10977,N_9668,N_10317);
xnor U10978 (N_10978,N_10195,N_10360);
or U10979 (N_10979,N_10496,N_10016);
and U10980 (N_10980,N_9590,N_9699);
xnor U10981 (N_10981,N_10477,N_10257);
and U10982 (N_10982,N_9504,N_9469);
or U10983 (N_10983,N_10386,N_9605);
nor U10984 (N_10984,N_9943,N_10084);
nand U10985 (N_10985,N_9303,N_9527);
and U10986 (N_10986,N_9116,N_10178);
xor U10987 (N_10987,N_10101,N_10066);
nor U10988 (N_10988,N_9751,N_10345);
and U10989 (N_10989,N_9333,N_9216);
xnor U10990 (N_10990,N_9345,N_10266);
or U10991 (N_10991,N_9948,N_10111);
or U10992 (N_10992,N_9911,N_9301);
and U10993 (N_10993,N_9887,N_10194);
or U10994 (N_10994,N_9464,N_9462);
nand U10995 (N_10995,N_9385,N_9039);
nand U10996 (N_10996,N_10108,N_10273);
and U10997 (N_10997,N_9931,N_10205);
xor U10998 (N_10998,N_9365,N_9875);
or U10999 (N_10999,N_10253,N_9825);
and U11000 (N_11000,N_9793,N_9057);
nor U11001 (N_11001,N_10115,N_9378);
or U11002 (N_11002,N_9087,N_9395);
nand U11003 (N_11003,N_9537,N_9472);
xnor U11004 (N_11004,N_10026,N_10277);
xnor U11005 (N_11005,N_10306,N_9338);
xor U11006 (N_11006,N_10459,N_9403);
xnor U11007 (N_11007,N_9430,N_10020);
nor U11008 (N_11008,N_9178,N_9698);
or U11009 (N_11009,N_9407,N_10439);
xnor U11010 (N_11010,N_9941,N_10267);
nor U11011 (N_11011,N_9566,N_9584);
xor U11012 (N_11012,N_9143,N_9613);
nand U11013 (N_11013,N_10341,N_9432);
xor U11014 (N_11014,N_9053,N_10061);
nor U11015 (N_11015,N_9985,N_9737);
nor U11016 (N_11016,N_9654,N_9135);
xnor U11017 (N_11017,N_9489,N_10220);
xor U11018 (N_11018,N_9770,N_10431);
nor U11019 (N_11019,N_9522,N_9230);
xor U11020 (N_11020,N_10283,N_10056);
nand U11021 (N_11021,N_9122,N_10037);
nor U11022 (N_11022,N_10475,N_10123);
and U11023 (N_11023,N_9263,N_9786);
xnor U11024 (N_11024,N_9007,N_9090);
and U11025 (N_11025,N_9703,N_9785);
or U11026 (N_11026,N_9031,N_9707);
or U11027 (N_11027,N_10450,N_10452);
or U11028 (N_11028,N_9084,N_9015);
xor U11029 (N_11029,N_9554,N_10193);
and U11030 (N_11030,N_9175,N_10086);
xnor U11031 (N_11031,N_10403,N_10499);
xor U11032 (N_11032,N_10465,N_9638);
nor U11033 (N_11033,N_9957,N_9436);
nor U11034 (N_11034,N_10408,N_10278);
nand U11035 (N_11035,N_10447,N_9842);
and U11036 (N_11036,N_10036,N_9099);
xor U11037 (N_11037,N_9695,N_9490);
nand U11038 (N_11038,N_9893,N_9731);
and U11039 (N_11039,N_10192,N_10156);
and U11040 (N_11040,N_9646,N_9548);
xor U11041 (N_11041,N_9362,N_10203);
xor U11042 (N_11042,N_9317,N_9346);
or U11043 (N_11043,N_10304,N_9900);
nor U11044 (N_11044,N_9225,N_9380);
and U11045 (N_11045,N_9824,N_9650);
and U11046 (N_11046,N_10414,N_9860);
and U11047 (N_11047,N_9423,N_10303);
xor U11048 (N_11048,N_10180,N_9496);
nand U11049 (N_11049,N_9949,N_9947);
or U11050 (N_11050,N_10288,N_9743);
nand U11051 (N_11051,N_10410,N_10177);
nor U11052 (N_11052,N_10265,N_9902);
or U11053 (N_11053,N_9800,N_9110);
xor U11054 (N_11054,N_9253,N_10008);
or U11055 (N_11055,N_9336,N_9295);
nand U11056 (N_11056,N_10270,N_10458);
nor U11057 (N_11057,N_9827,N_9744);
or U11058 (N_11058,N_10207,N_10454);
or U11059 (N_11059,N_9771,N_9664);
or U11060 (N_11060,N_9012,N_9237);
and U11061 (N_11061,N_10467,N_9579);
nand U11062 (N_11062,N_10244,N_10097);
or U11063 (N_11063,N_9416,N_9709);
and U11064 (N_11064,N_9787,N_9132);
xor U11065 (N_11065,N_9528,N_9854);
nor U11066 (N_11066,N_10478,N_10189);
nand U11067 (N_11067,N_9559,N_9444);
or U11068 (N_11068,N_9687,N_10284);
and U11069 (N_11069,N_10226,N_9656);
nand U11070 (N_11070,N_9035,N_9187);
xnor U11071 (N_11071,N_9512,N_9156);
nor U11072 (N_11072,N_10314,N_9058);
nor U11073 (N_11073,N_10132,N_9536);
xor U11074 (N_11074,N_10363,N_9269);
nand U11075 (N_11075,N_9050,N_9812);
nor U11076 (N_11076,N_9836,N_9136);
nand U11077 (N_11077,N_9840,N_10425);
and U11078 (N_11078,N_9886,N_9635);
or U11079 (N_11079,N_9151,N_10149);
xor U11080 (N_11080,N_9042,N_9051);
or U11081 (N_11081,N_9932,N_10172);
xnor U11082 (N_11082,N_9724,N_10120);
or U11083 (N_11083,N_10079,N_9287);
xor U11084 (N_11084,N_9693,N_9901);
nor U11085 (N_11085,N_10311,N_10071);
nor U11086 (N_11086,N_9394,N_10495);
and U11087 (N_11087,N_9942,N_10197);
or U11088 (N_11088,N_9200,N_9182);
xor U11089 (N_11089,N_9665,N_9597);
or U11090 (N_11090,N_10188,N_9859);
and U11091 (N_11091,N_9879,N_10344);
or U11092 (N_11092,N_9041,N_10483);
or U11093 (N_11093,N_9917,N_9331);
nor U11094 (N_11094,N_9515,N_10356);
and U11095 (N_11095,N_10143,N_10124);
nor U11096 (N_11096,N_9526,N_10413);
xor U11097 (N_11097,N_9549,N_10215);
or U11098 (N_11098,N_9292,N_9798);
nor U11099 (N_11099,N_10249,N_9993);
or U11100 (N_11100,N_10206,N_9124);
nand U11101 (N_11101,N_10210,N_9272);
or U11102 (N_11102,N_9681,N_9611);
xor U11103 (N_11103,N_10059,N_10481);
nor U11104 (N_11104,N_10175,N_9915);
xnor U11105 (N_11105,N_9906,N_9642);
xnor U11106 (N_11106,N_9215,N_10289);
and U11107 (N_11107,N_10087,N_9980);
xor U11108 (N_11108,N_10227,N_10462);
nand U11109 (N_11109,N_9560,N_9523);
and U11110 (N_11110,N_10234,N_10009);
and U11111 (N_11111,N_9601,N_9888);
and U11112 (N_11112,N_9189,N_10131);
nand U11113 (N_11113,N_9285,N_9494);
nor U11114 (N_11114,N_9563,N_9518);
and U11115 (N_11115,N_10053,N_9252);
nand U11116 (N_11116,N_9183,N_9339);
nand U11117 (N_11117,N_9781,N_9027);
or U11118 (N_11118,N_9390,N_9298);
and U11119 (N_11119,N_9064,N_9583);
nand U11120 (N_11120,N_10377,N_9924);
or U11121 (N_11121,N_9047,N_9329);
and U11122 (N_11122,N_9764,N_10058);
nor U11123 (N_11123,N_10242,N_9091);
and U11124 (N_11124,N_10011,N_9370);
nor U11125 (N_11125,N_10001,N_9672);
or U11126 (N_11126,N_9534,N_9323);
or U11127 (N_11127,N_9354,N_9874);
nand U11128 (N_11128,N_9779,N_10337);
or U11129 (N_11129,N_10324,N_10296);
and U11130 (N_11130,N_9437,N_9278);
nand U11131 (N_11131,N_9689,N_9872);
and U11132 (N_11132,N_9297,N_10098);
nor U11133 (N_11133,N_9680,N_10438);
and U11134 (N_11134,N_9467,N_9763);
xnor U11135 (N_11135,N_9492,N_9564);
nor U11136 (N_11136,N_9865,N_9071);
nor U11137 (N_11137,N_9944,N_9670);
and U11138 (N_11138,N_10251,N_9450);
nor U11139 (N_11139,N_9277,N_9977);
or U11140 (N_11140,N_9289,N_10313);
and U11141 (N_11141,N_9310,N_9290);
and U11142 (N_11142,N_9660,N_9280);
and U11143 (N_11143,N_10114,N_9926);
or U11144 (N_11144,N_9478,N_10262);
xor U11145 (N_11145,N_9713,N_10484);
nand U11146 (N_11146,N_9056,N_10271);
or U11147 (N_11147,N_10230,N_9710);
nor U11148 (N_11148,N_9889,N_9177);
nor U11149 (N_11149,N_10294,N_10365);
nand U11150 (N_11150,N_9696,N_10157);
xnor U11151 (N_11151,N_10440,N_9552);
or U11152 (N_11152,N_10285,N_9194);
nor U11153 (N_11153,N_9463,N_9409);
nor U11154 (N_11154,N_10094,N_9857);
and U11155 (N_11155,N_10343,N_9953);
nor U11156 (N_11156,N_10264,N_9322);
nand U11157 (N_11157,N_10051,N_10201);
and U11158 (N_11158,N_9335,N_10065);
and U11159 (N_11159,N_9233,N_10057);
nand U11160 (N_11160,N_9647,N_9150);
and U11161 (N_11161,N_9532,N_9199);
or U11162 (N_11162,N_10067,N_10369);
xnor U11163 (N_11163,N_10030,N_9261);
xnor U11164 (N_11164,N_9455,N_10247);
nor U11165 (N_11165,N_10198,N_9334);
nand U11166 (N_11166,N_9777,N_9816);
or U11167 (N_11167,N_10453,N_9626);
nand U11168 (N_11168,N_9034,N_9621);
xnor U11169 (N_11169,N_10170,N_10385);
nand U11170 (N_11170,N_9968,N_10375);
xnor U11171 (N_11171,N_10274,N_9419);
and U11172 (N_11172,N_9839,N_10050);
and U11173 (N_11173,N_9758,N_9592);
or U11174 (N_11174,N_9651,N_9706);
nor U11175 (N_11175,N_9984,N_9420);
and U11176 (N_11176,N_10301,N_9677);
nor U11177 (N_11177,N_10146,N_9599);
or U11178 (N_11178,N_9556,N_9172);
nor U11179 (N_11179,N_9026,N_9098);
xor U11180 (N_11180,N_9181,N_9421);
xnor U11181 (N_11181,N_9059,N_9759);
and U11182 (N_11182,N_9822,N_9821);
xnor U11183 (N_11183,N_9342,N_10395);
nand U11184 (N_11184,N_9107,N_10334);
nand U11185 (N_11185,N_9094,N_9176);
or U11186 (N_11186,N_9799,N_9373);
nand U11187 (N_11187,N_10019,N_9228);
xnor U11188 (N_11188,N_9808,N_10015);
or U11189 (N_11189,N_10308,N_10388);
xnor U11190 (N_11190,N_10093,N_9688);
and U11191 (N_11191,N_10320,N_10366);
or U11192 (N_11192,N_9959,N_10038);
nand U11193 (N_11193,N_9236,N_9048);
nand U11194 (N_11194,N_9279,N_10406);
nor U11195 (N_11195,N_9636,N_9198);
and U11196 (N_11196,N_9264,N_9965);
and U11197 (N_11197,N_10228,N_9870);
or U11198 (N_11198,N_9453,N_10418);
or U11199 (N_11199,N_10480,N_10033);
xor U11200 (N_11200,N_9312,N_9067);
nor U11201 (N_11201,N_10415,N_9833);
nor U11202 (N_11202,N_9374,N_9040);
and U11203 (N_11203,N_9466,N_10391);
nor U11204 (N_11204,N_9033,N_9645);
nor U11205 (N_11205,N_9757,N_9608);
nand U11206 (N_11206,N_9596,N_9281);
nand U11207 (N_11207,N_9262,N_9897);
nand U11208 (N_11208,N_10268,N_10110);
nor U11209 (N_11209,N_9316,N_9330);
nor U11210 (N_11210,N_9481,N_9364);
or U11211 (N_11211,N_9209,N_10166);
nor U11212 (N_11212,N_9547,N_9641);
or U11213 (N_11213,N_9009,N_9885);
nor U11214 (N_11214,N_10433,N_9914);
xor U11215 (N_11215,N_10340,N_9142);
and U11216 (N_11216,N_9553,N_9483);
xor U11217 (N_11217,N_10113,N_10309);
or U11218 (N_11218,N_10402,N_10060);
and U11219 (N_11219,N_9234,N_9046);
xnor U11220 (N_11220,N_9392,N_9460);
or U11221 (N_11221,N_9245,N_10346);
nor U11222 (N_11222,N_9231,N_10005);
or U11223 (N_11223,N_10209,N_10482);
xor U11224 (N_11224,N_10291,N_10003);
xor U11225 (N_11225,N_9856,N_9939);
or U11226 (N_11226,N_10152,N_9814);
nand U11227 (N_11227,N_10144,N_9095);
xnor U11228 (N_11228,N_9029,N_9864);
nand U11229 (N_11229,N_9103,N_9402);
or U11230 (N_11230,N_9721,N_9783);
or U11231 (N_11231,N_9282,N_10404);
nor U11232 (N_11232,N_9456,N_9192);
and U11233 (N_11233,N_9408,N_9167);
xnor U11234 (N_11234,N_10436,N_9992);
xnor U11235 (N_11235,N_9016,N_9694);
and U11236 (N_11236,N_9975,N_9400);
or U11237 (N_11237,N_10181,N_10394);
nand U11238 (N_11238,N_10214,N_10254);
xor U11239 (N_11239,N_9038,N_10351);
and U11240 (N_11240,N_9662,N_9991);
xnor U11241 (N_11241,N_9718,N_10432);
or U11242 (N_11242,N_10082,N_9963);
or U11243 (N_11243,N_9441,N_10044);
nor U11244 (N_11244,N_9684,N_9235);
nor U11245 (N_11245,N_9361,N_10034);
nand U11246 (N_11246,N_9008,N_9866);
xnor U11247 (N_11247,N_10445,N_9631);
or U11248 (N_11248,N_9147,N_9128);
xnor U11249 (N_11249,N_9607,N_9070);
xnor U11250 (N_11250,N_9622,N_9647);
xnor U11251 (N_11251,N_9423,N_9598);
nand U11252 (N_11252,N_9073,N_9892);
nand U11253 (N_11253,N_9705,N_9847);
nor U11254 (N_11254,N_10472,N_9824);
nand U11255 (N_11255,N_9339,N_10377);
and U11256 (N_11256,N_9281,N_9062);
nand U11257 (N_11257,N_9312,N_10017);
nor U11258 (N_11258,N_10495,N_10239);
nor U11259 (N_11259,N_9278,N_9609);
and U11260 (N_11260,N_10470,N_9451);
and U11261 (N_11261,N_10210,N_10492);
nor U11262 (N_11262,N_10010,N_10458);
xor U11263 (N_11263,N_9419,N_9403);
xor U11264 (N_11264,N_9898,N_9318);
xnor U11265 (N_11265,N_10233,N_9679);
or U11266 (N_11266,N_10416,N_9291);
nor U11267 (N_11267,N_10306,N_9272);
and U11268 (N_11268,N_10048,N_10360);
nor U11269 (N_11269,N_9880,N_9977);
or U11270 (N_11270,N_9759,N_9541);
and U11271 (N_11271,N_9880,N_10009);
and U11272 (N_11272,N_9966,N_9744);
nor U11273 (N_11273,N_10080,N_10069);
or U11274 (N_11274,N_10312,N_10141);
nor U11275 (N_11275,N_10329,N_9071);
and U11276 (N_11276,N_10477,N_9587);
nand U11277 (N_11277,N_9991,N_9179);
and U11278 (N_11278,N_9464,N_9965);
and U11279 (N_11279,N_9456,N_9870);
and U11280 (N_11280,N_9207,N_10260);
nor U11281 (N_11281,N_9734,N_9776);
or U11282 (N_11282,N_9880,N_10143);
and U11283 (N_11283,N_9051,N_9480);
and U11284 (N_11284,N_9461,N_10005);
and U11285 (N_11285,N_10345,N_9718);
nor U11286 (N_11286,N_10370,N_9685);
nand U11287 (N_11287,N_9517,N_10415);
or U11288 (N_11288,N_9820,N_9923);
nor U11289 (N_11289,N_10333,N_10463);
and U11290 (N_11290,N_10433,N_10093);
nand U11291 (N_11291,N_9245,N_10238);
nor U11292 (N_11292,N_9869,N_9609);
nand U11293 (N_11293,N_9406,N_9195);
and U11294 (N_11294,N_10230,N_10425);
nand U11295 (N_11295,N_9222,N_10387);
or U11296 (N_11296,N_9326,N_9005);
xor U11297 (N_11297,N_9336,N_10381);
nand U11298 (N_11298,N_9215,N_10009);
or U11299 (N_11299,N_9708,N_10147);
nand U11300 (N_11300,N_9028,N_9034);
nor U11301 (N_11301,N_10201,N_10412);
xnor U11302 (N_11302,N_9864,N_9161);
and U11303 (N_11303,N_9977,N_9828);
nand U11304 (N_11304,N_9124,N_9731);
and U11305 (N_11305,N_9338,N_9767);
nand U11306 (N_11306,N_9420,N_9293);
or U11307 (N_11307,N_10482,N_10190);
xor U11308 (N_11308,N_9322,N_9797);
nand U11309 (N_11309,N_9818,N_9417);
xnor U11310 (N_11310,N_9580,N_10389);
nand U11311 (N_11311,N_9597,N_9687);
nor U11312 (N_11312,N_9403,N_9424);
and U11313 (N_11313,N_9963,N_10319);
nand U11314 (N_11314,N_9303,N_10259);
nor U11315 (N_11315,N_9104,N_9774);
nor U11316 (N_11316,N_10247,N_10377);
nor U11317 (N_11317,N_9359,N_9807);
nor U11318 (N_11318,N_9805,N_10383);
and U11319 (N_11319,N_10210,N_9313);
or U11320 (N_11320,N_9681,N_10435);
nor U11321 (N_11321,N_9975,N_9887);
and U11322 (N_11322,N_9665,N_9230);
or U11323 (N_11323,N_9524,N_10291);
nor U11324 (N_11324,N_10300,N_10160);
nand U11325 (N_11325,N_10131,N_9627);
and U11326 (N_11326,N_9138,N_9932);
or U11327 (N_11327,N_9948,N_10274);
xnor U11328 (N_11328,N_10488,N_9001);
and U11329 (N_11329,N_9174,N_9702);
xnor U11330 (N_11330,N_9150,N_9106);
nor U11331 (N_11331,N_9952,N_10033);
nor U11332 (N_11332,N_9158,N_10297);
nand U11333 (N_11333,N_9673,N_10428);
or U11334 (N_11334,N_10498,N_9697);
and U11335 (N_11335,N_10135,N_9985);
and U11336 (N_11336,N_9921,N_9392);
and U11337 (N_11337,N_9203,N_9798);
nor U11338 (N_11338,N_9220,N_9459);
nand U11339 (N_11339,N_9310,N_10386);
xor U11340 (N_11340,N_9307,N_9935);
or U11341 (N_11341,N_10318,N_9284);
nor U11342 (N_11342,N_10427,N_10476);
nor U11343 (N_11343,N_9442,N_10333);
nand U11344 (N_11344,N_10303,N_9877);
and U11345 (N_11345,N_9876,N_9914);
nand U11346 (N_11346,N_9666,N_10491);
or U11347 (N_11347,N_9942,N_10201);
nand U11348 (N_11348,N_9181,N_10471);
and U11349 (N_11349,N_10110,N_9513);
and U11350 (N_11350,N_9300,N_9669);
nor U11351 (N_11351,N_9866,N_9643);
or U11352 (N_11352,N_9975,N_10118);
nor U11353 (N_11353,N_9313,N_9074);
or U11354 (N_11354,N_9000,N_9186);
nand U11355 (N_11355,N_9272,N_10414);
xnor U11356 (N_11356,N_10415,N_9220);
nand U11357 (N_11357,N_9886,N_9505);
xor U11358 (N_11358,N_10396,N_10495);
xor U11359 (N_11359,N_10050,N_10436);
nor U11360 (N_11360,N_10127,N_9941);
nand U11361 (N_11361,N_9746,N_10207);
nor U11362 (N_11362,N_9110,N_9347);
nand U11363 (N_11363,N_9167,N_9164);
or U11364 (N_11364,N_9073,N_9925);
and U11365 (N_11365,N_9449,N_10447);
xor U11366 (N_11366,N_10165,N_9526);
nand U11367 (N_11367,N_9549,N_9578);
nand U11368 (N_11368,N_9160,N_9761);
xor U11369 (N_11369,N_9838,N_9704);
nor U11370 (N_11370,N_9514,N_10095);
or U11371 (N_11371,N_9000,N_9691);
xor U11372 (N_11372,N_10272,N_9865);
and U11373 (N_11373,N_9526,N_9998);
nand U11374 (N_11374,N_10101,N_9621);
or U11375 (N_11375,N_10196,N_10208);
nor U11376 (N_11376,N_9933,N_9310);
nor U11377 (N_11377,N_10404,N_10027);
nand U11378 (N_11378,N_9728,N_10195);
xor U11379 (N_11379,N_9316,N_10261);
nor U11380 (N_11380,N_10211,N_10422);
nor U11381 (N_11381,N_10278,N_10375);
nand U11382 (N_11382,N_9353,N_9358);
and U11383 (N_11383,N_9713,N_10392);
xor U11384 (N_11384,N_9079,N_10239);
xor U11385 (N_11385,N_9596,N_9932);
nor U11386 (N_11386,N_9290,N_9317);
xnor U11387 (N_11387,N_9821,N_9289);
nand U11388 (N_11388,N_10474,N_9697);
xnor U11389 (N_11389,N_10320,N_9976);
nor U11390 (N_11390,N_9204,N_10402);
and U11391 (N_11391,N_9218,N_9355);
nand U11392 (N_11392,N_9982,N_10005);
nor U11393 (N_11393,N_9638,N_10369);
and U11394 (N_11394,N_10314,N_9356);
nand U11395 (N_11395,N_9490,N_10491);
xnor U11396 (N_11396,N_9794,N_9018);
nand U11397 (N_11397,N_9469,N_9219);
nor U11398 (N_11398,N_9193,N_9842);
and U11399 (N_11399,N_9636,N_10338);
and U11400 (N_11400,N_9242,N_9719);
nor U11401 (N_11401,N_9963,N_9162);
nor U11402 (N_11402,N_9469,N_9335);
and U11403 (N_11403,N_10287,N_10414);
or U11404 (N_11404,N_10431,N_9330);
and U11405 (N_11405,N_10403,N_10232);
and U11406 (N_11406,N_9441,N_9720);
nand U11407 (N_11407,N_9318,N_10169);
or U11408 (N_11408,N_9941,N_9749);
xnor U11409 (N_11409,N_10007,N_9582);
xnor U11410 (N_11410,N_10019,N_10191);
nor U11411 (N_11411,N_10250,N_10277);
nand U11412 (N_11412,N_10312,N_9604);
or U11413 (N_11413,N_9955,N_10221);
nand U11414 (N_11414,N_10488,N_10414);
nand U11415 (N_11415,N_9989,N_9675);
nor U11416 (N_11416,N_9438,N_10168);
nand U11417 (N_11417,N_9530,N_9082);
or U11418 (N_11418,N_9988,N_9670);
nor U11419 (N_11419,N_9717,N_9604);
nor U11420 (N_11420,N_9973,N_9069);
nand U11421 (N_11421,N_9750,N_9159);
nand U11422 (N_11422,N_10251,N_10070);
xor U11423 (N_11423,N_9411,N_10352);
nand U11424 (N_11424,N_9857,N_9273);
and U11425 (N_11425,N_9943,N_9681);
xnor U11426 (N_11426,N_9019,N_10351);
nand U11427 (N_11427,N_9415,N_9409);
nand U11428 (N_11428,N_10153,N_9674);
xor U11429 (N_11429,N_9387,N_9682);
and U11430 (N_11430,N_9369,N_10398);
or U11431 (N_11431,N_9390,N_9417);
nand U11432 (N_11432,N_10401,N_10333);
or U11433 (N_11433,N_10395,N_9534);
or U11434 (N_11434,N_10117,N_10202);
and U11435 (N_11435,N_9226,N_9273);
nor U11436 (N_11436,N_10431,N_9005);
xor U11437 (N_11437,N_9387,N_9394);
nor U11438 (N_11438,N_9756,N_10172);
or U11439 (N_11439,N_9252,N_9580);
or U11440 (N_11440,N_9708,N_9645);
or U11441 (N_11441,N_9789,N_9949);
nor U11442 (N_11442,N_9498,N_9389);
xor U11443 (N_11443,N_9982,N_9241);
and U11444 (N_11444,N_9967,N_10373);
nand U11445 (N_11445,N_9384,N_10253);
nor U11446 (N_11446,N_10019,N_10489);
or U11447 (N_11447,N_9725,N_10330);
or U11448 (N_11448,N_9755,N_10311);
or U11449 (N_11449,N_9979,N_10400);
or U11450 (N_11450,N_10277,N_9904);
and U11451 (N_11451,N_9310,N_9186);
or U11452 (N_11452,N_9229,N_10200);
and U11453 (N_11453,N_10417,N_9013);
and U11454 (N_11454,N_9857,N_9255);
xnor U11455 (N_11455,N_10462,N_9077);
and U11456 (N_11456,N_9148,N_9223);
and U11457 (N_11457,N_9536,N_9734);
or U11458 (N_11458,N_9836,N_10257);
nand U11459 (N_11459,N_9611,N_10167);
or U11460 (N_11460,N_9009,N_10333);
xor U11461 (N_11461,N_9383,N_9749);
nor U11462 (N_11462,N_9953,N_10230);
nor U11463 (N_11463,N_10185,N_10400);
nand U11464 (N_11464,N_9330,N_10204);
and U11465 (N_11465,N_10420,N_9053);
xor U11466 (N_11466,N_9823,N_9461);
nor U11467 (N_11467,N_9364,N_9050);
nand U11468 (N_11468,N_9740,N_9469);
and U11469 (N_11469,N_10225,N_9089);
and U11470 (N_11470,N_10362,N_10251);
nor U11471 (N_11471,N_9015,N_10116);
nand U11472 (N_11472,N_10085,N_10050);
nor U11473 (N_11473,N_9839,N_10414);
or U11474 (N_11474,N_10070,N_10186);
nor U11475 (N_11475,N_9519,N_10317);
and U11476 (N_11476,N_9331,N_9086);
xnor U11477 (N_11477,N_9531,N_10292);
and U11478 (N_11478,N_9969,N_10366);
xor U11479 (N_11479,N_9896,N_10432);
nor U11480 (N_11480,N_9818,N_9142);
xnor U11481 (N_11481,N_9829,N_9033);
nand U11482 (N_11482,N_10314,N_9478);
and U11483 (N_11483,N_10465,N_9843);
nand U11484 (N_11484,N_9683,N_9571);
or U11485 (N_11485,N_10471,N_10115);
or U11486 (N_11486,N_10278,N_9978);
nor U11487 (N_11487,N_9960,N_9573);
xnor U11488 (N_11488,N_9665,N_9776);
and U11489 (N_11489,N_10361,N_9347);
and U11490 (N_11490,N_9873,N_9549);
xor U11491 (N_11491,N_10238,N_10482);
nand U11492 (N_11492,N_10473,N_9358);
nor U11493 (N_11493,N_9594,N_9259);
and U11494 (N_11494,N_9842,N_9103);
nor U11495 (N_11495,N_9211,N_10084);
nor U11496 (N_11496,N_9352,N_10125);
or U11497 (N_11497,N_9618,N_9406);
nor U11498 (N_11498,N_10256,N_10425);
nand U11499 (N_11499,N_9058,N_10373);
and U11500 (N_11500,N_9211,N_9160);
and U11501 (N_11501,N_9548,N_10369);
nand U11502 (N_11502,N_10069,N_9882);
nor U11503 (N_11503,N_10254,N_9142);
xnor U11504 (N_11504,N_9373,N_9099);
and U11505 (N_11505,N_10277,N_10334);
or U11506 (N_11506,N_9025,N_9427);
xor U11507 (N_11507,N_10461,N_9122);
xor U11508 (N_11508,N_9920,N_9150);
and U11509 (N_11509,N_10393,N_9792);
and U11510 (N_11510,N_9483,N_9857);
nor U11511 (N_11511,N_9850,N_10287);
and U11512 (N_11512,N_9234,N_9092);
xor U11513 (N_11513,N_9729,N_9414);
xnor U11514 (N_11514,N_9325,N_9776);
and U11515 (N_11515,N_9085,N_9652);
or U11516 (N_11516,N_10011,N_10193);
nand U11517 (N_11517,N_10116,N_9076);
nand U11518 (N_11518,N_10264,N_9774);
and U11519 (N_11519,N_10315,N_9914);
xor U11520 (N_11520,N_9244,N_9124);
nor U11521 (N_11521,N_9680,N_9355);
nand U11522 (N_11522,N_9226,N_9977);
nor U11523 (N_11523,N_9176,N_9777);
nand U11524 (N_11524,N_9244,N_9608);
xnor U11525 (N_11525,N_10232,N_9248);
nor U11526 (N_11526,N_9285,N_9422);
nor U11527 (N_11527,N_9740,N_10309);
nor U11528 (N_11528,N_10480,N_9565);
nand U11529 (N_11529,N_9806,N_10003);
or U11530 (N_11530,N_10303,N_10339);
and U11531 (N_11531,N_9908,N_9307);
or U11532 (N_11532,N_9178,N_9320);
xnor U11533 (N_11533,N_9838,N_10296);
or U11534 (N_11534,N_9502,N_9700);
xor U11535 (N_11535,N_9148,N_9059);
nor U11536 (N_11536,N_10107,N_10301);
xor U11537 (N_11537,N_9582,N_9252);
and U11538 (N_11538,N_9709,N_10478);
xnor U11539 (N_11539,N_9572,N_9389);
or U11540 (N_11540,N_9329,N_9750);
and U11541 (N_11541,N_10481,N_9317);
and U11542 (N_11542,N_9370,N_9561);
or U11543 (N_11543,N_10149,N_9061);
xor U11544 (N_11544,N_10182,N_10211);
and U11545 (N_11545,N_9088,N_10412);
or U11546 (N_11546,N_10059,N_9827);
nand U11547 (N_11547,N_9214,N_10256);
nand U11548 (N_11548,N_9833,N_9168);
nand U11549 (N_11549,N_9367,N_9218);
nor U11550 (N_11550,N_9342,N_10299);
or U11551 (N_11551,N_9094,N_9045);
xnor U11552 (N_11552,N_10372,N_10165);
nand U11553 (N_11553,N_9139,N_9084);
nor U11554 (N_11554,N_10076,N_10091);
nand U11555 (N_11555,N_10412,N_10385);
nor U11556 (N_11556,N_9567,N_9490);
and U11557 (N_11557,N_9259,N_10317);
nor U11558 (N_11558,N_9551,N_10313);
xnor U11559 (N_11559,N_9753,N_9873);
xor U11560 (N_11560,N_9570,N_9806);
or U11561 (N_11561,N_9302,N_9886);
and U11562 (N_11562,N_9205,N_9672);
and U11563 (N_11563,N_9039,N_9945);
nand U11564 (N_11564,N_9919,N_9055);
nor U11565 (N_11565,N_10496,N_9957);
nand U11566 (N_11566,N_10244,N_10231);
and U11567 (N_11567,N_9835,N_9834);
xnor U11568 (N_11568,N_9417,N_9996);
xnor U11569 (N_11569,N_10223,N_9426);
or U11570 (N_11570,N_9849,N_9424);
and U11571 (N_11571,N_9082,N_9253);
or U11572 (N_11572,N_10419,N_9078);
xnor U11573 (N_11573,N_10160,N_10047);
xnor U11574 (N_11574,N_9296,N_9508);
xor U11575 (N_11575,N_10428,N_10338);
nor U11576 (N_11576,N_9276,N_9315);
and U11577 (N_11577,N_10324,N_10102);
nand U11578 (N_11578,N_10114,N_10378);
nor U11579 (N_11579,N_9839,N_10017);
nand U11580 (N_11580,N_9647,N_9550);
nor U11581 (N_11581,N_10285,N_9074);
and U11582 (N_11582,N_9246,N_9581);
and U11583 (N_11583,N_10021,N_9054);
or U11584 (N_11584,N_10120,N_9230);
nor U11585 (N_11585,N_9724,N_10324);
nand U11586 (N_11586,N_9464,N_9636);
xor U11587 (N_11587,N_9295,N_9712);
nand U11588 (N_11588,N_9663,N_10175);
or U11589 (N_11589,N_9543,N_9664);
or U11590 (N_11590,N_9167,N_9701);
nor U11591 (N_11591,N_10061,N_10371);
and U11592 (N_11592,N_10285,N_10051);
xor U11593 (N_11593,N_10356,N_10298);
nor U11594 (N_11594,N_9696,N_9743);
and U11595 (N_11595,N_10286,N_9077);
or U11596 (N_11596,N_9554,N_9952);
nand U11597 (N_11597,N_9827,N_9959);
and U11598 (N_11598,N_10039,N_10495);
nand U11599 (N_11599,N_10213,N_10237);
xor U11600 (N_11600,N_10376,N_9642);
xor U11601 (N_11601,N_9870,N_10477);
nand U11602 (N_11602,N_9855,N_9565);
xor U11603 (N_11603,N_10394,N_9677);
xnor U11604 (N_11604,N_10450,N_9183);
nor U11605 (N_11605,N_9048,N_10130);
nand U11606 (N_11606,N_9955,N_9676);
and U11607 (N_11607,N_10093,N_10235);
nand U11608 (N_11608,N_9379,N_10454);
xnor U11609 (N_11609,N_10119,N_9739);
xor U11610 (N_11610,N_9648,N_10240);
and U11611 (N_11611,N_10132,N_9012);
nand U11612 (N_11612,N_9315,N_10130);
and U11613 (N_11613,N_9261,N_9914);
or U11614 (N_11614,N_9274,N_9010);
and U11615 (N_11615,N_9419,N_10407);
and U11616 (N_11616,N_9716,N_9031);
nor U11617 (N_11617,N_9969,N_9353);
nor U11618 (N_11618,N_9954,N_10489);
xnor U11619 (N_11619,N_9285,N_9154);
and U11620 (N_11620,N_9944,N_9107);
and U11621 (N_11621,N_9900,N_9484);
and U11622 (N_11622,N_9909,N_9690);
nand U11623 (N_11623,N_9533,N_10078);
and U11624 (N_11624,N_10337,N_9977);
nor U11625 (N_11625,N_10341,N_9996);
or U11626 (N_11626,N_9194,N_10278);
or U11627 (N_11627,N_9924,N_9416);
nand U11628 (N_11628,N_10379,N_10014);
nor U11629 (N_11629,N_10127,N_10025);
or U11630 (N_11630,N_9187,N_9338);
or U11631 (N_11631,N_10015,N_10126);
nor U11632 (N_11632,N_9196,N_9203);
xor U11633 (N_11633,N_10478,N_9935);
or U11634 (N_11634,N_9413,N_9981);
nand U11635 (N_11635,N_10252,N_9736);
nand U11636 (N_11636,N_10137,N_9985);
nand U11637 (N_11637,N_9337,N_9359);
or U11638 (N_11638,N_10111,N_9867);
nor U11639 (N_11639,N_9162,N_10427);
or U11640 (N_11640,N_10268,N_10301);
and U11641 (N_11641,N_9706,N_9648);
and U11642 (N_11642,N_9292,N_9970);
and U11643 (N_11643,N_9717,N_10150);
nor U11644 (N_11644,N_10475,N_9883);
nand U11645 (N_11645,N_9058,N_9036);
xor U11646 (N_11646,N_10265,N_9385);
nor U11647 (N_11647,N_9042,N_9773);
xnor U11648 (N_11648,N_9571,N_9134);
xnor U11649 (N_11649,N_9706,N_9120);
nor U11650 (N_11650,N_9538,N_10155);
and U11651 (N_11651,N_9516,N_9413);
nor U11652 (N_11652,N_10486,N_10483);
xnor U11653 (N_11653,N_10355,N_9285);
nand U11654 (N_11654,N_9551,N_9478);
nor U11655 (N_11655,N_9972,N_10213);
nand U11656 (N_11656,N_9813,N_9758);
xnor U11657 (N_11657,N_9973,N_9048);
xnor U11658 (N_11658,N_9744,N_10248);
nand U11659 (N_11659,N_9576,N_9880);
and U11660 (N_11660,N_9333,N_9840);
nand U11661 (N_11661,N_9560,N_9665);
or U11662 (N_11662,N_9449,N_9777);
xnor U11663 (N_11663,N_9702,N_10234);
or U11664 (N_11664,N_10258,N_9876);
and U11665 (N_11665,N_9193,N_9474);
xor U11666 (N_11666,N_9793,N_9321);
nor U11667 (N_11667,N_10332,N_9942);
or U11668 (N_11668,N_9435,N_9894);
xor U11669 (N_11669,N_9994,N_9065);
or U11670 (N_11670,N_9488,N_9301);
or U11671 (N_11671,N_9866,N_10080);
and U11672 (N_11672,N_10204,N_9012);
and U11673 (N_11673,N_9897,N_9724);
and U11674 (N_11674,N_9682,N_9725);
or U11675 (N_11675,N_9467,N_9672);
and U11676 (N_11676,N_9030,N_10013);
nor U11677 (N_11677,N_9272,N_9982);
nor U11678 (N_11678,N_9941,N_10444);
and U11679 (N_11679,N_9481,N_10117);
xor U11680 (N_11680,N_9459,N_10326);
or U11681 (N_11681,N_9299,N_9047);
and U11682 (N_11682,N_9436,N_10179);
xnor U11683 (N_11683,N_9834,N_10091);
nor U11684 (N_11684,N_9044,N_10385);
nand U11685 (N_11685,N_9282,N_9590);
nor U11686 (N_11686,N_9522,N_9763);
and U11687 (N_11687,N_9045,N_9844);
and U11688 (N_11688,N_9558,N_9965);
and U11689 (N_11689,N_9845,N_10388);
and U11690 (N_11690,N_9078,N_9839);
nand U11691 (N_11691,N_9448,N_9093);
nor U11692 (N_11692,N_9372,N_10102);
or U11693 (N_11693,N_10033,N_10083);
or U11694 (N_11694,N_9043,N_9369);
nor U11695 (N_11695,N_10442,N_10391);
nand U11696 (N_11696,N_9423,N_10086);
xnor U11697 (N_11697,N_9969,N_9179);
or U11698 (N_11698,N_9267,N_9742);
nand U11699 (N_11699,N_9025,N_9319);
or U11700 (N_11700,N_9102,N_9816);
nand U11701 (N_11701,N_9207,N_9895);
and U11702 (N_11702,N_9579,N_9677);
xnor U11703 (N_11703,N_9938,N_9534);
or U11704 (N_11704,N_9418,N_10446);
and U11705 (N_11705,N_9606,N_9787);
or U11706 (N_11706,N_9318,N_9844);
and U11707 (N_11707,N_9764,N_9726);
nor U11708 (N_11708,N_10038,N_9799);
or U11709 (N_11709,N_10474,N_10059);
xnor U11710 (N_11710,N_9185,N_10080);
and U11711 (N_11711,N_10335,N_9867);
nor U11712 (N_11712,N_9218,N_9090);
or U11713 (N_11713,N_10231,N_9683);
nor U11714 (N_11714,N_9212,N_9748);
xor U11715 (N_11715,N_9620,N_10357);
nand U11716 (N_11716,N_10395,N_9920);
and U11717 (N_11717,N_10379,N_9912);
xnor U11718 (N_11718,N_9880,N_9166);
nand U11719 (N_11719,N_9698,N_9492);
and U11720 (N_11720,N_9928,N_9677);
and U11721 (N_11721,N_10408,N_10433);
nor U11722 (N_11722,N_9873,N_9340);
nor U11723 (N_11723,N_9443,N_9326);
or U11724 (N_11724,N_9194,N_9636);
nand U11725 (N_11725,N_10411,N_10407);
nand U11726 (N_11726,N_9679,N_10039);
or U11727 (N_11727,N_9635,N_9137);
nor U11728 (N_11728,N_9813,N_10216);
or U11729 (N_11729,N_10126,N_9739);
xor U11730 (N_11730,N_9906,N_9791);
nor U11731 (N_11731,N_9970,N_9625);
or U11732 (N_11732,N_9295,N_9122);
and U11733 (N_11733,N_9197,N_10117);
and U11734 (N_11734,N_10238,N_10432);
nand U11735 (N_11735,N_9041,N_9986);
nor U11736 (N_11736,N_9004,N_9477);
nand U11737 (N_11737,N_10499,N_9852);
nand U11738 (N_11738,N_10399,N_10211);
and U11739 (N_11739,N_10064,N_9697);
or U11740 (N_11740,N_9867,N_10170);
or U11741 (N_11741,N_9534,N_9696);
xnor U11742 (N_11742,N_10096,N_10055);
and U11743 (N_11743,N_10206,N_10193);
xnor U11744 (N_11744,N_9499,N_9035);
xor U11745 (N_11745,N_10468,N_9306);
nand U11746 (N_11746,N_9398,N_9735);
nand U11747 (N_11747,N_10011,N_9585);
nand U11748 (N_11748,N_10330,N_9721);
or U11749 (N_11749,N_10180,N_9215);
nor U11750 (N_11750,N_9663,N_9846);
nand U11751 (N_11751,N_10119,N_9124);
or U11752 (N_11752,N_9776,N_10079);
nor U11753 (N_11753,N_10310,N_10145);
xor U11754 (N_11754,N_10265,N_9225);
nand U11755 (N_11755,N_9138,N_10072);
nand U11756 (N_11756,N_9849,N_9139);
nor U11757 (N_11757,N_10347,N_10191);
nor U11758 (N_11758,N_10264,N_10056);
and U11759 (N_11759,N_9290,N_10041);
or U11760 (N_11760,N_9985,N_9099);
nand U11761 (N_11761,N_9502,N_9488);
or U11762 (N_11762,N_9711,N_10183);
or U11763 (N_11763,N_10078,N_10447);
and U11764 (N_11764,N_9197,N_9456);
or U11765 (N_11765,N_9443,N_9327);
xor U11766 (N_11766,N_9040,N_10006);
xor U11767 (N_11767,N_10310,N_10247);
xor U11768 (N_11768,N_10058,N_10241);
nor U11769 (N_11769,N_10182,N_9925);
or U11770 (N_11770,N_9628,N_10460);
or U11771 (N_11771,N_9278,N_9257);
nor U11772 (N_11772,N_9781,N_10441);
nand U11773 (N_11773,N_9584,N_9161);
or U11774 (N_11774,N_9558,N_10147);
nor U11775 (N_11775,N_10078,N_9714);
and U11776 (N_11776,N_9331,N_10043);
nand U11777 (N_11777,N_9258,N_9781);
or U11778 (N_11778,N_9612,N_10178);
or U11779 (N_11779,N_9340,N_10265);
or U11780 (N_11780,N_9988,N_9964);
or U11781 (N_11781,N_9907,N_10405);
and U11782 (N_11782,N_9244,N_10472);
or U11783 (N_11783,N_9507,N_10023);
nor U11784 (N_11784,N_10055,N_9370);
nand U11785 (N_11785,N_10036,N_9046);
and U11786 (N_11786,N_9667,N_9574);
nor U11787 (N_11787,N_9697,N_10030);
and U11788 (N_11788,N_10233,N_10389);
nor U11789 (N_11789,N_9132,N_9463);
and U11790 (N_11790,N_9079,N_9972);
and U11791 (N_11791,N_9844,N_10151);
xnor U11792 (N_11792,N_9286,N_9675);
or U11793 (N_11793,N_10422,N_9503);
xor U11794 (N_11794,N_10144,N_9084);
and U11795 (N_11795,N_9314,N_10329);
or U11796 (N_11796,N_9745,N_9828);
xnor U11797 (N_11797,N_10117,N_9911);
or U11798 (N_11798,N_9383,N_10259);
nand U11799 (N_11799,N_9103,N_9244);
xnor U11800 (N_11800,N_9259,N_9012);
or U11801 (N_11801,N_9529,N_9139);
nor U11802 (N_11802,N_9337,N_9358);
nand U11803 (N_11803,N_9989,N_9266);
xnor U11804 (N_11804,N_10143,N_9590);
and U11805 (N_11805,N_9515,N_9014);
or U11806 (N_11806,N_10431,N_9448);
nor U11807 (N_11807,N_10263,N_10445);
and U11808 (N_11808,N_10358,N_9025);
xor U11809 (N_11809,N_10478,N_9197);
nor U11810 (N_11810,N_10007,N_10293);
and U11811 (N_11811,N_9731,N_9596);
and U11812 (N_11812,N_9934,N_10351);
nor U11813 (N_11813,N_9513,N_9295);
nand U11814 (N_11814,N_9940,N_10426);
and U11815 (N_11815,N_9772,N_9902);
nand U11816 (N_11816,N_10490,N_9505);
nor U11817 (N_11817,N_9414,N_9718);
nor U11818 (N_11818,N_9623,N_9920);
and U11819 (N_11819,N_10221,N_10462);
or U11820 (N_11820,N_9624,N_9529);
and U11821 (N_11821,N_9828,N_10120);
nand U11822 (N_11822,N_9294,N_9931);
xnor U11823 (N_11823,N_9265,N_9117);
nor U11824 (N_11824,N_10392,N_9877);
or U11825 (N_11825,N_9627,N_9377);
xor U11826 (N_11826,N_9506,N_9008);
nor U11827 (N_11827,N_9072,N_9182);
nor U11828 (N_11828,N_9305,N_9431);
and U11829 (N_11829,N_10404,N_10093);
nand U11830 (N_11830,N_10355,N_9328);
nand U11831 (N_11831,N_9249,N_9855);
nand U11832 (N_11832,N_9856,N_9460);
or U11833 (N_11833,N_10008,N_9934);
xor U11834 (N_11834,N_9886,N_10461);
nand U11835 (N_11835,N_9273,N_9517);
and U11836 (N_11836,N_9719,N_9181);
nor U11837 (N_11837,N_10130,N_10388);
nand U11838 (N_11838,N_9089,N_9771);
xor U11839 (N_11839,N_9339,N_9732);
nor U11840 (N_11840,N_10443,N_10137);
or U11841 (N_11841,N_9450,N_9646);
or U11842 (N_11842,N_9747,N_9068);
xnor U11843 (N_11843,N_9988,N_9154);
or U11844 (N_11844,N_9425,N_10144);
nand U11845 (N_11845,N_9421,N_9524);
nand U11846 (N_11846,N_10495,N_9491);
or U11847 (N_11847,N_9599,N_9643);
and U11848 (N_11848,N_9568,N_10043);
nand U11849 (N_11849,N_9855,N_9763);
or U11850 (N_11850,N_9069,N_10051);
nand U11851 (N_11851,N_10389,N_10226);
nand U11852 (N_11852,N_9344,N_10031);
and U11853 (N_11853,N_10470,N_9753);
xnor U11854 (N_11854,N_10193,N_9116);
or U11855 (N_11855,N_9480,N_9136);
xnor U11856 (N_11856,N_9697,N_9814);
nand U11857 (N_11857,N_9934,N_9823);
nand U11858 (N_11858,N_9669,N_9142);
nand U11859 (N_11859,N_9909,N_10458);
xnor U11860 (N_11860,N_10484,N_10319);
xor U11861 (N_11861,N_9160,N_9611);
or U11862 (N_11862,N_9804,N_9131);
nand U11863 (N_11863,N_9010,N_9432);
nand U11864 (N_11864,N_9675,N_10166);
xnor U11865 (N_11865,N_9128,N_9056);
xor U11866 (N_11866,N_9728,N_10495);
and U11867 (N_11867,N_9115,N_10427);
or U11868 (N_11868,N_10317,N_9096);
nor U11869 (N_11869,N_9907,N_9130);
xnor U11870 (N_11870,N_9647,N_9694);
xor U11871 (N_11871,N_9694,N_9038);
nor U11872 (N_11872,N_9356,N_9227);
or U11873 (N_11873,N_9581,N_10147);
nor U11874 (N_11874,N_10280,N_9418);
and U11875 (N_11875,N_10367,N_9215);
nand U11876 (N_11876,N_9852,N_9535);
xor U11877 (N_11877,N_10464,N_9234);
xnor U11878 (N_11878,N_9319,N_10285);
nor U11879 (N_11879,N_9875,N_10016);
xor U11880 (N_11880,N_9531,N_10371);
and U11881 (N_11881,N_9070,N_9066);
and U11882 (N_11882,N_10430,N_9282);
and U11883 (N_11883,N_9557,N_10362);
and U11884 (N_11884,N_9602,N_9884);
and U11885 (N_11885,N_9652,N_9222);
or U11886 (N_11886,N_10060,N_9726);
and U11887 (N_11887,N_9295,N_10396);
nor U11888 (N_11888,N_9636,N_10379);
nor U11889 (N_11889,N_10006,N_10249);
nor U11890 (N_11890,N_10238,N_9433);
xor U11891 (N_11891,N_9251,N_10477);
nor U11892 (N_11892,N_9019,N_9289);
xnor U11893 (N_11893,N_9995,N_9930);
and U11894 (N_11894,N_10353,N_9947);
or U11895 (N_11895,N_10343,N_10482);
nor U11896 (N_11896,N_9645,N_9252);
xor U11897 (N_11897,N_9313,N_9042);
and U11898 (N_11898,N_9908,N_10495);
and U11899 (N_11899,N_9915,N_9184);
xor U11900 (N_11900,N_10139,N_9823);
nor U11901 (N_11901,N_9141,N_9126);
and U11902 (N_11902,N_10226,N_9097);
nand U11903 (N_11903,N_10299,N_9359);
xnor U11904 (N_11904,N_9894,N_10001);
nor U11905 (N_11905,N_9477,N_10080);
xnor U11906 (N_11906,N_9901,N_9924);
nor U11907 (N_11907,N_9879,N_9887);
nor U11908 (N_11908,N_10111,N_9171);
nand U11909 (N_11909,N_9264,N_9100);
and U11910 (N_11910,N_9039,N_9488);
xor U11911 (N_11911,N_10036,N_9621);
nor U11912 (N_11912,N_10182,N_9050);
and U11913 (N_11913,N_9496,N_9143);
xor U11914 (N_11914,N_9203,N_10476);
nor U11915 (N_11915,N_9936,N_9210);
nor U11916 (N_11916,N_10115,N_10181);
nor U11917 (N_11917,N_9382,N_9408);
nand U11918 (N_11918,N_9400,N_10135);
nand U11919 (N_11919,N_9456,N_9383);
or U11920 (N_11920,N_10182,N_10263);
xnor U11921 (N_11921,N_9526,N_10496);
or U11922 (N_11922,N_10001,N_10122);
nor U11923 (N_11923,N_10004,N_9371);
nor U11924 (N_11924,N_9026,N_9926);
or U11925 (N_11925,N_9975,N_9233);
xnor U11926 (N_11926,N_9214,N_10283);
nor U11927 (N_11927,N_10204,N_10473);
nor U11928 (N_11928,N_9744,N_9793);
or U11929 (N_11929,N_9031,N_9854);
nor U11930 (N_11930,N_9258,N_10089);
and U11931 (N_11931,N_9558,N_9734);
nor U11932 (N_11932,N_9480,N_9552);
xnor U11933 (N_11933,N_10453,N_9166);
nor U11934 (N_11934,N_10306,N_9969);
and U11935 (N_11935,N_10109,N_9309);
or U11936 (N_11936,N_9257,N_10005);
or U11937 (N_11937,N_9596,N_9572);
and U11938 (N_11938,N_9050,N_10211);
nand U11939 (N_11939,N_9015,N_9559);
xor U11940 (N_11940,N_9905,N_9668);
nand U11941 (N_11941,N_10163,N_9661);
nor U11942 (N_11942,N_9349,N_9557);
nor U11943 (N_11943,N_10491,N_10493);
and U11944 (N_11944,N_9682,N_9728);
and U11945 (N_11945,N_9869,N_10286);
and U11946 (N_11946,N_9257,N_10080);
nor U11947 (N_11947,N_10007,N_9851);
or U11948 (N_11948,N_9286,N_9471);
xnor U11949 (N_11949,N_9371,N_9654);
and U11950 (N_11950,N_10123,N_10412);
nand U11951 (N_11951,N_9950,N_10439);
nand U11952 (N_11952,N_9715,N_10404);
and U11953 (N_11953,N_9230,N_10499);
nand U11954 (N_11954,N_10227,N_10173);
xor U11955 (N_11955,N_9935,N_10465);
and U11956 (N_11956,N_10249,N_10347);
nand U11957 (N_11957,N_9234,N_9718);
or U11958 (N_11958,N_9813,N_9806);
and U11959 (N_11959,N_9046,N_9515);
nor U11960 (N_11960,N_9002,N_9380);
nor U11961 (N_11961,N_9032,N_9975);
or U11962 (N_11962,N_10496,N_9989);
xor U11963 (N_11963,N_9182,N_10062);
nand U11964 (N_11964,N_10445,N_9101);
or U11965 (N_11965,N_9748,N_9722);
xnor U11966 (N_11966,N_10229,N_9733);
xor U11967 (N_11967,N_9315,N_9988);
or U11968 (N_11968,N_10337,N_9481);
nand U11969 (N_11969,N_9531,N_9892);
nor U11970 (N_11970,N_9215,N_9879);
and U11971 (N_11971,N_9898,N_9137);
or U11972 (N_11972,N_10116,N_10149);
or U11973 (N_11973,N_10227,N_9801);
or U11974 (N_11974,N_9262,N_9015);
nand U11975 (N_11975,N_9228,N_9625);
or U11976 (N_11976,N_9462,N_9842);
nor U11977 (N_11977,N_9838,N_9835);
or U11978 (N_11978,N_9534,N_10082);
and U11979 (N_11979,N_9027,N_10327);
nand U11980 (N_11980,N_9921,N_9552);
nand U11981 (N_11981,N_9713,N_10114);
nand U11982 (N_11982,N_9275,N_10096);
xnor U11983 (N_11983,N_9266,N_10402);
and U11984 (N_11984,N_10298,N_9924);
nand U11985 (N_11985,N_10226,N_9570);
and U11986 (N_11986,N_9864,N_10050);
nand U11987 (N_11987,N_10012,N_9236);
nor U11988 (N_11988,N_9581,N_10363);
nor U11989 (N_11989,N_9968,N_9287);
xor U11990 (N_11990,N_10146,N_10447);
and U11991 (N_11991,N_9862,N_9165);
nor U11992 (N_11992,N_10477,N_9703);
nand U11993 (N_11993,N_9129,N_9138);
nand U11994 (N_11994,N_10170,N_10113);
nand U11995 (N_11995,N_10299,N_9142);
nor U11996 (N_11996,N_9895,N_9905);
xor U11997 (N_11997,N_10277,N_9543);
xnor U11998 (N_11998,N_9254,N_10390);
nor U11999 (N_11999,N_10433,N_10026);
or U12000 (N_12000,N_10953,N_11478);
xor U12001 (N_12001,N_11440,N_11551);
nand U12002 (N_12002,N_11616,N_10686);
or U12003 (N_12003,N_11162,N_11891);
or U12004 (N_12004,N_10558,N_11837);
xnor U12005 (N_12005,N_11627,N_11861);
nand U12006 (N_12006,N_10844,N_11914);
nor U12007 (N_12007,N_10882,N_11302);
nor U12008 (N_12008,N_11421,N_11495);
and U12009 (N_12009,N_11393,N_11946);
or U12010 (N_12010,N_11783,N_11282);
xor U12011 (N_12011,N_11986,N_11945);
or U12012 (N_12012,N_11787,N_11492);
xor U12013 (N_12013,N_10752,N_10502);
and U12014 (N_12014,N_11933,N_11909);
nand U12015 (N_12015,N_11655,N_10889);
xnor U12016 (N_12016,N_10636,N_11696);
nor U12017 (N_12017,N_11605,N_10571);
and U12018 (N_12018,N_11143,N_11506);
xor U12019 (N_12019,N_10907,N_10512);
xor U12020 (N_12020,N_10591,N_11033);
or U12021 (N_12021,N_10744,N_11342);
or U12022 (N_12022,N_11180,N_11124);
xor U12023 (N_12023,N_11754,N_11164);
xor U12024 (N_12024,N_10992,N_10981);
xor U12025 (N_12025,N_10829,N_11738);
xor U12026 (N_12026,N_10964,N_11568);
nand U12027 (N_12027,N_11536,N_10707);
xnor U12028 (N_12028,N_11064,N_10709);
xor U12029 (N_12029,N_11157,N_10818);
and U12030 (N_12030,N_11392,N_11087);
nor U12031 (N_12031,N_10903,N_11792);
nor U12032 (N_12032,N_11223,N_11182);
or U12033 (N_12033,N_11177,N_10904);
and U12034 (N_12034,N_11541,N_11363);
xnor U12035 (N_12035,N_11802,N_10792);
and U12036 (N_12036,N_11053,N_11035);
nor U12037 (N_12037,N_11594,N_10837);
nor U12038 (N_12038,N_10627,N_11472);
nor U12039 (N_12039,N_11467,N_11831);
or U12040 (N_12040,N_11714,N_10513);
or U12041 (N_12041,N_11537,N_11431);
nand U12042 (N_12042,N_10532,N_10740);
nor U12043 (N_12043,N_11334,N_11899);
xnor U12044 (N_12044,N_11731,N_11242);
and U12045 (N_12045,N_11309,N_10618);
or U12046 (N_12046,N_10834,N_11084);
or U12047 (N_12047,N_11694,N_10958);
nor U12048 (N_12048,N_11343,N_11148);
or U12049 (N_12049,N_11960,N_11181);
or U12050 (N_12050,N_10548,N_10746);
nor U12051 (N_12051,N_11331,N_11746);
or U12052 (N_12052,N_11367,N_11189);
nor U12053 (N_12053,N_11310,N_10683);
xnor U12054 (N_12054,N_10613,N_11489);
nand U12055 (N_12055,N_11679,N_10612);
nand U12056 (N_12056,N_11398,N_11370);
nand U12057 (N_12057,N_11298,N_10971);
or U12058 (N_12058,N_11482,N_11847);
nor U12059 (N_12059,N_10664,N_11790);
xnor U12060 (N_12060,N_11739,N_11815);
and U12061 (N_12061,N_10638,N_10701);
or U12062 (N_12062,N_11453,N_11761);
nor U12063 (N_12063,N_11598,N_10867);
nand U12064 (N_12064,N_10935,N_10514);
xor U12065 (N_12065,N_10576,N_11144);
xnor U12066 (N_12066,N_10741,N_10602);
and U12067 (N_12067,N_11606,N_11689);
nand U12068 (N_12068,N_11906,N_11400);
xnor U12069 (N_12069,N_11000,N_10812);
nand U12070 (N_12070,N_11968,N_11828);
or U12071 (N_12071,N_11789,N_10911);
xnor U12072 (N_12072,N_11785,N_11722);
xnor U12073 (N_12073,N_11580,N_11257);
xnor U12074 (N_12074,N_11179,N_11592);
or U12075 (N_12075,N_10601,N_11254);
nand U12076 (N_12076,N_11108,N_11522);
nor U12077 (N_12077,N_11122,N_11697);
nor U12078 (N_12078,N_11003,N_11997);
nand U12079 (N_12079,N_11077,N_10519);
or U12080 (N_12080,N_11947,N_10585);
xor U12081 (N_12081,N_11207,N_11813);
nor U12082 (N_12082,N_10861,N_10830);
or U12083 (N_12083,N_11127,N_11500);
xnor U12084 (N_12084,N_11823,N_10542);
nor U12085 (N_12085,N_11676,N_10962);
nand U12086 (N_12086,N_11626,N_11280);
xor U12087 (N_12087,N_10939,N_11666);
xor U12088 (N_12088,N_10906,N_11865);
xnor U12089 (N_12089,N_11415,N_11459);
xnor U12090 (N_12090,N_10766,N_11653);
nor U12091 (N_12091,N_10743,N_11633);
xor U12092 (N_12092,N_11566,N_10771);
or U12093 (N_12093,N_11644,N_10778);
and U12094 (N_12094,N_11229,N_11981);
or U12095 (N_12095,N_11481,N_11951);
nand U12096 (N_12096,N_10891,N_10530);
xnor U12097 (N_12097,N_10719,N_10804);
and U12098 (N_12098,N_11337,N_11272);
nor U12099 (N_12099,N_11215,N_11235);
or U12100 (N_12100,N_11455,N_11405);
or U12101 (N_12101,N_10692,N_11126);
nor U12102 (N_12102,N_10643,N_10648);
nor U12103 (N_12103,N_10808,N_10950);
nand U12104 (N_12104,N_10751,N_10641);
and U12105 (N_12105,N_10634,N_11677);
nor U12106 (N_12106,N_11692,N_10913);
xor U12107 (N_12107,N_11137,N_11401);
or U12108 (N_12108,N_11059,N_10553);
xor U12109 (N_12109,N_11186,N_10736);
nor U12110 (N_12110,N_11289,N_11065);
xor U12111 (N_12111,N_10816,N_11602);
or U12112 (N_12112,N_11420,N_10619);
or U12113 (N_12113,N_11493,N_11161);
and U12114 (N_12114,N_11438,N_11718);
xnor U12115 (N_12115,N_11917,N_10592);
nor U12116 (N_12116,N_11197,N_11276);
and U12117 (N_12117,N_11388,N_11973);
and U12118 (N_12118,N_11526,N_11674);
or U12119 (N_12119,N_11665,N_11972);
nor U12120 (N_12120,N_11520,N_10948);
or U12121 (N_12121,N_11700,N_10956);
and U12122 (N_12122,N_11525,N_11563);
and U12123 (N_12123,N_10959,N_11678);
or U12124 (N_12124,N_11199,N_10520);
or U12125 (N_12125,N_10857,N_10811);
nor U12126 (N_12126,N_11114,N_11572);
nand U12127 (N_12127,N_10824,N_10713);
nand U12128 (N_12128,N_11394,N_10960);
and U12129 (N_12129,N_10989,N_10782);
xor U12130 (N_12130,N_11673,N_10842);
and U12131 (N_12131,N_11275,N_10783);
xor U12132 (N_12132,N_11066,N_11086);
or U12133 (N_12133,N_10846,N_11695);
nor U12134 (N_12134,N_11043,N_11376);
and U12135 (N_12135,N_11936,N_11095);
or U12136 (N_12136,N_10767,N_10657);
or U12137 (N_12137,N_11646,N_11573);
nand U12138 (N_12138,N_11436,N_11717);
nor U12139 (N_12139,N_11292,N_10995);
nor U12140 (N_12140,N_11886,N_10915);
xor U12141 (N_12141,N_10908,N_11527);
and U12142 (N_12142,N_10863,N_11117);
xor U12143 (N_12143,N_10787,N_10756);
xnor U12144 (N_12144,N_11976,N_11921);
xor U12145 (N_12145,N_11191,N_10968);
and U12146 (N_12146,N_10931,N_11332);
or U12147 (N_12147,N_11120,N_11397);
and U12148 (N_12148,N_11217,N_11227);
and U12149 (N_12149,N_10801,N_10796);
xor U12150 (N_12150,N_11470,N_11390);
or U12151 (N_12151,N_11950,N_11725);
and U12152 (N_12152,N_11608,N_10626);
or U12153 (N_12153,N_11011,N_11067);
nor U12154 (N_12154,N_10825,N_11957);
xnor U12155 (N_12155,N_11051,N_10758);
or U12156 (N_12156,N_11039,N_11726);
nand U12157 (N_12157,N_10506,N_11962);
and U12158 (N_12158,N_10933,N_11629);
or U12159 (N_12159,N_10587,N_11359);
xnor U12160 (N_12160,N_10644,N_11709);
xor U12161 (N_12161,N_11680,N_11021);
nand U12162 (N_12162,N_11918,N_11544);
nor U12163 (N_12163,N_11928,N_11028);
or U12164 (N_12164,N_11875,N_10533);
nor U12165 (N_12165,N_11872,N_10902);
and U12166 (N_12166,N_11371,N_11924);
and U12167 (N_12167,N_10625,N_11859);
and U12168 (N_12168,N_11328,N_11412);
or U12169 (N_12169,N_10930,N_11588);
xor U12170 (N_12170,N_11348,N_10504);
xor U12171 (N_12171,N_11958,N_10870);
xnor U12172 (N_12172,N_10859,N_10828);
or U12173 (N_12173,N_10578,N_11850);
xor U12174 (N_12174,N_11346,N_11032);
xor U12175 (N_12175,N_11821,N_11931);
nand U12176 (N_12176,N_11411,N_11360);
xnor U12177 (N_12177,N_11867,N_10848);
nand U12178 (N_12178,N_11615,N_11675);
or U12179 (N_12179,N_11545,N_10656);
xor U12180 (N_12180,N_10773,N_11024);
and U12181 (N_12181,N_10645,N_10862);
nand U12182 (N_12182,N_11693,N_11351);
xor U12183 (N_12183,N_11168,N_10755);
or U12184 (N_12184,N_11839,N_10975);
or U12185 (N_12185,N_11613,N_11905);
or U12186 (N_12186,N_11897,N_11538);
or U12187 (N_12187,N_11132,N_10674);
nand U12188 (N_12188,N_10528,N_11940);
xnor U12189 (N_12189,N_10681,N_11840);
xor U12190 (N_12190,N_11660,N_11515);
nor U12191 (N_12191,N_11702,N_10984);
xnor U12192 (N_12192,N_11251,N_10869);
nand U12193 (N_12193,N_11979,N_11093);
or U12194 (N_12194,N_11050,N_10689);
xnor U12195 (N_12195,N_10919,N_11820);
nor U12196 (N_12196,N_10819,N_10775);
or U12197 (N_12197,N_11012,N_11582);
xor U12198 (N_12198,N_11650,N_11510);
nor U12199 (N_12199,N_11112,N_10853);
nand U12200 (N_12200,N_10742,N_10724);
or U12201 (N_12201,N_11423,N_11829);
and U12202 (N_12202,N_10652,N_11686);
nor U12203 (N_12203,N_11433,N_11099);
nand U12204 (N_12204,N_10607,N_11892);
xnor U12205 (N_12205,N_11183,N_11002);
nor U12206 (N_12206,N_11599,N_11381);
and U12207 (N_12207,N_10753,N_10604);
or U12208 (N_12208,N_10716,N_10665);
and U12209 (N_12209,N_10759,N_11955);
xnor U12210 (N_12210,N_11110,N_11497);
xor U12211 (N_12211,N_11920,N_11980);
and U12212 (N_12212,N_11073,N_11068);
and U12213 (N_12213,N_11333,N_11504);
and U12214 (N_12214,N_10895,N_11218);
xor U12215 (N_12215,N_11378,N_11637);
xor U12216 (N_12216,N_11652,N_10865);
nor U12217 (N_12217,N_11836,N_11311);
and U12218 (N_12218,N_10518,N_10609);
nor U12219 (N_12219,N_11712,N_10888);
and U12220 (N_12220,N_11911,N_10874);
nor U12221 (N_12221,N_11904,N_11741);
xor U12222 (N_12222,N_11873,N_11454);
xnor U12223 (N_12223,N_11221,N_11935);
and U12224 (N_12224,N_11442,N_11387);
xnor U12225 (N_12225,N_11006,N_11667);
nand U12226 (N_12226,N_11427,N_10810);
nand U12227 (N_12227,N_10581,N_11779);
xor U12228 (N_12228,N_11877,N_11888);
nand U12229 (N_12229,N_11944,N_11408);
nor U12230 (N_12230,N_10509,N_10708);
nor U12231 (N_12231,N_11794,N_10599);
nor U12232 (N_12232,N_11540,N_11170);
nand U12233 (N_12233,N_10552,N_11611);
or U12234 (N_12234,N_11410,N_11552);
xor U12235 (N_12235,N_11358,N_11542);
xor U12236 (N_12236,N_11042,N_11446);
or U12237 (N_12237,N_11547,N_11303);
and U12238 (N_12238,N_11476,N_11341);
nand U12239 (N_12239,N_10997,N_11038);
nor U12240 (N_12240,N_11304,N_11305);
and U12241 (N_12241,N_11462,N_11034);
and U12242 (N_12242,N_10507,N_11817);
and U12243 (N_12243,N_10925,N_11879);
xor U12244 (N_12244,N_11954,N_10815);
nor U12245 (N_12245,N_11621,N_11317);
xor U12246 (N_12246,N_10963,N_11092);
xnor U12247 (N_12247,N_11096,N_11742);
nor U12248 (N_12248,N_11187,N_11245);
and U12249 (N_12249,N_11017,N_10832);
or U12250 (N_12250,N_11880,N_11138);
and U12251 (N_12251,N_11659,N_11581);
nor U12252 (N_12252,N_10957,N_11314);
xnor U12253 (N_12253,N_11457,N_10823);
xor U12254 (N_12254,N_11558,N_10589);
and U12255 (N_12255,N_11784,N_11239);
and U12256 (N_12256,N_11844,N_11636);
nand U12257 (N_12257,N_11283,N_11031);
nor U12258 (N_12258,N_11361,N_11721);
nand U12259 (N_12259,N_11372,N_11374);
nand U12260 (N_12260,N_11174,N_10880);
or U12261 (N_12261,N_11103,N_10640);
or U12262 (N_12262,N_11151,N_10871);
and U12263 (N_12263,N_11971,N_10614);
nor U12264 (N_12264,N_11009,N_11001);
nand U12265 (N_12265,N_11238,N_10590);
nor U12266 (N_12266,N_10556,N_11444);
nand U12267 (N_12267,N_10761,N_11163);
and U12268 (N_12268,N_10800,N_11728);
or U12269 (N_12269,N_11424,N_10790);
xnor U12270 (N_12270,N_11115,N_10769);
nor U12271 (N_12271,N_11969,N_10910);
xnor U12272 (N_12272,N_11733,N_10595);
nor U12273 (N_12273,N_10517,N_10788);
or U12274 (N_12274,N_11713,N_11641);
xnor U12275 (N_12275,N_11403,N_11715);
xor U12276 (N_12276,N_11209,N_11494);
xor U12277 (N_12277,N_10723,N_11811);
nand U12278 (N_12278,N_11777,N_10588);
nor U12279 (N_12279,N_11325,N_10580);
and U12280 (N_12280,N_11070,N_10500);
nor U12281 (N_12281,N_10765,N_11796);
nand U12282 (N_12282,N_10879,N_11628);
nor U12283 (N_12283,N_11135,N_10917);
or U12284 (N_12284,N_10924,N_11827);
xnor U12285 (N_12285,N_11255,N_10999);
nor U12286 (N_12286,N_11736,N_11805);
nand U12287 (N_12287,N_10986,N_11727);
nand U12288 (N_12288,N_11452,N_10623);
nand U12289 (N_12289,N_10985,N_10762);
xnor U12290 (N_12290,N_10515,N_11324);
nor U12291 (N_12291,N_11630,N_11595);
xor U12292 (N_12292,N_11664,N_11952);
nand U12293 (N_12293,N_11752,N_11123);
nor U12294 (N_12294,N_11903,N_11668);
or U12295 (N_12295,N_11262,N_11434);
nand U12296 (N_12296,N_10797,N_11845);
nor U12297 (N_12297,N_10941,N_10596);
xor U12298 (N_12298,N_11425,N_11826);
or U12299 (N_12299,N_11090,N_10951);
and U12300 (N_12300,N_10661,N_11767);
xnor U12301 (N_12301,N_11804,N_11720);
and U12302 (N_12302,N_10539,N_10566);
or U12303 (N_12303,N_11048,N_10653);
nor U12304 (N_12304,N_11856,N_11670);
and U12305 (N_12305,N_11364,N_11091);
and U12306 (N_12306,N_11149,N_10983);
nand U12307 (N_12307,N_11716,N_11188);
nand U12308 (N_12308,N_11825,N_11499);
xnor U12309 (N_12309,N_11406,N_11601);
xor U12310 (N_12310,N_11756,N_11194);
or U12311 (N_12311,N_10991,N_10593);
nand U12312 (N_12312,N_10568,N_11838);
and U12313 (N_12313,N_11740,N_11270);
or U12314 (N_12314,N_10702,N_10600);
or U12315 (N_12315,N_11535,N_11576);
nor U12316 (N_12316,N_11147,N_11878);
nand U12317 (N_12317,N_10894,N_11672);
xnor U12318 (N_12318,N_10858,N_11391);
nand U12319 (N_12319,N_10923,N_10864);
xnor U12320 (N_12320,N_10563,N_11432);
or U12321 (N_12321,N_11205,N_11172);
and U12322 (N_12322,N_11632,N_11548);
xor U12323 (N_12323,N_11232,N_11249);
and U12324 (N_12324,N_11154,N_11498);
nor U12325 (N_12325,N_11208,N_11041);
and U12326 (N_12326,N_10734,N_10791);
and U12327 (N_12327,N_11669,N_10901);
nor U12328 (N_12328,N_11516,N_11071);
nand U12329 (N_12329,N_11587,N_11513);
nand U12330 (N_12330,N_11926,N_11220);
and U12331 (N_12331,N_11801,N_10764);
and U12332 (N_12332,N_11369,N_11037);
nor U12333 (N_12333,N_10955,N_10586);
nor U12334 (N_12334,N_10892,N_11529);
nand U12335 (N_12335,N_10916,N_11166);
and U12336 (N_12336,N_11835,N_10521);
or U12337 (N_12337,N_10667,N_11266);
nor U12338 (N_12338,N_11966,N_11167);
or U12339 (N_12339,N_11943,N_11244);
nor U12340 (N_12340,N_11141,N_11556);
and U12341 (N_12341,N_11810,N_11977);
nor U12342 (N_12342,N_11338,N_10727);
nor U12343 (N_12343,N_11795,N_11743);
nand U12344 (N_12344,N_10573,N_11340);
and U12345 (N_12345,N_11019,N_11623);
or U12346 (N_12346,N_10620,N_11569);
or U12347 (N_12347,N_11539,N_10711);
or U12348 (N_12348,N_10575,N_11922);
nand U12349 (N_12349,N_10905,N_11876);
xor U12350 (N_12350,N_11448,N_11014);
nor U12351 (N_12351,N_11948,N_10726);
and U12352 (N_12352,N_10881,N_11225);
nand U12353 (N_12353,N_11080,N_10898);
or U12354 (N_12354,N_10884,N_11354);
or U12355 (N_12355,N_11414,N_10763);
nor U12356 (N_12356,N_10546,N_11648);
nand U12357 (N_12357,N_11322,N_11708);
and U12358 (N_12358,N_11047,N_11871);
xor U12359 (N_12359,N_10505,N_11748);
nand U12360 (N_12360,N_11890,N_11176);
nand U12361 (N_12361,N_11040,N_11816);
nor U12362 (N_12362,N_10560,N_11134);
nor U12363 (N_12363,N_10739,N_11895);
nor U12364 (N_12364,N_11158,N_11550);
or U12365 (N_12365,N_11557,N_11119);
or U12366 (N_12366,N_10803,N_11543);
and U12367 (N_12367,N_11060,N_11368);
xor U12368 (N_12368,N_10845,N_10749);
nand U12369 (N_12369,N_11316,N_10703);
and U12370 (N_12370,N_10817,N_11081);
nand U12371 (N_12371,N_10990,N_11638);
nand U12372 (N_12372,N_11130,N_11076);
and U12373 (N_12373,N_11356,N_10650);
nor U12374 (N_12374,N_10946,N_10760);
xor U12375 (N_12375,N_11734,N_11773);
nor U12376 (N_12376,N_11583,N_10809);
and U12377 (N_12377,N_11849,N_10524);
and U12378 (N_12378,N_10608,N_10712);
nor U12379 (N_12379,N_11999,N_11780);
nand U12380 (N_12380,N_11990,N_11584);
nand U12381 (N_12381,N_11927,N_11910);
nand U12382 (N_12382,N_11604,N_11111);
or U12383 (N_12383,N_11213,N_11932);
xnor U12384 (N_12384,N_11320,N_11479);
nand U12385 (N_12385,N_11056,N_11524);
nand U12386 (N_12386,N_11681,N_11706);
and U12387 (N_12387,N_11030,N_11285);
xnor U12388 (N_12388,N_11770,N_11514);
nor U12389 (N_12389,N_11247,N_11993);
xor U12390 (N_12390,N_11671,N_10691);
nand U12391 (N_12391,N_11508,N_11246);
and U12392 (N_12392,N_11812,N_10526);
xor U12393 (N_12393,N_10993,N_11750);
xnor U12394 (N_12394,N_11206,N_11078);
xnor U12395 (N_12395,N_11869,N_10972);
xor U12396 (N_12396,N_11121,N_10969);
xnor U12397 (N_12397,N_10511,N_11152);
and U12398 (N_12398,N_10660,N_11384);
and U12399 (N_12399,N_10970,N_11488);
and U12400 (N_12400,N_11842,N_10840);
nand U12401 (N_12401,N_11778,N_10615);
nand U12402 (N_12402,N_11422,N_11362);
or U12403 (N_12403,N_11234,N_11153);
or U12404 (N_12404,N_10738,N_10503);
nand U12405 (N_12405,N_10714,N_11685);
and U12406 (N_12406,N_11062,N_11916);
nor U12407 (N_12407,N_11214,N_11509);
and U12408 (N_12408,N_11710,N_10883);
xor U12409 (N_12409,N_10843,N_11465);
nor U12410 (N_12410,N_11760,N_11564);
nand U12411 (N_12411,N_11241,N_11466);
nand U12412 (N_12412,N_10662,N_10821);
xnor U12413 (N_12413,N_11451,N_11596);
nor U12414 (N_12414,N_11203,N_11279);
and U12415 (N_12415,N_11737,N_10680);
or U12416 (N_12416,N_11730,N_11998);
nor U12417 (N_12417,N_10543,N_11365);
xor U12418 (N_12418,N_11061,N_11991);
and U12419 (N_12419,N_11758,N_11724);
and U12420 (N_12420,N_10710,N_11445);
nor U12421 (N_12421,N_11683,N_11355);
or U12422 (N_12422,N_11768,N_11243);
xor U12423 (N_12423,N_10729,N_10860);
and U12424 (N_12424,N_11159,N_10733);
or U12425 (N_12425,N_11854,N_11894);
and U12426 (N_12426,N_10732,N_11271);
xnor U12427 (N_12427,N_11069,N_10777);
or U12428 (N_12428,N_11774,N_11864);
nand U12429 (N_12429,N_11301,N_11639);
and U12430 (N_12430,N_11487,N_10577);
and U12431 (N_12431,N_11491,N_10831);
nand U12432 (N_12432,N_11389,N_10754);
and U12433 (N_12433,N_11079,N_10676);
and U12434 (N_12434,N_11647,N_10875);
and U12435 (N_12435,N_10582,N_11399);
nand U12436 (N_12436,N_11575,N_11049);
nand U12437 (N_12437,N_11377,N_11306);
or U12438 (N_12438,N_11469,N_10555);
and U12439 (N_12439,N_11763,N_11128);
nand U12440 (N_12440,N_10748,N_11978);
nand U12441 (N_12441,N_11764,N_11866);
and U12442 (N_12442,N_11352,N_11942);
xor U12443 (N_12443,N_11819,N_10536);
nand U12444 (N_12444,N_11413,N_11256);
nor U12445 (N_12445,N_11657,N_11753);
nand U12446 (N_12446,N_10541,N_11766);
nor U12447 (N_12447,N_10569,N_10899);
nand U12448 (N_12448,N_10926,N_10594);
xor U12449 (N_12449,N_10929,N_11586);
and U12450 (N_12450,N_11312,N_11101);
xor U12451 (N_12451,N_11008,N_11449);
and U12452 (N_12452,N_11222,N_11959);
nand U12453 (N_12453,N_10605,N_10693);
and U12454 (N_12454,N_11326,N_11344);
xnor U12455 (N_12455,N_11719,N_10942);
or U12456 (N_12456,N_10918,N_11435);
xor U12457 (N_12457,N_10943,N_10730);
xor U12458 (N_12458,N_11983,N_11624);
or U12459 (N_12459,N_11426,N_10531);
or U12460 (N_12460,N_11938,N_10833);
or U12461 (N_12461,N_11461,N_11382);
nand U12462 (N_12462,N_10720,N_11691);
or U12463 (N_12463,N_11456,N_10670);
and U12464 (N_12464,N_10651,N_11441);
nand U12465 (N_12465,N_11089,N_11882);
or U12466 (N_12466,N_10666,N_11661);
nor U12467 (N_12467,N_11518,N_10647);
and U12468 (N_12468,N_11236,N_11202);
nand U12469 (N_12469,N_11631,N_11104);
and U12470 (N_12470,N_11887,N_11313);
xor U12471 (N_12471,N_10570,N_10706);
xnor U12472 (N_12472,N_10885,N_10976);
and U12473 (N_12473,N_11765,N_11025);
and U12474 (N_12474,N_10822,N_10633);
nand U12475 (N_12475,N_11807,N_11085);
and U12476 (N_12476,N_11267,N_10798);
nor U12477 (N_12477,N_11546,N_11105);
xor U12478 (N_12478,N_11902,N_11614);
nor U12479 (N_12479,N_11142,N_11704);
or U12480 (N_12480,N_11567,N_11329);
xnor U12481 (N_12481,N_11925,N_11965);
nand U12482 (N_12482,N_11803,N_10565);
or U12483 (N_12483,N_10937,N_10735);
and U12484 (N_12484,N_11443,N_10852);
or U12485 (N_12485,N_10649,N_11125);
xor U12486 (N_12486,N_11184,N_10938);
xor U12487 (N_12487,N_11204,N_11800);
xor U12488 (N_12488,N_11230,N_11484);
xor U12489 (N_12489,N_11964,N_11759);
nor U12490 (N_12490,N_10772,N_11437);
nor U12491 (N_12491,N_10934,N_11511);
and U12492 (N_12492,N_11862,N_11559);
nor U12493 (N_12493,N_11597,N_10658);
or U12494 (N_12494,N_10725,N_11318);
or U12495 (N_12495,N_10722,N_11045);
nand U12496 (N_12496,N_11195,N_10682);
nand U12497 (N_12497,N_11155,N_10947);
or U12498 (N_12498,N_11345,N_11027);
nand U12499 (N_12499,N_11074,N_11949);
nand U12500 (N_12500,N_11475,N_11610);
nand U12501 (N_12501,N_11129,N_11417);
xnor U12502 (N_12502,N_11769,N_10685);
and U12503 (N_12503,N_10688,N_10806);
nand U12504 (N_12504,N_11323,N_11395);
nand U12505 (N_12505,N_11622,N_11521);
xnor U12506 (N_12506,N_11463,N_11335);
xor U12507 (N_12507,N_11591,N_11269);
nor U12508 (N_12508,N_10642,N_10814);
nor U12509 (N_12509,N_11160,N_11200);
xor U12510 (N_12510,N_10704,N_11956);
or U12511 (N_12511,N_10731,N_11707);
xor U12512 (N_12512,N_11350,N_10522);
xnor U12513 (N_12513,N_11502,N_10617);
and U12514 (N_12514,N_11822,N_11620);
and U12515 (N_12515,N_11458,N_10501);
or U12516 (N_12516,N_11744,N_11923);
or U12517 (N_12517,N_10785,N_11635);
or U12518 (N_12518,N_10768,N_11786);
and U12519 (N_12519,N_11732,N_11989);
or U12520 (N_12520,N_11347,N_11645);
xnor U12521 (N_12521,N_10551,N_11201);
nand U12522 (N_12522,N_10598,N_11775);
or U12523 (N_12523,N_10554,N_10646);
or U12524 (N_12524,N_11941,N_11643);
xor U12525 (N_12525,N_11321,N_10550);
or U12526 (N_12526,N_11982,N_11150);
or U12527 (N_12527,N_10516,N_11336);
and U12528 (N_12528,N_11253,N_11553);
nor U12529 (N_12529,N_10728,N_11261);
and U12530 (N_12530,N_11471,N_11211);
nor U12531 (N_12531,N_11259,N_11618);
and U12532 (N_12532,N_11855,N_11029);
nand U12533 (N_12533,N_11519,N_11533);
nand U12534 (N_12534,N_11330,N_10673);
nor U12535 (N_12535,N_11116,N_10663);
nor U12536 (N_12536,N_10897,N_11219);
nor U12537 (N_12537,N_11286,N_11824);
xor U12538 (N_12538,N_11404,N_11649);
and U12539 (N_12539,N_10980,N_10827);
or U12540 (N_12540,N_11995,N_11987);
and U12541 (N_12541,N_11113,N_11771);
and U12542 (N_12542,N_10921,N_10928);
nand U12543 (N_12543,N_11703,N_11531);
nand U12544 (N_12544,N_11853,N_10718);
xor U12545 (N_12545,N_10813,N_10781);
and U12546 (N_12546,N_11380,N_10974);
or U12547 (N_12547,N_11797,N_11609);
or U12548 (N_12548,N_11145,N_10538);
xor U12549 (N_12549,N_10836,N_11705);
or U12550 (N_12550,N_11554,N_11762);
xnor U12551 (N_12551,N_11688,N_10632);
nand U12552 (N_12552,N_11165,N_11353);
xnor U12553 (N_12553,N_10579,N_10545);
nor U12554 (N_12554,N_11701,N_11402);
and U12555 (N_12555,N_11052,N_11315);
nand U12556 (N_12556,N_11022,N_11843);
nor U12557 (N_12557,N_11258,N_11711);
xnor U12558 (N_12558,N_10705,N_10622);
nand U12559 (N_12559,N_10559,N_10789);
and U12560 (N_12560,N_10893,N_10557);
nand U12561 (N_12561,N_10996,N_11486);
and U12562 (N_12562,N_10994,N_10988);
nor U12563 (N_12563,N_10597,N_10606);
nor U12564 (N_12564,N_11439,N_11970);
and U12565 (N_12565,N_10873,N_11658);
and U12566 (N_12566,N_10544,N_11781);
nor U12567 (N_12567,N_11233,N_10690);
xor U12568 (N_12568,N_10886,N_11593);
or U12569 (N_12569,N_10978,N_11383);
and U12570 (N_12570,N_11961,N_11260);
nand U12571 (N_12571,N_11901,N_11994);
or U12572 (N_12572,N_11885,N_11578);
nor U12573 (N_12573,N_10655,N_10847);
nand U12574 (N_12574,N_11570,N_11357);
nor U12575 (N_12575,N_11532,N_10841);
nor U12576 (N_12576,N_11490,N_11485);
and U12577 (N_12577,N_10696,N_11349);
xor U12578 (N_12578,N_11848,N_11224);
nor U12579 (N_12579,N_11503,N_10624);
nor U12580 (N_12580,N_10629,N_11097);
nor U12581 (N_12581,N_11507,N_11654);
and U12582 (N_12582,N_11687,N_11818);
nor U12583 (N_12583,N_10687,N_11007);
or U12584 (N_12584,N_11881,N_10855);
or U12585 (N_12585,N_10672,N_11268);
or U12586 (N_12586,N_11600,N_10807);
nand U12587 (N_12587,N_10574,N_10774);
xnor U12588 (N_12588,N_11418,N_11102);
or U12589 (N_12589,N_11870,N_11967);
or U12590 (N_12590,N_10851,N_11013);
xnor U12591 (N_12591,N_10979,N_11793);
xnor U12592 (N_12592,N_11619,N_11133);
nor U12593 (N_12593,N_10610,N_10896);
and U12594 (N_12594,N_11996,N_11171);
or U12595 (N_12595,N_11058,N_10998);
xor U12596 (N_12596,N_10630,N_11178);
nand U12597 (N_12597,N_11118,N_11930);
and U12598 (N_12598,N_11295,N_11379);
nand U12599 (N_12599,N_11833,N_10679);
and U12600 (N_12600,N_11517,N_11216);
xnor U12601 (N_12601,N_11240,N_11934);
nand U12602 (N_12602,N_10794,N_11814);
and U12603 (N_12603,N_10961,N_11300);
and U12604 (N_12604,N_11020,N_11075);
nor U12605 (N_12605,N_11974,N_10920);
nor U12606 (N_12606,N_11898,N_11293);
nor U12607 (N_12607,N_10776,N_10561);
and U12608 (N_12608,N_10698,N_11589);
nand U12609 (N_12609,N_11429,N_10877);
or U12610 (N_12610,N_11963,N_11294);
or U12611 (N_12611,N_11284,N_10944);
nand U12612 (N_12612,N_11860,N_11791);
nor U12613 (N_12613,N_10932,N_11231);
or U12614 (N_12614,N_11830,N_10564);
nor U12615 (N_12615,N_10856,N_10780);
nand U12616 (N_12616,N_11975,N_11281);
and U12617 (N_12617,N_11757,N_11291);
or U12618 (N_12618,N_10793,N_10949);
xor U12619 (N_12619,N_11988,N_11480);
nor U12620 (N_12620,N_11735,N_11562);
or U12621 (N_12621,N_11094,N_11146);
xnor U12622 (N_12622,N_10876,N_11139);
nand U12623 (N_12623,N_11483,N_11858);
xor U12624 (N_12624,N_10878,N_11874);
and U12625 (N_12625,N_11296,N_11264);
and U12626 (N_12626,N_11366,N_10849);
xnor U12627 (N_12627,N_10639,N_11010);
and U12628 (N_12628,N_10936,N_11782);
or U12629 (N_12629,N_10534,N_11939);
or U12630 (N_12630,N_11863,N_11063);
or U12631 (N_12631,N_11106,N_11908);
or U12632 (N_12632,N_10525,N_10745);
and U12633 (N_12633,N_11193,N_10621);
xor U12634 (N_12634,N_11212,N_11192);
nor U12635 (N_12635,N_11016,N_11634);
nor U12636 (N_12636,N_10535,N_11561);
and U12637 (N_12637,N_10547,N_11985);
xor U12638 (N_12638,N_10802,N_11190);
and U12639 (N_12639,N_10872,N_10784);
or U12640 (N_12640,N_11884,N_11549);
nand U12641 (N_12641,N_11290,N_10900);
nor U12642 (N_12642,N_11460,N_10694);
nand U12643 (N_12643,N_10805,N_10868);
nor U12644 (N_12644,N_10671,N_11026);
nor U12645 (N_12645,N_11799,N_11603);
xnor U12646 (N_12646,N_11937,N_11023);
or U12647 (N_12647,N_10982,N_11288);
xor U12648 (N_12648,N_11430,N_10684);
nor U12649 (N_12649,N_11560,N_10747);
or U12650 (N_12650,N_10757,N_10890);
nor U12651 (N_12651,N_11136,N_11868);
and U12652 (N_12652,N_11477,N_10914);
nand U12653 (N_12653,N_11083,N_10603);
or U12654 (N_12654,N_10584,N_10952);
nor U12655 (N_12655,N_11319,N_11055);
nor U12656 (N_12656,N_11252,N_11501);
xor U12657 (N_12657,N_11841,N_11912);
and U12658 (N_12658,N_10717,N_11088);
nor U12659 (N_12659,N_11642,N_11992);
xor U12660 (N_12660,N_11169,N_11684);
and U12661 (N_12661,N_11907,N_11585);
nand U12662 (N_12662,N_10678,N_11044);
xnor U12663 (N_12663,N_11297,N_11237);
nor U12664 (N_12664,N_10850,N_11751);
xnor U12665 (N_12665,N_10839,N_11036);
or U12666 (N_12666,N_11409,N_11747);
nor U12667 (N_12667,N_11107,N_11809);
or U12668 (N_12668,N_10677,N_11373);
and U12669 (N_12669,N_11250,N_11651);
nor U12670 (N_12670,N_10583,N_11386);
or U12671 (N_12671,N_11832,N_11929);
nand U12672 (N_12672,N_11919,N_10508);
and U12673 (N_12673,N_11512,N_11699);
xor U12674 (N_12674,N_10700,N_10523);
nor U12675 (N_12675,N_11131,N_10795);
nor U12676 (N_12676,N_11776,N_11447);
xnor U12677 (N_12677,N_10669,N_11375);
xor U12678 (N_12678,N_10779,N_11893);
nand U12679 (N_12679,N_11098,N_11307);
or U12680 (N_12680,N_10737,N_11396);
nor U12681 (N_12681,N_11729,N_11496);
xor U12682 (N_12682,N_11530,N_11698);
or U12683 (N_12683,N_11755,N_11590);
nand U12684 (N_12684,N_10697,N_10940);
and U12685 (N_12685,N_11896,N_10695);
nand U12686 (N_12686,N_10912,N_11607);
xnor U12687 (N_12687,N_11015,N_11474);
or U12688 (N_12688,N_11617,N_11851);
nor U12689 (N_12689,N_11883,N_11772);
nand U12690 (N_12690,N_11407,N_11857);
and U12691 (N_12691,N_10965,N_11846);
nor U12692 (N_12692,N_11723,N_11749);
or U12693 (N_12693,N_11915,N_10838);
nor U12694 (N_12694,N_11745,N_10549);
or U12695 (N_12695,N_11528,N_11953);
nor U12696 (N_12696,N_11662,N_11082);
and U12697 (N_12697,N_11265,N_11682);
or U12698 (N_12698,N_11278,N_11625);
and U12699 (N_12699,N_11834,N_11140);
nor U12700 (N_12700,N_11198,N_11428);
nor U12701 (N_12701,N_10715,N_10699);
xnor U12702 (N_12702,N_11156,N_10966);
or U12703 (N_12703,N_11004,N_11057);
nor U12704 (N_12704,N_10675,N_11534);
nand U12705 (N_12705,N_11913,N_11579);
and U12706 (N_12706,N_11900,N_10540);
xnor U12707 (N_12707,N_10967,N_10945);
nand U12708 (N_12708,N_11273,N_11788);
nor U12709 (N_12709,N_10654,N_10977);
nand U12710 (N_12710,N_10631,N_11798);
or U12711 (N_12711,N_11263,N_11308);
nor U12712 (N_12712,N_10562,N_10616);
nand U12713 (N_12713,N_11185,N_11505);
and U12714 (N_12714,N_10799,N_11806);
nand U12715 (N_12715,N_10973,N_10854);
nand U12716 (N_12716,N_11984,N_10659);
and U12717 (N_12717,N_10611,N_11054);
xnor U12718 (N_12718,N_11228,N_11339);
nor U12719 (N_12719,N_11274,N_11523);
nor U12720 (N_12720,N_10567,N_10668);
and U12721 (N_12721,N_10887,N_11327);
xnor U12722 (N_12722,N_10770,N_11287);
or U12723 (N_12723,N_11464,N_11196);
nand U12724 (N_12724,N_10750,N_11046);
xor U12725 (N_12725,N_10866,N_11419);
and U12726 (N_12726,N_11656,N_11612);
and U12727 (N_12727,N_11277,N_10572);
or U12728 (N_12728,N_10987,N_11072);
and U12729 (N_12729,N_11100,N_11210);
and U12730 (N_12730,N_11690,N_10527);
xnor U12731 (N_12731,N_11555,N_10537);
nand U12732 (N_12732,N_11175,N_11450);
nor U12733 (N_12733,N_10927,N_11663);
or U12734 (N_12734,N_10635,N_10628);
nand U12735 (N_12735,N_11565,N_10835);
or U12736 (N_12736,N_10786,N_10826);
or U12737 (N_12737,N_11018,N_10529);
nor U12738 (N_12738,N_11005,N_10954);
or U12739 (N_12739,N_11577,N_11416);
nor U12740 (N_12740,N_11640,N_10637);
or U12741 (N_12741,N_11248,N_10820);
or U12742 (N_12742,N_11109,N_11571);
nand U12743 (N_12743,N_11173,N_11473);
nor U12744 (N_12744,N_10922,N_11226);
and U12745 (N_12745,N_10909,N_11852);
or U12746 (N_12746,N_11808,N_11468);
or U12747 (N_12747,N_11299,N_11574);
nand U12748 (N_12748,N_11889,N_10510);
xor U12749 (N_12749,N_11385,N_10721);
and U12750 (N_12750,N_10733,N_10727);
nor U12751 (N_12751,N_11155,N_11827);
nand U12752 (N_12752,N_11763,N_11708);
xor U12753 (N_12753,N_11311,N_10621);
and U12754 (N_12754,N_10736,N_10611);
xor U12755 (N_12755,N_10804,N_11622);
or U12756 (N_12756,N_10977,N_11737);
or U12757 (N_12757,N_11547,N_11224);
nand U12758 (N_12758,N_10992,N_11879);
and U12759 (N_12759,N_11640,N_11881);
nand U12760 (N_12760,N_11646,N_10541);
or U12761 (N_12761,N_10658,N_11835);
nor U12762 (N_12762,N_10925,N_11980);
or U12763 (N_12763,N_11888,N_11452);
or U12764 (N_12764,N_10689,N_11558);
xor U12765 (N_12765,N_10958,N_11293);
or U12766 (N_12766,N_11835,N_10558);
nand U12767 (N_12767,N_11080,N_11499);
xnor U12768 (N_12768,N_11590,N_10861);
and U12769 (N_12769,N_11005,N_11293);
or U12770 (N_12770,N_10880,N_10966);
and U12771 (N_12771,N_10854,N_11712);
or U12772 (N_12772,N_10724,N_11473);
nor U12773 (N_12773,N_11850,N_11183);
or U12774 (N_12774,N_11480,N_11487);
and U12775 (N_12775,N_11795,N_11863);
nor U12776 (N_12776,N_11153,N_10771);
or U12777 (N_12777,N_10663,N_10568);
nor U12778 (N_12778,N_11563,N_10644);
and U12779 (N_12779,N_11104,N_10752);
or U12780 (N_12780,N_11189,N_10933);
nor U12781 (N_12781,N_11512,N_11315);
nor U12782 (N_12782,N_10733,N_10893);
xnor U12783 (N_12783,N_11668,N_11030);
and U12784 (N_12784,N_11486,N_10989);
and U12785 (N_12785,N_10584,N_10673);
xor U12786 (N_12786,N_10599,N_11042);
xnor U12787 (N_12787,N_11131,N_11922);
or U12788 (N_12788,N_11106,N_10750);
and U12789 (N_12789,N_11985,N_11079);
xnor U12790 (N_12790,N_11680,N_11280);
and U12791 (N_12791,N_11498,N_10535);
and U12792 (N_12792,N_11306,N_10638);
or U12793 (N_12793,N_11728,N_11167);
nand U12794 (N_12794,N_11644,N_11479);
or U12795 (N_12795,N_10605,N_11167);
or U12796 (N_12796,N_11831,N_11004);
or U12797 (N_12797,N_11735,N_11415);
and U12798 (N_12798,N_11919,N_10712);
xor U12799 (N_12799,N_10831,N_11424);
and U12800 (N_12800,N_11051,N_11770);
nor U12801 (N_12801,N_10891,N_11618);
nand U12802 (N_12802,N_10913,N_11413);
nand U12803 (N_12803,N_10816,N_11473);
and U12804 (N_12804,N_11859,N_11417);
or U12805 (N_12805,N_11846,N_10980);
xor U12806 (N_12806,N_11250,N_10550);
nor U12807 (N_12807,N_11741,N_11931);
and U12808 (N_12808,N_10577,N_11095);
or U12809 (N_12809,N_11981,N_10812);
or U12810 (N_12810,N_11713,N_11616);
nand U12811 (N_12811,N_10713,N_11128);
or U12812 (N_12812,N_10536,N_11258);
xor U12813 (N_12813,N_11496,N_10774);
xor U12814 (N_12814,N_11064,N_10684);
and U12815 (N_12815,N_11548,N_11232);
or U12816 (N_12816,N_11404,N_11914);
and U12817 (N_12817,N_10885,N_11246);
xnor U12818 (N_12818,N_11079,N_11757);
or U12819 (N_12819,N_11254,N_11132);
and U12820 (N_12820,N_11618,N_10554);
or U12821 (N_12821,N_10516,N_11192);
and U12822 (N_12822,N_11382,N_10967);
xor U12823 (N_12823,N_11207,N_11682);
nor U12824 (N_12824,N_10774,N_11702);
or U12825 (N_12825,N_11371,N_11136);
and U12826 (N_12826,N_11146,N_11565);
xor U12827 (N_12827,N_10524,N_11433);
nand U12828 (N_12828,N_11741,N_10627);
nor U12829 (N_12829,N_11546,N_11812);
and U12830 (N_12830,N_11287,N_10523);
nor U12831 (N_12831,N_10643,N_11427);
nor U12832 (N_12832,N_11546,N_11583);
or U12833 (N_12833,N_10985,N_11644);
nor U12834 (N_12834,N_10894,N_11210);
and U12835 (N_12835,N_10568,N_11489);
and U12836 (N_12836,N_11330,N_11361);
nor U12837 (N_12837,N_10943,N_11257);
and U12838 (N_12838,N_10557,N_10687);
xnor U12839 (N_12839,N_11295,N_11052);
and U12840 (N_12840,N_11245,N_11552);
nand U12841 (N_12841,N_10978,N_10852);
xor U12842 (N_12842,N_10728,N_11333);
and U12843 (N_12843,N_11636,N_11469);
nand U12844 (N_12844,N_11015,N_11080);
or U12845 (N_12845,N_10616,N_11012);
nand U12846 (N_12846,N_11038,N_11352);
xor U12847 (N_12847,N_10711,N_11044);
xnor U12848 (N_12848,N_10668,N_11019);
xor U12849 (N_12849,N_11482,N_11461);
nor U12850 (N_12850,N_10711,N_11448);
nor U12851 (N_12851,N_11015,N_11894);
and U12852 (N_12852,N_11271,N_10837);
nand U12853 (N_12853,N_11147,N_11217);
and U12854 (N_12854,N_10614,N_10635);
nor U12855 (N_12855,N_11869,N_11273);
nand U12856 (N_12856,N_10562,N_11281);
or U12857 (N_12857,N_11831,N_10682);
and U12858 (N_12858,N_10954,N_10916);
nor U12859 (N_12859,N_11840,N_11330);
or U12860 (N_12860,N_11662,N_10703);
or U12861 (N_12861,N_10766,N_11295);
or U12862 (N_12862,N_11359,N_11245);
and U12863 (N_12863,N_11652,N_10649);
and U12864 (N_12864,N_10542,N_11818);
nand U12865 (N_12865,N_11994,N_10831);
nor U12866 (N_12866,N_11134,N_10563);
xnor U12867 (N_12867,N_11278,N_10651);
nor U12868 (N_12868,N_11228,N_11611);
nor U12869 (N_12869,N_11008,N_11994);
and U12870 (N_12870,N_11775,N_11134);
or U12871 (N_12871,N_11959,N_10703);
nor U12872 (N_12872,N_11392,N_11090);
and U12873 (N_12873,N_11422,N_10622);
nor U12874 (N_12874,N_10632,N_11216);
nand U12875 (N_12875,N_11969,N_10946);
or U12876 (N_12876,N_11606,N_10550);
xnor U12877 (N_12877,N_11715,N_11579);
or U12878 (N_12878,N_11050,N_10747);
and U12879 (N_12879,N_11922,N_10676);
xor U12880 (N_12880,N_10774,N_11794);
xnor U12881 (N_12881,N_11878,N_10890);
and U12882 (N_12882,N_11755,N_11248);
nor U12883 (N_12883,N_11784,N_11688);
and U12884 (N_12884,N_11821,N_10765);
nor U12885 (N_12885,N_11363,N_11001);
xnor U12886 (N_12886,N_11770,N_11812);
and U12887 (N_12887,N_11798,N_11400);
nor U12888 (N_12888,N_11634,N_10812);
and U12889 (N_12889,N_11946,N_11647);
nor U12890 (N_12890,N_11094,N_11748);
or U12891 (N_12891,N_10843,N_11148);
xor U12892 (N_12892,N_10891,N_11736);
nand U12893 (N_12893,N_11340,N_11093);
nand U12894 (N_12894,N_11833,N_11851);
nand U12895 (N_12895,N_11132,N_11674);
xor U12896 (N_12896,N_11527,N_11113);
and U12897 (N_12897,N_11551,N_11384);
and U12898 (N_12898,N_10677,N_11523);
and U12899 (N_12899,N_11336,N_11484);
nor U12900 (N_12900,N_11873,N_10508);
xor U12901 (N_12901,N_10718,N_11571);
nor U12902 (N_12902,N_11217,N_11400);
and U12903 (N_12903,N_11413,N_11134);
xor U12904 (N_12904,N_11733,N_11757);
nand U12905 (N_12905,N_11971,N_10802);
xor U12906 (N_12906,N_10789,N_11008);
xor U12907 (N_12907,N_11554,N_11964);
nand U12908 (N_12908,N_10542,N_11167);
nand U12909 (N_12909,N_11130,N_10949);
and U12910 (N_12910,N_11292,N_10778);
and U12911 (N_12911,N_10662,N_10796);
xnor U12912 (N_12912,N_11042,N_10860);
xor U12913 (N_12913,N_11593,N_10875);
xor U12914 (N_12914,N_11366,N_10682);
nor U12915 (N_12915,N_11598,N_11185);
or U12916 (N_12916,N_10724,N_11467);
and U12917 (N_12917,N_11686,N_11420);
nand U12918 (N_12918,N_11279,N_11127);
or U12919 (N_12919,N_11755,N_10608);
and U12920 (N_12920,N_11175,N_11868);
nor U12921 (N_12921,N_10953,N_10682);
or U12922 (N_12922,N_11961,N_11703);
xor U12923 (N_12923,N_11690,N_10825);
nor U12924 (N_12924,N_11237,N_10961);
xor U12925 (N_12925,N_11685,N_10799);
nor U12926 (N_12926,N_11619,N_11841);
nand U12927 (N_12927,N_11427,N_11278);
xor U12928 (N_12928,N_11705,N_11372);
nor U12929 (N_12929,N_10677,N_11292);
nor U12930 (N_12930,N_11322,N_11631);
or U12931 (N_12931,N_11693,N_10595);
nor U12932 (N_12932,N_10889,N_10500);
or U12933 (N_12933,N_10598,N_10700);
and U12934 (N_12934,N_11340,N_11557);
nand U12935 (N_12935,N_10905,N_10721);
and U12936 (N_12936,N_10827,N_11814);
nor U12937 (N_12937,N_11177,N_11621);
xor U12938 (N_12938,N_11383,N_11654);
xor U12939 (N_12939,N_10734,N_10563);
and U12940 (N_12940,N_11150,N_10572);
or U12941 (N_12941,N_11493,N_11736);
xnor U12942 (N_12942,N_10569,N_11215);
nand U12943 (N_12943,N_11340,N_11435);
xor U12944 (N_12944,N_10700,N_11803);
nor U12945 (N_12945,N_10754,N_11234);
xor U12946 (N_12946,N_10617,N_11013);
nand U12947 (N_12947,N_10936,N_11213);
or U12948 (N_12948,N_10569,N_10643);
and U12949 (N_12949,N_10758,N_10999);
or U12950 (N_12950,N_10868,N_10734);
nor U12951 (N_12951,N_10515,N_11943);
and U12952 (N_12952,N_10967,N_10629);
and U12953 (N_12953,N_10563,N_10792);
nand U12954 (N_12954,N_11587,N_10716);
nor U12955 (N_12955,N_10742,N_11015);
nor U12956 (N_12956,N_11453,N_11547);
nor U12957 (N_12957,N_11099,N_11881);
nor U12958 (N_12958,N_11386,N_10769);
nand U12959 (N_12959,N_10848,N_11744);
and U12960 (N_12960,N_11603,N_10503);
nand U12961 (N_12961,N_10843,N_10811);
nor U12962 (N_12962,N_11051,N_11154);
nor U12963 (N_12963,N_11149,N_11838);
nor U12964 (N_12964,N_10647,N_10646);
nor U12965 (N_12965,N_11025,N_11569);
nand U12966 (N_12966,N_11632,N_11359);
and U12967 (N_12967,N_10588,N_11659);
nand U12968 (N_12968,N_10831,N_10847);
xor U12969 (N_12969,N_10834,N_11583);
nand U12970 (N_12970,N_11807,N_10765);
xnor U12971 (N_12971,N_11990,N_10901);
nand U12972 (N_12972,N_11970,N_11066);
and U12973 (N_12973,N_11088,N_11484);
xor U12974 (N_12974,N_10634,N_11317);
and U12975 (N_12975,N_11411,N_11896);
nor U12976 (N_12976,N_10950,N_11022);
nand U12977 (N_12977,N_11371,N_10580);
xor U12978 (N_12978,N_10909,N_11186);
nor U12979 (N_12979,N_11330,N_11690);
xnor U12980 (N_12980,N_11149,N_11395);
nor U12981 (N_12981,N_11823,N_10518);
and U12982 (N_12982,N_11555,N_11567);
and U12983 (N_12983,N_10931,N_11847);
nand U12984 (N_12984,N_11804,N_11164);
or U12985 (N_12985,N_11362,N_10615);
and U12986 (N_12986,N_11606,N_10707);
xnor U12987 (N_12987,N_11049,N_11265);
xor U12988 (N_12988,N_11889,N_10973);
xor U12989 (N_12989,N_11536,N_11645);
and U12990 (N_12990,N_10903,N_11662);
nand U12991 (N_12991,N_11276,N_10835);
nand U12992 (N_12992,N_11394,N_11133);
and U12993 (N_12993,N_11694,N_11821);
nand U12994 (N_12994,N_11688,N_10600);
and U12995 (N_12995,N_10597,N_11181);
nor U12996 (N_12996,N_11300,N_11268);
and U12997 (N_12997,N_11897,N_11853);
nand U12998 (N_12998,N_10747,N_10885);
nor U12999 (N_12999,N_10708,N_11270);
and U13000 (N_13000,N_11926,N_10679);
nand U13001 (N_13001,N_11931,N_11383);
or U13002 (N_13002,N_11006,N_10741);
xnor U13003 (N_13003,N_10568,N_11719);
nor U13004 (N_13004,N_11455,N_11960);
or U13005 (N_13005,N_10738,N_10758);
xnor U13006 (N_13006,N_11058,N_10790);
xnor U13007 (N_13007,N_11181,N_11215);
nand U13008 (N_13008,N_10888,N_11727);
and U13009 (N_13009,N_11308,N_11032);
and U13010 (N_13010,N_10815,N_11374);
or U13011 (N_13011,N_11754,N_11632);
or U13012 (N_13012,N_11835,N_11481);
nor U13013 (N_13013,N_11948,N_11129);
nor U13014 (N_13014,N_11440,N_11953);
nand U13015 (N_13015,N_11663,N_11664);
and U13016 (N_13016,N_11317,N_10551);
and U13017 (N_13017,N_11421,N_11979);
nand U13018 (N_13018,N_10886,N_11023);
nand U13019 (N_13019,N_10852,N_10933);
nand U13020 (N_13020,N_10670,N_11363);
nand U13021 (N_13021,N_11116,N_11585);
or U13022 (N_13022,N_11080,N_10512);
nand U13023 (N_13023,N_11355,N_11532);
nand U13024 (N_13024,N_11036,N_10514);
nand U13025 (N_13025,N_11271,N_11017);
and U13026 (N_13026,N_11066,N_11809);
nand U13027 (N_13027,N_11590,N_10879);
or U13028 (N_13028,N_10944,N_11430);
or U13029 (N_13029,N_10591,N_10817);
nand U13030 (N_13030,N_10859,N_11940);
nand U13031 (N_13031,N_11263,N_11203);
and U13032 (N_13032,N_11692,N_11929);
or U13033 (N_13033,N_10548,N_11309);
and U13034 (N_13034,N_11749,N_11237);
nor U13035 (N_13035,N_11575,N_11886);
xor U13036 (N_13036,N_10872,N_11881);
nand U13037 (N_13037,N_11156,N_11308);
nor U13038 (N_13038,N_11307,N_11072);
nand U13039 (N_13039,N_11538,N_11425);
nor U13040 (N_13040,N_10640,N_11467);
nor U13041 (N_13041,N_11630,N_11576);
and U13042 (N_13042,N_11762,N_11372);
or U13043 (N_13043,N_10645,N_10870);
nor U13044 (N_13044,N_10660,N_11633);
nor U13045 (N_13045,N_11867,N_11389);
and U13046 (N_13046,N_11433,N_10780);
xor U13047 (N_13047,N_11407,N_11968);
and U13048 (N_13048,N_11916,N_11952);
nor U13049 (N_13049,N_10654,N_11412);
nor U13050 (N_13050,N_10873,N_11165);
xor U13051 (N_13051,N_11235,N_11336);
xor U13052 (N_13052,N_11601,N_11545);
nand U13053 (N_13053,N_10959,N_11019);
or U13054 (N_13054,N_11909,N_11070);
and U13055 (N_13055,N_11207,N_10653);
or U13056 (N_13056,N_10600,N_10539);
xnor U13057 (N_13057,N_11574,N_11672);
and U13058 (N_13058,N_10956,N_10839);
and U13059 (N_13059,N_11584,N_10654);
and U13060 (N_13060,N_10534,N_10961);
or U13061 (N_13061,N_11502,N_10562);
nor U13062 (N_13062,N_11633,N_10722);
or U13063 (N_13063,N_10579,N_10945);
nand U13064 (N_13064,N_11046,N_10927);
nor U13065 (N_13065,N_11235,N_10869);
and U13066 (N_13066,N_11940,N_11189);
nand U13067 (N_13067,N_11511,N_10616);
xor U13068 (N_13068,N_11460,N_10558);
nand U13069 (N_13069,N_10850,N_11085);
xor U13070 (N_13070,N_11079,N_11175);
xor U13071 (N_13071,N_10794,N_11957);
nand U13072 (N_13072,N_10588,N_11813);
xor U13073 (N_13073,N_11761,N_11880);
nor U13074 (N_13074,N_11370,N_11047);
and U13075 (N_13075,N_11121,N_11189);
nor U13076 (N_13076,N_11970,N_11457);
and U13077 (N_13077,N_11252,N_11994);
and U13078 (N_13078,N_11996,N_11552);
and U13079 (N_13079,N_11209,N_11378);
xnor U13080 (N_13080,N_11043,N_11490);
xnor U13081 (N_13081,N_11861,N_11908);
xnor U13082 (N_13082,N_11043,N_11703);
and U13083 (N_13083,N_10839,N_10678);
nor U13084 (N_13084,N_10924,N_11505);
and U13085 (N_13085,N_11709,N_11393);
and U13086 (N_13086,N_11158,N_10894);
xnor U13087 (N_13087,N_11674,N_10666);
nor U13088 (N_13088,N_11229,N_11739);
nor U13089 (N_13089,N_10548,N_11607);
nand U13090 (N_13090,N_11255,N_11422);
or U13091 (N_13091,N_11822,N_11362);
nand U13092 (N_13092,N_11783,N_11673);
or U13093 (N_13093,N_11060,N_11870);
and U13094 (N_13094,N_11297,N_11042);
xnor U13095 (N_13095,N_11519,N_11890);
xnor U13096 (N_13096,N_10590,N_11843);
or U13097 (N_13097,N_11924,N_10819);
or U13098 (N_13098,N_11122,N_11760);
and U13099 (N_13099,N_10954,N_11343);
or U13100 (N_13100,N_10886,N_11524);
nand U13101 (N_13101,N_11065,N_10978);
and U13102 (N_13102,N_11079,N_11584);
and U13103 (N_13103,N_10960,N_11938);
and U13104 (N_13104,N_11726,N_11077);
or U13105 (N_13105,N_10555,N_10723);
and U13106 (N_13106,N_11802,N_10511);
and U13107 (N_13107,N_10766,N_10926);
or U13108 (N_13108,N_11953,N_10662);
nand U13109 (N_13109,N_11882,N_10896);
nor U13110 (N_13110,N_11556,N_11404);
and U13111 (N_13111,N_11939,N_11398);
and U13112 (N_13112,N_11459,N_11962);
nand U13113 (N_13113,N_10779,N_11107);
and U13114 (N_13114,N_11279,N_11540);
and U13115 (N_13115,N_11134,N_11504);
or U13116 (N_13116,N_11316,N_11499);
nand U13117 (N_13117,N_11295,N_11666);
nand U13118 (N_13118,N_10868,N_11022);
nand U13119 (N_13119,N_11889,N_11026);
or U13120 (N_13120,N_10544,N_11457);
nor U13121 (N_13121,N_10857,N_10647);
and U13122 (N_13122,N_10681,N_11678);
or U13123 (N_13123,N_10541,N_11991);
and U13124 (N_13124,N_10522,N_11470);
or U13125 (N_13125,N_10795,N_10755);
nor U13126 (N_13126,N_11358,N_11863);
and U13127 (N_13127,N_10502,N_11515);
or U13128 (N_13128,N_10848,N_11714);
nand U13129 (N_13129,N_10640,N_11162);
or U13130 (N_13130,N_11393,N_10532);
or U13131 (N_13131,N_11849,N_11165);
nand U13132 (N_13132,N_11707,N_11866);
and U13133 (N_13133,N_11204,N_11004);
nor U13134 (N_13134,N_11261,N_10704);
or U13135 (N_13135,N_11588,N_11683);
nor U13136 (N_13136,N_11386,N_11259);
nand U13137 (N_13137,N_11868,N_11594);
or U13138 (N_13138,N_10712,N_11245);
xor U13139 (N_13139,N_10971,N_11481);
nand U13140 (N_13140,N_11232,N_11401);
and U13141 (N_13141,N_11213,N_11431);
or U13142 (N_13142,N_11676,N_11888);
xnor U13143 (N_13143,N_10840,N_11383);
and U13144 (N_13144,N_10909,N_10633);
nor U13145 (N_13145,N_10672,N_10823);
xnor U13146 (N_13146,N_11976,N_10502);
nor U13147 (N_13147,N_11691,N_11826);
or U13148 (N_13148,N_11804,N_11778);
xnor U13149 (N_13149,N_10727,N_10503);
and U13150 (N_13150,N_11128,N_11245);
nand U13151 (N_13151,N_11843,N_10646);
xnor U13152 (N_13152,N_11763,N_11934);
and U13153 (N_13153,N_11409,N_10690);
xor U13154 (N_13154,N_11415,N_10868);
or U13155 (N_13155,N_11544,N_11715);
or U13156 (N_13156,N_11685,N_11526);
or U13157 (N_13157,N_10745,N_11527);
or U13158 (N_13158,N_10807,N_11188);
nand U13159 (N_13159,N_11134,N_10938);
nand U13160 (N_13160,N_11283,N_11784);
and U13161 (N_13161,N_11061,N_11682);
or U13162 (N_13162,N_11650,N_11503);
or U13163 (N_13163,N_11464,N_10741);
nor U13164 (N_13164,N_11833,N_10848);
and U13165 (N_13165,N_10789,N_10879);
nand U13166 (N_13166,N_11808,N_11588);
xor U13167 (N_13167,N_11521,N_11118);
xnor U13168 (N_13168,N_11395,N_11910);
nor U13169 (N_13169,N_11555,N_11955);
or U13170 (N_13170,N_11252,N_11081);
nand U13171 (N_13171,N_11649,N_11953);
xor U13172 (N_13172,N_11102,N_11466);
nand U13173 (N_13173,N_11155,N_10519);
or U13174 (N_13174,N_11812,N_10664);
nand U13175 (N_13175,N_10607,N_11882);
or U13176 (N_13176,N_10955,N_11729);
nor U13177 (N_13177,N_11566,N_10531);
nor U13178 (N_13178,N_10938,N_10614);
nor U13179 (N_13179,N_11328,N_10718);
xor U13180 (N_13180,N_10845,N_11911);
xor U13181 (N_13181,N_10597,N_10779);
nor U13182 (N_13182,N_10885,N_10722);
xor U13183 (N_13183,N_11735,N_11731);
nor U13184 (N_13184,N_10512,N_11911);
nor U13185 (N_13185,N_11641,N_11702);
nor U13186 (N_13186,N_11146,N_11779);
and U13187 (N_13187,N_11285,N_10904);
nand U13188 (N_13188,N_11836,N_11060);
nand U13189 (N_13189,N_10925,N_11379);
or U13190 (N_13190,N_10969,N_10770);
nor U13191 (N_13191,N_10624,N_10970);
or U13192 (N_13192,N_10982,N_11819);
or U13193 (N_13193,N_11662,N_10734);
nand U13194 (N_13194,N_11740,N_10508);
nand U13195 (N_13195,N_11610,N_11468);
xor U13196 (N_13196,N_11949,N_10866);
and U13197 (N_13197,N_11757,N_10719);
nor U13198 (N_13198,N_11122,N_11533);
xnor U13199 (N_13199,N_11897,N_11629);
nand U13200 (N_13200,N_10891,N_11251);
nor U13201 (N_13201,N_10870,N_11716);
nor U13202 (N_13202,N_10677,N_10631);
nand U13203 (N_13203,N_11663,N_11738);
or U13204 (N_13204,N_11420,N_11288);
or U13205 (N_13205,N_11373,N_11990);
nor U13206 (N_13206,N_10533,N_11262);
or U13207 (N_13207,N_11228,N_11096);
nor U13208 (N_13208,N_11184,N_10892);
nor U13209 (N_13209,N_11312,N_10585);
and U13210 (N_13210,N_11518,N_10599);
and U13211 (N_13211,N_11474,N_11082);
nor U13212 (N_13212,N_10728,N_11510);
or U13213 (N_13213,N_10875,N_11868);
nand U13214 (N_13214,N_10647,N_10743);
nand U13215 (N_13215,N_11959,N_10986);
nor U13216 (N_13216,N_11761,N_11823);
nor U13217 (N_13217,N_10641,N_11349);
nand U13218 (N_13218,N_11059,N_11798);
and U13219 (N_13219,N_10971,N_11671);
nand U13220 (N_13220,N_11016,N_11788);
xnor U13221 (N_13221,N_11253,N_11488);
xnor U13222 (N_13222,N_11928,N_11672);
or U13223 (N_13223,N_11669,N_10766);
nor U13224 (N_13224,N_11881,N_10937);
nor U13225 (N_13225,N_11734,N_11245);
xnor U13226 (N_13226,N_10858,N_11917);
nand U13227 (N_13227,N_11495,N_11472);
or U13228 (N_13228,N_11497,N_11648);
nor U13229 (N_13229,N_11450,N_11178);
and U13230 (N_13230,N_11795,N_11787);
nand U13231 (N_13231,N_10652,N_11437);
nand U13232 (N_13232,N_10786,N_10906);
and U13233 (N_13233,N_10590,N_11756);
xor U13234 (N_13234,N_10674,N_11749);
nor U13235 (N_13235,N_11286,N_10929);
xor U13236 (N_13236,N_11650,N_10970);
and U13237 (N_13237,N_11432,N_11786);
nand U13238 (N_13238,N_11537,N_10742);
and U13239 (N_13239,N_11123,N_10942);
or U13240 (N_13240,N_11732,N_11707);
and U13241 (N_13241,N_11680,N_10524);
xor U13242 (N_13242,N_11075,N_11821);
nor U13243 (N_13243,N_11940,N_11878);
xor U13244 (N_13244,N_10901,N_11342);
and U13245 (N_13245,N_10765,N_11613);
and U13246 (N_13246,N_11857,N_11080);
xnor U13247 (N_13247,N_11233,N_10613);
or U13248 (N_13248,N_11199,N_11694);
nor U13249 (N_13249,N_11101,N_11237);
and U13250 (N_13250,N_11117,N_11489);
nor U13251 (N_13251,N_11206,N_11470);
nand U13252 (N_13252,N_10975,N_11272);
xnor U13253 (N_13253,N_11797,N_11168);
or U13254 (N_13254,N_11165,N_11046);
or U13255 (N_13255,N_11209,N_11219);
or U13256 (N_13256,N_10852,N_10820);
xor U13257 (N_13257,N_11482,N_10789);
or U13258 (N_13258,N_10877,N_11847);
nand U13259 (N_13259,N_10831,N_11307);
and U13260 (N_13260,N_10773,N_11501);
or U13261 (N_13261,N_11184,N_11239);
nand U13262 (N_13262,N_11086,N_11336);
xnor U13263 (N_13263,N_11926,N_11518);
xor U13264 (N_13264,N_11578,N_11824);
xor U13265 (N_13265,N_11752,N_11338);
nand U13266 (N_13266,N_10671,N_11355);
xnor U13267 (N_13267,N_11482,N_10844);
and U13268 (N_13268,N_10673,N_11775);
nand U13269 (N_13269,N_10924,N_11221);
xnor U13270 (N_13270,N_11403,N_10839);
nor U13271 (N_13271,N_11563,N_11925);
xnor U13272 (N_13272,N_11390,N_11623);
nand U13273 (N_13273,N_10576,N_11427);
nor U13274 (N_13274,N_11820,N_10552);
and U13275 (N_13275,N_11097,N_10835);
nor U13276 (N_13276,N_11445,N_10870);
nor U13277 (N_13277,N_11392,N_11010);
xnor U13278 (N_13278,N_11468,N_11221);
or U13279 (N_13279,N_10535,N_11221);
or U13280 (N_13280,N_11703,N_11591);
nor U13281 (N_13281,N_11395,N_10941);
and U13282 (N_13282,N_10750,N_10534);
and U13283 (N_13283,N_10741,N_11880);
nand U13284 (N_13284,N_10546,N_11996);
and U13285 (N_13285,N_11496,N_10594);
nand U13286 (N_13286,N_11860,N_11309);
nor U13287 (N_13287,N_11547,N_11942);
nor U13288 (N_13288,N_11978,N_10933);
or U13289 (N_13289,N_11615,N_10529);
nor U13290 (N_13290,N_11808,N_10581);
xnor U13291 (N_13291,N_11702,N_11367);
nor U13292 (N_13292,N_11751,N_11882);
nor U13293 (N_13293,N_10820,N_11680);
nor U13294 (N_13294,N_11987,N_10615);
nand U13295 (N_13295,N_11334,N_10615);
or U13296 (N_13296,N_11151,N_11698);
xor U13297 (N_13297,N_11912,N_11164);
nand U13298 (N_13298,N_11153,N_11222);
or U13299 (N_13299,N_11527,N_10845);
nor U13300 (N_13300,N_10842,N_11756);
xnor U13301 (N_13301,N_11317,N_11458);
nand U13302 (N_13302,N_11153,N_10537);
or U13303 (N_13303,N_11732,N_10724);
or U13304 (N_13304,N_11525,N_10720);
nor U13305 (N_13305,N_11694,N_10952);
or U13306 (N_13306,N_10527,N_10653);
nand U13307 (N_13307,N_10526,N_11352);
or U13308 (N_13308,N_11773,N_11980);
nor U13309 (N_13309,N_11904,N_10782);
xor U13310 (N_13310,N_10717,N_10921);
xor U13311 (N_13311,N_11300,N_11040);
nor U13312 (N_13312,N_11495,N_11402);
nand U13313 (N_13313,N_10851,N_10737);
xor U13314 (N_13314,N_10822,N_10837);
nor U13315 (N_13315,N_11986,N_10569);
xor U13316 (N_13316,N_11854,N_11183);
or U13317 (N_13317,N_11923,N_11583);
xor U13318 (N_13318,N_11763,N_11805);
nor U13319 (N_13319,N_11798,N_11521);
and U13320 (N_13320,N_11877,N_11663);
nand U13321 (N_13321,N_10531,N_11891);
and U13322 (N_13322,N_11302,N_11984);
nand U13323 (N_13323,N_10540,N_10513);
xor U13324 (N_13324,N_11385,N_10822);
or U13325 (N_13325,N_10945,N_11202);
xnor U13326 (N_13326,N_11471,N_10852);
or U13327 (N_13327,N_11660,N_10867);
or U13328 (N_13328,N_11061,N_11233);
and U13329 (N_13329,N_11879,N_11273);
or U13330 (N_13330,N_10782,N_10871);
xor U13331 (N_13331,N_11618,N_11633);
nand U13332 (N_13332,N_11194,N_10504);
and U13333 (N_13333,N_10961,N_11545);
xor U13334 (N_13334,N_11806,N_11260);
nand U13335 (N_13335,N_11695,N_10907);
nor U13336 (N_13336,N_10834,N_10870);
or U13337 (N_13337,N_10746,N_11209);
nand U13338 (N_13338,N_11803,N_11722);
nand U13339 (N_13339,N_10828,N_11668);
xnor U13340 (N_13340,N_11070,N_11316);
xnor U13341 (N_13341,N_11865,N_11722);
nor U13342 (N_13342,N_11890,N_11624);
or U13343 (N_13343,N_11679,N_11189);
and U13344 (N_13344,N_10729,N_11798);
nor U13345 (N_13345,N_11751,N_11894);
nand U13346 (N_13346,N_11637,N_11258);
or U13347 (N_13347,N_11423,N_10688);
and U13348 (N_13348,N_10839,N_10996);
xor U13349 (N_13349,N_11088,N_11899);
nand U13350 (N_13350,N_11413,N_11310);
or U13351 (N_13351,N_11253,N_10999);
and U13352 (N_13352,N_11585,N_10955);
or U13353 (N_13353,N_11879,N_10587);
or U13354 (N_13354,N_11599,N_10811);
xor U13355 (N_13355,N_11758,N_10981);
nor U13356 (N_13356,N_11962,N_11752);
or U13357 (N_13357,N_11284,N_11914);
nand U13358 (N_13358,N_11605,N_10720);
nand U13359 (N_13359,N_11519,N_11118);
nor U13360 (N_13360,N_11074,N_11730);
nor U13361 (N_13361,N_11157,N_11711);
xor U13362 (N_13362,N_10740,N_10877);
nor U13363 (N_13363,N_11703,N_10632);
nor U13364 (N_13364,N_11421,N_11294);
or U13365 (N_13365,N_10820,N_11020);
and U13366 (N_13366,N_11195,N_11523);
nand U13367 (N_13367,N_10540,N_10530);
xnor U13368 (N_13368,N_11021,N_11718);
or U13369 (N_13369,N_11207,N_11072);
nor U13370 (N_13370,N_10530,N_10649);
and U13371 (N_13371,N_11442,N_11816);
nor U13372 (N_13372,N_11744,N_11721);
nor U13373 (N_13373,N_10530,N_11471);
nor U13374 (N_13374,N_11369,N_11196);
nor U13375 (N_13375,N_10573,N_11066);
or U13376 (N_13376,N_11932,N_10908);
xor U13377 (N_13377,N_11752,N_10995);
nand U13378 (N_13378,N_10572,N_10650);
and U13379 (N_13379,N_10690,N_11283);
and U13380 (N_13380,N_11713,N_11283);
nor U13381 (N_13381,N_11590,N_11434);
nand U13382 (N_13382,N_10771,N_10523);
nor U13383 (N_13383,N_11186,N_10921);
and U13384 (N_13384,N_11667,N_11110);
nand U13385 (N_13385,N_11985,N_11816);
nand U13386 (N_13386,N_11288,N_11768);
and U13387 (N_13387,N_11136,N_11650);
or U13388 (N_13388,N_11438,N_10503);
or U13389 (N_13389,N_11155,N_11315);
xnor U13390 (N_13390,N_11885,N_10686);
xor U13391 (N_13391,N_10639,N_11909);
nand U13392 (N_13392,N_11905,N_11110);
nand U13393 (N_13393,N_11017,N_11513);
or U13394 (N_13394,N_10868,N_10848);
nand U13395 (N_13395,N_10749,N_10539);
or U13396 (N_13396,N_10922,N_11396);
nor U13397 (N_13397,N_10770,N_11622);
nand U13398 (N_13398,N_10520,N_11165);
and U13399 (N_13399,N_11894,N_10698);
or U13400 (N_13400,N_11596,N_10810);
and U13401 (N_13401,N_10703,N_10556);
xnor U13402 (N_13402,N_11970,N_10738);
xnor U13403 (N_13403,N_10718,N_10845);
nor U13404 (N_13404,N_11060,N_11807);
or U13405 (N_13405,N_11914,N_10715);
and U13406 (N_13406,N_11917,N_10760);
nand U13407 (N_13407,N_10781,N_11471);
nor U13408 (N_13408,N_10815,N_11824);
nand U13409 (N_13409,N_10655,N_11507);
or U13410 (N_13410,N_11448,N_10845);
nor U13411 (N_13411,N_11902,N_11435);
nor U13412 (N_13412,N_11126,N_10954);
nor U13413 (N_13413,N_11251,N_11427);
or U13414 (N_13414,N_11669,N_11967);
or U13415 (N_13415,N_11393,N_10740);
xnor U13416 (N_13416,N_11690,N_11029);
and U13417 (N_13417,N_11552,N_11361);
nand U13418 (N_13418,N_11427,N_10917);
nor U13419 (N_13419,N_11784,N_11213);
xor U13420 (N_13420,N_11791,N_11420);
or U13421 (N_13421,N_11035,N_11060);
or U13422 (N_13422,N_11644,N_10552);
nor U13423 (N_13423,N_10929,N_11541);
nor U13424 (N_13424,N_11828,N_11380);
nor U13425 (N_13425,N_11930,N_11150);
nor U13426 (N_13426,N_11331,N_11847);
and U13427 (N_13427,N_11465,N_11710);
nand U13428 (N_13428,N_11249,N_10926);
nand U13429 (N_13429,N_10852,N_10731);
nand U13430 (N_13430,N_11235,N_11906);
nor U13431 (N_13431,N_11007,N_11904);
nand U13432 (N_13432,N_11552,N_10557);
nand U13433 (N_13433,N_11057,N_10760);
nand U13434 (N_13434,N_10507,N_11077);
nor U13435 (N_13435,N_11761,N_11866);
or U13436 (N_13436,N_10790,N_10524);
or U13437 (N_13437,N_10718,N_10899);
xnor U13438 (N_13438,N_10546,N_11880);
nor U13439 (N_13439,N_10721,N_11974);
and U13440 (N_13440,N_11636,N_11814);
nand U13441 (N_13441,N_11018,N_11200);
xor U13442 (N_13442,N_11672,N_10716);
or U13443 (N_13443,N_10595,N_11524);
xnor U13444 (N_13444,N_11657,N_10539);
and U13445 (N_13445,N_10771,N_11743);
nor U13446 (N_13446,N_11959,N_11647);
nand U13447 (N_13447,N_11484,N_11172);
or U13448 (N_13448,N_11074,N_11814);
or U13449 (N_13449,N_10517,N_11661);
or U13450 (N_13450,N_10586,N_10589);
and U13451 (N_13451,N_11386,N_11153);
or U13452 (N_13452,N_11618,N_10699);
or U13453 (N_13453,N_11354,N_11579);
or U13454 (N_13454,N_11843,N_11424);
nand U13455 (N_13455,N_11826,N_11011);
xor U13456 (N_13456,N_11691,N_11184);
nand U13457 (N_13457,N_11932,N_11778);
nor U13458 (N_13458,N_11719,N_11607);
nor U13459 (N_13459,N_11387,N_10604);
or U13460 (N_13460,N_11654,N_11460);
nand U13461 (N_13461,N_11767,N_11893);
and U13462 (N_13462,N_10938,N_11201);
nand U13463 (N_13463,N_11661,N_11512);
xnor U13464 (N_13464,N_10505,N_11319);
and U13465 (N_13465,N_11239,N_11788);
nand U13466 (N_13466,N_10901,N_10836);
nor U13467 (N_13467,N_10782,N_11155);
nor U13468 (N_13468,N_10749,N_11048);
nor U13469 (N_13469,N_11701,N_10545);
and U13470 (N_13470,N_11758,N_11511);
nand U13471 (N_13471,N_10927,N_11684);
and U13472 (N_13472,N_11681,N_11016);
and U13473 (N_13473,N_11389,N_11078);
or U13474 (N_13474,N_11081,N_11095);
or U13475 (N_13475,N_10957,N_11223);
nor U13476 (N_13476,N_11965,N_10721);
nand U13477 (N_13477,N_11985,N_11763);
nand U13478 (N_13478,N_11765,N_11989);
and U13479 (N_13479,N_11394,N_11391);
nor U13480 (N_13480,N_10914,N_11958);
or U13481 (N_13481,N_10533,N_10748);
nand U13482 (N_13482,N_11965,N_10638);
nor U13483 (N_13483,N_11911,N_10936);
nor U13484 (N_13484,N_11016,N_10836);
nand U13485 (N_13485,N_11084,N_11901);
xor U13486 (N_13486,N_11251,N_11019);
or U13487 (N_13487,N_11146,N_11678);
xnor U13488 (N_13488,N_11200,N_11977);
nor U13489 (N_13489,N_10877,N_10776);
and U13490 (N_13490,N_11874,N_10749);
nor U13491 (N_13491,N_11536,N_10633);
nand U13492 (N_13492,N_10609,N_10532);
nor U13493 (N_13493,N_10774,N_10599);
nand U13494 (N_13494,N_11125,N_10944);
or U13495 (N_13495,N_11623,N_11160);
and U13496 (N_13496,N_10858,N_10834);
nand U13497 (N_13497,N_11593,N_11293);
or U13498 (N_13498,N_10596,N_10651);
nand U13499 (N_13499,N_10965,N_11852);
or U13500 (N_13500,N_12297,N_13395);
nand U13501 (N_13501,N_13220,N_12856);
and U13502 (N_13502,N_12109,N_13437);
nand U13503 (N_13503,N_12027,N_12438);
nand U13504 (N_13504,N_12202,N_12200);
and U13505 (N_13505,N_12127,N_12686);
or U13506 (N_13506,N_12428,N_13269);
nand U13507 (N_13507,N_12245,N_13007);
xnor U13508 (N_13508,N_13108,N_12595);
or U13509 (N_13509,N_12383,N_13093);
xor U13510 (N_13510,N_13258,N_13085);
and U13511 (N_13511,N_12650,N_12267);
xnor U13512 (N_13512,N_13243,N_13058);
or U13513 (N_13513,N_12400,N_12249);
nand U13514 (N_13514,N_12450,N_12862);
and U13515 (N_13515,N_12560,N_12179);
xor U13516 (N_13516,N_12644,N_13281);
nand U13517 (N_13517,N_12948,N_12557);
nor U13518 (N_13518,N_12011,N_12633);
or U13519 (N_13519,N_12725,N_12454);
and U13520 (N_13520,N_13337,N_12547);
xnor U13521 (N_13521,N_13128,N_13231);
or U13522 (N_13522,N_13286,N_13390);
nand U13523 (N_13523,N_13248,N_13009);
and U13524 (N_13524,N_12531,N_12185);
nand U13525 (N_13525,N_13347,N_13252);
nor U13526 (N_13526,N_12281,N_13104);
nor U13527 (N_13527,N_12268,N_13278);
nand U13528 (N_13528,N_13371,N_12242);
nand U13529 (N_13529,N_13367,N_13134);
or U13530 (N_13530,N_13218,N_13228);
or U13531 (N_13531,N_13124,N_12887);
xnor U13532 (N_13532,N_13296,N_12558);
and U13533 (N_13533,N_13202,N_13022);
xor U13534 (N_13534,N_13436,N_12133);
xnor U13535 (N_13535,N_12324,N_12512);
and U13536 (N_13536,N_13010,N_12304);
nand U13537 (N_13537,N_12715,N_12660);
or U13538 (N_13538,N_13451,N_12535);
nand U13539 (N_13539,N_13335,N_13234);
xnor U13540 (N_13540,N_13315,N_12357);
nand U13541 (N_13541,N_12780,N_12192);
nor U13542 (N_13542,N_13447,N_13377);
nand U13543 (N_13543,N_13191,N_12243);
nand U13544 (N_13544,N_12565,N_12571);
and U13545 (N_13545,N_13097,N_13397);
or U13546 (N_13546,N_12122,N_13272);
or U13547 (N_13547,N_13055,N_13485);
xnor U13548 (N_13548,N_13496,N_12797);
nor U13549 (N_13549,N_12128,N_12718);
nor U13550 (N_13550,N_12890,N_12076);
and U13551 (N_13551,N_13380,N_13419);
and U13552 (N_13552,N_13440,N_12012);
nand U13553 (N_13553,N_13090,N_12375);
and U13554 (N_13554,N_12629,N_12951);
nor U13555 (N_13555,N_12619,N_12177);
xor U13556 (N_13556,N_12017,N_12716);
and U13557 (N_13557,N_13136,N_13471);
nand U13558 (N_13558,N_12618,N_13458);
or U13559 (N_13559,N_12740,N_13235);
nand U13560 (N_13560,N_12988,N_13098);
nor U13561 (N_13561,N_13382,N_12298);
xor U13562 (N_13562,N_13219,N_12624);
nor U13563 (N_13563,N_12223,N_12980);
and U13564 (N_13564,N_12572,N_12782);
or U13565 (N_13565,N_12908,N_12150);
and U13566 (N_13566,N_13265,N_12730);
nor U13567 (N_13567,N_12592,N_12671);
and U13568 (N_13568,N_12057,N_12478);
nand U13569 (N_13569,N_12878,N_12498);
or U13570 (N_13570,N_12308,N_12462);
or U13571 (N_13571,N_12749,N_13432);
xor U13572 (N_13572,N_13161,N_12599);
and U13573 (N_13573,N_12032,N_13037);
xor U13574 (N_13574,N_12670,N_13307);
xor U13575 (N_13575,N_12882,N_12938);
nor U13576 (N_13576,N_12879,N_12141);
or U13577 (N_13577,N_13147,N_12616);
or U13578 (N_13578,N_12313,N_12186);
or U13579 (N_13579,N_12374,N_12861);
xor U13580 (N_13580,N_12175,N_12905);
nor U13581 (N_13581,N_13130,N_13329);
and U13582 (N_13582,N_12679,N_12501);
nand U13583 (N_13583,N_13424,N_13207);
and U13584 (N_13584,N_12408,N_13308);
nor U13585 (N_13585,N_12567,N_12528);
nand U13586 (N_13586,N_13160,N_12802);
xor U13587 (N_13587,N_12292,N_13164);
and U13588 (N_13588,N_12077,N_12800);
and U13589 (N_13589,N_12659,N_12404);
nand U13590 (N_13590,N_12845,N_12098);
nand U13591 (N_13591,N_12522,N_12411);
and U13592 (N_13592,N_12350,N_12822);
and U13593 (N_13593,N_12700,N_13166);
xor U13594 (N_13594,N_12688,N_13123);
nand U13595 (N_13595,N_12351,N_13324);
nor U13596 (N_13596,N_13443,N_12915);
nor U13597 (N_13597,N_12423,N_12663);
nor U13598 (N_13598,N_12162,N_12135);
and U13599 (N_13599,N_12768,N_12341);
xor U13600 (N_13600,N_12702,N_12452);
xnor U13601 (N_13601,N_12164,N_12804);
nor U13602 (N_13602,N_12769,N_12369);
nor U13603 (N_13603,N_12446,N_12442);
and U13604 (N_13604,N_13088,N_13226);
and U13605 (N_13605,N_12262,N_12503);
xor U13606 (N_13606,N_13195,N_12614);
xnor U13607 (N_13607,N_12643,N_12919);
nor U13608 (N_13608,N_12854,N_13035);
xnor U13609 (N_13609,N_12068,N_12414);
nand U13610 (N_13610,N_12950,N_13407);
nor U13611 (N_13611,N_13043,N_12534);
and U13612 (N_13612,N_12778,N_12847);
nor U13613 (N_13613,N_12604,N_13215);
nand U13614 (N_13614,N_13423,N_13473);
nor U13615 (N_13615,N_13455,N_12859);
and U13616 (N_13616,N_13211,N_12646);
nand U13617 (N_13617,N_12934,N_12603);
nor U13618 (N_13618,N_13236,N_13000);
xor U13619 (N_13619,N_12367,N_13205);
and U13620 (N_13620,N_12445,N_12582);
and U13621 (N_13621,N_12259,N_12566);
nand U13622 (N_13622,N_12347,N_12102);
nand U13623 (N_13623,N_13177,N_12026);
and U13624 (N_13624,N_12568,N_13071);
and U13625 (N_13625,N_13498,N_12140);
or U13626 (N_13626,N_12244,N_13320);
nand U13627 (N_13627,N_12353,N_13312);
and U13628 (N_13628,N_13421,N_12721);
or U13629 (N_13629,N_12342,N_12286);
xor U13630 (N_13630,N_13273,N_12987);
nand U13631 (N_13631,N_12540,N_12507);
nand U13632 (N_13632,N_12332,N_12349);
nand U13633 (N_13633,N_12830,N_12553);
or U13634 (N_13634,N_13365,N_12429);
and U13635 (N_13635,N_13227,N_12902);
and U13636 (N_13636,N_13404,N_12387);
nor U13637 (N_13637,N_13012,N_13350);
and U13638 (N_13638,N_13334,N_12738);
xnor U13639 (N_13639,N_13045,N_13003);
nor U13640 (N_13640,N_13261,N_12230);
nor U13641 (N_13641,N_12527,N_12166);
nor U13642 (N_13642,N_12711,N_13360);
nor U13643 (N_13643,N_13185,N_12380);
or U13644 (N_13644,N_12046,N_13398);
xor U13645 (N_13645,N_12877,N_12471);
and U13646 (N_13646,N_12481,N_12636);
nor U13647 (N_13647,N_12723,N_12838);
and U13648 (N_13648,N_12194,N_12783);
or U13649 (N_13649,N_13260,N_12699);
nor U13650 (N_13650,N_12279,N_12080);
or U13651 (N_13651,N_13283,N_12969);
xor U13652 (N_13652,N_12170,N_13196);
or U13653 (N_13653,N_12470,N_12779);
nand U13654 (N_13654,N_12147,N_12682);
xnor U13655 (N_13655,N_13490,N_12536);
and U13656 (N_13656,N_13370,N_12745);
or U13657 (N_13657,N_12271,N_12248);
or U13658 (N_13658,N_12791,N_12755);
nand U13659 (N_13659,N_12295,N_12456);
nor U13660 (N_13660,N_12921,N_12417);
or U13661 (N_13661,N_12863,N_12519);
nor U13662 (N_13662,N_12918,N_12649);
xor U13663 (N_13663,N_12786,N_12897);
or U13664 (N_13664,N_12421,N_12287);
and U13665 (N_13665,N_12216,N_12504);
or U13666 (N_13666,N_13294,N_12597);
or U13667 (N_13667,N_12168,N_12656);
xor U13668 (N_13668,N_12072,N_12666);
or U13669 (N_13669,N_12899,N_12541);
nand U13670 (N_13670,N_13024,N_13415);
or U13671 (N_13671,N_13408,N_12117);
nor U13672 (N_13672,N_12161,N_12479);
nor U13673 (N_13673,N_13379,N_12864);
or U13674 (N_13674,N_12484,N_12420);
or U13675 (N_13675,N_12215,N_13494);
nor U13676 (N_13676,N_13391,N_12173);
and U13677 (N_13677,N_12491,N_12895);
or U13678 (N_13678,N_12195,N_12538);
nor U13679 (N_13679,N_13306,N_13246);
or U13680 (N_13680,N_12187,N_12761);
and U13681 (N_13681,N_12600,N_12178);
and U13682 (N_13682,N_12336,N_13348);
nor U13683 (N_13683,N_13204,N_12205);
xor U13684 (N_13684,N_12952,N_12632);
nor U13685 (N_13685,N_13345,N_13210);
or U13686 (N_13686,N_12517,N_12589);
nand U13687 (N_13687,N_12240,N_12916);
nand U13688 (N_13688,N_13461,N_13474);
xnor U13689 (N_13689,N_13146,N_12118);
or U13690 (N_13690,N_13254,N_13300);
nor U13691 (N_13691,N_13028,N_13291);
and U13692 (N_13692,N_12196,N_12078);
nand U13693 (N_13693,N_13141,N_13378);
or U13694 (N_13694,N_12044,N_13113);
or U13695 (N_13695,N_13358,N_13425);
nand U13696 (N_13696,N_12193,N_12056);
and U13697 (N_13697,N_12169,N_12967);
xnor U13698 (N_13698,N_13107,N_12826);
and U13699 (N_13699,N_12494,N_13499);
nand U13700 (N_13700,N_12767,N_12326);
nand U13701 (N_13701,N_13187,N_12555);
nand U13702 (N_13702,N_12627,N_12642);
or U13703 (N_13703,N_13478,N_13014);
xor U13704 (N_13704,N_12694,N_13288);
and U13705 (N_13705,N_12440,N_12208);
xnor U13706 (N_13706,N_12941,N_12100);
and U13707 (N_13707,N_12285,N_13285);
xor U13708 (N_13708,N_13302,N_12924);
and U13709 (N_13709,N_12110,N_12134);
nor U13710 (N_13710,N_12483,N_13322);
or U13711 (N_13711,N_12562,N_12070);
or U13712 (N_13712,N_13148,N_12319);
and U13713 (N_13713,N_12638,N_13033);
and U13714 (N_13714,N_12805,N_12485);
xnor U13715 (N_13715,N_13433,N_12777);
and U13716 (N_13716,N_12698,N_12739);
nor U13717 (N_13717,N_12042,N_12338);
or U13718 (N_13718,N_12385,N_12238);
nand U13719 (N_13719,N_12611,N_12872);
and U13720 (N_13720,N_12453,N_13198);
nor U13721 (N_13721,N_12690,N_12418);
xor U13722 (N_13722,N_12296,N_12183);
xor U13723 (N_13723,N_12576,N_12607);
or U13724 (N_13724,N_12628,N_13282);
nor U13725 (N_13725,N_12706,N_13075);
or U13726 (N_13726,N_12900,N_13344);
or U13727 (N_13727,N_12551,N_13495);
nor U13728 (N_13728,N_12419,N_12676);
xor U13729 (N_13729,N_13165,N_13080);
or U13730 (N_13730,N_13118,N_12167);
nand U13731 (N_13731,N_12224,N_12620);
and U13732 (N_13732,N_12731,N_12957);
xor U13733 (N_13733,N_12697,N_12505);
or U13734 (N_13734,N_12305,N_13116);
xor U13735 (N_13735,N_13190,N_12691);
or U13736 (N_13736,N_12831,N_13483);
and U13737 (N_13737,N_12953,N_12325);
nand U13738 (N_13738,N_13405,N_12554);
and U13739 (N_13739,N_12047,N_12609);
nand U13740 (N_13740,N_12065,N_12762);
and U13741 (N_13741,N_12180,N_13083);
and U13742 (N_13742,N_12823,N_13135);
xnor U13743 (N_13743,N_12019,N_12149);
nand U13744 (N_13744,N_13456,N_12358);
nor U13745 (N_13745,N_13073,N_12641);
nor U13746 (N_13746,N_12490,N_12801);
or U13747 (N_13747,N_12596,N_12280);
and U13748 (N_13748,N_12940,N_12311);
or U13749 (N_13749,N_12949,N_12138);
and U13750 (N_13750,N_12055,N_12307);
nor U13751 (N_13751,N_13152,N_12502);
nor U13752 (N_13752,N_13127,N_12947);
nand U13753 (N_13753,N_12278,N_12093);
nand U13754 (N_13754,N_12943,N_13062);
nor U13755 (N_13755,N_12371,N_12997);
nor U13756 (N_13756,N_12936,N_12549);
or U13757 (N_13757,N_13042,N_13289);
nand U13758 (N_13758,N_12018,N_12159);
or U13759 (N_13759,N_12766,N_12008);
xor U13760 (N_13760,N_12964,N_13364);
xnor U13761 (N_13761,N_13239,N_12376);
nor U13762 (N_13762,N_13318,N_13102);
nand U13763 (N_13763,N_13203,N_12929);
or U13764 (N_13764,N_13132,N_12293);
and U13765 (N_13765,N_12561,N_12913);
or U13766 (N_13766,N_13048,N_12069);
xor U13767 (N_13767,N_12868,N_13287);
xor U13768 (N_13768,N_13067,N_12984);
xnor U13769 (N_13769,N_12747,N_12867);
and U13770 (N_13770,N_12724,N_12335);
nand U13771 (N_13771,N_12412,N_12040);
xor U13772 (N_13772,N_13326,N_12584);
xnor U13773 (N_13773,N_12955,N_12130);
nand U13774 (N_13774,N_13137,N_13275);
xnor U13775 (N_13775,N_12765,N_12617);
xnor U13776 (N_13776,N_12894,N_12962);
xor U13777 (N_13777,N_13303,N_13180);
nor U13778 (N_13778,N_12651,N_12521);
or U13779 (N_13779,N_13394,N_12689);
and U13780 (N_13780,N_13212,N_13155);
or U13781 (N_13781,N_12207,N_12045);
xor U13782 (N_13782,N_12085,N_12492);
xor U13783 (N_13783,N_12733,N_12709);
and U13784 (N_13784,N_13004,N_12086);
nor U13785 (N_13785,N_12935,N_13050);
xnor U13786 (N_13786,N_12577,N_13120);
nor U13787 (N_13787,N_13341,N_12382);
xnor U13788 (N_13788,N_13056,N_12105);
nor U13789 (N_13789,N_13078,N_13016);
nor U13790 (N_13790,N_13030,N_12737);
or U13791 (N_13791,N_12090,N_12920);
nor U13792 (N_13792,N_12493,N_12214);
nor U13793 (N_13793,N_13053,N_12707);
and U13794 (N_13794,N_12129,N_12176);
xor U13795 (N_13795,N_13314,N_12436);
nor U13796 (N_13796,N_12610,N_12282);
or U13797 (N_13797,N_12966,N_13416);
and U13798 (N_13798,N_12330,N_13027);
xor U13799 (N_13799,N_12869,N_13091);
and U13800 (N_13800,N_12875,N_12379);
or U13801 (N_13801,N_12811,N_12972);
or U13802 (N_13802,N_12398,N_13089);
nor U13803 (N_13803,N_12291,N_13178);
nand U13804 (N_13804,N_12089,N_13256);
and U13805 (N_13805,N_13001,N_13163);
nand U13806 (N_13806,N_12104,N_12836);
and U13807 (N_13807,N_13145,N_13167);
and U13808 (N_13808,N_13121,N_12874);
and U13809 (N_13809,N_12960,N_12235);
or U13810 (N_13810,N_12959,N_12579);
and U13811 (N_13811,N_12099,N_12746);
xor U13812 (N_13812,N_12225,N_13115);
nor U13813 (N_13813,N_13376,N_12833);
or U13814 (N_13814,N_12386,N_12909);
and U13815 (N_13815,N_12684,N_12322);
nand U13816 (N_13816,N_12263,N_12622);
xor U13817 (N_13817,N_13353,N_13065);
nand U13818 (N_13818,N_12635,N_12601);
or U13819 (N_13819,N_13438,N_12648);
nor U13820 (N_13820,N_13293,N_13125);
or U13821 (N_13821,N_12820,N_13122);
or U13822 (N_13822,N_13414,N_12209);
xor U13823 (N_13823,N_12630,N_12486);
or U13824 (N_13824,N_12662,N_12081);
or U13825 (N_13825,N_12356,N_12933);
and U13826 (N_13826,N_12981,N_12763);
nand U13827 (N_13827,N_12570,N_12665);
xnor U13828 (N_13828,N_12539,N_13156);
nor U13829 (N_13829,N_12865,N_13331);
nor U13830 (N_13830,N_12111,N_13020);
and U13831 (N_13831,N_12669,N_12946);
or U13832 (N_13832,N_13222,N_12405);
xor U13833 (N_13833,N_13117,N_13460);
and U13834 (N_13834,N_13343,N_12273);
nand U13835 (N_13835,N_12254,N_12160);
nand U13836 (N_13836,N_12719,N_12073);
xnor U13837 (N_13837,N_12548,N_12526);
and U13838 (N_13838,N_13295,N_13412);
nor U13839 (N_13839,N_12043,N_13181);
nand U13840 (N_13840,N_13441,N_13032);
nor U13841 (N_13841,N_12082,N_12321);
or U13842 (N_13842,N_12667,N_13214);
and U13843 (N_13843,N_13319,N_12664);
nor U13844 (N_13844,N_13284,N_12563);
or U13845 (N_13845,N_13084,N_12142);
xnor U13846 (N_13846,N_12229,N_12732);
or U13847 (N_13847,N_13270,N_13352);
xnor U13848 (N_13848,N_12006,N_12153);
and U13849 (N_13849,N_13488,N_13470);
and U13850 (N_13850,N_12144,N_13355);
or U13851 (N_13851,N_12255,N_12828);
and U13852 (N_13852,N_13096,N_12693);
or U13853 (N_13853,N_12067,N_12758);
or U13854 (N_13854,N_13277,N_12289);
and U13855 (N_13855,N_12002,N_13373);
xor U13856 (N_13856,N_12817,N_13479);
nor U13857 (N_13857,N_12720,N_12303);
or U13858 (N_13858,N_12965,N_12655);
or U13859 (N_13859,N_12218,N_13069);
nand U13860 (N_13860,N_12051,N_12896);
and U13861 (N_13861,N_12359,N_13230);
xor U13862 (N_13862,N_13229,N_12393);
and U13863 (N_13863,N_12776,N_13375);
nor U13864 (N_13864,N_12252,N_13486);
nor U13865 (N_13865,N_12425,N_12515);
nor U13866 (N_13866,N_12850,N_12256);
nand U13867 (N_13867,N_13428,N_12808);
or U13868 (N_13868,N_13262,N_13192);
nor U13869 (N_13869,N_12329,N_12904);
and U13870 (N_13870,N_12615,N_12365);
xnor U13871 (N_13871,N_12968,N_12283);
xor U13872 (N_13872,N_12204,N_13184);
xnor U13873 (N_13873,N_12424,N_13025);
nor U13874 (N_13874,N_13276,N_12574);
nand U13875 (N_13875,N_12829,N_13026);
nor U13876 (N_13876,N_13013,N_12059);
or U13877 (N_13877,N_12994,N_13119);
and U13878 (N_13878,N_12583,N_13330);
and U13879 (N_13879,N_12654,N_12703);
xnor U13880 (N_13880,N_13366,N_12126);
and U13881 (N_13881,N_13386,N_12165);
nand U13882 (N_13882,N_12020,N_12228);
nand U13883 (N_13883,N_13031,N_12550);
and U13884 (N_13884,N_12198,N_12401);
nor U13885 (N_13885,N_13074,N_13356);
or U13886 (N_13886,N_12340,N_12683);
or U13887 (N_13887,N_12288,N_13427);
nand U13888 (N_13888,N_12370,N_13142);
xnor U13889 (N_13889,N_12985,N_12809);
or U13890 (N_13890,N_12741,N_13401);
xnor U13891 (N_13891,N_13186,N_13472);
or U13892 (N_13892,N_12236,N_12318);
or U13893 (N_13893,N_12657,N_13063);
and U13894 (N_13894,N_13129,N_12511);
nand U13895 (N_13895,N_13340,N_12451);
and U13896 (N_13896,N_12033,N_12625);
or U13897 (N_13897,N_13388,N_12923);
nand U13898 (N_13898,N_13223,N_12163);
and U13899 (N_13899,N_13493,N_12775);
nand U13900 (N_13900,N_12488,N_12269);
and U13901 (N_13901,N_12672,N_12714);
nand U13902 (N_13902,N_13150,N_13209);
nor U13903 (N_13903,N_12088,N_12391);
nand U13904 (N_13904,N_13271,N_12513);
xor U13905 (N_13905,N_13413,N_12639);
xnor U13906 (N_13906,N_12005,N_12378);
and U13907 (N_13907,N_12925,N_12937);
or U13908 (N_13908,N_12095,N_12197);
or U13909 (N_13909,N_12131,N_12784);
or U13910 (N_13910,N_13411,N_12556);
and U13911 (N_13911,N_12813,N_12468);
nand U13912 (N_13912,N_12982,N_13465);
or U13913 (N_13913,N_13359,N_12912);
nor U13914 (N_13914,N_13086,N_12674);
or U13915 (N_13915,N_12132,N_12101);
nor U13916 (N_13916,N_12366,N_13457);
nor U13917 (N_13917,N_13109,N_12372);
nand U13918 (N_13918,N_12233,N_12007);
nor U13919 (N_13919,N_12781,N_12407);
nand U13920 (N_13920,N_12063,N_13453);
and U13921 (N_13921,N_13305,N_12397);
and U13922 (N_13922,N_12989,N_13019);
nand U13923 (N_13923,N_13481,N_13021);
or U13924 (N_13924,N_12807,N_13240);
xor U13925 (N_13925,N_13057,N_12343);
nor U13926 (N_13926,N_13492,N_12284);
nand U13927 (N_13927,N_13049,N_12750);
or U13928 (N_13928,N_12681,N_12096);
nand U13929 (N_13929,N_12480,N_12928);
xnor U13930 (N_13930,N_13051,N_13018);
and U13931 (N_13931,N_13105,N_12514);
and U13932 (N_13932,N_13144,N_13446);
or U13933 (N_13933,N_12125,N_13110);
nor U13934 (N_13934,N_13444,N_12328);
and U13935 (N_13935,N_12181,N_12508);
and U13936 (N_13936,N_12062,N_12309);
nand U13937 (N_13937,N_12814,N_12107);
or U13938 (N_13938,N_13101,N_13208);
or U13939 (N_13939,N_12961,N_12029);
nor U13940 (N_13940,N_13072,N_12839);
xnor U13941 (N_13941,N_13233,N_12678);
xor U13942 (N_13942,N_12631,N_13197);
nor U13943 (N_13943,N_13422,N_13462);
nor U13944 (N_13944,N_12337,N_13140);
xor U13945 (N_13945,N_13225,N_13374);
nand U13946 (N_13946,N_12990,N_12785);
nor U13947 (N_13947,N_12523,N_13046);
or U13948 (N_13948,N_13323,N_12573);
xor U13949 (N_13949,N_12154,N_12075);
nand U13950 (N_13950,N_12748,N_12866);
or U13951 (N_13951,N_12014,N_12294);
nand U13952 (N_13952,N_12203,N_13298);
or U13953 (N_13953,N_12647,N_12210);
nor U13954 (N_13954,N_12061,N_13174);
nor U13955 (N_13955,N_12860,N_12155);
nand U13956 (N_13956,N_12497,N_12482);
nor U13957 (N_13957,N_12368,N_13159);
nand U13958 (N_13958,N_12053,N_12474);
nor U13959 (N_13959,N_12250,N_13131);
nor U13960 (N_13960,N_12464,N_12048);
or U13961 (N_13961,N_13429,N_12835);
nor U13962 (N_13962,N_13468,N_13299);
nor U13963 (N_13963,N_12520,N_12352);
nand U13964 (N_13964,N_13487,N_12136);
xnor U13965 (N_13965,N_12301,N_12270);
and U13966 (N_13966,N_13339,N_12416);
nor U13967 (N_13967,N_12516,N_12145);
and U13968 (N_13968,N_12911,N_13342);
nand U13969 (N_13969,N_12637,N_13464);
and U13970 (N_13970,N_12092,N_12983);
nor U13971 (N_13971,N_12751,N_12885);
xnor U13972 (N_13972,N_13176,N_12016);
or U13973 (N_13973,N_13193,N_13194);
nor U13974 (N_13974,N_12692,N_13426);
or U13975 (N_13975,N_13354,N_12315);
nor U13976 (N_13976,N_13237,N_12710);
or U13977 (N_13977,N_12906,N_12873);
xnor U13978 (N_13978,N_12434,N_13351);
xor U13979 (N_13979,N_12432,N_13316);
or U13980 (N_13980,N_12832,N_13224);
nand U13981 (N_13981,N_12586,N_12844);
nand U13982 (N_13982,N_13321,N_13357);
nand U13983 (N_13983,N_13077,N_13153);
nand U13984 (N_13984,N_12277,N_12206);
xor U13985 (N_13985,N_13466,N_13362);
nand U13986 (N_13986,N_12518,N_13420);
nand U13987 (N_13987,N_12564,N_12500);
nand U13988 (N_13988,N_13094,N_12103);
nand U13989 (N_13989,N_12883,N_12712);
and U13990 (N_13990,N_13311,N_13201);
nand U13991 (N_13991,N_12608,N_12590);
nor U13992 (N_13992,N_12190,N_12588);
and U13993 (N_13993,N_13182,N_12760);
and U13994 (N_13994,N_12806,N_12487);
nor U13995 (N_13995,N_12979,N_12182);
nand U13996 (N_13996,N_13126,N_12898);
and U13997 (N_13997,N_12752,N_12932);
nand U13998 (N_13998,N_12593,N_12246);
and U13999 (N_13999,N_12704,N_12123);
nand U14000 (N_14000,N_12010,N_12792);
nand U14001 (N_14001,N_12903,N_13023);
and U14002 (N_14002,N_12930,N_13157);
or U14003 (N_14003,N_13216,N_12334);
nor U14004 (N_14004,N_12362,N_13034);
and U14005 (N_14005,N_12858,N_12158);
or U14006 (N_14006,N_12992,N_12695);
nor U14007 (N_14007,N_12771,N_13309);
nor U14008 (N_14008,N_12439,N_12467);
or U14009 (N_14009,N_13213,N_12717);
nand U14010 (N_14010,N_12355,N_13092);
or U14011 (N_14011,N_12108,N_12986);
or U14012 (N_14012,N_12037,N_13173);
and U14013 (N_14013,N_12677,N_12757);
and U14014 (N_14014,N_12024,N_12469);
and U14015 (N_14015,N_12217,N_13217);
nand U14016 (N_14016,N_12821,N_12036);
and U14017 (N_14017,N_13399,N_12410);
nor U14018 (N_14018,N_13480,N_12455);
nand U14019 (N_14019,N_13060,N_12849);
and U14020 (N_14020,N_12696,N_12354);
xnor U14021 (N_14021,N_12713,N_13442);
or U14022 (N_14022,N_12146,N_12734);
nand U14023 (N_14023,N_13402,N_12300);
or U14024 (N_14024,N_12079,N_12119);
xnor U14025 (N_14025,N_13036,N_12661);
and U14026 (N_14026,N_12594,N_12064);
or U14027 (N_14027,N_13434,N_12753);
nor U14028 (N_14028,N_13445,N_12939);
nor U14029 (N_14029,N_13044,N_12234);
xnor U14030 (N_14030,N_13002,N_13008);
xnor U14031 (N_14031,N_12533,N_12460);
nor U14032 (N_14032,N_12264,N_13431);
nor U14033 (N_14033,N_12087,N_12658);
nand U14034 (N_14034,N_12995,N_12316);
nor U14035 (N_14035,N_12422,N_13400);
or U14036 (N_14036,N_12172,N_12171);
xor U14037 (N_14037,N_12430,N_12841);
and U14038 (N_14038,N_12035,N_12640);
or U14039 (N_14039,N_12199,N_12816);
and U14040 (N_14040,N_12687,N_13418);
or U14041 (N_14041,N_12459,N_12634);
and U14042 (N_14042,N_12323,N_12031);
and U14043 (N_14043,N_12736,N_12041);
xnor U14044 (N_14044,N_12028,N_12058);
nor U14045 (N_14045,N_12074,N_12348);
or U14046 (N_14046,N_13103,N_12827);
and U14047 (N_14047,N_13381,N_12143);
nor U14048 (N_14048,N_12810,N_13232);
nand U14049 (N_14049,N_13061,N_12598);
or U14050 (N_14050,N_13241,N_12212);
xnor U14051 (N_14051,N_13459,N_12587);
xnor U14052 (N_14052,N_12705,N_12189);
or U14053 (N_14053,N_13064,N_12039);
xnor U14054 (N_14054,N_12466,N_12893);
and U14055 (N_14055,N_13029,N_12444);
nor U14056 (N_14056,N_13082,N_13006);
xnor U14057 (N_14057,N_12174,N_12842);
nor U14058 (N_14058,N_12116,N_13168);
nand U14059 (N_14059,N_12299,N_12364);
xor U14060 (N_14060,N_12722,N_13385);
and U14061 (N_14061,N_12232,N_12114);
nor U14062 (N_14062,N_12124,N_13384);
nand U14063 (N_14063,N_12544,N_12772);
nor U14064 (N_14064,N_13396,N_12013);
nand U14065 (N_14065,N_12977,N_12773);
or U14066 (N_14066,N_12954,N_12360);
and U14067 (N_14067,N_12834,N_13040);
xnor U14068 (N_14068,N_13169,N_12889);
xnor U14069 (N_14069,N_12437,N_13138);
or U14070 (N_14070,N_12402,N_12591);
nor U14071 (N_14071,N_12956,N_12901);
or U14072 (N_14072,N_13491,N_13154);
or U14073 (N_14073,N_12000,N_13274);
or U14074 (N_14074,N_13244,N_12066);
nor U14075 (N_14075,N_13475,N_12458);
nor U14076 (N_14076,N_12219,N_13076);
nand U14077 (N_14077,N_12052,N_12793);
or U14078 (N_14078,N_13041,N_12840);
and U14079 (N_14079,N_12754,N_12310);
nand U14080 (N_14080,N_12094,N_12743);
nand U14081 (N_14081,N_12764,N_13435);
nor U14082 (N_14082,N_12030,N_13452);
or U14083 (N_14083,N_13133,N_12226);
and U14084 (N_14084,N_12770,N_12022);
and U14085 (N_14085,N_12257,N_12237);
and U14086 (N_14086,N_13257,N_12306);
or U14087 (N_14087,N_13439,N_12958);
nor U14088 (N_14088,N_12509,N_13047);
and U14089 (N_14089,N_12524,N_12266);
and U14090 (N_14090,N_12602,N_12871);
nor U14091 (N_14091,N_12396,N_12457);
xor U14092 (N_14092,N_12701,N_12465);
nand U14093 (N_14093,N_12312,N_12148);
or U14094 (N_14094,N_12552,N_12927);
and U14095 (N_14095,N_12999,N_12049);
nor U14096 (N_14096,N_12998,N_13250);
nand U14097 (N_14097,N_12819,N_12213);
xor U14098 (N_14098,N_12435,N_12496);
and U14099 (N_14099,N_13383,N_13417);
nand U14100 (N_14100,N_12942,N_12803);
xnor U14101 (N_14101,N_12050,N_12097);
or U14102 (N_14102,N_13392,N_13387);
xor U14103 (N_14103,N_12545,N_12139);
nand U14104 (N_14104,N_12384,N_13327);
nor U14105 (N_14105,N_12227,N_13249);
xnor U14106 (N_14106,N_12413,N_13297);
and U14107 (N_14107,N_12975,N_13039);
or U14108 (N_14108,N_12978,N_13406);
and U14109 (N_14109,N_13139,N_12060);
or U14110 (N_14110,N_13317,N_13304);
nand U14111 (N_14111,N_12001,N_13463);
and U14112 (N_14112,N_12477,N_12626);
nand U14113 (N_14113,N_12537,N_12115);
xor U14114 (N_14114,N_12034,N_12870);
and U14115 (N_14115,N_13106,N_13253);
and U14116 (N_14116,N_13389,N_12449);
nand U14117 (N_14117,N_12499,N_12447);
and U14118 (N_14118,N_13279,N_12188);
and U14119 (N_14119,N_13363,N_12473);
nor U14120 (N_14120,N_12009,N_13264);
nor U14121 (N_14121,N_12403,N_12852);
or U14122 (N_14122,N_13242,N_13255);
or U14123 (N_14123,N_12275,N_12015);
and U14124 (N_14124,N_13005,N_12084);
nand U14125 (N_14125,N_12433,N_12156);
or U14126 (N_14126,N_12363,N_12971);
nor U14127 (N_14127,N_13070,N_12530);
or U14128 (N_14128,N_12812,N_13454);
and U14129 (N_14129,N_12580,N_13332);
and U14130 (N_14130,N_13054,N_13430);
nor U14131 (N_14131,N_12532,N_13143);
nor U14132 (N_14132,N_13267,N_12621);
or U14133 (N_14133,N_12744,N_13245);
or U14134 (N_14134,N_12025,N_12726);
nor U14135 (N_14135,N_12113,N_12996);
and U14136 (N_14136,N_13052,N_13170);
nor U14137 (N_14137,N_12395,N_12708);
and U14138 (N_14138,N_13361,N_13247);
nor U14139 (N_14139,N_12525,N_12851);
nand U14140 (N_14140,N_12542,N_12931);
or U14141 (N_14141,N_12756,N_13079);
nand U14142 (N_14142,N_13251,N_13151);
nor U14143 (N_14143,N_12653,N_13238);
xnor U14144 (N_14144,N_12443,N_12222);
nand U14145 (N_14145,N_13467,N_12253);
or U14146 (N_14146,N_13266,N_13325);
nand U14147 (N_14147,N_13484,N_12569);
nand U14148 (N_14148,N_12258,N_13189);
or U14149 (N_14149,N_12327,N_12728);
and U14150 (N_14150,N_12974,N_13263);
nor U14151 (N_14151,N_12794,N_12320);
xor U14152 (N_14152,N_12848,N_13292);
xor U14153 (N_14153,N_12394,N_12645);
nor U14154 (N_14154,N_12463,N_12489);
xor U14155 (N_14155,N_12837,N_12973);
and U14156 (N_14156,N_12945,N_13015);
and U14157 (N_14157,N_12910,N_13100);
or U14158 (N_14158,N_12623,N_13336);
xor U14159 (N_14159,N_12578,N_13179);
nor U14160 (N_14160,N_12038,N_12675);
and U14161 (N_14161,N_13410,N_13349);
nor U14162 (N_14162,N_12729,N_12506);
xor U14163 (N_14163,N_13489,N_13403);
nand U14164 (N_14164,N_13068,N_12795);
and U14165 (N_14165,N_12605,N_12390);
or U14166 (N_14166,N_12825,N_12241);
xor U14167 (N_14167,N_12265,N_12191);
nor U14168 (N_14168,N_13372,N_12613);
nand U14169 (N_14169,N_13369,N_12201);
and U14170 (N_14170,N_12774,N_13059);
xnor U14171 (N_14171,N_12926,N_12231);
xnor U14172 (N_14172,N_13328,N_12798);
and U14173 (N_14173,N_12331,N_12003);
nand U14174 (N_14174,N_12083,N_12559);
xor U14175 (N_14175,N_13338,N_12843);
nand U14176 (N_14176,N_12409,N_12472);
xor U14177 (N_14177,N_12381,N_13450);
and U14178 (N_14178,N_12260,N_12475);
or U14179 (N_14179,N_13393,N_12071);
and U14180 (N_14180,N_12976,N_12585);
nor U14181 (N_14181,N_12922,N_12211);
or U14182 (N_14182,N_12846,N_13290);
and U14183 (N_14183,N_13038,N_12091);
or U14184 (N_14184,N_12727,N_12993);
xnor U14185 (N_14185,N_12884,N_12963);
nor U14186 (N_14186,N_12415,N_12392);
xor U14187 (N_14187,N_12891,N_12759);
or U14188 (N_14188,N_12389,N_12220);
nor U14189 (N_14189,N_13188,N_12886);
xor U14190 (N_14190,N_12510,N_12317);
nor U14191 (N_14191,N_13448,N_12685);
nor U14192 (N_14192,N_12991,N_12818);
xor U14193 (N_14193,N_12261,N_12495);
nor U14194 (N_14194,N_12796,N_12251);
or U14195 (N_14195,N_12799,N_12855);
nand U14196 (N_14196,N_13333,N_13221);
xnor U14197 (N_14197,N_13095,N_12652);
nor U14198 (N_14198,N_12023,N_12824);
xnor U14199 (N_14199,N_13476,N_13114);
nor U14200 (N_14200,N_13111,N_13469);
nor U14201 (N_14201,N_12880,N_12274);
nand U14202 (N_14202,N_12021,N_12333);
nand U14203 (N_14203,N_12680,N_12673);
and U14204 (N_14204,N_12461,N_12892);
or U14205 (N_14205,N_12112,N_13346);
nor U14206 (N_14206,N_12789,N_13011);
or U14207 (N_14207,N_12944,N_13497);
nor U14208 (N_14208,N_12345,N_12344);
xor U14209 (N_14209,N_13172,N_13087);
or U14210 (N_14210,N_13259,N_12581);
or U14211 (N_14211,N_12151,N_12742);
nor U14212 (N_14212,N_13206,N_13199);
nor U14213 (N_14213,N_12426,N_12120);
nor U14214 (N_14214,N_12221,N_12917);
nand U14215 (N_14215,N_12857,N_13449);
and U14216 (N_14216,N_13081,N_12377);
nor U14217 (N_14217,N_12668,N_13112);
xor U14218 (N_14218,N_13183,N_12448);
and U14219 (N_14219,N_12137,N_13280);
nand U14220 (N_14220,N_13149,N_12339);
and U14221 (N_14221,N_13313,N_12302);
or U14222 (N_14222,N_12399,N_13477);
nor U14223 (N_14223,N_13171,N_13310);
xnor U14224 (N_14224,N_12054,N_13175);
or U14225 (N_14225,N_13301,N_13368);
nor U14226 (N_14226,N_12815,N_12612);
nor U14227 (N_14227,N_12914,N_12361);
nor U14228 (N_14228,N_12346,N_12543);
and U14229 (N_14229,N_13158,N_12276);
nand U14230 (N_14230,N_12247,N_13482);
nand U14231 (N_14231,N_12184,N_13017);
nand U14232 (N_14232,N_13409,N_12907);
xor U14233 (N_14233,N_12239,N_12441);
or U14234 (N_14234,N_13066,N_12476);
nor U14235 (N_14235,N_12431,N_12152);
xnor U14236 (N_14236,N_12004,N_12881);
or U14237 (N_14237,N_13268,N_12427);
nor U14238 (N_14238,N_12373,N_12529);
and U14239 (N_14239,N_12406,N_12314);
nand U14240 (N_14240,N_12735,N_12888);
or U14241 (N_14241,N_12121,N_12876);
nand U14242 (N_14242,N_12546,N_13200);
xor U14243 (N_14243,N_12575,N_13162);
xnor U14244 (N_14244,N_12157,N_12853);
and U14245 (N_14245,N_12606,N_12788);
or U14246 (N_14246,N_12272,N_12388);
or U14247 (N_14247,N_12290,N_12790);
or U14248 (N_14248,N_12106,N_12787);
nor U14249 (N_14249,N_12970,N_13099);
xor U14250 (N_14250,N_12007,N_13092);
and U14251 (N_14251,N_13151,N_12610);
xnor U14252 (N_14252,N_12587,N_13070);
nand U14253 (N_14253,N_12429,N_13181);
and U14254 (N_14254,N_13446,N_12811);
nand U14255 (N_14255,N_12762,N_12502);
and U14256 (N_14256,N_12913,N_13018);
nor U14257 (N_14257,N_13080,N_12482);
or U14258 (N_14258,N_12380,N_13270);
or U14259 (N_14259,N_12780,N_12265);
and U14260 (N_14260,N_12984,N_13285);
xor U14261 (N_14261,N_12790,N_13106);
xor U14262 (N_14262,N_13479,N_13421);
or U14263 (N_14263,N_13301,N_13460);
and U14264 (N_14264,N_12262,N_12507);
and U14265 (N_14265,N_13099,N_12935);
xor U14266 (N_14266,N_12724,N_12211);
or U14267 (N_14267,N_12433,N_12752);
or U14268 (N_14268,N_12624,N_12693);
and U14269 (N_14269,N_12608,N_12635);
or U14270 (N_14270,N_13221,N_12916);
nor U14271 (N_14271,N_12472,N_12852);
nand U14272 (N_14272,N_12406,N_12232);
or U14273 (N_14273,N_12223,N_13123);
and U14274 (N_14274,N_12203,N_13308);
nand U14275 (N_14275,N_13093,N_12491);
nand U14276 (N_14276,N_12040,N_12942);
and U14277 (N_14277,N_12657,N_12599);
nand U14278 (N_14278,N_13305,N_12432);
xor U14279 (N_14279,N_12546,N_12694);
nand U14280 (N_14280,N_13498,N_12744);
xor U14281 (N_14281,N_13315,N_12116);
nor U14282 (N_14282,N_12187,N_12344);
or U14283 (N_14283,N_12685,N_12400);
nand U14284 (N_14284,N_13094,N_13304);
or U14285 (N_14285,N_13321,N_13290);
and U14286 (N_14286,N_13339,N_12079);
nand U14287 (N_14287,N_12917,N_12023);
nand U14288 (N_14288,N_12184,N_12710);
and U14289 (N_14289,N_12665,N_12559);
and U14290 (N_14290,N_12816,N_12838);
and U14291 (N_14291,N_12608,N_12704);
nand U14292 (N_14292,N_13450,N_13112);
and U14293 (N_14293,N_13368,N_13001);
or U14294 (N_14294,N_13239,N_13333);
or U14295 (N_14295,N_13157,N_12695);
nor U14296 (N_14296,N_12883,N_13116);
xor U14297 (N_14297,N_12321,N_12489);
xor U14298 (N_14298,N_12131,N_12065);
and U14299 (N_14299,N_12730,N_12785);
nor U14300 (N_14300,N_13269,N_12046);
nand U14301 (N_14301,N_12851,N_12437);
and U14302 (N_14302,N_13395,N_12158);
or U14303 (N_14303,N_13390,N_13171);
and U14304 (N_14304,N_12684,N_12797);
xnor U14305 (N_14305,N_13044,N_12008);
nor U14306 (N_14306,N_12681,N_12419);
or U14307 (N_14307,N_12812,N_12078);
xor U14308 (N_14308,N_12488,N_13148);
or U14309 (N_14309,N_13358,N_13031);
nand U14310 (N_14310,N_12134,N_13155);
nor U14311 (N_14311,N_12786,N_13031);
or U14312 (N_14312,N_12786,N_13298);
nor U14313 (N_14313,N_13375,N_12694);
nor U14314 (N_14314,N_12563,N_12823);
or U14315 (N_14315,N_13190,N_12956);
or U14316 (N_14316,N_12569,N_13382);
nor U14317 (N_14317,N_12072,N_12645);
and U14318 (N_14318,N_12886,N_12491);
xor U14319 (N_14319,N_12673,N_12993);
nand U14320 (N_14320,N_12776,N_12198);
or U14321 (N_14321,N_13061,N_13417);
or U14322 (N_14322,N_12834,N_13105);
and U14323 (N_14323,N_12491,N_13298);
nand U14324 (N_14324,N_12920,N_12248);
and U14325 (N_14325,N_13345,N_13270);
xor U14326 (N_14326,N_12688,N_13218);
nand U14327 (N_14327,N_12339,N_12956);
and U14328 (N_14328,N_13434,N_13472);
and U14329 (N_14329,N_12396,N_12517);
or U14330 (N_14330,N_12850,N_12135);
nor U14331 (N_14331,N_12215,N_12300);
nor U14332 (N_14332,N_13467,N_13206);
xnor U14333 (N_14333,N_12556,N_13463);
xnor U14334 (N_14334,N_12250,N_12848);
nor U14335 (N_14335,N_12778,N_12482);
nor U14336 (N_14336,N_13187,N_12312);
xor U14337 (N_14337,N_13161,N_13113);
and U14338 (N_14338,N_12508,N_12025);
xor U14339 (N_14339,N_13375,N_12999);
nand U14340 (N_14340,N_12056,N_12577);
and U14341 (N_14341,N_12334,N_12081);
nor U14342 (N_14342,N_12615,N_12716);
nand U14343 (N_14343,N_13013,N_12492);
and U14344 (N_14344,N_12930,N_13438);
or U14345 (N_14345,N_12476,N_12488);
nand U14346 (N_14346,N_12844,N_12233);
and U14347 (N_14347,N_12001,N_12416);
or U14348 (N_14348,N_13240,N_13448);
or U14349 (N_14349,N_13117,N_12619);
and U14350 (N_14350,N_13484,N_12893);
nor U14351 (N_14351,N_13456,N_12732);
or U14352 (N_14352,N_12060,N_12002);
nand U14353 (N_14353,N_13075,N_13426);
xnor U14354 (N_14354,N_12897,N_12094);
nand U14355 (N_14355,N_13333,N_13404);
nand U14356 (N_14356,N_13455,N_12704);
or U14357 (N_14357,N_12156,N_12843);
xor U14358 (N_14358,N_12915,N_12894);
nand U14359 (N_14359,N_12326,N_12429);
or U14360 (N_14360,N_12954,N_12811);
nand U14361 (N_14361,N_12361,N_12593);
nand U14362 (N_14362,N_12852,N_12903);
nand U14363 (N_14363,N_12973,N_13196);
nand U14364 (N_14364,N_13334,N_12945);
or U14365 (N_14365,N_12318,N_13030);
nand U14366 (N_14366,N_12362,N_12676);
nor U14367 (N_14367,N_13222,N_12687);
nand U14368 (N_14368,N_12130,N_12651);
nor U14369 (N_14369,N_12324,N_12403);
nor U14370 (N_14370,N_13127,N_13049);
xor U14371 (N_14371,N_12410,N_12450);
and U14372 (N_14372,N_12164,N_12297);
and U14373 (N_14373,N_13041,N_13496);
nor U14374 (N_14374,N_12964,N_12474);
and U14375 (N_14375,N_13038,N_13226);
or U14376 (N_14376,N_13417,N_12641);
or U14377 (N_14377,N_13440,N_12071);
xor U14378 (N_14378,N_12352,N_12539);
nand U14379 (N_14379,N_13368,N_13372);
nand U14380 (N_14380,N_12536,N_12514);
or U14381 (N_14381,N_12615,N_12717);
and U14382 (N_14382,N_13411,N_12460);
or U14383 (N_14383,N_13393,N_12545);
nor U14384 (N_14384,N_12141,N_12723);
nand U14385 (N_14385,N_12107,N_12323);
nand U14386 (N_14386,N_13075,N_13143);
xnor U14387 (N_14387,N_12522,N_12770);
nor U14388 (N_14388,N_13031,N_12905);
nor U14389 (N_14389,N_12533,N_13220);
xor U14390 (N_14390,N_12236,N_12502);
and U14391 (N_14391,N_12067,N_13103);
or U14392 (N_14392,N_13411,N_13050);
xor U14393 (N_14393,N_13345,N_12228);
nor U14394 (N_14394,N_13375,N_12843);
nand U14395 (N_14395,N_12716,N_13463);
nor U14396 (N_14396,N_12759,N_12525);
or U14397 (N_14397,N_13469,N_13150);
nor U14398 (N_14398,N_12971,N_13107);
or U14399 (N_14399,N_13123,N_12859);
nand U14400 (N_14400,N_12922,N_12652);
nor U14401 (N_14401,N_12151,N_12497);
and U14402 (N_14402,N_12859,N_13424);
nor U14403 (N_14403,N_12060,N_12228);
and U14404 (N_14404,N_12131,N_12600);
xor U14405 (N_14405,N_12830,N_12268);
or U14406 (N_14406,N_12719,N_13309);
and U14407 (N_14407,N_12122,N_13207);
nand U14408 (N_14408,N_13168,N_12250);
and U14409 (N_14409,N_13088,N_12410);
and U14410 (N_14410,N_13415,N_12491);
xor U14411 (N_14411,N_13226,N_13341);
nor U14412 (N_14412,N_13495,N_12567);
xor U14413 (N_14413,N_12078,N_12686);
or U14414 (N_14414,N_12417,N_13212);
and U14415 (N_14415,N_12244,N_13069);
nand U14416 (N_14416,N_13285,N_12552);
nor U14417 (N_14417,N_12168,N_12079);
xnor U14418 (N_14418,N_13009,N_12954);
nor U14419 (N_14419,N_12827,N_12526);
or U14420 (N_14420,N_12514,N_12634);
or U14421 (N_14421,N_12483,N_13310);
nor U14422 (N_14422,N_13473,N_13145);
nand U14423 (N_14423,N_12113,N_13057);
nand U14424 (N_14424,N_12235,N_12349);
and U14425 (N_14425,N_12548,N_13411);
xnor U14426 (N_14426,N_12745,N_13291);
and U14427 (N_14427,N_13163,N_12266);
nor U14428 (N_14428,N_13189,N_12738);
and U14429 (N_14429,N_12927,N_13358);
xor U14430 (N_14430,N_12469,N_13413);
or U14431 (N_14431,N_12750,N_13032);
and U14432 (N_14432,N_13226,N_12414);
nand U14433 (N_14433,N_12462,N_12211);
nor U14434 (N_14434,N_12118,N_12787);
xor U14435 (N_14435,N_12504,N_12107);
or U14436 (N_14436,N_12802,N_13087);
xor U14437 (N_14437,N_12343,N_13048);
and U14438 (N_14438,N_13207,N_12182);
nand U14439 (N_14439,N_12997,N_12755);
nand U14440 (N_14440,N_12492,N_12315);
or U14441 (N_14441,N_12772,N_13074);
xor U14442 (N_14442,N_12753,N_12716);
and U14443 (N_14443,N_13005,N_13367);
and U14444 (N_14444,N_13213,N_12263);
nand U14445 (N_14445,N_12827,N_13005);
and U14446 (N_14446,N_12088,N_13349);
xor U14447 (N_14447,N_12659,N_12120);
or U14448 (N_14448,N_12851,N_13094);
nand U14449 (N_14449,N_12378,N_12754);
nand U14450 (N_14450,N_13170,N_12137);
xor U14451 (N_14451,N_13342,N_12410);
nand U14452 (N_14452,N_12324,N_13419);
or U14453 (N_14453,N_13299,N_12771);
nand U14454 (N_14454,N_12552,N_12349);
nand U14455 (N_14455,N_12080,N_12310);
nor U14456 (N_14456,N_13092,N_13495);
xnor U14457 (N_14457,N_12931,N_13386);
xor U14458 (N_14458,N_12398,N_13022);
and U14459 (N_14459,N_12541,N_13246);
and U14460 (N_14460,N_12046,N_13197);
nand U14461 (N_14461,N_12652,N_12360);
and U14462 (N_14462,N_13471,N_12954);
nand U14463 (N_14463,N_12680,N_13229);
or U14464 (N_14464,N_12436,N_12121);
and U14465 (N_14465,N_13062,N_13495);
nand U14466 (N_14466,N_12452,N_13048);
or U14467 (N_14467,N_12454,N_12370);
nand U14468 (N_14468,N_12427,N_12991);
xnor U14469 (N_14469,N_12638,N_12475);
xnor U14470 (N_14470,N_13411,N_12440);
and U14471 (N_14471,N_12975,N_12033);
xnor U14472 (N_14472,N_13444,N_12879);
nor U14473 (N_14473,N_12263,N_13287);
nor U14474 (N_14474,N_13231,N_12331);
xnor U14475 (N_14475,N_13345,N_12141);
and U14476 (N_14476,N_12556,N_12829);
and U14477 (N_14477,N_13168,N_13146);
nor U14478 (N_14478,N_12860,N_12923);
nand U14479 (N_14479,N_12225,N_13150);
or U14480 (N_14480,N_12122,N_13158);
and U14481 (N_14481,N_12954,N_12355);
xnor U14482 (N_14482,N_12324,N_13402);
and U14483 (N_14483,N_13005,N_12166);
and U14484 (N_14484,N_12808,N_13171);
or U14485 (N_14485,N_12979,N_12545);
or U14486 (N_14486,N_13053,N_12673);
nand U14487 (N_14487,N_12553,N_12939);
xnor U14488 (N_14488,N_13319,N_13455);
nor U14489 (N_14489,N_12091,N_13087);
xor U14490 (N_14490,N_13278,N_12272);
and U14491 (N_14491,N_13366,N_13223);
nand U14492 (N_14492,N_13231,N_13154);
nand U14493 (N_14493,N_12729,N_12745);
and U14494 (N_14494,N_13362,N_13230);
and U14495 (N_14495,N_13101,N_12463);
nand U14496 (N_14496,N_12252,N_12344);
and U14497 (N_14497,N_13111,N_12188);
nand U14498 (N_14498,N_13329,N_12554);
or U14499 (N_14499,N_12564,N_13072);
nand U14500 (N_14500,N_13076,N_12099);
xnor U14501 (N_14501,N_12661,N_12069);
or U14502 (N_14502,N_12374,N_13207);
or U14503 (N_14503,N_12977,N_13250);
xor U14504 (N_14504,N_12877,N_12412);
and U14505 (N_14505,N_13324,N_12407);
nand U14506 (N_14506,N_13027,N_12547);
xnor U14507 (N_14507,N_12984,N_12927);
xnor U14508 (N_14508,N_13198,N_12851);
or U14509 (N_14509,N_12071,N_12554);
and U14510 (N_14510,N_12392,N_13178);
nor U14511 (N_14511,N_12052,N_13289);
and U14512 (N_14512,N_13210,N_12557);
xnor U14513 (N_14513,N_12860,N_12897);
xnor U14514 (N_14514,N_12567,N_12478);
nand U14515 (N_14515,N_12674,N_12929);
nor U14516 (N_14516,N_13186,N_12836);
xor U14517 (N_14517,N_12101,N_12966);
nand U14518 (N_14518,N_12191,N_13433);
nand U14519 (N_14519,N_12586,N_13332);
xor U14520 (N_14520,N_13268,N_13128);
nor U14521 (N_14521,N_12699,N_13409);
xor U14522 (N_14522,N_12089,N_12275);
nand U14523 (N_14523,N_12531,N_12461);
nor U14524 (N_14524,N_13281,N_12360);
xnor U14525 (N_14525,N_12554,N_12083);
nand U14526 (N_14526,N_13319,N_13422);
nand U14527 (N_14527,N_12692,N_12110);
or U14528 (N_14528,N_12307,N_13289);
and U14529 (N_14529,N_13133,N_12959);
or U14530 (N_14530,N_12603,N_12247);
nor U14531 (N_14531,N_13472,N_13369);
and U14532 (N_14532,N_13051,N_12537);
nor U14533 (N_14533,N_12950,N_12687);
and U14534 (N_14534,N_12067,N_12060);
and U14535 (N_14535,N_13215,N_12826);
nand U14536 (N_14536,N_12108,N_12029);
nor U14537 (N_14537,N_12028,N_12083);
and U14538 (N_14538,N_12162,N_12715);
xor U14539 (N_14539,N_12882,N_12169);
nor U14540 (N_14540,N_13278,N_13017);
and U14541 (N_14541,N_12438,N_12326);
xnor U14542 (N_14542,N_13013,N_13134);
xor U14543 (N_14543,N_12774,N_12881);
or U14544 (N_14544,N_12624,N_12126);
nand U14545 (N_14545,N_12313,N_12684);
or U14546 (N_14546,N_12583,N_12626);
and U14547 (N_14547,N_12879,N_12218);
or U14548 (N_14548,N_12499,N_12109);
and U14549 (N_14549,N_12035,N_12705);
and U14550 (N_14550,N_12111,N_13171);
nand U14551 (N_14551,N_12379,N_12258);
xor U14552 (N_14552,N_13178,N_12771);
xor U14553 (N_14553,N_12242,N_12845);
or U14554 (N_14554,N_13053,N_13241);
and U14555 (N_14555,N_12369,N_12097);
or U14556 (N_14556,N_12061,N_13358);
or U14557 (N_14557,N_13456,N_12000);
and U14558 (N_14558,N_12079,N_12012);
and U14559 (N_14559,N_12166,N_13055);
xnor U14560 (N_14560,N_12868,N_12693);
or U14561 (N_14561,N_12891,N_12651);
and U14562 (N_14562,N_12132,N_12472);
nor U14563 (N_14563,N_13445,N_12550);
nand U14564 (N_14564,N_13116,N_13133);
or U14565 (N_14565,N_12573,N_12077);
and U14566 (N_14566,N_12245,N_12862);
xor U14567 (N_14567,N_12648,N_13071);
xor U14568 (N_14568,N_13335,N_12340);
or U14569 (N_14569,N_13021,N_12261);
nand U14570 (N_14570,N_12067,N_12439);
xnor U14571 (N_14571,N_13014,N_12636);
or U14572 (N_14572,N_13383,N_13187);
xnor U14573 (N_14573,N_12291,N_12096);
nand U14574 (N_14574,N_13478,N_12387);
nand U14575 (N_14575,N_12127,N_12895);
or U14576 (N_14576,N_12326,N_12996);
and U14577 (N_14577,N_12596,N_12377);
or U14578 (N_14578,N_12212,N_13300);
xnor U14579 (N_14579,N_12687,N_12604);
and U14580 (N_14580,N_13316,N_13288);
nor U14581 (N_14581,N_12595,N_12777);
xnor U14582 (N_14582,N_12048,N_13273);
and U14583 (N_14583,N_13168,N_12897);
or U14584 (N_14584,N_12764,N_12224);
xnor U14585 (N_14585,N_12741,N_12446);
and U14586 (N_14586,N_13467,N_13068);
or U14587 (N_14587,N_13268,N_12832);
nand U14588 (N_14588,N_12833,N_12098);
nor U14589 (N_14589,N_13275,N_12409);
nand U14590 (N_14590,N_12294,N_13476);
nand U14591 (N_14591,N_12177,N_12638);
xor U14592 (N_14592,N_12625,N_12814);
nor U14593 (N_14593,N_13431,N_12017);
nand U14594 (N_14594,N_12643,N_12233);
nor U14595 (N_14595,N_13303,N_12051);
and U14596 (N_14596,N_13049,N_12513);
and U14597 (N_14597,N_12108,N_12965);
and U14598 (N_14598,N_12863,N_13179);
or U14599 (N_14599,N_13164,N_13341);
and U14600 (N_14600,N_12174,N_12990);
or U14601 (N_14601,N_12445,N_12483);
nand U14602 (N_14602,N_12934,N_12874);
or U14603 (N_14603,N_13132,N_12927);
or U14604 (N_14604,N_12170,N_12273);
or U14605 (N_14605,N_12292,N_13448);
and U14606 (N_14606,N_13488,N_12652);
xor U14607 (N_14607,N_12948,N_12467);
or U14608 (N_14608,N_12146,N_13303);
xnor U14609 (N_14609,N_12000,N_12178);
and U14610 (N_14610,N_12339,N_12530);
nand U14611 (N_14611,N_13295,N_12943);
nand U14612 (N_14612,N_12396,N_12536);
nor U14613 (N_14613,N_12400,N_12307);
and U14614 (N_14614,N_13056,N_12356);
xnor U14615 (N_14615,N_12998,N_12802);
nor U14616 (N_14616,N_12179,N_12646);
nand U14617 (N_14617,N_12008,N_12369);
nand U14618 (N_14618,N_12682,N_13013);
xor U14619 (N_14619,N_13300,N_12871);
nor U14620 (N_14620,N_12274,N_13214);
or U14621 (N_14621,N_13379,N_12723);
and U14622 (N_14622,N_13214,N_12158);
or U14623 (N_14623,N_12631,N_12214);
or U14624 (N_14624,N_13211,N_13375);
nor U14625 (N_14625,N_12804,N_12999);
xor U14626 (N_14626,N_12896,N_12401);
and U14627 (N_14627,N_12485,N_12951);
nor U14628 (N_14628,N_12728,N_12078);
and U14629 (N_14629,N_13352,N_13038);
xor U14630 (N_14630,N_13113,N_13175);
nor U14631 (N_14631,N_12753,N_12193);
or U14632 (N_14632,N_13440,N_12655);
xor U14633 (N_14633,N_12004,N_13155);
or U14634 (N_14634,N_12292,N_13368);
xnor U14635 (N_14635,N_12223,N_12704);
and U14636 (N_14636,N_12471,N_12263);
and U14637 (N_14637,N_12242,N_13110);
xor U14638 (N_14638,N_12722,N_12818);
nand U14639 (N_14639,N_12602,N_12414);
nand U14640 (N_14640,N_12986,N_12001);
nand U14641 (N_14641,N_12574,N_12024);
xor U14642 (N_14642,N_12863,N_12389);
and U14643 (N_14643,N_13437,N_12916);
nand U14644 (N_14644,N_12825,N_12295);
nand U14645 (N_14645,N_13416,N_12711);
nor U14646 (N_14646,N_12895,N_13444);
nand U14647 (N_14647,N_12414,N_12556);
and U14648 (N_14648,N_12120,N_13487);
xnor U14649 (N_14649,N_13081,N_12893);
xnor U14650 (N_14650,N_12650,N_12427);
and U14651 (N_14651,N_12608,N_12293);
and U14652 (N_14652,N_12657,N_12010);
nor U14653 (N_14653,N_12681,N_12218);
or U14654 (N_14654,N_12608,N_12224);
or U14655 (N_14655,N_12961,N_13361);
xnor U14656 (N_14656,N_12031,N_13147);
nor U14657 (N_14657,N_12938,N_12816);
xor U14658 (N_14658,N_13452,N_13401);
xnor U14659 (N_14659,N_12655,N_13413);
nand U14660 (N_14660,N_13474,N_12603);
xnor U14661 (N_14661,N_12049,N_12842);
xor U14662 (N_14662,N_13035,N_12801);
xor U14663 (N_14663,N_12456,N_12276);
nand U14664 (N_14664,N_13471,N_13033);
nand U14665 (N_14665,N_12127,N_12355);
nor U14666 (N_14666,N_12883,N_13434);
or U14667 (N_14667,N_12383,N_12789);
nand U14668 (N_14668,N_12016,N_12064);
and U14669 (N_14669,N_13476,N_12826);
xor U14670 (N_14670,N_12478,N_12972);
xor U14671 (N_14671,N_13202,N_12220);
nand U14672 (N_14672,N_13458,N_12465);
nand U14673 (N_14673,N_12037,N_13412);
nor U14674 (N_14674,N_12709,N_12865);
nor U14675 (N_14675,N_12064,N_13134);
nand U14676 (N_14676,N_12352,N_12005);
or U14677 (N_14677,N_12800,N_13159);
and U14678 (N_14678,N_12307,N_12843);
and U14679 (N_14679,N_12758,N_13123);
nor U14680 (N_14680,N_13382,N_12231);
nor U14681 (N_14681,N_12020,N_12892);
nand U14682 (N_14682,N_13246,N_13059);
and U14683 (N_14683,N_12657,N_12481);
and U14684 (N_14684,N_12718,N_12827);
nor U14685 (N_14685,N_13352,N_13264);
and U14686 (N_14686,N_12831,N_12676);
and U14687 (N_14687,N_13242,N_12214);
xnor U14688 (N_14688,N_13365,N_12166);
nand U14689 (N_14689,N_13461,N_12541);
or U14690 (N_14690,N_13211,N_12392);
or U14691 (N_14691,N_12974,N_13296);
xor U14692 (N_14692,N_12126,N_13071);
and U14693 (N_14693,N_12020,N_13403);
and U14694 (N_14694,N_12022,N_12873);
or U14695 (N_14695,N_12094,N_12562);
xor U14696 (N_14696,N_12587,N_13083);
xor U14697 (N_14697,N_13033,N_12576);
nor U14698 (N_14698,N_12865,N_13489);
nor U14699 (N_14699,N_13481,N_12278);
nand U14700 (N_14700,N_13233,N_12287);
nor U14701 (N_14701,N_12309,N_12291);
nand U14702 (N_14702,N_12445,N_12844);
and U14703 (N_14703,N_12876,N_12930);
or U14704 (N_14704,N_12965,N_12157);
nor U14705 (N_14705,N_13071,N_12307);
nand U14706 (N_14706,N_12077,N_13287);
or U14707 (N_14707,N_12864,N_12266);
nand U14708 (N_14708,N_13393,N_12078);
or U14709 (N_14709,N_12629,N_12717);
and U14710 (N_14710,N_13089,N_12219);
and U14711 (N_14711,N_12247,N_12688);
or U14712 (N_14712,N_12873,N_13219);
nand U14713 (N_14713,N_12367,N_13162);
or U14714 (N_14714,N_13213,N_12855);
nor U14715 (N_14715,N_12418,N_13285);
nor U14716 (N_14716,N_12371,N_13232);
or U14717 (N_14717,N_12344,N_12729);
and U14718 (N_14718,N_12574,N_12321);
xnor U14719 (N_14719,N_13063,N_13004);
nor U14720 (N_14720,N_12451,N_12608);
nor U14721 (N_14721,N_12384,N_12023);
nor U14722 (N_14722,N_12849,N_12192);
nor U14723 (N_14723,N_12604,N_12823);
xnor U14724 (N_14724,N_12225,N_12739);
nand U14725 (N_14725,N_12814,N_12669);
xor U14726 (N_14726,N_12378,N_13329);
and U14727 (N_14727,N_13166,N_12837);
xor U14728 (N_14728,N_12078,N_12560);
xor U14729 (N_14729,N_13229,N_12047);
nor U14730 (N_14730,N_12305,N_12310);
xor U14731 (N_14731,N_13170,N_12775);
nand U14732 (N_14732,N_13458,N_12474);
and U14733 (N_14733,N_12272,N_12561);
nand U14734 (N_14734,N_12487,N_13018);
or U14735 (N_14735,N_12854,N_13288);
xor U14736 (N_14736,N_12688,N_12099);
xnor U14737 (N_14737,N_12122,N_12924);
nor U14738 (N_14738,N_12408,N_12377);
xnor U14739 (N_14739,N_13318,N_13073);
and U14740 (N_14740,N_13252,N_13226);
nor U14741 (N_14741,N_12561,N_12681);
or U14742 (N_14742,N_12337,N_12572);
xnor U14743 (N_14743,N_13150,N_13276);
xnor U14744 (N_14744,N_12362,N_12364);
nor U14745 (N_14745,N_13286,N_12536);
and U14746 (N_14746,N_12428,N_12165);
xor U14747 (N_14747,N_12757,N_12220);
and U14748 (N_14748,N_12589,N_13245);
xor U14749 (N_14749,N_12149,N_12830);
nor U14750 (N_14750,N_13039,N_12464);
nor U14751 (N_14751,N_12521,N_12915);
and U14752 (N_14752,N_12662,N_12313);
and U14753 (N_14753,N_12899,N_12382);
and U14754 (N_14754,N_12624,N_12277);
nand U14755 (N_14755,N_13475,N_12706);
xnor U14756 (N_14756,N_12546,N_12927);
and U14757 (N_14757,N_13250,N_12186);
or U14758 (N_14758,N_12961,N_12204);
or U14759 (N_14759,N_12983,N_13451);
or U14760 (N_14760,N_12684,N_12038);
xor U14761 (N_14761,N_13288,N_12188);
nor U14762 (N_14762,N_13352,N_12807);
and U14763 (N_14763,N_12379,N_12309);
xor U14764 (N_14764,N_13482,N_13012);
nor U14765 (N_14765,N_12721,N_13073);
nor U14766 (N_14766,N_12835,N_12744);
nor U14767 (N_14767,N_12242,N_13082);
nor U14768 (N_14768,N_13364,N_13058);
nand U14769 (N_14769,N_12046,N_12707);
or U14770 (N_14770,N_12563,N_12714);
nor U14771 (N_14771,N_12340,N_12465);
nand U14772 (N_14772,N_12636,N_12381);
nand U14773 (N_14773,N_12631,N_12177);
nor U14774 (N_14774,N_12972,N_12503);
xnor U14775 (N_14775,N_12477,N_12354);
nand U14776 (N_14776,N_12946,N_13119);
or U14777 (N_14777,N_12014,N_12278);
or U14778 (N_14778,N_12362,N_12918);
and U14779 (N_14779,N_12464,N_12813);
or U14780 (N_14780,N_12319,N_12280);
nor U14781 (N_14781,N_12529,N_13073);
xnor U14782 (N_14782,N_12026,N_12045);
nand U14783 (N_14783,N_12153,N_13305);
or U14784 (N_14784,N_12025,N_13359);
nand U14785 (N_14785,N_13056,N_13239);
or U14786 (N_14786,N_12964,N_13286);
xnor U14787 (N_14787,N_12956,N_13175);
and U14788 (N_14788,N_12662,N_12344);
xnor U14789 (N_14789,N_12082,N_12038);
xnor U14790 (N_14790,N_12318,N_12501);
xor U14791 (N_14791,N_12560,N_12171);
nand U14792 (N_14792,N_12133,N_12940);
nand U14793 (N_14793,N_12796,N_13039);
nor U14794 (N_14794,N_13343,N_12786);
and U14795 (N_14795,N_12269,N_13162);
nor U14796 (N_14796,N_13286,N_12587);
and U14797 (N_14797,N_13068,N_13331);
nand U14798 (N_14798,N_13041,N_12131);
and U14799 (N_14799,N_12638,N_13433);
or U14800 (N_14800,N_12222,N_12396);
xor U14801 (N_14801,N_12856,N_12536);
xor U14802 (N_14802,N_13102,N_13494);
nor U14803 (N_14803,N_13069,N_12727);
and U14804 (N_14804,N_12250,N_12469);
xor U14805 (N_14805,N_13074,N_13068);
or U14806 (N_14806,N_13097,N_13386);
and U14807 (N_14807,N_13335,N_12861);
and U14808 (N_14808,N_12520,N_13400);
or U14809 (N_14809,N_12244,N_12195);
and U14810 (N_14810,N_12941,N_12537);
or U14811 (N_14811,N_12399,N_12055);
nand U14812 (N_14812,N_12606,N_13251);
nor U14813 (N_14813,N_12155,N_13137);
nand U14814 (N_14814,N_12371,N_13496);
or U14815 (N_14815,N_12793,N_12622);
or U14816 (N_14816,N_13369,N_12035);
xnor U14817 (N_14817,N_13039,N_12938);
xnor U14818 (N_14818,N_12956,N_13379);
or U14819 (N_14819,N_13212,N_12599);
or U14820 (N_14820,N_12322,N_12383);
nor U14821 (N_14821,N_12405,N_13103);
or U14822 (N_14822,N_12041,N_12476);
xor U14823 (N_14823,N_13234,N_13495);
and U14824 (N_14824,N_12084,N_12312);
or U14825 (N_14825,N_13444,N_12721);
nand U14826 (N_14826,N_12274,N_12781);
nor U14827 (N_14827,N_12564,N_13308);
or U14828 (N_14828,N_12067,N_12415);
nand U14829 (N_14829,N_12989,N_12253);
or U14830 (N_14830,N_13121,N_13438);
nand U14831 (N_14831,N_13434,N_12160);
nand U14832 (N_14832,N_13111,N_12098);
xnor U14833 (N_14833,N_12657,N_13042);
xor U14834 (N_14834,N_12283,N_13442);
xnor U14835 (N_14835,N_12728,N_12950);
or U14836 (N_14836,N_12434,N_13421);
nor U14837 (N_14837,N_13094,N_12711);
and U14838 (N_14838,N_13413,N_12478);
nor U14839 (N_14839,N_12263,N_12316);
and U14840 (N_14840,N_12001,N_12720);
or U14841 (N_14841,N_13064,N_13021);
xnor U14842 (N_14842,N_13436,N_12776);
and U14843 (N_14843,N_13353,N_13445);
nand U14844 (N_14844,N_12858,N_12225);
or U14845 (N_14845,N_12194,N_12129);
or U14846 (N_14846,N_13231,N_13473);
xor U14847 (N_14847,N_13397,N_12937);
and U14848 (N_14848,N_13422,N_12167);
nor U14849 (N_14849,N_12224,N_12088);
or U14850 (N_14850,N_12280,N_12963);
nor U14851 (N_14851,N_12058,N_12331);
and U14852 (N_14852,N_13398,N_12416);
nand U14853 (N_14853,N_12285,N_12278);
xnor U14854 (N_14854,N_13221,N_12095);
or U14855 (N_14855,N_12700,N_12343);
and U14856 (N_14856,N_12782,N_13344);
or U14857 (N_14857,N_12789,N_12773);
nor U14858 (N_14858,N_12188,N_12754);
nand U14859 (N_14859,N_12416,N_13094);
nand U14860 (N_14860,N_13136,N_12761);
or U14861 (N_14861,N_12017,N_12645);
xor U14862 (N_14862,N_12924,N_12350);
xor U14863 (N_14863,N_12288,N_13434);
or U14864 (N_14864,N_12993,N_12705);
or U14865 (N_14865,N_12545,N_12716);
nand U14866 (N_14866,N_13408,N_12073);
nand U14867 (N_14867,N_12910,N_13494);
or U14868 (N_14868,N_13457,N_13008);
nand U14869 (N_14869,N_12349,N_12211);
or U14870 (N_14870,N_12850,N_13217);
and U14871 (N_14871,N_13440,N_12576);
nand U14872 (N_14872,N_12702,N_12432);
nand U14873 (N_14873,N_12632,N_13368);
xor U14874 (N_14874,N_13074,N_13114);
nor U14875 (N_14875,N_12433,N_12936);
nand U14876 (N_14876,N_12620,N_12829);
and U14877 (N_14877,N_12528,N_12095);
nand U14878 (N_14878,N_12227,N_13424);
and U14879 (N_14879,N_13250,N_12815);
or U14880 (N_14880,N_13498,N_13425);
or U14881 (N_14881,N_12238,N_12453);
xnor U14882 (N_14882,N_12007,N_12438);
nand U14883 (N_14883,N_12084,N_12972);
xor U14884 (N_14884,N_12864,N_12990);
or U14885 (N_14885,N_12167,N_12744);
nor U14886 (N_14886,N_12910,N_12608);
or U14887 (N_14887,N_12970,N_12500);
xor U14888 (N_14888,N_12920,N_12259);
nor U14889 (N_14889,N_12141,N_13337);
and U14890 (N_14890,N_12725,N_12262);
or U14891 (N_14891,N_13414,N_12404);
or U14892 (N_14892,N_12165,N_12257);
and U14893 (N_14893,N_13143,N_12913);
or U14894 (N_14894,N_12693,N_13483);
or U14895 (N_14895,N_12879,N_12066);
and U14896 (N_14896,N_13410,N_13466);
nor U14897 (N_14897,N_13021,N_12266);
or U14898 (N_14898,N_13162,N_12737);
or U14899 (N_14899,N_13178,N_12303);
xor U14900 (N_14900,N_12566,N_12505);
nor U14901 (N_14901,N_12693,N_13255);
xnor U14902 (N_14902,N_12292,N_12602);
nand U14903 (N_14903,N_13265,N_12146);
or U14904 (N_14904,N_12574,N_13004);
xnor U14905 (N_14905,N_12697,N_13002);
and U14906 (N_14906,N_12515,N_12082);
and U14907 (N_14907,N_12952,N_12157);
xor U14908 (N_14908,N_12317,N_12066);
or U14909 (N_14909,N_12022,N_12465);
xor U14910 (N_14910,N_12314,N_13245);
or U14911 (N_14911,N_12167,N_13405);
and U14912 (N_14912,N_12957,N_12024);
and U14913 (N_14913,N_12359,N_12023);
nor U14914 (N_14914,N_12253,N_13264);
xor U14915 (N_14915,N_13285,N_12815);
xor U14916 (N_14916,N_13352,N_13408);
nor U14917 (N_14917,N_12069,N_13381);
nor U14918 (N_14918,N_13152,N_12868);
and U14919 (N_14919,N_12466,N_13232);
nor U14920 (N_14920,N_12321,N_12626);
and U14921 (N_14921,N_12563,N_12730);
nand U14922 (N_14922,N_12045,N_13109);
nand U14923 (N_14923,N_13499,N_12836);
nand U14924 (N_14924,N_12557,N_12205);
or U14925 (N_14925,N_12291,N_12667);
nor U14926 (N_14926,N_12576,N_12916);
nand U14927 (N_14927,N_12265,N_12070);
nor U14928 (N_14928,N_12019,N_12398);
and U14929 (N_14929,N_12562,N_12591);
xnor U14930 (N_14930,N_13104,N_12305);
nor U14931 (N_14931,N_12081,N_12482);
and U14932 (N_14932,N_12033,N_13316);
nand U14933 (N_14933,N_13043,N_13036);
or U14934 (N_14934,N_13484,N_13299);
and U14935 (N_14935,N_12942,N_12005);
or U14936 (N_14936,N_12526,N_12303);
and U14937 (N_14937,N_12936,N_12370);
nor U14938 (N_14938,N_12910,N_13442);
xnor U14939 (N_14939,N_13483,N_13117);
or U14940 (N_14940,N_12536,N_12728);
and U14941 (N_14941,N_12188,N_12142);
nand U14942 (N_14942,N_12783,N_13083);
nand U14943 (N_14943,N_13176,N_13259);
or U14944 (N_14944,N_12799,N_13258);
and U14945 (N_14945,N_12198,N_12788);
or U14946 (N_14946,N_12117,N_12617);
and U14947 (N_14947,N_13331,N_13457);
xor U14948 (N_14948,N_12415,N_13404);
nand U14949 (N_14949,N_13409,N_12821);
nand U14950 (N_14950,N_12250,N_12232);
xor U14951 (N_14951,N_13476,N_13177);
nor U14952 (N_14952,N_13491,N_12027);
nor U14953 (N_14953,N_13498,N_13304);
xnor U14954 (N_14954,N_13354,N_12691);
nor U14955 (N_14955,N_13216,N_12287);
nand U14956 (N_14956,N_12730,N_12853);
nand U14957 (N_14957,N_13182,N_12661);
nand U14958 (N_14958,N_12953,N_13472);
nand U14959 (N_14959,N_12866,N_13102);
xor U14960 (N_14960,N_13194,N_12477);
and U14961 (N_14961,N_12887,N_12443);
or U14962 (N_14962,N_13102,N_13080);
nand U14963 (N_14963,N_13497,N_13155);
xnor U14964 (N_14964,N_12960,N_12054);
xor U14965 (N_14965,N_13098,N_13466);
or U14966 (N_14966,N_12212,N_13208);
and U14967 (N_14967,N_12182,N_12279);
nand U14968 (N_14968,N_12764,N_12964);
or U14969 (N_14969,N_12942,N_12935);
nand U14970 (N_14970,N_12645,N_12682);
or U14971 (N_14971,N_12672,N_13478);
nor U14972 (N_14972,N_12969,N_12356);
nor U14973 (N_14973,N_13104,N_13368);
nand U14974 (N_14974,N_12494,N_12267);
nor U14975 (N_14975,N_12828,N_13189);
nor U14976 (N_14976,N_13138,N_12629);
and U14977 (N_14977,N_13356,N_13032);
or U14978 (N_14978,N_13068,N_12151);
and U14979 (N_14979,N_13074,N_12343);
and U14980 (N_14980,N_13200,N_12089);
nand U14981 (N_14981,N_13403,N_13471);
nor U14982 (N_14982,N_12175,N_13246);
nor U14983 (N_14983,N_13301,N_13113);
xnor U14984 (N_14984,N_13074,N_12736);
or U14985 (N_14985,N_13358,N_12120);
nor U14986 (N_14986,N_12170,N_12640);
and U14987 (N_14987,N_13370,N_12520);
and U14988 (N_14988,N_13012,N_12549);
nor U14989 (N_14989,N_12641,N_12220);
xor U14990 (N_14990,N_12680,N_12975);
and U14991 (N_14991,N_13077,N_12438);
or U14992 (N_14992,N_13298,N_12487);
or U14993 (N_14993,N_12228,N_13124);
or U14994 (N_14994,N_13174,N_13223);
nand U14995 (N_14995,N_13148,N_13459);
nand U14996 (N_14996,N_12222,N_13107);
nor U14997 (N_14997,N_12904,N_13031);
xor U14998 (N_14998,N_12290,N_12250);
and U14999 (N_14999,N_13494,N_12281);
or U15000 (N_15000,N_14240,N_13794);
nor U15001 (N_15001,N_14607,N_13859);
or U15002 (N_15002,N_14663,N_14371);
xor U15003 (N_15003,N_14766,N_13834);
nor U15004 (N_15004,N_14850,N_14703);
and U15005 (N_15005,N_14427,N_14504);
nand U15006 (N_15006,N_13547,N_13832);
xor U15007 (N_15007,N_13927,N_14890);
nor U15008 (N_15008,N_13621,N_14405);
or U15009 (N_15009,N_14856,N_14748);
or U15010 (N_15010,N_14138,N_14997);
and U15011 (N_15011,N_14712,N_14666);
nor U15012 (N_15012,N_13803,N_13671);
and U15013 (N_15013,N_14625,N_13963);
and U15014 (N_15014,N_14631,N_13508);
and U15015 (N_15015,N_14550,N_14602);
nor U15016 (N_15016,N_14932,N_14070);
nand U15017 (N_15017,N_14260,N_14589);
nor U15018 (N_15018,N_14769,N_13975);
and U15019 (N_15019,N_13573,N_14894);
and U15020 (N_15020,N_14606,N_14746);
xnor U15021 (N_15021,N_14077,N_14081);
and U15022 (N_15022,N_13601,N_14252);
and U15023 (N_15023,N_14941,N_14216);
or U15024 (N_15024,N_13555,N_13983);
or U15025 (N_15025,N_13749,N_14593);
nor U15026 (N_15026,N_13883,N_13937);
and U15027 (N_15027,N_14868,N_14858);
xnor U15028 (N_15028,N_13625,N_13928);
or U15029 (N_15029,N_14226,N_14721);
xnor U15030 (N_15030,N_14053,N_14379);
and U15031 (N_15031,N_13747,N_14755);
or U15032 (N_15032,N_14425,N_14463);
nand U15033 (N_15033,N_14477,N_14847);
xnor U15034 (N_15034,N_14954,N_13609);
nor U15035 (N_15035,N_13602,N_14416);
nand U15036 (N_15036,N_13929,N_14322);
nand U15037 (N_15037,N_13936,N_14760);
nor U15038 (N_15038,N_14713,N_14392);
nand U15039 (N_15039,N_14943,N_14601);
and U15040 (N_15040,N_14604,N_14571);
and U15041 (N_15041,N_14153,N_14182);
nor U15042 (N_15042,N_13908,N_13824);
or U15043 (N_15043,N_13754,N_13896);
xor U15044 (N_15044,N_14878,N_14638);
and U15045 (N_15045,N_13528,N_13751);
nand U15046 (N_15046,N_13953,N_14750);
or U15047 (N_15047,N_14636,N_13798);
or U15048 (N_15048,N_14978,N_13562);
or U15049 (N_15049,N_14553,N_13713);
nor U15050 (N_15050,N_13505,N_14591);
and U15051 (N_15051,N_14213,N_14711);
xor U15052 (N_15052,N_14318,N_13695);
and U15053 (N_15053,N_14643,N_13990);
xnor U15054 (N_15054,N_14612,N_14520);
or U15055 (N_15055,N_13629,N_14268);
nor U15056 (N_15056,N_14651,N_13652);
xnor U15057 (N_15057,N_13698,N_13513);
xor U15058 (N_15058,N_14101,N_14585);
nor U15059 (N_15059,N_14447,N_13603);
or U15060 (N_15060,N_14881,N_14287);
xnor U15061 (N_15061,N_14333,N_14764);
or U15062 (N_15062,N_13781,N_14278);
and U15063 (N_15063,N_14300,N_14465);
nor U15064 (N_15064,N_14166,N_14665);
nand U15065 (N_15065,N_14420,N_14279);
nand U15066 (N_15066,N_14142,N_14562);
and U15067 (N_15067,N_14446,N_14084);
nand U15068 (N_15068,N_14738,N_14920);
nor U15069 (N_15069,N_14293,N_14782);
nor U15070 (N_15070,N_14702,N_14829);
or U15071 (N_15071,N_13897,N_14029);
nand U15072 (N_15072,N_13947,N_14451);
or U15073 (N_15073,N_14546,N_13767);
nand U15074 (N_15074,N_13768,N_13819);
or U15075 (N_15075,N_13626,N_14384);
xnor U15076 (N_15076,N_14376,N_14343);
or U15077 (N_15077,N_13575,N_13899);
nor U15078 (N_15078,N_14256,N_14164);
xnor U15079 (N_15079,N_13660,N_13790);
nor U15080 (N_15080,N_14910,N_14875);
xor U15081 (N_15081,N_13665,N_13782);
nor U15082 (N_15082,N_14295,N_14179);
or U15083 (N_15083,N_14310,N_14802);
xnor U15084 (N_15084,N_14987,N_13958);
xnor U15085 (N_15085,N_14127,N_14125);
or U15086 (N_15086,N_14065,N_13709);
xnor U15087 (N_15087,N_13820,N_14060);
nand U15088 (N_15088,N_14599,N_14397);
or U15089 (N_15089,N_13735,N_14285);
xnor U15090 (N_15090,N_14752,N_14440);
xnor U15091 (N_15091,N_14202,N_14656);
xor U15092 (N_15092,N_13526,N_14233);
or U15093 (N_15093,N_14388,N_14745);
nand U15094 (N_15094,N_13812,N_13599);
xor U15095 (N_15095,N_14778,N_14298);
xor U15096 (N_15096,N_14921,N_14382);
and U15097 (N_15097,N_14303,N_14496);
xnor U15098 (N_15098,N_13679,N_14935);
nand U15099 (N_15099,N_14556,N_13613);
nor U15100 (N_15100,N_13595,N_13616);
nand U15101 (N_15101,N_14775,N_13539);
nor U15102 (N_15102,N_14709,N_13909);
nand U15103 (N_15103,N_14234,N_13814);
and U15104 (N_15104,N_14359,N_14590);
xnor U15105 (N_15105,N_13638,N_14598);
and U15106 (N_15106,N_14444,N_14594);
or U15107 (N_15107,N_14937,N_13580);
nand U15108 (N_15108,N_13576,N_14885);
nand U15109 (N_15109,N_14035,N_14386);
nor U15110 (N_15110,N_13887,N_13653);
and U15111 (N_15111,N_14021,N_14025);
nand U15112 (N_15112,N_14646,N_14100);
and U15113 (N_15113,N_14966,N_14939);
xnor U15114 (N_15114,N_14434,N_13736);
nor U15115 (N_15115,N_14308,N_14493);
nand U15116 (N_15116,N_14089,N_14495);
or U15117 (N_15117,N_13755,N_14369);
nor U15118 (N_15118,N_14522,N_13942);
nor U15119 (N_15119,N_13651,N_14799);
nand U15120 (N_15120,N_14326,N_14759);
or U15121 (N_15121,N_14820,N_14246);
nor U15122 (N_15122,N_13657,N_14616);
or U15123 (N_15123,N_14879,N_13825);
xor U15124 (N_15124,N_13729,N_13787);
or U15125 (N_15125,N_13615,N_14902);
nand U15126 (N_15126,N_14149,N_13699);
nor U15127 (N_15127,N_14155,N_14706);
nand U15128 (N_15128,N_13639,N_14767);
xnor U15129 (N_15129,N_13804,N_14154);
xor U15130 (N_15130,N_14030,N_14803);
and U15131 (N_15131,N_14860,N_14812);
or U15132 (N_15132,N_14160,N_14331);
or U15133 (N_15133,N_13740,N_14524);
xor U15134 (N_15134,N_14112,N_14561);
and U15135 (N_15135,N_13635,N_13966);
and U15136 (N_15136,N_14510,N_14691);
nor U15137 (N_15137,N_14050,N_13907);
nor U15138 (N_15138,N_13588,N_14049);
nand U15139 (N_15139,N_14985,N_13822);
and U15140 (N_15140,N_14854,N_13543);
and U15141 (N_15141,N_14757,N_14309);
nand U15142 (N_15142,N_14972,N_14302);
and U15143 (N_15143,N_13659,N_14058);
nor U15144 (N_15144,N_14227,N_14664);
nor U15145 (N_15145,N_13962,N_14000);
nor U15146 (N_15146,N_14042,N_13873);
nor U15147 (N_15147,N_14649,N_13731);
xnor U15148 (N_15148,N_13581,N_13989);
nand U15149 (N_15149,N_14611,N_13536);
nand U15150 (N_15150,N_14412,N_13944);
or U15151 (N_15151,N_13501,N_14063);
xnor U15152 (N_15152,N_14175,N_13850);
nand U15153 (N_15153,N_13813,N_14041);
or U15154 (N_15154,N_13727,N_13745);
nand U15155 (N_15155,N_14116,N_14032);
xnor U15156 (N_15156,N_14187,N_14549);
xor U15157 (N_15157,N_13673,N_14507);
nor U15158 (N_15158,N_14689,N_14265);
nand U15159 (N_15159,N_14099,N_14040);
nand U15160 (N_15160,N_13622,N_14635);
xnor U15161 (N_15161,N_14765,N_14066);
and U15162 (N_15162,N_14873,N_14708);
nor U15163 (N_15163,N_14626,N_13807);
and U15164 (N_15164,N_13821,N_14443);
nor U15165 (N_15165,N_14271,N_14110);
and U15166 (N_15166,N_14837,N_13750);
and U15167 (N_15167,N_13548,N_14121);
nor U15168 (N_15168,N_14224,N_14565);
and U15169 (N_15169,N_13567,N_14918);
xnor U15170 (N_15170,N_14010,N_14073);
nand U15171 (N_15171,N_13738,N_13707);
or U15172 (N_15172,N_14705,N_14316);
xnor U15173 (N_15173,N_14104,N_14413);
and U15174 (N_15174,N_14483,N_13586);
and U15175 (N_15175,N_14450,N_13847);
nand U15176 (N_15176,N_14617,N_14418);
nor U15177 (N_15177,N_13633,N_14117);
nand U15178 (N_15178,N_14952,N_14011);
xnor U15179 (N_15179,N_14682,N_14056);
or U15180 (N_15180,N_14675,N_14807);
nor U15181 (N_15181,N_14292,N_14022);
and U15182 (N_15182,N_14317,N_14904);
and U15183 (N_15183,N_14909,N_13943);
xnor U15184 (N_15184,N_14728,N_13996);
and U15185 (N_15185,N_14068,N_13714);
xor U15186 (N_15186,N_14961,N_13972);
and U15187 (N_15187,N_13668,N_14845);
or U15188 (N_15188,N_14124,N_13677);
nand U15189 (N_15189,N_14018,N_14603);
and U15190 (N_15190,N_14658,N_13796);
nand U15191 (N_15191,N_13620,N_14628);
nand U15192 (N_15192,N_14136,N_13866);
or U15193 (N_15193,N_13565,N_14901);
nand U15194 (N_15194,N_14481,N_14560);
and U15195 (N_15195,N_13988,N_14869);
and U15196 (N_15196,N_14639,N_13889);
xnor U15197 (N_15197,N_14683,N_14687);
nor U15198 (N_15198,N_13941,N_14215);
and U15199 (N_15199,N_14681,N_14428);
nand U15200 (N_15200,N_14176,N_14061);
xor U15201 (N_15201,N_14335,N_13788);
and U15202 (N_15202,N_14171,N_14338);
and U15203 (N_15203,N_14743,N_13886);
xnor U15204 (N_15204,N_14431,N_14484);
and U15205 (N_15205,N_14119,N_14406);
nor U15206 (N_15206,N_13596,N_14788);
nor U15207 (N_15207,N_14357,N_14389);
and U15208 (N_15208,N_14783,N_14533);
or U15209 (N_15209,N_14632,N_14963);
nand U15210 (N_15210,N_14690,N_14844);
and U15211 (N_15211,N_14395,N_13959);
xnor U15212 (N_15212,N_13758,N_14181);
nor U15213 (N_15213,N_13828,N_14716);
nand U15214 (N_15214,N_14334,N_13518);
xor U15215 (N_15215,N_14732,N_13946);
nand U15216 (N_15216,N_14355,N_14544);
or U15217 (N_15217,N_13503,N_14538);
or U15218 (N_15218,N_14079,N_13678);
xor U15219 (N_15219,N_13840,N_14194);
or U15220 (N_15220,N_14055,N_14367);
nand U15221 (N_15221,N_14086,N_13692);
nand U15222 (N_15222,N_14016,N_14156);
xnor U15223 (N_15223,N_14509,N_14051);
xor U15224 (N_15224,N_14211,N_14014);
xor U15225 (N_15225,N_13512,N_14796);
and U15226 (N_15226,N_14914,N_13845);
or U15227 (N_15227,N_13534,N_14087);
xnor U15228 (N_15228,N_13656,N_14259);
or U15229 (N_15229,N_14903,N_13835);
nor U15230 (N_15230,N_14401,N_14193);
nand U15231 (N_15231,N_14830,N_13545);
and U15232 (N_15232,N_14015,N_13711);
xor U15233 (N_15233,N_14971,N_14973);
nand U15234 (N_15234,N_14170,N_14286);
and U15235 (N_15235,N_14196,N_14685);
xor U15236 (N_15236,N_14185,N_14059);
or U15237 (N_15237,N_14177,N_13506);
and U15238 (N_15238,N_13570,N_14002);
or U15239 (N_15239,N_14995,N_14186);
or U15240 (N_15240,N_14623,N_13862);
and U15241 (N_15241,N_14569,N_13974);
and U15242 (N_15242,N_14573,N_13921);
nor U15243 (N_15243,N_14884,N_14669);
nor U15244 (N_15244,N_14109,N_14809);
and U15245 (N_15245,N_14169,N_13888);
or U15246 (N_15246,N_14365,N_14661);
xnor U15247 (N_15247,N_14008,N_14487);
nand U15248 (N_15248,N_14892,N_13885);
or U15249 (N_15249,N_14818,N_14518);
nand U15250 (N_15250,N_14624,N_14784);
nand U15251 (N_15251,N_14574,N_13724);
xor U15252 (N_15252,N_14276,N_14974);
nor U15253 (N_15253,N_13611,N_13705);
and U15254 (N_15254,N_13637,N_13871);
xor U15255 (N_15255,N_14387,N_14724);
nand U15256 (N_15256,N_13805,N_14861);
xnor U15257 (N_15257,N_13895,N_13893);
nand U15258 (N_15258,N_14654,N_14200);
and U15259 (N_15259,N_13721,N_14848);
and U15260 (N_15260,N_14859,N_14426);
or U15261 (N_15261,N_14173,N_14323);
and U15262 (N_15262,N_13979,N_13710);
or U15263 (N_15263,N_14208,N_13510);
and U15264 (N_15264,N_14733,N_14304);
nor U15265 (N_15265,N_14964,N_14871);
nor U15266 (N_15266,N_14137,N_13589);
or U15267 (N_15267,N_13708,N_14763);
nor U15268 (N_15268,N_13892,N_14588);
or U15269 (N_15269,N_13900,N_14078);
or U15270 (N_15270,N_13702,N_14189);
nand U15271 (N_15271,N_14870,N_14991);
or U15272 (N_15272,N_14835,N_13655);
and U15273 (N_15273,N_14969,N_14877);
or U15274 (N_15274,N_14122,N_13761);
nor U15275 (N_15275,N_13522,N_14301);
nor U15276 (N_15276,N_13981,N_14673);
or U15277 (N_15277,N_13786,N_14057);
or U15278 (N_15278,N_14191,N_14960);
or U15279 (N_15279,N_14223,N_14003);
or U15280 (N_15280,N_14980,N_13682);
xor U15281 (N_15281,N_14229,N_13507);
xnor U15282 (N_15282,N_14751,N_13956);
nand U15283 (N_15283,N_14773,N_13583);
xor U15284 (N_15284,N_14648,N_14494);
nand U15285 (N_15285,N_14576,N_14126);
nand U15286 (N_15286,N_13864,N_14797);
xor U15287 (N_15287,N_13823,N_14393);
xor U15288 (N_15288,N_13879,N_14699);
nand U15289 (N_15289,N_14422,N_14324);
xor U15290 (N_15290,N_14356,N_14421);
nor U15291 (N_15291,N_14929,N_13760);
and U15292 (N_15292,N_13771,N_14069);
or U15293 (N_15293,N_14325,N_14471);
xor U15294 (N_15294,N_13756,N_14619);
xnor U15295 (N_15295,N_13955,N_14620);
nand U15296 (N_15296,N_14836,N_13569);
xor U15297 (N_15297,N_13774,N_13872);
or U15298 (N_15298,N_14466,N_14965);
nand U15299 (N_15299,N_14151,N_14183);
and U15300 (N_15300,N_13500,N_13865);
nor U15301 (N_15301,N_14828,N_13687);
nand U15302 (N_15302,N_13757,N_14740);
or U15303 (N_15303,N_13770,N_14345);
or U15304 (N_15304,N_14147,N_14207);
nor U15305 (N_15305,N_14314,N_14558);
nor U15306 (N_15306,N_14106,N_14131);
nand U15307 (N_15307,N_14092,N_14157);
nor U15308 (N_15308,N_13627,N_14097);
and U15309 (N_15309,N_13725,N_13644);
or U15310 (N_15310,N_14178,N_13739);
xor U15311 (N_15311,N_14795,N_13894);
nand U15312 (N_15312,N_14158,N_14103);
nor U15313 (N_15313,N_13610,N_13723);
nand U15314 (N_15314,N_13982,N_14714);
and U15315 (N_15315,N_14248,N_13667);
nor U15316 (N_15316,N_14277,N_13560);
and U15317 (N_15317,N_14013,N_14190);
nor U15318 (N_15318,N_14354,N_14517);
xor U15319 (N_15319,N_14793,N_13577);
or U15320 (N_15320,N_13861,N_14439);
nor U15321 (N_15321,N_14218,N_14288);
and U15322 (N_15322,N_14575,N_13641);
xor U15323 (N_15323,N_14402,N_14956);
and U15324 (N_15324,N_13561,N_14230);
and U15325 (N_15325,N_14542,N_13511);
xor U15326 (N_15326,N_14459,N_13915);
or U15327 (N_15327,N_14129,N_13792);
and U15328 (N_15328,N_14250,N_14243);
xor U15329 (N_15329,N_13516,N_14534);
xnor U15330 (N_15330,N_14266,N_13780);
and U15331 (N_15331,N_13715,N_14584);
or U15332 (N_15332,N_14815,N_14414);
xnor U15333 (N_15333,N_14486,N_13604);
xnor U15334 (N_15334,N_14238,N_13848);
and U15335 (N_15335,N_14315,N_14373);
xnor U15336 (N_15336,N_14919,N_14851);
nand U15337 (N_15337,N_14916,N_14957);
and U15338 (N_15338,N_13697,N_13933);
and U15339 (N_15339,N_14707,N_14726);
or U15340 (N_15340,N_14174,N_14228);
nor U15341 (N_15341,N_14697,N_14120);
nand U15342 (N_15342,N_14536,N_13808);
and U15343 (N_15343,N_13614,N_14415);
and U15344 (N_15344,N_14306,N_14786);
or U15345 (N_15345,N_14653,N_14905);
nor U15346 (N_15346,N_14291,N_14197);
nor U15347 (N_15347,N_14811,N_14236);
nor U15348 (N_15348,N_13965,N_14201);
or U15349 (N_15349,N_13954,N_14727);
and U15350 (N_15350,N_14461,N_14470);
and U15351 (N_15351,N_14841,N_13579);
nand U15352 (N_15352,N_14672,N_13919);
and U15353 (N_15353,N_13619,N_14363);
xor U15354 (N_15354,N_14254,N_14482);
nand U15355 (N_15355,N_14381,N_13732);
or U15356 (N_15356,N_13997,N_14044);
xnor U15357 (N_15357,N_14284,N_13618);
or U15358 (N_15358,N_13546,N_14614);
nand U15359 (N_15359,N_14358,N_13951);
xnor U15360 (N_15360,N_14134,N_13878);
or U15361 (N_15361,N_14438,N_14351);
nand U15362 (N_15362,N_14052,N_14258);
xor U15363 (N_15363,N_13945,N_14630);
nor U15364 (N_15364,N_14776,N_13931);
nor U15365 (N_15365,N_13830,N_14489);
nand U15366 (N_15366,N_14474,N_14513);
nand U15367 (N_15367,N_14693,N_14080);
xor U15368 (N_15368,N_13791,N_14380);
and U15369 (N_15369,N_13875,N_14977);
nor U15370 (N_15370,N_14328,N_13612);
nand U15371 (N_15371,N_13591,N_14390);
nand U15372 (N_15372,N_13863,N_14305);
nand U15373 (N_15373,N_13765,N_14548);
xor U15374 (N_15374,N_14475,N_14020);
nand U15375 (N_15375,N_14814,N_14742);
nand U15376 (N_15376,N_13606,N_14953);
xor U15377 (N_15377,N_14383,N_13901);
or U15378 (N_15378,N_14959,N_14054);
nand U15379 (N_15379,N_13844,N_13906);
nand U15380 (N_15380,N_14255,N_14928);
and U15381 (N_15381,N_14852,N_13789);
nand U15382 (N_15382,N_14645,N_13818);
xor U15383 (N_15383,N_13891,N_13842);
nor U15384 (N_15384,N_13874,N_14251);
and U15385 (N_15385,N_13557,N_14735);
and U15386 (N_15386,N_14955,N_14088);
and U15387 (N_15387,N_13759,N_14912);
nand U15388 (N_15388,N_14777,N_14942);
xnor U15389 (N_15389,N_14168,N_14867);
xor U15390 (N_15390,N_13593,N_14994);
xnor U15391 (N_15391,N_13992,N_14378);
or U15392 (N_15392,N_14102,N_13999);
xnor U15393 (N_15393,N_14568,N_14514);
nor U15394 (N_15394,N_14700,N_14801);
or U15395 (N_15395,N_14172,N_13742);
nand U15396 (N_15396,N_14167,N_13960);
nand U15397 (N_15397,N_13530,N_14453);
nand U15398 (N_15398,N_14281,N_14846);
xnor U15399 (N_15399,N_13645,N_13925);
nand U15400 (N_15400,N_13689,N_14033);
or U15401 (N_15401,N_14640,N_14849);
or U15402 (N_15402,N_13672,N_14608);
nor U15403 (N_15403,N_13741,N_13504);
and U15404 (N_15404,N_13597,N_14794);
nand U15405 (N_15405,N_14272,N_14113);
nand U15406 (N_15406,N_13552,N_14949);
and U15407 (N_15407,N_13957,N_14537);
and U15408 (N_15408,N_13867,N_14241);
or U15409 (N_15409,N_14822,N_14899);
xor U15410 (N_15410,N_14898,N_14307);
or U15411 (N_15411,N_14789,N_14637);
or U15412 (N_15412,N_13647,N_14992);
nor U15413 (N_15413,N_14083,N_13683);
xnor U15414 (N_15414,N_13775,N_13802);
or U15415 (N_15415,N_14289,N_13681);
and U15416 (N_15416,N_14135,N_14660);
xnor U15417 (N_15417,N_13926,N_13712);
nor U15418 (N_15418,N_14294,N_14855);
xnor U15419 (N_15419,N_13795,N_14618);
or U15420 (N_15420,N_14214,N_13809);
nor U15421 (N_15421,N_14970,N_14749);
nand U15422 (N_15422,N_14543,N_13726);
and U15423 (N_15423,N_14722,N_14979);
xnor U15424 (N_15424,N_13829,N_14586);
or U15425 (N_15425,N_14621,N_14128);
xnor U15426 (N_15426,N_14417,N_14865);
nor U15427 (N_15427,N_13924,N_14332);
nor U15428 (N_15428,N_13949,N_14296);
nand U15429 (N_15429,N_14827,N_14824);
nor U15430 (N_15430,N_14813,N_14924);
and U15431 (N_15431,N_13664,N_13554);
xor U15432 (N_15432,N_13806,N_13592);
or U15433 (N_15433,N_14600,N_14261);
and U15434 (N_15434,N_14976,N_13800);
and U15435 (N_15435,N_14212,N_14445);
and U15436 (N_15436,N_14968,N_14529);
xor U15437 (N_15437,N_13799,N_14832);
nand U15438 (N_15438,N_14244,N_14350);
nor U15439 (N_15439,N_14046,N_14671);
nand U15440 (N_15440,N_14290,N_14579);
and U15441 (N_15441,N_13985,N_14981);
nor U15442 (N_15442,N_14831,N_14161);
nor U15443 (N_15443,N_14988,N_14944);
and U15444 (N_15444,N_14516,N_13854);
xnor U15445 (N_15445,N_14499,N_14090);
or U15446 (N_15446,N_13841,N_14017);
or U15447 (N_15447,N_14432,N_13935);
xnor U15448 (N_15448,N_14715,N_14026);
nand U15449 (N_15449,N_14876,N_14950);
xnor U15450 (N_15450,N_14922,N_14269);
or U15451 (N_15451,N_14497,N_14729);
and U15452 (N_15452,N_13662,N_14001);
xor U15453 (N_15453,N_14990,N_13764);
and U15454 (N_15454,N_13632,N_13624);
xor U15455 (N_15455,N_14679,N_14774);
nand U15456 (N_15456,N_14037,N_14231);
xnor U15457 (N_15457,N_13532,N_13696);
or U15458 (N_15458,N_13922,N_13521);
xnor U15459 (N_15459,N_13568,N_13833);
nand U15460 (N_15460,N_14490,N_13515);
or U15461 (N_15461,N_14886,N_13544);
xnor U15462 (N_15462,N_13753,N_14398);
nand U15463 (N_15463,N_13533,N_14734);
nor U15464 (N_15464,N_14840,N_14622);
or U15465 (N_15465,N_13704,N_14834);
xor U15466 (N_15466,N_14578,N_13826);
or U15467 (N_15467,N_14580,N_14491);
and U15468 (N_15468,N_14429,N_14337);
and U15469 (N_15469,N_14423,N_14882);
and U15470 (N_15470,N_14821,N_14436);
nor U15471 (N_15471,N_14843,N_14864);
and U15472 (N_15472,N_14915,N_13661);
and U15473 (N_15473,N_13855,N_14555);
or U15474 (N_15474,N_14460,N_14024);
nand U15475 (N_15475,N_13884,N_14771);
xnor U15476 (N_15476,N_13779,N_14720);
nor U15477 (N_15477,N_14132,N_13571);
and U15478 (N_15478,N_14476,N_13553);
and U15479 (N_15479,N_13607,N_14019);
nor U15480 (N_15480,N_13769,N_14893);
xor U15481 (N_15481,N_14696,N_14874);
or U15482 (N_15482,N_14435,N_14264);
xnor U15483 (N_15483,N_13703,N_14982);
nor U15484 (N_15484,N_13793,N_14396);
or U15485 (N_15485,N_14634,N_14552);
nor U15486 (N_15486,N_14808,N_14344);
and U15487 (N_15487,N_13973,N_14004);
nand U15488 (N_15488,N_14933,N_14975);
and U15489 (N_15489,N_14780,N_14094);
xnor U15490 (N_15490,N_14195,N_14838);
or U15491 (N_15491,N_13849,N_14140);
or U15492 (N_15492,N_13811,N_13932);
nand U15493 (N_15493,N_13853,N_14857);
and U15494 (N_15494,N_14062,N_14005);
or U15495 (N_15495,N_13914,N_14374);
or U15496 (N_15496,N_14217,N_13984);
or U15497 (N_15497,N_13572,N_14889);
nand U15498 (N_15498,N_14442,N_13675);
xnor U15499 (N_15499,N_13509,N_14452);
or U15500 (N_15500,N_13977,N_14816);
and U15501 (N_15501,N_14237,N_14045);
nor U15502 (N_15502,N_13970,N_14772);
nand U15503 (N_15503,N_14887,N_13628);
nor U15504 (N_15504,N_14863,N_14688);
or U15505 (N_15505,N_13994,N_14242);
nand U15506 (N_15506,N_14564,N_13882);
nor U15507 (N_15507,N_14093,N_14572);
or U15508 (N_15508,N_13691,N_14430);
xor U15509 (N_15509,N_14409,N_14360);
xnor U15510 (N_15510,N_14592,N_14647);
or U15511 (N_15511,N_13594,N_13658);
and U15512 (N_15512,N_14947,N_14152);
or U15513 (N_15513,N_14023,N_14123);
and U15514 (N_15514,N_14133,N_13716);
or U15515 (N_15515,N_14114,N_14948);
nand U15516 (N_15516,N_13690,N_14043);
xor U15517 (N_15517,N_14670,N_14523);
xnor U15518 (N_15518,N_14519,N_14512);
or U15519 (N_15519,N_14551,N_14377);
or U15520 (N_15520,N_14785,N_13519);
xnor U15521 (N_15521,N_13541,N_13674);
nand U15522 (N_15522,N_14521,N_14725);
or U15523 (N_15523,N_14411,N_13890);
or U15524 (N_15524,N_14547,N_14336);
nand U15525 (N_15525,N_13550,N_14826);
and U15526 (N_15526,N_13752,N_13964);
nor U15527 (N_15527,N_14498,N_14506);
nand U15528 (N_15528,N_13762,N_14370);
nand U15529 (N_15529,N_14515,N_14257);
and U15530 (N_15530,N_13952,N_14330);
and U15531 (N_15531,N_14209,N_13701);
xnor U15532 (N_15532,N_14888,N_13810);
and U15533 (N_15533,N_14686,N_13538);
nand U15534 (N_15534,N_14754,N_13531);
and U15535 (N_15535,N_13558,N_14270);
or U15536 (N_15536,N_14199,N_14232);
nand U15537 (N_15537,N_14613,N_14719);
xnor U15538 (N_15538,N_14853,N_14931);
and U15539 (N_15539,N_14404,N_13920);
xnor U15540 (N_15540,N_13590,N_13608);
and U15541 (N_15541,N_14945,N_13587);
nand U15542 (N_15542,N_14203,N_13670);
nand U15543 (N_15543,N_13514,N_13930);
xnor U15544 (N_15544,N_13563,N_14641);
or U15545 (N_15545,N_14508,N_14321);
and U15546 (N_15546,N_14235,N_13578);
nor U15547 (N_15547,N_14804,N_13584);
or U15548 (N_15548,N_14701,N_14692);
nor U15549 (N_15549,N_14605,N_14680);
nor U15550 (N_15550,N_14946,N_14473);
nor U15551 (N_15551,N_14781,N_13870);
and U15552 (N_15552,N_13831,N_14221);
and U15553 (N_15553,N_13815,N_14327);
and U15554 (N_15554,N_14747,N_14839);
or U15555 (N_15555,N_13600,N_13642);
and U15556 (N_15556,N_14076,N_14403);
and U15557 (N_15557,N_13717,N_14723);
nor U15558 (N_15558,N_13934,N_14741);
or U15559 (N_15559,N_14989,N_14282);
nor U15560 (N_15560,N_13917,N_13858);
or U15561 (N_15561,N_14454,N_13904);
nand U15562 (N_15562,N_14245,N_14262);
nand U15563 (N_15563,N_14342,N_14570);
xnor U15564 (N_15564,N_14031,N_14455);
and U15565 (N_15565,N_13784,N_14698);
or U15566 (N_15566,N_14394,N_14895);
nand U15567 (N_15567,N_14610,N_13772);
and U15568 (N_15568,N_13730,N_14349);
nor U15569 (N_15569,N_13910,N_14609);
nor U15570 (N_15570,N_14267,N_14501);
nand U15571 (N_15571,N_14275,N_14677);
nand U15572 (N_15572,N_14348,N_13916);
and U15573 (N_15573,N_13763,N_13881);
xor U15574 (N_15574,N_14999,N_14934);
and U15575 (N_15575,N_13913,N_13938);
or U15576 (N_15576,N_13971,N_14312);
or U15577 (N_15577,N_14996,N_14940);
nor U15578 (N_15578,N_14180,N_13991);
and U15579 (N_15579,N_14710,N_13556);
nand U15580 (N_15580,N_13744,N_13525);
xor U15581 (N_15581,N_13631,N_14525);
nor U15582 (N_15582,N_13585,N_13903);
nand U15583 (N_15583,N_13783,N_14472);
and U15584 (N_15584,N_14539,N_14247);
nand U15585 (N_15585,N_13851,N_13993);
nand U15586 (N_15586,N_13816,N_13846);
nor U15587 (N_15587,N_14530,N_13838);
xnor U15588 (N_15588,N_14400,N_13636);
xnor U15589 (N_15589,N_13719,N_14911);
and U15590 (N_15590,N_14833,N_13986);
nand U15591 (N_15591,N_14039,N_14668);
nand U15592 (N_15592,N_14198,N_14205);
nand U15593 (N_15593,N_13574,N_14437);
or U15594 (N_15594,N_14184,N_14441);
xor U15595 (N_15595,N_13746,N_14297);
and U15596 (N_15596,N_14192,N_14718);
nor U15597 (N_15597,N_14792,N_14249);
nand U15598 (N_15598,N_14798,N_13648);
or U15599 (N_15599,N_13734,N_13968);
nor U15600 (N_15600,N_13827,N_14737);
or U15601 (N_15601,N_14009,N_14341);
nand U15602 (N_15602,N_14111,N_13654);
and U15603 (N_15603,N_14372,N_14075);
nor U15604 (N_15604,N_13676,N_14457);
and U15605 (N_15605,N_14141,N_14143);
xor U15606 (N_15606,N_13773,N_13857);
xor U15607 (N_15607,N_14652,N_13634);
and U15608 (N_15608,N_13797,N_14115);
xor U15609 (N_15609,N_14503,N_14883);
nand U15610 (N_15610,N_14038,N_13948);
or U15611 (N_15611,N_14930,N_13918);
nor U15612 (N_15612,N_14532,N_14926);
or U15613 (N_15613,N_14566,N_13978);
nand U15614 (N_15614,N_13649,N_14210);
and U15615 (N_15615,N_14962,N_14082);
nor U15616 (N_15616,N_14540,N_13777);
and U15617 (N_15617,N_14162,N_14758);
and U15618 (N_15618,N_14627,N_14554);
nand U15619 (N_15619,N_13663,N_13877);
xor U15620 (N_15620,N_14165,N_14583);
xnor U15621 (N_15621,N_14449,N_13950);
or U15622 (N_15622,N_14842,N_13980);
or U15623 (N_15623,N_13643,N_13693);
xor U15624 (N_15624,N_13839,N_14007);
nand U15625 (N_15625,N_13520,N_13912);
or U15626 (N_15626,N_13785,N_13527);
or U15627 (N_15627,N_13733,N_14787);
or U15628 (N_15628,N_14385,N_14399);
nor U15629 (N_15629,N_13523,N_13535);
xor U15630 (N_15630,N_14225,N_13998);
nand U15631 (N_15631,N_14644,N_14913);
nor U15632 (N_15632,N_14074,N_14790);
xor U15633 (N_15633,N_14047,N_14067);
and U15634 (N_15634,N_14559,N_14917);
or U15635 (N_15635,N_14938,N_14219);
nand U15636 (N_15636,N_14819,N_14048);
nand U15637 (N_15637,N_14615,N_14577);
nor U15638 (N_15638,N_14655,N_14925);
nor U15639 (N_15639,N_14967,N_14433);
or U15640 (N_15640,N_14587,N_13961);
xor U15641 (N_15641,N_14467,N_14872);
and U15642 (N_15642,N_13549,N_14526);
nor U15643 (N_15643,N_14704,N_14505);
nand U15644 (N_15644,N_14694,N_14163);
nor U15645 (N_15645,N_14145,N_14206);
xnor U15646 (N_15646,N_13540,N_14253);
nand U15647 (N_15647,N_14028,N_14419);
nand U15648 (N_15648,N_14146,N_13559);
or U15649 (N_15649,N_13776,N_14464);
or U15650 (N_15650,N_14339,N_14958);
or U15651 (N_15651,N_14072,N_13564);
and U15652 (N_15652,N_13685,N_13801);
or U15653 (N_15653,N_14364,N_13868);
xor U15654 (N_15654,N_14805,N_14375);
nor U15655 (N_15655,N_14034,N_14468);
xnor U15656 (N_15656,N_14500,N_14071);
nand U15657 (N_15657,N_14313,N_14511);
xor U15658 (N_15658,N_13623,N_14880);
xor U15659 (N_15659,N_13969,N_13684);
and U15660 (N_15660,N_14105,N_14762);
or U15661 (N_15661,N_14353,N_13939);
xor U15662 (N_15662,N_13700,N_14361);
nor U15663 (N_15663,N_14329,N_13617);
nand U15664 (N_15664,N_14993,N_14347);
nor U15665 (N_15665,N_14366,N_14891);
nand U15666 (N_15666,N_13630,N_14667);
or U15667 (N_15667,N_14036,N_14362);
xor U15668 (N_15668,N_14012,N_14064);
xnor U15669 (N_15669,N_14108,N_13905);
nor U15670 (N_15670,N_14779,N_14407);
or U15671 (N_15671,N_14674,N_13837);
or U15672 (N_15672,N_14770,N_14936);
or U15673 (N_15673,N_14791,N_14204);
or U15674 (N_15674,N_14159,N_14998);
xor U15675 (N_15675,N_14107,N_14424);
nand U15676 (N_15676,N_14263,N_13680);
nand U15677 (N_15677,N_14485,N_13817);
and U15678 (N_15678,N_14391,N_14462);
xor U15679 (N_15679,N_13706,N_14695);
nand U15680 (N_15680,N_14091,N_14557);
xor U15681 (N_15681,N_14581,N_14027);
xor U15682 (N_15682,N_14085,N_14239);
or U15683 (N_15683,N_13718,N_14545);
xnor U15684 (N_15684,N_14098,N_14736);
nand U15685 (N_15685,N_14130,N_14006);
xor U15686 (N_15686,N_13967,N_13876);
nor U15687 (N_15687,N_14678,N_14118);
xor U15688 (N_15688,N_14096,N_14642);
and U15689 (N_15689,N_14352,N_14567);
nand U15690 (N_15690,N_14823,N_13766);
nor U15691 (N_15691,N_14768,N_13688);
or U15692 (N_15692,N_14448,N_13843);
or U15693 (N_15693,N_14563,N_14761);
and U15694 (N_15694,N_14340,N_13940);
xnor U15695 (N_15695,N_14825,N_13722);
nand U15696 (N_15696,N_14469,N_14662);
or U15697 (N_15697,N_13551,N_13836);
nor U15698 (N_15698,N_14188,N_13694);
or U15699 (N_15699,N_13902,N_14456);
or U15700 (N_15700,N_14800,N_13737);
nand U15701 (N_15701,N_14753,N_14657);
or U15702 (N_15702,N_14144,N_14346);
and U15703 (N_15703,N_14717,N_14900);
and U15704 (N_15704,N_14908,N_14150);
nor U15705 (N_15705,N_14923,N_14595);
nor U15706 (N_15706,N_14983,N_14458);
nor U15707 (N_15707,N_13524,N_13605);
or U15708 (N_15708,N_13646,N_13860);
or U15709 (N_15709,N_14810,N_13987);
nand U15710 (N_15710,N_13856,N_13517);
or U15711 (N_15711,N_13669,N_14596);
nand U15712 (N_15712,N_14951,N_14320);
nor U15713 (N_15713,N_14629,N_14597);
and U15714 (N_15714,N_14488,N_14896);
nand U15715 (N_15715,N_13686,N_14528);
nor U15716 (N_15716,N_13743,N_14319);
or U15717 (N_15717,N_14684,N_13923);
xor U15718 (N_15718,N_13728,N_14220);
xnor U15719 (N_15719,N_13778,N_14756);
xnor U15720 (N_15720,N_14731,N_14897);
xor U15721 (N_15721,N_14408,N_14139);
xnor U15722 (N_15722,N_14479,N_14478);
or U15723 (N_15723,N_13976,N_13720);
nor U15724 (N_15724,N_14817,N_14535);
or U15725 (N_15725,N_14273,N_14866);
and U15726 (N_15726,N_14986,N_13748);
nor U15727 (N_15727,N_14744,N_13852);
or U15728 (N_15728,N_14502,N_13542);
or U15729 (N_15729,N_14650,N_14531);
nor U15730 (N_15730,N_14862,N_14984);
nor U15731 (N_15731,N_14280,N_13582);
and U15732 (N_15732,N_14676,N_14633);
xor U15733 (N_15733,N_13529,N_14541);
or U15734 (N_15734,N_13869,N_14095);
nor U15735 (N_15735,N_13640,N_14806);
xnor U15736 (N_15736,N_14906,N_13911);
nor U15737 (N_15737,N_14311,N_13650);
and U15738 (N_15738,N_14527,N_14148);
nand U15739 (N_15739,N_14283,N_14730);
xnor U15740 (N_15740,N_13898,N_14659);
or U15741 (N_15741,N_14480,N_14274);
nand U15742 (N_15742,N_13995,N_13666);
xnor U15743 (N_15743,N_14368,N_13537);
and U15744 (N_15744,N_13566,N_14927);
nor U15745 (N_15745,N_14739,N_13598);
or U15746 (N_15746,N_14907,N_14410);
or U15747 (N_15747,N_13880,N_14582);
or U15748 (N_15748,N_14492,N_14299);
xor U15749 (N_15749,N_14222,N_13502);
and U15750 (N_15750,N_13898,N_13560);
nand U15751 (N_15751,N_14120,N_13754);
or U15752 (N_15752,N_13934,N_14055);
and U15753 (N_15753,N_13898,N_14939);
and U15754 (N_15754,N_14614,N_14455);
xor U15755 (N_15755,N_13845,N_13983);
or U15756 (N_15756,N_14497,N_14466);
nand U15757 (N_15757,N_14048,N_14754);
xnor U15758 (N_15758,N_14946,N_14120);
or U15759 (N_15759,N_14088,N_13569);
nand U15760 (N_15760,N_14245,N_14472);
or U15761 (N_15761,N_14385,N_14621);
or U15762 (N_15762,N_14428,N_14044);
nand U15763 (N_15763,N_14258,N_14231);
xnor U15764 (N_15764,N_14252,N_14463);
and U15765 (N_15765,N_14849,N_14168);
and U15766 (N_15766,N_14531,N_14883);
or U15767 (N_15767,N_13616,N_14440);
and U15768 (N_15768,N_14044,N_14194);
or U15769 (N_15769,N_14897,N_14068);
or U15770 (N_15770,N_13554,N_14792);
nor U15771 (N_15771,N_13794,N_13518);
and U15772 (N_15772,N_14393,N_14480);
and U15773 (N_15773,N_13806,N_14016);
and U15774 (N_15774,N_14205,N_13635);
xor U15775 (N_15775,N_13864,N_14886);
nand U15776 (N_15776,N_13623,N_13842);
or U15777 (N_15777,N_14704,N_14121);
nand U15778 (N_15778,N_14388,N_14585);
or U15779 (N_15779,N_14210,N_13983);
nand U15780 (N_15780,N_14042,N_13540);
xnor U15781 (N_15781,N_14319,N_14546);
nand U15782 (N_15782,N_14209,N_14288);
nand U15783 (N_15783,N_14557,N_14264);
or U15784 (N_15784,N_13894,N_13820);
nor U15785 (N_15785,N_13724,N_13556);
nand U15786 (N_15786,N_14789,N_13894);
and U15787 (N_15787,N_13681,N_14723);
xnor U15788 (N_15788,N_13814,N_14211);
nand U15789 (N_15789,N_14423,N_13661);
nand U15790 (N_15790,N_13574,N_14672);
and U15791 (N_15791,N_14470,N_14943);
and U15792 (N_15792,N_14737,N_13539);
or U15793 (N_15793,N_14947,N_14913);
xnor U15794 (N_15794,N_13724,N_14967);
and U15795 (N_15795,N_14529,N_14378);
and U15796 (N_15796,N_14708,N_14016);
nand U15797 (N_15797,N_14438,N_14172);
and U15798 (N_15798,N_14666,N_14910);
nor U15799 (N_15799,N_14577,N_13816);
or U15800 (N_15800,N_14931,N_14505);
xnor U15801 (N_15801,N_14192,N_14175);
nor U15802 (N_15802,N_14869,N_14142);
and U15803 (N_15803,N_14017,N_14014);
nor U15804 (N_15804,N_13717,N_13615);
and U15805 (N_15805,N_14013,N_13903);
or U15806 (N_15806,N_14686,N_13750);
nor U15807 (N_15807,N_14775,N_14652);
nand U15808 (N_15808,N_14708,N_13979);
xor U15809 (N_15809,N_14848,N_14184);
nor U15810 (N_15810,N_13884,N_14626);
and U15811 (N_15811,N_13722,N_14096);
nand U15812 (N_15812,N_14612,N_14537);
or U15813 (N_15813,N_14365,N_14122);
or U15814 (N_15814,N_13508,N_14762);
or U15815 (N_15815,N_14462,N_13722);
nor U15816 (N_15816,N_14901,N_13629);
nand U15817 (N_15817,N_14308,N_14769);
and U15818 (N_15818,N_13510,N_13631);
nand U15819 (N_15819,N_14387,N_14931);
xnor U15820 (N_15820,N_14435,N_14347);
or U15821 (N_15821,N_14802,N_13711);
nor U15822 (N_15822,N_14512,N_14109);
nand U15823 (N_15823,N_13520,N_14446);
or U15824 (N_15824,N_14611,N_14957);
xnor U15825 (N_15825,N_14960,N_13692);
or U15826 (N_15826,N_14304,N_13501);
and U15827 (N_15827,N_13613,N_14242);
xnor U15828 (N_15828,N_14944,N_14808);
nor U15829 (N_15829,N_14152,N_13655);
and U15830 (N_15830,N_14025,N_14238);
xnor U15831 (N_15831,N_13902,N_13694);
xnor U15832 (N_15832,N_14292,N_14910);
and U15833 (N_15833,N_13691,N_14928);
and U15834 (N_15834,N_14270,N_14574);
or U15835 (N_15835,N_14793,N_14014);
xnor U15836 (N_15836,N_14480,N_13621);
nor U15837 (N_15837,N_14094,N_14131);
and U15838 (N_15838,N_14468,N_14937);
or U15839 (N_15839,N_14280,N_13546);
nor U15840 (N_15840,N_13611,N_13825);
or U15841 (N_15841,N_14323,N_14349);
xor U15842 (N_15842,N_13587,N_14403);
and U15843 (N_15843,N_14701,N_14143);
nor U15844 (N_15844,N_14458,N_14238);
nor U15845 (N_15845,N_14378,N_14677);
nor U15846 (N_15846,N_14847,N_14485);
nor U15847 (N_15847,N_13994,N_14771);
nor U15848 (N_15848,N_14148,N_14152);
nand U15849 (N_15849,N_13785,N_14283);
nand U15850 (N_15850,N_13855,N_14771);
nand U15851 (N_15851,N_14567,N_13991);
and U15852 (N_15852,N_14113,N_13995);
and U15853 (N_15853,N_13810,N_14484);
xor U15854 (N_15854,N_14081,N_14311);
and U15855 (N_15855,N_14810,N_13617);
or U15856 (N_15856,N_14029,N_13681);
xor U15857 (N_15857,N_14735,N_14654);
nand U15858 (N_15858,N_13536,N_13655);
or U15859 (N_15859,N_14666,N_14148);
xnor U15860 (N_15860,N_13790,N_13864);
and U15861 (N_15861,N_14854,N_13745);
nand U15862 (N_15862,N_14685,N_13773);
nand U15863 (N_15863,N_13837,N_14898);
xor U15864 (N_15864,N_14748,N_13633);
xnor U15865 (N_15865,N_14222,N_14624);
xnor U15866 (N_15866,N_14766,N_14795);
nor U15867 (N_15867,N_14325,N_14575);
nand U15868 (N_15868,N_14062,N_14903);
nand U15869 (N_15869,N_13838,N_14202);
xor U15870 (N_15870,N_14093,N_14744);
xor U15871 (N_15871,N_14919,N_14178);
nand U15872 (N_15872,N_14061,N_14686);
and U15873 (N_15873,N_13528,N_14934);
nor U15874 (N_15874,N_13945,N_13814);
and U15875 (N_15875,N_14116,N_13927);
or U15876 (N_15876,N_13979,N_14995);
nand U15877 (N_15877,N_14138,N_13805);
nor U15878 (N_15878,N_14155,N_13532);
and U15879 (N_15879,N_14466,N_14209);
and U15880 (N_15880,N_14463,N_13801);
nor U15881 (N_15881,N_13671,N_13753);
xnor U15882 (N_15882,N_13595,N_14065);
nand U15883 (N_15883,N_13731,N_13843);
nand U15884 (N_15884,N_13548,N_14597);
or U15885 (N_15885,N_13724,N_13769);
nand U15886 (N_15886,N_13982,N_14177);
or U15887 (N_15887,N_14362,N_14155);
and U15888 (N_15888,N_13898,N_14982);
nand U15889 (N_15889,N_13660,N_14560);
and U15890 (N_15890,N_13854,N_14880);
or U15891 (N_15891,N_14171,N_14304);
nand U15892 (N_15892,N_14516,N_14956);
nand U15893 (N_15893,N_14903,N_14633);
xor U15894 (N_15894,N_13680,N_14634);
nor U15895 (N_15895,N_14108,N_14313);
nand U15896 (N_15896,N_14319,N_13911);
nand U15897 (N_15897,N_13516,N_13930);
or U15898 (N_15898,N_13635,N_14388);
xnor U15899 (N_15899,N_13563,N_14373);
xor U15900 (N_15900,N_14620,N_14455);
nor U15901 (N_15901,N_14299,N_13583);
nor U15902 (N_15902,N_14504,N_14762);
nor U15903 (N_15903,N_14238,N_14094);
xor U15904 (N_15904,N_13765,N_14142);
nand U15905 (N_15905,N_14206,N_14878);
and U15906 (N_15906,N_14353,N_14243);
nor U15907 (N_15907,N_14126,N_14621);
or U15908 (N_15908,N_14199,N_14304);
nand U15909 (N_15909,N_14889,N_14855);
and U15910 (N_15910,N_14626,N_14562);
nand U15911 (N_15911,N_13517,N_14279);
xor U15912 (N_15912,N_14097,N_14966);
and U15913 (N_15913,N_14883,N_14983);
nor U15914 (N_15914,N_14822,N_14294);
or U15915 (N_15915,N_14292,N_14359);
nand U15916 (N_15916,N_14299,N_14800);
nand U15917 (N_15917,N_14538,N_14896);
xor U15918 (N_15918,N_14243,N_13655);
nand U15919 (N_15919,N_14397,N_13628);
or U15920 (N_15920,N_14315,N_14092);
xor U15921 (N_15921,N_14266,N_14620);
and U15922 (N_15922,N_14522,N_14166);
and U15923 (N_15923,N_14726,N_14700);
nand U15924 (N_15924,N_13850,N_14517);
and U15925 (N_15925,N_14085,N_13682);
and U15926 (N_15926,N_14383,N_14372);
xor U15927 (N_15927,N_14239,N_14005);
or U15928 (N_15928,N_13682,N_14163);
nor U15929 (N_15929,N_13817,N_14392);
nand U15930 (N_15930,N_14312,N_14223);
nor U15931 (N_15931,N_14347,N_14621);
nand U15932 (N_15932,N_14890,N_14448);
or U15933 (N_15933,N_14599,N_13687);
or U15934 (N_15934,N_13621,N_14336);
xnor U15935 (N_15935,N_14994,N_13820);
nor U15936 (N_15936,N_14842,N_14767);
or U15937 (N_15937,N_14059,N_14948);
xor U15938 (N_15938,N_14186,N_13950);
nor U15939 (N_15939,N_13926,N_13600);
nor U15940 (N_15940,N_14544,N_13517);
nor U15941 (N_15941,N_13938,N_14855);
nor U15942 (N_15942,N_14907,N_14463);
or U15943 (N_15943,N_14183,N_13933);
or U15944 (N_15944,N_14772,N_13635);
nand U15945 (N_15945,N_14934,N_14138);
and U15946 (N_15946,N_13559,N_13698);
xor U15947 (N_15947,N_14338,N_14287);
xnor U15948 (N_15948,N_13765,N_13842);
nand U15949 (N_15949,N_13513,N_13717);
and U15950 (N_15950,N_14600,N_14011);
xnor U15951 (N_15951,N_14837,N_13909);
or U15952 (N_15952,N_13678,N_13912);
or U15953 (N_15953,N_14817,N_14108);
nor U15954 (N_15954,N_14175,N_14675);
xnor U15955 (N_15955,N_13563,N_14668);
nand U15956 (N_15956,N_13885,N_14523);
nor U15957 (N_15957,N_14240,N_14241);
nand U15958 (N_15958,N_13652,N_13538);
nand U15959 (N_15959,N_14241,N_14046);
nand U15960 (N_15960,N_14275,N_14055);
xnor U15961 (N_15961,N_14319,N_14872);
nand U15962 (N_15962,N_13682,N_13980);
and U15963 (N_15963,N_13706,N_13608);
xor U15964 (N_15964,N_14056,N_13654);
or U15965 (N_15965,N_14814,N_14700);
or U15966 (N_15966,N_13583,N_14335);
xnor U15967 (N_15967,N_14292,N_14696);
or U15968 (N_15968,N_13743,N_13545);
nor U15969 (N_15969,N_13558,N_14338);
nand U15970 (N_15970,N_13902,N_14439);
nand U15971 (N_15971,N_14551,N_14211);
nand U15972 (N_15972,N_14552,N_14553);
xnor U15973 (N_15973,N_13991,N_13918);
or U15974 (N_15974,N_14040,N_13838);
nor U15975 (N_15975,N_14537,N_14623);
or U15976 (N_15976,N_14079,N_14266);
xor U15977 (N_15977,N_14857,N_13590);
xnor U15978 (N_15978,N_13590,N_14081);
nand U15979 (N_15979,N_14695,N_13642);
or U15980 (N_15980,N_14393,N_14565);
or U15981 (N_15981,N_13792,N_13715);
nand U15982 (N_15982,N_13621,N_14214);
or U15983 (N_15983,N_14481,N_13602);
or U15984 (N_15984,N_14882,N_14472);
and U15985 (N_15985,N_14048,N_13511);
or U15986 (N_15986,N_14066,N_14791);
and U15987 (N_15987,N_13860,N_14193);
and U15988 (N_15988,N_14757,N_14024);
xnor U15989 (N_15989,N_13544,N_14096);
nor U15990 (N_15990,N_14647,N_14371);
nor U15991 (N_15991,N_14660,N_13820);
nor U15992 (N_15992,N_14817,N_13654);
or U15993 (N_15993,N_14951,N_13514);
xor U15994 (N_15994,N_14804,N_13759);
xnor U15995 (N_15995,N_13615,N_14339);
or U15996 (N_15996,N_14934,N_14367);
and U15997 (N_15997,N_13892,N_14633);
nand U15998 (N_15998,N_14291,N_14555);
nor U15999 (N_15999,N_13879,N_14345);
nand U16000 (N_16000,N_14208,N_14504);
or U16001 (N_16001,N_14154,N_14684);
nor U16002 (N_16002,N_14447,N_14886);
nand U16003 (N_16003,N_13972,N_14353);
nand U16004 (N_16004,N_13837,N_13962);
or U16005 (N_16005,N_14879,N_14558);
xnor U16006 (N_16006,N_14322,N_13900);
and U16007 (N_16007,N_13800,N_13776);
nand U16008 (N_16008,N_14385,N_14521);
and U16009 (N_16009,N_14812,N_14587);
nand U16010 (N_16010,N_13629,N_14918);
nand U16011 (N_16011,N_14466,N_14223);
or U16012 (N_16012,N_13876,N_13878);
xnor U16013 (N_16013,N_13923,N_14913);
nor U16014 (N_16014,N_14740,N_13616);
and U16015 (N_16015,N_14077,N_14668);
xnor U16016 (N_16016,N_14783,N_14920);
and U16017 (N_16017,N_13659,N_13690);
nor U16018 (N_16018,N_14142,N_14847);
xor U16019 (N_16019,N_14437,N_13855);
and U16020 (N_16020,N_14952,N_14898);
nor U16021 (N_16021,N_14067,N_13996);
nor U16022 (N_16022,N_13693,N_14497);
xor U16023 (N_16023,N_13781,N_14607);
nor U16024 (N_16024,N_14237,N_14833);
nor U16025 (N_16025,N_13530,N_14685);
xnor U16026 (N_16026,N_14733,N_13938);
or U16027 (N_16027,N_14334,N_14372);
or U16028 (N_16028,N_13977,N_13677);
nor U16029 (N_16029,N_14752,N_14720);
and U16030 (N_16030,N_14251,N_14217);
and U16031 (N_16031,N_14280,N_13918);
or U16032 (N_16032,N_14238,N_14483);
nor U16033 (N_16033,N_14195,N_14508);
nor U16034 (N_16034,N_13647,N_14028);
and U16035 (N_16035,N_14024,N_14404);
nand U16036 (N_16036,N_14967,N_14782);
xnor U16037 (N_16037,N_14585,N_14517);
or U16038 (N_16038,N_14614,N_14310);
and U16039 (N_16039,N_13866,N_14495);
nor U16040 (N_16040,N_14733,N_13910);
nor U16041 (N_16041,N_14295,N_13883);
and U16042 (N_16042,N_14069,N_14189);
and U16043 (N_16043,N_14420,N_13688);
nand U16044 (N_16044,N_14322,N_14834);
or U16045 (N_16045,N_14486,N_14229);
nor U16046 (N_16046,N_14774,N_14798);
nor U16047 (N_16047,N_13717,N_13584);
nand U16048 (N_16048,N_14131,N_14458);
nand U16049 (N_16049,N_13769,N_14065);
and U16050 (N_16050,N_14963,N_14161);
and U16051 (N_16051,N_14066,N_14221);
xnor U16052 (N_16052,N_14779,N_13967);
or U16053 (N_16053,N_14086,N_13756);
and U16054 (N_16054,N_13581,N_14335);
or U16055 (N_16055,N_14447,N_14213);
nand U16056 (N_16056,N_13833,N_14959);
xor U16057 (N_16057,N_14479,N_14277);
xnor U16058 (N_16058,N_14511,N_14146);
or U16059 (N_16059,N_13648,N_14269);
nand U16060 (N_16060,N_14742,N_14886);
xnor U16061 (N_16061,N_14485,N_13943);
xnor U16062 (N_16062,N_14413,N_14282);
nand U16063 (N_16063,N_14747,N_14318);
nor U16064 (N_16064,N_13528,N_14246);
nand U16065 (N_16065,N_14156,N_13599);
or U16066 (N_16066,N_14108,N_14018);
xnor U16067 (N_16067,N_14847,N_13571);
and U16068 (N_16068,N_14324,N_14968);
xor U16069 (N_16069,N_14092,N_14053);
and U16070 (N_16070,N_14944,N_14061);
nand U16071 (N_16071,N_13888,N_14888);
and U16072 (N_16072,N_13775,N_14839);
xor U16073 (N_16073,N_14327,N_14749);
nand U16074 (N_16074,N_13533,N_13503);
or U16075 (N_16075,N_13665,N_14286);
xor U16076 (N_16076,N_14635,N_13965);
or U16077 (N_16077,N_14264,N_13579);
and U16078 (N_16078,N_14807,N_14586);
nand U16079 (N_16079,N_13986,N_13711);
xnor U16080 (N_16080,N_14222,N_14035);
and U16081 (N_16081,N_14083,N_13980);
nor U16082 (N_16082,N_14414,N_14015);
or U16083 (N_16083,N_14208,N_13949);
or U16084 (N_16084,N_13784,N_14667);
xnor U16085 (N_16085,N_14021,N_13503);
or U16086 (N_16086,N_14998,N_13570);
nor U16087 (N_16087,N_14221,N_14627);
xnor U16088 (N_16088,N_14796,N_14704);
or U16089 (N_16089,N_14097,N_13880);
nand U16090 (N_16090,N_14060,N_14803);
and U16091 (N_16091,N_14098,N_14199);
xnor U16092 (N_16092,N_14750,N_14514);
and U16093 (N_16093,N_14839,N_14425);
and U16094 (N_16094,N_14803,N_14154);
and U16095 (N_16095,N_13710,N_13615);
nor U16096 (N_16096,N_14258,N_13612);
nor U16097 (N_16097,N_14648,N_13654);
or U16098 (N_16098,N_13647,N_14679);
nand U16099 (N_16099,N_13926,N_13954);
nand U16100 (N_16100,N_14981,N_14256);
xor U16101 (N_16101,N_13943,N_13557);
nor U16102 (N_16102,N_14525,N_14809);
xnor U16103 (N_16103,N_13895,N_14868);
nor U16104 (N_16104,N_14379,N_14788);
xnor U16105 (N_16105,N_14859,N_13975);
nand U16106 (N_16106,N_14726,N_14163);
nand U16107 (N_16107,N_13726,N_13505);
nor U16108 (N_16108,N_14014,N_14891);
nor U16109 (N_16109,N_13565,N_14776);
or U16110 (N_16110,N_13723,N_14631);
xnor U16111 (N_16111,N_14274,N_14052);
or U16112 (N_16112,N_14731,N_13522);
nor U16113 (N_16113,N_14928,N_14802);
and U16114 (N_16114,N_14703,N_14378);
or U16115 (N_16115,N_13642,N_14924);
xor U16116 (N_16116,N_14914,N_13798);
and U16117 (N_16117,N_14256,N_14244);
xor U16118 (N_16118,N_14123,N_14587);
nor U16119 (N_16119,N_14361,N_13526);
nor U16120 (N_16120,N_14165,N_14966);
or U16121 (N_16121,N_13510,N_14687);
or U16122 (N_16122,N_13953,N_14254);
nor U16123 (N_16123,N_14187,N_13884);
or U16124 (N_16124,N_14580,N_13678);
xnor U16125 (N_16125,N_14923,N_14446);
or U16126 (N_16126,N_14669,N_13937);
xnor U16127 (N_16127,N_14417,N_13849);
nand U16128 (N_16128,N_14319,N_14300);
xor U16129 (N_16129,N_14465,N_14215);
or U16130 (N_16130,N_13810,N_14637);
or U16131 (N_16131,N_14621,N_14470);
or U16132 (N_16132,N_14537,N_14889);
xnor U16133 (N_16133,N_14238,N_14897);
and U16134 (N_16134,N_13888,N_13813);
xor U16135 (N_16135,N_14894,N_14227);
nor U16136 (N_16136,N_14894,N_13927);
nand U16137 (N_16137,N_13595,N_13734);
nor U16138 (N_16138,N_14582,N_13657);
nand U16139 (N_16139,N_13942,N_14767);
or U16140 (N_16140,N_14108,N_13688);
and U16141 (N_16141,N_14879,N_13728);
or U16142 (N_16142,N_14909,N_13559);
nor U16143 (N_16143,N_14136,N_13996);
xor U16144 (N_16144,N_13771,N_13676);
or U16145 (N_16145,N_14832,N_14086);
nor U16146 (N_16146,N_13538,N_14779);
and U16147 (N_16147,N_13836,N_14981);
nand U16148 (N_16148,N_14396,N_13654);
nor U16149 (N_16149,N_14830,N_13982);
nor U16150 (N_16150,N_13732,N_14213);
or U16151 (N_16151,N_13690,N_13737);
xnor U16152 (N_16152,N_14299,N_14498);
nor U16153 (N_16153,N_14936,N_14239);
xor U16154 (N_16154,N_13565,N_14354);
nand U16155 (N_16155,N_14474,N_14450);
nand U16156 (N_16156,N_14280,N_13524);
xnor U16157 (N_16157,N_14971,N_13586);
nor U16158 (N_16158,N_14887,N_14824);
and U16159 (N_16159,N_14115,N_13933);
or U16160 (N_16160,N_14477,N_13853);
or U16161 (N_16161,N_14753,N_14339);
xor U16162 (N_16162,N_14689,N_14535);
nor U16163 (N_16163,N_13541,N_14389);
nor U16164 (N_16164,N_14833,N_14945);
nand U16165 (N_16165,N_14097,N_13833);
xnor U16166 (N_16166,N_14733,N_14440);
xnor U16167 (N_16167,N_14032,N_14861);
nand U16168 (N_16168,N_13870,N_14214);
xnor U16169 (N_16169,N_14226,N_13878);
and U16170 (N_16170,N_14581,N_13855);
or U16171 (N_16171,N_13638,N_14146);
or U16172 (N_16172,N_14517,N_13807);
nand U16173 (N_16173,N_14433,N_14976);
nor U16174 (N_16174,N_13918,N_14192);
or U16175 (N_16175,N_14163,N_14916);
nand U16176 (N_16176,N_13751,N_14280);
nand U16177 (N_16177,N_14676,N_14118);
nor U16178 (N_16178,N_14310,N_13988);
nand U16179 (N_16179,N_14133,N_13711);
nand U16180 (N_16180,N_14841,N_13773);
or U16181 (N_16181,N_13564,N_14436);
or U16182 (N_16182,N_14089,N_14368);
nand U16183 (N_16183,N_14664,N_14140);
and U16184 (N_16184,N_14770,N_14881);
xnor U16185 (N_16185,N_14289,N_14380);
nand U16186 (N_16186,N_13899,N_13896);
and U16187 (N_16187,N_14569,N_14171);
xnor U16188 (N_16188,N_14985,N_13825);
or U16189 (N_16189,N_13590,N_13844);
and U16190 (N_16190,N_14856,N_14229);
and U16191 (N_16191,N_14711,N_14282);
xor U16192 (N_16192,N_14264,N_14207);
or U16193 (N_16193,N_14328,N_14054);
nand U16194 (N_16194,N_13935,N_14746);
xor U16195 (N_16195,N_14250,N_14471);
and U16196 (N_16196,N_14786,N_14059);
nor U16197 (N_16197,N_14188,N_14958);
nand U16198 (N_16198,N_14573,N_13506);
and U16199 (N_16199,N_14729,N_14610);
nand U16200 (N_16200,N_13916,N_14757);
nor U16201 (N_16201,N_14252,N_14669);
or U16202 (N_16202,N_13922,N_14264);
and U16203 (N_16203,N_14686,N_14578);
xor U16204 (N_16204,N_14108,N_13969);
xnor U16205 (N_16205,N_13936,N_13679);
or U16206 (N_16206,N_14169,N_14433);
or U16207 (N_16207,N_13646,N_14836);
xnor U16208 (N_16208,N_14341,N_14034);
or U16209 (N_16209,N_13711,N_13821);
nand U16210 (N_16210,N_13999,N_13936);
xnor U16211 (N_16211,N_14311,N_13881);
nor U16212 (N_16212,N_13978,N_14260);
or U16213 (N_16213,N_14628,N_14168);
xnor U16214 (N_16214,N_14197,N_14656);
and U16215 (N_16215,N_13712,N_14513);
nand U16216 (N_16216,N_14646,N_14223);
and U16217 (N_16217,N_13525,N_13978);
or U16218 (N_16218,N_14083,N_13905);
and U16219 (N_16219,N_13754,N_13932);
or U16220 (N_16220,N_14243,N_14722);
nand U16221 (N_16221,N_13681,N_14260);
nor U16222 (N_16222,N_14594,N_14194);
or U16223 (N_16223,N_13710,N_14497);
or U16224 (N_16224,N_14594,N_14946);
xnor U16225 (N_16225,N_13757,N_13670);
nor U16226 (N_16226,N_13801,N_14997);
nand U16227 (N_16227,N_14069,N_13548);
and U16228 (N_16228,N_14120,N_14622);
nor U16229 (N_16229,N_14830,N_14860);
or U16230 (N_16230,N_14994,N_14415);
nand U16231 (N_16231,N_14766,N_14617);
nand U16232 (N_16232,N_13735,N_14608);
xnor U16233 (N_16233,N_14874,N_14997);
xnor U16234 (N_16234,N_14869,N_14677);
and U16235 (N_16235,N_14975,N_14863);
nand U16236 (N_16236,N_14730,N_14993);
xor U16237 (N_16237,N_14579,N_13613);
or U16238 (N_16238,N_13994,N_14321);
nand U16239 (N_16239,N_13639,N_14600);
xnor U16240 (N_16240,N_14372,N_14958);
xor U16241 (N_16241,N_14144,N_14564);
or U16242 (N_16242,N_14112,N_14113);
or U16243 (N_16243,N_13679,N_14899);
nor U16244 (N_16244,N_14391,N_14829);
or U16245 (N_16245,N_14718,N_14687);
and U16246 (N_16246,N_14361,N_14477);
or U16247 (N_16247,N_13905,N_13639);
or U16248 (N_16248,N_14538,N_14961);
and U16249 (N_16249,N_14787,N_13908);
nand U16250 (N_16250,N_13665,N_14574);
or U16251 (N_16251,N_14649,N_14547);
xor U16252 (N_16252,N_14671,N_13571);
nor U16253 (N_16253,N_13834,N_14823);
xnor U16254 (N_16254,N_14714,N_14676);
xnor U16255 (N_16255,N_14418,N_14484);
and U16256 (N_16256,N_14824,N_13780);
xnor U16257 (N_16257,N_14822,N_14422);
or U16258 (N_16258,N_13960,N_14371);
nand U16259 (N_16259,N_14476,N_14348);
xnor U16260 (N_16260,N_14474,N_14904);
xnor U16261 (N_16261,N_13662,N_14467);
xnor U16262 (N_16262,N_14927,N_13876);
or U16263 (N_16263,N_14775,N_14114);
nor U16264 (N_16264,N_14337,N_14656);
or U16265 (N_16265,N_14828,N_14856);
or U16266 (N_16266,N_13817,N_14514);
xnor U16267 (N_16267,N_14411,N_14020);
nor U16268 (N_16268,N_14566,N_13555);
or U16269 (N_16269,N_13622,N_14282);
nand U16270 (N_16270,N_14316,N_14494);
nand U16271 (N_16271,N_13506,N_13671);
xor U16272 (N_16272,N_13528,N_14967);
xnor U16273 (N_16273,N_13879,N_13736);
xnor U16274 (N_16274,N_14473,N_13656);
or U16275 (N_16275,N_13831,N_14244);
and U16276 (N_16276,N_13823,N_14151);
or U16277 (N_16277,N_13542,N_14940);
xor U16278 (N_16278,N_13582,N_14941);
and U16279 (N_16279,N_14086,N_14010);
nand U16280 (N_16280,N_14689,N_14041);
nand U16281 (N_16281,N_13975,N_14930);
or U16282 (N_16282,N_14328,N_14742);
nand U16283 (N_16283,N_14359,N_13967);
nand U16284 (N_16284,N_14600,N_14062);
and U16285 (N_16285,N_13930,N_13829);
nand U16286 (N_16286,N_14930,N_14676);
nor U16287 (N_16287,N_14286,N_14780);
and U16288 (N_16288,N_14158,N_14272);
nand U16289 (N_16289,N_13762,N_14726);
nor U16290 (N_16290,N_14315,N_14672);
xor U16291 (N_16291,N_13807,N_13688);
nor U16292 (N_16292,N_14538,N_14136);
nor U16293 (N_16293,N_14447,N_13818);
and U16294 (N_16294,N_14587,N_14521);
or U16295 (N_16295,N_13881,N_13646);
nand U16296 (N_16296,N_13754,N_13885);
and U16297 (N_16297,N_13563,N_13954);
nor U16298 (N_16298,N_13915,N_14746);
nor U16299 (N_16299,N_13523,N_14586);
or U16300 (N_16300,N_14201,N_14867);
and U16301 (N_16301,N_14857,N_13949);
xnor U16302 (N_16302,N_14866,N_14320);
or U16303 (N_16303,N_13642,N_13904);
or U16304 (N_16304,N_14373,N_14659);
or U16305 (N_16305,N_14557,N_13768);
nand U16306 (N_16306,N_14074,N_14171);
nand U16307 (N_16307,N_13753,N_14798);
and U16308 (N_16308,N_14094,N_13608);
or U16309 (N_16309,N_14770,N_14908);
nand U16310 (N_16310,N_13881,N_13544);
nor U16311 (N_16311,N_14701,N_14538);
nand U16312 (N_16312,N_14717,N_14536);
nor U16313 (N_16313,N_14531,N_14703);
nand U16314 (N_16314,N_14792,N_14242);
or U16315 (N_16315,N_13926,N_14323);
xor U16316 (N_16316,N_14664,N_13822);
or U16317 (N_16317,N_13727,N_14736);
and U16318 (N_16318,N_14044,N_13664);
nor U16319 (N_16319,N_14132,N_13550);
xnor U16320 (N_16320,N_13927,N_14864);
and U16321 (N_16321,N_14955,N_14233);
nor U16322 (N_16322,N_13877,N_14143);
nand U16323 (N_16323,N_13744,N_14752);
nand U16324 (N_16324,N_13626,N_13681);
nor U16325 (N_16325,N_13838,N_13574);
nand U16326 (N_16326,N_14433,N_14251);
nand U16327 (N_16327,N_14327,N_14280);
and U16328 (N_16328,N_14762,N_13687);
or U16329 (N_16329,N_13614,N_14668);
xnor U16330 (N_16330,N_13763,N_13690);
nand U16331 (N_16331,N_14849,N_14280);
nand U16332 (N_16332,N_14688,N_13525);
or U16333 (N_16333,N_13508,N_14239);
and U16334 (N_16334,N_13532,N_13961);
nor U16335 (N_16335,N_13599,N_13718);
nand U16336 (N_16336,N_14163,N_14908);
nand U16337 (N_16337,N_14523,N_14744);
xnor U16338 (N_16338,N_13572,N_14783);
nor U16339 (N_16339,N_14169,N_14045);
and U16340 (N_16340,N_14505,N_13801);
xnor U16341 (N_16341,N_14782,N_14416);
xor U16342 (N_16342,N_14861,N_14116);
nor U16343 (N_16343,N_14273,N_13928);
xnor U16344 (N_16344,N_13727,N_14659);
or U16345 (N_16345,N_14850,N_14021);
or U16346 (N_16346,N_13815,N_14904);
nand U16347 (N_16347,N_14514,N_14347);
nor U16348 (N_16348,N_13945,N_13562);
or U16349 (N_16349,N_14805,N_14410);
nand U16350 (N_16350,N_14473,N_14831);
xor U16351 (N_16351,N_14741,N_14505);
nor U16352 (N_16352,N_14442,N_14549);
or U16353 (N_16353,N_14349,N_14056);
nand U16354 (N_16354,N_14598,N_13903);
nor U16355 (N_16355,N_13641,N_13766);
nand U16356 (N_16356,N_14972,N_14607);
nor U16357 (N_16357,N_14485,N_14346);
nor U16358 (N_16358,N_14816,N_14526);
xnor U16359 (N_16359,N_14784,N_13929);
nand U16360 (N_16360,N_13719,N_13818);
xnor U16361 (N_16361,N_14185,N_13938);
nand U16362 (N_16362,N_13878,N_14083);
nand U16363 (N_16363,N_14865,N_14488);
or U16364 (N_16364,N_13952,N_14596);
nand U16365 (N_16365,N_13884,N_13804);
or U16366 (N_16366,N_14178,N_13532);
and U16367 (N_16367,N_14655,N_14691);
or U16368 (N_16368,N_14018,N_14857);
or U16369 (N_16369,N_14088,N_14901);
and U16370 (N_16370,N_14881,N_14095);
nor U16371 (N_16371,N_14821,N_13554);
xor U16372 (N_16372,N_14167,N_13559);
nor U16373 (N_16373,N_13688,N_14318);
xnor U16374 (N_16374,N_14459,N_13904);
xor U16375 (N_16375,N_14658,N_14151);
and U16376 (N_16376,N_14033,N_14359);
nor U16377 (N_16377,N_14856,N_14568);
or U16378 (N_16378,N_13517,N_13747);
or U16379 (N_16379,N_13733,N_13883);
xnor U16380 (N_16380,N_14354,N_14707);
xor U16381 (N_16381,N_14468,N_13797);
nor U16382 (N_16382,N_14262,N_14114);
nand U16383 (N_16383,N_14953,N_14464);
xor U16384 (N_16384,N_13546,N_13555);
and U16385 (N_16385,N_14875,N_14445);
or U16386 (N_16386,N_14291,N_14233);
or U16387 (N_16387,N_14270,N_14036);
xor U16388 (N_16388,N_14099,N_13678);
or U16389 (N_16389,N_14007,N_14071);
xor U16390 (N_16390,N_13864,N_14869);
nand U16391 (N_16391,N_14027,N_14907);
xnor U16392 (N_16392,N_14729,N_13682);
nand U16393 (N_16393,N_13615,N_14965);
xnor U16394 (N_16394,N_14161,N_14788);
nand U16395 (N_16395,N_13794,N_14910);
xnor U16396 (N_16396,N_14660,N_14852);
or U16397 (N_16397,N_14129,N_13874);
nand U16398 (N_16398,N_14883,N_14011);
and U16399 (N_16399,N_13741,N_13848);
xnor U16400 (N_16400,N_14239,N_14692);
xor U16401 (N_16401,N_14984,N_13726);
and U16402 (N_16402,N_13777,N_14867);
or U16403 (N_16403,N_13611,N_14174);
and U16404 (N_16404,N_14955,N_14868);
or U16405 (N_16405,N_14608,N_13940);
xnor U16406 (N_16406,N_14718,N_14970);
nand U16407 (N_16407,N_13772,N_14847);
nor U16408 (N_16408,N_14433,N_14557);
nand U16409 (N_16409,N_14467,N_13843);
and U16410 (N_16410,N_13801,N_14460);
and U16411 (N_16411,N_14788,N_13712);
and U16412 (N_16412,N_14291,N_13626);
xnor U16413 (N_16413,N_13548,N_14255);
and U16414 (N_16414,N_14924,N_14796);
or U16415 (N_16415,N_14297,N_14188);
nor U16416 (N_16416,N_14557,N_14287);
and U16417 (N_16417,N_14250,N_14509);
nor U16418 (N_16418,N_13655,N_14807);
nand U16419 (N_16419,N_14672,N_13702);
nor U16420 (N_16420,N_14419,N_14159);
or U16421 (N_16421,N_13822,N_14843);
or U16422 (N_16422,N_14580,N_14983);
xnor U16423 (N_16423,N_14219,N_14257);
or U16424 (N_16424,N_14357,N_14359);
and U16425 (N_16425,N_13891,N_13745);
or U16426 (N_16426,N_14094,N_14182);
or U16427 (N_16427,N_14752,N_14343);
and U16428 (N_16428,N_13524,N_14955);
nand U16429 (N_16429,N_14231,N_14691);
nand U16430 (N_16430,N_13658,N_13909);
and U16431 (N_16431,N_14076,N_14995);
xor U16432 (N_16432,N_13738,N_13843);
nand U16433 (N_16433,N_14229,N_13718);
nand U16434 (N_16434,N_14875,N_13851);
or U16435 (N_16435,N_14985,N_13976);
xnor U16436 (N_16436,N_14465,N_14779);
xor U16437 (N_16437,N_14205,N_13577);
and U16438 (N_16438,N_14647,N_14164);
xnor U16439 (N_16439,N_14745,N_14271);
and U16440 (N_16440,N_14023,N_14536);
xor U16441 (N_16441,N_14695,N_14653);
nor U16442 (N_16442,N_14532,N_14031);
nor U16443 (N_16443,N_14482,N_14148);
xnor U16444 (N_16444,N_14194,N_13505);
nor U16445 (N_16445,N_13759,N_14068);
nor U16446 (N_16446,N_13919,N_13552);
or U16447 (N_16447,N_13894,N_13887);
nand U16448 (N_16448,N_13666,N_14663);
and U16449 (N_16449,N_13761,N_14071);
xor U16450 (N_16450,N_14043,N_13535);
xnor U16451 (N_16451,N_14194,N_14051);
and U16452 (N_16452,N_14724,N_13554);
nor U16453 (N_16453,N_14655,N_13515);
nand U16454 (N_16454,N_14544,N_14545);
or U16455 (N_16455,N_14201,N_13551);
nand U16456 (N_16456,N_13875,N_14315);
or U16457 (N_16457,N_13558,N_14230);
xnor U16458 (N_16458,N_14537,N_13550);
xor U16459 (N_16459,N_13649,N_14183);
nor U16460 (N_16460,N_14066,N_14252);
nor U16461 (N_16461,N_13673,N_14564);
or U16462 (N_16462,N_14542,N_14350);
xnor U16463 (N_16463,N_14808,N_14745);
or U16464 (N_16464,N_14535,N_14992);
or U16465 (N_16465,N_14017,N_13686);
or U16466 (N_16466,N_13841,N_14086);
and U16467 (N_16467,N_13798,N_14345);
or U16468 (N_16468,N_14736,N_14162);
nor U16469 (N_16469,N_14878,N_14500);
nand U16470 (N_16470,N_14948,N_14079);
nor U16471 (N_16471,N_14469,N_14875);
and U16472 (N_16472,N_14670,N_14706);
nand U16473 (N_16473,N_13876,N_14001);
nor U16474 (N_16474,N_14256,N_14778);
nand U16475 (N_16475,N_14166,N_14747);
nand U16476 (N_16476,N_13719,N_13866);
nand U16477 (N_16477,N_14074,N_14476);
or U16478 (N_16478,N_14938,N_14513);
or U16479 (N_16479,N_13527,N_14001);
nor U16480 (N_16480,N_14126,N_14981);
nand U16481 (N_16481,N_13931,N_13730);
xor U16482 (N_16482,N_13571,N_14167);
nand U16483 (N_16483,N_14832,N_13793);
xnor U16484 (N_16484,N_14159,N_14827);
or U16485 (N_16485,N_14802,N_13506);
nor U16486 (N_16486,N_13589,N_13756);
or U16487 (N_16487,N_14275,N_14854);
xor U16488 (N_16488,N_13949,N_13690);
nand U16489 (N_16489,N_14020,N_14859);
or U16490 (N_16490,N_13714,N_13569);
xnor U16491 (N_16491,N_14443,N_14947);
and U16492 (N_16492,N_14665,N_13579);
xor U16493 (N_16493,N_13536,N_13777);
and U16494 (N_16494,N_14025,N_14985);
nor U16495 (N_16495,N_14864,N_14017);
xor U16496 (N_16496,N_14567,N_13558);
nand U16497 (N_16497,N_14293,N_14084);
nand U16498 (N_16498,N_14984,N_13810);
nand U16499 (N_16499,N_14193,N_14255);
xnor U16500 (N_16500,N_15623,N_16105);
xnor U16501 (N_16501,N_15730,N_15009);
xor U16502 (N_16502,N_16046,N_15327);
nand U16503 (N_16503,N_15513,N_15966);
nand U16504 (N_16504,N_16477,N_15818);
xnor U16505 (N_16505,N_16069,N_15346);
nand U16506 (N_16506,N_15599,N_15900);
nand U16507 (N_16507,N_15469,N_16313);
xor U16508 (N_16508,N_15530,N_15662);
and U16509 (N_16509,N_16248,N_15988);
nand U16510 (N_16510,N_15452,N_15103);
nand U16511 (N_16511,N_15773,N_15203);
and U16512 (N_16512,N_16018,N_15028);
nor U16513 (N_16513,N_15932,N_15864);
or U16514 (N_16514,N_15952,N_15410);
and U16515 (N_16515,N_15618,N_15797);
and U16516 (N_16516,N_15057,N_16485);
and U16517 (N_16517,N_15369,N_15181);
and U16518 (N_16518,N_15584,N_15225);
xor U16519 (N_16519,N_16489,N_15881);
nor U16520 (N_16520,N_15617,N_15381);
or U16521 (N_16521,N_15986,N_15411);
nand U16522 (N_16522,N_15726,N_15373);
xor U16523 (N_16523,N_15575,N_15833);
nor U16524 (N_16524,N_15074,N_15206);
and U16525 (N_16525,N_15482,N_15859);
or U16526 (N_16526,N_15983,N_15012);
xor U16527 (N_16527,N_15837,N_15788);
xnor U16528 (N_16528,N_16093,N_15880);
nor U16529 (N_16529,N_16463,N_16049);
and U16530 (N_16530,N_16051,N_15865);
xnor U16531 (N_16531,N_15263,N_16307);
or U16532 (N_16532,N_15945,N_15685);
nand U16533 (N_16533,N_15613,N_15075);
and U16534 (N_16534,N_16487,N_15435);
xor U16535 (N_16535,N_15071,N_15349);
and U16536 (N_16536,N_16175,N_16262);
xnor U16537 (N_16537,N_15426,N_16382);
or U16538 (N_16538,N_15630,N_15389);
nor U16539 (N_16539,N_16261,N_16215);
and U16540 (N_16540,N_15669,N_15016);
nand U16541 (N_16541,N_15590,N_15271);
or U16542 (N_16542,N_15616,N_15388);
xor U16543 (N_16543,N_15468,N_16245);
or U16544 (N_16544,N_15596,N_15046);
or U16545 (N_16545,N_15425,N_15632);
nand U16546 (N_16546,N_16462,N_16232);
nand U16547 (N_16547,N_15387,N_15149);
xnor U16548 (N_16548,N_15417,N_15912);
or U16549 (N_16549,N_15278,N_16298);
nand U16550 (N_16550,N_16392,N_16317);
or U16551 (N_16551,N_15000,N_15519);
and U16552 (N_16552,N_15858,N_16324);
nand U16553 (N_16553,N_16475,N_16138);
and U16554 (N_16554,N_15884,N_15133);
xnor U16555 (N_16555,N_15649,N_15031);
nor U16556 (N_16556,N_15446,N_16383);
nand U16557 (N_16557,N_15922,N_15556);
and U16558 (N_16558,N_16476,N_16423);
nand U16559 (N_16559,N_16084,N_16001);
and U16560 (N_16560,N_16253,N_15476);
and U16561 (N_16561,N_15989,N_15041);
nand U16562 (N_16562,N_15154,N_15760);
and U16563 (N_16563,N_15115,N_15246);
and U16564 (N_16564,N_15363,N_16082);
nor U16565 (N_16565,N_15549,N_16243);
or U16566 (N_16566,N_16181,N_15241);
or U16567 (N_16567,N_15051,N_15238);
or U16568 (N_16568,N_16096,N_16086);
nand U16569 (N_16569,N_16499,N_15412);
xnor U16570 (N_16570,N_15076,N_15847);
nor U16571 (N_16571,N_15113,N_15708);
nand U16572 (N_16572,N_15364,N_15734);
and U16573 (N_16573,N_15737,N_15130);
nand U16574 (N_16574,N_15689,N_15407);
or U16575 (N_16575,N_16179,N_16309);
and U16576 (N_16576,N_15215,N_15594);
or U16577 (N_16577,N_15368,N_16474);
or U16578 (N_16578,N_16202,N_15505);
and U16579 (N_16579,N_15904,N_16007);
and U16580 (N_16580,N_15905,N_15501);
nor U16581 (N_16581,N_15895,N_15370);
nor U16582 (N_16582,N_16268,N_15845);
nand U16583 (N_16583,N_16438,N_15933);
or U16584 (N_16584,N_16065,N_16155);
or U16585 (N_16585,N_16042,N_16210);
nor U16586 (N_16586,N_15072,N_16106);
nand U16587 (N_16587,N_16174,N_15047);
xor U16588 (N_16588,N_15844,N_15559);
and U16589 (N_16589,N_15699,N_15109);
or U16590 (N_16590,N_15896,N_16297);
xnor U16591 (N_16591,N_15860,N_15286);
and U16592 (N_16592,N_15261,N_15080);
xor U16593 (N_16593,N_16408,N_16095);
xnor U16594 (N_16594,N_16094,N_16368);
and U16595 (N_16595,N_16230,N_15420);
nand U16596 (N_16596,N_16184,N_15344);
nand U16597 (N_16597,N_15185,N_15258);
nand U16598 (N_16598,N_15114,N_15676);
or U16599 (N_16599,N_15638,N_16025);
xnor U16600 (N_16600,N_16244,N_15179);
and U16601 (N_16601,N_15715,N_15650);
nand U16602 (N_16602,N_15752,N_15729);
nand U16603 (N_16603,N_15867,N_16389);
nand U16604 (N_16604,N_15320,N_15897);
or U16605 (N_16605,N_16258,N_15621);
xor U16606 (N_16606,N_16347,N_15331);
or U16607 (N_16607,N_15520,N_15485);
and U16608 (N_16608,N_15529,N_15736);
nor U16609 (N_16609,N_15800,N_15902);
nand U16610 (N_16610,N_16342,N_16402);
and U16611 (N_16611,N_16461,N_16098);
or U16612 (N_16612,N_15776,N_16235);
nor U16613 (N_16613,N_15558,N_15637);
nand U16614 (N_16614,N_15068,N_16400);
or U16615 (N_16615,N_16306,N_15947);
or U16616 (N_16616,N_15043,N_16102);
nand U16617 (N_16617,N_15444,N_16172);
xnor U16618 (N_16618,N_15703,N_15307);
xnor U16619 (N_16619,N_16166,N_15913);
nand U16620 (N_16620,N_15088,N_15840);
or U16621 (N_16621,N_15438,N_15538);
and U16622 (N_16622,N_15508,N_16149);
and U16623 (N_16623,N_15005,N_15450);
nor U16624 (N_16624,N_16206,N_15570);
or U16625 (N_16625,N_16440,N_16439);
and U16626 (N_16626,N_16471,N_15832);
xnor U16627 (N_16627,N_16355,N_16087);
or U16628 (N_16628,N_15318,N_15159);
xor U16629 (N_16629,N_15757,N_15089);
nor U16630 (N_16630,N_16053,N_15661);
and U16631 (N_16631,N_15950,N_15394);
and U16632 (N_16632,N_15173,N_16110);
nand U16633 (N_16633,N_16050,N_15968);
xnor U16634 (N_16634,N_16331,N_16497);
and U16635 (N_16635,N_16020,N_16308);
and U16636 (N_16636,N_16249,N_15494);
and U16637 (N_16637,N_15144,N_15545);
nor U16638 (N_16638,N_15978,N_15402);
nand U16639 (N_16639,N_15082,N_15995);
nor U16640 (N_16640,N_15323,N_15775);
nor U16641 (N_16641,N_16144,N_15487);
and U16642 (N_16642,N_15316,N_16374);
and U16643 (N_16643,N_15150,N_15583);
and U16644 (N_16644,N_16256,N_16036);
and U16645 (N_16645,N_15062,N_15667);
xnor U16646 (N_16646,N_16335,N_15335);
nor U16647 (N_16647,N_16490,N_15595);
nor U16648 (N_16648,N_16254,N_15834);
and U16649 (N_16649,N_15121,N_16164);
xnor U16650 (N_16650,N_15248,N_16427);
xnor U16651 (N_16651,N_15714,N_15447);
or U16652 (N_16652,N_15112,N_15565);
nand U16653 (N_16653,N_16023,N_15798);
nor U16654 (N_16654,N_16178,N_15615);
xnor U16655 (N_16655,N_15522,N_16425);
nand U16656 (N_16656,N_15284,N_16109);
and U16657 (N_16657,N_16193,N_16078);
nor U16658 (N_16658,N_15517,N_16039);
xnor U16659 (N_16659,N_15213,N_16246);
xnor U16660 (N_16660,N_16449,N_15014);
nor U16661 (N_16661,N_15648,N_15564);
xor U16662 (N_16662,N_16472,N_15568);
nor U16663 (N_16663,N_16395,N_15518);
nor U16664 (N_16664,N_15674,N_16452);
xnor U16665 (N_16665,N_16371,N_15526);
nand U16666 (N_16666,N_16424,N_15682);
or U16667 (N_16667,N_15807,N_15531);
nand U16668 (N_16668,N_15610,N_15211);
nand U16669 (N_16669,N_16115,N_15537);
nand U16670 (N_16670,N_15756,N_15493);
nand U16671 (N_16671,N_15345,N_16219);
xnor U16672 (N_16672,N_16118,N_15955);
or U16673 (N_16673,N_15378,N_16085);
or U16674 (N_16674,N_15256,N_16220);
nor U16675 (N_16675,N_15941,N_16430);
xnor U16676 (N_16676,N_15162,N_16151);
and U16677 (N_16677,N_16296,N_15360);
nand U16678 (N_16678,N_16266,N_15108);
or U16679 (N_16679,N_16074,N_16072);
and U16680 (N_16680,N_15290,N_15557);
nand U16681 (N_16681,N_16458,N_15287);
xor U16682 (N_16682,N_15274,N_16008);
or U16683 (N_16683,N_15477,N_15755);
nor U16684 (N_16684,N_16337,N_15489);
or U16685 (N_16685,N_15145,N_16496);
or U16686 (N_16686,N_15790,N_15333);
or U16687 (N_16687,N_15392,N_15534);
or U16688 (N_16688,N_16136,N_15355);
nor U16689 (N_16689,N_16047,N_15742);
xor U16690 (N_16690,N_16121,N_15193);
and U16691 (N_16691,N_16414,N_16457);
or U16692 (N_16692,N_15939,N_16428);
and U16693 (N_16693,N_15500,N_15868);
xnor U16694 (N_16694,N_16429,N_15257);
nor U16695 (N_16695,N_16446,N_15111);
and U16696 (N_16696,N_16140,N_15045);
and U16697 (N_16697,N_15843,N_15754);
xnor U16698 (N_16698,N_15972,N_15021);
and U16699 (N_16699,N_15151,N_15190);
nand U16700 (N_16700,N_16068,N_16017);
and U16701 (N_16701,N_15107,N_16401);
nor U16702 (N_16702,N_15358,N_15740);
and U16703 (N_16703,N_16404,N_16290);
nand U16704 (N_16704,N_15971,N_15453);
nand U16705 (N_16705,N_15543,N_16279);
nor U16706 (N_16706,N_16029,N_16067);
or U16707 (N_16707,N_15391,N_15044);
xnor U16708 (N_16708,N_15455,N_15289);
nor U16709 (N_16709,N_15770,N_15901);
xor U16710 (N_16710,N_15208,N_15872);
nor U16711 (N_16711,N_16228,N_15054);
nand U16712 (N_16712,N_15786,N_16189);
nand U16713 (N_16713,N_16259,N_15242);
and U16714 (N_16714,N_15254,N_15930);
and U16715 (N_16715,N_15384,N_15496);
or U16716 (N_16716,N_15499,N_16070);
nor U16717 (N_16717,N_16344,N_15359);
xnor U16718 (N_16718,N_16080,N_16079);
nand U16719 (N_16719,N_15228,N_15914);
and U16720 (N_16720,N_15163,N_16165);
xnor U16721 (N_16721,N_15440,N_16183);
xnor U16722 (N_16722,N_15633,N_16146);
or U16723 (N_16723,N_15727,N_15343);
and U16724 (N_16724,N_15198,N_15970);
or U16725 (N_16725,N_16329,N_15116);
nor U16726 (N_16726,N_15507,N_15758);
nand U16727 (N_16727,N_15251,N_15092);
and U16728 (N_16728,N_16417,N_15723);
xnor U16729 (N_16729,N_16300,N_15684);
nor U16730 (N_16730,N_16168,N_15696);
and U16731 (N_16731,N_16208,N_16269);
xnor U16732 (N_16732,N_15294,N_16161);
nand U16733 (N_16733,N_15663,N_16294);
nand U16734 (N_16734,N_15999,N_16274);
and U16735 (N_16735,N_15183,N_15132);
and U16736 (N_16736,N_16407,N_16455);
and U16737 (N_16737,N_15361,N_15974);
nand U16738 (N_16738,N_15161,N_16469);
xor U16739 (N_16739,N_15552,N_15413);
nor U16740 (N_16740,N_15078,N_15953);
nor U16741 (N_16741,N_15958,N_15509);
nor U16742 (N_16742,N_15553,N_15229);
and U16743 (N_16743,N_16338,N_15069);
nor U16744 (N_16744,N_15996,N_15406);
nor U16745 (N_16745,N_15448,N_16024);
xnor U16746 (N_16746,N_15937,N_16000);
xor U16747 (N_16747,N_15470,N_16257);
or U16748 (N_16748,N_16104,N_15421);
and U16749 (N_16749,N_15460,N_15400);
and U16750 (N_16750,N_15659,N_15218);
or U16751 (N_16751,N_15017,N_16358);
xor U16752 (N_16752,N_15512,N_15525);
nor U16753 (N_16753,N_15184,N_15332);
or U16754 (N_16754,N_16169,N_15137);
nand U16755 (N_16755,N_15465,N_16247);
xnor U16756 (N_16756,N_15437,N_15015);
and U16757 (N_16757,N_16167,N_15611);
nor U16758 (N_16758,N_15140,N_16127);
xnor U16759 (N_16759,N_15677,N_15504);
or U16760 (N_16760,N_15772,N_16302);
or U16761 (N_16761,N_16340,N_16363);
xnor U16762 (N_16762,N_16479,N_15252);
and U16763 (N_16763,N_15027,N_16147);
nand U16764 (N_16764,N_15102,N_15510);
and U16765 (N_16765,N_15521,N_15502);
nor U16766 (N_16766,N_15093,N_15574);
or U16767 (N_16767,N_15820,N_16037);
xnor U16768 (N_16768,N_16375,N_16066);
or U16769 (N_16769,N_16227,N_16356);
nand U16770 (N_16770,N_15277,N_15805);
and U16771 (N_16771,N_15990,N_15227);
xnor U16772 (N_16772,N_16445,N_15516);
and U16773 (N_16773,N_15802,N_16460);
xor U16774 (N_16774,N_16378,N_16346);
and U16775 (N_16775,N_15224,N_16353);
nand U16776 (N_16776,N_16061,N_15281);
nand U16777 (N_16777,N_16216,N_16162);
nor U16778 (N_16778,N_16250,N_16453);
xnor U16779 (N_16779,N_15724,N_15835);
or U16780 (N_16780,N_16432,N_15276);
nand U16781 (N_16781,N_15812,N_15928);
nand U16782 (N_16782,N_15533,N_15657);
xor U16783 (N_16783,N_15329,N_15681);
nand U16784 (N_16784,N_16350,N_15809);
or U16785 (N_16785,N_16128,N_15924);
nand U16786 (N_16786,N_15993,N_15070);
xnor U16787 (N_16787,N_15925,N_15918);
nor U16788 (N_16788,N_16034,N_16191);
nand U16789 (N_16789,N_15831,N_16170);
nor U16790 (N_16790,N_16014,N_15602);
or U16791 (N_16791,N_15910,N_15886);
xor U16792 (N_16792,N_16071,N_15957);
nand U16793 (N_16793,N_15490,N_15003);
xnor U16794 (N_16794,N_15739,N_15334);
nand U16795 (N_16795,N_15182,N_15541);
and U16796 (N_16796,N_15687,N_16211);
nand U16797 (N_16797,N_16270,N_16077);
or U16798 (N_16798,N_15608,N_15239);
xnor U16799 (N_16799,N_15635,N_16122);
or U16800 (N_16800,N_15964,N_16101);
nand U16801 (N_16801,N_15087,N_16241);
and U16802 (N_16802,N_15780,N_16240);
and U16803 (N_16803,N_15707,N_15365);
and U16804 (N_16804,N_15055,N_15793);
nor U16805 (N_16805,N_15457,N_16311);
nand U16806 (N_16806,N_16099,N_16410);
nor U16807 (N_16807,N_15838,N_15328);
xnor U16808 (N_16808,N_15155,N_16495);
and U16809 (N_16809,N_15878,N_16040);
or U16810 (N_16810,N_15836,N_15824);
and U16811 (N_16811,N_15842,N_15486);
xnor U16812 (N_16812,N_15869,N_16376);
or U16813 (N_16813,N_15641,N_15295);
or U16814 (N_16814,N_15934,N_16030);
and U16815 (N_16815,N_15600,N_16081);
xnor U16816 (N_16816,N_15245,N_16433);
nor U16817 (N_16817,N_15819,N_15326);
and U16818 (N_16818,N_15168,N_16394);
nor U16819 (N_16819,N_15383,N_16285);
and U16820 (N_16820,N_15459,N_15769);
nand U16821 (N_16821,N_15419,N_15826);
or U16822 (N_16822,N_15624,N_15963);
nor U16823 (N_16823,N_16176,N_16027);
nand U16824 (N_16824,N_16016,N_16186);
or U16825 (N_16825,N_15985,N_15646);
nor U16826 (N_16826,N_16273,N_15273);
xnor U16827 (N_16827,N_15700,N_15704);
nor U16828 (N_16828,N_16359,N_16325);
nand U16829 (N_16829,N_15322,N_15375);
and U16830 (N_16830,N_15713,N_15298);
or U16831 (N_16831,N_16075,N_15603);
or U16832 (N_16832,N_16252,N_16332);
and U16833 (N_16833,N_15721,N_15299);
and U16834 (N_16834,N_15622,N_15305);
nand U16835 (N_16835,N_15550,N_16190);
and U16836 (N_16836,N_16205,N_15199);
and U16837 (N_16837,N_15866,N_15804);
or U16838 (N_16838,N_16203,N_16058);
and U16839 (N_16839,N_16237,N_16188);
and U16840 (N_16840,N_15965,N_15214);
or U16841 (N_16841,N_16013,N_15588);
and U16842 (N_16842,N_15170,N_16117);
xnor U16843 (N_16843,N_15207,N_15266);
nand U16844 (N_16844,N_16365,N_15692);
nor U16845 (N_16845,N_15100,N_15722);
or U16846 (N_16846,N_15546,N_16073);
nor U16847 (N_16847,N_15129,N_15023);
xnor U16848 (N_16848,N_15127,N_16343);
nand U16849 (N_16849,N_15982,N_16345);
nand U16850 (N_16850,N_15774,N_16141);
xnor U16851 (N_16851,N_15434,N_15167);
xnor U16852 (N_16852,N_15936,N_16187);
or U16853 (N_16853,N_15401,N_16009);
nor U16854 (N_16854,N_16207,N_15341);
and U16855 (N_16855,N_15451,N_16348);
nor U16856 (N_16856,N_16357,N_15589);
nor U16857 (N_16857,N_15441,N_16336);
xor U16858 (N_16858,N_15415,N_16278);
and U16859 (N_16859,N_15099,N_15551);
or U16860 (N_16860,N_16441,N_16492);
nor U16861 (N_16861,N_15422,N_15039);
nor U16862 (N_16862,N_16059,N_15377);
or U16863 (N_16863,N_15042,N_16366);
or U16864 (N_16864,N_15196,N_16015);
nand U16865 (N_16865,N_16021,N_16287);
nor U16866 (N_16866,N_15823,N_15429);
and U16867 (N_16867,N_16041,N_15815);
xor U16868 (N_16868,N_16354,N_16312);
and U16869 (N_16869,N_15883,N_15827);
nand U16870 (N_16870,N_15577,N_15861);
and U16871 (N_16871,N_15586,N_16131);
nand U16872 (N_16872,N_15956,N_16484);
nor U16873 (N_16873,N_15002,N_15313);
or U16874 (N_16874,N_15197,N_16396);
and U16875 (N_16875,N_15876,N_16139);
nor U16876 (N_16876,N_15171,N_15579);
or U16877 (N_16877,N_15702,N_16480);
and U16878 (N_16878,N_16421,N_15612);
nand U16879 (N_16879,N_16316,N_15338);
or U16880 (N_16880,N_15428,N_16416);
and U16881 (N_16881,N_15348,N_15119);
nand U16882 (N_16882,N_15857,N_15125);
and U16883 (N_16883,N_15711,N_15220);
xor U16884 (N_16884,N_15544,N_15506);
and U16885 (N_16885,N_15741,N_15732);
and U16886 (N_16886,N_16004,N_15097);
nor U16887 (N_16887,N_16043,N_15706);
xnor U16888 (N_16888,N_16114,N_15779);
or U16889 (N_16889,N_15572,N_16379);
xnor U16890 (N_16890,N_15073,N_15135);
xnor U16891 (N_16891,N_15454,N_15660);
nor U16892 (N_16892,N_15236,N_15718);
xnor U16893 (N_16893,N_15735,N_16134);
xnor U16894 (N_16894,N_15582,N_15157);
nor U16895 (N_16895,N_15795,N_16314);
or U16896 (N_16896,N_15743,N_16442);
xnor U16897 (N_16897,N_15614,N_15139);
and U16898 (N_16898,N_15853,N_15398);
xnor U16899 (N_16899,N_15024,N_15601);
nand U16900 (N_16900,N_15160,N_16434);
nor U16901 (N_16901,N_16163,N_16448);
or U16902 (N_16902,N_16217,N_15312);
or U16903 (N_16903,N_16288,N_15606);
or U16904 (N_16904,N_15124,N_15604);
and U16905 (N_16905,N_16238,N_16038);
and U16906 (N_16906,N_16156,N_16265);
or U16907 (N_16907,N_15644,N_15792);
nor U16908 (N_16908,N_16415,N_15018);
xnor U16909 (N_16909,N_15794,N_15656);
nand U16910 (N_16910,N_16411,N_15035);
and U16911 (N_16911,N_15688,N_16289);
and U16912 (N_16912,N_16204,N_15882);
nor U16913 (N_16913,N_15709,N_15423);
or U16914 (N_16914,N_16351,N_15466);
and U16915 (N_16915,N_16223,N_15464);
or U16916 (N_16916,N_15061,N_16054);
nor U16917 (N_16917,N_15973,N_15352);
nand U16918 (N_16918,N_15048,N_15849);
xnor U16919 (N_16919,N_15153,N_15156);
nor U16920 (N_16920,N_16470,N_15250);
and U16921 (N_16921,N_15719,N_16310);
nor U16922 (N_16922,N_16148,N_16035);
nor U16923 (N_16923,N_16224,N_15785);
and U16924 (N_16924,N_16291,N_15535);
nand U16925 (N_16925,N_16052,N_15488);
xor U16926 (N_16926,N_16133,N_16334);
xor U16927 (N_16927,N_15960,N_15580);
nand U16928 (N_16928,N_15008,N_15456);
xnor U16929 (N_16929,N_15079,N_15701);
xnor U16930 (N_16930,N_16242,N_15777);
or U16931 (N_16931,N_16456,N_15350);
xnor U16932 (N_16932,N_15306,N_15977);
xnor U16933 (N_16933,N_15554,N_16108);
and U16934 (N_16934,N_16192,N_15698);
nand U16935 (N_16935,N_15050,N_15462);
nand U16936 (N_16936,N_16126,N_16467);
nand U16937 (N_16937,N_15759,N_16003);
nor U16938 (N_16938,N_16280,N_16321);
xor U16939 (N_16939,N_16326,N_15458);
xnor U16940 (N_16940,N_15852,N_15767);
and U16941 (N_16941,N_16437,N_16319);
nor U16942 (N_16942,N_15569,N_15879);
or U16943 (N_16943,N_15848,N_16318);
or U16944 (N_16944,N_16177,N_15191);
and U16945 (N_16945,N_16234,N_16406);
xnor U16946 (N_16946,N_15483,N_16195);
xor U16947 (N_16947,N_16171,N_15480);
and U16948 (N_16948,N_15386,N_15146);
and U16949 (N_16949,N_16255,N_15059);
xor U16950 (N_16950,N_16137,N_15782);
nor U16951 (N_16951,N_16130,N_15060);
nand U16952 (N_16952,N_15110,N_16212);
and U16953 (N_16953,N_15762,N_16125);
or U16954 (N_16954,N_15309,N_16360);
and U16955 (N_16955,N_16493,N_15796);
nor U16956 (N_16956,N_15929,N_16180);
nor U16957 (N_16957,N_15347,N_16111);
or U16958 (N_16958,N_15766,N_15524);
nand U16959 (N_16959,N_16045,N_16391);
xnor U16960 (N_16960,N_15117,N_15143);
xor U16961 (N_16961,N_15268,N_16239);
nand U16962 (N_16962,N_16091,N_15065);
and U16963 (N_16963,N_15404,N_15926);
nand U16964 (N_16964,N_15673,N_16465);
and U16965 (N_16965,N_15189,N_16362);
and U16966 (N_16966,N_16390,N_15169);
xor U16967 (N_16967,N_15814,N_15372);
nand U16968 (N_16968,N_15176,N_15249);
nor U16969 (N_16969,N_16281,N_15025);
and U16970 (N_16970,N_15801,N_16483);
or U16971 (N_16971,N_15201,N_16158);
xnor U16972 (N_16972,N_15279,N_16129);
and U16973 (N_16973,N_15086,N_15651);
nand U16974 (N_16974,N_16494,N_15094);
xnor U16975 (N_16975,N_15562,N_15625);
nand U16976 (N_16976,N_16159,N_16263);
nand U16977 (N_16977,N_15272,N_16327);
or U16978 (N_16978,N_15104,N_16409);
and U16979 (N_16979,N_15056,N_15136);
nand U16980 (N_16980,N_16222,N_15037);
or U16981 (N_16981,N_15026,N_16473);
nand U16982 (N_16982,N_16010,N_15498);
nor U16983 (N_16983,N_16028,N_15314);
nand U16984 (N_16984,N_15336,N_15232);
and U16985 (N_16985,N_15474,N_15237);
nor U16986 (N_16986,N_15255,N_15567);
xor U16987 (N_16987,N_15888,N_15885);
nand U16988 (N_16988,N_16226,N_15944);
and U16989 (N_16989,N_15898,N_16283);
nand U16990 (N_16990,N_16083,N_16482);
and U16991 (N_16991,N_15781,N_15479);
nand U16992 (N_16992,N_16367,N_16218);
nand U16993 (N_16993,N_16276,N_15907);
nor U16994 (N_16994,N_16057,N_16090);
nor U16995 (N_16995,N_16032,N_15892);
nor U16996 (N_16996,N_15763,N_15851);
or U16997 (N_16997,N_16398,N_15695);
nor U16998 (N_16998,N_16272,N_15324);
and U16999 (N_16999,N_16200,N_16182);
xor U17000 (N_17000,N_15642,N_15032);
nand U17001 (N_17001,N_15319,N_15503);
xor U17002 (N_17002,N_16100,N_15230);
or U17003 (N_17003,N_15855,N_16388);
nor U17004 (N_17004,N_15204,N_15750);
nand U17005 (N_17005,N_15219,N_15850);
and U17006 (N_17006,N_16201,N_15856);
nand U17007 (N_17007,N_15396,N_15511);
nand U17008 (N_17008,N_15951,N_15013);
or U17009 (N_17009,N_15969,N_15301);
and U17010 (N_17010,N_16286,N_15120);
and U17011 (N_17011,N_15473,N_16451);
nor U17012 (N_17012,N_15122,N_16486);
nand U17013 (N_17013,N_16373,N_15906);
nor U17014 (N_17014,N_15547,N_15174);
xor U17015 (N_17015,N_15084,N_15096);
and U17016 (N_17016,N_15038,N_15783);
and U17017 (N_17017,N_15374,N_16113);
nor U17018 (N_17018,N_15192,N_15158);
nand U17019 (N_17019,N_15655,N_16385);
nor U17020 (N_17020,N_15416,N_15175);
and U17021 (N_17021,N_15475,N_15292);
or U17022 (N_17022,N_15931,N_15816);
or U17023 (N_17023,N_15427,N_16064);
xnor U17024 (N_17024,N_16293,N_15751);
or U17025 (N_17025,N_15935,N_15683);
or U17026 (N_17026,N_15619,N_15948);
and U17027 (N_17027,N_15609,N_15994);
and U17028 (N_17028,N_15234,N_15984);
nor U17029 (N_17029,N_15874,N_16277);
nand U17030 (N_17030,N_15787,N_15063);
or U17031 (N_17031,N_15260,N_15397);
nand U17032 (N_17032,N_15822,N_15262);
nor U17033 (N_17033,N_15862,N_16418);
xor U17034 (N_17034,N_15414,N_15403);
nor U17035 (N_17035,N_16119,N_15591);
and U17036 (N_17036,N_15300,N_16413);
nand U17037 (N_17037,N_15870,N_15040);
or U17038 (N_17038,N_15675,N_15765);
xnor U17039 (N_17039,N_15366,N_16107);
nor U17040 (N_17040,N_15653,N_15216);
nand U17041 (N_17041,N_15491,N_15471);
xor U17042 (N_17042,N_15259,N_16236);
or U17043 (N_17043,N_16459,N_15961);
and U17044 (N_17044,N_15919,N_16349);
or U17045 (N_17045,N_16422,N_15917);
or U17046 (N_17046,N_15385,N_16026);
nand U17047 (N_17047,N_15987,N_15321);
nand U17048 (N_17048,N_15748,N_15705);
nand U17049 (N_17049,N_15064,N_15390);
and U17050 (N_17050,N_16328,N_16142);
nand U17051 (N_17051,N_16320,N_15222);
and U17052 (N_17052,N_16303,N_16120);
nor U17053 (N_17053,N_16124,N_16123);
xnor U17054 (N_17054,N_15267,N_16478);
nand U17055 (N_17055,N_15066,N_15409);
nor U17056 (N_17056,N_15461,N_15909);
or U17057 (N_17057,N_15979,N_15821);
or U17058 (N_17058,N_15379,N_15353);
nor U17059 (N_17059,N_15172,N_15679);
and U17060 (N_17060,N_15325,N_15645);
or U17061 (N_17061,N_15808,N_15576);
xnor U17062 (N_17062,N_16213,N_15915);
and U17063 (N_17063,N_15001,N_16299);
xor U17064 (N_17064,N_15636,N_15010);
and U17065 (N_17065,N_15029,N_16229);
nor U17066 (N_17066,N_15717,N_15640);
and U17067 (N_17067,N_15920,N_15253);
xor U17068 (N_17068,N_16225,N_16381);
xor U17069 (N_17069,N_15725,N_15371);
nand U17070 (N_17070,N_15105,N_15877);
nand U17071 (N_17071,N_15210,N_15889);
xor U17072 (N_17072,N_15540,N_16260);
and U17073 (N_17073,N_15927,N_15691);
xor U17074 (N_17074,N_16352,N_15654);
nor U17075 (N_17075,N_15004,N_15943);
or U17076 (N_17076,N_15893,N_15916);
and U17077 (N_17077,N_16384,N_16002);
nor U17078 (N_17078,N_15539,N_15817);
and U17079 (N_17079,N_15753,N_16431);
nor U17080 (N_17080,N_16315,N_16160);
xor U17081 (N_17081,N_15188,N_15810);
or U17082 (N_17082,N_16491,N_16295);
nand U17083 (N_17083,N_15631,N_15686);
and U17084 (N_17084,N_15959,N_16304);
or U17085 (N_17085,N_15315,N_15672);
xor U17086 (N_17086,N_15830,N_15283);
and U17087 (N_17087,N_15166,N_16275);
and U17088 (N_17088,N_16197,N_15745);
nor U17089 (N_17089,N_16076,N_15693);
or U17090 (N_17090,N_15131,N_15598);
and U17091 (N_17091,N_15052,N_15764);
or U17092 (N_17092,N_16063,N_16154);
and U17093 (N_17093,N_16436,N_15431);
xnor U17094 (N_17094,N_15846,N_15991);
nor U17095 (N_17095,N_15226,N_15652);
nand U17096 (N_17096,N_15747,N_16060);
or U17097 (N_17097,N_15463,N_15006);
and U17098 (N_17098,N_16399,N_15998);
and U17099 (N_17099,N_16420,N_15472);
nor U17100 (N_17100,N_15484,N_15894);
nor U17101 (N_17101,N_15235,N_16005);
and U17102 (N_17102,N_16292,N_15720);
nor U17103 (N_17103,N_15095,N_16132);
and U17104 (N_17104,N_15478,N_15716);
and U17105 (N_17105,N_16426,N_15304);
and U17106 (N_17106,N_15828,N_15442);
and U17107 (N_17107,N_16194,N_15247);
and U17108 (N_17108,N_16152,N_15240);
nor U17109 (N_17109,N_16019,N_16231);
nand U17110 (N_17110,N_15288,N_16033);
nor U17111 (N_17111,N_15946,N_15223);
nor U17112 (N_17112,N_15678,N_15164);
xnor U17113 (N_17113,N_15542,N_15908);
xnor U17114 (N_17114,N_15528,N_15138);
nand U17115 (N_17115,N_15342,N_15581);
nor U17116 (N_17116,N_15620,N_15134);
xnor U17117 (N_17117,N_15875,N_15200);
and U17118 (N_17118,N_15180,N_15658);
nor U17119 (N_17119,N_15280,N_15497);
and U17120 (N_17120,N_16450,N_16372);
nor U17121 (N_17121,N_16488,N_15761);
nand U17122 (N_17122,N_15670,N_15269);
nand U17123 (N_17123,N_15561,N_15081);
nand U17124 (N_17124,N_15311,N_15011);
nor U17125 (N_17125,N_16380,N_15712);
nand U17126 (N_17126,N_16361,N_15049);
and U17127 (N_17127,N_15587,N_15841);
xnor U17128 (N_17128,N_16282,N_15085);
or U17129 (N_17129,N_15147,N_15467);
or U17130 (N_17130,N_16443,N_15264);
or U17131 (N_17131,N_16405,N_16209);
nand U17132 (N_17132,N_16301,N_15091);
or U17133 (N_17133,N_15432,N_16403);
xnor U17134 (N_17134,N_15548,N_16092);
and U17135 (N_17135,N_15405,N_15436);
xnor U17136 (N_17136,N_15445,N_15997);
nor U17137 (N_17137,N_15694,N_16284);
xnor U17138 (N_17138,N_15668,N_16185);
or U17139 (N_17139,N_16006,N_15899);
xnor U17140 (N_17140,N_15746,N_16097);
and U17141 (N_17141,N_16397,N_16444);
or U17142 (N_17142,N_15514,N_15231);
or U17143 (N_17143,N_15209,N_16322);
or U17144 (N_17144,N_16454,N_15666);
xor U17145 (N_17145,N_15710,N_15597);
nand U17146 (N_17146,N_15690,N_16370);
xor U17147 (N_17147,N_15560,N_15282);
or U17148 (N_17148,N_16088,N_15217);
or U17149 (N_17149,N_15890,N_16323);
and U17150 (N_17150,N_15923,N_15036);
nor U17151 (N_17151,N_15233,N_15418);
nor U17152 (N_17152,N_16369,N_15339);
nand U17153 (N_17153,N_16419,N_15784);
nor U17154 (N_17154,N_15007,N_15954);
xnor U17155 (N_17155,N_15310,N_15424);
and U17156 (N_17156,N_16112,N_15106);
nand U17157 (N_17157,N_15165,N_15430);
nand U17158 (N_17158,N_15243,N_16377);
and U17159 (N_17159,N_15992,N_15142);
nor U17160 (N_17160,N_15340,N_16011);
xor U17161 (N_17161,N_15302,N_15643);
nor U17162 (N_17162,N_15067,N_15408);
xnor U17163 (N_17163,N_16267,N_16062);
nand U17164 (N_17164,N_16435,N_15357);
nor U17165 (N_17165,N_15555,N_15585);
and U17166 (N_17166,N_16056,N_15020);
nand U17167 (N_17167,N_15330,N_15665);
xnor U17168 (N_17168,N_15433,N_15629);
or U17169 (N_17169,N_15962,N_16116);
nand U17170 (N_17170,N_16153,N_16386);
or U17171 (N_17171,N_15789,N_16251);
nor U17172 (N_17172,N_15439,N_16447);
nor U17173 (N_17173,N_15523,N_15592);
nor U17174 (N_17174,N_15186,N_15778);
nor U17175 (N_17175,N_15033,N_15627);
or U17176 (N_17176,N_15118,N_15628);
and U17177 (N_17177,N_15195,N_15098);
xor U17178 (N_17178,N_15178,N_15938);
or U17179 (N_17179,N_15634,N_15303);
and U17180 (N_17180,N_15605,N_15495);
nor U17181 (N_17181,N_15799,N_15152);
or U17182 (N_17182,N_16089,N_15697);
xnor U17183 (N_17183,N_15285,N_15293);
or U17184 (N_17184,N_16466,N_16481);
nor U17185 (N_17185,N_15077,N_15317);
and U17186 (N_17186,N_16412,N_15873);
nand U17187 (N_17187,N_15593,N_16031);
nand U17188 (N_17188,N_15376,N_15871);
and U17189 (N_17189,N_15270,N_16173);
nor U17190 (N_17190,N_15813,N_16339);
and U17191 (N_17191,N_15980,N_15680);
or U17192 (N_17192,N_15337,N_15356);
or U17193 (N_17193,N_15664,N_15101);
xor U17194 (N_17194,N_15022,N_15351);
nand U17195 (N_17195,N_15265,N_15806);
and U17196 (N_17196,N_15141,N_15731);
nand U17197 (N_17197,N_15803,N_15887);
nand U17198 (N_17198,N_15123,N_15090);
nor U17199 (N_17199,N_15863,N_15744);
and U17200 (N_17200,N_15393,N_15921);
xnor U17201 (N_17201,N_15571,N_15839);
or U17202 (N_17202,N_15976,N_15515);
or U17203 (N_17203,N_15671,N_15297);
or U17204 (N_17204,N_16196,N_16498);
nor U17205 (N_17205,N_15205,N_15083);
nor U17206 (N_17206,N_16199,N_16150);
xor U17207 (N_17207,N_15399,N_15291);
and U17208 (N_17208,N_16012,N_15829);
nor U17209 (N_17209,N_15527,N_15563);
xor U17210 (N_17210,N_15578,N_15749);
nor U17211 (N_17211,N_16145,N_15949);
and U17212 (N_17212,N_16044,N_15942);
and U17213 (N_17213,N_15053,N_15296);
nor U17214 (N_17214,N_16468,N_15380);
and U17215 (N_17215,N_15647,N_15981);
nor U17216 (N_17216,N_16364,N_15532);
and U17217 (N_17217,N_15975,N_15244);
nand U17218 (N_17218,N_15492,N_16198);
xor U17219 (N_17219,N_15177,N_16055);
and U17220 (N_17220,N_16157,N_15382);
and U17221 (N_17221,N_15275,N_16214);
xor U17222 (N_17222,N_16135,N_15626);
or U17223 (N_17223,N_15940,N_15443);
or U17224 (N_17224,N_15019,N_15771);
and U17225 (N_17225,N_15194,N_15607);
or U17226 (N_17226,N_15573,N_15967);
xor U17227 (N_17227,N_15449,N_16393);
or U17228 (N_17228,N_15395,N_15058);
xor U17229 (N_17229,N_16221,N_15148);
xnor U17230 (N_17230,N_16387,N_15891);
nand U17231 (N_17231,N_16464,N_15030);
or U17232 (N_17232,N_15768,N_15126);
xor U17233 (N_17233,N_15221,N_15854);
or U17234 (N_17234,N_15903,N_15362);
xnor U17235 (N_17235,N_15187,N_16022);
nand U17236 (N_17236,N_15639,N_16330);
and U17237 (N_17237,N_15308,N_15733);
nor U17238 (N_17238,N_15354,N_15536);
or U17239 (N_17239,N_16048,N_15481);
or U17240 (N_17240,N_16264,N_15212);
or U17241 (N_17241,N_15825,N_15034);
nand U17242 (N_17242,N_16341,N_15728);
or U17243 (N_17243,N_15911,N_15566);
xor U17244 (N_17244,N_15738,N_15811);
xnor U17245 (N_17245,N_15367,N_16333);
and U17246 (N_17246,N_16271,N_16103);
xnor U17247 (N_17247,N_15791,N_16233);
or U17248 (N_17248,N_15202,N_16143);
xnor U17249 (N_17249,N_16305,N_15128);
or U17250 (N_17250,N_15659,N_15044);
nor U17251 (N_17251,N_16405,N_16278);
or U17252 (N_17252,N_16286,N_16282);
xor U17253 (N_17253,N_15579,N_16389);
xor U17254 (N_17254,N_15610,N_15469);
and U17255 (N_17255,N_15453,N_16193);
and U17256 (N_17256,N_15835,N_15816);
xnor U17257 (N_17257,N_15368,N_16279);
and U17258 (N_17258,N_15155,N_15394);
nor U17259 (N_17259,N_15868,N_16011);
nor U17260 (N_17260,N_15769,N_15231);
nor U17261 (N_17261,N_15849,N_16222);
nor U17262 (N_17262,N_15793,N_16202);
nand U17263 (N_17263,N_16416,N_15068);
and U17264 (N_17264,N_15419,N_16254);
xor U17265 (N_17265,N_15080,N_16124);
nand U17266 (N_17266,N_16026,N_15344);
xor U17267 (N_17267,N_15033,N_16196);
and U17268 (N_17268,N_16122,N_16077);
xnor U17269 (N_17269,N_15838,N_15008);
or U17270 (N_17270,N_15009,N_16078);
and U17271 (N_17271,N_16133,N_16304);
nand U17272 (N_17272,N_15244,N_15291);
nor U17273 (N_17273,N_15578,N_16443);
or U17274 (N_17274,N_15827,N_15424);
and U17275 (N_17275,N_15934,N_16244);
and U17276 (N_17276,N_15190,N_16225);
xor U17277 (N_17277,N_15928,N_15338);
and U17278 (N_17278,N_15037,N_15471);
or U17279 (N_17279,N_15920,N_16245);
nor U17280 (N_17280,N_15247,N_15184);
nor U17281 (N_17281,N_15197,N_15624);
nor U17282 (N_17282,N_16255,N_15230);
nand U17283 (N_17283,N_15727,N_16232);
nor U17284 (N_17284,N_15211,N_16145);
nor U17285 (N_17285,N_15824,N_15108);
xor U17286 (N_17286,N_15100,N_15687);
or U17287 (N_17287,N_16112,N_16073);
and U17288 (N_17288,N_16179,N_16173);
xnor U17289 (N_17289,N_16350,N_15192);
nor U17290 (N_17290,N_16401,N_15957);
and U17291 (N_17291,N_15730,N_16177);
or U17292 (N_17292,N_15442,N_16078);
nor U17293 (N_17293,N_15471,N_15740);
xor U17294 (N_17294,N_15996,N_16247);
or U17295 (N_17295,N_16039,N_15672);
nor U17296 (N_17296,N_16432,N_15804);
and U17297 (N_17297,N_15068,N_15817);
nand U17298 (N_17298,N_16078,N_15548);
xor U17299 (N_17299,N_16116,N_15766);
and U17300 (N_17300,N_16094,N_16400);
nor U17301 (N_17301,N_15455,N_15766);
nor U17302 (N_17302,N_15726,N_15930);
and U17303 (N_17303,N_16374,N_15013);
nand U17304 (N_17304,N_15562,N_16384);
nand U17305 (N_17305,N_15928,N_15146);
nor U17306 (N_17306,N_16038,N_15043);
nand U17307 (N_17307,N_16141,N_16149);
nand U17308 (N_17308,N_15912,N_16453);
nor U17309 (N_17309,N_15713,N_15269);
or U17310 (N_17310,N_15622,N_15443);
or U17311 (N_17311,N_16278,N_15939);
xor U17312 (N_17312,N_15352,N_15516);
nor U17313 (N_17313,N_16408,N_15645);
nor U17314 (N_17314,N_16142,N_15390);
xnor U17315 (N_17315,N_16050,N_15132);
nor U17316 (N_17316,N_15801,N_15118);
and U17317 (N_17317,N_15994,N_15049);
nand U17318 (N_17318,N_15583,N_15547);
nor U17319 (N_17319,N_15940,N_15427);
nand U17320 (N_17320,N_15607,N_15464);
xnor U17321 (N_17321,N_15003,N_15917);
nor U17322 (N_17322,N_16253,N_16201);
or U17323 (N_17323,N_15407,N_15419);
and U17324 (N_17324,N_15787,N_15330);
and U17325 (N_17325,N_15692,N_15431);
or U17326 (N_17326,N_15665,N_16483);
nand U17327 (N_17327,N_15835,N_15820);
nand U17328 (N_17328,N_15742,N_15255);
and U17329 (N_17329,N_16197,N_15778);
nand U17330 (N_17330,N_15999,N_15878);
and U17331 (N_17331,N_15231,N_15448);
nor U17332 (N_17332,N_15066,N_15647);
nand U17333 (N_17333,N_15897,N_16065);
nor U17334 (N_17334,N_15238,N_15844);
nor U17335 (N_17335,N_16410,N_15117);
xor U17336 (N_17336,N_15942,N_15714);
nor U17337 (N_17337,N_15976,N_16116);
or U17338 (N_17338,N_16378,N_15698);
nor U17339 (N_17339,N_16187,N_15246);
and U17340 (N_17340,N_15902,N_15203);
and U17341 (N_17341,N_15150,N_15738);
nand U17342 (N_17342,N_16253,N_15441);
nor U17343 (N_17343,N_15366,N_15018);
and U17344 (N_17344,N_16448,N_15059);
nor U17345 (N_17345,N_15157,N_15982);
and U17346 (N_17346,N_15182,N_15458);
nand U17347 (N_17347,N_15601,N_15986);
or U17348 (N_17348,N_15041,N_16032);
or U17349 (N_17349,N_15180,N_15581);
nand U17350 (N_17350,N_16161,N_15745);
and U17351 (N_17351,N_16098,N_15790);
xnor U17352 (N_17352,N_16401,N_15095);
and U17353 (N_17353,N_15955,N_16445);
nor U17354 (N_17354,N_16437,N_15792);
and U17355 (N_17355,N_15069,N_15163);
nor U17356 (N_17356,N_15692,N_16162);
or U17357 (N_17357,N_15632,N_15158);
nand U17358 (N_17358,N_16002,N_16162);
nor U17359 (N_17359,N_16046,N_15019);
or U17360 (N_17360,N_15329,N_15060);
nand U17361 (N_17361,N_15927,N_15973);
nand U17362 (N_17362,N_16379,N_15541);
and U17363 (N_17363,N_15464,N_15025);
xnor U17364 (N_17364,N_15927,N_16064);
nand U17365 (N_17365,N_16205,N_15255);
nor U17366 (N_17366,N_16499,N_15076);
or U17367 (N_17367,N_15339,N_16478);
nand U17368 (N_17368,N_15797,N_16425);
and U17369 (N_17369,N_15629,N_15717);
nand U17370 (N_17370,N_15632,N_15369);
nand U17371 (N_17371,N_16410,N_15778);
nand U17372 (N_17372,N_16060,N_15729);
and U17373 (N_17373,N_16281,N_15298);
nor U17374 (N_17374,N_15034,N_16264);
xor U17375 (N_17375,N_16334,N_15035);
nand U17376 (N_17376,N_16306,N_16049);
xnor U17377 (N_17377,N_15822,N_15811);
nand U17378 (N_17378,N_16377,N_15657);
nor U17379 (N_17379,N_15956,N_15455);
or U17380 (N_17380,N_16056,N_15323);
xor U17381 (N_17381,N_15921,N_15626);
or U17382 (N_17382,N_15147,N_15879);
xor U17383 (N_17383,N_15341,N_16345);
nand U17384 (N_17384,N_15027,N_15754);
xnor U17385 (N_17385,N_16024,N_15098);
xnor U17386 (N_17386,N_15763,N_15838);
and U17387 (N_17387,N_15869,N_16163);
xor U17388 (N_17388,N_15373,N_15659);
nor U17389 (N_17389,N_16493,N_16111);
xnor U17390 (N_17390,N_15713,N_16337);
nand U17391 (N_17391,N_15312,N_16130);
and U17392 (N_17392,N_15249,N_15299);
and U17393 (N_17393,N_15841,N_16201);
nor U17394 (N_17394,N_15750,N_16449);
or U17395 (N_17395,N_15583,N_15870);
nor U17396 (N_17396,N_16284,N_16228);
nand U17397 (N_17397,N_16391,N_15641);
xor U17398 (N_17398,N_16445,N_16004);
xnor U17399 (N_17399,N_16300,N_15689);
nand U17400 (N_17400,N_16374,N_15692);
xor U17401 (N_17401,N_15162,N_15332);
or U17402 (N_17402,N_16261,N_15489);
and U17403 (N_17403,N_16483,N_15237);
and U17404 (N_17404,N_15213,N_15854);
and U17405 (N_17405,N_15358,N_15647);
and U17406 (N_17406,N_16287,N_15258);
nand U17407 (N_17407,N_16240,N_15644);
and U17408 (N_17408,N_15563,N_16396);
nand U17409 (N_17409,N_15358,N_16314);
or U17410 (N_17410,N_16030,N_15917);
nand U17411 (N_17411,N_16027,N_15485);
and U17412 (N_17412,N_15223,N_15466);
xor U17413 (N_17413,N_15564,N_15642);
or U17414 (N_17414,N_15248,N_15410);
nand U17415 (N_17415,N_16057,N_15132);
and U17416 (N_17416,N_15910,N_16168);
and U17417 (N_17417,N_15887,N_15640);
nor U17418 (N_17418,N_15338,N_15128);
xor U17419 (N_17419,N_16240,N_15382);
and U17420 (N_17420,N_16450,N_15482);
xnor U17421 (N_17421,N_15525,N_15777);
nor U17422 (N_17422,N_15872,N_15055);
nor U17423 (N_17423,N_15033,N_15416);
xor U17424 (N_17424,N_16472,N_15404);
nor U17425 (N_17425,N_16129,N_15793);
xor U17426 (N_17426,N_15061,N_15245);
and U17427 (N_17427,N_16448,N_15478);
nor U17428 (N_17428,N_16157,N_15042);
nor U17429 (N_17429,N_16217,N_15547);
nand U17430 (N_17430,N_15599,N_16084);
or U17431 (N_17431,N_15468,N_15509);
xnor U17432 (N_17432,N_16048,N_15631);
nand U17433 (N_17433,N_15135,N_15395);
and U17434 (N_17434,N_15610,N_15319);
and U17435 (N_17435,N_16387,N_16017);
or U17436 (N_17436,N_15060,N_15683);
nor U17437 (N_17437,N_16073,N_15624);
or U17438 (N_17438,N_15720,N_15108);
nor U17439 (N_17439,N_15156,N_15321);
and U17440 (N_17440,N_16338,N_16041);
and U17441 (N_17441,N_16476,N_16200);
or U17442 (N_17442,N_16398,N_16363);
and U17443 (N_17443,N_15680,N_16351);
nand U17444 (N_17444,N_15318,N_15243);
nor U17445 (N_17445,N_15993,N_15759);
xor U17446 (N_17446,N_16241,N_15120);
xnor U17447 (N_17447,N_15714,N_16174);
or U17448 (N_17448,N_15889,N_16480);
nand U17449 (N_17449,N_16423,N_15660);
nor U17450 (N_17450,N_16294,N_16085);
and U17451 (N_17451,N_16489,N_16409);
or U17452 (N_17452,N_16168,N_15633);
nor U17453 (N_17453,N_15310,N_15236);
nand U17454 (N_17454,N_15115,N_15231);
nor U17455 (N_17455,N_16010,N_15467);
xor U17456 (N_17456,N_16493,N_15814);
xnor U17457 (N_17457,N_15461,N_16400);
nand U17458 (N_17458,N_15727,N_15068);
nand U17459 (N_17459,N_16409,N_16257);
nor U17460 (N_17460,N_15664,N_15475);
nor U17461 (N_17461,N_15927,N_15014);
nor U17462 (N_17462,N_15412,N_16490);
and U17463 (N_17463,N_16026,N_15152);
nor U17464 (N_17464,N_16482,N_15133);
nor U17465 (N_17465,N_16263,N_15397);
nand U17466 (N_17466,N_15459,N_16113);
nor U17467 (N_17467,N_16212,N_16352);
or U17468 (N_17468,N_15408,N_15080);
or U17469 (N_17469,N_16278,N_15400);
nor U17470 (N_17470,N_16351,N_16393);
and U17471 (N_17471,N_16494,N_15120);
or U17472 (N_17472,N_15964,N_15023);
xor U17473 (N_17473,N_16264,N_15367);
nor U17474 (N_17474,N_16323,N_15684);
nor U17475 (N_17475,N_15676,N_15242);
and U17476 (N_17476,N_15527,N_15873);
xor U17477 (N_17477,N_16164,N_16284);
or U17478 (N_17478,N_16192,N_15089);
nand U17479 (N_17479,N_15984,N_16048);
or U17480 (N_17480,N_15085,N_15166);
nand U17481 (N_17481,N_15386,N_15812);
and U17482 (N_17482,N_16346,N_15603);
nor U17483 (N_17483,N_15803,N_16392);
nand U17484 (N_17484,N_15928,N_16444);
nor U17485 (N_17485,N_15125,N_16313);
xor U17486 (N_17486,N_15383,N_16286);
nor U17487 (N_17487,N_15091,N_15323);
and U17488 (N_17488,N_15728,N_15711);
nand U17489 (N_17489,N_16328,N_15416);
nand U17490 (N_17490,N_15683,N_15303);
xor U17491 (N_17491,N_15509,N_15517);
nand U17492 (N_17492,N_15891,N_15037);
or U17493 (N_17493,N_15893,N_16106);
or U17494 (N_17494,N_16093,N_15237);
or U17495 (N_17495,N_15051,N_16106);
or U17496 (N_17496,N_16452,N_15981);
or U17497 (N_17497,N_15795,N_16436);
and U17498 (N_17498,N_15303,N_16131);
or U17499 (N_17499,N_16172,N_16028);
xor U17500 (N_17500,N_16398,N_15592);
or U17501 (N_17501,N_15299,N_16195);
or U17502 (N_17502,N_16251,N_16203);
and U17503 (N_17503,N_15408,N_15295);
and U17504 (N_17504,N_15131,N_15704);
and U17505 (N_17505,N_16065,N_16223);
and U17506 (N_17506,N_15587,N_15376);
nand U17507 (N_17507,N_16367,N_15787);
nand U17508 (N_17508,N_16150,N_15419);
xor U17509 (N_17509,N_15884,N_15184);
xnor U17510 (N_17510,N_16336,N_16350);
xnor U17511 (N_17511,N_15467,N_15246);
or U17512 (N_17512,N_15654,N_15429);
nand U17513 (N_17513,N_16352,N_15040);
or U17514 (N_17514,N_16405,N_16266);
nand U17515 (N_17515,N_15252,N_16435);
nand U17516 (N_17516,N_16271,N_16129);
or U17517 (N_17517,N_16221,N_15083);
nor U17518 (N_17518,N_15150,N_15312);
or U17519 (N_17519,N_16484,N_15023);
xnor U17520 (N_17520,N_16380,N_16251);
xor U17521 (N_17521,N_15654,N_15436);
nand U17522 (N_17522,N_16323,N_15517);
and U17523 (N_17523,N_15603,N_16366);
nand U17524 (N_17524,N_15043,N_15694);
and U17525 (N_17525,N_16380,N_15925);
nand U17526 (N_17526,N_15668,N_16101);
and U17527 (N_17527,N_16231,N_16316);
and U17528 (N_17528,N_15219,N_16394);
or U17529 (N_17529,N_15911,N_16287);
nor U17530 (N_17530,N_16464,N_16003);
xor U17531 (N_17531,N_15548,N_16429);
and U17532 (N_17532,N_15895,N_15715);
and U17533 (N_17533,N_15687,N_15297);
xor U17534 (N_17534,N_15993,N_15042);
nand U17535 (N_17535,N_15009,N_16159);
or U17536 (N_17536,N_15760,N_16346);
nand U17537 (N_17537,N_16410,N_15646);
nor U17538 (N_17538,N_16079,N_16423);
nand U17539 (N_17539,N_15305,N_15486);
xor U17540 (N_17540,N_15787,N_15378);
and U17541 (N_17541,N_15218,N_16262);
and U17542 (N_17542,N_15168,N_15183);
xor U17543 (N_17543,N_16387,N_15256);
nor U17544 (N_17544,N_15894,N_15192);
xnor U17545 (N_17545,N_15216,N_16025);
and U17546 (N_17546,N_16127,N_15275);
nand U17547 (N_17547,N_15516,N_16425);
and U17548 (N_17548,N_16111,N_15178);
or U17549 (N_17549,N_16096,N_15722);
xor U17550 (N_17550,N_15749,N_15893);
or U17551 (N_17551,N_16223,N_16414);
xnor U17552 (N_17552,N_15250,N_15303);
nor U17553 (N_17553,N_15685,N_15739);
xor U17554 (N_17554,N_16020,N_15185);
or U17555 (N_17555,N_15231,N_16327);
xor U17556 (N_17556,N_15291,N_16122);
xor U17557 (N_17557,N_15213,N_16026);
xnor U17558 (N_17558,N_15646,N_15662);
nor U17559 (N_17559,N_16104,N_15524);
nand U17560 (N_17560,N_15578,N_15526);
nand U17561 (N_17561,N_15650,N_15742);
xor U17562 (N_17562,N_16371,N_15237);
xnor U17563 (N_17563,N_16480,N_15095);
or U17564 (N_17564,N_15843,N_15670);
xor U17565 (N_17565,N_15400,N_15387);
nand U17566 (N_17566,N_15260,N_15435);
nor U17567 (N_17567,N_15325,N_16386);
or U17568 (N_17568,N_15546,N_15614);
or U17569 (N_17569,N_15470,N_15074);
nor U17570 (N_17570,N_15585,N_15966);
or U17571 (N_17571,N_15004,N_16265);
nor U17572 (N_17572,N_15542,N_15023);
or U17573 (N_17573,N_15883,N_15370);
or U17574 (N_17574,N_15728,N_16493);
nand U17575 (N_17575,N_15371,N_15272);
and U17576 (N_17576,N_16478,N_16481);
and U17577 (N_17577,N_15999,N_15439);
nand U17578 (N_17578,N_16363,N_15466);
nor U17579 (N_17579,N_15693,N_15349);
nand U17580 (N_17580,N_16225,N_15967);
xnor U17581 (N_17581,N_15915,N_15347);
nor U17582 (N_17582,N_16356,N_15496);
nor U17583 (N_17583,N_16187,N_16206);
xnor U17584 (N_17584,N_16297,N_16084);
nor U17585 (N_17585,N_15270,N_15566);
xor U17586 (N_17586,N_16454,N_15068);
or U17587 (N_17587,N_15703,N_15482);
nor U17588 (N_17588,N_15825,N_15183);
or U17589 (N_17589,N_16066,N_15799);
xnor U17590 (N_17590,N_15698,N_15373);
xor U17591 (N_17591,N_15948,N_15186);
or U17592 (N_17592,N_15394,N_15065);
nand U17593 (N_17593,N_15248,N_15799);
or U17594 (N_17594,N_15385,N_15262);
nor U17595 (N_17595,N_15905,N_16403);
and U17596 (N_17596,N_15020,N_15516);
nand U17597 (N_17597,N_15370,N_16425);
nand U17598 (N_17598,N_15059,N_15641);
and U17599 (N_17599,N_15536,N_15606);
nand U17600 (N_17600,N_15590,N_16225);
or U17601 (N_17601,N_16331,N_16084);
nor U17602 (N_17602,N_15835,N_15597);
xnor U17603 (N_17603,N_15107,N_15880);
xor U17604 (N_17604,N_15352,N_15329);
nor U17605 (N_17605,N_16126,N_15598);
nor U17606 (N_17606,N_15058,N_15112);
xnor U17607 (N_17607,N_15449,N_15222);
nor U17608 (N_17608,N_16121,N_15664);
and U17609 (N_17609,N_15455,N_15077);
nor U17610 (N_17610,N_16183,N_15411);
nor U17611 (N_17611,N_15628,N_16245);
xor U17612 (N_17612,N_15724,N_15972);
xor U17613 (N_17613,N_15288,N_16111);
or U17614 (N_17614,N_15581,N_16477);
or U17615 (N_17615,N_16499,N_15837);
nor U17616 (N_17616,N_16227,N_15994);
and U17617 (N_17617,N_16484,N_16146);
or U17618 (N_17618,N_15827,N_16446);
nor U17619 (N_17619,N_15821,N_15721);
nand U17620 (N_17620,N_16335,N_16214);
nor U17621 (N_17621,N_15148,N_16404);
nor U17622 (N_17622,N_15101,N_15441);
nand U17623 (N_17623,N_16107,N_15603);
nand U17624 (N_17624,N_15692,N_15890);
nor U17625 (N_17625,N_16162,N_16402);
xor U17626 (N_17626,N_15717,N_15100);
xor U17627 (N_17627,N_15209,N_15014);
nor U17628 (N_17628,N_16438,N_15028);
xor U17629 (N_17629,N_16155,N_15199);
nor U17630 (N_17630,N_16120,N_15324);
nand U17631 (N_17631,N_16115,N_15050);
nor U17632 (N_17632,N_16195,N_16238);
nor U17633 (N_17633,N_15876,N_15433);
nor U17634 (N_17634,N_15450,N_15558);
and U17635 (N_17635,N_15984,N_15260);
xnor U17636 (N_17636,N_15171,N_16248);
and U17637 (N_17637,N_15317,N_15102);
and U17638 (N_17638,N_15406,N_16109);
or U17639 (N_17639,N_15465,N_15728);
and U17640 (N_17640,N_15993,N_16438);
nor U17641 (N_17641,N_15970,N_16224);
nor U17642 (N_17642,N_16219,N_15422);
nor U17643 (N_17643,N_15565,N_16453);
xor U17644 (N_17644,N_15483,N_16385);
xnor U17645 (N_17645,N_15802,N_15115);
or U17646 (N_17646,N_15970,N_16178);
and U17647 (N_17647,N_15565,N_15606);
nand U17648 (N_17648,N_16001,N_15535);
xnor U17649 (N_17649,N_15471,N_15884);
nor U17650 (N_17650,N_15507,N_16396);
and U17651 (N_17651,N_15997,N_15130);
nand U17652 (N_17652,N_15742,N_15814);
and U17653 (N_17653,N_15296,N_16175);
nor U17654 (N_17654,N_16195,N_15954);
nand U17655 (N_17655,N_15218,N_16231);
nand U17656 (N_17656,N_15472,N_15053);
xor U17657 (N_17657,N_15431,N_15996);
xor U17658 (N_17658,N_15618,N_16492);
nand U17659 (N_17659,N_16420,N_16337);
nor U17660 (N_17660,N_15631,N_15851);
or U17661 (N_17661,N_15859,N_15577);
nand U17662 (N_17662,N_15548,N_16077);
nand U17663 (N_17663,N_15661,N_15093);
or U17664 (N_17664,N_15026,N_15760);
nand U17665 (N_17665,N_15771,N_16277);
xor U17666 (N_17666,N_15935,N_15058);
nor U17667 (N_17667,N_15306,N_16313);
nand U17668 (N_17668,N_15183,N_16423);
or U17669 (N_17669,N_15911,N_15691);
nand U17670 (N_17670,N_16435,N_15251);
or U17671 (N_17671,N_16267,N_15555);
nand U17672 (N_17672,N_15650,N_16398);
or U17673 (N_17673,N_15667,N_15741);
or U17674 (N_17674,N_15358,N_15451);
and U17675 (N_17675,N_15758,N_15594);
nand U17676 (N_17676,N_16309,N_15991);
xor U17677 (N_17677,N_16238,N_15786);
nor U17678 (N_17678,N_15833,N_16416);
nor U17679 (N_17679,N_15043,N_15311);
nor U17680 (N_17680,N_15802,N_16166);
and U17681 (N_17681,N_16449,N_15165);
or U17682 (N_17682,N_15777,N_15814);
nand U17683 (N_17683,N_15765,N_15531);
nand U17684 (N_17684,N_15388,N_15731);
or U17685 (N_17685,N_15932,N_15072);
nor U17686 (N_17686,N_15834,N_15084);
nor U17687 (N_17687,N_15142,N_15990);
nor U17688 (N_17688,N_16308,N_15247);
and U17689 (N_17689,N_15571,N_16096);
or U17690 (N_17690,N_15977,N_16306);
xor U17691 (N_17691,N_15444,N_16126);
or U17692 (N_17692,N_15779,N_15818);
or U17693 (N_17693,N_15705,N_15262);
nor U17694 (N_17694,N_15460,N_16296);
nor U17695 (N_17695,N_15892,N_16003);
or U17696 (N_17696,N_15430,N_16002);
nor U17697 (N_17697,N_15320,N_15528);
nor U17698 (N_17698,N_16487,N_15803);
xor U17699 (N_17699,N_15962,N_15560);
nand U17700 (N_17700,N_16285,N_15979);
and U17701 (N_17701,N_16402,N_15947);
xor U17702 (N_17702,N_15604,N_15431);
nand U17703 (N_17703,N_16015,N_15805);
nor U17704 (N_17704,N_15442,N_15531);
nor U17705 (N_17705,N_15111,N_16129);
nor U17706 (N_17706,N_15011,N_15892);
or U17707 (N_17707,N_15882,N_16274);
nor U17708 (N_17708,N_16355,N_15295);
and U17709 (N_17709,N_15747,N_16152);
xor U17710 (N_17710,N_15293,N_15502);
xnor U17711 (N_17711,N_15589,N_15619);
nand U17712 (N_17712,N_15200,N_15411);
nand U17713 (N_17713,N_16171,N_15652);
xor U17714 (N_17714,N_15946,N_15017);
and U17715 (N_17715,N_16437,N_15610);
or U17716 (N_17716,N_15801,N_15170);
xnor U17717 (N_17717,N_15439,N_15688);
nand U17718 (N_17718,N_15990,N_16457);
or U17719 (N_17719,N_16078,N_15447);
nor U17720 (N_17720,N_16451,N_15699);
and U17721 (N_17721,N_15189,N_15369);
and U17722 (N_17722,N_15148,N_15724);
nand U17723 (N_17723,N_15643,N_15110);
nand U17724 (N_17724,N_15725,N_15058);
xnor U17725 (N_17725,N_15706,N_15087);
nor U17726 (N_17726,N_16410,N_16156);
and U17727 (N_17727,N_16005,N_15659);
xnor U17728 (N_17728,N_15546,N_16478);
or U17729 (N_17729,N_15073,N_15877);
or U17730 (N_17730,N_15212,N_15374);
or U17731 (N_17731,N_16453,N_15094);
xnor U17732 (N_17732,N_16280,N_15137);
xnor U17733 (N_17733,N_15947,N_16285);
or U17734 (N_17734,N_15464,N_16272);
xnor U17735 (N_17735,N_15088,N_16205);
nor U17736 (N_17736,N_16219,N_15070);
or U17737 (N_17737,N_16006,N_15403);
xor U17738 (N_17738,N_15344,N_15876);
nor U17739 (N_17739,N_15262,N_15788);
nor U17740 (N_17740,N_15514,N_16111);
or U17741 (N_17741,N_15684,N_15509);
nand U17742 (N_17742,N_15261,N_15666);
xor U17743 (N_17743,N_15339,N_15904);
nor U17744 (N_17744,N_15654,N_15671);
or U17745 (N_17745,N_16290,N_16422);
or U17746 (N_17746,N_16485,N_15061);
and U17747 (N_17747,N_16283,N_16188);
and U17748 (N_17748,N_15692,N_15079);
nor U17749 (N_17749,N_15575,N_15713);
xor U17750 (N_17750,N_16089,N_16334);
xnor U17751 (N_17751,N_15237,N_16051);
nor U17752 (N_17752,N_15740,N_15234);
xor U17753 (N_17753,N_16276,N_15452);
and U17754 (N_17754,N_16357,N_16468);
or U17755 (N_17755,N_16491,N_15421);
and U17756 (N_17756,N_15655,N_15011);
or U17757 (N_17757,N_15730,N_15514);
nor U17758 (N_17758,N_15291,N_16099);
nand U17759 (N_17759,N_16299,N_15814);
and U17760 (N_17760,N_15768,N_15022);
or U17761 (N_17761,N_15038,N_16264);
nand U17762 (N_17762,N_15487,N_15006);
nor U17763 (N_17763,N_15526,N_15349);
xnor U17764 (N_17764,N_15473,N_16301);
and U17765 (N_17765,N_15280,N_15094);
xnor U17766 (N_17766,N_16294,N_15164);
or U17767 (N_17767,N_15483,N_15993);
or U17768 (N_17768,N_15067,N_15972);
nor U17769 (N_17769,N_15386,N_15787);
nand U17770 (N_17770,N_15477,N_15702);
or U17771 (N_17771,N_15050,N_16188);
or U17772 (N_17772,N_16012,N_15056);
and U17773 (N_17773,N_16493,N_15806);
nand U17774 (N_17774,N_16338,N_16357);
and U17775 (N_17775,N_16495,N_15158);
nor U17776 (N_17776,N_15968,N_16103);
nand U17777 (N_17777,N_15097,N_15966);
nand U17778 (N_17778,N_16184,N_15416);
nor U17779 (N_17779,N_16093,N_15857);
xnor U17780 (N_17780,N_15515,N_15654);
xor U17781 (N_17781,N_15318,N_15936);
nand U17782 (N_17782,N_15400,N_15270);
nor U17783 (N_17783,N_15704,N_16389);
nor U17784 (N_17784,N_15887,N_15299);
xnor U17785 (N_17785,N_15608,N_15310);
and U17786 (N_17786,N_15069,N_15125);
xor U17787 (N_17787,N_15422,N_15808);
and U17788 (N_17788,N_16039,N_15914);
or U17789 (N_17789,N_15251,N_15146);
and U17790 (N_17790,N_16019,N_16406);
nand U17791 (N_17791,N_15186,N_16188);
or U17792 (N_17792,N_15131,N_15094);
xnor U17793 (N_17793,N_15129,N_15849);
nand U17794 (N_17794,N_16244,N_15108);
nand U17795 (N_17795,N_15843,N_15546);
xor U17796 (N_17796,N_15477,N_15717);
nand U17797 (N_17797,N_15707,N_16051);
nand U17798 (N_17798,N_15460,N_15945);
and U17799 (N_17799,N_15166,N_15145);
or U17800 (N_17800,N_15614,N_15981);
nor U17801 (N_17801,N_16369,N_16022);
and U17802 (N_17802,N_15265,N_15863);
nand U17803 (N_17803,N_15375,N_16047);
and U17804 (N_17804,N_15697,N_15601);
and U17805 (N_17805,N_15730,N_16277);
nor U17806 (N_17806,N_15223,N_15117);
nor U17807 (N_17807,N_15549,N_15621);
xor U17808 (N_17808,N_15564,N_15832);
nand U17809 (N_17809,N_15455,N_16102);
xnor U17810 (N_17810,N_16172,N_15260);
xor U17811 (N_17811,N_16371,N_16077);
and U17812 (N_17812,N_16282,N_15536);
nor U17813 (N_17813,N_15373,N_16365);
xor U17814 (N_17814,N_15298,N_15639);
nor U17815 (N_17815,N_16261,N_15609);
xor U17816 (N_17816,N_15472,N_15096);
and U17817 (N_17817,N_16359,N_15035);
nor U17818 (N_17818,N_15533,N_15136);
nor U17819 (N_17819,N_16293,N_16109);
nand U17820 (N_17820,N_15670,N_15794);
or U17821 (N_17821,N_15268,N_15801);
nor U17822 (N_17822,N_16293,N_16233);
nor U17823 (N_17823,N_15923,N_15251);
and U17824 (N_17824,N_15445,N_16209);
or U17825 (N_17825,N_15353,N_15555);
nor U17826 (N_17826,N_16003,N_15120);
nand U17827 (N_17827,N_15756,N_16117);
nor U17828 (N_17828,N_15472,N_16492);
and U17829 (N_17829,N_16083,N_15301);
xor U17830 (N_17830,N_15175,N_15124);
xnor U17831 (N_17831,N_15025,N_15207);
or U17832 (N_17832,N_15084,N_16285);
nor U17833 (N_17833,N_16017,N_15528);
and U17834 (N_17834,N_15505,N_15052);
nand U17835 (N_17835,N_15987,N_15113);
or U17836 (N_17836,N_15965,N_15610);
and U17837 (N_17837,N_15739,N_15920);
nand U17838 (N_17838,N_15014,N_15136);
xnor U17839 (N_17839,N_16367,N_15979);
nor U17840 (N_17840,N_15751,N_16134);
xor U17841 (N_17841,N_15131,N_15610);
nand U17842 (N_17842,N_15391,N_15046);
nand U17843 (N_17843,N_15861,N_16230);
and U17844 (N_17844,N_15409,N_15147);
and U17845 (N_17845,N_15741,N_15778);
and U17846 (N_17846,N_15810,N_16265);
or U17847 (N_17847,N_16263,N_15652);
nand U17848 (N_17848,N_16486,N_16198);
xnor U17849 (N_17849,N_16268,N_16118);
or U17850 (N_17850,N_15015,N_15885);
nor U17851 (N_17851,N_15480,N_15836);
nand U17852 (N_17852,N_16441,N_16035);
or U17853 (N_17853,N_15584,N_15554);
nor U17854 (N_17854,N_16427,N_15958);
xor U17855 (N_17855,N_16476,N_15037);
nand U17856 (N_17856,N_16263,N_16428);
and U17857 (N_17857,N_16056,N_15178);
xor U17858 (N_17858,N_15105,N_15819);
nor U17859 (N_17859,N_15519,N_15241);
nand U17860 (N_17860,N_15708,N_16147);
nor U17861 (N_17861,N_15614,N_15989);
and U17862 (N_17862,N_15593,N_16216);
nand U17863 (N_17863,N_15206,N_16262);
xnor U17864 (N_17864,N_15735,N_15436);
nand U17865 (N_17865,N_16173,N_15107);
nand U17866 (N_17866,N_16319,N_15075);
nand U17867 (N_17867,N_16006,N_16452);
nor U17868 (N_17868,N_15912,N_15795);
or U17869 (N_17869,N_15541,N_15051);
xnor U17870 (N_17870,N_16028,N_16275);
or U17871 (N_17871,N_15868,N_15245);
xor U17872 (N_17872,N_15355,N_15944);
nor U17873 (N_17873,N_15350,N_15948);
xnor U17874 (N_17874,N_16369,N_16432);
or U17875 (N_17875,N_16301,N_16137);
and U17876 (N_17876,N_15891,N_15491);
nor U17877 (N_17877,N_15494,N_16016);
nor U17878 (N_17878,N_16139,N_16252);
or U17879 (N_17879,N_15761,N_15464);
and U17880 (N_17880,N_16020,N_15326);
and U17881 (N_17881,N_16164,N_16288);
xor U17882 (N_17882,N_15972,N_15717);
nor U17883 (N_17883,N_15724,N_15293);
nor U17884 (N_17884,N_15766,N_15877);
or U17885 (N_17885,N_16404,N_15114);
and U17886 (N_17886,N_16336,N_16141);
xnor U17887 (N_17887,N_15783,N_15678);
nand U17888 (N_17888,N_15690,N_15659);
nor U17889 (N_17889,N_15987,N_16335);
and U17890 (N_17890,N_15011,N_15441);
and U17891 (N_17891,N_15905,N_16000);
xnor U17892 (N_17892,N_15735,N_15967);
nor U17893 (N_17893,N_16137,N_16034);
nand U17894 (N_17894,N_16323,N_15635);
and U17895 (N_17895,N_15773,N_15975);
or U17896 (N_17896,N_15881,N_15132);
or U17897 (N_17897,N_16071,N_15929);
nand U17898 (N_17898,N_15453,N_16261);
or U17899 (N_17899,N_15892,N_16448);
and U17900 (N_17900,N_15370,N_16362);
nor U17901 (N_17901,N_16482,N_15561);
xnor U17902 (N_17902,N_15760,N_15964);
or U17903 (N_17903,N_15429,N_15307);
and U17904 (N_17904,N_15897,N_15836);
nand U17905 (N_17905,N_15411,N_16064);
xnor U17906 (N_17906,N_16005,N_16315);
or U17907 (N_17907,N_16097,N_15639);
nand U17908 (N_17908,N_16313,N_15948);
nor U17909 (N_17909,N_15523,N_15836);
or U17910 (N_17910,N_15660,N_15625);
nand U17911 (N_17911,N_15655,N_15039);
nand U17912 (N_17912,N_15373,N_16488);
nor U17913 (N_17913,N_16056,N_15205);
nor U17914 (N_17914,N_15278,N_15359);
xnor U17915 (N_17915,N_15973,N_15219);
nand U17916 (N_17916,N_16360,N_16252);
xor U17917 (N_17917,N_16394,N_16129);
nor U17918 (N_17918,N_15782,N_15106);
nor U17919 (N_17919,N_15722,N_15981);
nor U17920 (N_17920,N_15462,N_15658);
nor U17921 (N_17921,N_15204,N_15962);
nor U17922 (N_17922,N_15689,N_15916);
and U17923 (N_17923,N_15891,N_16154);
and U17924 (N_17924,N_15844,N_15562);
nor U17925 (N_17925,N_15869,N_16073);
xnor U17926 (N_17926,N_15984,N_15570);
and U17927 (N_17927,N_15888,N_15823);
and U17928 (N_17928,N_16065,N_15478);
nor U17929 (N_17929,N_15500,N_15093);
nand U17930 (N_17930,N_15477,N_16006);
nor U17931 (N_17931,N_15064,N_15428);
and U17932 (N_17932,N_16148,N_15101);
or U17933 (N_17933,N_15700,N_15744);
nor U17934 (N_17934,N_15508,N_15629);
xor U17935 (N_17935,N_15291,N_15709);
and U17936 (N_17936,N_16383,N_16021);
or U17937 (N_17937,N_15314,N_15278);
nand U17938 (N_17938,N_15968,N_16359);
and U17939 (N_17939,N_15392,N_15648);
nor U17940 (N_17940,N_16453,N_16146);
nand U17941 (N_17941,N_15190,N_16452);
or U17942 (N_17942,N_15986,N_15831);
nand U17943 (N_17943,N_16237,N_15884);
nor U17944 (N_17944,N_15729,N_15755);
or U17945 (N_17945,N_16261,N_15560);
nor U17946 (N_17946,N_16276,N_16043);
nand U17947 (N_17947,N_15888,N_16297);
or U17948 (N_17948,N_15935,N_16215);
and U17949 (N_17949,N_16265,N_15858);
nand U17950 (N_17950,N_15372,N_15643);
and U17951 (N_17951,N_15893,N_16365);
nand U17952 (N_17952,N_15359,N_15451);
nand U17953 (N_17953,N_16335,N_16252);
and U17954 (N_17954,N_15210,N_15525);
nor U17955 (N_17955,N_15916,N_16186);
nor U17956 (N_17956,N_15967,N_16024);
or U17957 (N_17957,N_15771,N_15331);
and U17958 (N_17958,N_16078,N_15728);
or U17959 (N_17959,N_16244,N_16170);
nand U17960 (N_17960,N_15248,N_15549);
nand U17961 (N_17961,N_15907,N_15196);
nand U17962 (N_17962,N_15212,N_16054);
nor U17963 (N_17963,N_16103,N_16295);
nand U17964 (N_17964,N_15220,N_15395);
nand U17965 (N_17965,N_16180,N_15117);
nand U17966 (N_17966,N_16292,N_15862);
or U17967 (N_17967,N_16078,N_16167);
nor U17968 (N_17968,N_15203,N_15413);
xnor U17969 (N_17969,N_15531,N_15861);
xnor U17970 (N_17970,N_15136,N_15782);
and U17971 (N_17971,N_15008,N_16088);
xnor U17972 (N_17972,N_15426,N_15663);
or U17973 (N_17973,N_16356,N_15391);
nor U17974 (N_17974,N_16256,N_15456);
or U17975 (N_17975,N_15661,N_15903);
or U17976 (N_17976,N_15198,N_15044);
or U17977 (N_17977,N_16058,N_15709);
nand U17978 (N_17978,N_15850,N_15309);
xor U17979 (N_17979,N_15329,N_15791);
nand U17980 (N_17980,N_16294,N_15064);
nor U17981 (N_17981,N_16006,N_15629);
nor U17982 (N_17982,N_15267,N_16308);
or U17983 (N_17983,N_15116,N_15602);
or U17984 (N_17984,N_16108,N_15279);
or U17985 (N_17985,N_15090,N_15691);
xor U17986 (N_17986,N_15696,N_15548);
or U17987 (N_17987,N_16432,N_16426);
and U17988 (N_17988,N_15361,N_15223);
or U17989 (N_17989,N_16466,N_16496);
and U17990 (N_17990,N_15782,N_16218);
nand U17991 (N_17991,N_15325,N_16103);
nor U17992 (N_17992,N_16293,N_15539);
and U17993 (N_17993,N_16308,N_16005);
nand U17994 (N_17994,N_15398,N_15721);
or U17995 (N_17995,N_16188,N_15170);
nor U17996 (N_17996,N_15972,N_16176);
and U17997 (N_17997,N_15054,N_16280);
and U17998 (N_17998,N_15461,N_15264);
and U17999 (N_17999,N_16273,N_15867);
nor U18000 (N_18000,N_17451,N_17954);
and U18001 (N_18001,N_16640,N_17643);
and U18002 (N_18002,N_17253,N_17407);
nand U18003 (N_18003,N_17932,N_17634);
nor U18004 (N_18004,N_17546,N_17023);
or U18005 (N_18005,N_17547,N_17068);
nand U18006 (N_18006,N_17359,N_16712);
xor U18007 (N_18007,N_17102,N_17840);
or U18008 (N_18008,N_17138,N_17197);
and U18009 (N_18009,N_16677,N_16780);
or U18010 (N_18010,N_17944,N_16846);
nor U18011 (N_18011,N_16593,N_17737);
nor U18012 (N_18012,N_17849,N_16675);
or U18013 (N_18013,N_16632,N_17041);
and U18014 (N_18014,N_16832,N_16786);
and U18015 (N_18015,N_17838,N_16917);
nand U18016 (N_18016,N_16743,N_17566);
nor U18017 (N_18017,N_16788,N_17416);
nand U18018 (N_18018,N_17446,N_17015);
xnor U18019 (N_18019,N_16643,N_17523);
or U18020 (N_18020,N_17894,N_16967);
nand U18021 (N_18021,N_16560,N_16611);
and U18022 (N_18022,N_17286,N_17484);
or U18023 (N_18023,N_17163,N_17714);
or U18024 (N_18024,N_17482,N_17221);
and U18025 (N_18025,N_17135,N_17788);
or U18026 (N_18026,N_17623,N_17209);
and U18027 (N_18027,N_16623,N_17987);
nor U18028 (N_18028,N_16886,N_16584);
nor U18029 (N_18029,N_16888,N_16730);
nor U18030 (N_18030,N_17669,N_16918);
nand U18031 (N_18031,N_17156,N_17252);
and U18032 (N_18032,N_16987,N_16607);
xnor U18033 (N_18033,N_17474,N_17294);
and U18034 (N_18034,N_17240,N_17909);
nor U18035 (N_18035,N_16581,N_17401);
nor U18036 (N_18036,N_17131,N_17734);
and U18037 (N_18037,N_17116,N_17191);
xor U18038 (N_18038,N_17193,N_17939);
nand U18039 (N_18039,N_17267,N_17848);
and U18040 (N_18040,N_16760,N_16538);
and U18041 (N_18041,N_17605,N_17236);
or U18042 (N_18042,N_17897,N_17347);
and U18043 (N_18043,N_17481,N_17445);
nor U18044 (N_18044,N_16842,N_17383);
xnor U18045 (N_18045,N_16983,N_17828);
nand U18046 (N_18046,N_17364,N_17542);
xor U18047 (N_18047,N_17980,N_16506);
xor U18048 (N_18048,N_17952,N_16847);
nor U18049 (N_18049,N_17914,N_16951);
xnor U18050 (N_18050,N_17146,N_17958);
or U18051 (N_18051,N_17915,N_17504);
xor U18052 (N_18052,N_16613,N_17260);
and U18053 (N_18053,N_16570,N_17560);
and U18054 (N_18054,N_17567,N_17083);
xor U18055 (N_18055,N_16541,N_16817);
nand U18056 (N_18056,N_16668,N_17646);
nor U18057 (N_18057,N_17405,N_16891);
nor U18058 (N_18058,N_17493,N_17895);
nand U18059 (N_18059,N_17893,N_16910);
and U18060 (N_18060,N_17033,N_17762);
xor U18061 (N_18061,N_16756,N_16678);
and U18062 (N_18062,N_17403,N_17164);
xnor U18063 (N_18063,N_17730,N_16901);
and U18064 (N_18064,N_17208,N_16770);
nor U18065 (N_18065,N_16664,N_17469);
nor U18066 (N_18066,N_17871,N_17192);
and U18067 (N_18067,N_16665,N_17820);
nor U18068 (N_18068,N_16954,N_17650);
xor U18069 (N_18069,N_16695,N_16543);
nor U18070 (N_18070,N_17532,N_17630);
or U18071 (N_18071,N_16572,N_16993);
and U18072 (N_18072,N_16911,N_16592);
nand U18073 (N_18073,N_16723,N_16673);
nand U18074 (N_18074,N_17076,N_17534);
and U18075 (N_18075,N_16682,N_17761);
and U18076 (N_18076,N_16648,N_17779);
and U18077 (N_18077,N_17308,N_17908);
and U18078 (N_18078,N_17512,N_17262);
and U18079 (N_18079,N_17603,N_16858);
and U18080 (N_18080,N_17463,N_17419);
and U18081 (N_18081,N_16588,N_17886);
nor U18082 (N_18082,N_17077,N_17212);
xor U18083 (N_18083,N_17148,N_17637);
xnor U18084 (N_18084,N_17806,N_17591);
or U18085 (N_18085,N_17925,N_17723);
and U18086 (N_18086,N_16729,N_17214);
nand U18087 (N_18087,N_17654,N_17042);
nor U18088 (N_18088,N_16562,N_17215);
nor U18089 (N_18089,N_17781,N_17257);
nand U18090 (N_18090,N_16551,N_16809);
xnor U18091 (N_18091,N_17398,N_17689);
and U18092 (N_18092,N_17856,N_17425);
nor U18093 (N_18093,N_17506,N_17049);
nor U18094 (N_18094,N_16616,N_17985);
nand U18095 (N_18095,N_17736,N_17622);
or U18096 (N_18096,N_17843,N_17518);
nor U18097 (N_18097,N_17079,N_17786);
and U18098 (N_18098,N_16844,N_17947);
nor U18099 (N_18099,N_16948,N_17489);
xor U18100 (N_18100,N_17485,N_16594);
nand U18101 (N_18101,N_17675,N_16652);
nand U18102 (N_18102,N_16973,N_16773);
and U18103 (N_18103,N_17767,N_17242);
or U18104 (N_18104,N_17016,N_17683);
nand U18105 (N_18105,N_17115,N_17804);
nor U18106 (N_18106,N_16827,N_16900);
nor U18107 (N_18107,N_17237,N_17072);
and U18108 (N_18108,N_17390,N_17353);
nor U18109 (N_18109,N_17306,N_17065);
nor U18110 (N_18110,N_17576,N_17352);
and U18111 (N_18111,N_16864,N_17964);
nand U18112 (N_18112,N_17845,N_16564);
xor U18113 (N_18113,N_16565,N_17552);
nand U18114 (N_18114,N_16889,N_17662);
nor U18115 (N_18115,N_17497,N_16772);
and U18116 (N_18116,N_16676,N_16526);
or U18117 (N_18117,N_17619,N_17855);
nand U18118 (N_18118,N_16843,N_17300);
and U18119 (N_18119,N_17176,N_17219);
nand U18120 (N_18120,N_17344,N_17968);
nand U18121 (N_18121,N_17113,N_17125);
nor U18122 (N_18122,N_16749,N_16792);
xnor U18123 (N_18123,N_17002,N_17269);
nand U18124 (N_18124,N_17872,N_16708);
or U18125 (N_18125,N_16956,N_17022);
or U18126 (N_18126,N_17074,N_17367);
xor U18127 (N_18127,N_17942,N_17490);
and U18128 (N_18128,N_16826,N_16599);
and U18129 (N_18129,N_16688,N_16833);
nand U18130 (N_18130,N_16503,N_17165);
and U18131 (N_18131,N_17168,N_17741);
nand U18132 (N_18132,N_16720,N_16801);
or U18133 (N_18133,N_17608,N_17513);
and U18134 (N_18134,N_17284,N_17177);
nor U18135 (N_18135,N_17655,N_16566);
xnor U18136 (N_18136,N_17205,N_16701);
nand U18137 (N_18137,N_16898,N_16812);
xnor U18138 (N_18138,N_16573,N_17647);
nor U18139 (N_18139,N_16602,N_16816);
xor U18140 (N_18140,N_16968,N_17038);
xor U18141 (N_18141,N_17004,N_17449);
xor U18142 (N_18142,N_16975,N_17140);
nor U18143 (N_18143,N_17509,N_16995);
and U18144 (N_18144,N_17568,N_17812);
or U18145 (N_18145,N_17333,N_16965);
nand U18146 (N_18146,N_16627,N_16776);
nand U18147 (N_18147,N_17617,N_16742);
and U18148 (N_18148,N_16717,N_17027);
nand U18149 (N_18149,N_17050,N_17951);
nand U18150 (N_18150,N_17424,N_17198);
nand U18151 (N_18151,N_17412,N_17147);
nand U18152 (N_18152,N_17747,N_17919);
xnor U18153 (N_18153,N_17765,N_17001);
and U18154 (N_18154,N_16798,N_16774);
and U18155 (N_18155,N_16721,N_17020);
and U18156 (N_18156,N_17644,N_17230);
or U18157 (N_18157,N_17107,N_16750);
and U18158 (N_18158,N_17305,N_16582);
xnor U18159 (N_18159,N_16763,N_16872);
xor U18160 (N_18160,N_16785,N_17764);
and U18161 (N_18161,N_17733,N_16986);
xnor U18162 (N_18162,N_17317,N_17393);
and U18163 (N_18163,N_16765,N_17217);
nand U18164 (N_18164,N_17834,N_17226);
or U18165 (N_18165,N_17320,N_17210);
or U18166 (N_18166,N_17061,N_16806);
nand U18167 (N_18167,N_16852,N_16795);
xnor U18168 (N_18168,N_17385,N_17447);
nor U18169 (N_18169,N_17372,N_17880);
and U18170 (N_18170,N_17956,N_17883);
nand U18171 (N_18171,N_16681,N_17461);
nor U18172 (N_18172,N_16571,N_16981);
or U18173 (N_18173,N_17373,N_17090);
nand U18174 (N_18174,N_16764,N_17105);
xnor U18175 (N_18175,N_17720,N_17615);
nand U18176 (N_18176,N_17151,N_17776);
and U18177 (N_18177,N_17108,N_17099);
or U18178 (N_18178,N_17078,N_17955);
xor U18179 (N_18179,N_17480,N_17274);
xor U18180 (N_18180,N_17235,N_17564);
xnor U18181 (N_18181,N_17745,N_17249);
xnor U18182 (N_18182,N_17624,N_17738);
xnor U18183 (N_18183,N_16713,N_17940);
nand U18184 (N_18184,N_17064,N_17415);
and U18185 (N_18185,N_17303,N_17429);
and U18186 (N_18186,N_17960,N_17441);
or U18187 (N_18187,N_17790,N_17611);
and U18188 (N_18188,N_17013,N_17690);
nor U18189 (N_18189,N_17340,N_17578);
or U18190 (N_18190,N_16778,N_16950);
or U18191 (N_18191,N_17247,N_16614);
xnor U18192 (N_18192,N_16610,N_16869);
xor U18193 (N_18193,N_17255,N_16529);
or U18194 (N_18194,N_17450,N_16545);
nor U18195 (N_18195,N_17595,N_16793);
nand U18196 (N_18196,N_16969,N_17335);
nand U18197 (N_18197,N_16881,N_17783);
and U18198 (N_18198,N_17103,N_16892);
nand U18199 (N_18199,N_16794,N_16929);
xnor U18200 (N_18200,N_17561,N_17739);
and U18201 (N_18201,N_16521,N_16567);
xor U18202 (N_18202,N_17931,N_17460);
and U18203 (N_18203,N_16909,N_17477);
or U18204 (N_18204,N_17473,N_17711);
or U18205 (N_18205,N_17659,N_16662);
and U18206 (N_18206,N_17256,N_16552);
nand U18207 (N_18207,N_17316,N_17997);
and U18208 (N_18208,N_17133,N_17059);
and U18209 (N_18209,N_17837,N_17978);
nand U18210 (N_18210,N_17825,N_16800);
xnor U18211 (N_18211,N_17979,N_17858);
nor U18212 (N_18212,N_17826,N_17218);
nand U18213 (N_18213,N_17819,N_17973);
xnor U18214 (N_18214,N_16690,N_16639);
nor U18215 (N_18215,N_17996,N_17898);
nand U18216 (N_18216,N_17321,N_16893);
or U18217 (N_18217,N_17012,N_17427);
and U18218 (N_18218,N_17860,N_16600);
nand U18219 (N_18219,N_17376,N_17992);
and U18220 (N_18220,N_16976,N_17189);
nand U18221 (N_18221,N_17588,N_17999);
xnor U18222 (N_18222,N_17586,N_17453);
nor U18223 (N_18223,N_17440,N_17727);
nor U18224 (N_18224,N_16885,N_17904);
and U18225 (N_18225,N_16530,N_16904);
xor U18226 (N_18226,N_17713,N_17876);
or U18227 (N_18227,N_16789,N_16884);
and U18228 (N_18228,N_17551,N_17058);
xor U18229 (N_18229,N_17370,N_17297);
or U18230 (N_18230,N_17454,N_17599);
nand U18231 (N_18231,N_16738,N_17428);
nor U18232 (N_18232,N_16849,N_17098);
nand U18233 (N_18233,N_17649,N_17044);
nand U18234 (N_18234,N_17232,N_17961);
and U18235 (N_18235,N_17500,N_17043);
nand U18236 (N_18236,N_16554,N_17106);
nand U18237 (N_18237,N_17196,N_16906);
or U18238 (N_18238,N_17291,N_17807);
nor U18239 (N_18239,N_16934,N_16609);
or U18240 (N_18240,N_17859,N_17363);
nor U18241 (N_18241,N_17081,N_17332);
and U18242 (N_18242,N_16779,N_16622);
nand U18243 (N_18243,N_17533,N_16861);
and U18244 (N_18244,N_16595,N_17417);
nand U18245 (N_18245,N_17963,N_17742);
and U18246 (N_18246,N_16865,N_16907);
and U18247 (N_18247,N_17793,N_17063);
or U18248 (N_18248,N_16533,N_17271);
nand U18249 (N_18249,N_17657,N_16509);
nor U18250 (N_18250,N_17562,N_17696);
or U18251 (N_18251,N_17970,N_17094);
and U18252 (N_18252,N_17642,N_16796);
or U18253 (N_18253,N_17379,N_17035);
xnor U18254 (N_18254,N_16957,N_17318);
or U18255 (N_18255,N_17361,N_17557);
and U18256 (N_18256,N_16870,N_17527);
nor U18257 (N_18257,N_17167,N_17170);
and U18258 (N_18258,N_16755,N_16875);
nor U18259 (N_18259,N_16985,N_17206);
xnor U18260 (N_18260,N_17005,N_17648);
and U18261 (N_18261,N_17935,N_17254);
and U18262 (N_18262,N_17540,N_17854);
nand U18263 (N_18263,N_16860,N_16590);
and U18264 (N_18264,N_16645,N_16558);
nand U18265 (N_18265,N_17682,N_16555);
nor U18266 (N_18266,N_17055,N_17857);
and U18267 (N_18267,N_17844,N_17991);
nand U18268 (N_18268,N_16697,N_17368);
nor U18269 (N_18269,N_17937,N_17651);
or U18270 (N_18270,N_17350,N_17088);
and U18271 (N_18271,N_17414,N_16807);
nand U18272 (N_18272,N_17345,N_17132);
xor U18273 (N_18273,N_16597,N_16687);
xor U18274 (N_18274,N_16994,N_17162);
nor U18275 (N_18275,N_16962,N_17635);
and U18276 (N_18276,N_17275,N_17025);
nand U18277 (N_18277,N_17057,N_17281);
or U18278 (N_18278,N_17459,N_16728);
xor U18279 (N_18279,N_17029,N_17965);
xor U18280 (N_18280,N_17906,N_16947);
nand U18281 (N_18281,N_16857,N_17080);
xnor U18282 (N_18282,N_17128,N_16699);
xor U18283 (N_18283,N_17516,N_17550);
and U18284 (N_18284,N_17520,N_17680);
nand U18285 (N_18285,N_16641,N_17531);
or U18286 (N_18286,N_17452,N_17929);
nor U18287 (N_18287,N_17465,N_17716);
xnor U18288 (N_18288,N_16838,N_17143);
and U18289 (N_18289,N_17822,N_17541);
nand U18290 (N_18290,N_16820,N_17549);
nor U18291 (N_18291,N_17095,N_17123);
xnor U18292 (N_18292,N_17943,N_16739);
or U18293 (N_18293,N_17186,N_17348);
and U18294 (N_18294,N_16502,N_17671);
nor U18295 (N_18295,N_16504,N_17325);
xnor U18296 (N_18296,N_16859,N_16867);
xnor U18297 (N_18297,N_16671,N_17674);
nor U18298 (N_18298,N_16630,N_17902);
xor U18299 (N_18299,N_17225,N_17111);
and U18300 (N_18300,N_17778,N_17019);
nand U18301 (N_18301,N_17693,N_16598);
and U18302 (N_18302,N_16810,N_16575);
and U18303 (N_18303,N_17977,N_16549);
nand U18304 (N_18304,N_16821,N_17548);
nand U18305 (N_18305,N_17927,N_17290);
nand U18306 (N_18306,N_17075,N_16928);
xor U18307 (N_18307,N_16922,N_17334);
nor U18308 (N_18308,N_17101,N_17270);
nor U18309 (N_18309,N_16633,N_17701);
or U18310 (N_18310,N_16762,N_17584);
nand U18311 (N_18311,N_17688,N_16932);
or U18312 (N_18312,N_17375,N_17323);
xnor U18313 (N_18313,N_16718,N_17666);
and U18314 (N_18314,N_17056,N_17472);
xnor U18315 (N_18315,N_17673,N_16658);
xnor U18316 (N_18316,N_17545,N_17342);
or U18317 (N_18317,N_17604,N_17182);
nor U18318 (N_18318,N_16577,N_17507);
and U18319 (N_18319,N_17406,N_16596);
nor U18320 (N_18320,N_17633,N_16784);
xnor U18321 (N_18321,N_17863,N_17136);
and U18322 (N_18322,N_16899,N_17795);
nor U18323 (N_18323,N_17621,N_16915);
or U18324 (N_18324,N_17338,N_16510);
xor U18325 (N_18325,N_17556,N_16710);
or U18326 (N_18326,N_17686,N_16505);
or U18327 (N_18327,N_16589,N_17559);
nand U18328 (N_18328,N_16725,N_17918);
or U18329 (N_18329,N_17744,N_16876);
nor U18330 (N_18330,N_17468,N_17870);
and U18331 (N_18331,N_16923,N_17581);
nand U18332 (N_18332,N_16656,N_17749);
and U18333 (N_18333,N_16719,N_17729);
nor U18334 (N_18334,N_17708,N_17360);
xor U18335 (N_18335,N_17010,N_17458);
and U18336 (N_18336,N_16831,N_17264);
or U18337 (N_18337,N_17171,N_16926);
nor U18338 (N_18338,N_17528,N_17582);
nand U18339 (N_18339,N_17705,N_17014);
and U18340 (N_18340,N_17246,N_17339);
nand U18341 (N_18341,N_16659,N_16525);
xor U18342 (N_18342,N_16706,N_16635);
and U18343 (N_18343,N_17413,N_17530);
nor U18344 (N_18344,N_16603,N_16925);
nor U18345 (N_18345,N_17658,N_16912);
nand U18346 (N_18346,N_16657,N_17821);
xnor U18347 (N_18347,N_17295,N_17455);
nand U18348 (N_18348,N_17718,N_16568);
nand U18349 (N_18349,N_17910,N_17157);
and U18350 (N_18350,N_17382,N_17715);
nand U18351 (N_18351,N_17652,N_17994);
nor U18352 (N_18352,N_17879,N_17137);
or U18353 (N_18353,N_17250,N_17535);
xnor U18354 (N_18354,N_17972,N_17593);
nor U18355 (N_18355,N_17684,N_16920);
and U18356 (N_18356,N_17231,N_16548);
or U18357 (N_18357,N_17831,N_17847);
or U18358 (N_18358,N_16921,N_17104);
nor U18359 (N_18359,N_17957,N_17846);
nand U18360 (N_18360,N_17791,N_17031);
nor U18361 (N_18361,N_17354,N_17488);
nor U18362 (N_18362,N_17261,N_17492);
nor U18363 (N_18363,N_17073,N_17725);
nand U18364 (N_18364,N_16650,N_17687);
xnor U18365 (N_18365,N_17503,N_17558);
or U18366 (N_18366,N_17572,N_16601);
nand U18367 (N_18367,N_17202,N_17802);
xnor U18368 (N_18368,N_17830,N_17620);
xor U18369 (N_18369,N_16866,N_17313);
or U18370 (N_18370,N_17122,N_16724);
nor U18371 (N_18371,N_16705,N_16804);
nor U18372 (N_18372,N_16823,N_16963);
nand U18373 (N_18373,N_17054,N_16946);
nor U18374 (N_18374,N_17378,N_16685);
xor U18375 (N_18375,N_16716,N_16797);
or U18376 (N_18376,N_17695,N_17989);
or U18377 (N_18377,N_16781,N_17755);
nor U18378 (N_18378,N_16539,N_17810);
nand U18379 (N_18379,N_17850,N_17501);
nor U18380 (N_18380,N_17636,N_17975);
xor U18381 (N_18381,N_17607,N_17888);
nand U18382 (N_18382,N_17431,N_16734);
nand U18383 (N_18383,N_17948,N_17200);
and U18384 (N_18384,N_16841,N_16692);
nor U18385 (N_18385,N_16970,N_16583);
or U18386 (N_18386,N_17923,N_17362);
nand U18387 (N_18387,N_16837,N_16580);
and U18388 (N_18388,N_16534,N_16767);
xor U18389 (N_18389,N_16751,N_17722);
nand U18390 (N_18390,N_17134,N_17172);
nor U18391 (N_18391,N_16972,N_16523);
nand U18392 (N_18392,N_17051,N_17011);
nor U18393 (N_18393,N_16752,N_17962);
nor U18394 (N_18394,N_17905,N_16544);
and U18395 (N_18395,N_17203,N_17084);
xor U18396 (N_18396,N_17238,N_17495);
nor U18397 (N_18397,N_17769,N_16989);
xnor U18398 (N_18398,N_17502,N_17155);
and U18399 (N_18399,N_17190,N_16937);
and U18400 (N_18400,N_16887,N_17173);
nand U18401 (N_18401,N_17438,N_17435);
nand U18402 (N_18402,N_17048,N_17357);
xnor U18403 (N_18403,N_17663,N_16653);
nor U18404 (N_18404,N_17785,N_17187);
or U18405 (N_18405,N_17456,N_17945);
nor U18406 (N_18406,N_16514,N_17265);
xor U18407 (N_18407,N_16945,N_17109);
nand U18408 (N_18408,N_17224,N_17579);
or U18409 (N_18409,N_17832,N_17371);
nor U18410 (N_18410,N_17752,N_16722);
nand U18411 (N_18411,N_17126,N_16615);
nand U18412 (N_18412,N_16988,N_16711);
xor U18413 (N_18413,N_17117,N_17211);
or U18414 (N_18414,N_16908,N_17865);
nor U18415 (N_18415,N_17796,N_17841);
nor U18416 (N_18416,N_17381,N_16996);
nor U18417 (N_18417,N_17327,N_16941);
or U18418 (N_18418,N_17891,N_16698);
xnor U18419 (N_18419,N_17921,N_17312);
nand U18420 (N_18420,N_17784,N_16740);
and U18421 (N_18421,N_16579,N_16830);
or U18422 (N_18422,N_16894,N_17066);
and U18423 (N_18423,N_17139,N_17096);
nor U18424 (N_18424,N_16938,N_16748);
or U18425 (N_18425,N_17032,N_17422);
nand U18426 (N_18426,N_17158,N_17008);
or U18427 (N_18427,N_17719,N_16927);
and U18428 (N_18428,N_17439,N_17301);
xnor U18429 (N_18429,N_17600,N_16576);
nor U18430 (N_18430,N_17580,N_16815);
and U18431 (N_18431,N_17037,N_17349);
xor U18432 (N_18432,N_17307,N_16873);
xnor U18433 (N_18433,N_17288,N_17803);
nor U18434 (N_18434,N_17366,N_17751);
or U18435 (N_18435,N_17887,N_17178);
xor U18436 (N_18436,N_16782,N_17437);
nor U18437 (N_18437,N_17543,N_17248);
nand U18438 (N_18438,N_17750,N_17780);
nand U18439 (N_18439,N_16990,N_17154);
nor U18440 (N_18440,N_17901,N_17587);
nor U18441 (N_18441,N_17602,N_17569);
or U18442 (N_18442,N_17628,N_17656);
nand U18443 (N_18443,N_16625,N_16546);
nand U18444 (N_18444,N_17694,N_17092);
nand U18445 (N_18445,N_17526,N_16661);
xor U18446 (N_18446,N_16914,N_17724);
and U18447 (N_18447,N_17400,N_17610);
nor U18448 (N_18448,N_17896,N_17967);
nor U18449 (N_18449,N_16537,N_17241);
nand U18450 (N_18450,N_17946,N_17071);
and U18451 (N_18451,N_17279,N_17553);
xnor U18452 (N_18452,N_17585,N_17388);
nor U18453 (N_18453,N_17315,N_16977);
nand U18454 (N_18454,N_17930,N_17142);
or U18455 (N_18455,N_17377,N_17285);
and U18456 (N_18456,N_17629,N_16618);
and U18457 (N_18457,N_17772,N_17959);
and U18458 (N_18458,N_16850,N_17920);
nand U18459 (N_18459,N_17185,N_17598);
xnor U18460 (N_18460,N_16768,N_17861);
xor U18461 (N_18461,N_17982,N_17748);
xor U18462 (N_18462,N_17983,N_17322);
or U18463 (N_18463,N_17047,N_16997);
nand U18464 (N_18464,N_16811,N_17478);
xor U18465 (N_18465,N_16933,N_17021);
nor U18466 (N_18466,N_16984,N_17799);
or U18467 (N_18467,N_17276,N_17774);
nand U18468 (N_18468,N_17805,N_17852);
or U18469 (N_18469,N_16703,N_17691);
xor U18470 (N_18470,N_17233,N_17302);
or U18471 (N_18471,N_17777,N_16879);
nor U18472 (N_18472,N_16636,N_16839);
nand U18473 (N_18473,N_17386,N_17789);
and U18474 (N_18474,N_17036,N_17756);
and U18475 (N_18475,N_16655,N_17510);
xor U18476 (N_18476,N_17258,N_17326);
xor U18477 (N_18477,N_17152,N_17287);
xor U18478 (N_18478,N_17199,N_17692);
and U18479 (N_18479,N_17356,N_17119);
xnor U18480 (N_18480,N_17184,N_17129);
or U18481 (N_18481,N_17678,N_17766);
nor U18482 (N_18482,N_17763,N_17869);
nor U18483 (N_18483,N_17702,N_17836);
or U18484 (N_18484,N_17709,N_17299);
xnor U18485 (N_18485,N_17928,N_17792);
nor U18486 (N_18486,N_17809,N_16855);
nand U18487 (N_18487,N_17645,N_16761);
xnor U18488 (N_18488,N_16591,N_16949);
and U18489 (N_18489,N_16644,N_17800);
nand U18490 (N_18490,N_16709,N_16727);
or U18491 (N_18491,N_16629,N_17827);
and U18492 (N_18492,N_17003,N_16634);
or U18493 (N_18493,N_16535,N_17726);
xnor U18494 (N_18494,N_17007,N_17627);
nor U18495 (N_18495,N_16757,N_17950);
nor U18496 (N_18496,N_16999,N_17505);
and U18497 (N_18497,N_17746,N_17862);
nand U18498 (N_18498,N_16802,N_17570);
or U18499 (N_18499,N_17913,N_16853);
nor U18500 (N_18500,N_17907,N_17679);
nor U18501 (N_18501,N_16836,N_16845);
or U18502 (N_18502,N_17521,N_16683);
or U18503 (N_18503,N_17638,N_17434);
and U18504 (N_18504,N_17220,N_16878);
nand U18505 (N_18505,N_17430,N_17544);
or U18506 (N_18506,N_16825,N_17758);
nand U18507 (N_18507,N_16744,N_16696);
and U18508 (N_18508,N_17341,N_17293);
or U18509 (N_18509,N_16998,N_16512);
nor U18510 (N_18510,N_17421,N_16787);
or U18511 (N_18511,N_17974,N_17053);
and U18512 (N_18512,N_17272,N_16874);
and U18513 (N_18513,N_17743,N_16672);
nand U18514 (N_18514,N_17900,N_16732);
and U18515 (N_18515,N_16515,N_17426);
nor U18516 (N_18516,N_17522,N_16619);
nand U18517 (N_18517,N_17864,N_16979);
nor U18518 (N_18518,N_17467,N_17583);
xnor U18519 (N_18519,N_17922,N_17175);
nor U18520 (N_18520,N_16822,N_17319);
nand U18521 (N_18521,N_16769,N_16513);
nor U18522 (N_18522,N_17384,N_17677);
or U18523 (N_18523,N_17229,N_16517);
xor U18524 (N_18524,N_17995,N_17195);
or U18525 (N_18525,N_17494,N_17571);
nor U18526 (N_18526,N_17612,N_16704);
nor U18527 (N_18527,N_17017,N_16771);
nor U18528 (N_18528,N_17402,N_16882);
xor U18529 (N_18529,N_17818,N_17771);
nor U18530 (N_18530,N_17292,N_16578);
xor U18531 (N_18531,N_17912,N_16902);
nand U18532 (N_18532,N_16519,N_16516);
nor U18533 (N_18533,N_17601,N_17984);
nand U18534 (N_18534,N_16741,N_16903);
nand U18535 (N_18535,N_17498,N_17130);
xor U18536 (N_18536,N_17089,N_17775);
or U18537 (N_18537,N_17590,N_17087);
nand U18538 (N_18538,N_17577,N_16654);
and U18539 (N_18539,N_17277,N_16674);
xnor U18540 (N_18540,N_17525,N_17877);
nor U18541 (N_18541,N_16960,N_16758);
or U18542 (N_18542,N_17903,N_17731);
nand U18543 (N_18543,N_16895,N_17597);
nand U18544 (N_18544,N_17380,N_17770);
nor U18545 (N_18545,N_17814,N_16574);
nor U18546 (N_18546,N_17085,N_17483);
and U18547 (N_18547,N_16966,N_17517);
xor U18548 (N_18548,N_17149,N_16670);
and U18549 (N_18549,N_17120,N_16803);
and U18550 (N_18550,N_16943,N_16527);
xnor U18551 (N_18551,N_17660,N_16936);
nand U18552 (N_18552,N_17853,N_17976);
nor U18553 (N_18553,N_16992,N_17815);
and U18554 (N_18554,N_17668,N_16829);
nand U18555 (N_18555,N_17890,N_16814);
nor U18556 (N_18556,N_17153,N_16766);
nor U18557 (N_18557,N_16563,N_17222);
nand U18558 (N_18558,N_17759,N_17993);
xor U18559 (N_18559,N_17062,N_17470);
or U18560 (N_18560,N_17309,N_17916);
and U18561 (N_18561,N_17889,N_16606);
and U18562 (N_18562,N_17911,N_16731);
nand U18563 (N_18563,N_16585,N_17273);
and U18564 (N_18564,N_16935,N_16542);
or U18565 (N_18565,N_16799,N_16835);
nor U18566 (N_18566,N_16532,N_16508);
nand U18567 (N_18567,N_17251,N_16862);
xor U18568 (N_18568,N_17851,N_17626);
or U18569 (N_18569,N_17884,N_16746);
nor U18570 (N_18570,N_16714,N_17487);
nor U18571 (N_18571,N_17444,N_17538);
xor U18572 (N_18572,N_17926,N_16883);
nand U18573 (N_18573,N_17337,N_17304);
or U18574 (N_18574,N_17329,N_17392);
nand U18575 (N_18575,N_16547,N_17728);
nor U18576 (N_18576,N_17787,N_17245);
and U18577 (N_18577,N_17740,N_17632);
nor U18578 (N_18578,N_17676,N_16931);
or U18579 (N_18579,N_17592,N_17801);
xor U18580 (N_18580,N_17127,N_17179);
or U18581 (N_18581,N_16818,N_17259);
or U18582 (N_18582,N_17418,N_17408);
nand U18583 (N_18583,N_17554,N_17039);
or U18584 (N_18584,N_17710,N_17613);
nand U18585 (N_18585,N_16553,N_17892);
xnor U18586 (N_18586,N_17699,N_16689);
and U18587 (N_18587,N_17515,N_16702);
nor U18588 (N_18588,N_17466,N_17310);
xor U18589 (N_18589,N_17462,N_17816);
xnor U18590 (N_18590,N_16608,N_17511);
nand U18591 (N_18591,N_17698,N_17881);
and U18592 (N_18592,N_16686,N_16851);
nand U18593 (N_18593,N_17409,N_16569);
and U18594 (N_18594,N_17009,N_16586);
nor U18595 (N_18595,N_16775,N_16754);
xor U18596 (N_18596,N_17296,N_16637);
or U18597 (N_18597,N_17213,N_17589);
nor U18598 (N_18598,N_17144,N_17735);
and U18599 (N_18599,N_16626,N_17389);
xor U18600 (N_18600,N_16663,N_17732);
xnor U18601 (N_18601,N_16991,N_17018);
and U18602 (N_18602,N_17717,N_16561);
or U18603 (N_18603,N_16790,N_17443);
nor U18604 (N_18604,N_16550,N_17491);
nor U18605 (N_18605,N_16735,N_17124);
and U18606 (N_18606,N_16647,N_17933);
or U18607 (N_18607,N_17024,N_16856);
xor U18608 (N_18608,N_16557,N_17082);
or U18609 (N_18609,N_16939,N_17873);
nor U18610 (N_18610,N_17665,N_16924);
or U18611 (N_18611,N_17829,N_17263);
xor U18612 (N_18612,N_16819,N_17343);
nand U18613 (N_18613,N_17365,N_17969);
xor U18614 (N_18614,N_16733,N_17040);
xor U18615 (N_18615,N_17432,N_17216);
and U18616 (N_18616,N_17704,N_17324);
nor U18617 (N_18617,N_17808,N_17596);
and U18618 (N_18618,N_17953,N_17000);
nor U18619 (N_18619,N_17391,N_17006);
nand U18620 (N_18620,N_16694,N_17374);
and U18621 (N_18621,N_17070,N_16500);
nor U18622 (N_18622,N_16805,N_17998);
nand U18623 (N_18623,N_17697,N_16964);
nor U18624 (N_18624,N_17574,N_17314);
or U18625 (N_18625,N_16854,N_16540);
xor U18626 (N_18626,N_17411,N_17625);
nand U18627 (N_18627,N_16646,N_17201);
xor U18628 (N_18628,N_16890,N_17183);
nor U18629 (N_18629,N_16507,N_16834);
nand U18630 (N_18630,N_16961,N_17824);
and U18631 (N_18631,N_16679,N_17399);
and U18632 (N_18632,N_17150,N_17986);
xnor U18633 (N_18633,N_16959,N_17112);
or U18634 (N_18634,N_17536,N_17594);
xor U18635 (N_18635,N_16955,N_16896);
and U18636 (N_18636,N_16522,N_17966);
or U18637 (N_18637,N_16624,N_17046);
or U18638 (N_18638,N_16919,N_16971);
and U18639 (N_18639,N_16974,N_16736);
and U18640 (N_18640,N_17283,N_16813);
and U18641 (N_18641,N_16691,N_16669);
xnor U18642 (N_18642,N_16982,N_17575);
nor U18643 (N_18643,N_17614,N_17653);
nand U18644 (N_18644,N_16684,N_16617);
and U18645 (N_18645,N_16913,N_17086);
or U18646 (N_18646,N_17941,N_17529);
xnor U18647 (N_18647,N_17028,N_17754);
nand U18648 (N_18648,N_17110,N_16715);
and U18649 (N_18649,N_17797,N_17410);
or U18650 (N_18650,N_17813,N_16520);
nor U18651 (N_18651,N_16700,N_17331);
nand U18652 (N_18652,N_17244,N_16824);
or U18653 (N_18653,N_17145,N_17387);
nand U18654 (N_18654,N_17936,N_17631);
nand U18655 (N_18655,N_17433,N_17067);
nand U18656 (N_18656,N_17166,N_17336);
or U18657 (N_18657,N_17311,N_17060);
nor U18658 (N_18658,N_17706,N_17981);
and U18659 (N_18659,N_16877,N_17681);
or U18660 (N_18660,N_17882,N_17874);
or U18661 (N_18661,N_16944,N_17700);
and U18662 (N_18662,N_16518,N_16880);
xor U18663 (N_18663,N_17369,N_17757);
and U18664 (N_18664,N_17639,N_17464);
and U18665 (N_18665,N_17833,N_17811);
nor U18666 (N_18666,N_16759,N_17330);
nand U18667 (N_18667,N_17223,N_17358);
xnor U18668 (N_18668,N_16649,N_17169);
nand U18669 (N_18669,N_16726,N_16863);
xnor U18670 (N_18670,N_17519,N_17794);
and U18671 (N_18671,N_17100,N_17773);
xnor U18672 (N_18672,N_17181,N_16660);
nand U18673 (N_18673,N_17239,N_17159);
or U18674 (N_18674,N_17685,N_17423);
nor U18675 (N_18675,N_17924,N_17457);
nand U18676 (N_18676,N_17712,N_16612);
or U18677 (N_18677,N_17207,N_16605);
xor U18678 (N_18678,N_17034,N_17475);
xor U18679 (N_18679,N_17282,N_16621);
nand U18680 (N_18680,N_17875,N_17355);
xnor U18681 (N_18681,N_17760,N_17990);
xnor U18682 (N_18682,N_17664,N_16905);
nand U18683 (N_18683,N_16559,N_17878);
nand U18684 (N_18684,N_16958,N_17661);
nand U18685 (N_18685,N_17141,N_16871);
and U18686 (N_18686,N_17641,N_17514);
and U18687 (N_18687,N_17486,N_17835);
nand U18688 (N_18688,N_17508,N_17988);
and U18689 (N_18689,N_17606,N_17565);
nor U18690 (N_18690,N_16667,N_16680);
xor U18691 (N_18691,N_16942,N_17188);
or U18692 (N_18692,N_17667,N_16638);
nand U18693 (N_18693,N_17204,N_16828);
and U18694 (N_18694,N_16940,N_17121);
or U18695 (N_18695,N_17045,N_17234);
and U18696 (N_18696,N_17026,N_17328);
and U18697 (N_18697,N_17069,N_17823);
or U18698 (N_18698,N_16737,N_17616);
and U18699 (N_18699,N_16666,N_16531);
and U18700 (N_18700,N_16953,N_17524);
and U18701 (N_18701,N_17114,N_16840);
xnor U18702 (N_18702,N_17174,N_17537);
and U18703 (N_18703,N_16777,N_16707);
nor U18704 (N_18704,N_16808,N_16511);
and U18705 (N_18705,N_16791,N_17097);
xnor U18706 (N_18706,N_16642,N_17496);
and U18707 (N_18707,N_17753,N_16753);
or U18708 (N_18708,N_17420,N_17938);
and U18709 (N_18709,N_17476,N_16745);
and U18710 (N_18710,N_17160,N_17396);
and U18711 (N_18711,N_17842,N_17640);
nor U18712 (N_18712,N_17346,N_17093);
or U18713 (N_18713,N_17091,N_17471);
xnor U18714 (N_18714,N_17670,N_17030);
nand U18715 (N_18715,N_16628,N_16651);
nor U18716 (N_18716,N_16980,N_17298);
xnor U18717 (N_18717,N_17394,N_17351);
nor U18718 (N_18718,N_17867,N_17268);
nor U18719 (N_18719,N_17609,N_17278);
or U18720 (N_18720,N_16747,N_17949);
nand U18721 (N_18721,N_17555,N_16978);
xor U18722 (N_18722,N_16524,N_16631);
and U18723 (N_18723,N_17442,N_16620);
or U18724 (N_18724,N_16868,N_17227);
and U18725 (N_18725,N_17289,N_17672);
nor U18726 (N_18726,N_16848,N_17798);
nor U18727 (N_18727,N_17885,N_17397);
and U18728 (N_18728,N_17180,N_16930);
and U18729 (N_18729,N_17703,N_17817);
xnor U18730 (N_18730,N_17499,N_17479);
nor U18731 (N_18731,N_17573,N_17539);
xnor U18732 (N_18732,N_17194,N_16501);
nor U18733 (N_18733,N_17266,N_17618);
or U18734 (N_18734,N_17707,N_16604);
nor U18735 (N_18735,N_16587,N_17782);
and U18736 (N_18736,N_16556,N_16693);
or U18737 (N_18737,N_17768,N_17395);
xor U18738 (N_18738,N_16952,N_17721);
and U18739 (N_18739,N_16536,N_17563);
nand U18740 (N_18740,N_17161,N_17866);
and U18741 (N_18741,N_17052,N_17971);
or U18742 (N_18742,N_17436,N_17934);
xnor U18743 (N_18743,N_17868,N_17917);
nor U18744 (N_18744,N_17228,N_17404);
xor U18745 (N_18745,N_17118,N_17243);
and U18746 (N_18746,N_17448,N_17899);
nor U18747 (N_18747,N_17280,N_16916);
and U18748 (N_18748,N_16528,N_16783);
nand U18749 (N_18749,N_17839,N_16897);
and U18750 (N_18750,N_16832,N_17056);
or U18751 (N_18751,N_17566,N_17971);
and U18752 (N_18752,N_17923,N_17382);
and U18753 (N_18753,N_16570,N_17670);
or U18754 (N_18754,N_16573,N_17434);
nor U18755 (N_18755,N_17053,N_17739);
nand U18756 (N_18756,N_16568,N_16660);
or U18757 (N_18757,N_17269,N_17422);
or U18758 (N_18758,N_16865,N_16628);
or U18759 (N_18759,N_16680,N_17813);
nor U18760 (N_18760,N_17325,N_16555);
nand U18761 (N_18761,N_17785,N_17954);
nand U18762 (N_18762,N_16939,N_17702);
nor U18763 (N_18763,N_17897,N_17050);
xnor U18764 (N_18764,N_17461,N_17882);
xor U18765 (N_18765,N_17022,N_17887);
nand U18766 (N_18766,N_16671,N_17523);
xor U18767 (N_18767,N_16778,N_17950);
and U18768 (N_18768,N_16711,N_17907);
nor U18769 (N_18769,N_16895,N_16751);
nor U18770 (N_18770,N_17757,N_17993);
xor U18771 (N_18771,N_17802,N_16747);
nor U18772 (N_18772,N_16978,N_16807);
nor U18773 (N_18773,N_16781,N_17869);
nand U18774 (N_18774,N_17386,N_17187);
or U18775 (N_18775,N_16869,N_16760);
xor U18776 (N_18776,N_17551,N_16664);
xnor U18777 (N_18777,N_17735,N_17927);
and U18778 (N_18778,N_17094,N_16575);
xnor U18779 (N_18779,N_16987,N_16525);
and U18780 (N_18780,N_17538,N_17542);
or U18781 (N_18781,N_17913,N_17129);
and U18782 (N_18782,N_16569,N_17241);
and U18783 (N_18783,N_17039,N_17530);
xor U18784 (N_18784,N_17518,N_17945);
or U18785 (N_18785,N_16569,N_17140);
and U18786 (N_18786,N_17187,N_17305);
xor U18787 (N_18787,N_16998,N_17535);
nor U18788 (N_18788,N_16812,N_17867);
nand U18789 (N_18789,N_16971,N_16998);
xor U18790 (N_18790,N_16598,N_17223);
xnor U18791 (N_18791,N_17561,N_17801);
nor U18792 (N_18792,N_17258,N_16538);
xor U18793 (N_18793,N_16779,N_17563);
and U18794 (N_18794,N_16875,N_17542);
xnor U18795 (N_18795,N_16513,N_17646);
xnor U18796 (N_18796,N_17118,N_16996);
nand U18797 (N_18797,N_16689,N_17053);
and U18798 (N_18798,N_16790,N_17590);
or U18799 (N_18799,N_17381,N_17551);
nor U18800 (N_18800,N_17614,N_16787);
nor U18801 (N_18801,N_17392,N_17114);
and U18802 (N_18802,N_17130,N_17014);
nor U18803 (N_18803,N_16724,N_17324);
and U18804 (N_18804,N_16666,N_16590);
nand U18805 (N_18805,N_17737,N_17249);
xnor U18806 (N_18806,N_16706,N_17102);
xnor U18807 (N_18807,N_17843,N_17274);
or U18808 (N_18808,N_16587,N_16542);
nor U18809 (N_18809,N_17347,N_17295);
xor U18810 (N_18810,N_16643,N_16552);
xnor U18811 (N_18811,N_17363,N_16893);
nor U18812 (N_18812,N_16948,N_17423);
or U18813 (N_18813,N_17549,N_17188);
and U18814 (N_18814,N_16911,N_17624);
or U18815 (N_18815,N_17370,N_17203);
and U18816 (N_18816,N_17628,N_16569);
nor U18817 (N_18817,N_17135,N_17050);
nand U18818 (N_18818,N_16627,N_16558);
or U18819 (N_18819,N_17592,N_17342);
nor U18820 (N_18820,N_17939,N_17186);
and U18821 (N_18821,N_16772,N_17083);
and U18822 (N_18822,N_17056,N_17617);
nand U18823 (N_18823,N_16767,N_16698);
nor U18824 (N_18824,N_16785,N_17039);
xnor U18825 (N_18825,N_17982,N_16848);
nand U18826 (N_18826,N_17524,N_17958);
and U18827 (N_18827,N_17698,N_16761);
or U18828 (N_18828,N_17862,N_17413);
xnor U18829 (N_18829,N_16596,N_17716);
and U18830 (N_18830,N_17837,N_17114);
xnor U18831 (N_18831,N_17598,N_17594);
xnor U18832 (N_18832,N_17841,N_16541);
nor U18833 (N_18833,N_17831,N_16783);
xor U18834 (N_18834,N_17730,N_16701);
or U18835 (N_18835,N_17387,N_16554);
nand U18836 (N_18836,N_17006,N_16603);
nand U18837 (N_18837,N_17353,N_17742);
nand U18838 (N_18838,N_16765,N_17865);
nor U18839 (N_18839,N_16749,N_16645);
nand U18840 (N_18840,N_17715,N_17733);
and U18841 (N_18841,N_16519,N_16601);
or U18842 (N_18842,N_17699,N_17277);
xnor U18843 (N_18843,N_17703,N_17054);
nand U18844 (N_18844,N_16835,N_17964);
nor U18845 (N_18845,N_17464,N_17726);
or U18846 (N_18846,N_16553,N_16614);
and U18847 (N_18847,N_17236,N_16556);
nand U18848 (N_18848,N_17280,N_17313);
xnor U18849 (N_18849,N_16902,N_17632);
or U18850 (N_18850,N_17954,N_17767);
nor U18851 (N_18851,N_17351,N_17115);
nand U18852 (N_18852,N_17130,N_17666);
nand U18853 (N_18853,N_17528,N_17037);
or U18854 (N_18854,N_17662,N_17702);
or U18855 (N_18855,N_17974,N_16810);
or U18856 (N_18856,N_17620,N_17717);
and U18857 (N_18857,N_16540,N_17866);
nor U18858 (N_18858,N_17717,N_16982);
xnor U18859 (N_18859,N_16908,N_17730);
nor U18860 (N_18860,N_17659,N_17845);
and U18861 (N_18861,N_16866,N_16608);
xnor U18862 (N_18862,N_17650,N_16706);
xor U18863 (N_18863,N_16991,N_16958);
nor U18864 (N_18864,N_16759,N_16894);
and U18865 (N_18865,N_16553,N_17107);
or U18866 (N_18866,N_17262,N_17464);
nor U18867 (N_18867,N_16648,N_17851);
or U18868 (N_18868,N_16779,N_17059);
or U18869 (N_18869,N_17985,N_16702);
and U18870 (N_18870,N_17305,N_17784);
nand U18871 (N_18871,N_17583,N_17591);
xor U18872 (N_18872,N_17099,N_17859);
nand U18873 (N_18873,N_17187,N_17129);
xor U18874 (N_18874,N_17780,N_16566);
nand U18875 (N_18875,N_16640,N_16961);
nand U18876 (N_18876,N_17512,N_17659);
nor U18877 (N_18877,N_17603,N_16598);
and U18878 (N_18878,N_16702,N_16753);
nand U18879 (N_18879,N_16610,N_17522);
nor U18880 (N_18880,N_17482,N_16859);
or U18881 (N_18881,N_17904,N_16677);
and U18882 (N_18882,N_17696,N_17991);
nor U18883 (N_18883,N_16768,N_16751);
or U18884 (N_18884,N_16755,N_17780);
and U18885 (N_18885,N_17766,N_17480);
xor U18886 (N_18886,N_16971,N_17983);
or U18887 (N_18887,N_17930,N_16891);
nand U18888 (N_18888,N_17472,N_17712);
or U18889 (N_18889,N_17060,N_17457);
xor U18890 (N_18890,N_17714,N_17671);
and U18891 (N_18891,N_17796,N_17822);
xor U18892 (N_18892,N_17929,N_17316);
nand U18893 (N_18893,N_16594,N_16596);
xor U18894 (N_18894,N_17108,N_16561);
and U18895 (N_18895,N_17896,N_16517);
and U18896 (N_18896,N_17525,N_17308);
nand U18897 (N_18897,N_17056,N_16881);
xnor U18898 (N_18898,N_16918,N_16982);
nand U18899 (N_18899,N_17534,N_16705);
nor U18900 (N_18900,N_16612,N_17156);
or U18901 (N_18901,N_17420,N_17441);
nor U18902 (N_18902,N_16799,N_17955);
or U18903 (N_18903,N_17204,N_17304);
xnor U18904 (N_18904,N_16788,N_17903);
and U18905 (N_18905,N_16792,N_16974);
nand U18906 (N_18906,N_17095,N_17389);
nand U18907 (N_18907,N_16981,N_16876);
xor U18908 (N_18908,N_16988,N_16894);
xnor U18909 (N_18909,N_16809,N_16889);
or U18910 (N_18910,N_16573,N_16896);
or U18911 (N_18911,N_17235,N_17026);
or U18912 (N_18912,N_17171,N_17515);
nand U18913 (N_18913,N_17124,N_17921);
nor U18914 (N_18914,N_17046,N_17664);
or U18915 (N_18915,N_17607,N_17673);
nor U18916 (N_18916,N_16636,N_16903);
xnor U18917 (N_18917,N_16571,N_17221);
xor U18918 (N_18918,N_17681,N_16530);
xor U18919 (N_18919,N_16843,N_16730);
or U18920 (N_18920,N_17879,N_16891);
nor U18921 (N_18921,N_17242,N_16974);
or U18922 (N_18922,N_17478,N_17144);
and U18923 (N_18923,N_16983,N_16550);
and U18924 (N_18924,N_17491,N_17931);
nand U18925 (N_18925,N_16597,N_17104);
nor U18926 (N_18926,N_17813,N_17067);
nor U18927 (N_18927,N_17332,N_16613);
nand U18928 (N_18928,N_16770,N_16860);
nand U18929 (N_18929,N_16794,N_16721);
xor U18930 (N_18930,N_16732,N_17624);
or U18931 (N_18931,N_16606,N_17954);
nor U18932 (N_18932,N_16656,N_17750);
nand U18933 (N_18933,N_16799,N_16903);
xor U18934 (N_18934,N_17710,N_16691);
or U18935 (N_18935,N_16782,N_17658);
and U18936 (N_18936,N_17070,N_17501);
nand U18937 (N_18937,N_17828,N_16735);
or U18938 (N_18938,N_16773,N_17267);
nor U18939 (N_18939,N_17204,N_17775);
nand U18940 (N_18940,N_17141,N_17888);
or U18941 (N_18941,N_16778,N_16983);
nor U18942 (N_18942,N_17845,N_17685);
or U18943 (N_18943,N_16501,N_17953);
or U18944 (N_18944,N_17490,N_17886);
or U18945 (N_18945,N_16837,N_16918);
and U18946 (N_18946,N_17211,N_17286);
nor U18947 (N_18947,N_17298,N_17929);
xnor U18948 (N_18948,N_16656,N_17044);
nand U18949 (N_18949,N_17618,N_17477);
nor U18950 (N_18950,N_17383,N_16893);
nand U18951 (N_18951,N_17887,N_16518);
nor U18952 (N_18952,N_17813,N_16712);
xor U18953 (N_18953,N_16665,N_17442);
nor U18954 (N_18954,N_17722,N_16541);
and U18955 (N_18955,N_17720,N_17581);
nand U18956 (N_18956,N_17789,N_16918);
nand U18957 (N_18957,N_16898,N_17262);
nand U18958 (N_18958,N_16529,N_17138);
nand U18959 (N_18959,N_17429,N_17957);
xnor U18960 (N_18960,N_17153,N_16693);
and U18961 (N_18961,N_17855,N_17261);
nand U18962 (N_18962,N_17826,N_17245);
nor U18963 (N_18963,N_17707,N_17832);
nand U18964 (N_18964,N_16679,N_17001);
xnor U18965 (N_18965,N_16849,N_17163);
nor U18966 (N_18966,N_16725,N_16840);
or U18967 (N_18967,N_16983,N_17608);
nor U18968 (N_18968,N_17489,N_17752);
nand U18969 (N_18969,N_16714,N_17425);
and U18970 (N_18970,N_16555,N_16814);
xor U18971 (N_18971,N_17894,N_16859);
xnor U18972 (N_18972,N_16863,N_17393);
xnor U18973 (N_18973,N_16607,N_17913);
or U18974 (N_18974,N_17412,N_17944);
xor U18975 (N_18975,N_17596,N_17694);
nand U18976 (N_18976,N_17456,N_16591);
nand U18977 (N_18977,N_16856,N_17927);
or U18978 (N_18978,N_17007,N_17531);
xnor U18979 (N_18979,N_17235,N_16673);
nand U18980 (N_18980,N_17333,N_17739);
nor U18981 (N_18981,N_17563,N_17024);
or U18982 (N_18982,N_17487,N_17332);
or U18983 (N_18983,N_17845,N_16788);
or U18984 (N_18984,N_16628,N_17907);
and U18985 (N_18985,N_17664,N_17936);
xor U18986 (N_18986,N_17754,N_16976);
xor U18987 (N_18987,N_17148,N_17612);
nand U18988 (N_18988,N_16508,N_16685);
xor U18989 (N_18989,N_16644,N_17516);
nand U18990 (N_18990,N_17458,N_17348);
xnor U18991 (N_18991,N_17282,N_17848);
or U18992 (N_18992,N_17885,N_17497);
and U18993 (N_18993,N_17610,N_16696);
xor U18994 (N_18994,N_16624,N_17451);
xnor U18995 (N_18995,N_17123,N_17280);
xor U18996 (N_18996,N_16537,N_17192);
nor U18997 (N_18997,N_17621,N_16961);
nor U18998 (N_18998,N_17440,N_17203);
or U18999 (N_18999,N_16630,N_17941);
nand U19000 (N_19000,N_17557,N_16678);
nand U19001 (N_19001,N_17748,N_17245);
nor U19002 (N_19002,N_16611,N_17718);
nor U19003 (N_19003,N_16690,N_16757);
xnor U19004 (N_19004,N_16508,N_17280);
nor U19005 (N_19005,N_17789,N_17443);
xnor U19006 (N_19006,N_17583,N_16858);
xor U19007 (N_19007,N_17692,N_16962);
nor U19008 (N_19008,N_17458,N_17451);
and U19009 (N_19009,N_17556,N_17326);
nand U19010 (N_19010,N_17142,N_16515);
or U19011 (N_19011,N_17898,N_17845);
xnor U19012 (N_19012,N_17596,N_17599);
xnor U19013 (N_19013,N_17461,N_17006);
nand U19014 (N_19014,N_17957,N_17345);
nand U19015 (N_19015,N_16745,N_16731);
xor U19016 (N_19016,N_16562,N_17014);
and U19017 (N_19017,N_17278,N_16726);
nand U19018 (N_19018,N_16901,N_16783);
nor U19019 (N_19019,N_17854,N_17441);
xnor U19020 (N_19020,N_17500,N_16642);
xnor U19021 (N_19021,N_17420,N_17046);
xnor U19022 (N_19022,N_17458,N_17907);
and U19023 (N_19023,N_17664,N_17186);
or U19024 (N_19024,N_17802,N_17151);
and U19025 (N_19025,N_17356,N_17262);
xnor U19026 (N_19026,N_16593,N_17930);
and U19027 (N_19027,N_17375,N_17706);
or U19028 (N_19028,N_17377,N_17331);
nor U19029 (N_19029,N_16868,N_16689);
or U19030 (N_19030,N_17946,N_17417);
nor U19031 (N_19031,N_16774,N_16893);
nor U19032 (N_19032,N_17633,N_16649);
and U19033 (N_19033,N_17508,N_17797);
nand U19034 (N_19034,N_17030,N_17038);
xnor U19035 (N_19035,N_17142,N_17998);
xnor U19036 (N_19036,N_16511,N_16617);
and U19037 (N_19037,N_17658,N_17934);
or U19038 (N_19038,N_16739,N_16945);
or U19039 (N_19039,N_17120,N_17602);
nor U19040 (N_19040,N_17765,N_16919);
or U19041 (N_19041,N_17185,N_17918);
and U19042 (N_19042,N_17128,N_17113);
xnor U19043 (N_19043,N_17487,N_17804);
or U19044 (N_19044,N_17747,N_17340);
and U19045 (N_19045,N_17749,N_17833);
or U19046 (N_19046,N_16652,N_17631);
and U19047 (N_19047,N_17163,N_17042);
and U19048 (N_19048,N_17374,N_16717);
or U19049 (N_19049,N_17864,N_17220);
nand U19050 (N_19050,N_17308,N_17935);
nor U19051 (N_19051,N_16940,N_17249);
nand U19052 (N_19052,N_16648,N_17418);
or U19053 (N_19053,N_17329,N_16768);
nand U19054 (N_19054,N_16594,N_17710);
nand U19055 (N_19055,N_17619,N_17080);
nand U19056 (N_19056,N_17446,N_17914);
or U19057 (N_19057,N_16617,N_16659);
nor U19058 (N_19058,N_17942,N_17450);
nand U19059 (N_19059,N_17922,N_17136);
or U19060 (N_19060,N_17865,N_16923);
nor U19061 (N_19061,N_17872,N_16722);
xor U19062 (N_19062,N_17617,N_17381);
or U19063 (N_19063,N_17331,N_17232);
nor U19064 (N_19064,N_17288,N_17549);
nor U19065 (N_19065,N_17148,N_17821);
xor U19066 (N_19066,N_17922,N_17613);
nor U19067 (N_19067,N_16588,N_17881);
or U19068 (N_19068,N_16685,N_17628);
and U19069 (N_19069,N_17919,N_16787);
nand U19070 (N_19070,N_17808,N_17229);
and U19071 (N_19071,N_16653,N_17472);
nor U19072 (N_19072,N_17906,N_17718);
xnor U19073 (N_19073,N_17984,N_17724);
nor U19074 (N_19074,N_17983,N_17092);
xor U19075 (N_19075,N_16602,N_16519);
nor U19076 (N_19076,N_17527,N_17209);
nand U19077 (N_19077,N_16720,N_17801);
xnor U19078 (N_19078,N_17618,N_17629);
and U19079 (N_19079,N_16792,N_17832);
nand U19080 (N_19080,N_17375,N_17962);
xor U19081 (N_19081,N_16688,N_17632);
nand U19082 (N_19082,N_16873,N_17378);
or U19083 (N_19083,N_17946,N_16759);
nor U19084 (N_19084,N_17500,N_17383);
nor U19085 (N_19085,N_17332,N_17717);
xnor U19086 (N_19086,N_16671,N_17896);
xnor U19087 (N_19087,N_16523,N_16543);
nand U19088 (N_19088,N_17353,N_17532);
nand U19089 (N_19089,N_17010,N_17668);
nor U19090 (N_19090,N_17846,N_16806);
and U19091 (N_19091,N_17543,N_17244);
and U19092 (N_19092,N_17009,N_17958);
and U19093 (N_19093,N_16518,N_17817);
xor U19094 (N_19094,N_17223,N_17189);
nor U19095 (N_19095,N_17481,N_17714);
or U19096 (N_19096,N_17369,N_17641);
xnor U19097 (N_19097,N_17067,N_17782);
nor U19098 (N_19098,N_16783,N_17238);
and U19099 (N_19099,N_17422,N_17553);
nor U19100 (N_19100,N_17285,N_17554);
nand U19101 (N_19101,N_17350,N_16747);
nor U19102 (N_19102,N_16967,N_16662);
nand U19103 (N_19103,N_17015,N_17011);
and U19104 (N_19104,N_16800,N_17303);
nor U19105 (N_19105,N_16537,N_17743);
xor U19106 (N_19106,N_17922,N_17706);
and U19107 (N_19107,N_17900,N_17157);
nor U19108 (N_19108,N_17411,N_16843);
nor U19109 (N_19109,N_17931,N_17324);
xor U19110 (N_19110,N_17245,N_17564);
and U19111 (N_19111,N_17417,N_16544);
xor U19112 (N_19112,N_17982,N_17820);
nand U19113 (N_19113,N_17030,N_17469);
or U19114 (N_19114,N_17426,N_17155);
or U19115 (N_19115,N_17566,N_17530);
nand U19116 (N_19116,N_16852,N_17953);
or U19117 (N_19117,N_17690,N_17838);
xnor U19118 (N_19118,N_17690,N_17705);
and U19119 (N_19119,N_16900,N_17833);
and U19120 (N_19120,N_17199,N_16624);
or U19121 (N_19121,N_17326,N_16799);
or U19122 (N_19122,N_17000,N_17033);
nor U19123 (N_19123,N_17316,N_17443);
and U19124 (N_19124,N_16895,N_17576);
nor U19125 (N_19125,N_16600,N_16783);
xor U19126 (N_19126,N_16560,N_17007);
nand U19127 (N_19127,N_17090,N_16817);
nand U19128 (N_19128,N_17832,N_17365);
or U19129 (N_19129,N_17292,N_17936);
and U19130 (N_19130,N_17933,N_17308);
and U19131 (N_19131,N_16925,N_17530);
and U19132 (N_19132,N_17742,N_17155);
and U19133 (N_19133,N_16698,N_17738);
nand U19134 (N_19134,N_17372,N_17389);
xor U19135 (N_19135,N_17358,N_16750);
or U19136 (N_19136,N_17523,N_17623);
and U19137 (N_19137,N_17617,N_16677);
nor U19138 (N_19138,N_17049,N_17579);
nor U19139 (N_19139,N_16701,N_17816);
nand U19140 (N_19140,N_17465,N_17538);
nand U19141 (N_19141,N_17158,N_17592);
nor U19142 (N_19142,N_17033,N_16947);
xnor U19143 (N_19143,N_17754,N_17298);
or U19144 (N_19144,N_16752,N_17890);
nand U19145 (N_19145,N_17924,N_17184);
nand U19146 (N_19146,N_16768,N_17211);
nand U19147 (N_19147,N_16859,N_16606);
and U19148 (N_19148,N_16717,N_17889);
xnor U19149 (N_19149,N_17060,N_17198);
nor U19150 (N_19150,N_17850,N_17091);
or U19151 (N_19151,N_16626,N_17591);
nand U19152 (N_19152,N_17754,N_17326);
nand U19153 (N_19153,N_16651,N_16890);
nor U19154 (N_19154,N_17901,N_17324);
xor U19155 (N_19155,N_17519,N_17939);
nand U19156 (N_19156,N_17126,N_17534);
nand U19157 (N_19157,N_16787,N_17639);
nor U19158 (N_19158,N_17899,N_17717);
nand U19159 (N_19159,N_17008,N_17241);
nand U19160 (N_19160,N_17075,N_17809);
and U19161 (N_19161,N_17297,N_17229);
nand U19162 (N_19162,N_16711,N_16675);
nand U19163 (N_19163,N_16743,N_16606);
or U19164 (N_19164,N_17107,N_17801);
or U19165 (N_19165,N_17294,N_16713);
or U19166 (N_19166,N_16969,N_17570);
and U19167 (N_19167,N_17416,N_16928);
or U19168 (N_19168,N_16645,N_17735);
and U19169 (N_19169,N_17006,N_17738);
nand U19170 (N_19170,N_17066,N_17514);
nor U19171 (N_19171,N_16735,N_17127);
or U19172 (N_19172,N_17057,N_17660);
xnor U19173 (N_19173,N_16969,N_17942);
xnor U19174 (N_19174,N_16971,N_17993);
and U19175 (N_19175,N_17092,N_17250);
and U19176 (N_19176,N_17791,N_17029);
xor U19177 (N_19177,N_17067,N_17494);
and U19178 (N_19178,N_17854,N_17658);
nor U19179 (N_19179,N_16841,N_17067);
or U19180 (N_19180,N_16922,N_16604);
xnor U19181 (N_19181,N_17544,N_16917);
nor U19182 (N_19182,N_17990,N_17769);
or U19183 (N_19183,N_17484,N_16813);
nor U19184 (N_19184,N_17945,N_17484);
nor U19185 (N_19185,N_16949,N_16527);
nand U19186 (N_19186,N_17583,N_17277);
nor U19187 (N_19187,N_17696,N_17961);
nand U19188 (N_19188,N_16867,N_17699);
and U19189 (N_19189,N_17760,N_17749);
nor U19190 (N_19190,N_17309,N_17941);
or U19191 (N_19191,N_16712,N_17538);
nand U19192 (N_19192,N_17685,N_17006);
or U19193 (N_19193,N_17034,N_17222);
nand U19194 (N_19194,N_16651,N_17580);
or U19195 (N_19195,N_17239,N_17827);
nand U19196 (N_19196,N_16865,N_17356);
and U19197 (N_19197,N_17912,N_17169);
or U19198 (N_19198,N_17613,N_17645);
xor U19199 (N_19199,N_17147,N_17310);
nor U19200 (N_19200,N_16626,N_17958);
nand U19201 (N_19201,N_16645,N_17602);
nor U19202 (N_19202,N_17625,N_17058);
and U19203 (N_19203,N_17085,N_17408);
and U19204 (N_19204,N_17433,N_17866);
nand U19205 (N_19205,N_17081,N_17980);
and U19206 (N_19206,N_17521,N_17482);
nor U19207 (N_19207,N_17958,N_16856);
nor U19208 (N_19208,N_17967,N_17550);
or U19209 (N_19209,N_17551,N_17867);
and U19210 (N_19210,N_17057,N_17806);
nor U19211 (N_19211,N_17327,N_17311);
nand U19212 (N_19212,N_17960,N_17828);
and U19213 (N_19213,N_16719,N_17795);
nand U19214 (N_19214,N_16720,N_17670);
xnor U19215 (N_19215,N_17779,N_17636);
nor U19216 (N_19216,N_17730,N_16566);
and U19217 (N_19217,N_16959,N_17031);
nor U19218 (N_19218,N_16837,N_17382);
nand U19219 (N_19219,N_17368,N_16609);
xnor U19220 (N_19220,N_16982,N_17628);
xnor U19221 (N_19221,N_17819,N_17907);
and U19222 (N_19222,N_17117,N_16777);
nand U19223 (N_19223,N_17420,N_16669);
nor U19224 (N_19224,N_17792,N_17406);
nor U19225 (N_19225,N_16710,N_17843);
xnor U19226 (N_19226,N_17811,N_17301);
and U19227 (N_19227,N_16569,N_16591);
nand U19228 (N_19228,N_17921,N_17118);
nor U19229 (N_19229,N_17181,N_17888);
or U19230 (N_19230,N_17784,N_17425);
nor U19231 (N_19231,N_17382,N_17904);
and U19232 (N_19232,N_17015,N_17574);
or U19233 (N_19233,N_17560,N_16754);
and U19234 (N_19234,N_17078,N_17351);
and U19235 (N_19235,N_17472,N_17926);
nor U19236 (N_19236,N_17885,N_16783);
nand U19237 (N_19237,N_17167,N_17609);
nor U19238 (N_19238,N_16726,N_16624);
or U19239 (N_19239,N_17378,N_16661);
nand U19240 (N_19240,N_17054,N_17062);
and U19241 (N_19241,N_17403,N_16532);
xnor U19242 (N_19242,N_17137,N_17000);
nand U19243 (N_19243,N_16798,N_17028);
nand U19244 (N_19244,N_17109,N_17253);
or U19245 (N_19245,N_17742,N_16561);
and U19246 (N_19246,N_17602,N_16734);
or U19247 (N_19247,N_16961,N_16544);
or U19248 (N_19248,N_17657,N_16611);
and U19249 (N_19249,N_17289,N_17020);
or U19250 (N_19250,N_17756,N_16674);
and U19251 (N_19251,N_16581,N_17291);
nand U19252 (N_19252,N_17186,N_17959);
or U19253 (N_19253,N_17618,N_17016);
nand U19254 (N_19254,N_16524,N_16873);
xnor U19255 (N_19255,N_17448,N_16647);
and U19256 (N_19256,N_16878,N_16818);
xor U19257 (N_19257,N_16639,N_17199);
and U19258 (N_19258,N_17738,N_16879);
nor U19259 (N_19259,N_17564,N_17477);
xnor U19260 (N_19260,N_17998,N_17310);
xnor U19261 (N_19261,N_16880,N_16637);
nor U19262 (N_19262,N_17391,N_17269);
xnor U19263 (N_19263,N_16588,N_17301);
and U19264 (N_19264,N_16897,N_17359);
nor U19265 (N_19265,N_16662,N_17361);
or U19266 (N_19266,N_17128,N_17725);
xor U19267 (N_19267,N_16761,N_17518);
nand U19268 (N_19268,N_17472,N_17053);
or U19269 (N_19269,N_16752,N_17672);
or U19270 (N_19270,N_17120,N_16828);
or U19271 (N_19271,N_17242,N_16684);
nor U19272 (N_19272,N_16572,N_17508);
xnor U19273 (N_19273,N_16741,N_17297);
xnor U19274 (N_19274,N_16579,N_16533);
or U19275 (N_19275,N_16751,N_16823);
and U19276 (N_19276,N_16673,N_17712);
or U19277 (N_19277,N_16869,N_16537);
nor U19278 (N_19278,N_17401,N_17061);
nor U19279 (N_19279,N_17239,N_17098);
nor U19280 (N_19280,N_17026,N_17077);
xnor U19281 (N_19281,N_17728,N_17623);
nand U19282 (N_19282,N_16727,N_16733);
or U19283 (N_19283,N_17936,N_17299);
nor U19284 (N_19284,N_17719,N_16859);
nor U19285 (N_19285,N_17432,N_17455);
or U19286 (N_19286,N_17383,N_17906);
nand U19287 (N_19287,N_17741,N_17848);
nand U19288 (N_19288,N_17979,N_16961);
and U19289 (N_19289,N_17446,N_17972);
nor U19290 (N_19290,N_16858,N_16689);
nand U19291 (N_19291,N_17725,N_17228);
nor U19292 (N_19292,N_17833,N_17995);
and U19293 (N_19293,N_17065,N_17840);
nor U19294 (N_19294,N_17915,N_17622);
xnor U19295 (N_19295,N_16653,N_17453);
xnor U19296 (N_19296,N_17711,N_16581);
nor U19297 (N_19297,N_17609,N_16820);
and U19298 (N_19298,N_17910,N_17300);
xor U19299 (N_19299,N_16920,N_17429);
and U19300 (N_19300,N_17513,N_17029);
nor U19301 (N_19301,N_17067,N_17097);
nand U19302 (N_19302,N_17092,N_16738);
or U19303 (N_19303,N_17976,N_16689);
nand U19304 (N_19304,N_17915,N_17954);
nand U19305 (N_19305,N_16780,N_17318);
nand U19306 (N_19306,N_17505,N_16791);
nand U19307 (N_19307,N_17831,N_17573);
nand U19308 (N_19308,N_16538,N_17480);
or U19309 (N_19309,N_16503,N_16616);
nand U19310 (N_19310,N_17455,N_17680);
nor U19311 (N_19311,N_17386,N_16736);
and U19312 (N_19312,N_17858,N_17664);
nor U19313 (N_19313,N_17242,N_16971);
nand U19314 (N_19314,N_17238,N_17418);
or U19315 (N_19315,N_17733,N_17573);
or U19316 (N_19316,N_17849,N_16936);
nand U19317 (N_19317,N_17954,N_17918);
or U19318 (N_19318,N_16786,N_17668);
nor U19319 (N_19319,N_16588,N_16802);
nor U19320 (N_19320,N_17244,N_17127);
or U19321 (N_19321,N_17621,N_17966);
nand U19322 (N_19322,N_17544,N_17150);
or U19323 (N_19323,N_16918,N_17453);
xnor U19324 (N_19324,N_17038,N_16717);
and U19325 (N_19325,N_17331,N_17429);
and U19326 (N_19326,N_17004,N_17235);
xor U19327 (N_19327,N_16657,N_17168);
and U19328 (N_19328,N_16510,N_17058);
nor U19329 (N_19329,N_16661,N_17814);
or U19330 (N_19330,N_17088,N_16576);
nand U19331 (N_19331,N_16975,N_17441);
nor U19332 (N_19332,N_17598,N_17061);
or U19333 (N_19333,N_16568,N_17253);
nor U19334 (N_19334,N_17636,N_16930);
or U19335 (N_19335,N_16849,N_16972);
xor U19336 (N_19336,N_16928,N_17454);
nor U19337 (N_19337,N_16592,N_17721);
nor U19338 (N_19338,N_17139,N_17403);
and U19339 (N_19339,N_17358,N_16808);
xor U19340 (N_19340,N_17122,N_17227);
nand U19341 (N_19341,N_17283,N_17580);
and U19342 (N_19342,N_17915,N_17853);
or U19343 (N_19343,N_17162,N_17530);
xor U19344 (N_19344,N_17658,N_17140);
or U19345 (N_19345,N_16996,N_16792);
and U19346 (N_19346,N_17617,N_17177);
or U19347 (N_19347,N_17552,N_17114);
xor U19348 (N_19348,N_17813,N_16796);
xnor U19349 (N_19349,N_17227,N_17767);
or U19350 (N_19350,N_17028,N_17041);
and U19351 (N_19351,N_16671,N_17081);
or U19352 (N_19352,N_17675,N_17274);
nor U19353 (N_19353,N_17329,N_16959);
or U19354 (N_19354,N_16673,N_17182);
or U19355 (N_19355,N_17916,N_17772);
xnor U19356 (N_19356,N_17556,N_17982);
nand U19357 (N_19357,N_17192,N_17069);
nor U19358 (N_19358,N_16694,N_17202);
nor U19359 (N_19359,N_17703,N_17218);
nand U19360 (N_19360,N_16689,N_17504);
or U19361 (N_19361,N_17035,N_16692);
nand U19362 (N_19362,N_16883,N_17590);
or U19363 (N_19363,N_16865,N_17740);
nor U19364 (N_19364,N_17626,N_17065);
nor U19365 (N_19365,N_17684,N_17810);
or U19366 (N_19366,N_16604,N_16916);
xnor U19367 (N_19367,N_17438,N_16550);
or U19368 (N_19368,N_16588,N_17803);
nor U19369 (N_19369,N_16985,N_16856);
nand U19370 (N_19370,N_17514,N_17827);
or U19371 (N_19371,N_17253,N_16910);
nor U19372 (N_19372,N_16559,N_17308);
and U19373 (N_19373,N_17025,N_17519);
xnor U19374 (N_19374,N_17398,N_16894);
nand U19375 (N_19375,N_17645,N_17796);
nand U19376 (N_19376,N_17293,N_16792);
xnor U19377 (N_19377,N_17141,N_17227);
nand U19378 (N_19378,N_17341,N_17062);
or U19379 (N_19379,N_17286,N_16635);
and U19380 (N_19380,N_17784,N_17355);
or U19381 (N_19381,N_16738,N_16964);
nand U19382 (N_19382,N_17741,N_17262);
nand U19383 (N_19383,N_17775,N_16815);
xnor U19384 (N_19384,N_16690,N_16610);
xnor U19385 (N_19385,N_17081,N_16600);
xor U19386 (N_19386,N_17110,N_16521);
nor U19387 (N_19387,N_17898,N_17191);
and U19388 (N_19388,N_17184,N_17960);
nand U19389 (N_19389,N_16831,N_17078);
nand U19390 (N_19390,N_17859,N_16920);
nor U19391 (N_19391,N_17971,N_17078);
and U19392 (N_19392,N_16803,N_16532);
xor U19393 (N_19393,N_17704,N_17678);
xnor U19394 (N_19394,N_16644,N_17458);
and U19395 (N_19395,N_17284,N_17051);
and U19396 (N_19396,N_16650,N_17532);
or U19397 (N_19397,N_16757,N_17491);
or U19398 (N_19398,N_16584,N_17036);
nor U19399 (N_19399,N_17945,N_17387);
and U19400 (N_19400,N_17045,N_17975);
and U19401 (N_19401,N_17398,N_16929);
and U19402 (N_19402,N_16834,N_17038);
xnor U19403 (N_19403,N_17326,N_16660);
or U19404 (N_19404,N_16739,N_16514);
xnor U19405 (N_19405,N_17147,N_17229);
and U19406 (N_19406,N_17735,N_17928);
nor U19407 (N_19407,N_16728,N_17046);
nand U19408 (N_19408,N_17298,N_17030);
nor U19409 (N_19409,N_17196,N_16720);
nor U19410 (N_19410,N_16755,N_17457);
nand U19411 (N_19411,N_17237,N_17211);
xnor U19412 (N_19412,N_17472,N_17798);
or U19413 (N_19413,N_17518,N_16889);
nand U19414 (N_19414,N_17716,N_16975);
or U19415 (N_19415,N_17185,N_17427);
or U19416 (N_19416,N_17856,N_16869);
and U19417 (N_19417,N_17399,N_17975);
or U19418 (N_19418,N_16508,N_16774);
nor U19419 (N_19419,N_16838,N_17392);
nand U19420 (N_19420,N_17659,N_17886);
nand U19421 (N_19421,N_17175,N_17506);
xnor U19422 (N_19422,N_17815,N_16854);
and U19423 (N_19423,N_17481,N_17937);
and U19424 (N_19424,N_17861,N_16846);
nor U19425 (N_19425,N_17474,N_17756);
nand U19426 (N_19426,N_17191,N_16961);
or U19427 (N_19427,N_17787,N_17166);
or U19428 (N_19428,N_16813,N_16924);
xnor U19429 (N_19429,N_17703,N_17251);
or U19430 (N_19430,N_17957,N_17588);
and U19431 (N_19431,N_16653,N_17843);
xnor U19432 (N_19432,N_17189,N_17420);
nand U19433 (N_19433,N_17026,N_17278);
and U19434 (N_19434,N_17981,N_17566);
nand U19435 (N_19435,N_16813,N_17147);
and U19436 (N_19436,N_17808,N_17571);
and U19437 (N_19437,N_17675,N_17106);
xnor U19438 (N_19438,N_16598,N_17098);
and U19439 (N_19439,N_17964,N_16616);
and U19440 (N_19440,N_16631,N_16944);
nand U19441 (N_19441,N_17867,N_17340);
and U19442 (N_19442,N_17690,N_17275);
xor U19443 (N_19443,N_17061,N_17437);
xnor U19444 (N_19444,N_16808,N_17194);
or U19445 (N_19445,N_17649,N_17948);
xnor U19446 (N_19446,N_16529,N_17954);
nand U19447 (N_19447,N_16703,N_16883);
xnor U19448 (N_19448,N_16918,N_17877);
or U19449 (N_19449,N_16667,N_16785);
and U19450 (N_19450,N_17446,N_17998);
nand U19451 (N_19451,N_17136,N_16984);
nor U19452 (N_19452,N_16662,N_17144);
nand U19453 (N_19453,N_16658,N_16627);
and U19454 (N_19454,N_16896,N_16671);
nand U19455 (N_19455,N_17417,N_16710);
or U19456 (N_19456,N_16880,N_17492);
and U19457 (N_19457,N_17415,N_16903);
nand U19458 (N_19458,N_17657,N_17699);
xnor U19459 (N_19459,N_17918,N_17362);
and U19460 (N_19460,N_17683,N_17186);
nand U19461 (N_19461,N_17829,N_17639);
xor U19462 (N_19462,N_17792,N_16957);
or U19463 (N_19463,N_17450,N_16660);
and U19464 (N_19464,N_17661,N_17583);
xnor U19465 (N_19465,N_16551,N_17209);
or U19466 (N_19466,N_17279,N_17155);
or U19467 (N_19467,N_17200,N_16975);
nor U19468 (N_19468,N_17720,N_16841);
and U19469 (N_19469,N_17170,N_16991);
and U19470 (N_19470,N_17667,N_17527);
and U19471 (N_19471,N_16528,N_17087);
xnor U19472 (N_19472,N_17766,N_16646);
nand U19473 (N_19473,N_16846,N_17304);
nand U19474 (N_19474,N_16666,N_17415);
nand U19475 (N_19475,N_17255,N_17018);
or U19476 (N_19476,N_17504,N_17951);
xor U19477 (N_19477,N_17820,N_17428);
and U19478 (N_19478,N_17957,N_17559);
and U19479 (N_19479,N_17886,N_16873);
and U19480 (N_19480,N_17925,N_17871);
xnor U19481 (N_19481,N_16927,N_16665);
xor U19482 (N_19482,N_16531,N_17396);
nor U19483 (N_19483,N_17495,N_17602);
or U19484 (N_19484,N_17285,N_17317);
nor U19485 (N_19485,N_17074,N_16791);
or U19486 (N_19486,N_17152,N_17160);
nor U19487 (N_19487,N_17964,N_17644);
xnor U19488 (N_19488,N_17059,N_17904);
and U19489 (N_19489,N_16726,N_16987);
and U19490 (N_19490,N_16944,N_16690);
nor U19491 (N_19491,N_17121,N_17967);
and U19492 (N_19492,N_16630,N_17461);
and U19493 (N_19493,N_17208,N_17190);
or U19494 (N_19494,N_16758,N_16854);
nand U19495 (N_19495,N_17451,N_17423);
and U19496 (N_19496,N_16500,N_17159);
xnor U19497 (N_19497,N_17524,N_17183);
xor U19498 (N_19498,N_17257,N_16533);
and U19499 (N_19499,N_17957,N_16878);
or U19500 (N_19500,N_19224,N_18724);
and U19501 (N_19501,N_18091,N_18036);
or U19502 (N_19502,N_18159,N_18321);
or U19503 (N_19503,N_18116,N_19375);
xnor U19504 (N_19504,N_18610,N_19373);
xnor U19505 (N_19505,N_19489,N_18692);
nor U19506 (N_19506,N_18951,N_19490);
or U19507 (N_19507,N_18837,N_18120);
nand U19508 (N_19508,N_19040,N_19353);
xnor U19509 (N_19509,N_19210,N_18217);
or U19510 (N_19510,N_18569,N_18126);
xnor U19511 (N_19511,N_19173,N_19300);
or U19512 (N_19512,N_18398,N_18288);
xor U19513 (N_19513,N_18051,N_19333);
nand U19514 (N_19514,N_18609,N_19116);
nand U19515 (N_19515,N_18850,N_18546);
and U19516 (N_19516,N_18156,N_18967);
xor U19517 (N_19517,N_19176,N_18028);
nand U19518 (N_19518,N_18515,N_18768);
or U19519 (N_19519,N_19365,N_18987);
or U19520 (N_19520,N_18138,N_19229);
or U19521 (N_19521,N_18928,N_18027);
xor U19522 (N_19522,N_19039,N_19352);
or U19523 (N_19523,N_18806,N_19385);
nor U19524 (N_19524,N_19114,N_19471);
or U19525 (N_19525,N_18137,N_18244);
or U19526 (N_19526,N_18705,N_19394);
nand U19527 (N_19527,N_18127,N_18170);
or U19528 (N_19528,N_18521,N_18256);
and U19529 (N_19529,N_18479,N_18102);
nor U19530 (N_19530,N_19052,N_18275);
xnor U19531 (N_19531,N_19191,N_19477);
or U19532 (N_19532,N_18016,N_19446);
nand U19533 (N_19533,N_18828,N_18079);
and U19534 (N_19534,N_19348,N_18838);
xnor U19535 (N_19535,N_18171,N_18240);
and U19536 (N_19536,N_19188,N_18961);
nand U19537 (N_19537,N_18442,N_19262);
or U19538 (N_19538,N_18204,N_19170);
and U19539 (N_19539,N_18225,N_18548);
nor U19540 (N_19540,N_18203,N_19174);
xor U19541 (N_19541,N_18110,N_18432);
xor U19542 (N_19542,N_18011,N_19053);
or U19543 (N_19543,N_18878,N_18501);
and U19544 (N_19544,N_19054,N_19387);
nor U19545 (N_19545,N_19214,N_18387);
xor U19546 (N_19546,N_18982,N_18884);
or U19547 (N_19547,N_18721,N_19302);
nor U19548 (N_19548,N_18318,N_19288);
and U19549 (N_19549,N_18090,N_18894);
or U19550 (N_19550,N_19343,N_18871);
xor U19551 (N_19551,N_18050,N_19131);
xor U19552 (N_19552,N_19480,N_19047);
nand U19553 (N_19553,N_18260,N_18731);
xnor U19554 (N_19554,N_18042,N_18931);
xor U19555 (N_19555,N_19185,N_19265);
nand U19556 (N_19556,N_18397,N_18346);
nor U19557 (N_19557,N_19140,N_18075);
and U19558 (N_19558,N_18406,N_18486);
xor U19559 (N_19559,N_18094,N_18816);
xor U19560 (N_19560,N_18697,N_18584);
xnor U19561 (N_19561,N_18617,N_19208);
and U19562 (N_19562,N_18269,N_19382);
nand U19563 (N_19563,N_18463,N_18445);
nand U19564 (N_19564,N_18134,N_18183);
nor U19565 (N_19565,N_18720,N_18762);
or U19566 (N_19566,N_18284,N_18498);
xnor U19567 (N_19567,N_19290,N_18349);
and U19568 (N_19568,N_18219,N_18458);
nor U19569 (N_19569,N_18934,N_18921);
nand U19570 (N_19570,N_19198,N_18258);
nor U19571 (N_19571,N_18930,N_18178);
nor U19572 (N_19572,N_18968,N_19487);
nand U19573 (N_19573,N_18020,N_18672);
nor U19574 (N_19574,N_19313,N_19318);
nand U19575 (N_19575,N_18497,N_18210);
xor U19576 (N_19576,N_18136,N_18162);
nand U19577 (N_19577,N_18723,N_18709);
and U19578 (N_19578,N_18339,N_18821);
or U19579 (N_19579,N_18427,N_19351);
or U19580 (N_19580,N_19000,N_18669);
and U19581 (N_19581,N_18952,N_18566);
or U19582 (N_19582,N_18543,N_18074);
or U19583 (N_19583,N_19150,N_18717);
xor U19584 (N_19584,N_18071,N_18531);
xnor U19585 (N_19585,N_18009,N_18022);
nand U19586 (N_19586,N_18511,N_18229);
xnor U19587 (N_19587,N_19400,N_19325);
nor U19588 (N_19588,N_19079,N_18940);
nor U19589 (N_19589,N_18337,N_19263);
and U19590 (N_19590,N_19127,N_18804);
and U19591 (N_19591,N_18603,N_19392);
nand U19592 (N_19592,N_19217,N_18765);
or U19593 (N_19593,N_18499,N_18274);
nand U19594 (N_19594,N_18294,N_18144);
nand U19595 (N_19595,N_18865,N_19416);
nand U19596 (N_19596,N_18508,N_19013);
xnor U19597 (N_19597,N_19247,N_19018);
nand U19598 (N_19598,N_18907,N_18914);
or U19599 (N_19599,N_18323,N_18909);
nor U19600 (N_19600,N_18629,N_19415);
and U19601 (N_19601,N_19323,N_18819);
and U19602 (N_19602,N_18446,N_18883);
xnor U19603 (N_19603,N_19028,N_18303);
nand U19604 (N_19604,N_18745,N_18836);
and U19605 (N_19605,N_18895,N_18668);
and U19606 (N_19606,N_19051,N_19164);
or U19607 (N_19607,N_19007,N_19494);
nand U19608 (N_19608,N_19275,N_18747);
and U19609 (N_19609,N_18946,N_18992);
or U19610 (N_19610,N_18786,N_19221);
nor U19611 (N_19611,N_18797,N_18621);
xnor U19612 (N_19612,N_18311,N_18021);
or U19613 (N_19613,N_19431,N_18718);
xnor U19614 (N_19614,N_19134,N_19468);
nor U19615 (N_19615,N_18250,N_18341);
and U19616 (N_19616,N_18333,N_18553);
nand U19617 (N_19617,N_18157,N_18176);
nor U19618 (N_19618,N_18695,N_19078);
nor U19619 (N_19619,N_18099,N_18848);
nor U19620 (N_19620,N_18018,N_19082);
xor U19621 (N_19621,N_19100,N_18782);
or U19622 (N_19622,N_18593,N_18614);
nand U19623 (N_19623,N_18000,N_18971);
nor U19624 (N_19624,N_18661,N_18866);
or U19625 (N_19625,N_18639,N_18007);
and U19626 (N_19626,N_18885,N_18017);
nand U19627 (N_19627,N_18057,N_19293);
nor U19628 (N_19628,N_18599,N_18759);
and U19629 (N_19629,N_18988,N_18033);
nand U19630 (N_19630,N_19278,N_19182);
or U19631 (N_19631,N_18361,N_19228);
nor U19632 (N_19632,N_18773,N_19239);
xnor U19633 (N_19633,N_19337,N_18925);
nand U19634 (N_19634,N_19199,N_18464);
or U19635 (N_19635,N_18409,N_19350);
nor U19636 (N_19636,N_19284,N_18932);
xor U19637 (N_19637,N_19080,N_18675);
xnor U19638 (N_19638,N_19447,N_18495);
and U19639 (N_19639,N_18671,N_18585);
or U19640 (N_19640,N_18182,N_18864);
nor U19641 (N_19641,N_19027,N_18518);
nor U19642 (N_19642,N_19335,N_18025);
and U19643 (N_19643,N_19042,N_18662);
nand U19644 (N_19644,N_18913,N_19465);
and U19645 (N_19645,N_19254,N_18522);
nand U19646 (N_19646,N_18840,N_18960);
or U19647 (N_19647,N_18935,N_18826);
or U19648 (N_19648,N_18350,N_18942);
and U19649 (N_19649,N_18264,N_18876);
and U19650 (N_19650,N_19336,N_18291);
and U19651 (N_19651,N_18010,N_18667);
xnor U19652 (N_19652,N_18257,N_18334);
or U19653 (N_19653,N_19488,N_18608);
nand U19654 (N_19654,N_18161,N_18381);
nor U19655 (N_19655,N_18282,N_19359);
nor U19656 (N_19656,N_18468,N_18135);
xor U19657 (N_19657,N_18820,N_18933);
or U19658 (N_19658,N_18410,N_18371);
and U19659 (N_19659,N_18435,N_18754);
xor U19660 (N_19660,N_19307,N_18858);
xnor U19661 (N_19661,N_18336,N_18873);
xor U19662 (N_19662,N_19376,N_18981);
or U19663 (N_19663,N_19380,N_18324);
xnor U19664 (N_19664,N_19384,N_18150);
or U19665 (N_19665,N_19259,N_18317);
nand U19666 (N_19666,N_18312,N_18173);
nand U19667 (N_19667,N_18038,N_18143);
nor U19668 (N_19668,N_18998,N_19237);
nand U19669 (N_19669,N_18474,N_18117);
xor U19670 (N_19670,N_18713,N_19094);
nor U19671 (N_19671,N_18802,N_18119);
and U19672 (N_19672,N_19156,N_18347);
and U19673 (N_19673,N_18460,N_18107);
and U19674 (N_19674,N_18148,N_19186);
nor U19675 (N_19675,N_18476,N_19092);
nand U19676 (N_19676,N_18947,N_19222);
or U19677 (N_19677,N_18646,N_18673);
nand U19678 (N_19678,N_18362,N_19363);
or U19679 (N_19679,N_18519,N_19440);
or U19680 (N_19680,N_19157,N_19364);
nor U19681 (N_19681,N_19383,N_18122);
xnor U19682 (N_19682,N_18073,N_18367);
xor U19683 (N_19683,N_18001,N_18623);
nand U19684 (N_19684,N_18375,N_18657);
nor U19685 (N_19685,N_19154,N_19061);
nor U19686 (N_19686,N_19104,N_18087);
nor U19687 (N_19687,N_19066,N_18910);
nor U19688 (N_19688,N_19169,N_18401);
nor U19689 (N_19689,N_18533,N_19171);
nand U19690 (N_19690,N_18253,N_19204);
or U19691 (N_19691,N_18287,N_18366);
nand U19692 (N_19692,N_19112,N_19123);
and U19693 (N_19693,N_18449,N_18627);
nor U19694 (N_19694,N_18979,N_18405);
nor U19695 (N_19695,N_18123,N_18354);
nor U19696 (N_19696,N_19202,N_19212);
or U19697 (N_19697,N_18554,N_19396);
and U19698 (N_19698,N_18165,N_18155);
and U19699 (N_19699,N_18927,N_18985);
xnor U19700 (N_19700,N_19009,N_18444);
xnor U19701 (N_19701,N_19160,N_18777);
xor U19702 (N_19702,N_18579,N_19417);
nor U19703 (N_19703,N_18564,N_18631);
nand U19704 (N_19704,N_19338,N_19441);
xnor U19705 (N_19705,N_18491,N_18844);
xnor U19706 (N_19706,N_19058,N_18535);
and U19707 (N_19707,N_19161,N_18887);
nand U19708 (N_19708,N_18413,N_19409);
nand U19709 (N_19709,N_18113,N_18950);
nand U19710 (N_19710,N_18624,N_18592);
xnor U19711 (N_19711,N_19143,N_19057);
xor U19712 (N_19712,N_18897,N_18456);
xnor U19713 (N_19713,N_19425,N_18562);
xor U19714 (N_19714,N_18748,N_18976);
xor U19715 (N_19715,N_18300,N_18310);
and U19716 (N_19716,N_18213,N_18746);
and U19717 (N_19717,N_19450,N_19461);
nand U19718 (N_19718,N_19277,N_19410);
xor U19719 (N_19719,N_19460,N_18728);
or U19720 (N_19720,N_19287,N_18849);
nand U19721 (N_19721,N_18023,N_19455);
or U19722 (N_19722,N_19495,N_18815);
xor U19723 (N_19723,N_18761,N_19452);
xor U19724 (N_19724,N_18586,N_18047);
or U19725 (N_19725,N_19218,N_18239);
and U19726 (N_19726,N_18466,N_18489);
nor U19727 (N_19727,N_18167,N_18649);
nand U19728 (N_19728,N_19436,N_18309);
nor U19729 (N_19729,N_19266,N_19141);
nand U19730 (N_19730,N_18039,N_19073);
nand U19731 (N_19731,N_19473,N_18228);
xnor U19732 (N_19732,N_18271,N_18902);
xor U19733 (N_19733,N_19038,N_19421);
xnor U19734 (N_19734,N_18083,N_18483);
and U19735 (N_19735,N_18642,N_19368);
xnor U19736 (N_19736,N_19304,N_18035);
or U19737 (N_19737,N_19366,N_19083);
xor U19738 (N_19738,N_18687,N_18899);
nor U19739 (N_19739,N_18049,N_18359);
xnor U19740 (N_19740,N_18787,N_19250);
xor U19741 (N_19741,N_19085,N_18212);
nor U19742 (N_19742,N_18360,N_18189);
xnor U19743 (N_19743,N_18776,N_18265);
and U19744 (N_19744,N_18622,N_18041);
or U19745 (N_19745,N_18395,N_18106);
nand U19746 (N_19746,N_18357,N_19005);
xnor U19747 (N_19747,N_18246,N_18529);
or U19748 (N_19748,N_19474,N_19068);
or U19749 (N_19749,N_19055,N_19379);
or U19750 (N_19750,N_18070,N_18740);
xnor U19751 (N_19751,N_18475,N_19200);
or U19752 (N_19752,N_19231,N_18462);
nand U19753 (N_19753,N_18735,N_18948);
and U19754 (N_19754,N_19483,N_18438);
nand U19755 (N_19755,N_18683,N_19469);
and U19756 (N_19756,N_18054,N_19486);
xor U19757 (N_19757,N_19152,N_18602);
xnor U19758 (N_19758,N_19391,N_18450);
or U19759 (N_19759,N_18242,N_19470);
and U19760 (N_19760,N_19482,N_18289);
or U19761 (N_19761,N_18571,N_18764);
nand U19762 (N_19762,N_18874,N_19330);
or U19763 (N_19763,N_18412,N_18175);
nor U19764 (N_19764,N_19306,N_18296);
xor U19765 (N_19765,N_18216,N_19423);
nand U19766 (N_19766,N_18984,N_18549);
nor U19767 (N_19767,N_19220,N_19075);
xor U19768 (N_19768,N_18612,N_18630);
nand U19769 (N_19769,N_18280,N_19479);
nand U19770 (N_19770,N_18986,N_18772);
or U19771 (N_19771,N_19476,N_19227);
nand U19772 (N_19772,N_19091,N_18898);
and U19773 (N_19773,N_18637,N_18506);
nor U19774 (N_19774,N_18488,N_19120);
nand U19775 (N_19775,N_18139,N_18513);
xnor U19776 (N_19776,N_19426,N_18243);
xnor U19777 (N_19777,N_18516,N_19126);
nor U19778 (N_19778,N_19438,N_18140);
xor U19779 (N_19779,N_19133,N_18537);
nor U19780 (N_19780,N_18108,N_19301);
xor U19781 (N_19781,N_18185,N_18852);
nor U19782 (N_19782,N_18390,N_18538);
nor U19783 (N_19783,N_18903,N_18251);
nand U19784 (N_19784,N_19031,N_19360);
nand U19785 (N_19785,N_18338,N_18247);
or U19786 (N_19786,N_18635,N_18812);
or U19787 (N_19787,N_19044,N_18040);
xnor U19788 (N_19788,N_18975,N_18404);
nor U19789 (N_19789,N_19475,N_18187);
or U19790 (N_19790,N_18358,N_18520);
nand U19791 (N_19791,N_19095,N_18965);
xor U19792 (N_19792,N_18620,N_18419);
or U19793 (N_19793,N_19015,N_18972);
and U19794 (N_19794,N_18158,N_18859);
nand U19795 (N_19795,N_19491,N_18278);
nor U19796 (N_19796,N_19084,N_18613);
or U19797 (N_19797,N_18273,N_18188);
and U19798 (N_19798,N_18417,N_19175);
or U19799 (N_19799,N_18628,N_19060);
nor U19800 (N_19800,N_18313,N_19187);
or U19801 (N_19801,N_18077,N_18149);
xnor U19802 (N_19802,N_19260,N_18220);
nand U19803 (N_19803,N_18693,N_18340);
xnor U19804 (N_19804,N_19381,N_19129);
nor U19805 (N_19805,N_18722,N_18550);
or U19806 (N_19806,N_18790,N_19178);
nand U19807 (N_19807,N_18307,N_18231);
xnor U19808 (N_19808,N_19388,N_18414);
or U19809 (N_19809,N_19011,N_18365);
xnor U19810 (N_19810,N_19430,N_18904);
xnor U19811 (N_19811,N_18298,N_18532);
nor U19812 (N_19812,N_18084,N_19238);
nand U19813 (N_19813,N_19063,N_18710);
or U19814 (N_19814,N_18238,N_19451);
or U19815 (N_19815,N_18104,N_18392);
nor U19816 (N_19816,N_18407,N_19132);
and U19817 (N_19817,N_18774,N_18378);
nor U19818 (N_19818,N_18180,N_19189);
or U19819 (N_19819,N_19349,N_18861);
nand U19820 (N_19820,N_18959,N_18448);
nand U19821 (N_19821,N_18095,N_18785);
nor U19822 (N_19822,N_18372,N_18207);
xor U19823 (N_19823,N_18201,N_18916);
xor U19824 (N_19824,N_19086,N_18262);
nand U19825 (N_19825,N_18974,N_18997);
xnor U19826 (N_19826,N_18478,N_18043);
xnor U19827 (N_19827,N_18736,N_19089);
nor U19828 (N_19828,N_19096,N_18425);
nor U19829 (N_19829,N_18461,N_18955);
nor U19830 (N_19830,N_18817,N_18471);
nor U19831 (N_19831,N_19032,N_19233);
and U19832 (N_19832,N_19101,N_18315);
and U19833 (N_19833,N_19347,N_18936);
nand U19834 (N_19834,N_19093,N_18174);
nand U19835 (N_19835,N_18026,N_18632);
nor U19836 (N_19836,N_19340,N_18682);
or U19837 (N_19837,N_19026,N_18744);
or U19838 (N_19838,N_18922,N_18918);
nor U19839 (N_19839,N_18781,N_19070);
nand U19840 (N_19840,N_19420,N_18293);
nor U19841 (N_19841,N_18160,N_18388);
and U19842 (N_19842,N_18666,N_19215);
and U19843 (N_19843,N_19294,N_18648);
and U19844 (N_19844,N_18002,N_18245);
nor U19845 (N_19845,N_18380,N_18956);
xor U19846 (N_19846,N_18373,N_19458);
nand U19847 (N_19847,N_18128,N_19484);
nand U19848 (N_19848,N_18943,N_19295);
nor U19849 (N_19849,N_18467,N_18881);
or U19850 (N_19850,N_18830,N_18939);
nand U19851 (N_19851,N_19168,N_19326);
xor U19852 (N_19852,N_19371,N_19356);
xnor U19853 (N_19853,N_19397,N_18004);
or U19854 (N_19854,N_19370,N_18568);
and U19855 (N_19855,N_18941,N_19201);
nand U19856 (N_19856,N_19405,N_18485);
or U19857 (N_19857,N_18575,N_18222);
xor U19858 (N_19858,N_19286,N_19243);
or U19859 (N_19859,N_19264,N_18527);
nor U19860 (N_19860,N_18330,N_18069);
nor U19861 (N_19861,N_19454,N_18302);
or U19862 (N_19862,N_18196,N_18580);
xor U19863 (N_19863,N_19437,N_19485);
or U19864 (N_19864,N_19322,N_18115);
nand U19865 (N_19865,N_18560,N_19435);
nand U19866 (N_19866,N_18044,N_18551);
xor U19867 (N_19867,N_18591,N_19401);
or U19868 (N_19868,N_19088,N_18389);
or U19869 (N_19869,N_18429,N_19390);
nor U19870 (N_19870,N_19308,N_18536);
or U19871 (N_19871,N_18234,N_19213);
nor U19872 (N_19872,N_18376,N_18507);
and U19873 (N_19873,N_18825,N_18784);
nand U19874 (N_19874,N_18594,N_18211);
and U19875 (N_19875,N_18472,N_19367);
and U19876 (N_19876,N_19389,N_18465);
nor U19877 (N_19877,N_18086,N_18232);
or U19878 (N_19878,N_18048,N_18879);
and U19879 (N_19879,N_18767,N_18872);
and U19880 (N_19880,N_18920,N_18595);
nand U19881 (N_19881,N_19466,N_18810);
xor U19882 (N_19882,N_18712,N_19464);
nand U19883 (N_19883,N_19179,N_18494);
nor U19884 (N_19884,N_18607,N_18556);
and U19885 (N_19885,N_18651,N_19177);
xor U19886 (N_19886,N_19022,N_19050);
and U19887 (N_19887,N_19107,N_18793);
nand U19888 (N_19888,N_19180,N_18418);
or U19889 (N_19889,N_18823,N_18809);
or U19890 (N_19890,N_19244,N_18750);
nor U19891 (N_19891,N_18072,N_18578);
or U19892 (N_19892,N_19467,N_18124);
nor U19893 (N_19893,N_19166,N_18345);
nand U19894 (N_19894,N_18698,N_19076);
xor U19895 (N_19895,N_18443,N_18484);
xnor U19896 (N_19896,N_18062,N_19339);
and U19897 (N_19897,N_18685,N_18295);
or U19898 (N_19898,N_18689,N_18179);
nor U19899 (N_19899,N_18431,N_18857);
or U19900 (N_19900,N_18800,N_18514);
nand U19901 (N_19901,N_18473,N_18202);
xor U19902 (N_19902,N_18868,N_18061);
nand U19903 (N_19903,N_18905,N_18596);
xor U19904 (N_19904,N_18915,N_19422);
or U19905 (N_19905,N_19269,N_19002);
xor U19906 (N_19906,N_18638,N_18386);
or U19907 (N_19907,N_18455,N_19117);
xor U19908 (N_19908,N_19404,N_18342);
nor U19909 (N_19909,N_18891,N_18803);
nand U19910 (N_19910,N_19130,N_18908);
and U19911 (N_19911,N_18290,N_18098);
and U19912 (N_19912,N_18503,N_18394);
nor U19913 (N_19913,N_19167,N_18964);
xor U19914 (N_19914,N_19449,N_19358);
nor U19915 (N_19915,N_19147,N_18487);
nand U19916 (N_19916,N_19443,N_19025);
nand U19917 (N_19917,N_19261,N_18991);
nor U19918 (N_19918,N_18132,N_18517);
xnor U19919 (N_19919,N_18558,N_18370);
nor U19920 (N_19920,N_18655,N_18436);
nand U19921 (N_19921,N_19242,N_18319);
xnor U19922 (N_19922,N_19030,N_18919);
or U19923 (N_19923,N_19297,N_19105);
nor U19924 (N_19924,N_18270,N_19142);
xor U19925 (N_19925,N_19008,N_18082);
nor U19926 (N_19926,N_19045,N_19273);
and U19927 (N_19927,N_18423,N_18272);
xnor U19928 (N_19928,N_18996,N_19069);
xor U19929 (N_19929,N_18500,N_18078);
and U19930 (N_19930,N_19241,N_19357);
or U19931 (N_19931,N_18505,N_18525);
nand U19932 (N_19932,N_18882,N_18654);
or U19933 (N_19933,N_18588,N_18818);
xnor U19934 (N_19934,N_19151,N_18055);
or U19935 (N_19935,N_18572,N_18215);
and U19936 (N_19936,N_18308,N_18194);
nor U19937 (N_19937,N_18428,N_18066);
or U19938 (N_19938,N_18912,N_19046);
nor U19939 (N_19939,N_18382,N_18037);
nand U19940 (N_19940,N_19492,N_18343);
and U19941 (N_19941,N_18733,N_19428);
xnor U19942 (N_19942,N_18197,N_18154);
nor U19943 (N_19943,N_18890,N_18938);
xnor U19944 (N_19944,N_18730,N_19344);
nor U19945 (N_19945,N_19226,N_18065);
nand U19946 (N_19946,N_19434,N_18177);
xor U19947 (N_19947,N_18316,N_18640);
or U19948 (N_19948,N_18670,N_18958);
nand U19949 (N_19949,N_18068,N_18147);
or U19950 (N_19950,N_19408,N_18034);
xnor U19951 (N_19951,N_18625,N_18510);
and U19952 (N_19952,N_19115,N_18504);
or U19953 (N_19953,N_19403,N_18853);
or U19954 (N_19954,N_18512,N_18542);
or U19955 (N_19955,N_18663,N_19109);
or U19956 (N_19956,N_18755,N_18589);
nand U19957 (N_19957,N_18453,N_18377);
nor U19958 (N_19958,N_18766,N_19206);
xor U19959 (N_19959,N_18681,N_18841);
or U19960 (N_19960,N_19271,N_18191);
xnor U19961 (N_19961,N_19499,N_18129);
nand U19962 (N_19962,N_19258,N_18252);
or U19963 (N_19963,N_19209,N_19125);
or U19964 (N_19964,N_18969,N_18598);
nand U19965 (N_19965,N_19412,N_19236);
or U19966 (N_19966,N_19194,N_18297);
nand U19967 (N_19967,N_19299,N_18164);
and U19968 (N_19968,N_18374,N_19327);
nand U19969 (N_19969,N_19372,N_18186);
nand U19970 (N_19970,N_18949,N_18798);
nor U19971 (N_19971,N_19137,N_18805);
or U19972 (N_19972,N_19081,N_18335);
xnor U19973 (N_19973,N_18081,N_18530);
and U19974 (N_19974,N_19362,N_18875);
xor U19975 (N_19975,N_18541,N_18353);
nand U19976 (N_19976,N_19149,N_18643);
nor U19977 (N_19977,N_18105,N_19004);
or U19978 (N_19978,N_18656,N_18789);
or U19979 (N_19979,N_18699,N_19291);
nor U19980 (N_19980,N_19424,N_19190);
nor U19981 (N_19981,N_18788,N_18711);
xor U19982 (N_19982,N_18408,N_19034);
and U19983 (N_19983,N_19249,N_19111);
or U19984 (N_19984,N_19378,N_18808);
nand U19985 (N_19985,N_19399,N_18304);
or U19986 (N_19986,N_18688,N_19234);
nand U19987 (N_19987,N_18056,N_19270);
nand U19988 (N_19988,N_18230,N_18109);
nand U19989 (N_19989,N_19138,N_19496);
or U19990 (N_19990,N_18565,N_18714);
nand U19991 (N_19991,N_18103,N_19312);
and U19992 (N_19992,N_18118,N_18402);
nand U19993 (N_19993,N_18901,N_18328);
or U19994 (N_19994,N_18753,N_19110);
xor U19995 (N_19995,N_18980,N_18172);
xor U19996 (N_19996,N_18329,N_18970);
or U19997 (N_19997,N_18605,N_19145);
or U19998 (N_19998,N_19163,N_19225);
nand U19999 (N_19999,N_19498,N_19049);
xor U20000 (N_20000,N_18719,N_19016);
and U20001 (N_20001,N_18888,N_18600);
xor U20002 (N_20002,N_18421,N_18814);
and U20003 (N_20003,N_18561,N_18824);
nand U20004 (N_20004,N_18707,N_18647);
nor U20005 (N_20005,N_18032,N_19102);
nor U20006 (N_20006,N_18917,N_19497);
xnor U20007 (N_20007,N_19248,N_18771);
nor U20008 (N_20008,N_18058,N_19087);
and U20009 (N_20009,N_19321,N_18769);
or U20010 (N_20010,N_18141,N_18447);
and U20011 (N_20011,N_19159,N_18944);
and U20012 (N_20012,N_19153,N_18259);
and U20013 (N_20013,N_18080,N_18540);
or U20014 (N_20014,N_18660,N_18101);
nand U20015 (N_20015,N_18223,N_18851);
nand U20016 (N_20016,N_18827,N_18459);
nand U20017 (N_20017,N_19329,N_18100);
and U20018 (N_20018,N_18440,N_18854);
xnor U20019 (N_20019,N_18552,N_19398);
nand U20020 (N_20020,N_19433,N_18792);
xnor U20021 (N_20021,N_19230,N_19135);
nand U20022 (N_20022,N_18325,N_19314);
or U20023 (N_20023,N_19256,N_19246);
or U20024 (N_20024,N_18439,N_18999);
or U20025 (N_20025,N_18758,N_18583);
nand U20026 (N_20026,N_18779,N_18995);
nand U20027 (N_20027,N_19041,N_18775);
nand U20028 (N_20028,N_19012,N_18701);
xor U20029 (N_20029,N_19067,N_18470);
nor U20030 (N_20030,N_18152,N_18426);
nand U20031 (N_20031,N_19207,N_18870);
or U20032 (N_20032,N_18266,N_18945);
and U20033 (N_20033,N_18254,N_18749);
nor U20034 (N_20034,N_19320,N_18833);
nand U20035 (N_20035,N_18184,N_18807);
or U20036 (N_20036,N_19411,N_19033);
xnor U20037 (N_20037,N_18725,N_19282);
or U20038 (N_20038,N_18422,N_18292);
and U20039 (N_20039,N_18249,N_18433);
xor U20040 (N_20040,N_18235,N_18559);
nand U20041 (N_20041,N_19144,N_18142);
xor U20042 (N_20042,N_18005,N_19283);
and U20043 (N_20043,N_18469,N_18299);
xnor U20044 (N_20044,N_19193,N_18570);
xnor U20045 (N_20045,N_18834,N_19106);
nor U20046 (N_20046,N_18702,N_19128);
or U20047 (N_20047,N_19442,N_18524);
or U20048 (N_20048,N_18121,N_18963);
or U20049 (N_20049,N_18990,N_18633);
nor U20050 (N_20050,N_18839,N_19406);
and U20051 (N_20051,N_18163,N_18477);
nand U20052 (N_20052,N_19219,N_18153);
or U20053 (N_20053,N_19303,N_18146);
xnor U20054 (N_20054,N_18261,N_18348);
nor U20055 (N_20055,N_19341,N_18190);
and U20056 (N_20056,N_18855,N_18399);
or U20057 (N_20057,N_18653,N_18544);
and U20058 (N_20058,N_18658,N_18973);
xor U20059 (N_20059,N_19478,N_18678);
or U20060 (N_20060,N_19407,N_19311);
or U20061 (N_20061,N_19457,N_19146);
and U20062 (N_20062,N_18267,N_18641);
and U20063 (N_20063,N_18218,N_18856);
nor U20064 (N_20064,N_19090,N_19418);
nand U20065 (N_20065,N_18659,N_18906);
xor U20066 (N_20066,N_19253,N_19232);
xnor U20067 (N_20067,N_18130,N_18411);
nor U20068 (N_20068,N_18539,N_18236);
and U20069 (N_20069,N_18024,N_18923);
nor U20070 (N_20070,N_18966,N_19427);
or U20071 (N_20071,N_18555,N_18111);
nor U20072 (N_20072,N_19334,N_19315);
or U20073 (N_20073,N_18567,N_18863);
nor U20074 (N_20074,N_18014,N_19098);
or U20075 (N_20075,N_18706,N_18114);
and U20076 (N_20076,N_19172,N_18030);
nand U20077 (N_20077,N_18618,N_18193);
xnor U20078 (N_20078,N_19310,N_18794);
nand U20079 (N_20079,N_18420,N_18994);
xor U20080 (N_20080,N_18604,N_18703);
nor U20081 (N_20081,N_19001,N_18509);
xnor U20082 (N_20082,N_18112,N_19071);
and U20083 (N_20083,N_18795,N_18208);
or U20084 (N_20084,N_19064,N_18125);
nand U20085 (N_20085,N_18206,N_19139);
xor U20086 (N_20086,N_18680,N_18492);
or U20087 (N_20087,N_18780,N_18214);
xnor U20088 (N_20088,N_19472,N_19413);
xor U20089 (N_20089,N_18481,N_18332);
or U20090 (N_20090,N_18285,N_19289);
or U20091 (N_20091,N_19023,N_18209);
nor U20092 (N_20092,N_18277,N_19056);
nor U20093 (N_20093,N_18846,N_18089);
or U20094 (N_20094,N_18351,N_19124);
and U20095 (N_20095,N_19155,N_19453);
xnor U20096 (N_20096,N_18224,N_18482);
nor U20097 (N_20097,N_18783,N_18847);
or U20098 (N_20098,N_18911,N_18181);
nor U20099 (N_20099,N_19223,N_18480);
nor U20100 (N_20100,N_19374,N_18822);
and U20101 (N_20101,N_18493,N_19342);
nor U20102 (N_20102,N_18327,N_18796);
nand U20103 (N_20103,N_18241,N_18726);
and U20104 (N_20104,N_18989,N_19035);
nand U20105 (N_20105,N_18029,N_19059);
xnor U20106 (N_20106,N_19216,N_18364);
and U20107 (N_20107,N_18742,N_19386);
nor U20108 (N_20108,N_19165,N_19245);
nor U20109 (N_20109,N_19196,N_18093);
nor U20110 (N_20110,N_18133,N_19037);
nor U20111 (N_20111,N_18665,N_18835);
or U20112 (N_20112,N_18145,N_19279);
nand U20113 (N_20113,N_18396,N_18845);
and U20114 (N_20114,N_18752,N_18059);
nand U20115 (N_20115,N_18019,N_18770);
nand U20116 (N_20116,N_18322,N_19108);
nor U20117 (N_20117,N_18169,N_19024);
nand U20118 (N_20118,N_19317,N_18451);
xnor U20119 (N_20119,N_18031,N_18526);
and U20120 (N_20120,N_18636,N_18199);
xnor U20121 (N_20121,N_19072,N_18060);
nor U20122 (N_20122,N_18233,N_18756);
and U20123 (N_20123,N_18743,N_19331);
nor U20124 (N_20124,N_18227,N_18502);
xnor U20125 (N_20125,N_19240,N_18192);
xor U20126 (N_20126,N_18587,N_18403);
and U20127 (N_20127,N_19235,N_19445);
nor U20128 (N_20128,N_18652,N_18434);
and U20129 (N_20129,N_19077,N_19393);
xor U20130 (N_20130,N_19113,N_19065);
nor U20131 (N_20131,N_18715,N_18331);
xnor U20132 (N_20132,N_19017,N_18097);
and U20133 (N_20133,N_19103,N_18811);
and U20134 (N_20134,N_18926,N_18619);
and U20135 (N_20135,N_19014,N_18385);
xnor U20136 (N_20136,N_19395,N_18283);
or U20137 (N_20137,N_19481,N_19121);
and U20138 (N_20138,N_18993,N_18813);
xor U20139 (N_20139,N_18320,N_18674);
xor U20140 (N_20140,N_19205,N_19043);
or U20141 (N_20141,N_18168,N_18574);
or U20142 (N_20142,N_18581,N_19402);
nor U20143 (N_20143,N_18355,N_18729);
nand U20144 (N_20144,N_18067,N_18008);
and U20145 (N_20145,N_18650,N_19119);
nor U20146 (N_20146,N_18843,N_18573);
nand U20147 (N_20147,N_18053,N_18741);
nor U20148 (N_20148,N_18221,N_19274);
nor U20149 (N_20149,N_19324,N_19148);
nand U20150 (N_20150,N_19019,N_18255);
xnor U20151 (N_20151,N_18978,N_18611);
nand U20152 (N_20152,N_18727,N_18195);
and U20153 (N_20153,N_18064,N_19020);
nor U20154 (N_20154,N_18454,N_18237);
nand U20155 (N_20155,N_18676,N_19292);
nand U20156 (N_20156,N_18305,N_18739);
and U20157 (N_20157,N_18791,N_18937);
nand U20158 (N_20158,N_18557,N_19251);
nor U20159 (N_20159,N_18679,N_19118);
and U20160 (N_20160,N_18896,N_19281);
nand U20161 (N_20161,N_18576,N_18778);
xnor U20162 (N_20162,N_18344,N_19162);
and U20163 (N_20163,N_19328,N_18738);
and U20164 (N_20164,N_18226,N_18634);
nand U20165 (N_20165,N_18352,N_19298);
and U20166 (N_20166,N_18799,N_19462);
nor U20167 (N_20167,N_18248,N_18760);
and U20168 (N_20168,N_19355,N_18953);
and U20169 (N_20169,N_18708,N_19316);
xor U20170 (N_20170,N_18301,N_18046);
or U20171 (N_20171,N_19272,N_19197);
nor U20172 (N_20172,N_18957,N_18877);
nor U20173 (N_20173,N_18045,N_19346);
and U20174 (N_20174,N_19448,N_18306);
nand U20175 (N_20175,N_18424,N_18088);
nand U20176 (N_20176,N_18684,N_19010);
and U20177 (N_20177,N_18601,N_18626);
nand U20178 (N_20178,N_19429,N_19463);
nand U20179 (N_20179,N_18694,N_19192);
and U20180 (N_20180,N_18400,N_18085);
nand U20181 (N_20181,N_19136,N_18716);
or U20182 (N_20182,N_18691,N_18279);
nor U20183 (N_20183,N_18954,N_18889);
or U20184 (N_20184,N_18862,N_18368);
nor U20185 (N_20185,N_19195,N_18384);
nor U20186 (N_20186,N_19432,N_19048);
and U20187 (N_20187,N_19493,N_18151);
xor U20188 (N_20188,N_18983,N_19036);
xor U20189 (N_20189,N_18416,N_18131);
nand U20190 (N_20190,N_19319,N_18391);
nand U20191 (N_20191,N_19280,N_18496);
xor U20192 (N_20192,N_19183,N_19257);
and U20193 (N_20193,N_18457,N_19305);
and U20194 (N_20194,N_18052,N_18686);
xor U20195 (N_20195,N_19296,N_18924);
or U20196 (N_20196,N_18880,N_18892);
nand U20197 (N_20197,N_18616,N_19332);
nor U20198 (N_20198,N_18013,N_19345);
and U20199 (N_20199,N_18867,N_19377);
nor U20200 (N_20200,N_18096,N_19099);
or U20201 (N_20201,N_18523,N_19003);
and U20202 (N_20202,N_18363,N_18452);
and U20203 (N_20203,N_18962,N_18757);
nor U20204 (N_20204,N_19439,N_18547);
nand U20205 (N_20205,N_18886,N_18198);
or U20206 (N_20206,N_18200,N_18860);
nand U20207 (N_20207,N_18166,N_18801);
nor U20208 (N_20208,N_18751,N_18700);
nand U20209 (N_20209,N_18829,N_18430);
and U20210 (N_20210,N_18534,N_18763);
nand U20211 (N_20211,N_18929,N_19276);
and U20212 (N_20212,N_18379,N_18383);
and U20213 (N_20213,N_19122,N_19285);
nand U20214 (N_20214,N_18076,N_18893);
xor U20215 (N_20215,N_19181,N_18900);
nor U20216 (N_20216,N_18006,N_18012);
nand U20217 (N_20217,N_18545,N_19252);
xor U20218 (N_20218,N_18977,N_19006);
nor U20219 (N_20219,N_19361,N_18696);
and U20220 (N_20220,N_19029,N_18582);
and U20221 (N_20221,N_18644,N_18326);
and U20222 (N_20222,N_18356,N_18314);
and U20223 (N_20223,N_18577,N_18563);
xor U20224 (N_20224,N_19021,N_18590);
nand U20225 (N_20225,N_18732,N_19184);
or U20226 (N_20226,N_18205,N_18734);
nand U20227 (N_20227,N_18606,N_19158);
nand U20228 (N_20228,N_18690,N_18003);
nand U20229 (N_20229,N_18268,N_19097);
xor U20230 (N_20230,N_19354,N_19203);
nor U20231 (N_20231,N_18645,N_18597);
and U20232 (N_20232,N_18869,N_19255);
xor U20233 (N_20233,N_18528,N_19309);
and U20234 (N_20234,N_18063,N_18831);
or U20235 (N_20235,N_18441,N_19369);
or U20236 (N_20236,N_18263,N_18664);
or U20237 (N_20237,N_18842,N_18015);
nor U20238 (N_20238,N_19419,N_18490);
nor U20239 (N_20239,N_19074,N_18615);
or U20240 (N_20240,N_19444,N_18415);
or U20241 (N_20241,N_18677,N_18281);
nor U20242 (N_20242,N_18393,N_18286);
or U20243 (N_20243,N_18737,N_18437);
or U20244 (N_20244,N_19459,N_18369);
or U20245 (N_20245,N_18704,N_18832);
or U20246 (N_20246,N_19456,N_19414);
nand U20247 (N_20247,N_19211,N_18092);
nand U20248 (N_20248,N_19267,N_19268);
and U20249 (N_20249,N_18276,N_19062);
and U20250 (N_20250,N_18414,N_19051);
xor U20251 (N_20251,N_18003,N_18879);
and U20252 (N_20252,N_18839,N_18102);
xor U20253 (N_20253,N_18757,N_18358);
xnor U20254 (N_20254,N_18357,N_18746);
nor U20255 (N_20255,N_19096,N_19301);
or U20256 (N_20256,N_18357,N_19179);
nor U20257 (N_20257,N_18202,N_19173);
xor U20258 (N_20258,N_19042,N_18598);
xnor U20259 (N_20259,N_18798,N_19079);
xor U20260 (N_20260,N_18824,N_19363);
and U20261 (N_20261,N_19122,N_18788);
nand U20262 (N_20262,N_18767,N_18015);
nand U20263 (N_20263,N_18322,N_19105);
nor U20264 (N_20264,N_18921,N_18989);
nand U20265 (N_20265,N_18114,N_18855);
nand U20266 (N_20266,N_18801,N_18991);
nand U20267 (N_20267,N_19220,N_19279);
or U20268 (N_20268,N_18053,N_19450);
and U20269 (N_20269,N_18399,N_18403);
and U20270 (N_20270,N_18996,N_19131);
nor U20271 (N_20271,N_18904,N_18364);
nor U20272 (N_20272,N_18953,N_19157);
nor U20273 (N_20273,N_18340,N_18558);
nand U20274 (N_20274,N_18360,N_19035);
nand U20275 (N_20275,N_18620,N_18909);
or U20276 (N_20276,N_18528,N_19381);
nand U20277 (N_20277,N_19143,N_18754);
nand U20278 (N_20278,N_19032,N_18025);
nand U20279 (N_20279,N_18465,N_18582);
xor U20280 (N_20280,N_19238,N_18168);
nand U20281 (N_20281,N_18719,N_18473);
and U20282 (N_20282,N_18900,N_18865);
and U20283 (N_20283,N_18572,N_18589);
or U20284 (N_20284,N_19229,N_18211);
and U20285 (N_20285,N_18797,N_18579);
nand U20286 (N_20286,N_18825,N_18054);
xnor U20287 (N_20287,N_18293,N_19445);
nor U20288 (N_20288,N_18061,N_18503);
and U20289 (N_20289,N_18664,N_19327);
xor U20290 (N_20290,N_18542,N_18928);
nand U20291 (N_20291,N_19051,N_18346);
or U20292 (N_20292,N_18483,N_18640);
nand U20293 (N_20293,N_18184,N_18017);
nor U20294 (N_20294,N_18601,N_18954);
or U20295 (N_20295,N_18341,N_18483);
xnor U20296 (N_20296,N_18780,N_18632);
nand U20297 (N_20297,N_18766,N_18004);
xnor U20298 (N_20298,N_18059,N_19235);
nor U20299 (N_20299,N_18652,N_19058);
nor U20300 (N_20300,N_19219,N_18944);
xnor U20301 (N_20301,N_18564,N_18088);
nor U20302 (N_20302,N_18174,N_18527);
xor U20303 (N_20303,N_18516,N_18913);
and U20304 (N_20304,N_19344,N_18781);
nor U20305 (N_20305,N_19489,N_19240);
nand U20306 (N_20306,N_19153,N_18805);
and U20307 (N_20307,N_18167,N_19151);
nor U20308 (N_20308,N_18891,N_19480);
nand U20309 (N_20309,N_19395,N_19112);
and U20310 (N_20310,N_19144,N_18338);
nor U20311 (N_20311,N_18251,N_19031);
and U20312 (N_20312,N_19163,N_18821);
and U20313 (N_20313,N_18036,N_18264);
and U20314 (N_20314,N_18810,N_19025);
xnor U20315 (N_20315,N_18424,N_18883);
or U20316 (N_20316,N_19188,N_18645);
nand U20317 (N_20317,N_18249,N_19147);
nand U20318 (N_20318,N_19170,N_19223);
nand U20319 (N_20319,N_18905,N_18891);
xnor U20320 (N_20320,N_18147,N_19359);
nand U20321 (N_20321,N_18429,N_18890);
nand U20322 (N_20322,N_19218,N_18713);
xor U20323 (N_20323,N_19111,N_19364);
nand U20324 (N_20324,N_18091,N_19265);
and U20325 (N_20325,N_19254,N_18895);
xor U20326 (N_20326,N_18482,N_18539);
nand U20327 (N_20327,N_18439,N_18310);
nand U20328 (N_20328,N_19182,N_18909);
nor U20329 (N_20329,N_19041,N_19176);
or U20330 (N_20330,N_18219,N_18941);
and U20331 (N_20331,N_18363,N_18417);
xnor U20332 (N_20332,N_19487,N_18371);
nand U20333 (N_20333,N_18161,N_18874);
xor U20334 (N_20334,N_18408,N_19323);
or U20335 (N_20335,N_19195,N_18069);
and U20336 (N_20336,N_18693,N_19255);
nor U20337 (N_20337,N_18718,N_18585);
and U20338 (N_20338,N_19136,N_18103);
or U20339 (N_20339,N_18377,N_19230);
xor U20340 (N_20340,N_19275,N_19438);
xnor U20341 (N_20341,N_18886,N_18371);
nand U20342 (N_20342,N_18501,N_18944);
nor U20343 (N_20343,N_18629,N_18754);
or U20344 (N_20344,N_19470,N_18841);
and U20345 (N_20345,N_19345,N_18890);
nand U20346 (N_20346,N_18807,N_18092);
or U20347 (N_20347,N_19453,N_18818);
nand U20348 (N_20348,N_18707,N_19291);
nor U20349 (N_20349,N_18911,N_18293);
xnor U20350 (N_20350,N_18351,N_19276);
nor U20351 (N_20351,N_18892,N_18800);
and U20352 (N_20352,N_18646,N_19368);
xor U20353 (N_20353,N_18829,N_18580);
nor U20354 (N_20354,N_18949,N_19433);
nand U20355 (N_20355,N_19250,N_18829);
nand U20356 (N_20356,N_18995,N_18096);
nor U20357 (N_20357,N_18364,N_18073);
or U20358 (N_20358,N_18330,N_19027);
or U20359 (N_20359,N_18169,N_18438);
or U20360 (N_20360,N_18048,N_18795);
or U20361 (N_20361,N_18608,N_19141);
nor U20362 (N_20362,N_18229,N_19488);
nand U20363 (N_20363,N_19299,N_18497);
nand U20364 (N_20364,N_18429,N_19473);
nand U20365 (N_20365,N_18855,N_18911);
nand U20366 (N_20366,N_18732,N_18857);
xor U20367 (N_20367,N_19262,N_19005);
xnor U20368 (N_20368,N_18725,N_19449);
xor U20369 (N_20369,N_18374,N_19450);
nor U20370 (N_20370,N_18247,N_18609);
nand U20371 (N_20371,N_18762,N_18429);
nand U20372 (N_20372,N_18333,N_18442);
and U20373 (N_20373,N_19407,N_18694);
or U20374 (N_20374,N_19234,N_18489);
nand U20375 (N_20375,N_18852,N_18810);
xor U20376 (N_20376,N_18116,N_19020);
nand U20377 (N_20377,N_19245,N_18539);
and U20378 (N_20378,N_18101,N_18737);
nand U20379 (N_20379,N_18162,N_18726);
nor U20380 (N_20380,N_18278,N_18721);
nand U20381 (N_20381,N_18069,N_18372);
nand U20382 (N_20382,N_18370,N_19087);
nand U20383 (N_20383,N_19264,N_18258);
xor U20384 (N_20384,N_19258,N_19454);
nand U20385 (N_20385,N_18293,N_19091);
and U20386 (N_20386,N_18003,N_18570);
nor U20387 (N_20387,N_19346,N_18524);
xor U20388 (N_20388,N_19245,N_18905);
or U20389 (N_20389,N_18607,N_18842);
nand U20390 (N_20390,N_18101,N_19027);
nor U20391 (N_20391,N_18466,N_19280);
nor U20392 (N_20392,N_18370,N_18983);
and U20393 (N_20393,N_19382,N_19074);
nor U20394 (N_20394,N_18042,N_18265);
and U20395 (N_20395,N_18120,N_18366);
nor U20396 (N_20396,N_18938,N_18323);
and U20397 (N_20397,N_18217,N_18185);
or U20398 (N_20398,N_19270,N_18292);
or U20399 (N_20399,N_18326,N_18968);
or U20400 (N_20400,N_18996,N_18942);
or U20401 (N_20401,N_18691,N_19302);
and U20402 (N_20402,N_19442,N_18291);
xor U20403 (N_20403,N_18506,N_18922);
nor U20404 (N_20404,N_18539,N_18507);
xnor U20405 (N_20405,N_18327,N_18397);
and U20406 (N_20406,N_19062,N_19464);
xnor U20407 (N_20407,N_19341,N_18077);
xnor U20408 (N_20408,N_18816,N_19019);
or U20409 (N_20409,N_19292,N_18991);
or U20410 (N_20410,N_18521,N_18972);
nand U20411 (N_20411,N_18348,N_18835);
xnor U20412 (N_20412,N_19117,N_18010);
nor U20413 (N_20413,N_19022,N_19162);
or U20414 (N_20414,N_18286,N_18041);
and U20415 (N_20415,N_18409,N_18303);
nand U20416 (N_20416,N_18286,N_19218);
or U20417 (N_20417,N_18745,N_18097);
xnor U20418 (N_20418,N_18339,N_19432);
xor U20419 (N_20419,N_18089,N_19221);
xnor U20420 (N_20420,N_19165,N_18523);
xnor U20421 (N_20421,N_19002,N_18768);
or U20422 (N_20422,N_19316,N_18958);
nand U20423 (N_20423,N_18920,N_19239);
or U20424 (N_20424,N_18614,N_18426);
or U20425 (N_20425,N_18736,N_18399);
xor U20426 (N_20426,N_18804,N_18125);
and U20427 (N_20427,N_19399,N_18093);
xnor U20428 (N_20428,N_18421,N_19135);
nor U20429 (N_20429,N_18815,N_18230);
nor U20430 (N_20430,N_19445,N_18888);
and U20431 (N_20431,N_18755,N_19153);
xnor U20432 (N_20432,N_18018,N_18064);
xnor U20433 (N_20433,N_18913,N_18479);
and U20434 (N_20434,N_19302,N_18447);
xor U20435 (N_20435,N_18717,N_18325);
or U20436 (N_20436,N_18743,N_19274);
or U20437 (N_20437,N_19183,N_18360);
or U20438 (N_20438,N_18672,N_19117);
nor U20439 (N_20439,N_18324,N_18451);
nand U20440 (N_20440,N_19220,N_18861);
xor U20441 (N_20441,N_19084,N_18980);
and U20442 (N_20442,N_19250,N_18156);
xnor U20443 (N_20443,N_18277,N_18932);
xnor U20444 (N_20444,N_18825,N_18226);
nand U20445 (N_20445,N_19373,N_18428);
nor U20446 (N_20446,N_18659,N_18418);
nor U20447 (N_20447,N_18798,N_18712);
and U20448 (N_20448,N_18183,N_18167);
nor U20449 (N_20449,N_18880,N_19190);
xnor U20450 (N_20450,N_19441,N_18389);
and U20451 (N_20451,N_18873,N_19215);
xor U20452 (N_20452,N_18723,N_18618);
and U20453 (N_20453,N_19270,N_18671);
or U20454 (N_20454,N_19035,N_18558);
or U20455 (N_20455,N_18871,N_18274);
and U20456 (N_20456,N_18162,N_19111);
xnor U20457 (N_20457,N_19105,N_18172);
and U20458 (N_20458,N_18652,N_18456);
xor U20459 (N_20459,N_18652,N_18256);
or U20460 (N_20460,N_18193,N_19389);
nand U20461 (N_20461,N_18804,N_19309);
and U20462 (N_20462,N_18681,N_18007);
nor U20463 (N_20463,N_18327,N_19163);
nand U20464 (N_20464,N_18010,N_19376);
and U20465 (N_20465,N_18702,N_19247);
xor U20466 (N_20466,N_19314,N_18983);
or U20467 (N_20467,N_18491,N_18965);
nor U20468 (N_20468,N_18333,N_18311);
nand U20469 (N_20469,N_18332,N_19483);
xnor U20470 (N_20470,N_18953,N_18559);
xnor U20471 (N_20471,N_18471,N_18798);
nor U20472 (N_20472,N_18649,N_19018);
and U20473 (N_20473,N_19023,N_19380);
nor U20474 (N_20474,N_18458,N_18400);
nand U20475 (N_20475,N_19451,N_19457);
xor U20476 (N_20476,N_18965,N_18357);
xor U20477 (N_20477,N_19388,N_18833);
nand U20478 (N_20478,N_18298,N_19037);
nor U20479 (N_20479,N_18620,N_18391);
xnor U20480 (N_20480,N_18296,N_18450);
nor U20481 (N_20481,N_18683,N_19454);
nand U20482 (N_20482,N_18571,N_19448);
or U20483 (N_20483,N_19274,N_18552);
or U20484 (N_20484,N_18800,N_18900);
nor U20485 (N_20485,N_18825,N_19052);
nand U20486 (N_20486,N_18478,N_19486);
nor U20487 (N_20487,N_18740,N_19335);
or U20488 (N_20488,N_19244,N_19295);
and U20489 (N_20489,N_19180,N_18748);
xnor U20490 (N_20490,N_18476,N_19319);
or U20491 (N_20491,N_19318,N_19188);
or U20492 (N_20492,N_18815,N_18160);
nor U20493 (N_20493,N_19375,N_18858);
or U20494 (N_20494,N_19286,N_19313);
xnor U20495 (N_20495,N_18663,N_18375);
or U20496 (N_20496,N_18518,N_19257);
nor U20497 (N_20497,N_19135,N_19495);
xor U20498 (N_20498,N_19134,N_18931);
xnor U20499 (N_20499,N_19155,N_18696);
xnor U20500 (N_20500,N_18875,N_18290);
nand U20501 (N_20501,N_18809,N_18395);
xnor U20502 (N_20502,N_19143,N_18289);
xor U20503 (N_20503,N_19162,N_18073);
or U20504 (N_20504,N_19358,N_18185);
xor U20505 (N_20505,N_18350,N_18590);
or U20506 (N_20506,N_18554,N_18971);
nand U20507 (N_20507,N_19406,N_18243);
and U20508 (N_20508,N_18496,N_18866);
xnor U20509 (N_20509,N_18419,N_19190);
nand U20510 (N_20510,N_19023,N_18894);
nand U20511 (N_20511,N_18386,N_19326);
nand U20512 (N_20512,N_19067,N_18994);
xor U20513 (N_20513,N_19034,N_18648);
nand U20514 (N_20514,N_18726,N_18465);
and U20515 (N_20515,N_19009,N_18172);
nand U20516 (N_20516,N_18963,N_18026);
xnor U20517 (N_20517,N_19136,N_18101);
xor U20518 (N_20518,N_18203,N_18762);
nor U20519 (N_20519,N_18361,N_18458);
nand U20520 (N_20520,N_19324,N_18752);
nand U20521 (N_20521,N_18543,N_18390);
and U20522 (N_20522,N_18899,N_19428);
nand U20523 (N_20523,N_18621,N_18695);
nor U20524 (N_20524,N_18269,N_18835);
and U20525 (N_20525,N_18745,N_18597);
or U20526 (N_20526,N_19461,N_18297);
xnor U20527 (N_20527,N_19276,N_19074);
and U20528 (N_20528,N_18006,N_18134);
and U20529 (N_20529,N_18818,N_18690);
nor U20530 (N_20530,N_18913,N_18463);
xnor U20531 (N_20531,N_18511,N_18232);
nor U20532 (N_20532,N_18786,N_18170);
and U20533 (N_20533,N_18199,N_19317);
or U20534 (N_20534,N_18809,N_18806);
xor U20535 (N_20535,N_18148,N_18869);
nor U20536 (N_20536,N_18207,N_18635);
nor U20537 (N_20537,N_18778,N_18963);
and U20538 (N_20538,N_18138,N_18679);
and U20539 (N_20539,N_18139,N_19124);
nand U20540 (N_20540,N_19400,N_18901);
nand U20541 (N_20541,N_18266,N_18946);
and U20542 (N_20542,N_18930,N_18660);
nand U20543 (N_20543,N_18602,N_19375);
nor U20544 (N_20544,N_18395,N_18808);
nor U20545 (N_20545,N_18503,N_19099);
and U20546 (N_20546,N_19162,N_18768);
xnor U20547 (N_20547,N_19287,N_18704);
nor U20548 (N_20548,N_19446,N_18656);
and U20549 (N_20549,N_18890,N_18374);
nor U20550 (N_20550,N_18733,N_18121);
nand U20551 (N_20551,N_18496,N_18730);
and U20552 (N_20552,N_19247,N_18586);
and U20553 (N_20553,N_19127,N_18547);
and U20554 (N_20554,N_18897,N_18503);
nand U20555 (N_20555,N_18382,N_19079);
and U20556 (N_20556,N_19083,N_18295);
xnor U20557 (N_20557,N_19457,N_18855);
xnor U20558 (N_20558,N_19271,N_18981);
nand U20559 (N_20559,N_18902,N_18259);
xnor U20560 (N_20560,N_18052,N_19386);
or U20561 (N_20561,N_19019,N_18335);
nand U20562 (N_20562,N_19208,N_18944);
xnor U20563 (N_20563,N_18792,N_18153);
and U20564 (N_20564,N_18036,N_18216);
nor U20565 (N_20565,N_19302,N_18096);
or U20566 (N_20566,N_18886,N_18611);
xnor U20567 (N_20567,N_18389,N_18139);
and U20568 (N_20568,N_19409,N_18596);
and U20569 (N_20569,N_18747,N_19414);
or U20570 (N_20570,N_18708,N_18825);
xnor U20571 (N_20571,N_18717,N_18131);
nor U20572 (N_20572,N_18401,N_18930);
nor U20573 (N_20573,N_19145,N_18617);
xnor U20574 (N_20574,N_18208,N_18402);
nor U20575 (N_20575,N_18417,N_18454);
xor U20576 (N_20576,N_19279,N_18413);
xor U20577 (N_20577,N_18199,N_19055);
or U20578 (N_20578,N_18141,N_18617);
xor U20579 (N_20579,N_18532,N_18869);
or U20580 (N_20580,N_18769,N_18243);
nand U20581 (N_20581,N_18780,N_18851);
xor U20582 (N_20582,N_19337,N_18224);
and U20583 (N_20583,N_18204,N_18453);
and U20584 (N_20584,N_18144,N_18338);
nand U20585 (N_20585,N_18704,N_18921);
or U20586 (N_20586,N_18497,N_18820);
or U20587 (N_20587,N_18480,N_18232);
and U20588 (N_20588,N_18599,N_18889);
nand U20589 (N_20589,N_18211,N_18476);
nor U20590 (N_20590,N_18794,N_18379);
nand U20591 (N_20591,N_18184,N_18457);
xor U20592 (N_20592,N_18830,N_18646);
nand U20593 (N_20593,N_19221,N_18141);
nor U20594 (N_20594,N_18687,N_18349);
or U20595 (N_20595,N_18738,N_18486);
nand U20596 (N_20596,N_19482,N_18208);
or U20597 (N_20597,N_18907,N_18071);
nor U20598 (N_20598,N_19209,N_18397);
and U20599 (N_20599,N_18820,N_18136);
nand U20600 (N_20600,N_18811,N_18830);
xnor U20601 (N_20601,N_18129,N_19404);
xor U20602 (N_20602,N_18578,N_19128);
nor U20603 (N_20603,N_19197,N_18444);
and U20604 (N_20604,N_18350,N_18746);
nand U20605 (N_20605,N_18700,N_18049);
and U20606 (N_20606,N_18058,N_18906);
and U20607 (N_20607,N_18519,N_18699);
xnor U20608 (N_20608,N_19221,N_18584);
xor U20609 (N_20609,N_18721,N_19140);
nor U20610 (N_20610,N_18192,N_18462);
or U20611 (N_20611,N_18803,N_19461);
xor U20612 (N_20612,N_19087,N_18282);
nor U20613 (N_20613,N_19233,N_18652);
or U20614 (N_20614,N_18555,N_19328);
nor U20615 (N_20615,N_18733,N_18876);
nand U20616 (N_20616,N_18746,N_19341);
nand U20617 (N_20617,N_18635,N_18918);
xor U20618 (N_20618,N_19092,N_19498);
nor U20619 (N_20619,N_19058,N_18799);
and U20620 (N_20620,N_19157,N_18293);
xnor U20621 (N_20621,N_18059,N_19048);
nand U20622 (N_20622,N_18483,N_18594);
xnor U20623 (N_20623,N_19049,N_18939);
and U20624 (N_20624,N_19293,N_18525);
nor U20625 (N_20625,N_18522,N_18886);
or U20626 (N_20626,N_19337,N_18983);
and U20627 (N_20627,N_19269,N_18674);
xnor U20628 (N_20628,N_18677,N_18119);
nor U20629 (N_20629,N_19246,N_19176);
and U20630 (N_20630,N_18872,N_19296);
or U20631 (N_20631,N_18726,N_18190);
nand U20632 (N_20632,N_18391,N_19111);
nor U20633 (N_20633,N_19207,N_18845);
or U20634 (N_20634,N_18620,N_18002);
xor U20635 (N_20635,N_18081,N_18375);
and U20636 (N_20636,N_18060,N_18460);
xor U20637 (N_20637,N_18649,N_18847);
xnor U20638 (N_20638,N_18276,N_18385);
and U20639 (N_20639,N_19489,N_18940);
nor U20640 (N_20640,N_18152,N_18633);
or U20641 (N_20641,N_18112,N_18231);
nand U20642 (N_20642,N_19009,N_18408);
or U20643 (N_20643,N_18265,N_18546);
nand U20644 (N_20644,N_18500,N_18210);
or U20645 (N_20645,N_18330,N_18043);
or U20646 (N_20646,N_18293,N_19348);
xnor U20647 (N_20647,N_18658,N_18364);
and U20648 (N_20648,N_18943,N_18200);
nor U20649 (N_20649,N_18345,N_18170);
or U20650 (N_20650,N_19176,N_18919);
and U20651 (N_20651,N_19393,N_18835);
nand U20652 (N_20652,N_18055,N_18799);
or U20653 (N_20653,N_18197,N_18337);
xnor U20654 (N_20654,N_18349,N_19098);
nand U20655 (N_20655,N_18594,N_19374);
nor U20656 (N_20656,N_18200,N_18140);
nand U20657 (N_20657,N_19316,N_18914);
xnor U20658 (N_20658,N_18765,N_18321);
nor U20659 (N_20659,N_18433,N_19087);
and U20660 (N_20660,N_18543,N_19290);
nor U20661 (N_20661,N_18737,N_18852);
nand U20662 (N_20662,N_19118,N_18970);
and U20663 (N_20663,N_19325,N_18659);
and U20664 (N_20664,N_19233,N_19178);
nor U20665 (N_20665,N_18494,N_18567);
nand U20666 (N_20666,N_18445,N_19260);
xnor U20667 (N_20667,N_19295,N_19109);
xnor U20668 (N_20668,N_18246,N_18732);
nor U20669 (N_20669,N_19182,N_18440);
nor U20670 (N_20670,N_18147,N_19091);
nand U20671 (N_20671,N_18172,N_18725);
and U20672 (N_20672,N_19338,N_18311);
nand U20673 (N_20673,N_18164,N_19300);
and U20674 (N_20674,N_18456,N_18144);
nand U20675 (N_20675,N_19379,N_19197);
xor U20676 (N_20676,N_18163,N_19000);
nor U20677 (N_20677,N_19320,N_18851);
and U20678 (N_20678,N_18920,N_18592);
or U20679 (N_20679,N_19310,N_19200);
nand U20680 (N_20680,N_18521,N_18903);
nand U20681 (N_20681,N_18124,N_18469);
or U20682 (N_20682,N_18337,N_18558);
or U20683 (N_20683,N_18058,N_19287);
nor U20684 (N_20684,N_19474,N_18996);
or U20685 (N_20685,N_18952,N_18826);
and U20686 (N_20686,N_18274,N_19003);
nor U20687 (N_20687,N_18286,N_19213);
and U20688 (N_20688,N_19278,N_19127);
nor U20689 (N_20689,N_18686,N_18474);
nand U20690 (N_20690,N_18780,N_19287);
and U20691 (N_20691,N_18215,N_18210);
or U20692 (N_20692,N_19120,N_18155);
nand U20693 (N_20693,N_18088,N_18471);
or U20694 (N_20694,N_19353,N_19032);
xor U20695 (N_20695,N_19430,N_19209);
or U20696 (N_20696,N_18157,N_18577);
nand U20697 (N_20697,N_18512,N_19154);
xnor U20698 (N_20698,N_19259,N_18686);
and U20699 (N_20699,N_18378,N_18648);
nand U20700 (N_20700,N_18471,N_19254);
and U20701 (N_20701,N_18538,N_19486);
nor U20702 (N_20702,N_19036,N_19001);
and U20703 (N_20703,N_18740,N_19069);
nand U20704 (N_20704,N_18281,N_18065);
nor U20705 (N_20705,N_18721,N_19083);
nand U20706 (N_20706,N_19299,N_19355);
or U20707 (N_20707,N_18321,N_19244);
and U20708 (N_20708,N_18503,N_18935);
nor U20709 (N_20709,N_19069,N_19231);
nor U20710 (N_20710,N_19168,N_18665);
nor U20711 (N_20711,N_19497,N_18640);
nand U20712 (N_20712,N_18344,N_19131);
or U20713 (N_20713,N_18244,N_19060);
or U20714 (N_20714,N_18501,N_19278);
or U20715 (N_20715,N_18377,N_19209);
nor U20716 (N_20716,N_19005,N_18576);
and U20717 (N_20717,N_19257,N_19162);
nand U20718 (N_20718,N_19051,N_18174);
or U20719 (N_20719,N_18225,N_18498);
nand U20720 (N_20720,N_18022,N_18992);
nand U20721 (N_20721,N_18324,N_18131);
nand U20722 (N_20722,N_18770,N_19375);
nand U20723 (N_20723,N_19424,N_19025);
nand U20724 (N_20724,N_18463,N_19413);
and U20725 (N_20725,N_18643,N_18727);
nor U20726 (N_20726,N_18073,N_18215);
xor U20727 (N_20727,N_18448,N_18727);
or U20728 (N_20728,N_19322,N_18710);
nand U20729 (N_20729,N_19351,N_19048);
or U20730 (N_20730,N_18743,N_19045);
xor U20731 (N_20731,N_18360,N_19469);
or U20732 (N_20732,N_18530,N_19052);
and U20733 (N_20733,N_18802,N_19423);
nor U20734 (N_20734,N_18940,N_18303);
nor U20735 (N_20735,N_19493,N_18024);
nand U20736 (N_20736,N_18295,N_18074);
nor U20737 (N_20737,N_18385,N_18892);
or U20738 (N_20738,N_18364,N_18947);
xor U20739 (N_20739,N_18460,N_19484);
nand U20740 (N_20740,N_18008,N_19067);
or U20741 (N_20741,N_18914,N_18287);
nand U20742 (N_20742,N_18136,N_18404);
nand U20743 (N_20743,N_18366,N_18117);
nor U20744 (N_20744,N_18344,N_18000);
or U20745 (N_20745,N_19065,N_18804);
nor U20746 (N_20746,N_18023,N_18225);
and U20747 (N_20747,N_18419,N_18936);
and U20748 (N_20748,N_19078,N_18165);
and U20749 (N_20749,N_18187,N_18349);
and U20750 (N_20750,N_19417,N_19459);
nand U20751 (N_20751,N_18820,N_18964);
or U20752 (N_20752,N_18970,N_18475);
and U20753 (N_20753,N_19343,N_18658);
and U20754 (N_20754,N_18615,N_18443);
nor U20755 (N_20755,N_18553,N_18789);
xor U20756 (N_20756,N_19411,N_19271);
nor U20757 (N_20757,N_19453,N_19307);
and U20758 (N_20758,N_18735,N_18932);
xnor U20759 (N_20759,N_18332,N_18637);
nand U20760 (N_20760,N_18116,N_19152);
xor U20761 (N_20761,N_18516,N_18520);
nand U20762 (N_20762,N_18976,N_19232);
nor U20763 (N_20763,N_19207,N_19089);
xnor U20764 (N_20764,N_18523,N_18326);
nor U20765 (N_20765,N_19111,N_19251);
xor U20766 (N_20766,N_18472,N_19152);
and U20767 (N_20767,N_18903,N_18787);
xor U20768 (N_20768,N_18281,N_18917);
or U20769 (N_20769,N_18781,N_19413);
nand U20770 (N_20770,N_18148,N_18122);
nand U20771 (N_20771,N_18319,N_19381);
nand U20772 (N_20772,N_18823,N_18429);
nor U20773 (N_20773,N_18440,N_18111);
or U20774 (N_20774,N_19321,N_19428);
or U20775 (N_20775,N_18618,N_18041);
nand U20776 (N_20776,N_18263,N_18896);
nand U20777 (N_20777,N_18454,N_18876);
and U20778 (N_20778,N_18365,N_18303);
or U20779 (N_20779,N_18033,N_18438);
and U20780 (N_20780,N_18588,N_18511);
nand U20781 (N_20781,N_18650,N_18217);
and U20782 (N_20782,N_18291,N_18244);
nor U20783 (N_20783,N_19178,N_18715);
or U20784 (N_20784,N_19057,N_19076);
or U20785 (N_20785,N_18558,N_18185);
and U20786 (N_20786,N_18784,N_18875);
nor U20787 (N_20787,N_19035,N_18653);
and U20788 (N_20788,N_19268,N_18527);
xnor U20789 (N_20789,N_18966,N_19364);
xnor U20790 (N_20790,N_18609,N_18426);
and U20791 (N_20791,N_18993,N_19419);
and U20792 (N_20792,N_18792,N_19477);
or U20793 (N_20793,N_18801,N_19200);
nor U20794 (N_20794,N_18506,N_19243);
xor U20795 (N_20795,N_18897,N_18562);
nor U20796 (N_20796,N_19402,N_18345);
and U20797 (N_20797,N_19064,N_18486);
nor U20798 (N_20798,N_18568,N_19033);
and U20799 (N_20799,N_18108,N_19264);
nand U20800 (N_20800,N_18301,N_19123);
nor U20801 (N_20801,N_18957,N_19083);
xor U20802 (N_20802,N_18420,N_18869);
and U20803 (N_20803,N_19309,N_18665);
nand U20804 (N_20804,N_18109,N_19040);
nor U20805 (N_20805,N_18926,N_18642);
and U20806 (N_20806,N_18245,N_19161);
xnor U20807 (N_20807,N_18530,N_18512);
xor U20808 (N_20808,N_19417,N_19292);
xnor U20809 (N_20809,N_19460,N_18409);
nand U20810 (N_20810,N_19366,N_18197);
nand U20811 (N_20811,N_19054,N_18520);
xnor U20812 (N_20812,N_18182,N_19346);
nand U20813 (N_20813,N_18032,N_18399);
nor U20814 (N_20814,N_19178,N_18653);
xor U20815 (N_20815,N_19039,N_18412);
nor U20816 (N_20816,N_18813,N_19309);
and U20817 (N_20817,N_19273,N_18753);
nand U20818 (N_20818,N_19265,N_19145);
nor U20819 (N_20819,N_18604,N_19101);
nand U20820 (N_20820,N_18366,N_18565);
nand U20821 (N_20821,N_19225,N_18907);
and U20822 (N_20822,N_18653,N_18804);
nand U20823 (N_20823,N_19219,N_18564);
xnor U20824 (N_20824,N_18679,N_18469);
nor U20825 (N_20825,N_18609,N_19030);
or U20826 (N_20826,N_19376,N_19135);
and U20827 (N_20827,N_18477,N_19423);
or U20828 (N_20828,N_18495,N_18311);
or U20829 (N_20829,N_18447,N_19179);
nor U20830 (N_20830,N_18271,N_18566);
or U20831 (N_20831,N_18131,N_19088);
and U20832 (N_20832,N_18460,N_18170);
nor U20833 (N_20833,N_18779,N_19217);
and U20834 (N_20834,N_18329,N_18656);
and U20835 (N_20835,N_18055,N_19113);
xor U20836 (N_20836,N_19332,N_18886);
nor U20837 (N_20837,N_18838,N_18583);
or U20838 (N_20838,N_18433,N_18330);
or U20839 (N_20839,N_18246,N_18747);
nor U20840 (N_20840,N_19490,N_18611);
nand U20841 (N_20841,N_18732,N_18597);
nor U20842 (N_20842,N_18845,N_18859);
nand U20843 (N_20843,N_18414,N_18007);
or U20844 (N_20844,N_19036,N_19032);
and U20845 (N_20845,N_18644,N_19041);
nor U20846 (N_20846,N_19118,N_18344);
nor U20847 (N_20847,N_18348,N_18012);
or U20848 (N_20848,N_19180,N_18383);
nand U20849 (N_20849,N_18848,N_18213);
and U20850 (N_20850,N_18475,N_18835);
xor U20851 (N_20851,N_19175,N_19361);
and U20852 (N_20852,N_19455,N_18384);
or U20853 (N_20853,N_18747,N_19060);
and U20854 (N_20854,N_19316,N_18916);
and U20855 (N_20855,N_18445,N_18983);
nor U20856 (N_20856,N_18401,N_18592);
and U20857 (N_20857,N_18921,N_18938);
or U20858 (N_20858,N_18632,N_19439);
nor U20859 (N_20859,N_18392,N_18318);
nand U20860 (N_20860,N_19380,N_19029);
and U20861 (N_20861,N_18646,N_18248);
xnor U20862 (N_20862,N_18150,N_18338);
or U20863 (N_20863,N_18672,N_18169);
and U20864 (N_20864,N_18398,N_18606);
and U20865 (N_20865,N_19005,N_19469);
xnor U20866 (N_20866,N_19085,N_18754);
nand U20867 (N_20867,N_19078,N_18184);
and U20868 (N_20868,N_18324,N_19482);
or U20869 (N_20869,N_18122,N_19295);
nand U20870 (N_20870,N_18655,N_18720);
nor U20871 (N_20871,N_18418,N_19078);
xor U20872 (N_20872,N_18086,N_18199);
and U20873 (N_20873,N_18329,N_19059);
and U20874 (N_20874,N_19233,N_18391);
nand U20875 (N_20875,N_18975,N_19425);
and U20876 (N_20876,N_18324,N_18763);
nor U20877 (N_20877,N_19305,N_19255);
xnor U20878 (N_20878,N_18646,N_18534);
nand U20879 (N_20879,N_19028,N_18381);
or U20880 (N_20880,N_18717,N_19387);
nand U20881 (N_20881,N_18259,N_19279);
xnor U20882 (N_20882,N_19112,N_18190);
xnor U20883 (N_20883,N_18910,N_18387);
or U20884 (N_20884,N_19487,N_19469);
nor U20885 (N_20885,N_19413,N_19299);
nor U20886 (N_20886,N_19349,N_19040);
nor U20887 (N_20887,N_19260,N_19175);
and U20888 (N_20888,N_18945,N_18046);
nand U20889 (N_20889,N_19179,N_18195);
nor U20890 (N_20890,N_19120,N_18171);
nor U20891 (N_20891,N_18259,N_18939);
or U20892 (N_20892,N_19115,N_19407);
and U20893 (N_20893,N_18919,N_18737);
and U20894 (N_20894,N_18433,N_18561);
and U20895 (N_20895,N_19322,N_18010);
nand U20896 (N_20896,N_18694,N_18810);
or U20897 (N_20897,N_18089,N_18816);
xor U20898 (N_20898,N_19383,N_19125);
or U20899 (N_20899,N_18802,N_19466);
xor U20900 (N_20900,N_18486,N_19336);
nand U20901 (N_20901,N_18804,N_18770);
xor U20902 (N_20902,N_18748,N_19135);
nand U20903 (N_20903,N_18571,N_19137);
nor U20904 (N_20904,N_19281,N_19195);
or U20905 (N_20905,N_18036,N_19025);
or U20906 (N_20906,N_18733,N_18192);
nand U20907 (N_20907,N_18672,N_19009);
nor U20908 (N_20908,N_18899,N_19452);
and U20909 (N_20909,N_18939,N_18609);
nand U20910 (N_20910,N_19453,N_18661);
nor U20911 (N_20911,N_18054,N_18748);
and U20912 (N_20912,N_19397,N_18440);
nand U20913 (N_20913,N_18265,N_19302);
nand U20914 (N_20914,N_19058,N_19227);
and U20915 (N_20915,N_19183,N_18410);
and U20916 (N_20916,N_18768,N_19305);
nand U20917 (N_20917,N_18703,N_19076);
nand U20918 (N_20918,N_19145,N_19070);
or U20919 (N_20919,N_18557,N_18809);
nand U20920 (N_20920,N_18619,N_18937);
nor U20921 (N_20921,N_19452,N_19350);
or U20922 (N_20922,N_18583,N_19209);
or U20923 (N_20923,N_18630,N_18574);
xnor U20924 (N_20924,N_18246,N_18787);
nor U20925 (N_20925,N_18882,N_18372);
xor U20926 (N_20926,N_18574,N_19201);
nor U20927 (N_20927,N_19186,N_18515);
or U20928 (N_20928,N_18045,N_18144);
xnor U20929 (N_20929,N_18874,N_18367);
xnor U20930 (N_20930,N_18278,N_18841);
nand U20931 (N_20931,N_18557,N_19190);
or U20932 (N_20932,N_18655,N_18557);
and U20933 (N_20933,N_18912,N_18528);
or U20934 (N_20934,N_18705,N_18917);
or U20935 (N_20935,N_18545,N_18484);
xor U20936 (N_20936,N_18126,N_19470);
or U20937 (N_20937,N_18401,N_19056);
and U20938 (N_20938,N_19181,N_18870);
or U20939 (N_20939,N_19146,N_18267);
or U20940 (N_20940,N_19085,N_18807);
nand U20941 (N_20941,N_18006,N_18387);
xnor U20942 (N_20942,N_18966,N_19113);
and U20943 (N_20943,N_18912,N_18443);
xor U20944 (N_20944,N_19187,N_19037);
nor U20945 (N_20945,N_19015,N_19278);
xnor U20946 (N_20946,N_18503,N_18838);
and U20947 (N_20947,N_18156,N_19063);
nand U20948 (N_20948,N_19419,N_19160);
nor U20949 (N_20949,N_18340,N_18291);
nand U20950 (N_20950,N_18174,N_18708);
nand U20951 (N_20951,N_19481,N_18120);
and U20952 (N_20952,N_18886,N_19278);
and U20953 (N_20953,N_18152,N_18361);
or U20954 (N_20954,N_19420,N_19356);
and U20955 (N_20955,N_18097,N_19479);
or U20956 (N_20956,N_19491,N_19169);
xnor U20957 (N_20957,N_18598,N_18389);
xor U20958 (N_20958,N_18425,N_18119);
xor U20959 (N_20959,N_18370,N_18526);
xor U20960 (N_20960,N_19289,N_18113);
or U20961 (N_20961,N_19400,N_18051);
or U20962 (N_20962,N_18066,N_19072);
or U20963 (N_20963,N_18132,N_18108);
and U20964 (N_20964,N_19456,N_19165);
or U20965 (N_20965,N_18086,N_18991);
or U20966 (N_20966,N_19221,N_19351);
and U20967 (N_20967,N_18616,N_18886);
nor U20968 (N_20968,N_19256,N_18718);
nand U20969 (N_20969,N_18564,N_18291);
or U20970 (N_20970,N_19118,N_18689);
nor U20971 (N_20971,N_19459,N_18516);
xnor U20972 (N_20972,N_19041,N_18789);
xor U20973 (N_20973,N_18901,N_18590);
nand U20974 (N_20974,N_18282,N_19053);
nand U20975 (N_20975,N_18817,N_18344);
nor U20976 (N_20976,N_18473,N_18387);
nor U20977 (N_20977,N_18406,N_18449);
nand U20978 (N_20978,N_18229,N_18908);
nand U20979 (N_20979,N_18541,N_18088);
nor U20980 (N_20980,N_19455,N_18149);
or U20981 (N_20981,N_18283,N_18032);
nand U20982 (N_20982,N_18419,N_19021);
and U20983 (N_20983,N_19262,N_18644);
nor U20984 (N_20984,N_19148,N_18434);
nand U20985 (N_20985,N_18641,N_18418);
nand U20986 (N_20986,N_18322,N_19052);
nor U20987 (N_20987,N_18539,N_19144);
nand U20988 (N_20988,N_19451,N_19178);
nor U20989 (N_20989,N_18580,N_18804);
xor U20990 (N_20990,N_18348,N_18459);
nand U20991 (N_20991,N_19048,N_18160);
xor U20992 (N_20992,N_18577,N_19265);
xnor U20993 (N_20993,N_18010,N_18042);
nor U20994 (N_20994,N_18267,N_18533);
nor U20995 (N_20995,N_18554,N_18866);
xor U20996 (N_20996,N_18200,N_18994);
xor U20997 (N_20997,N_19067,N_18809);
and U20998 (N_20998,N_19499,N_18641);
and U20999 (N_20999,N_18396,N_18881);
nor U21000 (N_21000,N_20983,N_19849);
xor U21001 (N_21001,N_20044,N_19534);
nor U21002 (N_21002,N_19928,N_19945);
or U21003 (N_21003,N_20318,N_20776);
xor U21004 (N_21004,N_20668,N_20370);
nand U21005 (N_21005,N_20274,N_20502);
nand U21006 (N_21006,N_20030,N_20036);
and U21007 (N_21007,N_20991,N_20489);
and U21008 (N_21008,N_20915,N_19854);
xor U21009 (N_21009,N_19605,N_20353);
and U21010 (N_21010,N_20658,N_20769);
and U21011 (N_21011,N_20172,N_20149);
nand U21012 (N_21012,N_19732,N_20236);
or U21013 (N_21013,N_19598,N_20610);
xor U21014 (N_21014,N_19552,N_19652);
or U21015 (N_21015,N_19774,N_20708);
xor U21016 (N_21016,N_20442,N_20001);
and U21017 (N_21017,N_20517,N_20351);
nand U21018 (N_21018,N_20386,N_20644);
xnor U21019 (N_21019,N_19847,N_20912);
xnor U21020 (N_21020,N_20560,N_19693);
nor U21021 (N_21021,N_19771,N_20949);
and U21022 (N_21022,N_20689,N_20378);
xor U21023 (N_21023,N_20816,N_20080);
or U21024 (N_21024,N_20262,N_20525);
nor U21025 (N_21025,N_20966,N_20215);
or U21026 (N_21026,N_20661,N_20791);
or U21027 (N_21027,N_20071,N_19805);
nor U21028 (N_21028,N_20028,N_20267);
nand U21029 (N_21029,N_19581,N_19957);
or U21030 (N_21030,N_20363,N_20112);
nor U21031 (N_21031,N_20040,N_19950);
and U21032 (N_21032,N_20298,N_20359);
nor U21033 (N_21033,N_19800,N_20847);
nor U21034 (N_21034,N_20210,N_20952);
nand U21035 (N_21035,N_19866,N_20812);
and U21036 (N_21036,N_20056,N_20093);
and U21037 (N_21037,N_20700,N_20259);
nor U21038 (N_21038,N_20367,N_20582);
xor U21039 (N_21039,N_20702,N_20813);
nand U21040 (N_21040,N_19955,N_19707);
or U21041 (N_21041,N_19891,N_20108);
and U21042 (N_21042,N_20483,N_20438);
or U21043 (N_21043,N_20960,N_19685);
and U21044 (N_21044,N_20592,N_20907);
or U21045 (N_21045,N_19617,N_19985);
xnor U21046 (N_21046,N_20023,N_19943);
xnor U21047 (N_21047,N_20929,N_20146);
nor U21048 (N_21048,N_20410,N_20959);
nand U21049 (N_21049,N_20555,N_20862);
or U21050 (N_21050,N_20406,N_19768);
or U21051 (N_21051,N_20356,N_20453);
nand U21052 (N_21052,N_19518,N_19616);
nor U21053 (N_21053,N_19748,N_20335);
nor U21054 (N_21054,N_20137,N_20885);
xor U21055 (N_21055,N_20109,N_19868);
nor U21056 (N_21056,N_19872,N_20435);
and U21057 (N_21057,N_20035,N_20784);
nand U21058 (N_21058,N_19627,N_19628);
nand U21059 (N_21059,N_19841,N_19833);
or U21060 (N_21060,N_19668,N_19753);
nand U21061 (N_21061,N_19728,N_20313);
nor U21062 (N_21062,N_20857,N_20740);
nor U21063 (N_21063,N_20581,N_19861);
nor U21064 (N_21064,N_20482,N_20166);
xor U21065 (N_21065,N_19824,N_19939);
nand U21066 (N_21066,N_20576,N_20797);
or U21067 (N_21067,N_20693,N_20147);
nand U21068 (N_21068,N_20711,N_20434);
xnor U21069 (N_21069,N_20189,N_20234);
and U21070 (N_21070,N_20466,N_20664);
or U21071 (N_21071,N_20452,N_19700);
nand U21072 (N_21072,N_20198,N_20691);
or U21073 (N_21073,N_20051,N_20894);
or U21074 (N_21074,N_19860,N_20395);
nor U21075 (N_21075,N_20543,N_19516);
nand U21076 (N_21076,N_19724,N_20004);
or U21077 (N_21077,N_20856,N_19907);
nor U21078 (N_21078,N_20654,N_20533);
nor U21079 (N_21079,N_19917,N_19525);
nand U21080 (N_21080,N_19618,N_20766);
and U21081 (N_21081,N_19530,N_19610);
nand U21082 (N_21082,N_19900,N_20834);
and U21083 (N_21083,N_19770,N_20311);
or U21084 (N_21084,N_19964,N_20032);
or U21085 (N_21085,N_20323,N_20314);
nor U21086 (N_21086,N_20900,N_20544);
xor U21087 (N_21087,N_20640,N_20387);
nand U21088 (N_21088,N_19689,N_20807);
nor U21089 (N_21089,N_20888,N_20542);
or U21090 (N_21090,N_20628,N_20195);
and U21091 (N_21091,N_19767,N_20104);
nand U21092 (N_21092,N_20814,N_20443);
xor U21093 (N_21093,N_20537,N_20403);
nand U21094 (N_21094,N_20346,N_19650);
nand U21095 (N_21095,N_19733,N_19521);
and U21096 (N_21096,N_19844,N_19745);
xnor U21097 (N_21097,N_20762,N_20496);
nor U21098 (N_21098,N_19877,N_20275);
xor U21099 (N_21099,N_19543,N_20958);
nand U21100 (N_21100,N_20278,N_20853);
or U21101 (N_21101,N_20871,N_20910);
nand U21102 (N_21102,N_20974,N_20160);
xnor U21103 (N_21103,N_20852,N_20755);
nand U21104 (N_21104,N_19704,N_20045);
and U21105 (N_21105,N_19554,N_20296);
nand U21106 (N_21106,N_20184,N_19665);
nor U21107 (N_21107,N_20264,N_19663);
nand U21108 (N_21108,N_20715,N_19880);
or U21109 (N_21109,N_19739,N_20240);
nand U21110 (N_21110,N_20709,N_19672);
or U21111 (N_21111,N_20439,N_19925);
nand U21112 (N_21112,N_19579,N_20993);
nand U21113 (N_21113,N_20696,N_20332);
and U21114 (N_21114,N_20519,N_19561);
xor U21115 (N_21115,N_19835,N_19836);
and U21116 (N_21116,N_20969,N_19750);
xor U21117 (N_21117,N_20380,N_19741);
xor U21118 (N_21118,N_20297,N_20244);
nor U21119 (N_21119,N_19811,N_20424);
xor U21120 (N_21120,N_20926,N_20577);
xor U21121 (N_21121,N_20136,N_20670);
xor U21122 (N_21122,N_20669,N_20065);
or U21123 (N_21123,N_20979,N_20680);
and U21124 (N_21124,N_20339,N_19933);
nor U21125 (N_21125,N_20786,N_19746);
and U21126 (N_21126,N_19954,N_20132);
or U21127 (N_21127,N_19649,N_20985);
xnor U21128 (N_21128,N_20428,N_19946);
xor U21129 (N_21129,N_20081,N_20887);
and U21130 (N_21130,N_20948,N_20790);
xor U21131 (N_21131,N_20638,N_20593);
nor U21132 (N_21132,N_20009,N_19548);
nand U21133 (N_21133,N_20598,N_20672);
xor U21134 (N_21134,N_20495,N_20650);
nor U21135 (N_21135,N_19978,N_20557);
nor U21136 (N_21136,N_20961,N_20315);
xor U21137 (N_21137,N_19619,N_19555);
and U21138 (N_21138,N_20687,N_20990);
nand U21139 (N_21139,N_19821,N_19603);
or U21140 (N_21140,N_20421,N_20761);
xnor U21141 (N_21141,N_20566,N_20682);
and U21142 (N_21142,N_19608,N_20013);
nor U21143 (N_21143,N_20545,N_19677);
or U21144 (N_21144,N_20425,N_19590);
nor U21145 (N_21145,N_20446,N_20733);
or U21146 (N_21146,N_20512,N_20381);
or U21147 (N_21147,N_19743,N_20225);
or U21148 (N_21148,N_20111,N_20678);
xor U21149 (N_21149,N_20142,N_19643);
nor U21150 (N_21150,N_20374,N_20076);
nor U21151 (N_21151,N_20605,N_19684);
or U21152 (N_21152,N_20667,N_20968);
xor U21153 (N_21153,N_20157,N_20735);
xnor U21154 (N_21154,N_20676,N_20526);
or U21155 (N_21155,N_20479,N_20930);
xnor U21156 (N_21156,N_20491,N_20456);
xor U21157 (N_21157,N_19640,N_20584);
and U21158 (N_21158,N_20033,N_20869);
nand U21159 (N_21159,N_20880,N_20747);
xor U21160 (N_21160,N_20083,N_20398);
xor U21161 (N_21161,N_20053,N_20192);
nand U21162 (N_21162,N_19820,N_20940);
or U21163 (N_21163,N_20389,N_19815);
xnor U21164 (N_21164,N_20587,N_19675);
and U21165 (N_21165,N_20103,N_19705);
and U21166 (N_21166,N_20532,N_20651);
xor U21167 (N_21167,N_20568,N_19511);
nor U21168 (N_21168,N_20569,N_20357);
xnor U21169 (N_21169,N_20097,N_20580);
and U21170 (N_21170,N_20271,N_19651);
and U21171 (N_21171,N_20607,N_20333);
xnor U21172 (N_21172,N_20202,N_19965);
and U21173 (N_21173,N_20105,N_19904);
nor U21174 (N_21174,N_19851,N_20704);
or U21175 (N_21175,N_19502,N_20261);
and U21176 (N_21176,N_20072,N_19926);
or U21177 (N_21177,N_19738,N_19698);
nand U21178 (N_21178,N_19512,N_19576);
and U21179 (N_21179,N_20882,N_19930);
xor U21180 (N_21180,N_20062,N_20694);
nand U21181 (N_21181,N_20904,N_19542);
or U21182 (N_21182,N_20655,N_19885);
nor U21183 (N_21183,N_20504,N_19895);
nor U21184 (N_21184,N_20705,N_20352);
nor U21185 (N_21185,N_20385,N_20874);
or U21186 (N_21186,N_20626,N_19823);
or U21187 (N_21187,N_20141,N_20469);
or U21188 (N_21188,N_19522,N_20501);
or U21189 (N_21189,N_19637,N_20127);
nor U21190 (N_21190,N_19974,N_19573);
or U21191 (N_21191,N_20746,N_20742);
and U21192 (N_21192,N_20879,N_19856);
xor U21193 (N_21193,N_20583,N_19865);
nand U21194 (N_21194,N_20795,N_20843);
xor U21195 (N_21195,N_20506,N_20154);
xor U21196 (N_21196,N_19842,N_20113);
xor U21197 (N_21197,N_20850,N_19818);
nand U21198 (N_21198,N_20712,N_19729);
xnor U21199 (N_21199,N_20050,N_20014);
nor U21200 (N_21200,N_19817,N_20269);
and U21201 (N_21201,N_20734,N_19621);
or U21202 (N_21202,N_20227,N_20535);
or U21203 (N_21203,N_20559,N_20409);
nor U21204 (N_21204,N_20486,N_20675);
xnor U21205 (N_21205,N_19929,N_19919);
or U21206 (N_21206,N_20753,N_19714);
and U21207 (N_21207,N_20055,N_19813);
nor U21208 (N_21208,N_20039,N_19690);
or U21209 (N_21209,N_20309,N_19655);
xor U21210 (N_21210,N_19592,N_20804);
or U21211 (N_21211,N_19881,N_20954);
and U21212 (N_21212,N_20806,N_20831);
xnor U21213 (N_21213,N_20052,N_20291);
and U21214 (N_21214,N_19898,N_19992);
nand U21215 (N_21215,N_19725,N_19683);
xor U21216 (N_21216,N_19807,N_20855);
nor U21217 (N_21217,N_20485,N_20413);
or U21218 (N_21218,N_19987,N_20823);
and U21219 (N_21219,N_20552,N_20467);
and U21220 (N_21220,N_19712,N_20006);
nand U21221 (N_21221,N_20858,N_20444);
or U21222 (N_21222,N_20523,N_20273);
or U21223 (N_21223,N_20170,N_19830);
and U21224 (N_21224,N_20738,N_20737);
nor U21225 (N_21225,N_20212,N_19659);
nand U21226 (N_21226,N_20931,N_19814);
nand U21227 (N_21227,N_20892,N_20860);
xnor U21228 (N_21228,N_20963,N_20138);
xnor U21229 (N_21229,N_20017,N_20938);
nor U21230 (N_21230,N_20515,N_20548);
or U21231 (N_21231,N_19503,N_20728);
nor U21232 (N_21232,N_19609,N_20690);
nand U21233 (N_21233,N_20376,N_20503);
nor U21234 (N_21234,N_20220,N_20509);
nand U21235 (N_21235,N_20868,N_19763);
nand U21236 (N_21236,N_20088,N_20956);
xor U21237 (N_21237,N_20665,N_19559);
and U21238 (N_21238,N_20263,N_19870);
nand U21239 (N_21239,N_20546,N_20794);
or U21240 (N_21240,N_20837,N_19638);
xor U21241 (N_21241,N_19762,N_20345);
or U21242 (N_21242,N_20919,N_20726);
nand U21243 (N_21243,N_20621,N_20152);
and U21244 (N_21244,N_20944,N_19852);
nand U21245 (N_21245,N_20206,N_20015);
and U21246 (N_21246,N_20787,N_20462);
and U21247 (N_21247,N_20480,N_20292);
xnor U21248 (N_21248,N_19966,N_20597);
xnor U21249 (N_21249,N_19843,N_19799);
and U21250 (N_21250,N_19706,N_20754);
nand U21251 (N_21251,N_20564,N_20947);
nor U21252 (N_21252,N_19873,N_20732);
xor U21253 (N_21253,N_20140,N_20833);
nand U21254 (N_21254,N_19508,N_20760);
nand U21255 (N_21255,N_20516,N_19892);
xnor U21256 (N_21256,N_20808,N_20348);
nor U21257 (N_21257,N_19859,N_20135);
nand U21258 (N_21258,N_20043,N_19959);
and U21259 (N_21259,N_20967,N_19757);
xor U21260 (N_21260,N_20233,N_20243);
xor U21261 (N_21261,N_20942,N_19888);
xor U21262 (N_21262,N_20350,N_20619);
xnor U21263 (N_21263,N_20599,N_20209);
and U21264 (N_21264,N_19641,N_19645);
nor U21265 (N_21265,N_20768,N_19789);
nand U21266 (N_21266,N_20624,N_20392);
nand U21267 (N_21267,N_20673,N_20686);
and U21268 (N_21268,N_20971,N_19654);
nand U21269 (N_21269,N_20102,N_19546);
xnor U21270 (N_21270,N_20107,N_20394);
and U21271 (N_21271,N_20204,N_20038);
nand U21272 (N_21272,N_20792,N_20437);
and U21273 (N_21273,N_20063,N_19695);
nor U21274 (N_21274,N_19614,N_19633);
nand U21275 (N_21275,N_20743,N_20299);
nand U21276 (N_21276,N_19827,N_20115);
nor U21277 (N_21277,N_19562,N_20415);
and U21278 (N_21278,N_19862,N_19995);
xnor U21279 (N_21279,N_19699,N_20100);
nor U21280 (N_21280,N_20241,N_19647);
xor U21281 (N_21281,N_20554,N_19878);
xnor U21282 (N_21282,N_19944,N_19994);
or U21283 (N_21283,N_19819,N_19653);
nand U21284 (N_21284,N_19718,N_19510);
or U21285 (N_21285,N_20326,N_19719);
nor U21286 (N_21286,N_19838,N_19906);
xnor U21287 (N_21287,N_20429,N_19781);
nand U21288 (N_21288,N_20224,N_19961);
and U21289 (N_21289,N_20422,N_20487);
xor U21290 (N_21290,N_19623,N_20481);
and U21291 (N_21291,N_20117,N_20563);
nor U21292 (N_21292,N_20763,N_19810);
or U21293 (N_21293,N_19551,N_20932);
nor U21294 (N_21294,N_19796,N_20632);
xnor U21295 (N_21295,N_20720,N_20986);
or U21296 (N_21296,N_19723,N_20237);
or U21297 (N_21297,N_20068,N_19526);
xor U21298 (N_21298,N_20729,N_20288);
xor U21299 (N_21299,N_20280,N_20802);
and U21300 (N_21300,N_19822,N_20550);
nand U21301 (N_21301,N_20404,N_20925);
xor U21302 (N_21302,N_20953,N_19674);
and U21303 (N_21303,N_19834,N_20134);
or U21304 (N_21304,N_19910,N_19890);
xnor U21305 (N_21305,N_20008,N_19997);
xnor U21306 (N_21306,N_19624,N_19515);
nand U21307 (N_21307,N_19752,N_20098);
nor U21308 (N_21308,N_20214,N_20114);
and U21309 (N_21309,N_20934,N_20499);
or U21310 (N_21310,N_20476,N_20945);
xor U21311 (N_21311,N_20228,N_20402);
xnor U21312 (N_21312,N_20364,N_19786);
and U21313 (N_21313,N_20301,N_20290);
and U21314 (N_21314,N_20645,N_20445);
nand U21315 (N_21315,N_20748,N_19636);
or U21316 (N_21316,N_19875,N_20375);
nor U21317 (N_21317,N_20764,N_19831);
and U21318 (N_21318,N_20612,N_20815);
nand U21319 (N_21319,N_20788,N_20069);
or U21320 (N_21320,N_19803,N_20937);
or U21321 (N_21321,N_20075,N_20901);
nand U21322 (N_21322,N_19912,N_20169);
and U21323 (N_21323,N_20153,N_20433);
nor U21324 (N_21324,N_20538,N_19973);
xnor U21325 (N_21325,N_20772,N_20739);
nand U21326 (N_21326,N_20358,N_20156);
nor U21327 (N_21327,N_20848,N_19801);
nand U21328 (N_21328,N_20475,N_20011);
xnor U21329 (N_21329,N_19858,N_19857);
xor U21330 (N_21330,N_20066,N_20270);
nor U21331 (N_21331,N_19626,N_20663);
nand U21332 (N_21332,N_20633,N_19541);
nand U21333 (N_21333,N_19710,N_19730);
nor U21334 (N_21334,N_20713,N_19788);
xor U21335 (N_21335,N_20471,N_20923);
or U21336 (N_21336,N_19635,N_19612);
or U21337 (N_21337,N_20027,N_20256);
nand U21338 (N_21338,N_19597,N_20617);
nor U21339 (N_21339,N_19622,N_19505);
xnor U21340 (N_21340,N_20251,N_19600);
and U21341 (N_21341,N_19918,N_20988);
xor U21342 (N_21342,N_20474,N_20671);
nand U21343 (N_21343,N_20253,N_20312);
or U21344 (N_21344,N_19599,N_20614);
and U21345 (N_21345,N_19701,N_20161);
and U21346 (N_21346,N_19751,N_20699);
xor U21347 (N_21347,N_19611,N_19527);
or U21348 (N_21348,N_20877,N_19691);
or U21349 (N_21349,N_20634,N_20167);
xnor U21350 (N_21350,N_20895,N_19931);
xnor U21351 (N_21351,N_20864,N_20886);
nor U21352 (N_21352,N_19514,N_19908);
nor U21353 (N_21353,N_20349,N_19960);
nor U21354 (N_21354,N_19897,N_20609);
xnor U21355 (N_21355,N_20125,N_19602);
or U21356 (N_21356,N_19634,N_20463);
xnor U21357 (N_21357,N_20631,N_20020);
nand U21358 (N_21358,N_19662,N_19924);
nor U21359 (N_21359,N_20637,N_20750);
and U21360 (N_21360,N_19631,N_20190);
nand U21361 (N_21361,N_20372,N_20765);
nor U21362 (N_21362,N_20606,N_20987);
nor U21363 (N_21363,N_19812,N_20148);
and U21364 (N_21364,N_20820,N_20447);
nor U21365 (N_21365,N_19953,N_19764);
nor U21366 (N_21366,N_20158,N_19916);
xnor U21367 (N_21367,N_20514,N_20426);
nor U21368 (N_21368,N_20078,N_19501);
nand U21369 (N_21369,N_20282,N_20641);
xnor U21370 (N_21370,N_20193,N_20723);
and U21371 (N_21371,N_19975,N_19720);
xor U21372 (N_21372,N_19596,N_20235);
or U21373 (N_21373,N_19517,N_20522);
nor U21374 (N_21374,N_20208,N_20889);
nand U21375 (N_21375,N_19703,N_19539);
and U21376 (N_21376,N_20286,N_20844);
nor U21377 (N_21377,N_20091,N_19556);
and U21378 (N_21378,N_19828,N_19571);
and U21379 (N_21379,N_20484,N_20681);
nand U21380 (N_21380,N_20547,N_19980);
nor U21381 (N_21381,N_20596,N_20354);
xnor U21382 (N_21382,N_19914,N_20121);
or U21383 (N_21383,N_20245,N_19721);
or U21384 (N_21384,N_20187,N_20841);
nor U21385 (N_21385,N_20377,N_20200);
nand U21386 (N_21386,N_19826,N_20449);
or U21387 (N_21387,N_20054,N_19670);
xor U21388 (N_21388,N_19523,N_20859);
and U21389 (N_21389,N_19915,N_20325);
nand U21390 (N_21390,N_20799,N_20412);
nand U21391 (N_21391,N_20845,N_19927);
nor U21392 (N_21392,N_20527,N_20336);
xnor U21393 (N_21393,N_19567,N_20838);
xor U21394 (N_21394,N_19970,N_20388);
nand U21395 (N_21395,N_20459,N_20477);
nand U21396 (N_21396,N_19845,N_20460);
and U21397 (N_21397,N_20414,N_19566);
nand U21398 (N_21398,N_20432,N_20721);
nand U21399 (N_21399,N_20316,N_20647);
or U21400 (N_21400,N_19936,N_20373);
xnor U21401 (N_21401,N_20034,N_20283);
or U21402 (N_21402,N_19742,N_19798);
or U21403 (N_21403,N_19879,N_20810);
nand U21404 (N_21404,N_19709,N_20830);
nand U21405 (N_21405,N_20355,N_20465);
xnor U21406 (N_21406,N_20997,N_20252);
and U21407 (N_21407,N_20989,N_19996);
nor U21408 (N_21408,N_19785,N_20741);
or U21409 (N_21409,N_19632,N_20219);
and U21410 (N_21410,N_20163,N_20846);
nor U21411 (N_21411,N_20774,N_20608);
and U21412 (N_21412,N_20706,N_19557);
nor U21413 (N_21413,N_20116,N_20419);
nand U21414 (N_21414,N_20457,N_19575);
xor U21415 (N_21415,N_20293,N_20400);
nor U21416 (N_21416,N_20981,N_19661);
xnor U21417 (N_21417,N_20551,N_20277);
or U21418 (N_21418,N_19754,N_19737);
nor U21419 (N_21419,N_20984,N_20005);
nor U21420 (N_21420,N_19666,N_20767);
xor U21421 (N_21421,N_19772,N_19568);
and U21422 (N_21422,N_20883,N_20994);
and U21423 (N_21423,N_20133,N_19948);
and U21424 (N_21424,N_20724,N_20041);
nor U21425 (N_21425,N_19864,N_19889);
and U21426 (N_21426,N_20805,N_20018);
and U21427 (N_21427,N_20232,N_20329);
and U21428 (N_21428,N_19792,N_19876);
nand U21429 (N_21429,N_20770,N_19528);
or U21430 (N_21430,N_20151,N_20284);
or U21431 (N_21431,N_20302,N_20785);
and U21432 (N_21432,N_20950,N_20077);
or U21433 (N_21433,N_20524,N_20829);
nor U21434 (N_21434,N_20371,N_20026);
nand U21435 (N_21435,N_19547,N_20397);
or U21436 (N_21436,N_20454,N_19582);
nor U21437 (N_21437,N_20317,N_19794);
and U21438 (N_21438,N_20570,N_20752);
or U21439 (N_21439,N_19962,N_19716);
nand U21440 (N_21440,N_20178,N_20319);
xor U21441 (N_21441,N_19667,N_20589);
and U21442 (N_21442,N_20123,N_20217);
or U21443 (N_21443,N_20058,N_20401);
nand U21444 (N_21444,N_20420,N_19646);
nand U21445 (N_21445,N_20222,N_19656);
and U21446 (N_21446,N_19923,N_20534);
or U21447 (N_21447,N_19545,N_19837);
and U21448 (N_21448,N_20455,N_20935);
xnor U21449 (N_21449,N_20529,N_19867);
nand U21450 (N_21450,N_20164,N_19639);
nor U21451 (N_21451,N_20927,N_20022);
and U21452 (N_21452,N_19809,N_19749);
and U21453 (N_21453,N_19593,N_20510);
nor U21454 (N_21454,N_20890,N_20150);
or U21455 (N_21455,N_20096,N_19583);
or U21456 (N_21456,N_20436,N_19871);
and U21457 (N_21457,N_19570,N_20221);
xnor U21458 (N_21458,N_20884,N_20165);
or U21459 (N_21459,N_20196,N_20007);
or U21460 (N_21460,N_20941,N_20223);
nor U21461 (N_21461,N_19901,N_20320);
and U21462 (N_21462,N_19620,N_20246);
and U21463 (N_21463,N_20703,N_20917);
and U21464 (N_21464,N_19529,N_20811);
nand U21465 (N_21465,N_19780,N_19832);
nor U21466 (N_21466,N_19644,N_20801);
or U21467 (N_21467,N_19673,N_19669);
nor U21468 (N_21468,N_20191,N_20337);
or U21469 (N_21469,N_19531,N_20588);
and U21470 (N_21470,N_20101,N_20891);
nor U21471 (N_21471,N_19580,N_20461);
or U21472 (N_21472,N_20490,N_20777);
nor U21473 (N_21473,N_20574,N_20579);
or U21474 (N_21474,N_20561,N_20783);
or U21475 (N_21475,N_20194,N_20897);
xnor U21476 (N_21476,N_20955,N_20648);
nor U21477 (N_21477,N_19572,N_20079);
or U21478 (N_21478,N_20186,N_20327);
or U21479 (N_21479,N_20684,N_19629);
nor U21480 (N_21480,N_19998,N_20488);
nor U21481 (N_21481,N_20881,N_20197);
nor U21482 (N_21482,N_20255,N_20870);
nand U21483 (N_21483,N_19591,N_20468);
and U21484 (N_21484,N_19601,N_19680);
nand U21485 (N_21485,N_20540,N_19671);
and U21486 (N_21486,N_20342,N_19983);
or U21487 (N_21487,N_20701,N_19769);
xor U21488 (N_21488,N_19896,N_19783);
nand U21489 (N_21489,N_20176,N_20340);
and U21490 (N_21490,N_19758,N_19564);
and U21491 (N_21491,N_19795,N_19642);
xnor U21492 (N_21492,N_20379,N_19941);
or U21493 (N_21493,N_20168,N_19500);
or U21494 (N_21494,N_20998,N_19999);
xnor U21495 (N_21495,N_20324,N_19736);
and U21496 (N_21496,N_19882,N_20511);
nor U21497 (N_21497,N_19696,N_20779);
nor U21498 (N_21498,N_19986,N_19884);
nand U21499 (N_21499,N_19952,N_20710);
nand U21500 (N_21500,N_20778,N_19678);
nor U21501 (N_21501,N_20306,N_20322);
or U21502 (N_21502,N_20231,N_20031);
xnor U21503 (N_21503,N_19886,N_19956);
and U21504 (N_21504,N_20558,N_19722);
or U21505 (N_21505,N_20876,N_19784);
and U21506 (N_21506,N_19779,N_20162);
and U21507 (N_21507,N_19968,N_19586);
or U21508 (N_21508,N_20674,N_19979);
xor U21509 (N_21509,N_20595,N_20666);
nand U21510 (N_21510,N_20308,N_19702);
nor U21511 (N_21511,N_20021,N_20578);
or U21512 (N_21512,N_20759,N_20727);
nor U21513 (N_21513,N_20369,N_20362);
or U21514 (N_21514,N_20338,N_20585);
and U21515 (N_21515,N_19938,N_20571);
nand U21516 (N_21516,N_20573,N_20092);
xnor U21517 (N_21517,N_20042,N_20285);
xor U21518 (N_21518,N_20183,N_20643);
and U21519 (N_21519,N_20590,N_19713);
xor U21520 (N_21520,N_20343,N_19544);
and U21521 (N_21521,N_19658,N_20916);
and U21522 (N_21522,N_19687,N_20174);
or U21523 (N_21523,N_20472,N_20908);
xnor U21524 (N_21524,N_20029,N_19657);
nor U21525 (N_21525,N_20800,N_19947);
or U21526 (N_21526,N_19506,N_19989);
nor U21527 (N_21527,N_19855,N_20085);
and U21528 (N_21528,N_20828,N_20498);
nand U21529 (N_21529,N_19940,N_20933);
nor U21530 (N_21530,N_20094,N_19778);
nand U21531 (N_21531,N_19903,N_20782);
and U21532 (N_21532,N_20798,N_20835);
or U21533 (N_21533,N_20060,N_20002);
or U21534 (N_21534,N_20059,N_20046);
xnor U21535 (N_21535,N_19569,N_20646);
xor U21536 (N_21536,N_20082,N_20321);
nor U21537 (N_21537,N_19760,N_20145);
or U21538 (N_21538,N_20268,N_20155);
and U21539 (N_21539,N_20898,N_20893);
and U21540 (N_21540,N_19708,N_19759);
and U21541 (N_21541,N_20144,N_20556);
nand U21542 (N_21542,N_19977,N_20242);
nand U21543 (N_21543,N_20936,N_20902);
nor U21544 (N_21544,N_20731,N_20139);
and U21545 (N_21545,N_19984,N_20718);
nor U21546 (N_21546,N_19804,N_20758);
nor U21547 (N_21547,N_20736,N_19971);
nand U21548 (N_21548,N_20616,N_20188);
xor U21549 (N_21549,N_20175,N_19949);
xnor U21550 (N_21550,N_20110,N_20656);
or U21551 (N_21551,N_19993,N_20304);
and U21552 (N_21552,N_20973,N_20536);
nand U21553 (N_21553,N_20618,N_20975);
and U21554 (N_21554,N_20218,N_20238);
xnor U21555 (N_21555,N_19887,N_20662);
nand U21556 (N_21556,N_19578,N_20396);
or U21557 (N_21557,N_19711,N_20716);
or U21558 (N_21558,N_20061,N_20048);
xor U21559 (N_21559,N_20513,N_20978);
and U21560 (N_21560,N_20287,N_20106);
or U21561 (N_21561,N_19615,N_20982);
or U21562 (N_21562,N_20920,N_20863);
or U21563 (N_21563,N_20430,N_20660);
nor U21564 (N_21564,N_19797,N_20128);
or U21565 (N_21565,N_20905,N_20827);
nor U21566 (N_21566,N_20565,N_20819);
and U21567 (N_21567,N_20365,N_20839);
xor U21568 (N_21568,N_20996,N_19840);
xnor U21569 (N_21569,N_20382,N_19697);
nand U21570 (N_21570,N_20260,N_19937);
or U21571 (N_21571,N_20003,N_20751);
nand U21572 (N_21572,N_20817,N_20591);
and U21573 (N_21573,N_20793,N_20600);
and U21574 (N_21574,N_20964,N_20130);
nand U21575 (N_21575,N_19744,N_20602);
or U21576 (N_21576,N_20070,N_19958);
and U21577 (N_21577,N_19905,N_19791);
and U21578 (N_21578,N_20464,N_20622);
nand U21579 (N_21579,N_19913,N_20980);
and U21580 (N_21580,N_20909,N_20207);
or U21581 (N_21581,N_20344,N_19537);
nor U21582 (N_21582,N_19727,N_19909);
xor U21583 (N_21583,N_20865,N_19853);
nand U21584 (N_21584,N_20972,N_20749);
nand U21585 (N_21585,N_20180,N_20620);
xnor U21586 (N_21586,N_20826,N_20331);
and U21587 (N_21587,N_20266,N_20677);
and U21588 (N_21588,N_20781,N_20289);
and U21589 (N_21589,N_20604,N_20549);
and U21590 (N_21590,N_20939,N_20249);
xnor U21591 (N_21591,N_19921,N_20272);
and U21592 (N_21592,N_20789,N_19942);
nor U21593 (N_21593,N_19806,N_20970);
xor U21594 (N_21594,N_20478,N_20341);
nor U21595 (N_21595,N_19613,N_20203);
nand U21596 (N_21596,N_19717,N_20611);
and U21597 (N_21597,N_20441,N_19558);
nand U21598 (N_21598,N_20541,N_20913);
nor U21599 (N_21599,N_19726,N_20659);
or U21600 (N_21600,N_20185,N_19967);
and U21601 (N_21601,N_20745,N_20411);
and U21602 (N_21602,N_19969,N_20796);
xor U21603 (N_21603,N_19734,N_20493);
or U21604 (N_21604,N_19607,N_20360);
or U21605 (N_21605,N_20976,N_19988);
xnor U21606 (N_21606,N_20416,N_20265);
nor U21607 (N_21607,N_19990,N_19991);
nor U21608 (N_21608,N_19584,N_20159);
nor U21609 (N_21609,N_20247,N_20832);
or U21610 (N_21610,N_19765,N_20057);
nand U21611 (N_21611,N_20179,N_20872);
xor U21612 (N_21612,N_19793,N_20064);
and U21613 (N_21613,N_20840,N_19740);
or U21614 (N_21614,N_19735,N_20818);
and U21615 (N_21615,N_20216,N_19520);
xor U21616 (N_21616,N_20281,N_19894);
or U21617 (N_21617,N_20368,N_20943);
nor U21618 (N_21618,N_20084,N_19790);
and U21619 (N_21619,N_19625,N_19761);
nand U21620 (N_21620,N_19755,N_19536);
nand U21621 (N_21621,N_20450,N_20899);
nor U21622 (N_21622,N_19802,N_20697);
or U21623 (N_21623,N_19731,N_20873);
nand U21624 (N_21624,N_20725,N_20572);
nor U21625 (N_21625,N_20867,N_20924);
nand U21626 (N_21626,N_20636,N_19563);
xnor U21627 (N_21627,N_19775,N_20257);
and U21628 (N_21628,N_20630,N_20201);
xnor U21629 (N_21629,N_20334,N_19899);
xor U21630 (N_21630,N_20276,N_19874);
and U21631 (N_21631,N_20047,N_20124);
xor U21632 (N_21632,N_20448,N_20383);
nand U21633 (N_21633,N_20181,N_19682);
nor U21634 (N_21634,N_19981,N_20119);
or U21635 (N_21635,N_19504,N_19848);
and U21636 (N_21636,N_20213,N_20010);
and U21637 (N_21637,N_19911,N_19560);
nand U21638 (N_21638,N_20250,N_20418);
xor U21639 (N_21639,N_20965,N_20294);
nand U21640 (N_21640,N_20122,N_20229);
or U21641 (N_21641,N_19513,N_20957);
nand U21642 (N_21642,N_20090,N_20000);
xor U21643 (N_21643,N_20427,N_19595);
xor U21644 (N_21644,N_20361,N_20239);
or U21645 (N_21645,N_20698,N_19787);
or U21646 (N_21646,N_20854,N_20730);
and U21647 (N_21647,N_20896,N_20649);
nand U21648 (N_21648,N_19679,N_19776);
and U21649 (N_21649,N_20530,N_20775);
nor U21650 (N_21650,N_20918,N_19839);
nand U21651 (N_21651,N_20505,N_19664);
or U21652 (N_21652,N_19660,N_20408);
xor U21653 (N_21653,N_20423,N_20129);
xor U21654 (N_21654,N_20625,N_20074);
or U21655 (N_21655,N_20143,N_20279);
and U21656 (N_21656,N_19550,N_20131);
nand U21657 (N_21657,N_19533,N_20492);
xor U21658 (N_21658,N_20330,N_20226);
nand U21659 (N_21659,N_20507,N_20906);
or U21660 (N_21660,N_19782,N_20836);
or U21661 (N_21661,N_20037,N_19535);
xor U21662 (N_21662,N_20773,N_20473);
and U21663 (N_21663,N_20756,N_20012);
nor U21664 (N_21664,N_20025,N_20431);
nand U21665 (N_21665,N_20878,N_19777);
or U21666 (N_21666,N_19951,N_20615);
or U21667 (N_21667,N_20470,N_20714);
and U21668 (N_21668,N_19585,N_19507);
or U21669 (N_21669,N_20295,N_19588);
xnor U21670 (N_21670,N_20120,N_19766);
and U21671 (N_21671,N_20305,N_20307);
nor U21672 (N_21672,N_20683,N_20531);
or U21673 (N_21673,N_20521,N_20205);
and U21674 (N_21674,N_19816,N_19630);
nor U21675 (N_21675,N_20508,N_20822);
nand U21676 (N_21676,N_20951,N_19524);
and U21677 (N_21677,N_20849,N_20962);
xor U21678 (N_21678,N_19540,N_19606);
nand U21679 (N_21679,N_20861,N_19538);
nand U21680 (N_21680,N_20300,N_19883);
nand U21681 (N_21681,N_20258,N_20328);
nor U21682 (N_21682,N_19681,N_20946);
or U21683 (N_21683,N_20635,N_20417);
or U21684 (N_21684,N_20875,N_19574);
or U21685 (N_21685,N_19920,N_20089);
xnor U21686 (N_21686,N_20230,N_20921);
and U21687 (N_21687,N_20407,N_19893);
or U21688 (N_21688,N_20722,N_20494);
nor U21689 (N_21689,N_20095,N_20500);
nor U21690 (N_21690,N_20440,N_19676);
xnor U21691 (N_21691,N_20707,N_19577);
nor U21692 (N_21692,N_19963,N_20347);
xor U21693 (N_21693,N_20199,N_20016);
nand U21694 (N_21694,N_20688,N_20539);
or U21695 (N_21695,N_19694,N_20757);
and U21696 (N_21696,N_20685,N_20126);
xnor U21697 (N_21697,N_20520,N_20692);
nor U21698 (N_21698,N_20451,N_20653);
nand U21699 (N_21699,N_20695,N_20629);
xor U21700 (N_21700,N_20024,N_20399);
or U21701 (N_21701,N_19688,N_20771);
nor U21702 (N_21702,N_19935,N_20809);
nand U21703 (N_21703,N_20248,N_20182);
and U21704 (N_21704,N_20842,N_20851);
and U21705 (N_21705,N_19519,N_19922);
or U21706 (N_21706,N_20518,N_19589);
xor U21707 (N_21707,N_20086,N_19846);
nand U21708 (N_21708,N_20553,N_20719);
and U21709 (N_21709,N_20067,N_20575);
or U21710 (N_21710,N_19825,N_19932);
nor U21711 (N_21711,N_19982,N_19549);
nand U21712 (N_21712,N_19756,N_20639);
or U21713 (N_21713,N_20393,N_19604);
xnor U21714 (N_21714,N_20118,N_19934);
and U21715 (N_21715,N_19773,N_20366);
nor U21716 (N_21716,N_20642,N_20613);
nor U21717 (N_21717,N_19976,N_19863);
or U21718 (N_21718,N_20562,N_19972);
nor U21719 (N_21719,N_20601,N_19648);
nor U21720 (N_21720,N_20603,N_20254);
xnor U21721 (N_21721,N_19686,N_20821);
and U21722 (N_21722,N_20019,N_20657);
nor U21723 (N_21723,N_20627,N_20977);
or U21724 (N_21724,N_20177,N_20049);
nor U21725 (N_21725,N_19850,N_20999);
xor U21726 (N_21726,N_19829,N_20594);
nor U21727 (N_21727,N_20914,N_20586);
nand U21728 (N_21728,N_19565,N_19747);
or U21729 (N_21729,N_20310,N_20211);
xor U21730 (N_21730,N_19902,N_19587);
nand U21731 (N_21731,N_20824,N_20922);
xnor U21732 (N_21732,N_20995,N_20911);
and U21733 (N_21733,N_20173,N_20744);
or U21734 (N_21734,N_20567,N_20652);
or U21735 (N_21735,N_20171,N_20780);
xnor U21736 (N_21736,N_19869,N_20623);
and U21737 (N_21737,N_19692,N_20405);
xor U21738 (N_21738,N_20073,N_20303);
and U21739 (N_21739,N_20391,N_19594);
xor U21740 (N_21740,N_19509,N_20903);
nor U21741 (N_21741,N_20497,N_20928);
xor U21742 (N_21742,N_20679,N_20992);
xor U21743 (N_21743,N_19715,N_20528);
nand U21744 (N_21744,N_20803,N_20866);
and U21745 (N_21745,N_20390,N_19553);
or U21746 (N_21746,N_20384,N_20099);
and U21747 (N_21747,N_19532,N_19808);
nor U21748 (N_21748,N_20717,N_20087);
nor U21749 (N_21749,N_20458,N_20825);
nor U21750 (N_21750,N_20101,N_20424);
and U21751 (N_21751,N_19961,N_19870);
nand U21752 (N_21752,N_20308,N_20143);
or U21753 (N_21753,N_19780,N_20912);
nand U21754 (N_21754,N_20355,N_20454);
and U21755 (N_21755,N_20757,N_19728);
and U21756 (N_21756,N_19714,N_20826);
nor U21757 (N_21757,N_20106,N_20384);
nor U21758 (N_21758,N_20479,N_20243);
or U21759 (N_21759,N_20649,N_20035);
nor U21760 (N_21760,N_19596,N_19682);
and U21761 (N_21761,N_20260,N_19590);
xnor U21762 (N_21762,N_19594,N_19544);
and U21763 (N_21763,N_20176,N_20064);
nor U21764 (N_21764,N_20079,N_20500);
nor U21765 (N_21765,N_19670,N_19902);
and U21766 (N_21766,N_19611,N_20014);
nand U21767 (N_21767,N_19801,N_19838);
and U21768 (N_21768,N_20699,N_20634);
nor U21769 (N_21769,N_19902,N_20495);
and U21770 (N_21770,N_20142,N_19504);
or U21771 (N_21771,N_19831,N_20644);
xnor U21772 (N_21772,N_20343,N_19608);
and U21773 (N_21773,N_19770,N_20351);
and U21774 (N_21774,N_20211,N_20550);
or U21775 (N_21775,N_20857,N_20045);
xnor U21776 (N_21776,N_20385,N_20777);
nand U21777 (N_21777,N_20974,N_19933);
nor U21778 (N_21778,N_20349,N_20159);
and U21779 (N_21779,N_20798,N_20171);
nand U21780 (N_21780,N_19564,N_19935);
xor U21781 (N_21781,N_20861,N_20820);
xnor U21782 (N_21782,N_20297,N_20955);
xnor U21783 (N_21783,N_19622,N_20086);
xor U21784 (N_21784,N_20892,N_20299);
nand U21785 (N_21785,N_20428,N_20347);
nor U21786 (N_21786,N_20724,N_20732);
nand U21787 (N_21787,N_20588,N_19523);
nand U21788 (N_21788,N_20854,N_20528);
nand U21789 (N_21789,N_20230,N_20470);
or U21790 (N_21790,N_19875,N_20014);
nand U21791 (N_21791,N_20293,N_20236);
xnor U21792 (N_21792,N_20605,N_20768);
or U21793 (N_21793,N_20157,N_20148);
xnor U21794 (N_21794,N_20958,N_19636);
nor U21795 (N_21795,N_19690,N_20963);
xor U21796 (N_21796,N_20113,N_20220);
nor U21797 (N_21797,N_19782,N_20177);
xor U21798 (N_21798,N_20813,N_20238);
or U21799 (N_21799,N_20316,N_20866);
or U21800 (N_21800,N_20619,N_20225);
or U21801 (N_21801,N_20373,N_20842);
and U21802 (N_21802,N_20071,N_20075);
and U21803 (N_21803,N_20816,N_20839);
nor U21804 (N_21804,N_19658,N_19547);
and U21805 (N_21805,N_20918,N_19531);
and U21806 (N_21806,N_20911,N_19777);
and U21807 (N_21807,N_20638,N_19644);
and U21808 (N_21808,N_20588,N_20892);
xor U21809 (N_21809,N_20891,N_19776);
or U21810 (N_21810,N_19719,N_19665);
nor U21811 (N_21811,N_20211,N_20488);
and U21812 (N_21812,N_20823,N_20971);
nor U21813 (N_21813,N_20881,N_20999);
nand U21814 (N_21814,N_20044,N_20549);
or U21815 (N_21815,N_20239,N_20754);
nor U21816 (N_21816,N_20062,N_20402);
or U21817 (N_21817,N_20718,N_19542);
and U21818 (N_21818,N_20979,N_20932);
and U21819 (N_21819,N_20034,N_19811);
or U21820 (N_21820,N_20429,N_20440);
xnor U21821 (N_21821,N_19931,N_20783);
and U21822 (N_21822,N_19523,N_20231);
and U21823 (N_21823,N_20599,N_20468);
and U21824 (N_21824,N_19572,N_20048);
nand U21825 (N_21825,N_20294,N_19629);
or U21826 (N_21826,N_20842,N_20091);
nand U21827 (N_21827,N_19509,N_20661);
nor U21828 (N_21828,N_20894,N_20361);
nor U21829 (N_21829,N_20747,N_19574);
and U21830 (N_21830,N_20608,N_19514);
or U21831 (N_21831,N_20496,N_20960);
nand U21832 (N_21832,N_19920,N_19846);
nor U21833 (N_21833,N_20791,N_19709);
nand U21834 (N_21834,N_20810,N_20661);
or U21835 (N_21835,N_20197,N_20841);
nor U21836 (N_21836,N_20013,N_20110);
or U21837 (N_21837,N_20949,N_19829);
and U21838 (N_21838,N_19981,N_19572);
xnor U21839 (N_21839,N_20203,N_19976);
xnor U21840 (N_21840,N_19959,N_20198);
xnor U21841 (N_21841,N_20825,N_19921);
or U21842 (N_21842,N_20093,N_20880);
and U21843 (N_21843,N_20992,N_19593);
and U21844 (N_21844,N_20072,N_19917);
and U21845 (N_21845,N_20655,N_19599);
and U21846 (N_21846,N_20704,N_19999);
or U21847 (N_21847,N_20982,N_20409);
and U21848 (N_21848,N_20312,N_19631);
xor U21849 (N_21849,N_19550,N_20648);
nand U21850 (N_21850,N_20542,N_20960);
nor U21851 (N_21851,N_19691,N_20128);
nor U21852 (N_21852,N_20038,N_20100);
nand U21853 (N_21853,N_20349,N_19971);
xor U21854 (N_21854,N_20747,N_19628);
nand U21855 (N_21855,N_19934,N_20106);
and U21856 (N_21856,N_20974,N_19885);
or U21857 (N_21857,N_20461,N_19789);
xnor U21858 (N_21858,N_20673,N_19886);
xnor U21859 (N_21859,N_20406,N_20523);
xor U21860 (N_21860,N_20262,N_20391);
nor U21861 (N_21861,N_19578,N_19627);
and U21862 (N_21862,N_20108,N_20009);
nand U21863 (N_21863,N_20175,N_20561);
nor U21864 (N_21864,N_19979,N_20647);
xnor U21865 (N_21865,N_20737,N_19729);
and U21866 (N_21866,N_20272,N_19959);
and U21867 (N_21867,N_20856,N_20439);
nor U21868 (N_21868,N_20157,N_20397);
nand U21869 (N_21869,N_20567,N_20656);
nand U21870 (N_21870,N_19980,N_20065);
or U21871 (N_21871,N_20890,N_20194);
and U21872 (N_21872,N_20140,N_19949);
nand U21873 (N_21873,N_19869,N_19933);
nand U21874 (N_21874,N_20674,N_20677);
nor U21875 (N_21875,N_20631,N_19690);
nor U21876 (N_21876,N_19647,N_19516);
or U21877 (N_21877,N_20245,N_20348);
nor U21878 (N_21878,N_20927,N_19626);
or U21879 (N_21879,N_20268,N_20334);
xor U21880 (N_21880,N_20203,N_20255);
nor U21881 (N_21881,N_20125,N_20835);
nor U21882 (N_21882,N_20096,N_19553);
or U21883 (N_21883,N_19780,N_20735);
and U21884 (N_21884,N_19510,N_19641);
nand U21885 (N_21885,N_20609,N_20576);
xnor U21886 (N_21886,N_20515,N_19857);
nand U21887 (N_21887,N_19763,N_20475);
nor U21888 (N_21888,N_20569,N_19895);
nand U21889 (N_21889,N_20995,N_19812);
or U21890 (N_21890,N_19990,N_19935);
xor U21891 (N_21891,N_20430,N_20637);
and U21892 (N_21892,N_20505,N_19751);
or U21893 (N_21893,N_20829,N_19735);
nand U21894 (N_21894,N_20058,N_20062);
nor U21895 (N_21895,N_20890,N_20940);
or U21896 (N_21896,N_20180,N_20182);
nor U21897 (N_21897,N_19515,N_19900);
and U21898 (N_21898,N_20040,N_20392);
and U21899 (N_21899,N_20565,N_19731);
or U21900 (N_21900,N_19887,N_20582);
and U21901 (N_21901,N_20756,N_20292);
or U21902 (N_21902,N_20066,N_19893);
nor U21903 (N_21903,N_20097,N_20686);
xnor U21904 (N_21904,N_19520,N_19943);
or U21905 (N_21905,N_20833,N_20486);
and U21906 (N_21906,N_20951,N_20339);
or U21907 (N_21907,N_19533,N_20340);
and U21908 (N_21908,N_20614,N_20924);
xnor U21909 (N_21909,N_20589,N_20445);
nor U21910 (N_21910,N_19896,N_20217);
xor U21911 (N_21911,N_20468,N_19986);
nand U21912 (N_21912,N_20413,N_20763);
nand U21913 (N_21913,N_19515,N_20793);
nand U21914 (N_21914,N_20675,N_20562);
and U21915 (N_21915,N_19620,N_20776);
or U21916 (N_21916,N_19686,N_20015);
and U21917 (N_21917,N_20334,N_19977);
or U21918 (N_21918,N_19724,N_20547);
or U21919 (N_21919,N_19739,N_19677);
nor U21920 (N_21920,N_20275,N_20433);
and U21921 (N_21921,N_20071,N_19772);
xnor U21922 (N_21922,N_20632,N_20290);
nand U21923 (N_21923,N_20686,N_19507);
nor U21924 (N_21924,N_19630,N_19663);
xnor U21925 (N_21925,N_20224,N_20174);
nor U21926 (N_21926,N_20600,N_20238);
nand U21927 (N_21927,N_20378,N_20779);
and U21928 (N_21928,N_20715,N_20253);
and U21929 (N_21929,N_20862,N_20304);
or U21930 (N_21930,N_20373,N_19826);
xnor U21931 (N_21931,N_19801,N_20225);
xor U21932 (N_21932,N_20006,N_20572);
nor U21933 (N_21933,N_20596,N_19530);
or U21934 (N_21934,N_20237,N_20190);
and U21935 (N_21935,N_20063,N_19641);
xor U21936 (N_21936,N_19806,N_20905);
and U21937 (N_21937,N_20382,N_20432);
nand U21938 (N_21938,N_20287,N_19763);
nand U21939 (N_21939,N_20573,N_20324);
or U21940 (N_21940,N_19934,N_20580);
nor U21941 (N_21941,N_20861,N_20218);
or U21942 (N_21942,N_19529,N_20242);
xor U21943 (N_21943,N_20570,N_20187);
and U21944 (N_21944,N_19871,N_19639);
xnor U21945 (N_21945,N_20977,N_19885);
or U21946 (N_21946,N_20745,N_20824);
and U21947 (N_21947,N_20957,N_20858);
nand U21948 (N_21948,N_20832,N_20088);
xnor U21949 (N_21949,N_19718,N_20407);
xor U21950 (N_21950,N_20516,N_20640);
or U21951 (N_21951,N_19585,N_20388);
nand U21952 (N_21952,N_19527,N_20871);
xor U21953 (N_21953,N_20100,N_19619);
and U21954 (N_21954,N_20076,N_20957);
nor U21955 (N_21955,N_19527,N_20618);
and U21956 (N_21956,N_20515,N_20584);
nand U21957 (N_21957,N_20488,N_20919);
or U21958 (N_21958,N_20276,N_20338);
nand U21959 (N_21959,N_19847,N_20910);
xor U21960 (N_21960,N_20479,N_20834);
xor U21961 (N_21961,N_19965,N_20635);
or U21962 (N_21962,N_20696,N_20074);
xor U21963 (N_21963,N_19638,N_20405);
nor U21964 (N_21964,N_19550,N_19695);
nor U21965 (N_21965,N_20961,N_19744);
xor U21966 (N_21966,N_20281,N_20304);
nand U21967 (N_21967,N_20253,N_20817);
nand U21968 (N_21968,N_20284,N_20925);
xor U21969 (N_21969,N_19910,N_20162);
nor U21970 (N_21970,N_20403,N_19727);
nand U21971 (N_21971,N_19852,N_19886);
xor U21972 (N_21972,N_19726,N_19798);
or U21973 (N_21973,N_20043,N_19613);
nand U21974 (N_21974,N_20033,N_20518);
xnor U21975 (N_21975,N_20197,N_20969);
or U21976 (N_21976,N_20638,N_19595);
nor U21977 (N_21977,N_19573,N_19733);
xor U21978 (N_21978,N_20068,N_19885);
or U21979 (N_21979,N_20845,N_19530);
nor U21980 (N_21980,N_20512,N_20468);
or U21981 (N_21981,N_19972,N_19575);
or U21982 (N_21982,N_20840,N_20270);
xor U21983 (N_21983,N_20489,N_20838);
or U21984 (N_21984,N_20842,N_19912);
and U21985 (N_21985,N_19792,N_20452);
or U21986 (N_21986,N_20689,N_20094);
nor U21987 (N_21987,N_20068,N_20315);
and U21988 (N_21988,N_19792,N_20298);
and U21989 (N_21989,N_19665,N_20690);
and U21990 (N_21990,N_20591,N_19808);
nand U21991 (N_21991,N_19808,N_20585);
or U21992 (N_21992,N_20428,N_20894);
nand U21993 (N_21993,N_20209,N_20120);
nor U21994 (N_21994,N_20717,N_20103);
nand U21995 (N_21995,N_20784,N_20537);
or U21996 (N_21996,N_20021,N_20628);
xnor U21997 (N_21997,N_20022,N_20220);
and U21998 (N_21998,N_20402,N_19990);
nand U21999 (N_21999,N_20936,N_19717);
nor U22000 (N_22000,N_20579,N_20917);
and U22001 (N_22001,N_20791,N_19975);
xor U22002 (N_22002,N_20898,N_19629);
xnor U22003 (N_22003,N_20457,N_20385);
or U22004 (N_22004,N_20587,N_19610);
xor U22005 (N_22005,N_20575,N_20026);
or U22006 (N_22006,N_19747,N_20141);
xnor U22007 (N_22007,N_20055,N_20573);
or U22008 (N_22008,N_20285,N_19813);
and U22009 (N_22009,N_19856,N_19695);
and U22010 (N_22010,N_20880,N_19828);
xnor U22011 (N_22011,N_20496,N_19934);
nand U22012 (N_22012,N_20276,N_20868);
xor U22013 (N_22013,N_20542,N_19955);
and U22014 (N_22014,N_19719,N_19966);
and U22015 (N_22015,N_19788,N_19946);
nor U22016 (N_22016,N_20116,N_19768);
xnor U22017 (N_22017,N_20661,N_19590);
xnor U22018 (N_22018,N_20540,N_19532);
and U22019 (N_22019,N_19965,N_19760);
nand U22020 (N_22020,N_19816,N_20862);
nor U22021 (N_22021,N_20170,N_20304);
and U22022 (N_22022,N_20398,N_19533);
or U22023 (N_22023,N_19635,N_20887);
nor U22024 (N_22024,N_20698,N_20860);
nand U22025 (N_22025,N_19964,N_19920);
nor U22026 (N_22026,N_20471,N_20299);
or U22027 (N_22027,N_20511,N_19791);
nor U22028 (N_22028,N_19860,N_20107);
nor U22029 (N_22029,N_20641,N_19883);
xor U22030 (N_22030,N_20421,N_20137);
nor U22031 (N_22031,N_20874,N_20802);
nand U22032 (N_22032,N_20905,N_20299);
xnor U22033 (N_22033,N_20769,N_20452);
nand U22034 (N_22034,N_19893,N_20489);
nor U22035 (N_22035,N_19916,N_20753);
nor U22036 (N_22036,N_20941,N_20363);
xnor U22037 (N_22037,N_20030,N_20258);
nor U22038 (N_22038,N_20840,N_20877);
nand U22039 (N_22039,N_20973,N_20884);
xnor U22040 (N_22040,N_20361,N_19761);
xnor U22041 (N_22041,N_19811,N_19903);
and U22042 (N_22042,N_19790,N_20809);
and U22043 (N_22043,N_19639,N_20506);
and U22044 (N_22044,N_19858,N_20056);
and U22045 (N_22045,N_20801,N_20909);
nor U22046 (N_22046,N_19816,N_19717);
xnor U22047 (N_22047,N_20988,N_19778);
nand U22048 (N_22048,N_20520,N_20166);
nor U22049 (N_22049,N_20681,N_20148);
xnor U22050 (N_22050,N_19805,N_19931);
or U22051 (N_22051,N_20997,N_20235);
nand U22052 (N_22052,N_20309,N_20426);
or U22053 (N_22053,N_20152,N_20877);
nand U22054 (N_22054,N_19832,N_20326);
nand U22055 (N_22055,N_20668,N_20444);
and U22056 (N_22056,N_19669,N_20809);
nor U22057 (N_22057,N_20049,N_20212);
nor U22058 (N_22058,N_20445,N_20551);
or U22059 (N_22059,N_20439,N_20473);
or U22060 (N_22060,N_20170,N_20462);
nor U22061 (N_22061,N_20483,N_20638);
or U22062 (N_22062,N_19613,N_19522);
xnor U22063 (N_22063,N_19545,N_20023);
nor U22064 (N_22064,N_20681,N_20437);
nor U22065 (N_22065,N_20418,N_20630);
or U22066 (N_22066,N_20659,N_20081);
nand U22067 (N_22067,N_19530,N_20358);
nand U22068 (N_22068,N_19924,N_20302);
and U22069 (N_22069,N_20996,N_20271);
xnor U22070 (N_22070,N_20127,N_19563);
and U22071 (N_22071,N_19508,N_20499);
nor U22072 (N_22072,N_20074,N_20067);
xor U22073 (N_22073,N_20015,N_20691);
and U22074 (N_22074,N_20183,N_19526);
xnor U22075 (N_22075,N_20476,N_20185);
and U22076 (N_22076,N_20196,N_19858);
or U22077 (N_22077,N_20824,N_20247);
nand U22078 (N_22078,N_20666,N_20414);
nor U22079 (N_22079,N_20980,N_20221);
nor U22080 (N_22080,N_20849,N_19906);
xor U22081 (N_22081,N_20390,N_20569);
xnor U22082 (N_22082,N_20257,N_20639);
xnor U22083 (N_22083,N_20814,N_20898);
xnor U22084 (N_22084,N_20128,N_20713);
or U22085 (N_22085,N_20871,N_19518);
or U22086 (N_22086,N_19839,N_20925);
xor U22087 (N_22087,N_20614,N_20362);
xor U22088 (N_22088,N_19869,N_20505);
xnor U22089 (N_22089,N_20639,N_20720);
or U22090 (N_22090,N_20213,N_19738);
or U22091 (N_22091,N_20533,N_19564);
and U22092 (N_22092,N_20517,N_20311);
xnor U22093 (N_22093,N_20859,N_19708);
nor U22094 (N_22094,N_20893,N_20749);
and U22095 (N_22095,N_19820,N_19911);
xnor U22096 (N_22096,N_19803,N_20413);
or U22097 (N_22097,N_19868,N_19554);
nor U22098 (N_22098,N_20811,N_20946);
nand U22099 (N_22099,N_19991,N_20804);
nand U22100 (N_22100,N_20929,N_20614);
nor U22101 (N_22101,N_20767,N_19791);
nor U22102 (N_22102,N_20619,N_20055);
nand U22103 (N_22103,N_19820,N_19626);
nor U22104 (N_22104,N_20602,N_20584);
and U22105 (N_22105,N_20935,N_19613);
nand U22106 (N_22106,N_20325,N_20687);
xor U22107 (N_22107,N_20872,N_19689);
nand U22108 (N_22108,N_19563,N_20475);
xnor U22109 (N_22109,N_19810,N_20214);
nor U22110 (N_22110,N_20110,N_19721);
or U22111 (N_22111,N_20276,N_20433);
nor U22112 (N_22112,N_19751,N_20447);
xor U22113 (N_22113,N_20984,N_20084);
and U22114 (N_22114,N_20536,N_19599);
nor U22115 (N_22115,N_19778,N_20252);
nand U22116 (N_22116,N_20096,N_20117);
xor U22117 (N_22117,N_19730,N_20084);
xnor U22118 (N_22118,N_20870,N_20728);
nor U22119 (N_22119,N_20098,N_20388);
nand U22120 (N_22120,N_20348,N_19653);
or U22121 (N_22121,N_19964,N_20414);
and U22122 (N_22122,N_20311,N_20658);
or U22123 (N_22123,N_20390,N_20753);
nand U22124 (N_22124,N_20650,N_19807);
and U22125 (N_22125,N_20736,N_19554);
nor U22126 (N_22126,N_20089,N_19631);
xor U22127 (N_22127,N_20864,N_20662);
or U22128 (N_22128,N_20127,N_20921);
nor U22129 (N_22129,N_19570,N_19504);
and U22130 (N_22130,N_20583,N_19814);
and U22131 (N_22131,N_20421,N_20185);
nor U22132 (N_22132,N_19672,N_20186);
xor U22133 (N_22133,N_20106,N_20718);
or U22134 (N_22134,N_20937,N_19817);
nand U22135 (N_22135,N_20922,N_19582);
nor U22136 (N_22136,N_20063,N_19891);
xor U22137 (N_22137,N_20944,N_20963);
or U22138 (N_22138,N_19821,N_19670);
xor U22139 (N_22139,N_20057,N_20707);
nor U22140 (N_22140,N_20257,N_20533);
nor U22141 (N_22141,N_20857,N_20213);
nand U22142 (N_22142,N_20381,N_20241);
or U22143 (N_22143,N_19670,N_20844);
or U22144 (N_22144,N_20996,N_20552);
nand U22145 (N_22145,N_19667,N_20956);
xnor U22146 (N_22146,N_20010,N_20144);
xnor U22147 (N_22147,N_20725,N_20672);
nand U22148 (N_22148,N_20006,N_20430);
nand U22149 (N_22149,N_20705,N_20521);
or U22150 (N_22150,N_19785,N_19539);
nand U22151 (N_22151,N_20564,N_20349);
nor U22152 (N_22152,N_20617,N_20990);
and U22153 (N_22153,N_20795,N_20484);
xnor U22154 (N_22154,N_20492,N_20284);
or U22155 (N_22155,N_20078,N_20802);
and U22156 (N_22156,N_20362,N_20104);
xnor U22157 (N_22157,N_19741,N_19890);
xnor U22158 (N_22158,N_20727,N_20270);
nand U22159 (N_22159,N_20780,N_20291);
nand U22160 (N_22160,N_19657,N_20116);
nand U22161 (N_22161,N_19551,N_19960);
nand U22162 (N_22162,N_20155,N_20123);
nor U22163 (N_22163,N_20465,N_20669);
or U22164 (N_22164,N_20286,N_20987);
and U22165 (N_22165,N_20782,N_19668);
or U22166 (N_22166,N_20408,N_20644);
and U22167 (N_22167,N_20840,N_20422);
xnor U22168 (N_22168,N_20404,N_19800);
nand U22169 (N_22169,N_19664,N_20122);
or U22170 (N_22170,N_20230,N_20979);
or U22171 (N_22171,N_19850,N_20740);
or U22172 (N_22172,N_20128,N_20412);
nand U22173 (N_22173,N_19969,N_19926);
nand U22174 (N_22174,N_19549,N_19867);
nor U22175 (N_22175,N_20381,N_20270);
nand U22176 (N_22176,N_20137,N_20334);
and U22177 (N_22177,N_20552,N_20433);
and U22178 (N_22178,N_19632,N_19979);
or U22179 (N_22179,N_20464,N_19929);
nand U22180 (N_22180,N_20598,N_20714);
or U22181 (N_22181,N_20183,N_20691);
nand U22182 (N_22182,N_20950,N_20889);
and U22183 (N_22183,N_19888,N_20569);
xor U22184 (N_22184,N_19703,N_20816);
and U22185 (N_22185,N_19839,N_20027);
and U22186 (N_22186,N_20481,N_20996);
and U22187 (N_22187,N_19757,N_20567);
nor U22188 (N_22188,N_19814,N_19508);
xor U22189 (N_22189,N_19748,N_20593);
or U22190 (N_22190,N_20051,N_20019);
or U22191 (N_22191,N_19994,N_20368);
and U22192 (N_22192,N_19813,N_19561);
nor U22193 (N_22193,N_20846,N_19542);
xnor U22194 (N_22194,N_20908,N_20723);
xor U22195 (N_22195,N_20661,N_20807);
and U22196 (N_22196,N_20563,N_20717);
nor U22197 (N_22197,N_20362,N_20703);
nand U22198 (N_22198,N_20885,N_20554);
xor U22199 (N_22199,N_20194,N_20123);
xor U22200 (N_22200,N_20605,N_20997);
nand U22201 (N_22201,N_19702,N_19813);
nor U22202 (N_22202,N_19729,N_20096);
xnor U22203 (N_22203,N_19804,N_19591);
or U22204 (N_22204,N_20120,N_20037);
nand U22205 (N_22205,N_20305,N_20506);
nand U22206 (N_22206,N_19662,N_20670);
and U22207 (N_22207,N_20694,N_20043);
and U22208 (N_22208,N_20576,N_20607);
nand U22209 (N_22209,N_20651,N_20880);
and U22210 (N_22210,N_19832,N_20620);
and U22211 (N_22211,N_20244,N_19861);
xor U22212 (N_22212,N_20167,N_19649);
or U22213 (N_22213,N_20588,N_19632);
and U22214 (N_22214,N_20120,N_20036);
or U22215 (N_22215,N_20706,N_20744);
xnor U22216 (N_22216,N_20197,N_19827);
nand U22217 (N_22217,N_20154,N_20892);
or U22218 (N_22218,N_19947,N_19827);
nor U22219 (N_22219,N_20904,N_20963);
and U22220 (N_22220,N_20248,N_20842);
or U22221 (N_22221,N_19774,N_20292);
nor U22222 (N_22222,N_19722,N_19650);
nand U22223 (N_22223,N_20045,N_20262);
xor U22224 (N_22224,N_19572,N_20348);
nor U22225 (N_22225,N_20976,N_20239);
nand U22226 (N_22226,N_19610,N_20106);
xor U22227 (N_22227,N_19844,N_19684);
or U22228 (N_22228,N_20253,N_20781);
nand U22229 (N_22229,N_19774,N_20681);
or U22230 (N_22230,N_20526,N_20943);
xor U22231 (N_22231,N_19924,N_20458);
and U22232 (N_22232,N_19568,N_20741);
nor U22233 (N_22233,N_20671,N_20605);
nand U22234 (N_22234,N_20657,N_20170);
nand U22235 (N_22235,N_19735,N_19736);
nor U22236 (N_22236,N_19579,N_19739);
nor U22237 (N_22237,N_19528,N_20768);
nor U22238 (N_22238,N_19677,N_20569);
xor U22239 (N_22239,N_20684,N_19541);
nand U22240 (N_22240,N_20510,N_20823);
xor U22241 (N_22241,N_20726,N_20264);
nand U22242 (N_22242,N_20476,N_20302);
nor U22243 (N_22243,N_20834,N_20979);
or U22244 (N_22244,N_20724,N_19692);
nand U22245 (N_22245,N_20231,N_20457);
and U22246 (N_22246,N_20418,N_20819);
and U22247 (N_22247,N_20329,N_20995);
xor U22248 (N_22248,N_19665,N_20132);
or U22249 (N_22249,N_20940,N_19536);
xor U22250 (N_22250,N_19931,N_19795);
nand U22251 (N_22251,N_19737,N_19983);
nand U22252 (N_22252,N_20763,N_20907);
nor U22253 (N_22253,N_20702,N_20168);
nand U22254 (N_22254,N_20620,N_20708);
nor U22255 (N_22255,N_20681,N_20795);
xor U22256 (N_22256,N_19705,N_20790);
or U22257 (N_22257,N_20765,N_19586);
and U22258 (N_22258,N_20208,N_19723);
and U22259 (N_22259,N_20391,N_20988);
nor U22260 (N_22260,N_19876,N_20377);
nor U22261 (N_22261,N_20108,N_20151);
nand U22262 (N_22262,N_20019,N_20269);
xnor U22263 (N_22263,N_19780,N_20165);
or U22264 (N_22264,N_20202,N_20433);
or U22265 (N_22265,N_19545,N_20398);
or U22266 (N_22266,N_19797,N_20052);
xor U22267 (N_22267,N_20739,N_20969);
xnor U22268 (N_22268,N_20636,N_20334);
or U22269 (N_22269,N_20418,N_20643);
xnor U22270 (N_22270,N_19817,N_20404);
or U22271 (N_22271,N_20444,N_20078);
nand U22272 (N_22272,N_20006,N_20136);
xnor U22273 (N_22273,N_19615,N_20239);
and U22274 (N_22274,N_20571,N_19592);
xnor U22275 (N_22275,N_20825,N_20852);
or U22276 (N_22276,N_19863,N_20802);
and U22277 (N_22277,N_20895,N_20314);
and U22278 (N_22278,N_19952,N_20328);
or U22279 (N_22279,N_19580,N_19735);
and U22280 (N_22280,N_19603,N_20902);
nor U22281 (N_22281,N_19814,N_20567);
nor U22282 (N_22282,N_20380,N_20887);
or U22283 (N_22283,N_19594,N_19506);
or U22284 (N_22284,N_20591,N_20053);
or U22285 (N_22285,N_19906,N_19820);
xor U22286 (N_22286,N_19969,N_19524);
nand U22287 (N_22287,N_20490,N_20459);
or U22288 (N_22288,N_20108,N_20239);
nand U22289 (N_22289,N_20736,N_19888);
nor U22290 (N_22290,N_19783,N_20466);
nor U22291 (N_22291,N_20912,N_20764);
nor U22292 (N_22292,N_20792,N_20430);
or U22293 (N_22293,N_20926,N_20244);
nand U22294 (N_22294,N_19954,N_20748);
and U22295 (N_22295,N_20523,N_19663);
and U22296 (N_22296,N_20193,N_19541);
nor U22297 (N_22297,N_20968,N_19894);
nand U22298 (N_22298,N_20489,N_19988);
xor U22299 (N_22299,N_20149,N_20646);
nand U22300 (N_22300,N_20045,N_20603);
or U22301 (N_22301,N_20088,N_20918);
nand U22302 (N_22302,N_20754,N_20284);
nor U22303 (N_22303,N_20831,N_19839);
and U22304 (N_22304,N_20789,N_20547);
nand U22305 (N_22305,N_20892,N_19518);
or U22306 (N_22306,N_20273,N_20348);
nand U22307 (N_22307,N_19609,N_19625);
and U22308 (N_22308,N_19982,N_20832);
or U22309 (N_22309,N_19671,N_19919);
or U22310 (N_22310,N_20605,N_19587);
nor U22311 (N_22311,N_19638,N_19859);
nor U22312 (N_22312,N_20817,N_20947);
nor U22313 (N_22313,N_19731,N_20286);
nand U22314 (N_22314,N_20854,N_19913);
nor U22315 (N_22315,N_19800,N_20618);
or U22316 (N_22316,N_19802,N_19734);
and U22317 (N_22317,N_19700,N_19905);
nor U22318 (N_22318,N_19718,N_19716);
xor U22319 (N_22319,N_20008,N_19572);
and U22320 (N_22320,N_20818,N_20809);
and U22321 (N_22321,N_19597,N_20442);
nand U22322 (N_22322,N_20191,N_20929);
nor U22323 (N_22323,N_19715,N_20412);
nand U22324 (N_22324,N_19938,N_19724);
or U22325 (N_22325,N_20229,N_20069);
or U22326 (N_22326,N_20743,N_20156);
nand U22327 (N_22327,N_19900,N_20385);
or U22328 (N_22328,N_20750,N_20096);
or U22329 (N_22329,N_19843,N_19951);
or U22330 (N_22330,N_20324,N_20546);
and U22331 (N_22331,N_20406,N_19887);
nor U22332 (N_22332,N_20454,N_20892);
nor U22333 (N_22333,N_20016,N_20845);
nor U22334 (N_22334,N_20377,N_19969);
and U22335 (N_22335,N_20604,N_19705);
nand U22336 (N_22336,N_20394,N_20407);
or U22337 (N_22337,N_20350,N_20674);
or U22338 (N_22338,N_19978,N_19938);
or U22339 (N_22339,N_20179,N_20526);
and U22340 (N_22340,N_20508,N_20339);
or U22341 (N_22341,N_20950,N_20691);
nand U22342 (N_22342,N_20395,N_20567);
nor U22343 (N_22343,N_20986,N_19751);
xnor U22344 (N_22344,N_19894,N_20454);
nor U22345 (N_22345,N_20082,N_19927);
xnor U22346 (N_22346,N_19806,N_20695);
xnor U22347 (N_22347,N_20521,N_20281);
or U22348 (N_22348,N_19701,N_20242);
nand U22349 (N_22349,N_20623,N_19553);
nand U22350 (N_22350,N_19588,N_20411);
and U22351 (N_22351,N_20873,N_19996);
nor U22352 (N_22352,N_19975,N_20333);
or U22353 (N_22353,N_20482,N_19714);
or U22354 (N_22354,N_20093,N_19569);
or U22355 (N_22355,N_20537,N_20249);
and U22356 (N_22356,N_19583,N_20764);
or U22357 (N_22357,N_20259,N_19744);
nor U22358 (N_22358,N_19582,N_20986);
and U22359 (N_22359,N_19904,N_20278);
or U22360 (N_22360,N_19552,N_19982);
or U22361 (N_22361,N_20909,N_20587);
nor U22362 (N_22362,N_19758,N_20919);
nor U22363 (N_22363,N_20853,N_20695);
xor U22364 (N_22364,N_20797,N_20245);
or U22365 (N_22365,N_20849,N_19521);
or U22366 (N_22366,N_19618,N_19525);
or U22367 (N_22367,N_20130,N_20246);
xnor U22368 (N_22368,N_20826,N_19914);
xnor U22369 (N_22369,N_20484,N_19684);
or U22370 (N_22370,N_20948,N_20679);
and U22371 (N_22371,N_20969,N_19659);
or U22372 (N_22372,N_19843,N_19562);
or U22373 (N_22373,N_20314,N_20237);
nor U22374 (N_22374,N_19838,N_20455);
nand U22375 (N_22375,N_20095,N_20914);
or U22376 (N_22376,N_20937,N_19647);
nand U22377 (N_22377,N_20499,N_20937);
nor U22378 (N_22378,N_19528,N_20159);
nor U22379 (N_22379,N_20786,N_19639);
nand U22380 (N_22380,N_20593,N_20063);
nand U22381 (N_22381,N_19705,N_20641);
or U22382 (N_22382,N_20964,N_19779);
or U22383 (N_22383,N_20695,N_20220);
nor U22384 (N_22384,N_20057,N_20007);
nand U22385 (N_22385,N_20495,N_20742);
and U22386 (N_22386,N_19826,N_20443);
and U22387 (N_22387,N_20196,N_20524);
nor U22388 (N_22388,N_19716,N_20891);
and U22389 (N_22389,N_20402,N_19558);
nand U22390 (N_22390,N_20927,N_20908);
xnor U22391 (N_22391,N_20381,N_20477);
xnor U22392 (N_22392,N_19997,N_20578);
nand U22393 (N_22393,N_19632,N_19520);
xnor U22394 (N_22394,N_20603,N_20756);
nor U22395 (N_22395,N_20482,N_20405);
nand U22396 (N_22396,N_19701,N_19501);
nor U22397 (N_22397,N_20923,N_20498);
nand U22398 (N_22398,N_19889,N_19791);
xnor U22399 (N_22399,N_20579,N_20471);
and U22400 (N_22400,N_20219,N_20380);
nand U22401 (N_22401,N_20783,N_19502);
or U22402 (N_22402,N_20335,N_20302);
nor U22403 (N_22403,N_20028,N_20218);
nor U22404 (N_22404,N_19982,N_19855);
nor U22405 (N_22405,N_20541,N_20871);
or U22406 (N_22406,N_20424,N_20741);
nand U22407 (N_22407,N_20547,N_20396);
xnor U22408 (N_22408,N_19818,N_19656);
xor U22409 (N_22409,N_20841,N_20618);
or U22410 (N_22410,N_19744,N_19730);
nor U22411 (N_22411,N_20710,N_19648);
xor U22412 (N_22412,N_20608,N_20644);
nand U22413 (N_22413,N_19702,N_19930);
or U22414 (N_22414,N_20652,N_20316);
and U22415 (N_22415,N_20593,N_19527);
nor U22416 (N_22416,N_20925,N_20732);
and U22417 (N_22417,N_20230,N_19793);
and U22418 (N_22418,N_20518,N_19657);
nand U22419 (N_22419,N_20366,N_20564);
and U22420 (N_22420,N_19531,N_20161);
nor U22421 (N_22421,N_19844,N_19601);
and U22422 (N_22422,N_19973,N_20097);
nor U22423 (N_22423,N_19759,N_19511);
xor U22424 (N_22424,N_20499,N_19630);
xor U22425 (N_22425,N_19756,N_20374);
xor U22426 (N_22426,N_19892,N_20746);
nand U22427 (N_22427,N_20199,N_20676);
and U22428 (N_22428,N_20507,N_19628);
nand U22429 (N_22429,N_19516,N_20562);
nand U22430 (N_22430,N_20745,N_20790);
nor U22431 (N_22431,N_20325,N_20995);
xor U22432 (N_22432,N_20114,N_19757);
nand U22433 (N_22433,N_19863,N_20609);
nor U22434 (N_22434,N_20648,N_19504);
nand U22435 (N_22435,N_20902,N_19916);
xnor U22436 (N_22436,N_20801,N_20243);
nand U22437 (N_22437,N_20716,N_20896);
and U22438 (N_22438,N_20580,N_20139);
and U22439 (N_22439,N_20829,N_20562);
or U22440 (N_22440,N_20962,N_20710);
and U22441 (N_22441,N_19532,N_20973);
xnor U22442 (N_22442,N_20085,N_19960);
xnor U22443 (N_22443,N_20709,N_19740);
xor U22444 (N_22444,N_19868,N_20143);
xnor U22445 (N_22445,N_19769,N_20337);
nand U22446 (N_22446,N_20323,N_20820);
nor U22447 (N_22447,N_20189,N_19797);
nor U22448 (N_22448,N_20432,N_20101);
or U22449 (N_22449,N_20845,N_19751);
xor U22450 (N_22450,N_20083,N_20130);
nor U22451 (N_22451,N_20243,N_20514);
and U22452 (N_22452,N_20517,N_20010);
nor U22453 (N_22453,N_20426,N_20573);
nor U22454 (N_22454,N_20070,N_19720);
xor U22455 (N_22455,N_20967,N_20036);
or U22456 (N_22456,N_20941,N_19587);
nand U22457 (N_22457,N_20286,N_20526);
nor U22458 (N_22458,N_20905,N_20043);
or U22459 (N_22459,N_20012,N_20897);
xor U22460 (N_22460,N_19990,N_19605);
nand U22461 (N_22461,N_20304,N_20733);
or U22462 (N_22462,N_20826,N_20957);
xnor U22463 (N_22463,N_20615,N_20513);
nor U22464 (N_22464,N_19823,N_20084);
nand U22465 (N_22465,N_19736,N_19711);
nor U22466 (N_22466,N_20917,N_19801);
or U22467 (N_22467,N_20606,N_19517);
xor U22468 (N_22468,N_19760,N_20658);
and U22469 (N_22469,N_20513,N_19778);
or U22470 (N_22470,N_20971,N_19620);
nor U22471 (N_22471,N_20785,N_19722);
nor U22472 (N_22472,N_19547,N_20718);
nand U22473 (N_22473,N_20256,N_20747);
and U22474 (N_22474,N_20677,N_19603);
nor U22475 (N_22475,N_20993,N_20435);
and U22476 (N_22476,N_19804,N_20762);
nor U22477 (N_22477,N_20832,N_20823);
or U22478 (N_22478,N_20319,N_19815);
nand U22479 (N_22479,N_19639,N_19662);
nand U22480 (N_22480,N_20534,N_19790);
xor U22481 (N_22481,N_19886,N_20800);
and U22482 (N_22482,N_19690,N_20101);
nand U22483 (N_22483,N_20613,N_19889);
nand U22484 (N_22484,N_20187,N_20938);
nand U22485 (N_22485,N_20067,N_19561);
xor U22486 (N_22486,N_20722,N_19603);
nor U22487 (N_22487,N_20373,N_20769);
and U22488 (N_22488,N_20587,N_19838);
or U22489 (N_22489,N_20224,N_20756);
or U22490 (N_22490,N_20995,N_19900);
xnor U22491 (N_22491,N_20761,N_20562);
nand U22492 (N_22492,N_20964,N_20857);
or U22493 (N_22493,N_20086,N_19842);
nand U22494 (N_22494,N_20465,N_20623);
and U22495 (N_22495,N_20512,N_20454);
nand U22496 (N_22496,N_20183,N_19914);
nand U22497 (N_22497,N_20361,N_20688);
or U22498 (N_22498,N_19506,N_19640);
xnor U22499 (N_22499,N_20913,N_20972);
nor U22500 (N_22500,N_21513,N_22393);
nor U22501 (N_22501,N_21181,N_21047);
and U22502 (N_22502,N_21432,N_21775);
nand U22503 (N_22503,N_22174,N_21711);
nand U22504 (N_22504,N_22351,N_22445);
or U22505 (N_22505,N_21304,N_21155);
nor U22506 (N_22506,N_22453,N_21769);
xor U22507 (N_22507,N_22415,N_22372);
nor U22508 (N_22508,N_21739,N_22151);
nor U22509 (N_22509,N_22127,N_21721);
nand U22510 (N_22510,N_22286,N_21274);
nand U22511 (N_22511,N_22167,N_21046);
or U22512 (N_22512,N_21367,N_22446);
nor U22513 (N_22513,N_21344,N_22325);
and U22514 (N_22514,N_21868,N_21714);
nand U22515 (N_22515,N_21616,N_21555);
nor U22516 (N_22516,N_21877,N_21416);
xnor U22517 (N_22517,N_21393,N_22479);
nand U22518 (N_22518,N_21875,N_21031);
or U22519 (N_22519,N_22419,N_22238);
nand U22520 (N_22520,N_21341,N_22305);
nor U22521 (N_22521,N_22191,N_22219);
nor U22522 (N_22522,N_21381,N_21850);
or U22523 (N_22523,N_22170,N_21576);
nand U22524 (N_22524,N_21136,N_21414);
xor U22525 (N_22525,N_21243,N_22413);
nand U22526 (N_22526,N_21614,N_21256);
nand U22527 (N_22527,N_22438,N_21268);
xnor U22528 (N_22528,N_22381,N_21949);
nand U22529 (N_22529,N_21002,N_21984);
nand U22530 (N_22530,N_21279,N_21222);
or U22531 (N_22531,N_22007,N_21434);
nor U22532 (N_22532,N_22148,N_21538);
nor U22533 (N_22533,N_22009,N_21307);
xnor U22534 (N_22534,N_21262,N_21605);
or U22535 (N_22535,N_21626,N_22296);
xor U22536 (N_22536,N_21643,N_21273);
or U22537 (N_22537,N_21910,N_21597);
xor U22538 (N_22538,N_21904,N_21437);
xnor U22539 (N_22539,N_21378,N_22205);
xnor U22540 (N_22540,N_22457,N_21923);
nand U22541 (N_22541,N_21417,N_21411);
xnor U22542 (N_22542,N_21718,N_22214);
nand U22543 (N_22543,N_21599,N_21329);
or U22544 (N_22544,N_22355,N_22134);
xor U22545 (N_22545,N_22078,N_21809);
or U22546 (N_22546,N_21685,N_21701);
xnor U22547 (N_22547,N_22137,N_22300);
nand U22548 (N_22548,N_21692,N_22276);
nor U22549 (N_22549,N_21717,N_21288);
nor U22550 (N_22550,N_21883,N_21921);
nor U22551 (N_22551,N_21937,N_21006);
nor U22552 (N_22552,N_21254,N_21255);
or U22553 (N_22553,N_21588,N_21052);
and U22554 (N_22554,N_22474,N_21746);
nor U22555 (N_22555,N_21996,N_22048);
and U22556 (N_22556,N_22408,N_22266);
and U22557 (N_22557,N_21025,N_21713);
and U22558 (N_22558,N_22357,N_21783);
nand U22559 (N_22559,N_21791,N_21546);
and U22560 (N_22560,N_21815,N_21287);
or U22561 (N_22561,N_21516,N_21798);
and U22562 (N_22562,N_22384,N_21527);
nand U22563 (N_22563,N_22039,N_21302);
and U22564 (N_22564,N_21689,N_22224);
and U22565 (N_22565,N_21011,N_21567);
or U22566 (N_22566,N_21821,N_21660);
nand U22567 (N_22567,N_22083,N_21976);
nand U22568 (N_22568,N_21228,N_22141);
xor U22569 (N_22569,N_21298,N_22118);
nor U22570 (N_22570,N_21270,N_21529);
or U22571 (N_22571,N_22467,N_21296);
and U22572 (N_22572,N_21966,N_21340);
xnor U22573 (N_22573,N_21332,N_21762);
nor U22574 (N_22574,N_21690,N_21051);
or U22575 (N_22575,N_21878,N_22179);
and U22576 (N_22576,N_22023,N_22129);
nand U22577 (N_22577,N_21184,N_22133);
or U22578 (N_22578,N_22051,N_22189);
xnor U22579 (N_22579,N_21142,N_21606);
nor U22580 (N_22580,N_21009,N_21370);
nand U22581 (N_22581,N_22405,N_21085);
and U22582 (N_22582,N_21869,N_21029);
and U22583 (N_22583,N_22335,N_21100);
and U22584 (N_22584,N_22016,N_21200);
nor U22585 (N_22585,N_21654,N_21147);
and U22586 (N_22586,N_21246,N_21895);
and U22587 (N_22587,N_21148,N_21125);
nand U22588 (N_22588,N_22387,N_21645);
and U22589 (N_22589,N_22215,N_21280);
or U22590 (N_22590,N_21568,N_22264);
nor U22591 (N_22591,N_21502,N_22211);
xor U22592 (N_22592,N_21013,N_21640);
nor U22593 (N_22593,N_21559,N_21366);
nand U22594 (N_22594,N_21382,N_21334);
or U22595 (N_22595,N_21446,N_22244);
nor U22596 (N_22596,N_22213,N_21102);
nor U22597 (N_22597,N_21308,N_22182);
and U22598 (N_22598,N_21731,N_22253);
nand U22599 (N_22599,N_22431,N_22280);
nor U22600 (N_22600,N_21540,N_22478);
and U22601 (N_22601,N_21350,N_22200);
nor U22602 (N_22602,N_22124,N_21232);
nor U22603 (N_22603,N_22242,N_21498);
nor U22604 (N_22604,N_21623,N_22043);
and U22605 (N_22605,N_21524,N_21755);
xnor U22606 (N_22606,N_21541,N_22397);
nand U22607 (N_22607,N_21741,N_22089);
or U22608 (N_22608,N_22092,N_21187);
or U22609 (N_22609,N_22435,N_22282);
xnor U22610 (N_22610,N_22140,N_21004);
or U22611 (N_22611,N_21892,N_22365);
and U22612 (N_22612,N_22011,N_22473);
and U22613 (N_22613,N_22323,N_21466);
xnor U22614 (N_22614,N_21406,N_21707);
or U22615 (N_22615,N_22394,N_22334);
or U22616 (N_22616,N_21844,N_22185);
nand U22617 (N_22617,N_21680,N_21832);
nand U22618 (N_22618,N_21140,N_21677);
xnor U22619 (N_22619,N_21508,N_21257);
xnor U22620 (N_22620,N_21843,N_22268);
xor U22621 (N_22621,N_22115,N_22454);
nand U22622 (N_22622,N_21276,N_21328);
and U22623 (N_22623,N_21777,N_21045);
xor U22624 (N_22624,N_21186,N_22256);
or U22625 (N_22625,N_21321,N_21807);
nor U22626 (N_22626,N_21804,N_22120);
and U22627 (N_22627,N_21915,N_22366);
nor U22628 (N_22628,N_21730,N_21986);
xor U22629 (N_22629,N_21343,N_21687);
or U22630 (N_22630,N_21259,N_22196);
and U22631 (N_22631,N_21162,N_21905);
or U22632 (N_22632,N_22038,N_21973);
nor U22633 (N_22633,N_21035,N_21441);
nor U22634 (N_22634,N_21969,N_21670);
xnor U22635 (N_22635,N_21722,N_21021);
and U22636 (N_22636,N_21445,N_21562);
nor U22637 (N_22637,N_21152,N_21453);
xnor U22638 (N_22638,N_22345,N_22055);
nor U22639 (N_22639,N_22019,N_21706);
xor U22640 (N_22640,N_21801,N_21790);
or U22641 (N_22641,N_21023,N_21865);
and U22642 (N_22642,N_21612,N_21547);
nor U22643 (N_22643,N_21129,N_21115);
xnor U22644 (N_22644,N_22432,N_22310);
or U22645 (N_22645,N_21324,N_22112);
nand U22646 (N_22646,N_22373,N_21153);
nand U22647 (N_22647,N_21475,N_22443);
nor U22648 (N_22648,N_21595,N_21965);
and U22649 (N_22649,N_21728,N_21585);
xnor U22650 (N_22650,N_21556,N_21942);
and U22651 (N_22651,N_22192,N_22107);
xnor U22652 (N_22652,N_22030,N_21063);
and U22653 (N_22653,N_21784,N_21374);
xor U22654 (N_22654,N_21693,N_22402);
nand U22655 (N_22655,N_21512,N_22220);
and U22656 (N_22656,N_21827,N_21533);
nand U22657 (N_22657,N_21579,N_21286);
and U22658 (N_22658,N_21771,N_22342);
nand U22659 (N_22659,N_22207,N_21097);
nor U22660 (N_22660,N_21931,N_21419);
xnor U22661 (N_22661,N_22150,N_22024);
nand U22662 (N_22662,N_21027,N_22404);
nor U22663 (N_22663,N_21300,N_22097);
nand U22664 (N_22664,N_21096,N_21899);
or U22665 (N_22665,N_21566,N_21483);
xnor U22666 (N_22666,N_21647,N_21413);
and U22667 (N_22667,N_21346,N_22370);
and U22668 (N_22668,N_21379,N_21348);
nand U22669 (N_22669,N_22401,N_22295);
and U22670 (N_22670,N_22159,N_22113);
nor U22671 (N_22671,N_21083,N_21810);
or U22672 (N_22672,N_21299,N_22313);
xor U22673 (N_22673,N_21918,N_21471);
nor U22674 (N_22674,N_21362,N_21008);
nand U22675 (N_22675,N_21825,N_22004);
xor U22676 (N_22676,N_22360,N_21111);
nand U22677 (N_22677,N_22066,N_21565);
nand U22678 (N_22678,N_22226,N_21294);
and U22679 (N_22679,N_22060,N_21853);
xnor U22680 (N_22680,N_22262,N_21487);
nor U22681 (N_22681,N_21174,N_21210);
nand U22682 (N_22682,N_22052,N_21390);
and U22683 (N_22683,N_21700,N_21916);
and U22684 (N_22684,N_21201,N_21743);
and U22685 (N_22685,N_21613,N_22314);
nand U22686 (N_22686,N_22161,N_21226);
xnor U22687 (N_22687,N_21688,N_21872);
nor U22688 (N_22688,N_21668,N_22385);
or U22689 (N_22689,N_21550,N_22143);
or U22690 (N_22690,N_22488,N_22424);
xnor U22691 (N_22691,N_21552,N_21506);
or U22692 (N_22692,N_21528,N_22079);
nand U22693 (N_22693,N_22311,N_21363);
xor U22694 (N_22694,N_21824,N_21767);
nand U22695 (N_22695,N_21816,N_22114);
and U22696 (N_22696,N_21238,N_21554);
or U22697 (N_22697,N_21805,N_21526);
nor U22698 (N_22698,N_21001,N_21387);
nand U22699 (N_22699,N_21042,N_21056);
or U22700 (N_22700,N_21456,N_21593);
xor U22701 (N_22701,N_22498,N_21799);
nand U22702 (N_22702,N_21808,N_22096);
nor U22703 (N_22703,N_22091,N_21880);
xnor U22704 (N_22704,N_22425,N_22106);
xnor U22705 (N_22705,N_22270,N_21972);
or U22706 (N_22706,N_22315,N_22495);
or U22707 (N_22707,N_21738,N_21846);
xor U22708 (N_22708,N_21427,N_22447);
xor U22709 (N_22709,N_21607,N_21830);
and U22710 (N_22710,N_22077,N_21269);
and U22711 (N_22711,N_22003,N_21520);
nor U22712 (N_22712,N_21069,N_21402);
xnor U22713 (N_22713,N_22202,N_21463);
xor U22714 (N_22714,N_21968,N_22391);
or U22715 (N_22715,N_21563,N_21514);
xor U22716 (N_22716,N_21442,N_21386);
nor U22717 (N_22717,N_21164,N_21503);
and U22718 (N_22718,N_21620,N_21289);
xor U22719 (N_22719,N_21311,N_21681);
xor U22720 (N_22720,N_21058,N_22010);
nor U22721 (N_22721,N_21855,N_22171);
nor U22722 (N_22722,N_22322,N_22257);
nand U22723 (N_22723,N_21234,N_22255);
or U22724 (N_22724,N_21231,N_21320);
xnor U22725 (N_22725,N_21837,N_21829);
nand U22726 (N_22726,N_21150,N_22483);
nor U22727 (N_22727,N_21823,N_21032);
and U22728 (N_22728,N_22285,N_21325);
nor U22729 (N_22729,N_21473,N_22426);
nor U22730 (N_22730,N_21209,N_21686);
or U22731 (N_22731,N_21763,N_21795);
and U22732 (N_22732,N_22098,N_21537);
xor U22733 (N_22733,N_22429,N_22153);
nor U22734 (N_22734,N_21486,N_22411);
nor U22735 (N_22735,N_22061,N_21397);
nor U22736 (N_22736,N_21128,N_21703);
nor U22737 (N_22737,N_21055,N_21188);
xor U22738 (N_22738,N_21663,N_22260);
nor U22739 (N_22739,N_21179,N_21342);
or U22740 (N_22740,N_22176,N_21927);
nor U22741 (N_22741,N_21138,N_21208);
xnor U22742 (N_22742,N_21636,N_22409);
xor U22743 (N_22743,N_21309,N_21926);
xor U22744 (N_22744,N_21998,N_22070);
and U22745 (N_22745,N_21662,N_22427);
nor U22746 (N_22746,N_22076,N_21444);
nor U22747 (N_22747,N_21871,N_21664);
xor U22748 (N_22748,N_21478,N_21589);
xor U22749 (N_22749,N_22216,N_21947);
xnor U22750 (N_22750,N_21283,N_21952);
and U22751 (N_22751,N_21840,N_21195);
nand U22752 (N_22752,N_22470,N_22247);
and U22753 (N_22753,N_21160,N_21617);
nor U22754 (N_22754,N_22309,N_22053);
xnor U22755 (N_22755,N_22054,N_21462);
nor U22756 (N_22756,N_22317,N_21678);
or U22757 (N_22757,N_21999,N_21183);
xnor U22758 (N_22758,N_21291,N_22085);
nand U22759 (N_22759,N_22390,N_22382);
and U22760 (N_22760,N_22469,N_22290);
or U22761 (N_22761,N_21053,N_22418);
nor U22762 (N_22762,N_22316,N_22031);
and U22763 (N_22763,N_21674,N_21776);
or U22764 (N_22764,N_22020,N_21098);
and U22765 (N_22765,N_21099,N_21591);
nor U22766 (N_22766,N_21696,N_22493);
nor U22767 (N_22767,N_22389,N_22341);
or U22768 (N_22768,N_21803,N_22364);
and U22769 (N_22769,N_21353,N_21876);
nand U22770 (N_22770,N_21322,N_21224);
and U22771 (N_22771,N_21260,N_21271);
or U22772 (N_22772,N_21395,N_22304);
xnor U22773 (N_22773,N_21683,N_21610);
nor U22774 (N_22774,N_22086,N_22459);
or U22775 (N_22775,N_21197,N_21974);
nor U22776 (N_22776,N_21492,N_21295);
xnor U22777 (N_22777,N_21542,N_22223);
and U22778 (N_22778,N_21770,N_21223);
nor U22779 (N_22779,N_21994,N_21331);
or U22780 (N_22780,N_21460,N_21505);
nor U22781 (N_22781,N_22146,N_22281);
xor U22782 (N_22782,N_22034,N_22386);
xnor U22783 (N_22783,N_22361,N_22040);
nand U22784 (N_22784,N_21326,N_22232);
nand U22785 (N_22785,N_22492,N_21034);
nor U22786 (N_22786,N_21146,N_21971);
nand U22787 (N_22787,N_21922,N_21472);
nor U22788 (N_22788,N_21394,N_21561);
or U22789 (N_22789,N_22354,N_21190);
xor U22790 (N_22790,N_21944,N_21422);
or U22791 (N_22791,N_21145,N_22486);
nand U22792 (N_22792,N_21191,N_22029);
or U22793 (N_22793,N_22117,N_22121);
xor U22794 (N_22794,N_21742,N_22152);
xnor U22795 (N_22795,N_21796,N_22297);
or U22796 (N_22796,N_21245,N_22221);
xor U22797 (N_22797,N_22198,N_21578);
or U22798 (N_22798,N_22450,N_21244);
or U22799 (N_22799,N_21773,N_21656);
and U22800 (N_22800,N_21319,N_22273);
nor U22801 (N_22801,N_21392,N_21793);
and U22802 (N_22802,N_22059,N_21089);
nor U22803 (N_22803,N_21977,N_21292);
and U22804 (N_22804,N_21253,N_22108);
nor U22805 (N_22805,N_21858,N_21980);
xor U22806 (N_22806,N_22484,N_21715);
nand U22807 (N_22807,N_22465,N_21504);
and U22808 (N_22808,N_21932,N_21822);
nor U22809 (N_22809,N_22058,N_22021);
nor U22810 (N_22810,N_21401,N_21560);
nand U22811 (N_22811,N_21836,N_21040);
and U22812 (N_22812,N_21806,N_22116);
nor U22813 (N_22813,N_22050,N_22173);
nor U22814 (N_22814,N_21780,N_21104);
or U22815 (N_22815,N_22230,N_21928);
and U22816 (N_22816,N_21519,N_21093);
xnor U22817 (N_22817,N_22452,N_21211);
or U22818 (N_22818,N_22487,N_22163);
xnor U22819 (N_22819,N_21819,N_21082);
nor U22820 (N_22820,N_22455,N_21007);
and U22821 (N_22821,N_21043,N_21615);
nand U22822 (N_22822,N_21699,N_21240);
xor U22823 (N_22823,N_21571,N_22275);
or U22824 (N_22824,N_21264,N_21684);
nand U22825 (N_22825,N_21631,N_21494);
xor U22826 (N_22826,N_21318,N_21124);
nor U22827 (N_22827,N_21134,N_21400);
or U22828 (N_22828,N_21206,N_21316);
nor U22829 (N_22829,N_21787,N_21592);
or U22830 (N_22830,N_22125,N_22002);
or U22831 (N_22831,N_22269,N_21365);
nor U22832 (N_22832,N_21539,N_21048);
or U22833 (N_22833,N_22331,N_21433);
or U22834 (N_22834,N_21691,N_21551);
and U22835 (N_22835,N_21768,N_21022);
and U22836 (N_22836,N_22068,N_22318);
nor U22837 (N_22837,N_22158,N_22037);
nand U22838 (N_22838,N_22292,N_21726);
and U22839 (N_22839,N_22128,N_21193);
and U22840 (N_22840,N_21018,N_22201);
xor U22841 (N_22841,N_22101,N_21758);
or U22842 (N_22842,N_21204,N_21587);
or U22843 (N_22843,N_22186,N_22245);
and U22844 (N_22844,N_22376,N_21424);
and U22845 (N_22845,N_22155,N_21648);
nor U22846 (N_22846,N_22087,N_21667);
nor U22847 (N_22847,N_21629,N_21525);
xor U22848 (N_22848,N_21313,N_22344);
and U22849 (N_22849,N_21092,N_22476);
nand U22850 (N_22850,N_22001,N_21112);
and U22851 (N_22851,N_22458,N_21451);
or U22852 (N_22852,N_21229,N_21012);
or U22853 (N_22853,N_22056,N_21515);
nor U22854 (N_22854,N_21194,N_22111);
xor U22855 (N_22855,N_22267,N_21133);
and U22856 (N_22856,N_22379,N_21026);
xnor U22857 (N_22857,N_22168,N_21549);
xnor U22858 (N_22858,N_22042,N_21061);
nor U22859 (N_22859,N_21275,N_21317);
xnor U22860 (N_22860,N_22288,N_22347);
xor U22861 (N_22861,N_21215,N_21870);
xnor U22862 (N_22862,N_22339,N_21163);
xnor U22863 (N_22863,N_21856,N_22352);
or U22864 (N_22864,N_22154,N_21054);
xor U22865 (N_22865,N_21250,N_21420);
nor U22866 (N_22866,N_22274,N_22271);
xor U22867 (N_22867,N_21137,N_21185);
nand U22868 (N_22868,N_22217,N_21608);
and U22869 (N_22869,N_21118,N_22022);
or U22870 (N_22870,N_21073,N_22358);
nand U22871 (N_22871,N_21580,N_21831);
xor U22872 (N_22872,N_21518,N_21992);
nor U22873 (N_22873,N_21067,N_22277);
nor U22874 (N_22874,N_21116,N_22399);
or U22875 (N_22875,N_21624,N_21960);
nor U22876 (N_22876,N_21600,N_21530);
xnor U22877 (N_22877,N_21785,N_22326);
and U22878 (N_22878,N_21015,N_21141);
xor U22879 (N_22879,N_21517,N_21781);
and U22880 (N_22880,N_21979,N_22017);
nor U22881 (N_22881,N_21898,N_22062);
nand U22882 (N_22882,N_21860,N_22222);
nand U22883 (N_22883,N_21101,N_21995);
and U22884 (N_22884,N_21491,N_21535);
nand U22885 (N_22885,N_21753,N_22289);
nor U22886 (N_22886,N_21946,N_22398);
nor U22887 (N_22887,N_21627,N_21178);
or U22888 (N_22888,N_21076,N_22239);
and U22889 (N_22889,N_21360,N_21988);
and U22890 (N_22890,N_21314,N_21448);
or U22891 (N_22891,N_22035,N_21737);
and U22892 (N_22892,N_21903,N_21500);
xnor U22893 (N_22893,N_21079,N_21151);
nand U22894 (N_22894,N_21709,N_22321);
nand U22895 (N_22895,N_21019,N_22307);
nand U22896 (N_22896,N_21584,N_22246);
nand U22897 (N_22897,N_21987,N_21282);
or U22898 (N_22898,N_22126,N_21057);
nor U22899 (N_22899,N_22284,N_22369);
nor U22900 (N_22900,N_21820,N_22359);
and U22901 (N_22901,N_21572,N_21852);
nand U22902 (N_22902,N_22279,N_21914);
and U22903 (N_22903,N_21900,N_21581);
nor U22904 (N_22904,N_21964,N_22396);
and U22905 (N_22905,N_21198,N_21789);
xnor U22906 (N_22906,N_21461,N_21418);
nand U22907 (N_22907,N_22188,N_21953);
nand U22908 (N_22908,N_21761,N_21488);
and U22909 (N_22909,N_21107,N_21658);
and U22910 (N_22910,N_21438,N_21169);
xnor U22911 (N_22911,N_21044,N_21041);
xor U22912 (N_22912,N_21315,N_21729);
or U22913 (N_22913,N_21956,N_22160);
nor U22914 (N_22914,N_21227,N_21786);
or U22915 (N_22915,N_21447,N_21747);
nor U22916 (N_22916,N_21881,N_22049);
nand U22917 (N_22917,N_21172,N_21225);
nor U22918 (N_22918,N_22368,N_22008);
and U22919 (N_22919,N_22451,N_22193);
nand U22920 (N_22920,N_22377,N_21220);
and U22921 (N_22921,N_22103,N_22348);
or U22922 (N_22922,N_21695,N_21235);
nor U22923 (N_22923,N_22175,N_22416);
xor U22924 (N_22924,N_21263,N_21864);
xnor U22925 (N_22925,N_21496,N_21217);
or U22926 (N_22926,N_21080,N_22063);
and U22927 (N_22927,N_21060,N_21156);
xnor U22928 (N_22928,N_21609,N_22180);
xnor U22929 (N_22929,N_21929,N_21358);
or U22930 (N_22930,N_21356,N_21997);
nand U22931 (N_22931,N_21754,N_22013);
nor U22932 (N_22932,N_21239,N_21564);
nor U22933 (N_22933,N_22371,N_21113);
xnor U22934 (N_22934,N_21301,N_21380);
nand U22935 (N_22935,N_22422,N_21545);
nand U22936 (N_22936,N_21765,N_22283);
xor U22937 (N_22937,N_22135,N_22464);
nor U22938 (N_22938,N_21602,N_21885);
and U22939 (N_22939,N_21642,N_21454);
or U22940 (N_22940,N_21725,N_21625);
nor U22941 (N_22941,N_22303,N_22000);
nor U22942 (N_22942,N_21499,N_21982);
xnor U22943 (N_22943,N_21170,N_21521);
nor U22944 (N_22944,N_21049,N_21575);
xnor U22945 (N_22945,N_21650,N_22461);
or U22946 (N_22946,N_21088,N_21712);
nand U22947 (N_22947,N_22233,N_22350);
or U22948 (N_22948,N_22184,N_22199);
xor U22949 (N_22949,N_21901,N_21961);
and U22950 (N_22950,N_22206,N_22420);
xnor U22951 (N_22951,N_22258,N_22123);
and U22952 (N_22952,N_21698,N_22243);
or U22953 (N_22953,N_21284,N_21764);
or U22954 (N_22954,N_21583,N_22356);
xor U22955 (N_22955,N_21385,N_22299);
and U22956 (N_22956,N_22084,N_21158);
nor U22957 (N_22957,N_21745,N_22212);
nand U22958 (N_22958,N_22250,N_21248);
or U22959 (N_22959,N_21957,N_22375);
and U22960 (N_22960,N_21531,N_21493);
nor U22961 (N_22961,N_21037,N_21351);
nor U22962 (N_22962,N_21272,N_21934);
or U22963 (N_22963,N_21017,N_21114);
and U22964 (N_22964,N_21024,N_22428);
nor U22965 (N_22965,N_22337,N_21373);
xnor U22966 (N_22966,N_21586,N_22104);
and U22967 (N_22967,N_21039,N_21180);
nor U22968 (N_22968,N_22157,N_21833);
nand U22969 (N_22969,N_21553,N_21161);
nor U22970 (N_22970,N_21105,N_21818);
xnor U22971 (N_22971,N_21218,N_22082);
nand U22972 (N_22972,N_21480,N_22410);
nor U22973 (N_22973,N_21501,N_21935);
and U22974 (N_22974,N_21888,N_21569);
and U22975 (N_22975,N_22105,N_21676);
nor U22976 (N_22976,N_22012,N_21590);
nor U22977 (N_22977,N_21774,N_22482);
xor U22978 (N_22978,N_21490,N_22249);
and U22979 (N_22979,N_21293,N_22190);
nor U22980 (N_22980,N_22294,N_22293);
or U22981 (N_22981,N_21857,N_21665);
xor U22982 (N_22982,N_22480,N_22237);
or U22983 (N_22983,N_21396,N_21065);
nand U22984 (N_22984,N_21192,N_21349);
nor U22985 (N_22985,N_21242,N_21740);
nand U22986 (N_22986,N_22466,N_21630);
nor U22987 (N_22987,N_21874,N_21435);
nor U22988 (N_22988,N_22324,N_22210);
nor U22989 (N_22989,N_22430,N_21077);
or U22990 (N_22990,N_21603,N_21772);
nor U22991 (N_22991,N_21467,N_21812);
nand U22992 (N_22992,N_21570,N_21216);
nand U22993 (N_22993,N_21144,N_21511);
or U22994 (N_22994,N_21132,N_21484);
and U22995 (N_22995,N_21306,N_21084);
nor U22996 (N_22996,N_21618,N_21659);
and U22997 (N_22997,N_21933,N_21265);
nor U22998 (N_22998,N_21882,N_21557);
and U22999 (N_22999,N_21861,N_21495);
nand U23000 (N_23000,N_21811,N_21970);
nand U23001 (N_23001,N_21838,N_21074);
nor U23002 (N_23002,N_21752,N_22434);
or U23003 (N_23003,N_22057,N_21258);
nor U23004 (N_23004,N_22392,N_22149);
nand U23005 (N_23005,N_21655,N_21963);
nor U23006 (N_23006,N_21369,N_21081);
nor U23007 (N_23007,N_21354,N_21159);
and U23008 (N_23008,N_21277,N_22353);
nand U23009 (N_23009,N_21207,N_22027);
xnor U23010 (N_23010,N_22259,N_21509);
nand U23011 (N_23011,N_21893,N_21628);
nor U23012 (N_23012,N_22093,N_21510);
nand U23013 (N_23013,N_22449,N_21720);
xnor U23014 (N_23014,N_22252,N_21281);
and U23015 (N_23015,N_21723,N_21748);
or U23016 (N_23016,N_22036,N_21523);
and U23017 (N_23017,N_22044,N_22448);
nand U23018 (N_23018,N_21794,N_21384);
and U23019 (N_23019,N_21489,N_21993);
and U23020 (N_23020,N_21110,N_21673);
xor U23021 (N_23021,N_22441,N_21005);
or U23022 (N_23022,N_22363,N_21574);
nand U23023 (N_23023,N_22187,N_21398);
nor U23024 (N_23024,N_21902,N_22162);
xor U23025 (N_23025,N_21958,N_22088);
nor U23026 (N_23026,N_21756,N_21464);
nand U23027 (N_23027,N_22308,N_22462);
and U23028 (N_23028,N_21033,N_21897);
nor U23029 (N_23029,N_22437,N_21455);
or U23030 (N_23030,N_21735,N_21267);
or U23031 (N_23031,N_22298,N_21357);
nor U23032 (N_23032,N_21534,N_22075);
nor U23033 (N_23033,N_21536,N_21835);
and U23034 (N_23034,N_21639,N_21403);
and U23035 (N_23035,N_21890,N_21168);
nor U23036 (N_23036,N_22349,N_21352);
and U23037 (N_23037,N_21702,N_21950);
and U23038 (N_23038,N_21219,N_21908);
xnor U23039 (N_23039,N_22225,N_22440);
or U23040 (N_23040,N_21884,N_22302);
nor U23041 (N_23041,N_21368,N_21633);
or U23042 (N_23042,N_22095,N_21337);
xor U23043 (N_23043,N_21679,N_22139);
xnor U23044 (N_23044,N_22439,N_21839);
xnor U23045 (N_23045,N_21652,N_21050);
nand U23046 (N_23046,N_21173,N_21879);
nand U23047 (N_23047,N_21886,N_21165);
and U23048 (N_23048,N_22287,N_21750);
nand U23049 (N_23049,N_22005,N_22018);
or U23050 (N_23050,N_22203,N_21449);
xor U23051 (N_23051,N_21948,N_22178);
and U23052 (N_23052,N_21985,N_21103);
and U23053 (N_23053,N_21704,N_22272);
or U23054 (N_23054,N_22130,N_21233);
nand U23055 (N_23055,N_21867,N_21176);
nand U23056 (N_23056,N_22485,N_22236);
xnor U23057 (N_23057,N_22362,N_21123);
xnor U23058 (N_23058,N_22026,N_21669);
nor U23059 (N_23059,N_21182,N_22374);
or U23060 (N_23060,N_22471,N_21457);
nand U23061 (N_23061,N_21028,N_21641);
and U23062 (N_23062,N_21653,N_21278);
nand U23063 (N_23063,N_21474,N_21310);
or U23064 (N_23064,N_21671,N_22033);
or U23065 (N_23065,N_21909,N_21062);
nand U23066 (N_23066,N_21649,N_22028);
and U23067 (N_23067,N_21802,N_21000);
and U23068 (N_23068,N_21938,N_21303);
and U23069 (N_23069,N_21335,N_21383);
and U23070 (N_23070,N_22301,N_22421);
xnor U23071 (N_23071,N_21862,N_21423);
and U23072 (N_23072,N_21312,N_22497);
or U23073 (N_23073,N_21930,N_21841);
nor U23074 (N_23074,N_21359,N_21759);
nor U23075 (N_23075,N_22472,N_21285);
and U23076 (N_23076,N_21845,N_22169);
and U23077 (N_23077,N_22380,N_21347);
or U23078 (N_23078,N_22460,N_21672);
or U23079 (N_23079,N_21727,N_21199);
and U23080 (N_23080,N_21733,N_22181);
or U23081 (N_23081,N_21339,N_21851);
nor U23082 (N_23082,N_22423,N_22014);
and U23083 (N_23083,N_21757,N_21800);
and U23084 (N_23084,N_21376,N_21666);
nand U23085 (N_23085,N_21371,N_21439);
or U23086 (N_23086,N_21450,N_21290);
nor U23087 (N_23087,N_21766,N_22204);
nor U23088 (N_23088,N_21030,N_21405);
nor U23089 (N_23089,N_21854,N_21476);
or U23090 (N_23090,N_21120,N_21779);
and U23091 (N_23091,N_21221,N_21782);
nand U23092 (N_23092,N_21205,N_22444);
nor U23093 (N_23093,N_21601,N_21911);
nand U23094 (N_23094,N_21940,N_21955);
xor U23095 (N_23095,N_21425,N_21887);
and U23096 (N_23096,N_21522,N_21788);
and U23097 (N_23097,N_21778,N_21991);
or U23098 (N_23098,N_21108,N_21305);
xnor U23099 (N_23099,N_21682,N_22132);
and U23100 (N_23100,N_21859,N_22240);
or U23101 (N_23101,N_22333,N_21323);
xor U23102 (N_23102,N_22491,N_21719);
xor U23103 (N_23103,N_21130,N_22346);
xnor U23104 (N_23104,N_22412,N_21064);
or U23105 (N_23105,N_21251,N_21889);
and U23106 (N_23106,N_22197,N_22338);
or U23107 (N_23107,N_21497,N_21436);
or U23108 (N_23108,N_21697,N_21760);
or U23109 (N_23109,N_22261,N_21355);
or U23110 (N_23110,N_21716,N_21241);
or U23111 (N_23111,N_22414,N_22228);
xnor U23112 (N_23112,N_22164,N_21951);
xor U23113 (N_23113,N_22071,N_21962);
xnor U23114 (N_23114,N_22094,N_21936);
and U23115 (N_23115,N_22147,N_21749);
and U23116 (N_23116,N_21143,N_21177);
and U23117 (N_23117,N_21485,N_21736);
nor U23118 (N_23118,N_21891,N_21622);
xor U23119 (N_23119,N_21020,N_22156);
or U23120 (N_23120,N_21482,N_22081);
and U23121 (N_23121,N_22265,N_21426);
nand U23122 (N_23122,N_21651,N_22172);
xnor U23123 (N_23123,N_21548,N_22463);
and U23124 (N_23124,N_21266,N_22388);
xnor U23125 (N_23125,N_21945,N_21010);
xor U23126 (N_23126,N_22218,N_21939);
nand U23127 (N_23127,N_22064,N_21038);
nor U23128 (N_23128,N_21213,N_22015);
xor U23129 (N_23129,N_21621,N_22433);
xnor U23130 (N_23130,N_22251,N_22183);
nor U23131 (N_23131,N_22194,N_21459);
nor U23132 (N_23132,N_21863,N_21611);
xnor U23133 (N_23133,N_21896,N_21109);
xnor U23134 (N_23134,N_22367,N_21415);
nor U23135 (N_23135,N_21131,N_21913);
and U23136 (N_23136,N_22110,N_21072);
xnor U23137 (N_23137,N_21236,N_21375);
nand U23138 (N_23138,N_21507,N_21261);
or U23139 (N_23139,N_21431,N_21594);
and U23140 (N_23140,N_21297,N_22340);
xnor U23141 (N_23141,N_22336,N_22074);
and U23142 (N_23142,N_22100,N_21171);
or U23143 (N_23143,N_21468,N_21388);
or U23144 (N_23144,N_21470,N_21917);
nand U23145 (N_23145,N_21967,N_21361);
or U23146 (N_23146,N_22041,N_22227);
xnor U23147 (N_23147,N_21330,N_21119);
nand U23148 (N_23148,N_21167,N_21941);
xor U23149 (N_23149,N_22456,N_22291);
nor U23150 (N_23150,N_21036,N_22144);
or U23151 (N_23151,N_22122,N_21675);
xnor U23152 (N_23152,N_21989,N_21661);
or U23153 (N_23153,N_21920,N_21106);
xnor U23154 (N_23154,N_22131,N_22400);
xor U23155 (N_23155,N_21657,N_22332);
and U23156 (N_23156,N_22477,N_21070);
nor U23157 (N_23157,N_21573,N_22395);
nand U23158 (N_23158,N_22138,N_21407);
or U23159 (N_23159,N_22378,N_21834);
nand U23160 (N_23160,N_21924,N_21087);
xor U23161 (N_23161,N_22235,N_21943);
or U23162 (N_23162,N_21440,N_21598);
xor U23163 (N_23163,N_21724,N_22263);
nand U23164 (N_23164,N_21452,N_21469);
or U23165 (N_23165,N_21203,N_21596);
or U23166 (N_23166,N_21404,N_21732);
and U23167 (N_23167,N_21635,N_22025);
or U23168 (N_23168,N_21126,N_21428);
nand U23169 (N_23169,N_22278,N_22403);
xor U23170 (N_23170,N_22442,N_21068);
nor U23171 (N_23171,N_21175,N_21646);
xnor U23172 (N_23172,N_21429,N_22099);
nand U23173 (N_23173,N_21558,N_21637);
xor U23174 (N_23174,N_21477,N_22241);
and U23175 (N_23175,N_22006,N_22343);
and U23176 (N_23176,N_22209,N_21075);
nor U23177 (N_23177,N_21212,N_21708);
nand U23178 (N_23178,N_21817,N_21644);
xor U23179 (N_23179,N_22490,N_22320);
nand U23180 (N_23180,N_21364,N_21196);
xor U23181 (N_23181,N_22046,N_21907);
nor U23182 (N_23182,N_21751,N_22417);
nand U23183 (N_23183,N_21619,N_22496);
or U23184 (N_23184,N_21734,N_21412);
xor U23185 (N_23185,N_21189,N_21078);
xor U23186 (N_23186,N_21959,N_21848);
xor U23187 (N_23187,N_21847,N_21135);
nor U23188 (N_23188,N_21252,N_21479);
nand U23189 (N_23189,N_21710,N_21744);
nand U23190 (N_23190,N_21247,N_21121);
and U23191 (N_23191,N_21338,N_22468);
xnor U23192 (N_23192,N_21122,N_21430);
xor U23193 (N_23193,N_21604,N_22254);
and U23194 (N_23194,N_22319,N_22329);
or U23195 (N_23195,N_21866,N_21978);
or U23196 (N_23196,N_21214,N_22231);
xnor U23197 (N_23197,N_21582,N_21532);
and U23198 (N_23198,N_21813,N_21814);
and U23199 (N_23199,N_21981,N_22067);
nand U23200 (N_23200,N_22406,N_21634);
nor U23201 (N_23201,N_22177,N_21391);
nor U23202 (N_23202,N_21202,N_22069);
xnor U23203 (N_23203,N_22166,N_22119);
xor U23204 (N_23204,N_22142,N_22032);
nand U23205 (N_23205,N_22090,N_22195);
or U23206 (N_23206,N_22080,N_22475);
nand U23207 (N_23207,N_21249,N_22102);
and U23208 (N_23208,N_21003,N_22494);
nor U23209 (N_23209,N_21912,N_22208);
nor U23210 (N_23210,N_22499,N_21066);
nor U23211 (N_23211,N_21139,N_21014);
or U23212 (N_23212,N_21694,N_21408);
xor U23213 (N_23213,N_21906,N_21983);
xnor U23214 (N_23214,N_21792,N_21059);
nor U23215 (N_23215,N_22328,N_21873);
xnor U23216 (N_23216,N_21849,N_22065);
and U23217 (N_23217,N_21094,N_21237);
nor U23218 (N_23218,N_21458,N_22045);
nand U23219 (N_23219,N_21327,N_21071);
nand U23220 (N_23220,N_21826,N_22145);
nand U23221 (N_23221,N_21086,N_21919);
or U23222 (N_23222,N_21577,N_21345);
nand U23223 (N_23223,N_22489,N_21481);
or U23224 (N_23224,N_21894,N_21705);
and U23225 (N_23225,N_21157,N_21127);
or U23226 (N_23226,N_21954,N_21389);
nor U23227 (N_23227,N_21016,N_21421);
nand U23228 (N_23228,N_21410,N_21399);
and U23229 (N_23229,N_22248,N_21638);
nor U23230 (N_23230,N_21443,N_21230);
or U23231 (N_23231,N_21333,N_21797);
nor U23232 (N_23232,N_21990,N_21632);
nor U23233 (N_23233,N_21377,N_21925);
nand U23234 (N_23234,N_22306,N_21842);
xnor U23235 (N_23235,N_22436,N_21117);
nor U23236 (N_23236,N_21409,N_22109);
or U23237 (N_23237,N_22383,N_21828);
nand U23238 (N_23238,N_22330,N_21465);
and U23239 (N_23239,N_22234,N_21975);
nand U23240 (N_23240,N_21166,N_22136);
or U23241 (N_23241,N_22481,N_22165);
or U23242 (N_23242,N_21544,N_22229);
nor U23243 (N_23243,N_22047,N_22407);
or U23244 (N_23244,N_22312,N_21336);
xnor U23245 (N_23245,N_22327,N_21372);
or U23246 (N_23246,N_21091,N_21095);
and U23247 (N_23247,N_22072,N_21149);
or U23248 (N_23248,N_22073,N_21154);
and U23249 (N_23249,N_21090,N_21543);
nor U23250 (N_23250,N_21128,N_21574);
or U23251 (N_23251,N_22455,N_22159);
and U23252 (N_23252,N_22199,N_22391);
xor U23253 (N_23253,N_22388,N_22382);
nor U23254 (N_23254,N_22302,N_21586);
and U23255 (N_23255,N_22023,N_21606);
nor U23256 (N_23256,N_21789,N_21936);
xnor U23257 (N_23257,N_22111,N_22433);
nand U23258 (N_23258,N_21999,N_21513);
nand U23259 (N_23259,N_21541,N_21033);
nor U23260 (N_23260,N_22392,N_22388);
xnor U23261 (N_23261,N_21437,N_21742);
nor U23262 (N_23262,N_21647,N_21122);
xnor U23263 (N_23263,N_21768,N_21532);
xnor U23264 (N_23264,N_22205,N_21044);
nor U23265 (N_23265,N_22470,N_22410);
or U23266 (N_23266,N_21083,N_22339);
xnor U23267 (N_23267,N_21993,N_22440);
or U23268 (N_23268,N_21179,N_21964);
nor U23269 (N_23269,N_22445,N_21042);
nand U23270 (N_23270,N_21527,N_21486);
nand U23271 (N_23271,N_21616,N_22159);
and U23272 (N_23272,N_22421,N_22358);
or U23273 (N_23273,N_21984,N_21887);
nor U23274 (N_23274,N_22287,N_21653);
and U23275 (N_23275,N_21966,N_22365);
nand U23276 (N_23276,N_22028,N_21192);
nor U23277 (N_23277,N_22079,N_21040);
xnor U23278 (N_23278,N_21026,N_21532);
xor U23279 (N_23279,N_22276,N_21539);
and U23280 (N_23280,N_21376,N_21456);
or U23281 (N_23281,N_21344,N_22444);
and U23282 (N_23282,N_21605,N_21351);
nor U23283 (N_23283,N_22408,N_22200);
nor U23284 (N_23284,N_21068,N_21930);
xor U23285 (N_23285,N_22014,N_21696);
nand U23286 (N_23286,N_21769,N_21668);
nor U23287 (N_23287,N_22325,N_21176);
or U23288 (N_23288,N_21141,N_22225);
nand U23289 (N_23289,N_22095,N_21993);
nand U23290 (N_23290,N_22324,N_22105);
or U23291 (N_23291,N_21062,N_21084);
nand U23292 (N_23292,N_21325,N_21780);
xnor U23293 (N_23293,N_22142,N_22348);
or U23294 (N_23294,N_21303,N_22132);
or U23295 (N_23295,N_21216,N_22437);
nor U23296 (N_23296,N_21190,N_21209);
or U23297 (N_23297,N_21506,N_21296);
nand U23298 (N_23298,N_21530,N_22034);
nor U23299 (N_23299,N_21152,N_21811);
nand U23300 (N_23300,N_21270,N_21472);
and U23301 (N_23301,N_21583,N_22331);
and U23302 (N_23302,N_21109,N_21509);
and U23303 (N_23303,N_22463,N_22158);
or U23304 (N_23304,N_21628,N_22207);
and U23305 (N_23305,N_21413,N_21522);
xnor U23306 (N_23306,N_21361,N_22442);
nand U23307 (N_23307,N_21022,N_22172);
nor U23308 (N_23308,N_22096,N_21598);
and U23309 (N_23309,N_21578,N_21140);
or U23310 (N_23310,N_21124,N_22230);
and U23311 (N_23311,N_22017,N_21047);
xor U23312 (N_23312,N_21833,N_21971);
and U23313 (N_23313,N_21525,N_21367);
and U23314 (N_23314,N_21436,N_22226);
nor U23315 (N_23315,N_22335,N_21625);
nor U23316 (N_23316,N_21860,N_21866);
or U23317 (N_23317,N_21685,N_22273);
nand U23318 (N_23318,N_21592,N_21685);
nor U23319 (N_23319,N_21550,N_22490);
nand U23320 (N_23320,N_22030,N_21407);
xor U23321 (N_23321,N_21191,N_22126);
xnor U23322 (N_23322,N_21643,N_22411);
or U23323 (N_23323,N_21946,N_22077);
xor U23324 (N_23324,N_21636,N_21087);
or U23325 (N_23325,N_21639,N_21771);
and U23326 (N_23326,N_22405,N_21568);
and U23327 (N_23327,N_22157,N_21995);
xnor U23328 (N_23328,N_22028,N_21691);
and U23329 (N_23329,N_22294,N_22384);
nand U23330 (N_23330,N_22370,N_21489);
xnor U23331 (N_23331,N_21464,N_21901);
xor U23332 (N_23332,N_22175,N_21835);
nor U23333 (N_23333,N_21999,N_22391);
xor U23334 (N_23334,N_22380,N_21014);
xor U23335 (N_23335,N_21597,N_21418);
and U23336 (N_23336,N_22304,N_21652);
nor U23337 (N_23337,N_21294,N_21803);
xor U23338 (N_23338,N_21817,N_21940);
or U23339 (N_23339,N_22047,N_21127);
nor U23340 (N_23340,N_21585,N_22155);
xnor U23341 (N_23341,N_21963,N_21736);
or U23342 (N_23342,N_22414,N_21640);
or U23343 (N_23343,N_21040,N_21424);
nand U23344 (N_23344,N_21162,N_21859);
nand U23345 (N_23345,N_21855,N_22481);
xnor U23346 (N_23346,N_21882,N_21222);
nand U23347 (N_23347,N_22098,N_21536);
and U23348 (N_23348,N_22274,N_22396);
nand U23349 (N_23349,N_22090,N_22206);
or U23350 (N_23350,N_21244,N_21612);
and U23351 (N_23351,N_21548,N_21614);
nor U23352 (N_23352,N_21012,N_21023);
and U23353 (N_23353,N_21245,N_22410);
nor U23354 (N_23354,N_22377,N_21280);
or U23355 (N_23355,N_22141,N_22037);
xnor U23356 (N_23356,N_22001,N_21654);
or U23357 (N_23357,N_21833,N_21263);
nand U23358 (N_23358,N_22270,N_22173);
xor U23359 (N_23359,N_21124,N_22017);
xnor U23360 (N_23360,N_21091,N_22026);
xnor U23361 (N_23361,N_21297,N_21542);
or U23362 (N_23362,N_21882,N_22390);
and U23363 (N_23363,N_21656,N_22383);
nand U23364 (N_23364,N_21070,N_21240);
xnor U23365 (N_23365,N_21943,N_21541);
nand U23366 (N_23366,N_21291,N_22264);
xor U23367 (N_23367,N_22049,N_21221);
nand U23368 (N_23368,N_21769,N_21396);
xnor U23369 (N_23369,N_21057,N_22332);
nand U23370 (N_23370,N_22174,N_21515);
nand U23371 (N_23371,N_21879,N_21512);
xnor U23372 (N_23372,N_21277,N_21527);
xnor U23373 (N_23373,N_21829,N_21552);
and U23374 (N_23374,N_21610,N_22074);
nor U23375 (N_23375,N_21730,N_21548);
nand U23376 (N_23376,N_21739,N_21856);
nand U23377 (N_23377,N_21597,N_21767);
nand U23378 (N_23378,N_22056,N_21568);
nor U23379 (N_23379,N_22298,N_22430);
nor U23380 (N_23380,N_21331,N_22371);
nor U23381 (N_23381,N_21362,N_22251);
nor U23382 (N_23382,N_21828,N_21973);
and U23383 (N_23383,N_21304,N_21217);
nor U23384 (N_23384,N_21927,N_22449);
nand U23385 (N_23385,N_22172,N_21110);
and U23386 (N_23386,N_21227,N_21011);
xor U23387 (N_23387,N_22341,N_22250);
xor U23388 (N_23388,N_21374,N_21422);
and U23389 (N_23389,N_22166,N_21778);
and U23390 (N_23390,N_21251,N_21882);
nor U23391 (N_23391,N_21774,N_21442);
nand U23392 (N_23392,N_22237,N_21464);
or U23393 (N_23393,N_22008,N_21762);
nor U23394 (N_23394,N_21108,N_21426);
nor U23395 (N_23395,N_21882,N_21855);
xor U23396 (N_23396,N_21462,N_21107);
or U23397 (N_23397,N_21971,N_21487);
nor U23398 (N_23398,N_21399,N_21921);
and U23399 (N_23399,N_21395,N_22319);
nor U23400 (N_23400,N_21438,N_22494);
and U23401 (N_23401,N_21637,N_21580);
or U23402 (N_23402,N_21199,N_21692);
and U23403 (N_23403,N_22199,N_21179);
or U23404 (N_23404,N_21732,N_22356);
xnor U23405 (N_23405,N_21603,N_21652);
and U23406 (N_23406,N_21271,N_21764);
nand U23407 (N_23407,N_21235,N_21568);
and U23408 (N_23408,N_22457,N_22195);
xor U23409 (N_23409,N_22086,N_21423);
nand U23410 (N_23410,N_21286,N_21986);
or U23411 (N_23411,N_22066,N_22477);
and U23412 (N_23412,N_22060,N_21064);
xor U23413 (N_23413,N_21621,N_21432);
and U23414 (N_23414,N_22196,N_21221);
nor U23415 (N_23415,N_21528,N_21804);
xor U23416 (N_23416,N_21405,N_21201);
nor U23417 (N_23417,N_21907,N_21602);
xor U23418 (N_23418,N_21118,N_21745);
xor U23419 (N_23419,N_21281,N_21503);
nor U23420 (N_23420,N_22441,N_21889);
nor U23421 (N_23421,N_22222,N_21201);
or U23422 (N_23422,N_21728,N_22342);
nor U23423 (N_23423,N_21173,N_21426);
xnor U23424 (N_23424,N_21575,N_22153);
nor U23425 (N_23425,N_21363,N_21617);
nor U23426 (N_23426,N_21010,N_21496);
and U23427 (N_23427,N_21698,N_22284);
and U23428 (N_23428,N_22474,N_21625);
and U23429 (N_23429,N_21671,N_22482);
xor U23430 (N_23430,N_22487,N_21573);
or U23431 (N_23431,N_21159,N_21503);
nor U23432 (N_23432,N_22358,N_22498);
or U23433 (N_23433,N_21585,N_22404);
and U23434 (N_23434,N_22128,N_21898);
or U23435 (N_23435,N_21939,N_22186);
or U23436 (N_23436,N_21624,N_21886);
or U23437 (N_23437,N_21419,N_21323);
nand U23438 (N_23438,N_21826,N_21263);
xor U23439 (N_23439,N_21719,N_21180);
and U23440 (N_23440,N_22054,N_22480);
nor U23441 (N_23441,N_21892,N_21302);
xnor U23442 (N_23442,N_22288,N_21733);
and U23443 (N_23443,N_21526,N_21325);
nand U23444 (N_23444,N_21500,N_22231);
or U23445 (N_23445,N_21518,N_21807);
and U23446 (N_23446,N_21735,N_22002);
or U23447 (N_23447,N_21968,N_21751);
nor U23448 (N_23448,N_21660,N_21330);
nor U23449 (N_23449,N_21958,N_21290);
nor U23450 (N_23450,N_22335,N_22029);
xnor U23451 (N_23451,N_21998,N_22269);
xnor U23452 (N_23452,N_21761,N_22118);
or U23453 (N_23453,N_21448,N_22210);
nor U23454 (N_23454,N_21786,N_21848);
xor U23455 (N_23455,N_21420,N_22005);
nand U23456 (N_23456,N_21486,N_21705);
xnor U23457 (N_23457,N_21667,N_21327);
and U23458 (N_23458,N_22207,N_21346);
nor U23459 (N_23459,N_21642,N_21877);
and U23460 (N_23460,N_22418,N_21406);
nand U23461 (N_23461,N_21808,N_21394);
nand U23462 (N_23462,N_21643,N_22495);
and U23463 (N_23463,N_21171,N_21520);
nand U23464 (N_23464,N_22010,N_21978);
or U23465 (N_23465,N_21842,N_21971);
nor U23466 (N_23466,N_22313,N_21579);
xnor U23467 (N_23467,N_21524,N_21150);
or U23468 (N_23468,N_22283,N_21607);
xor U23469 (N_23469,N_21651,N_21374);
or U23470 (N_23470,N_21080,N_22367);
and U23471 (N_23471,N_21474,N_21157);
nor U23472 (N_23472,N_21173,N_21006);
or U23473 (N_23473,N_21825,N_21483);
and U23474 (N_23474,N_22401,N_21833);
nor U23475 (N_23475,N_21348,N_21539);
or U23476 (N_23476,N_21111,N_21863);
nand U23477 (N_23477,N_21529,N_21935);
and U23478 (N_23478,N_22051,N_21943);
xor U23479 (N_23479,N_21479,N_22399);
xnor U23480 (N_23480,N_21782,N_21994);
nand U23481 (N_23481,N_22219,N_21179);
and U23482 (N_23482,N_21436,N_21487);
nand U23483 (N_23483,N_21534,N_22392);
nor U23484 (N_23484,N_21090,N_21989);
nor U23485 (N_23485,N_21572,N_21790);
or U23486 (N_23486,N_21479,N_21064);
and U23487 (N_23487,N_22456,N_21318);
and U23488 (N_23488,N_22104,N_21145);
xor U23489 (N_23489,N_22091,N_21688);
or U23490 (N_23490,N_21391,N_22065);
xnor U23491 (N_23491,N_21616,N_21904);
nor U23492 (N_23492,N_21608,N_21846);
or U23493 (N_23493,N_21521,N_21957);
xor U23494 (N_23494,N_21921,N_21970);
xnor U23495 (N_23495,N_22386,N_21944);
or U23496 (N_23496,N_21164,N_22393);
xnor U23497 (N_23497,N_21616,N_21869);
or U23498 (N_23498,N_21371,N_21943);
nor U23499 (N_23499,N_22238,N_21313);
nor U23500 (N_23500,N_21795,N_21765);
xor U23501 (N_23501,N_21764,N_22082);
nor U23502 (N_23502,N_21092,N_21414);
or U23503 (N_23503,N_21181,N_21672);
nor U23504 (N_23504,N_21834,N_21829);
and U23505 (N_23505,N_22164,N_21342);
nor U23506 (N_23506,N_21287,N_22329);
nand U23507 (N_23507,N_22102,N_22153);
nor U23508 (N_23508,N_21130,N_22085);
nor U23509 (N_23509,N_21014,N_21412);
xor U23510 (N_23510,N_22017,N_21296);
nor U23511 (N_23511,N_21645,N_21523);
or U23512 (N_23512,N_22023,N_21304);
nand U23513 (N_23513,N_21603,N_21447);
nand U23514 (N_23514,N_21485,N_21693);
and U23515 (N_23515,N_21353,N_21411);
nor U23516 (N_23516,N_21451,N_21914);
nor U23517 (N_23517,N_21719,N_22385);
nor U23518 (N_23518,N_22468,N_22001);
nor U23519 (N_23519,N_22038,N_21335);
and U23520 (N_23520,N_22393,N_22467);
and U23521 (N_23521,N_21600,N_21968);
and U23522 (N_23522,N_22051,N_22211);
and U23523 (N_23523,N_22182,N_21292);
or U23524 (N_23524,N_22188,N_22409);
xor U23525 (N_23525,N_21250,N_21410);
xor U23526 (N_23526,N_21307,N_21934);
or U23527 (N_23527,N_22447,N_21003);
xor U23528 (N_23528,N_22278,N_22424);
and U23529 (N_23529,N_21094,N_22161);
nor U23530 (N_23530,N_21549,N_21327);
or U23531 (N_23531,N_21723,N_21965);
and U23532 (N_23532,N_21497,N_21226);
and U23533 (N_23533,N_21638,N_21020);
xnor U23534 (N_23534,N_21567,N_21410);
xor U23535 (N_23535,N_21175,N_22144);
nor U23536 (N_23536,N_22297,N_21576);
nor U23537 (N_23537,N_21823,N_21174);
nor U23538 (N_23538,N_21267,N_21710);
or U23539 (N_23539,N_22161,N_21490);
and U23540 (N_23540,N_21768,N_21883);
or U23541 (N_23541,N_21521,N_21154);
and U23542 (N_23542,N_21361,N_21556);
nand U23543 (N_23543,N_21794,N_22018);
nand U23544 (N_23544,N_21117,N_21298);
nand U23545 (N_23545,N_21539,N_21510);
nand U23546 (N_23546,N_21796,N_22039);
nand U23547 (N_23547,N_22044,N_22138);
xor U23548 (N_23548,N_21768,N_21172);
xnor U23549 (N_23549,N_21184,N_22071);
nand U23550 (N_23550,N_21509,N_21460);
xnor U23551 (N_23551,N_21254,N_22357);
nor U23552 (N_23552,N_22034,N_22051);
nor U23553 (N_23553,N_22387,N_21521);
or U23554 (N_23554,N_21152,N_21208);
nor U23555 (N_23555,N_22275,N_21832);
nor U23556 (N_23556,N_21002,N_21254);
or U23557 (N_23557,N_22319,N_22219);
xnor U23558 (N_23558,N_22232,N_21667);
nand U23559 (N_23559,N_21439,N_21199);
nand U23560 (N_23560,N_22306,N_21644);
nand U23561 (N_23561,N_22099,N_21995);
and U23562 (N_23562,N_22240,N_21473);
xor U23563 (N_23563,N_21618,N_21340);
nor U23564 (N_23564,N_21962,N_21509);
and U23565 (N_23565,N_22450,N_21592);
nor U23566 (N_23566,N_21433,N_21302);
xnor U23567 (N_23567,N_21383,N_22008);
nand U23568 (N_23568,N_22382,N_21394);
nand U23569 (N_23569,N_21267,N_22161);
and U23570 (N_23570,N_21989,N_21242);
nor U23571 (N_23571,N_21500,N_21795);
nand U23572 (N_23572,N_21299,N_22238);
nand U23573 (N_23573,N_22176,N_21358);
or U23574 (N_23574,N_21078,N_21646);
and U23575 (N_23575,N_21024,N_21389);
nand U23576 (N_23576,N_21042,N_21004);
and U23577 (N_23577,N_21780,N_21026);
and U23578 (N_23578,N_22493,N_21499);
and U23579 (N_23579,N_21175,N_21074);
nor U23580 (N_23580,N_22371,N_21376);
xor U23581 (N_23581,N_21910,N_21958);
or U23582 (N_23582,N_21263,N_21466);
xnor U23583 (N_23583,N_22109,N_21742);
nand U23584 (N_23584,N_21833,N_22030);
and U23585 (N_23585,N_21878,N_21513);
xor U23586 (N_23586,N_21611,N_21628);
xor U23587 (N_23587,N_22299,N_21048);
nand U23588 (N_23588,N_21732,N_21627);
and U23589 (N_23589,N_22323,N_21707);
and U23590 (N_23590,N_21714,N_22483);
nand U23591 (N_23591,N_21964,N_21354);
or U23592 (N_23592,N_21066,N_21816);
xor U23593 (N_23593,N_21995,N_22294);
nand U23594 (N_23594,N_22365,N_22201);
nor U23595 (N_23595,N_22419,N_21503);
nand U23596 (N_23596,N_22072,N_22479);
or U23597 (N_23597,N_21057,N_22382);
nand U23598 (N_23598,N_21528,N_21386);
nor U23599 (N_23599,N_21667,N_21206);
xnor U23600 (N_23600,N_21711,N_21385);
nand U23601 (N_23601,N_21427,N_21329);
nand U23602 (N_23602,N_22125,N_22176);
or U23603 (N_23603,N_22264,N_22288);
or U23604 (N_23604,N_21835,N_21659);
nand U23605 (N_23605,N_21538,N_21792);
xnor U23606 (N_23606,N_21208,N_22172);
nor U23607 (N_23607,N_21314,N_21307);
xor U23608 (N_23608,N_21519,N_21459);
or U23609 (N_23609,N_21654,N_22309);
nor U23610 (N_23610,N_21293,N_22111);
nand U23611 (N_23611,N_21927,N_21969);
nand U23612 (N_23612,N_22160,N_22095);
xor U23613 (N_23613,N_21971,N_21083);
nor U23614 (N_23614,N_21049,N_21742);
xnor U23615 (N_23615,N_22449,N_22043);
or U23616 (N_23616,N_22008,N_21925);
or U23617 (N_23617,N_22390,N_22275);
nor U23618 (N_23618,N_21784,N_21494);
and U23619 (N_23619,N_21687,N_21683);
and U23620 (N_23620,N_21057,N_22213);
nand U23621 (N_23621,N_21841,N_22252);
nor U23622 (N_23622,N_21913,N_21734);
and U23623 (N_23623,N_21207,N_22436);
or U23624 (N_23624,N_21935,N_22376);
xor U23625 (N_23625,N_22161,N_22314);
nand U23626 (N_23626,N_21014,N_21000);
nand U23627 (N_23627,N_22437,N_21026);
nor U23628 (N_23628,N_21823,N_21980);
nand U23629 (N_23629,N_21590,N_22424);
nor U23630 (N_23630,N_21973,N_21035);
or U23631 (N_23631,N_21567,N_21564);
nand U23632 (N_23632,N_22243,N_21861);
and U23633 (N_23633,N_21725,N_21929);
and U23634 (N_23634,N_21863,N_21474);
and U23635 (N_23635,N_22482,N_22130);
nor U23636 (N_23636,N_21859,N_22344);
nor U23637 (N_23637,N_21266,N_22190);
nand U23638 (N_23638,N_21735,N_22004);
nand U23639 (N_23639,N_21197,N_21051);
nor U23640 (N_23640,N_21473,N_21818);
nand U23641 (N_23641,N_22345,N_21610);
xnor U23642 (N_23642,N_21830,N_22400);
or U23643 (N_23643,N_21477,N_21807);
nor U23644 (N_23644,N_21587,N_22066);
nand U23645 (N_23645,N_21049,N_21616);
nor U23646 (N_23646,N_21097,N_21890);
or U23647 (N_23647,N_21150,N_21213);
nand U23648 (N_23648,N_21023,N_21243);
or U23649 (N_23649,N_21924,N_21476);
or U23650 (N_23650,N_21790,N_22269);
and U23651 (N_23651,N_21404,N_21514);
or U23652 (N_23652,N_22468,N_21519);
xnor U23653 (N_23653,N_21577,N_21353);
nor U23654 (N_23654,N_22480,N_21309);
xnor U23655 (N_23655,N_22214,N_22386);
and U23656 (N_23656,N_21855,N_21565);
nor U23657 (N_23657,N_21138,N_22418);
nor U23658 (N_23658,N_21507,N_21099);
nand U23659 (N_23659,N_21892,N_22309);
or U23660 (N_23660,N_21390,N_22111);
xnor U23661 (N_23661,N_21442,N_22497);
nand U23662 (N_23662,N_21848,N_22405);
xor U23663 (N_23663,N_21632,N_21352);
or U23664 (N_23664,N_21540,N_21717);
xnor U23665 (N_23665,N_21370,N_21544);
or U23666 (N_23666,N_21034,N_21735);
and U23667 (N_23667,N_22149,N_22480);
and U23668 (N_23668,N_21919,N_21088);
xor U23669 (N_23669,N_21848,N_21256);
nor U23670 (N_23670,N_22246,N_22004);
or U23671 (N_23671,N_21386,N_21070);
xnor U23672 (N_23672,N_21041,N_22369);
or U23673 (N_23673,N_22417,N_21593);
nor U23674 (N_23674,N_21686,N_21951);
nor U23675 (N_23675,N_21849,N_21437);
and U23676 (N_23676,N_22336,N_21103);
nand U23677 (N_23677,N_22101,N_21179);
nand U23678 (N_23678,N_21455,N_21839);
nor U23679 (N_23679,N_21052,N_21428);
xor U23680 (N_23680,N_22368,N_21794);
or U23681 (N_23681,N_21434,N_22000);
xnor U23682 (N_23682,N_22451,N_22053);
and U23683 (N_23683,N_22264,N_22184);
and U23684 (N_23684,N_22301,N_21785);
and U23685 (N_23685,N_21608,N_21401);
or U23686 (N_23686,N_21733,N_21760);
nor U23687 (N_23687,N_21857,N_22204);
nand U23688 (N_23688,N_22022,N_21284);
nor U23689 (N_23689,N_21124,N_22470);
and U23690 (N_23690,N_22202,N_22097);
nor U23691 (N_23691,N_22330,N_22363);
nand U23692 (N_23692,N_22388,N_22162);
and U23693 (N_23693,N_21372,N_22275);
nand U23694 (N_23694,N_21746,N_21872);
nor U23695 (N_23695,N_21030,N_22246);
nand U23696 (N_23696,N_21230,N_21137);
nor U23697 (N_23697,N_21520,N_22270);
xnor U23698 (N_23698,N_22114,N_21035);
nor U23699 (N_23699,N_21719,N_21481);
xor U23700 (N_23700,N_22485,N_21769);
xnor U23701 (N_23701,N_21981,N_22381);
and U23702 (N_23702,N_21766,N_21704);
xor U23703 (N_23703,N_21250,N_21918);
xor U23704 (N_23704,N_21978,N_21010);
xnor U23705 (N_23705,N_21834,N_21652);
or U23706 (N_23706,N_21899,N_21163);
or U23707 (N_23707,N_21490,N_21380);
nand U23708 (N_23708,N_21250,N_21203);
nand U23709 (N_23709,N_22243,N_22483);
nor U23710 (N_23710,N_21008,N_22294);
nor U23711 (N_23711,N_22094,N_21274);
nor U23712 (N_23712,N_21240,N_21090);
nand U23713 (N_23713,N_21514,N_21160);
and U23714 (N_23714,N_21292,N_21415);
nand U23715 (N_23715,N_21847,N_21633);
nor U23716 (N_23716,N_21375,N_22002);
xnor U23717 (N_23717,N_22305,N_22284);
and U23718 (N_23718,N_21594,N_21077);
or U23719 (N_23719,N_22073,N_21720);
nor U23720 (N_23720,N_21985,N_22044);
nand U23721 (N_23721,N_21604,N_21508);
and U23722 (N_23722,N_21525,N_21002);
or U23723 (N_23723,N_22315,N_21933);
nand U23724 (N_23724,N_22323,N_21156);
and U23725 (N_23725,N_22319,N_21736);
xor U23726 (N_23726,N_21822,N_21009);
or U23727 (N_23727,N_21138,N_21502);
xnor U23728 (N_23728,N_21780,N_22057);
nand U23729 (N_23729,N_21815,N_21928);
nor U23730 (N_23730,N_21739,N_21990);
nand U23731 (N_23731,N_21885,N_22286);
and U23732 (N_23732,N_21670,N_22410);
nand U23733 (N_23733,N_22005,N_21682);
nand U23734 (N_23734,N_21142,N_21020);
nand U23735 (N_23735,N_21005,N_21099);
or U23736 (N_23736,N_21566,N_21109);
or U23737 (N_23737,N_22202,N_21327);
or U23738 (N_23738,N_21062,N_22279);
xnor U23739 (N_23739,N_21674,N_21994);
xor U23740 (N_23740,N_22023,N_22089);
nor U23741 (N_23741,N_22160,N_22004);
and U23742 (N_23742,N_21610,N_21496);
nand U23743 (N_23743,N_21635,N_22396);
and U23744 (N_23744,N_21642,N_21922);
nor U23745 (N_23745,N_21633,N_21487);
and U23746 (N_23746,N_21349,N_22467);
xnor U23747 (N_23747,N_22472,N_22231);
nand U23748 (N_23748,N_21701,N_21287);
xor U23749 (N_23749,N_22206,N_21909);
nor U23750 (N_23750,N_21015,N_21428);
nand U23751 (N_23751,N_21235,N_22052);
or U23752 (N_23752,N_21739,N_21453);
nand U23753 (N_23753,N_21195,N_21911);
xnor U23754 (N_23754,N_21332,N_22444);
nand U23755 (N_23755,N_22196,N_21389);
nand U23756 (N_23756,N_21570,N_21106);
or U23757 (N_23757,N_21837,N_22080);
and U23758 (N_23758,N_21246,N_21239);
and U23759 (N_23759,N_22461,N_22212);
xor U23760 (N_23760,N_22143,N_21028);
and U23761 (N_23761,N_21384,N_22047);
xnor U23762 (N_23762,N_21195,N_22338);
or U23763 (N_23763,N_21941,N_22204);
xor U23764 (N_23764,N_21261,N_22294);
nor U23765 (N_23765,N_22467,N_21224);
and U23766 (N_23766,N_21447,N_21125);
or U23767 (N_23767,N_21195,N_21065);
xor U23768 (N_23768,N_21697,N_21116);
and U23769 (N_23769,N_21035,N_21105);
nor U23770 (N_23770,N_21543,N_21003);
xnor U23771 (N_23771,N_21442,N_21780);
nand U23772 (N_23772,N_22119,N_21670);
nand U23773 (N_23773,N_22476,N_21415);
and U23774 (N_23774,N_22242,N_22005);
or U23775 (N_23775,N_22329,N_21980);
or U23776 (N_23776,N_21124,N_21727);
and U23777 (N_23777,N_21076,N_21364);
and U23778 (N_23778,N_21419,N_21937);
or U23779 (N_23779,N_22395,N_21392);
and U23780 (N_23780,N_21518,N_21724);
and U23781 (N_23781,N_22388,N_22285);
and U23782 (N_23782,N_21398,N_21265);
xor U23783 (N_23783,N_22256,N_21285);
xor U23784 (N_23784,N_21747,N_21724);
nand U23785 (N_23785,N_22445,N_21519);
nor U23786 (N_23786,N_21835,N_21839);
and U23787 (N_23787,N_22211,N_22363);
nor U23788 (N_23788,N_22121,N_21692);
nor U23789 (N_23789,N_21139,N_22324);
nor U23790 (N_23790,N_22328,N_22406);
and U23791 (N_23791,N_21012,N_21855);
nor U23792 (N_23792,N_21993,N_21421);
nor U23793 (N_23793,N_21121,N_21344);
nand U23794 (N_23794,N_22108,N_22213);
nor U23795 (N_23795,N_21029,N_22100);
xnor U23796 (N_23796,N_21491,N_22074);
xor U23797 (N_23797,N_21231,N_21946);
or U23798 (N_23798,N_21378,N_22368);
and U23799 (N_23799,N_21036,N_21338);
nand U23800 (N_23800,N_21656,N_21356);
xnor U23801 (N_23801,N_21308,N_21898);
nand U23802 (N_23802,N_21430,N_21729);
nor U23803 (N_23803,N_21982,N_21823);
and U23804 (N_23804,N_22365,N_22487);
or U23805 (N_23805,N_21793,N_22100);
xor U23806 (N_23806,N_21133,N_21254);
nor U23807 (N_23807,N_21716,N_21096);
nand U23808 (N_23808,N_21419,N_21862);
and U23809 (N_23809,N_22155,N_21361);
nand U23810 (N_23810,N_21828,N_21965);
nor U23811 (N_23811,N_22061,N_21149);
xnor U23812 (N_23812,N_21279,N_22213);
or U23813 (N_23813,N_22284,N_21284);
or U23814 (N_23814,N_21392,N_21146);
and U23815 (N_23815,N_22445,N_21081);
nand U23816 (N_23816,N_22431,N_22228);
xor U23817 (N_23817,N_22034,N_21536);
and U23818 (N_23818,N_21163,N_21592);
xnor U23819 (N_23819,N_21229,N_21848);
xnor U23820 (N_23820,N_21064,N_21125);
nor U23821 (N_23821,N_22388,N_21022);
and U23822 (N_23822,N_21691,N_21378);
or U23823 (N_23823,N_21606,N_21468);
or U23824 (N_23824,N_22360,N_22149);
nand U23825 (N_23825,N_22472,N_22467);
nand U23826 (N_23826,N_21598,N_21878);
or U23827 (N_23827,N_22293,N_21380);
nor U23828 (N_23828,N_21100,N_21617);
and U23829 (N_23829,N_21467,N_21386);
nor U23830 (N_23830,N_22289,N_21170);
or U23831 (N_23831,N_21939,N_21568);
xnor U23832 (N_23832,N_21803,N_21877);
or U23833 (N_23833,N_21525,N_21484);
nand U23834 (N_23834,N_21723,N_21355);
nor U23835 (N_23835,N_21390,N_21420);
or U23836 (N_23836,N_22176,N_21520);
or U23837 (N_23837,N_22267,N_22064);
xnor U23838 (N_23838,N_22174,N_22241);
nor U23839 (N_23839,N_21469,N_21645);
nand U23840 (N_23840,N_22011,N_22298);
xor U23841 (N_23841,N_21414,N_21497);
and U23842 (N_23842,N_21914,N_21132);
nor U23843 (N_23843,N_21788,N_22163);
nor U23844 (N_23844,N_21425,N_22113);
and U23845 (N_23845,N_22202,N_21702);
nand U23846 (N_23846,N_21732,N_21292);
nand U23847 (N_23847,N_21881,N_21135);
and U23848 (N_23848,N_21780,N_22156);
or U23849 (N_23849,N_22275,N_21096);
nor U23850 (N_23850,N_21313,N_21126);
nand U23851 (N_23851,N_22249,N_21388);
xnor U23852 (N_23852,N_21203,N_21948);
xor U23853 (N_23853,N_21866,N_21316);
nor U23854 (N_23854,N_21697,N_21246);
or U23855 (N_23855,N_21704,N_22294);
and U23856 (N_23856,N_21481,N_21800);
nor U23857 (N_23857,N_22354,N_21775);
and U23858 (N_23858,N_21195,N_22433);
and U23859 (N_23859,N_21082,N_21522);
xor U23860 (N_23860,N_21200,N_21619);
nand U23861 (N_23861,N_21342,N_21641);
nand U23862 (N_23862,N_21103,N_21741);
or U23863 (N_23863,N_21460,N_21355);
or U23864 (N_23864,N_22471,N_21578);
nand U23865 (N_23865,N_22089,N_21026);
xor U23866 (N_23866,N_22079,N_21273);
nand U23867 (N_23867,N_21232,N_22197);
and U23868 (N_23868,N_22329,N_21482);
nor U23869 (N_23869,N_21228,N_22096);
xor U23870 (N_23870,N_21159,N_22313);
nand U23871 (N_23871,N_21000,N_21026);
nand U23872 (N_23872,N_21098,N_21965);
nor U23873 (N_23873,N_21000,N_22259);
or U23874 (N_23874,N_21759,N_21266);
or U23875 (N_23875,N_22376,N_22180);
nand U23876 (N_23876,N_22251,N_21066);
nand U23877 (N_23877,N_21773,N_21636);
nor U23878 (N_23878,N_21567,N_21029);
nor U23879 (N_23879,N_21365,N_21618);
and U23880 (N_23880,N_22147,N_21178);
xor U23881 (N_23881,N_22083,N_21663);
nand U23882 (N_23882,N_22003,N_22436);
and U23883 (N_23883,N_22021,N_21699);
xnor U23884 (N_23884,N_21099,N_21843);
nand U23885 (N_23885,N_21677,N_21438);
nor U23886 (N_23886,N_21466,N_21149);
xor U23887 (N_23887,N_22384,N_22394);
nor U23888 (N_23888,N_22245,N_22390);
and U23889 (N_23889,N_22178,N_21409);
and U23890 (N_23890,N_22373,N_21999);
xor U23891 (N_23891,N_21381,N_22489);
xor U23892 (N_23892,N_21749,N_22492);
nand U23893 (N_23893,N_21630,N_21094);
or U23894 (N_23894,N_21397,N_22076);
or U23895 (N_23895,N_21438,N_22360);
nor U23896 (N_23896,N_22122,N_21844);
nor U23897 (N_23897,N_22427,N_22265);
and U23898 (N_23898,N_21134,N_21476);
or U23899 (N_23899,N_21962,N_22061);
nand U23900 (N_23900,N_22327,N_21804);
or U23901 (N_23901,N_21711,N_22011);
nor U23902 (N_23902,N_21776,N_21450);
and U23903 (N_23903,N_21234,N_21743);
or U23904 (N_23904,N_22441,N_21219);
nor U23905 (N_23905,N_22154,N_22296);
and U23906 (N_23906,N_22212,N_22483);
xor U23907 (N_23907,N_22133,N_22134);
nor U23908 (N_23908,N_21253,N_22242);
or U23909 (N_23909,N_21274,N_21890);
nor U23910 (N_23910,N_22006,N_22367);
and U23911 (N_23911,N_22150,N_22057);
nor U23912 (N_23912,N_21272,N_21116);
nand U23913 (N_23913,N_21473,N_22183);
or U23914 (N_23914,N_22392,N_22053);
or U23915 (N_23915,N_21558,N_21460);
xnor U23916 (N_23916,N_22185,N_22125);
xnor U23917 (N_23917,N_22033,N_21611);
nand U23918 (N_23918,N_21053,N_21162);
or U23919 (N_23919,N_21005,N_21490);
nor U23920 (N_23920,N_21431,N_21007);
and U23921 (N_23921,N_22075,N_21952);
nor U23922 (N_23922,N_21172,N_21251);
xnor U23923 (N_23923,N_22048,N_21862);
nand U23924 (N_23924,N_21808,N_21816);
and U23925 (N_23925,N_21558,N_22008);
nand U23926 (N_23926,N_21945,N_21586);
xnor U23927 (N_23927,N_21409,N_21008);
xnor U23928 (N_23928,N_22404,N_22131);
nand U23929 (N_23929,N_21122,N_21240);
and U23930 (N_23930,N_21712,N_22125);
nand U23931 (N_23931,N_21076,N_22082);
or U23932 (N_23932,N_21345,N_21981);
and U23933 (N_23933,N_21240,N_21641);
nor U23934 (N_23934,N_21736,N_22403);
or U23935 (N_23935,N_21907,N_21206);
and U23936 (N_23936,N_22233,N_22264);
or U23937 (N_23937,N_21274,N_21908);
and U23938 (N_23938,N_21810,N_21076);
xor U23939 (N_23939,N_21661,N_21423);
xnor U23940 (N_23940,N_22292,N_21196);
xor U23941 (N_23941,N_22185,N_21334);
nand U23942 (N_23942,N_22296,N_22120);
and U23943 (N_23943,N_22429,N_21595);
nand U23944 (N_23944,N_22392,N_21023);
xnor U23945 (N_23945,N_22005,N_21300);
nor U23946 (N_23946,N_21853,N_21689);
xnor U23947 (N_23947,N_21927,N_22058);
or U23948 (N_23948,N_22136,N_21509);
or U23949 (N_23949,N_22298,N_22353);
nor U23950 (N_23950,N_22213,N_21118);
and U23951 (N_23951,N_21485,N_21379);
nand U23952 (N_23952,N_22348,N_21705);
nor U23953 (N_23953,N_22319,N_21200);
nor U23954 (N_23954,N_21591,N_22389);
xnor U23955 (N_23955,N_21499,N_21401);
nor U23956 (N_23956,N_21930,N_22067);
or U23957 (N_23957,N_22486,N_21289);
nand U23958 (N_23958,N_21033,N_21986);
nand U23959 (N_23959,N_21138,N_21781);
nor U23960 (N_23960,N_22376,N_22394);
nand U23961 (N_23961,N_21288,N_22215);
xnor U23962 (N_23962,N_21632,N_21955);
nand U23963 (N_23963,N_21928,N_21534);
and U23964 (N_23964,N_21450,N_21203);
nor U23965 (N_23965,N_21510,N_21569);
nor U23966 (N_23966,N_21301,N_22241);
nor U23967 (N_23967,N_22143,N_22056);
nor U23968 (N_23968,N_21165,N_21961);
or U23969 (N_23969,N_22059,N_22131);
nand U23970 (N_23970,N_21698,N_22211);
or U23971 (N_23971,N_21371,N_21123);
xor U23972 (N_23972,N_22386,N_21305);
and U23973 (N_23973,N_22060,N_22065);
or U23974 (N_23974,N_21556,N_22132);
xnor U23975 (N_23975,N_21954,N_21767);
or U23976 (N_23976,N_21049,N_22149);
and U23977 (N_23977,N_22395,N_21711);
or U23978 (N_23978,N_21757,N_21871);
xor U23979 (N_23979,N_21665,N_21728);
nor U23980 (N_23980,N_21374,N_21974);
xor U23981 (N_23981,N_22453,N_21254);
and U23982 (N_23982,N_22318,N_21051);
nand U23983 (N_23983,N_22195,N_21085);
xor U23984 (N_23984,N_21769,N_21350);
and U23985 (N_23985,N_22211,N_21158);
and U23986 (N_23986,N_21403,N_22279);
nor U23987 (N_23987,N_21854,N_22338);
xnor U23988 (N_23988,N_21185,N_21129);
or U23989 (N_23989,N_21435,N_21423);
nand U23990 (N_23990,N_21604,N_21458);
nor U23991 (N_23991,N_21246,N_21455);
nand U23992 (N_23992,N_22224,N_22214);
nor U23993 (N_23993,N_21932,N_21726);
or U23994 (N_23994,N_22012,N_22237);
and U23995 (N_23995,N_21341,N_22083);
nor U23996 (N_23996,N_21347,N_22482);
nor U23997 (N_23997,N_22047,N_22036);
xor U23998 (N_23998,N_22283,N_22144);
and U23999 (N_23999,N_22049,N_21160);
xnor U24000 (N_24000,N_22731,N_22821);
or U24001 (N_24001,N_23344,N_23426);
xor U24002 (N_24002,N_22935,N_23392);
nor U24003 (N_24003,N_22625,N_23189);
or U24004 (N_24004,N_22699,N_22514);
nand U24005 (N_24005,N_23383,N_23384);
xnor U24006 (N_24006,N_23914,N_23273);
nand U24007 (N_24007,N_22739,N_22728);
and U24008 (N_24008,N_23543,N_23138);
xor U24009 (N_24009,N_23873,N_22761);
or U24010 (N_24010,N_23869,N_23193);
nand U24011 (N_24011,N_22620,N_23494);
nand U24012 (N_24012,N_22593,N_23429);
and U24013 (N_24013,N_23456,N_23249);
or U24014 (N_24014,N_22603,N_23902);
or U24015 (N_24015,N_23659,N_23988);
xnor U24016 (N_24016,N_22910,N_22693);
and U24017 (N_24017,N_23803,N_23350);
or U24018 (N_24018,N_23747,N_23602);
and U24019 (N_24019,N_23134,N_22845);
nor U24020 (N_24020,N_23728,N_22732);
xor U24021 (N_24021,N_22850,N_23776);
nand U24022 (N_24022,N_22720,N_23744);
nand U24023 (N_24023,N_22794,N_23632);
or U24024 (N_24024,N_23644,N_23047);
and U24025 (N_24025,N_23834,N_23578);
and U24026 (N_24026,N_22635,N_23029);
or U24027 (N_24027,N_23598,N_23748);
nand U24028 (N_24028,N_23656,N_23613);
or U24029 (N_24029,N_22674,N_23178);
xor U24030 (N_24030,N_23987,N_23974);
and U24031 (N_24031,N_22614,N_23830);
nor U24032 (N_24032,N_22504,N_23587);
nor U24033 (N_24033,N_22611,N_23582);
nor U24034 (N_24034,N_23805,N_23393);
xnor U24035 (N_24035,N_22616,N_23961);
and U24036 (N_24036,N_22663,N_23810);
or U24037 (N_24037,N_22531,N_22512);
and U24038 (N_24038,N_23733,N_23851);
nand U24039 (N_24039,N_22866,N_23993);
nand U24040 (N_24040,N_23146,N_22714);
xnor U24041 (N_24041,N_22719,N_23752);
nor U24042 (N_24042,N_23214,N_23625);
xnor U24043 (N_24043,N_23052,N_23419);
and U24044 (N_24044,N_23572,N_23895);
xnor U24045 (N_24045,N_23963,N_23048);
nand U24046 (N_24046,N_23142,N_22542);
or U24047 (N_24047,N_22785,N_22647);
or U24048 (N_24048,N_22579,N_23875);
nor U24049 (N_24049,N_23493,N_23511);
or U24050 (N_24050,N_22924,N_23700);
xnor U24051 (N_24051,N_22643,N_22993);
and U24052 (N_24052,N_23729,N_23418);
xnor U24053 (N_24053,N_22927,N_22586);
or U24054 (N_24054,N_22997,N_23413);
nand U24055 (N_24055,N_23755,N_23480);
or U24056 (N_24056,N_23476,N_22873);
nand U24057 (N_24057,N_23863,N_23595);
nor U24058 (N_24058,N_22560,N_23324);
nand U24059 (N_24059,N_22944,N_23443);
xnor U24060 (N_24060,N_23321,N_23486);
and U24061 (N_24061,N_22547,N_23329);
and U24062 (N_24062,N_23897,N_23514);
or U24063 (N_24063,N_23211,N_23622);
and U24064 (N_24064,N_22583,N_22994);
and U24065 (N_24065,N_22769,N_23018);
nand U24066 (N_24066,N_23753,N_23127);
nor U24067 (N_24067,N_23120,N_22533);
nand U24068 (N_24068,N_23280,N_23741);
and U24069 (N_24069,N_22640,N_22807);
nand U24070 (N_24070,N_23496,N_23591);
nand U24071 (N_24071,N_23742,N_23505);
and U24072 (N_24072,N_22961,N_22630);
nand U24073 (N_24073,N_22926,N_23635);
or U24074 (N_24074,N_23843,N_23703);
nand U24075 (N_24075,N_22931,N_22666);
or U24076 (N_24076,N_23633,N_23787);
nor U24077 (N_24077,N_23562,N_22860);
xnor U24078 (N_24078,N_22694,N_23121);
nand U24079 (N_24079,N_23888,N_22706);
and U24080 (N_24080,N_22517,N_23536);
or U24081 (N_24081,N_22851,N_23260);
nand U24082 (N_24082,N_22729,N_22650);
nor U24083 (N_24083,N_23570,N_22528);
and U24084 (N_24084,N_23947,N_23466);
and U24085 (N_24085,N_23720,N_22917);
and U24086 (N_24086,N_23802,N_23353);
nand U24087 (N_24087,N_22555,N_22816);
nand U24088 (N_24088,N_22790,N_22757);
nor U24089 (N_24089,N_23069,N_23906);
xor U24090 (N_24090,N_23933,N_23574);
and U24091 (N_24091,N_23290,N_22770);
or U24092 (N_24092,N_22691,N_22796);
nand U24093 (N_24093,N_23323,N_23432);
and U24094 (N_24094,N_23643,N_22559);
nand U24095 (N_24095,N_23959,N_22862);
nand U24096 (N_24096,N_22908,N_22569);
xor U24097 (N_24097,N_23735,N_22737);
nor U24098 (N_24098,N_23208,N_23594);
nand U24099 (N_24099,N_22686,N_22992);
or U24100 (N_24100,N_22557,N_22525);
xor U24101 (N_24101,N_22836,N_23083);
nand U24102 (N_24102,N_23016,N_22856);
xor U24103 (N_24103,N_23495,N_23637);
xnor U24104 (N_24104,N_23490,N_23979);
nand U24105 (N_24105,N_22967,N_23912);
and U24106 (N_24106,N_23874,N_22746);
nand U24107 (N_24107,N_23149,N_22823);
xnor U24108 (N_24108,N_23283,N_23313);
xor U24109 (N_24109,N_23746,N_23401);
or U24110 (N_24110,N_23183,N_23673);
or U24111 (N_24111,N_23770,N_23256);
nor U24112 (N_24112,N_23859,N_22985);
and U24113 (N_24113,N_22521,N_23998);
and U24114 (N_24114,N_23581,N_23475);
and U24115 (N_24115,N_23119,N_23679);
and U24116 (N_24116,N_23014,N_22957);
nor U24117 (N_24117,N_23856,N_22711);
nand U24118 (N_24118,N_23816,N_23206);
nand U24119 (N_24119,N_23345,N_23986);
and U24120 (N_24120,N_23568,N_22641);
xor U24121 (N_24121,N_22991,N_23235);
nand U24122 (N_24122,N_22612,N_22621);
and U24123 (N_24123,N_22825,N_23416);
xor U24124 (N_24124,N_23144,N_23564);
nand U24125 (N_24125,N_22655,N_23903);
or U24126 (N_24126,N_22610,N_23704);
nor U24127 (N_24127,N_22921,N_23448);
nor U24128 (N_24128,N_23558,N_23483);
nand U24129 (N_24129,N_22812,N_22881);
xor U24130 (N_24130,N_22544,N_23706);
or U24131 (N_24131,N_23117,N_23672);
nor U24132 (N_24132,N_23201,N_22932);
nand U24133 (N_24133,N_22580,N_22772);
xor U24134 (N_24134,N_23455,N_22918);
nand U24135 (N_24135,N_23525,N_23956);
or U24136 (N_24136,N_22638,N_22747);
and U24137 (N_24137,N_22507,N_23714);
or U24138 (N_24138,N_23698,N_22914);
xor U24139 (N_24139,N_22778,N_23093);
nand U24140 (N_24140,N_23388,N_23254);
or U24141 (N_24141,N_23630,N_23163);
nand U24142 (N_24142,N_23534,N_22636);
nor U24143 (N_24143,N_23327,N_22986);
and U24144 (N_24144,N_23583,N_23671);
or U24145 (N_24145,N_23920,N_23592);
or U24146 (N_24146,N_23529,N_23717);
nand U24147 (N_24147,N_22869,N_22791);
nand U24148 (N_24148,N_22752,N_23306);
nand U24149 (N_24149,N_23112,N_23867);
and U24150 (N_24150,N_23537,N_23515);
and U24151 (N_24151,N_23760,N_23182);
xnor U24152 (N_24152,N_23169,N_22852);
or U24153 (N_24153,N_23111,N_23964);
and U24154 (N_24154,N_23076,N_23167);
or U24155 (N_24155,N_22605,N_23757);
or U24156 (N_24156,N_23860,N_22510);
xnor U24157 (N_24157,N_22988,N_23996);
or U24158 (N_24158,N_23406,N_23571);
nor U24159 (N_24159,N_22783,N_22654);
nor U24160 (N_24160,N_23151,N_23921);
or U24161 (N_24161,N_23941,N_23621);
xor U24162 (N_24162,N_22795,N_23506);
nor U24163 (N_24163,N_23924,N_23056);
nor U24164 (N_24164,N_22946,N_23955);
nor U24165 (N_24165,N_23415,N_22965);
xnor U24166 (N_24166,N_23533,N_23944);
or U24167 (N_24167,N_23531,N_23122);
nor U24168 (N_24168,N_23210,N_22738);
nor U24169 (N_24169,N_22589,N_22842);
and U24170 (N_24170,N_23363,N_23911);
xnor U24171 (N_24171,N_23794,N_22971);
nor U24172 (N_24172,N_23243,N_23239);
and U24173 (N_24173,N_23464,N_22948);
nor U24174 (N_24174,N_22594,N_23523);
and U24175 (N_24175,N_22668,N_23864);
and U24176 (N_24176,N_23833,N_23614);
xnor U24177 (N_24177,N_23380,N_22895);
and U24178 (N_24178,N_23532,N_22697);
or U24179 (N_24179,N_22632,N_23715);
or U24180 (N_24180,N_23768,N_23693);
nand U24181 (N_24181,N_23553,N_23784);
xor U24182 (N_24182,N_22838,N_22964);
or U24183 (N_24183,N_23450,N_22519);
xor U24184 (N_24184,N_23772,N_23109);
xnor U24185 (N_24185,N_23627,N_22744);
or U24186 (N_24186,N_23736,N_23301);
and U24187 (N_24187,N_22526,N_23657);
nand U24188 (N_24188,N_23125,N_22853);
or U24189 (N_24189,N_22870,N_23796);
nor U24190 (N_24190,N_22634,N_23268);
and U24191 (N_24191,N_22859,N_22696);
nand U24192 (N_24192,N_23597,N_22892);
nor U24193 (N_24193,N_23829,N_22798);
nor U24194 (N_24194,N_23198,N_23187);
and U24195 (N_24195,N_23585,N_23152);
nand U24196 (N_24196,N_23428,N_23230);
or U24197 (N_24197,N_22886,N_23965);
and U24198 (N_24198,N_23909,N_23219);
nor U24199 (N_24199,N_23369,N_22960);
nand U24200 (N_24200,N_23130,N_23872);
nand U24201 (N_24201,N_22916,N_22658);
and U24202 (N_24202,N_22773,N_22609);
and U24203 (N_24203,N_23849,N_23050);
nand U24204 (N_24204,N_22767,N_23228);
nand U24205 (N_24205,N_23465,N_22867);
and U24206 (N_24206,N_23275,N_23177);
nand U24207 (N_24207,N_23293,N_23844);
xnor U24208 (N_24208,N_23368,N_23586);
or U24209 (N_24209,N_22736,N_22940);
nand U24210 (N_24210,N_22597,N_23894);
nand U24211 (N_24211,N_23205,N_23539);
xor U24212 (N_24212,N_22864,N_22628);
nor U24213 (N_24213,N_23173,N_23516);
nor U24214 (N_24214,N_23137,N_22585);
and U24215 (N_24215,N_23217,N_22802);
nor U24216 (N_24216,N_23269,N_23129);
xnor U24217 (N_24217,N_22561,N_23351);
or U24218 (N_24218,N_23164,N_22692);
xor U24219 (N_24219,N_22570,N_22680);
nand U24220 (N_24220,N_23017,N_22941);
nand U24221 (N_24221,N_22741,N_23054);
nand U24222 (N_24222,N_23446,N_23795);
xor U24223 (N_24223,N_23066,N_22690);
or U24224 (N_24224,N_22797,N_23139);
xor U24225 (N_24225,N_22846,N_22743);
xor U24226 (N_24226,N_23542,N_23030);
xnor U24227 (N_24227,N_23576,N_23241);
and U24228 (N_24228,N_23811,N_22565);
nand U24229 (N_24229,N_22750,N_23629);
nand U24230 (N_24230,N_23147,N_22820);
and U24231 (N_24231,N_23389,N_22899);
or U24232 (N_24232,N_23006,N_22800);
nor U24233 (N_24233,N_23404,N_23997);
xor U24234 (N_24234,N_23638,N_23412);
nand U24235 (N_24235,N_23407,N_22629);
and U24236 (N_24236,N_23391,N_23100);
nand U24237 (N_24237,N_23690,N_23482);
or U24238 (N_24238,N_23791,N_22751);
or U24239 (N_24239,N_23754,N_22677);
nor U24240 (N_24240,N_22541,N_23408);
nand U24241 (N_24241,N_23609,N_22806);
nor U24242 (N_24242,N_22534,N_22540);
and U24243 (N_24243,N_23799,N_22811);
or U24244 (N_24244,N_23341,N_23086);
nor U24245 (N_24245,N_23927,N_23234);
xnor U24246 (N_24246,N_22530,N_22513);
xor U24247 (N_24247,N_22676,N_23185);
xor U24248 (N_24248,N_22607,N_23326);
nand U24249 (N_24249,N_23981,N_22619);
and U24250 (N_24250,N_23232,N_22735);
nor U24251 (N_24251,N_22606,N_22522);
nor U24252 (N_24252,N_23781,N_22562);
nor U24253 (N_24253,N_23821,N_22813);
and U24254 (N_24254,N_23718,N_23618);
xnor U24255 (N_24255,N_23299,N_22553);
or U24256 (N_24256,N_23061,N_23347);
nor U24257 (N_24257,N_23689,N_22930);
xor U24258 (N_24258,N_23161,N_23552);
nor U24259 (N_24259,N_23454,N_22646);
and U24260 (N_24260,N_23108,N_23952);
nand U24261 (N_24261,N_23879,N_22656);
or U24262 (N_24262,N_23845,N_23291);
nor U24263 (N_24263,N_23145,N_23155);
xor U24264 (N_24264,N_23237,N_23267);
xnor U24265 (N_24265,N_23132,N_22575);
xnor U24266 (N_24266,N_23284,N_23611);
nor U24267 (N_24267,N_23584,N_23320);
and U24268 (N_24268,N_23190,N_22968);
nor U24269 (N_24269,N_23563,N_23910);
or U24270 (N_24270,N_23339,N_22536);
xnor U24271 (N_24271,N_23785,N_22716);
nand U24272 (N_24272,N_23855,N_23648);
or U24273 (N_24273,N_23491,N_23654);
or U24274 (N_24274,N_23010,N_23436);
or U24275 (N_24275,N_23352,N_22915);
nand U24276 (N_24276,N_23686,N_23527);
and U24277 (N_24277,N_23021,N_23362);
and U24278 (N_24278,N_22730,N_23946);
and U24279 (N_24279,N_23687,N_23213);
nand U24280 (N_24280,N_22573,N_22661);
or U24281 (N_24281,N_23890,N_23303);
nand U24282 (N_24282,N_23433,N_23257);
nor U24283 (N_24283,N_23786,N_23764);
nor U24284 (N_24284,N_23647,N_23898);
and U24285 (N_24285,N_23312,N_23364);
xor U24286 (N_24286,N_23042,N_23857);
nor U24287 (N_24287,N_22755,N_22937);
nand U24288 (N_24288,N_22774,N_22911);
or U24289 (N_24289,N_23423,N_23295);
nand U24290 (N_24290,N_23004,N_22854);
nand U24291 (N_24291,N_23503,N_23031);
nand U24292 (N_24292,N_23246,N_22984);
or U24293 (N_24293,N_22887,N_23440);
or U24294 (N_24294,N_23342,N_23188);
or U24295 (N_24295,N_23174,N_23469);
and U24296 (N_24296,N_23677,N_23800);
nor U24297 (N_24297,N_23904,N_22515);
and U24298 (N_24298,N_23215,N_23868);
nand U24299 (N_24299,N_22799,N_22618);
nand U24300 (N_24300,N_22524,N_22828);
or U24301 (N_24301,N_22718,N_22637);
or U24302 (N_24302,N_22703,N_23668);
nand U24303 (N_24303,N_23296,N_23601);
or U24304 (N_24304,N_22977,N_23750);
and U24305 (N_24305,N_23074,N_23285);
nor U24306 (N_24306,N_23925,N_22841);
and U24307 (N_24307,N_23024,N_23740);
xor U24308 (N_24308,N_23304,N_23058);
and U24309 (N_24309,N_23915,N_23624);
or U24310 (N_24310,N_23396,N_23658);
or U24311 (N_24311,N_23402,N_22602);
nand U24312 (N_24312,N_23682,N_23390);
and U24313 (N_24313,N_23953,N_23549);
and U24314 (N_24314,N_23308,N_23500);
nor U24315 (N_24315,N_23809,N_22775);
nor U24316 (N_24316,N_22554,N_23115);
and U24317 (N_24317,N_23634,N_23359);
xor U24318 (N_24318,N_23192,N_23937);
xor U24319 (N_24319,N_23039,N_22564);
nand U24320 (N_24320,N_23331,N_23261);
and U24321 (N_24321,N_23013,N_23360);
xnor U24322 (N_24322,N_23498,N_23073);
or U24323 (N_24323,N_23623,N_22893);
nor U24324 (N_24324,N_23691,N_22987);
xor U24325 (N_24325,N_23992,N_23097);
nand U24326 (N_24326,N_23950,N_23451);
and U24327 (N_24327,N_23288,N_23734);
and U24328 (N_24328,N_23832,N_23779);
nand U24329 (N_24329,N_23227,N_23271);
and U24330 (N_24330,N_23939,N_23015);
and U24331 (N_24331,N_23279,N_23887);
nand U24332 (N_24332,N_23355,N_23931);
or U24333 (N_24333,N_22883,N_23166);
nor U24334 (N_24334,N_23730,N_23431);
xor U24335 (N_24335,N_23991,N_22803);
nand U24336 (N_24336,N_23005,N_22506);
or U24337 (N_24337,N_23999,N_22576);
or U24338 (N_24338,N_22804,N_22546);
and U24339 (N_24339,N_23688,N_23639);
nor U24340 (N_24340,N_22702,N_22882);
or U24341 (N_24341,N_22644,N_23274);
or U24342 (N_24342,N_23699,N_23289);
nor U24343 (N_24343,N_23224,N_22532);
or U24344 (N_24344,N_23619,N_23540);
nor U24345 (N_24345,N_22815,N_22768);
nor U24346 (N_24346,N_23773,N_23510);
xnor U24347 (N_24347,N_23901,N_23798);
or U24348 (N_24348,N_22685,N_23348);
nor U24349 (N_24349,N_23171,N_23116);
or U24350 (N_24350,N_22981,N_23971);
or U24351 (N_24351,N_23528,N_22793);
and U24352 (N_24352,N_23819,N_23938);
nand U24353 (N_24353,N_23775,N_22724);
nor U24354 (N_24354,N_22669,N_22901);
xor U24355 (N_24355,N_22889,N_23445);
xnor U24356 (N_24356,N_22857,N_22518);
nor U24357 (N_24357,N_22884,N_23852);
nand U24358 (N_24358,N_22885,N_23333);
and U24359 (N_24359,N_23104,N_23535);
or U24360 (N_24360,N_22969,N_22776);
nor U24361 (N_24361,N_23970,N_23731);
or U24362 (N_24362,N_22558,N_23509);
xnor U24363 (N_24363,N_23447,N_22749);
nand U24364 (N_24364,N_23133,N_23761);
and U24365 (N_24365,N_22617,N_23172);
nor U24366 (N_24366,N_23221,N_22936);
or U24367 (N_24367,N_23881,N_23762);
xor U24368 (N_24368,N_23545,N_23878);
nor U24369 (N_24369,N_23573,N_23064);
xnor U24370 (N_24370,N_23685,N_23453);
or U24371 (N_24371,N_23756,N_23376);
nand U24372 (N_24372,N_22779,N_23989);
xnor U24373 (N_24373,N_23317,N_23410);
and U24374 (N_24374,N_23311,N_23826);
or U24375 (N_24375,N_23281,N_23732);
nor U24376 (N_24376,N_23272,N_23371);
and U24377 (N_24377,N_22649,N_23357);
nor U24378 (N_24378,N_22989,N_22976);
or U24379 (N_24379,N_23305,N_22626);
or U24380 (N_24380,N_22608,N_23943);
nor U24381 (N_24381,N_23969,N_23737);
nor U24382 (N_24382,N_23053,N_23660);
or U24383 (N_24383,N_22639,N_22912);
or U24384 (N_24384,N_23782,N_23470);
or U24385 (N_24385,N_23560,N_23365);
and U24386 (N_24386,N_23824,N_22789);
or U24387 (N_24387,N_23011,N_23608);
nor U24388 (N_24388,N_23695,N_23497);
xor U24389 (N_24389,N_23765,N_23425);
xor U24390 (N_24390,N_23936,N_23265);
nand U24391 (N_24391,N_23065,N_22837);
xor U24392 (N_24392,N_22704,N_22945);
xor U24393 (N_24393,N_23319,N_22900);
nand U24394 (N_24394,N_22786,N_23777);
xnor U24395 (N_24395,N_23663,N_22672);
or U24396 (N_24396,N_23107,N_22771);
and U24397 (N_24397,N_23136,N_23292);
xnor U24398 (N_24398,N_23049,N_22670);
and U24399 (N_24399,N_22721,N_23942);
nand U24400 (N_24400,N_23000,N_22698);
xor U24401 (N_24401,N_23814,N_23057);
nor U24402 (N_24402,N_23612,N_22966);
nor U24403 (N_24403,N_23322,N_23615);
xor U24404 (N_24404,N_23207,N_23876);
or U24405 (N_24405,N_23488,N_23278);
and U24406 (N_24406,N_23788,N_23244);
nand U24407 (N_24407,N_23579,N_23141);
or U24408 (N_24408,N_23973,N_23085);
nand U24409 (N_24409,N_23884,N_22662);
or U24410 (N_24410,N_23179,N_23835);
xor U24411 (N_24411,N_23094,N_23062);
nor U24412 (N_24412,N_22678,N_22500);
nand U24413 (N_24413,N_23526,N_23096);
xor U24414 (N_24414,N_23160,N_23398);
or U24415 (N_24415,N_23546,N_23945);
or U24416 (N_24416,N_23847,N_23727);
and U24417 (N_24417,N_22934,N_22923);
nor U24418 (N_24418,N_23655,N_22502);
xnor U24419 (N_24419,N_22613,N_22947);
xor U24420 (N_24420,N_22995,N_23520);
xor U24421 (N_24421,N_22578,N_23191);
nor U24422 (N_24422,N_23841,N_23087);
and U24423 (N_24423,N_22511,N_23837);
and U24424 (N_24424,N_23046,N_23403);
and U24425 (N_24425,N_22682,N_23951);
nor U24426 (N_24426,N_23458,N_22954);
or U24427 (N_24427,N_22942,N_23865);
xnor U24428 (N_24428,N_23547,N_22726);
nand U24429 (N_24429,N_23091,N_23131);
or U24430 (N_24430,N_23702,N_23896);
nor U24431 (N_24431,N_23665,N_23745);
nor U24432 (N_24432,N_23966,N_23180);
and U24433 (N_24433,N_22582,N_23170);
or U24434 (N_24434,N_22700,N_22835);
or U24435 (N_24435,N_22801,N_23675);
or U24436 (N_24436,N_23710,N_22764);
or U24437 (N_24437,N_23853,N_23033);
nand U24438 (N_24438,N_23967,N_22808);
or U24439 (N_24439,N_23502,N_22535);
or U24440 (N_24440,N_23681,N_23025);
nand U24441 (N_24441,N_23978,N_23580);
or U24442 (N_24442,N_23551,N_22727);
nand U24443 (N_24443,N_23110,N_22707);
xor U24444 (N_24444,N_23334,N_23070);
xnor U24445 (N_24445,N_23818,N_22958);
nor U24446 (N_24446,N_23457,N_22701);
and U24447 (N_24447,N_22834,N_22903);
nor U24448 (N_24448,N_23556,N_23705);
and U24449 (N_24449,N_23977,N_23653);
or U24450 (N_24450,N_22508,N_23538);
xnor U24451 (N_24451,N_23079,N_23492);
nand U24452 (N_24452,N_23007,N_23994);
nand U24453 (N_24453,N_23790,N_23009);
and U24454 (N_24454,N_22715,N_23315);
nand U24455 (N_24455,N_23519,N_23697);
and U24456 (N_24456,N_23157,N_23922);
nand U24457 (N_24457,N_22844,N_22827);
and U24458 (N_24458,N_23958,N_23589);
and U24459 (N_24459,N_22591,N_23680);
xor U24460 (N_24460,N_23893,N_23223);
xnor U24461 (N_24461,N_23354,N_22833);
and U24462 (N_24462,N_23815,N_23721);
and U24463 (N_24463,N_22933,N_23212);
nand U24464 (N_24464,N_23442,N_22868);
or U24465 (N_24465,N_22550,N_23128);
and U24466 (N_24466,N_22909,N_22861);
nor U24467 (N_24467,N_23176,N_23678);
and U24468 (N_24468,N_22734,N_22951);
nor U24469 (N_24469,N_23892,N_23566);
or U24470 (N_24470,N_23034,N_23825);
nand U24471 (N_24471,N_22843,N_23975);
nand U24472 (N_24472,N_22847,N_23692);
nor U24473 (N_24473,N_23330,N_23032);
nor U24474 (N_24474,N_23027,N_22998);
or U24475 (N_24475,N_23441,N_22505);
and U24476 (N_24476,N_23962,N_23780);
or U24477 (N_24477,N_23038,N_22596);
nand U24478 (N_24478,N_23225,N_22972);
nor U24479 (N_24479,N_22713,N_22955);
nand U24480 (N_24480,N_23381,N_23332);
nand U24481 (N_24481,N_23233,N_23508);
nand U24482 (N_24482,N_23374,N_22782);
or U24483 (N_24483,N_23544,N_23302);
and U24484 (N_24484,N_23738,N_23885);
or U24485 (N_24485,N_23485,N_23926);
xor U24486 (N_24486,N_23593,N_22710);
or U24487 (N_24487,N_23739,N_22717);
and U24488 (N_24488,N_22953,N_22982);
or U24489 (N_24489,N_22563,N_23968);
and U24490 (N_24490,N_23907,N_23262);
or U24491 (N_24491,N_22872,N_23603);
and U24492 (N_24492,N_23263,N_22759);
or U24493 (N_24493,N_23866,N_23077);
and U24494 (N_24494,N_23080,N_23793);
nand U24495 (N_24495,N_23471,N_23759);
or U24496 (N_24496,N_23850,N_23449);
nand U24497 (N_24497,N_22631,N_23026);
or U24498 (N_24498,N_23277,N_22826);
and U24499 (N_24499,N_23848,N_22863);
nor U24500 (N_24500,N_23719,N_22874);
nor U24501 (N_24501,N_23886,N_22667);
nor U24502 (N_24502,N_22571,N_23022);
nand U24503 (N_24503,N_23003,N_22577);
nor U24504 (N_24504,N_23590,N_23530);
or U24505 (N_24505,N_22879,N_22758);
nand U24506 (N_24506,N_23983,N_22651);
and U24507 (N_24507,N_23645,N_23328);
nand U24508 (N_24508,N_23518,N_22979);
xnor U24509 (N_24509,N_22840,N_23106);
and U24510 (N_24510,N_22659,N_23153);
nor U24511 (N_24511,N_23420,N_23250);
and U24512 (N_24512,N_23020,N_23995);
nand U24513 (N_24513,N_23023,N_22509);
or U24514 (N_24514,N_23238,N_22978);
or U24515 (N_24515,N_23438,N_23555);
or U24516 (N_24516,N_23186,N_23666);
nor U24517 (N_24517,N_22708,N_22983);
nand U24518 (N_24518,N_22622,N_23043);
and U24519 (N_24519,N_22814,N_23220);
xor U24520 (N_24520,N_22633,N_23199);
xor U24521 (N_24521,N_22980,N_23379);
nor U24522 (N_24522,N_23882,N_23916);
nor U24523 (N_24523,N_22598,N_22970);
and U24524 (N_24524,N_23806,N_23218);
or U24525 (N_24525,N_22645,N_23891);
and U24526 (N_24526,N_23708,N_23102);
or U24527 (N_24527,N_23366,N_22722);
nand U24528 (N_24528,N_23797,N_22890);
nand U24529 (N_24529,N_23694,N_23976);
and U24530 (N_24530,N_22523,N_22681);
nand U24531 (N_24531,N_23071,N_23674);
nand U24532 (N_24532,N_23828,N_23960);
nor U24533 (N_24533,N_23035,N_23044);
or U24534 (N_24534,N_22878,N_23245);
nand U24535 (N_24535,N_22805,N_22963);
nand U24536 (N_24536,N_23636,N_22929);
xor U24537 (N_24537,N_23934,N_23954);
xnor U24538 (N_24538,N_23118,N_22642);
and U24539 (N_24539,N_23567,N_23041);
nor U24540 (N_24540,N_23600,N_23055);
or U24541 (N_24541,N_23099,N_22817);
nor U24542 (N_24542,N_23474,N_23883);
nor U24543 (N_24543,N_23662,N_23631);
or U24544 (N_24544,N_22831,N_22660);
and U24545 (N_24545,N_22683,N_23184);
nor U24546 (N_24546,N_23051,N_23801);
or U24547 (N_24547,N_22830,N_23307);
nor U24548 (N_24548,N_23461,N_23287);
nor U24549 (N_24549,N_23930,N_22684);
nor U24550 (N_24550,N_23255,N_22538);
and U24551 (N_24551,N_23231,N_22529);
or U24552 (N_24552,N_22648,N_22865);
and U24553 (N_24553,N_23081,N_22552);
nor U24554 (N_24554,N_23463,N_23716);
xnor U24555 (N_24555,N_23378,N_23854);
nor U24556 (N_24556,N_23575,N_23550);
or U24557 (N_24557,N_23604,N_23820);
nand U24558 (N_24558,N_23373,N_23778);
xnor U24559 (N_24559,N_22787,N_23259);
nor U24560 (N_24560,N_23842,N_22832);
nor U24561 (N_24561,N_23616,N_22962);
nor U24562 (N_24562,N_23226,N_23338);
nand U24563 (N_24563,N_23222,N_22996);
and U24564 (N_24564,N_23124,N_23399);
nor U24565 (N_24565,N_23175,N_23282);
and U24566 (N_24566,N_22688,N_22876);
nor U24567 (N_24567,N_22974,N_22590);
or U24568 (N_24568,N_22766,N_23248);
nor U24569 (N_24569,N_23504,N_22990);
or U24570 (N_24570,N_22780,N_23276);
nand U24571 (N_24571,N_23871,N_22595);
or U24572 (N_24572,N_23628,N_22689);
or U24573 (N_24573,N_23807,N_22788);
and U24574 (N_24574,N_23652,N_23385);
nor U24575 (N_24575,N_23664,N_23711);
and U24576 (N_24576,N_23513,N_23229);
and U24577 (N_24577,N_23557,N_23068);
and U24578 (N_24578,N_23103,N_23928);
nor U24579 (N_24579,N_23067,N_23541);
nand U24580 (N_24580,N_22950,N_23763);
nand U24581 (N_24581,N_23985,N_22896);
and U24582 (N_24582,N_22549,N_23683);
xnor U24583 (N_24583,N_22712,N_23840);
or U24584 (N_24584,N_23372,N_22973);
nor U24585 (N_24585,N_22545,N_23707);
nand U24586 (N_24586,N_23913,N_22723);
or U24587 (N_24587,N_23661,N_22753);
xnor U24588 (N_24588,N_23019,N_23386);
and U24589 (N_24589,N_23252,N_23670);
or U24590 (N_24590,N_22566,N_23923);
xnor U24591 (N_24591,N_23467,N_22839);
xor U24592 (N_24592,N_23713,N_23427);
or U24593 (N_24593,N_23751,N_23251);
nand U24594 (N_24594,N_23297,N_23197);
nand U24595 (N_24595,N_22624,N_23861);
and U24596 (N_24596,N_23101,N_23478);
xor U24597 (N_24597,N_22919,N_22763);
nor U24598 (N_24598,N_23060,N_23387);
and U24599 (N_24599,N_23105,N_23195);
xnor U24600 (N_24600,N_23468,N_23487);
xnor U24601 (N_24601,N_23804,N_23517);
xnor U24602 (N_24602,N_22925,N_23340);
or U24603 (N_24603,N_23424,N_23696);
nor U24604 (N_24604,N_23375,N_22592);
or U24605 (N_24605,N_23484,N_22745);
or U24606 (N_24606,N_23148,N_23294);
or U24607 (N_24607,N_23726,N_22587);
xor U24608 (N_24608,N_23114,N_22907);
or U24609 (N_24609,N_22855,N_23247);
nor U24610 (N_24610,N_23253,N_23599);
and U24611 (N_24611,N_23088,N_22503);
xor U24612 (N_24612,N_23499,N_22849);
nor U24613 (N_24613,N_23001,N_22543);
nand U24614 (N_24614,N_22922,N_23749);
nor U24615 (N_24615,N_23554,N_23522);
and U24616 (N_24616,N_22653,N_23676);
and U24617 (N_24617,N_22537,N_23712);
nor U24618 (N_24618,N_23439,N_23501);
xnor U24619 (N_24619,N_22623,N_23789);
and U24620 (N_24620,N_23168,N_23150);
and U24621 (N_24621,N_23240,N_23045);
nor U24622 (N_24622,N_22765,N_23135);
xnor U24623 (N_24623,N_23889,N_23588);
xor U24624 (N_24624,N_22568,N_22810);
nand U24625 (N_24625,N_23336,N_22705);
nand U24626 (N_24626,N_23298,N_23846);
and U24627 (N_24627,N_23817,N_23343);
xnor U24628 (N_24628,N_23948,N_23565);
nand U24629 (N_24629,N_22740,N_22627);
xor U24630 (N_24630,N_23831,N_23669);
or U24631 (N_24631,N_23036,N_23434);
and U24632 (N_24632,N_23827,N_23642);
nand U24633 (N_24633,N_23908,N_23430);
nand U24634 (N_24634,N_22920,N_23900);
or U24635 (N_24635,N_23813,N_23349);
nand U24636 (N_24636,N_23400,N_23481);
nor U24637 (N_24637,N_22664,N_22581);
xnor U24638 (N_24638,N_22501,N_23200);
nand U24639 (N_24639,N_23489,N_23877);
nor U24640 (N_24640,N_22905,N_23310);
or U24641 (N_24641,N_22733,N_22975);
nor U24642 (N_24642,N_23918,N_23822);
and U24643 (N_24643,N_23382,N_23414);
xnor U24644 (N_24644,N_23258,N_23507);
xnor U24645 (N_24645,N_23409,N_23684);
or U24646 (N_24646,N_23316,N_23264);
xnor U24647 (N_24647,N_23990,N_22516);
or U24648 (N_24648,N_23335,N_23143);
and U24649 (N_24649,N_23156,N_23082);
and U24650 (N_24650,N_23090,N_23394);
and U24651 (N_24651,N_23159,N_22959);
xnor U24652 (N_24652,N_23722,N_23242);
nor U24653 (N_24653,N_22906,N_22657);
nand U24654 (N_24654,N_23361,N_23650);
xor U24655 (N_24655,N_23524,N_23709);
nand U24656 (N_24656,N_23008,N_23905);
nor U24657 (N_24657,N_23089,N_22551);
or U24658 (N_24658,N_23437,N_23949);
xnor U24659 (N_24659,N_23858,N_22880);
and U24660 (N_24660,N_22599,N_23367);
and U24661 (N_24661,N_22601,N_23377);
xor U24662 (N_24662,N_22679,N_22556);
xnor U24663 (N_24663,N_23626,N_23569);
nand U24664 (N_24664,N_23605,N_23640);
and U24665 (N_24665,N_23196,N_23012);
and U24666 (N_24666,N_23646,N_23561);
nand U24667 (N_24667,N_23641,N_22709);
nor U24668 (N_24668,N_23606,N_23078);
nand U24669 (N_24669,N_23607,N_23723);
xor U24670 (N_24670,N_23063,N_23422);
nor U24671 (N_24671,N_23899,N_23808);
and U24672 (N_24672,N_23405,N_23577);
and U24673 (N_24673,N_23957,N_23202);
xor U24674 (N_24674,N_22600,N_22897);
xnor U24675 (N_24675,N_23126,N_22858);
nand U24676 (N_24676,N_23204,N_22781);
and U24677 (N_24677,N_23459,N_23266);
and U24678 (N_24678,N_22898,N_22567);
xnor U24679 (N_24679,N_23521,N_22818);
nand U24680 (N_24680,N_23559,N_23870);
and U24681 (N_24681,N_23084,N_22687);
nand U24682 (N_24682,N_23370,N_23037);
nand U24683 (N_24683,N_23411,N_23783);
nor U24684 (N_24684,N_22894,N_23417);
xor U24685 (N_24685,N_22572,N_23984);
nand U24686 (N_24686,N_22695,N_23473);
nor U24687 (N_24687,N_22760,N_23158);
xnor U24688 (N_24688,N_23059,N_23203);
or U24689 (N_24689,N_22928,N_22809);
xnor U24690 (N_24690,N_23839,N_23452);
and U24691 (N_24691,N_22665,N_22822);
and U24692 (N_24692,N_22938,N_23919);
nand U24693 (N_24693,N_23397,N_22891);
nand U24694 (N_24694,N_22904,N_22673);
nand U24695 (N_24695,N_23935,N_23972);
xor U24696 (N_24696,N_23325,N_22829);
xnor U24697 (N_24697,N_23472,N_22824);
nor U24698 (N_24698,N_23462,N_23724);
nor U24699 (N_24699,N_23337,N_23838);
and U24700 (N_24700,N_23140,N_23075);
xnor U24701 (N_24701,N_23917,N_22902);
and U24702 (N_24702,N_22675,N_23300);
nand U24703 (N_24703,N_23358,N_22574);
xnor U24704 (N_24704,N_22875,N_22548);
nor U24705 (N_24705,N_22652,N_23620);
nand U24706 (N_24706,N_23098,N_23836);
nor U24707 (N_24707,N_23165,N_23286);
nor U24708 (N_24708,N_23477,N_22671);
and U24709 (N_24709,N_22584,N_22754);
and U24710 (N_24710,N_22939,N_23812);
nand U24711 (N_24711,N_23743,N_22952);
xor U24712 (N_24712,N_23460,N_23181);
or U24713 (N_24713,N_23610,N_22848);
nor U24714 (N_24714,N_22588,N_22762);
or U24715 (N_24715,N_23667,N_22792);
or U24716 (N_24716,N_22539,N_23940);
nand U24717 (N_24717,N_23649,N_23318);
or U24718 (N_24718,N_22527,N_23162);
nor U24719 (N_24719,N_23270,N_23309);
or U24720 (N_24720,N_23701,N_22784);
and U24721 (N_24721,N_22913,N_23216);
nand U24722 (N_24722,N_22956,N_23767);
and U24723 (N_24723,N_22520,N_23617);
and U24724 (N_24724,N_23002,N_23512);
nor U24725 (N_24725,N_23095,N_22877);
nand U24726 (N_24726,N_23651,N_22949);
xor U24727 (N_24727,N_23123,N_23880);
or U24728 (N_24728,N_23346,N_23823);
and U24729 (N_24729,N_23072,N_23236);
xnor U24730 (N_24730,N_23932,N_23548);
and U24731 (N_24731,N_23154,N_23479);
nor U24732 (N_24732,N_23435,N_23028);
xor U24733 (N_24733,N_22888,N_23792);
nor U24734 (N_24734,N_23092,N_23980);
nor U24735 (N_24735,N_23769,N_23113);
nand U24736 (N_24736,N_23774,N_23194);
nor U24737 (N_24737,N_22999,N_23421);
nor U24738 (N_24738,N_23395,N_22819);
xnor U24739 (N_24739,N_22756,N_22604);
or U24740 (N_24740,N_22615,N_23314);
nor U24741 (N_24741,N_22943,N_23725);
or U24742 (N_24742,N_23862,N_23444);
xor U24743 (N_24743,N_22777,N_23040);
or U24744 (N_24744,N_23209,N_22871);
nand U24745 (N_24745,N_23771,N_23596);
and U24746 (N_24746,N_23356,N_23758);
xnor U24747 (N_24747,N_22748,N_23982);
nand U24748 (N_24748,N_23766,N_23929);
or U24749 (N_24749,N_22725,N_22742);
nand U24750 (N_24750,N_23111,N_22830);
and U24751 (N_24751,N_22699,N_23588);
and U24752 (N_24752,N_22605,N_23909);
nand U24753 (N_24753,N_23828,N_22957);
nor U24754 (N_24754,N_23119,N_22780);
nor U24755 (N_24755,N_23879,N_23678);
xor U24756 (N_24756,N_23203,N_23943);
or U24757 (N_24757,N_23872,N_23259);
nand U24758 (N_24758,N_23977,N_23982);
or U24759 (N_24759,N_23054,N_23658);
or U24760 (N_24760,N_23142,N_23123);
and U24761 (N_24761,N_23018,N_22764);
nor U24762 (N_24762,N_22786,N_23958);
or U24763 (N_24763,N_22994,N_23416);
nand U24764 (N_24764,N_23856,N_22691);
nand U24765 (N_24765,N_23197,N_23192);
nor U24766 (N_24766,N_22982,N_23098);
and U24767 (N_24767,N_23538,N_23724);
xnor U24768 (N_24768,N_22972,N_23376);
nand U24769 (N_24769,N_23474,N_23880);
or U24770 (N_24770,N_23042,N_23983);
nor U24771 (N_24771,N_22684,N_23079);
and U24772 (N_24772,N_22969,N_22837);
nand U24773 (N_24773,N_23506,N_23749);
or U24774 (N_24774,N_23156,N_23453);
nand U24775 (N_24775,N_23853,N_23967);
or U24776 (N_24776,N_23425,N_23287);
nand U24777 (N_24777,N_22719,N_23587);
and U24778 (N_24778,N_23347,N_22516);
nand U24779 (N_24779,N_23697,N_23915);
xnor U24780 (N_24780,N_23639,N_23815);
xor U24781 (N_24781,N_23560,N_22989);
xor U24782 (N_24782,N_23056,N_23168);
nor U24783 (N_24783,N_23236,N_23614);
nand U24784 (N_24784,N_23586,N_23552);
nor U24785 (N_24785,N_22668,N_23223);
xor U24786 (N_24786,N_23062,N_23693);
and U24787 (N_24787,N_23008,N_22666);
nand U24788 (N_24788,N_23074,N_22831);
or U24789 (N_24789,N_22639,N_22636);
nand U24790 (N_24790,N_23275,N_23898);
and U24791 (N_24791,N_23742,N_23812);
or U24792 (N_24792,N_22616,N_23777);
xor U24793 (N_24793,N_22772,N_23237);
nand U24794 (N_24794,N_22873,N_22623);
or U24795 (N_24795,N_23222,N_22635);
or U24796 (N_24796,N_22817,N_22568);
or U24797 (N_24797,N_23695,N_22894);
and U24798 (N_24798,N_23366,N_22723);
nor U24799 (N_24799,N_23153,N_22983);
or U24800 (N_24800,N_23409,N_23892);
or U24801 (N_24801,N_23682,N_23933);
nor U24802 (N_24802,N_22906,N_23355);
or U24803 (N_24803,N_23150,N_23897);
nor U24804 (N_24804,N_23929,N_23803);
and U24805 (N_24805,N_22536,N_22547);
or U24806 (N_24806,N_23478,N_22633);
or U24807 (N_24807,N_22634,N_22881);
and U24808 (N_24808,N_23415,N_23840);
nand U24809 (N_24809,N_23872,N_23397);
nor U24810 (N_24810,N_23417,N_23842);
or U24811 (N_24811,N_23041,N_23319);
nand U24812 (N_24812,N_23796,N_22823);
nand U24813 (N_24813,N_23368,N_22812);
or U24814 (N_24814,N_22849,N_23555);
or U24815 (N_24815,N_23946,N_23518);
or U24816 (N_24816,N_23108,N_22823);
nor U24817 (N_24817,N_22894,N_22953);
and U24818 (N_24818,N_23539,N_23278);
nand U24819 (N_24819,N_22536,N_23790);
or U24820 (N_24820,N_23765,N_23883);
nor U24821 (N_24821,N_22915,N_23373);
nor U24822 (N_24822,N_23743,N_23196);
or U24823 (N_24823,N_23039,N_22898);
xnor U24824 (N_24824,N_23416,N_22745);
nand U24825 (N_24825,N_23030,N_23436);
nor U24826 (N_24826,N_23604,N_23069);
xnor U24827 (N_24827,N_23498,N_23884);
nor U24828 (N_24828,N_23885,N_22999);
xor U24829 (N_24829,N_23022,N_22750);
or U24830 (N_24830,N_23086,N_23537);
or U24831 (N_24831,N_22563,N_23447);
xnor U24832 (N_24832,N_23221,N_23232);
nor U24833 (N_24833,N_23511,N_23700);
xnor U24834 (N_24834,N_22670,N_23401);
nor U24835 (N_24835,N_22812,N_23792);
or U24836 (N_24836,N_22537,N_22670);
xnor U24837 (N_24837,N_23670,N_22783);
nand U24838 (N_24838,N_22571,N_23690);
and U24839 (N_24839,N_23250,N_23872);
nand U24840 (N_24840,N_23413,N_23658);
xor U24841 (N_24841,N_23217,N_23958);
nand U24842 (N_24842,N_23232,N_23379);
nor U24843 (N_24843,N_23919,N_22761);
xor U24844 (N_24844,N_22720,N_23198);
or U24845 (N_24845,N_22890,N_23322);
and U24846 (N_24846,N_23522,N_22542);
nand U24847 (N_24847,N_23348,N_23817);
xor U24848 (N_24848,N_22608,N_23532);
nand U24849 (N_24849,N_22808,N_23148);
nor U24850 (N_24850,N_23497,N_23125);
xor U24851 (N_24851,N_23991,N_23669);
nand U24852 (N_24852,N_23321,N_23818);
and U24853 (N_24853,N_23052,N_22735);
nand U24854 (N_24854,N_22817,N_22924);
nand U24855 (N_24855,N_23202,N_22625);
or U24856 (N_24856,N_22507,N_23921);
or U24857 (N_24857,N_23924,N_23970);
nor U24858 (N_24858,N_22917,N_22683);
or U24859 (N_24859,N_22557,N_22503);
or U24860 (N_24860,N_22793,N_22624);
nor U24861 (N_24861,N_23882,N_23371);
and U24862 (N_24862,N_23418,N_22695);
nor U24863 (N_24863,N_22738,N_23035);
xnor U24864 (N_24864,N_23351,N_23652);
or U24865 (N_24865,N_23126,N_23179);
and U24866 (N_24866,N_23684,N_23940);
nor U24867 (N_24867,N_23566,N_23800);
nor U24868 (N_24868,N_22551,N_23752);
nand U24869 (N_24869,N_22664,N_23308);
or U24870 (N_24870,N_22648,N_23515);
or U24871 (N_24871,N_23146,N_23498);
and U24872 (N_24872,N_22500,N_23232);
xor U24873 (N_24873,N_23826,N_23641);
or U24874 (N_24874,N_22604,N_22929);
or U24875 (N_24875,N_22979,N_23631);
or U24876 (N_24876,N_22715,N_23832);
and U24877 (N_24877,N_23126,N_23985);
xnor U24878 (N_24878,N_22784,N_22772);
or U24879 (N_24879,N_22749,N_23561);
nor U24880 (N_24880,N_23521,N_22659);
nand U24881 (N_24881,N_22609,N_23238);
nor U24882 (N_24882,N_23918,N_23855);
nand U24883 (N_24883,N_22718,N_23416);
xnor U24884 (N_24884,N_22905,N_23847);
nand U24885 (N_24885,N_22601,N_22858);
or U24886 (N_24886,N_22702,N_23928);
and U24887 (N_24887,N_23142,N_22743);
xnor U24888 (N_24888,N_23843,N_23550);
nand U24889 (N_24889,N_23548,N_22937);
nor U24890 (N_24890,N_22784,N_23476);
nand U24891 (N_24891,N_23008,N_23012);
nor U24892 (N_24892,N_22723,N_23007);
and U24893 (N_24893,N_23551,N_23266);
or U24894 (N_24894,N_23650,N_23859);
xor U24895 (N_24895,N_23698,N_23848);
nor U24896 (N_24896,N_23821,N_23397);
or U24897 (N_24897,N_23825,N_22613);
nor U24898 (N_24898,N_23727,N_23948);
xnor U24899 (N_24899,N_23171,N_23460);
nand U24900 (N_24900,N_22773,N_23240);
nand U24901 (N_24901,N_23820,N_23899);
or U24902 (N_24902,N_23758,N_23485);
nor U24903 (N_24903,N_22661,N_23078);
or U24904 (N_24904,N_22927,N_23783);
xnor U24905 (N_24905,N_22900,N_23276);
and U24906 (N_24906,N_23051,N_22645);
nand U24907 (N_24907,N_23598,N_23086);
nand U24908 (N_24908,N_22593,N_23832);
or U24909 (N_24909,N_23047,N_23752);
or U24910 (N_24910,N_23780,N_23930);
nand U24911 (N_24911,N_23778,N_23565);
and U24912 (N_24912,N_23578,N_22668);
and U24913 (N_24913,N_23059,N_23448);
xnor U24914 (N_24914,N_23101,N_22622);
nand U24915 (N_24915,N_22752,N_23059);
xor U24916 (N_24916,N_23230,N_22572);
nor U24917 (N_24917,N_23332,N_22540);
nand U24918 (N_24918,N_23039,N_22958);
xnor U24919 (N_24919,N_23755,N_22680);
nor U24920 (N_24920,N_22991,N_22684);
nand U24921 (N_24921,N_23608,N_22893);
xnor U24922 (N_24922,N_23235,N_23590);
nor U24923 (N_24923,N_23249,N_23381);
nor U24924 (N_24924,N_23295,N_23591);
and U24925 (N_24925,N_23765,N_23455);
nand U24926 (N_24926,N_23747,N_23059);
and U24927 (N_24927,N_23304,N_23450);
or U24928 (N_24928,N_23159,N_23378);
and U24929 (N_24929,N_23454,N_22998);
nand U24930 (N_24930,N_22934,N_23514);
nand U24931 (N_24931,N_23844,N_23617);
nor U24932 (N_24932,N_22541,N_22646);
nor U24933 (N_24933,N_22596,N_22569);
or U24934 (N_24934,N_23836,N_23064);
nor U24935 (N_24935,N_23137,N_22811);
xor U24936 (N_24936,N_23123,N_23541);
nor U24937 (N_24937,N_23451,N_22789);
nor U24938 (N_24938,N_23036,N_23103);
nand U24939 (N_24939,N_23057,N_23855);
nor U24940 (N_24940,N_22619,N_22699);
and U24941 (N_24941,N_23125,N_23333);
nand U24942 (N_24942,N_23066,N_23351);
xnor U24943 (N_24943,N_22766,N_23131);
and U24944 (N_24944,N_22502,N_23492);
or U24945 (N_24945,N_22859,N_23453);
or U24946 (N_24946,N_23254,N_22949);
nor U24947 (N_24947,N_23724,N_22858);
xnor U24948 (N_24948,N_22764,N_23040);
nand U24949 (N_24949,N_23682,N_23472);
nor U24950 (N_24950,N_23191,N_23706);
and U24951 (N_24951,N_23586,N_23086);
xnor U24952 (N_24952,N_23881,N_23645);
or U24953 (N_24953,N_23465,N_22590);
or U24954 (N_24954,N_23795,N_23549);
nand U24955 (N_24955,N_22612,N_23763);
xnor U24956 (N_24956,N_23279,N_23516);
xnor U24957 (N_24957,N_22795,N_23453);
and U24958 (N_24958,N_23684,N_22785);
nor U24959 (N_24959,N_22909,N_23760);
and U24960 (N_24960,N_23115,N_22812);
and U24961 (N_24961,N_22948,N_23031);
or U24962 (N_24962,N_23611,N_23688);
and U24963 (N_24963,N_22635,N_22667);
and U24964 (N_24964,N_22760,N_22661);
and U24965 (N_24965,N_22844,N_22586);
nor U24966 (N_24966,N_22951,N_23407);
nand U24967 (N_24967,N_23298,N_23946);
nor U24968 (N_24968,N_22806,N_23744);
nor U24969 (N_24969,N_23449,N_23294);
nand U24970 (N_24970,N_22697,N_23837);
nand U24971 (N_24971,N_23633,N_23882);
or U24972 (N_24972,N_22679,N_22810);
nand U24973 (N_24973,N_23017,N_23339);
nand U24974 (N_24974,N_22936,N_23514);
nand U24975 (N_24975,N_22500,N_22935);
nand U24976 (N_24976,N_23714,N_23753);
and U24977 (N_24977,N_22860,N_23756);
xnor U24978 (N_24978,N_23490,N_23986);
nand U24979 (N_24979,N_22666,N_23690);
or U24980 (N_24980,N_22634,N_23056);
and U24981 (N_24981,N_23340,N_22616);
xor U24982 (N_24982,N_22648,N_22736);
and U24983 (N_24983,N_22537,N_23569);
or U24984 (N_24984,N_23872,N_23374);
nand U24985 (N_24985,N_22548,N_23997);
or U24986 (N_24986,N_23176,N_22722);
nor U24987 (N_24987,N_23330,N_23731);
and U24988 (N_24988,N_23095,N_22836);
xnor U24989 (N_24989,N_23525,N_23571);
xnor U24990 (N_24990,N_23770,N_22631);
nand U24991 (N_24991,N_23597,N_22765);
or U24992 (N_24992,N_23761,N_22727);
nand U24993 (N_24993,N_22887,N_23235);
and U24994 (N_24994,N_23200,N_23403);
and U24995 (N_24995,N_23262,N_23336);
and U24996 (N_24996,N_22553,N_23057);
nor U24997 (N_24997,N_22805,N_23441);
or U24998 (N_24998,N_23605,N_22945);
xnor U24999 (N_24999,N_23704,N_23341);
nor U25000 (N_25000,N_23479,N_23545);
and U25001 (N_25001,N_23895,N_23446);
and U25002 (N_25002,N_23258,N_23883);
nor U25003 (N_25003,N_23539,N_23680);
or U25004 (N_25004,N_22958,N_23774);
and U25005 (N_25005,N_23758,N_22692);
nor U25006 (N_25006,N_23676,N_23402);
or U25007 (N_25007,N_22909,N_23143);
xnor U25008 (N_25008,N_23478,N_23871);
nand U25009 (N_25009,N_23242,N_22643);
xnor U25010 (N_25010,N_23703,N_23970);
nand U25011 (N_25011,N_23788,N_23780);
and U25012 (N_25012,N_22933,N_22814);
nand U25013 (N_25013,N_23505,N_23712);
nor U25014 (N_25014,N_22923,N_22855);
nor U25015 (N_25015,N_22896,N_22580);
xnor U25016 (N_25016,N_23904,N_22613);
and U25017 (N_25017,N_22951,N_22735);
or U25018 (N_25018,N_23457,N_22589);
or U25019 (N_25019,N_22635,N_23630);
xor U25020 (N_25020,N_22778,N_23647);
or U25021 (N_25021,N_22534,N_23559);
and U25022 (N_25022,N_23379,N_23570);
and U25023 (N_25023,N_23961,N_23993);
or U25024 (N_25024,N_23417,N_23125);
nor U25025 (N_25025,N_23295,N_23329);
and U25026 (N_25026,N_23668,N_23271);
nand U25027 (N_25027,N_23760,N_23568);
nor U25028 (N_25028,N_22637,N_22709);
xor U25029 (N_25029,N_23035,N_22584);
nand U25030 (N_25030,N_22685,N_22554);
and U25031 (N_25031,N_22774,N_22843);
nand U25032 (N_25032,N_23345,N_23343);
nor U25033 (N_25033,N_23316,N_22863);
xnor U25034 (N_25034,N_23544,N_22770);
nand U25035 (N_25035,N_23965,N_23197);
nand U25036 (N_25036,N_23162,N_22657);
and U25037 (N_25037,N_23964,N_23546);
and U25038 (N_25038,N_23529,N_22505);
or U25039 (N_25039,N_23874,N_23654);
xnor U25040 (N_25040,N_23844,N_23480);
xor U25041 (N_25041,N_23910,N_22834);
nand U25042 (N_25042,N_23692,N_22552);
and U25043 (N_25043,N_23060,N_22626);
and U25044 (N_25044,N_23966,N_22941);
xor U25045 (N_25045,N_22572,N_22941);
or U25046 (N_25046,N_23246,N_22675);
xor U25047 (N_25047,N_22936,N_23786);
nand U25048 (N_25048,N_23670,N_23832);
or U25049 (N_25049,N_22981,N_23489);
nor U25050 (N_25050,N_23011,N_23952);
and U25051 (N_25051,N_23905,N_23370);
xnor U25052 (N_25052,N_23654,N_23171);
or U25053 (N_25053,N_22706,N_23953);
nand U25054 (N_25054,N_23227,N_23348);
and U25055 (N_25055,N_23902,N_23947);
and U25056 (N_25056,N_23492,N_23937);
nor U25057 (N_25057,N_23318,N_23355);
xor U25058 (N_25058,N_23044,N_22693);
nor U25059 (N_25059,N_23326,N_23022);
xnor U25060 (N_25060,N_23192,N_23656);
nand U25061 (N_25061,N_23925,N_23652);
nor U25062 (N_25062,N_22763,N_23346);
or U25063 (N_25063,N_22559,N_23112);
xor U25064 (N_25064,N_23361,N_23204);
and U25065 (N_25065,N_23165,N_22856);
and U25066 (N_25066,N_23752,N_22662);
or U25067 (N_25067,N_23429,N_23394);
nor U25068 (N_25068,N_22566,N_23799);
nand U25069 (N_25069,N_23297,N_23458);
and U25070 (N_25070,N_22971,N_23999);
nor U25071 (N_25071,N_23068,N_23164);
nand U25072 (N_25072,N_23214,N_23680);
nand U25073 (N_25073,N_23425,N_22909);
xor U25074 (N_25074,N_23886,N_23686);
or U25075 (N_25075,N_23431,N_22814);
xnor U25076 (N_25076,N_22721,N_23770);
xor U25077 (N_25077,N_23643,N_23400);
xor U25078 (N_25078,N_22504,N_22788);
nor U25079 (N_25079,N_22571,N_22671);
or U25080 (N_25080,N_22729,N_23457);
nor U25081 (N_25081,N_23255,N_22523);
nor U25082 (N_25082,N_23937,N_23735);
or U25083 (N_25083,N_23189,N_23036);
or U25084 (N_25084,N_22511,N_22517);
nor U25085 (N_25085,N_22927,N_22678);
or U25086 (N_25086,N_23184,N_23455);
nand U25087 (N_25087,N_22951,N_22717);
and U25088 (N_25088,N_23493,N_23242);
nand U25089 (N_25089,N_23479,N_23331);
nor U25090 (N_25090,N_23540,N_22802);
nand U25091 (N_25091,N_23864,N_23729);
nand U25092 (N_25092,N_22611,N_23225);
or U25093 (N_25093,N_23136,N_23582);
or U25094 (N_25094,N_22834,N_22503);
and U25095 (N_25095,N_22711,N_22734);
and U25096 (N_25096,N_23029,N_23072);
or U25097 (N_25097,N_23577,N_23787);
nand U25098 (N_25098,N_23596,N_22629);
and U25099 (N_25099,N_22754,N_22701);
nor U25100 (N_25100,N_22634,N_23793);
and U25101 (N_25101,N_22949,N_23754);
or U25102 (N_25102,N_23591,N_23661);
or U25103 (N_25103,N_23812,N_23747);
nor U25104 (N_25104,N_22986,N_22884);
nor U25105 (N_25105,N_23424,N_23047);
nor U25106 (N_25106,N_22743,N_23373);
xnor U25107 (N_25107,N_23556,N_23242);
nor U25108 (N_25108,N_22530,N_22710);
or U25109 (N_25109,N_22920,N_23279);
or U25110 (N_25110,N_22588,N_23980);
nor U25111 (N_25111,N_22785,N_22720);
and U25112 (N_25112,N_23877,N_23772);
and U25113 (N_25113,N_22625,N_22947);
nand U25114 (N_25114,N_22877,N_23448);
xor U25115 (N_25115,N_23857,N_22989);
nand U25116 (N_25116,N_23913,N_22563);
and U25117 (N_25117,N_23896,N_23677);
or U25118 (N_25118,N_22588,N_22814);
and U25119 (N_25119,N_23557,N_23913);
nand U25120 (N_25120,N_22514,N_23670);
and U25121 (N_25121,N_23228,N_23157);
nor U25122 (N_25122,N_22729,N_23111);
nor U25123 (N_25123,N_23391,N_22898);
or U25124 (N_25124,N_22730,N_23049);
and U25125 (N_25125,N_23682,N_22815);
xor U25126 (N_25126,N_22623,N_22526);
and U25127 (N_25127,N_22585,N_23563);
or U25128 (N_25128,N_23885,N_23980);
or U25129 (N_25129,N_23510,N_23229);
or U25130 (N_25130,N_22689,N_23403);
or U25131 (N_25131,N_22908,N_22885);
or U25132 (N_25132,N_23245,N_23211);
nor U25133 (N_25133,N_22737,N_23944);
xnor U25134 (N_25134,N_22581,N_23013);
nand U25135 (N_25135,N_23940,N_22881);
xnor U25136 (N_25136,N_22612,N_23899);
and U25137 (N_25137,N_23390,N_22964);
xnor U25138 (N_25138,N_22770,N_22807);
nand U25139 (N_25139,N_23324,N_22698);
nor U25140 (N_25140,N_22753,N_23774);
xnor U25141 (N_25141,N_23883,N_22710);
nor U25142 (N_25142,N_23604,N_23098);
nor U25143 (N_25143,N_23720,N_23478);
or U25144 (N_25144,N_23636,N_22960);
or U25145 (N_25145,N_22822,N_23106);
or U25146 (N_25146,N_23338,N_23615);
nand U25147 (N_25147,N_23643,N_22548);
nand U25148 (N_25148,N_23993,N_22973);
xor U25149 (N_25149,N_23514,N_23281);
and U25150 (N_25150,N_23221,N_23195);
xor U25151 (N_25151,N_22830,N_23443);
xor U25152 (N_25152,N_22634,N_23575);
nor U25153 (N_25153,N_23921,N_23249);
xnor U25154 (N_25154,N_23010,N_23183);
xnor U25155 (N_25155,N_23676,N_22701);
and U25156 (N_25156,N_23485,N_22764);
nor U25157 (N_25157,N_22921,N_23180);
nor U25158 (N_25158,N_23100,N_23615);
nor U25159 (N_25159,N_22674,N_23721);
or U25160 (N_25160,N_23824,N_22590);
and U25161 (N_25161,N_23273,N_23608);
and U25162 (N_25162,N_22959,N_22743);
xor U25163 (N_25163,N_22825,N_23262);
or U25164 (N_25164,N_23286,N_22876);
nor U25165 (N_25165,N_23601,N_23972);
nor U25166 (N_25166,N_22684,N_23319);
nand U25167 (N_25167,N_22740,N_23703);
nor U25168 (N_25168,N_23515,N_23093);
and U25169 (N_25169,N_23824,N_23085);
xnor U25170 (N_25170,N_22998,N_23702);
or U25171 (N_25171,N_23387,N_23001);
and U25172 (N_25172,N_23232,N_23734);
nor U25173 (N_25173,N_22817,N_22915);
or U25174 (N_25174,N_22501,N_22909);
or U25175 (N_25175,N_22744,N_23574);
nand U25176 (N_25176,N_23886,N_23873);
xnor U25177 (N_25177,N_23719,N_22825);
or U25178 (N_25178,N_22825,N_23630);
xor U25179 (N_25179,N_22884,N_23761);
or U25180 (N_25180,N_23794,N_23297);
and U25181 (N_25181,N_22689,N_22560);
nand U25182 (N_25182,N_23154,N_23879);
nor U25183 (N_25183,N_23802,N_23107);
nor U25184 (N_25184,N_23951,N_23735);
nand U25185 (N_25185,N_23138,N_23617);
nand U25186 (N_25186,N_23927,N_22646);
nand U25187 (N_25187,N_22616,N_23189);
xnor U25188 (N_25188,N_22750,N_23261);
and U25189 (N_25189,N_23288,N_23454);
nor U25190 (N_25190,N_23543,N_22747);
nand U25191 (N_25191,N_22941,N_23930);
and U25192 (N_25192,N_22643,N_23192);
and U25193 (N_25193,N_23448,N_22831);
nor U25194 (N_25194,N_23280,N_23487);
or U25195 (N_25195,N_22682,N_23234);
and U25196 (N_25196,N_23741,N_22685);
nand U25197 (N_25197,N_23446,N_22577);
or U25198 (N_25198,N_22626,N_23263);
or U25199 (N_25199,N_23947,N_23866);
nand U25200 (N_25200,N_22817,N_23557);
nand U25201 (N_25201,N_22943,N_22963);
or U25202 (N_25202,N_22616,N_23187);
and U25203 (N_25203,N_23025,N_23068);
xor U25204 (N_25204,N_23909,N_23407);
xor U25205 (N_25205,N_23731,N_22771);
nand U25206 (N_25206,N_23911,N_23147);
xor U25207 (N_25207,N_22573,N_22649);
xor U25208 (N_25208,N_23178,N_23395);
and U25209 (N_25209,N_22988,N_22978);
nor U25210 (N_25210,N_23145,N_23339);
xor U25211 (N_25211,N_22964,N_23313);
nor U25212 (N_25212,N_23934,N_22679);
xor U25213 (N_25213,N_23295,N_22969);
or U25214 (N_25214,N_23974,N_23142);
and U25215 (N_25215,N_22678,N_23838);
and U25216 (N_25216,N_23955,N_23342);
or U25217 (N_25217,N_23656,N_23431);
or U25218 (N_25218,N_22943,N_23070);
nor U25219 (N_25219,N_23472,N_23869);
or U25220 (N_25220,N_23191,N_22796);
nand U25221 (N_25221,N_23596,N_22872);
xor U25222 (N_25222,N_23881,N_23381);
nor U25223 (N_25223,N_23650,N_23078);
nor U25224 (N_25224,N_23792,N_23627);
or U25225 (N_25225,N_22895,N_23394);
xor U25226 (N_25226,N_22614,N_23857);
nand U25227 (N_25227,N_23058,N_23624);
nand U25228 (N_25228,N_22946,N_23308);
nand U25229 (N_25229,N_23398,N_22836);
nor U25230 (N_25230,N_23801,N_23260);
or U25231 (N_25231,N_23091,N_23727);
and U25232 (N_25232,N_23934,N_23618);
xor U25233 (N_25233,N_22855,N_23763);
and U25234 (N_25234,N_22710,N_22760);
nand U25235 (N_25235,N_22622,N_22914);
xor U25236 (N_25236,N_22768,N_22812);
nor U25237 (N_25237,N_22742,N_23883);
nand U25238 (N_25238,N_23272,N_22631);
nor U25239 (N_25239,N_23045,N_23437);
nand U25240 (N_25240,N_23049,N_22824);
nand U25241 (N_25241,N_23391,N_23963);
and U25242 (N_25242,N_23328,N_23192);
nand U25243 (N_25243,N_23838,N_22996);
nand U25244 (N_25244,N_23692,N_23012);
nand U25245 (N_25245,N_23297,N_23329);
and U25246 (N_25246,N_22555,N_23994);
or U25247 (N_25247,N_23487,N_22823);
or U25248 (N_25248,N_23886,N_23277);
nand U25249 (N_25249,N_23545,N_23484);
nor U25250 (N_25250,N_23836,N_23477);
and U25251 (N_25251,N_23646,N_23960);
or U25252 (N_25252,N_23377,N_23655);
xnor U25253 (N_25253,N_23509,N_23031);
nor U25254 (N_25254,N_22610,N_23403);
or U25255 (N_25255,N_23742,N_23567);
nor U25256 (N_25256,N_23899,N_23602);
nor U25257 (N_25257,N_22758,N_23888);
nand U25258 (N_25258,N_22951,N_23901);
nand U25259 (N_25259,N_23752,N_22564);
and U25260 (N_25260,N_22607,N_23427);
nor U25261 (N_25261,N_23412,N_23683);
and U25262 (N_25262,N_23634,N_23797);
xor U25263 (N_25263,N_22729,N_23844);
nor U25264 (N_25264,N_22648,N_23641);
nor U25265 (N_25265,N_23843,N_22559);
nor U25266 (N_25266,N_23500,N_22504);
nand U25267 (N_25267,N_23304,N_23931);
and U25268 (N_25268,N_22934,N_23624);
nor U25269 (N_25269,N_22623,N_22604);
or U25270 (N_25270,N_23618,N_23410);
nor U25271 (N_25271,N_23618,N_23125);
nand U25272 (N_25272,N_23106,N_23016);
nor U25273 (N_25273,N_23201,N_23672);
and U25274 (N_25274,N_23298,N_23008);
and U25275 (N_25275,N_22615,N_23837);
nor U25276 (N_25276,N_23405,N_23838);
nand U25277 (N_25277,N_23696,N_23158);
nand U25278 (N_25278,N_23542,N_22815);
and U25279 (N_25279,N_23922,N_23508);
nor U25280 (N_25280,N_22999,N_22559);
or U25281 (N_25281,N_22869,N_22582);
xor U25282 (N_25282,N_23323,N_23634);
nor U25283 (N_25283,N_23795,N_23606);
nor U25284 (N_25284,N_23142,N_22689);
or U25285 (N_25285,N_22924,N_23297);
nor U25286 (N_25286,N_22729,N_23405);
or U25287 (N_25287,N_23201,N_22665);
xnor U25288 (N_25288,N_22593,N_23251);
and U25289 (N_25289,N_23038,N_23291);
nand U25290 (N_25290,N_22989,N_22610);
or U25291 (N_25291,N_23414,N_23768);
xor U25292 (N_25292,N_22501,N_23877);
and U25293 (N_25293,N_22852,N_23651);
or U25294 (N_25294,N_23526,N_23173);
nor U25295 (N_25295,N_22786,N_23523);
or U25296 (N_25296,N_23012,N_23860);
or U25297 (N_25297,N_22758,N_23932);
nor U25298 (N_25298,N_23128,N_23311);
or U25299 (N_25299,N_22895,N_23528);
xor U25300 (N_25300,N_23457,N_23410);
and U25301 (N_25301,N_23948,N_23693);
nand U25302 (N_25302,N_22906,N_23386);
and U25303 (N_25303,N_23888,N_23386);
xor U25304 (N_25304,N_23414,N_23079);
nor U25305 (N_25305,N_23799,N_23637);
nor U25306 (N_25306,N_23794,N_22533);
nor U25307 (N_25307,N_23896,N_23914);
or U25308 (N_25308,N_23257,N_22746);
xor U25309 (N_25309,N_23917,N_23927);
nand U25310 (N_25310,N_23870,N_23571);
nor U25311 (N_25311,N_22668,N_23862);
xnor U25312 (N_25312,N_23782,N_22962);
and U25313 (N_25313,N_23477,N_23571);
or U25314 (N_25314,N_23263,N_22902);
nor U25315 (N_25315,N_22522,N_23596);
nand U25316 (N_25316,N_23094,N_23723);
and U25317 (N_25317,N_23190,N_23917);
xor U25318 (N_25318,N_22822,N_22989);
nor U25319 (N_25319,N_23406,N_22511);
or U25320 (N_25320,N_22926,N_23738);
xnor U25321 (N_25321,N_23722,N_22593);
nand U25322 (N_25322,N_23737,N_22563);
xnor U25323 (N_25323,N_23257,N_22926);
or U25324 (N_25324,N_23250,N_23601);
and U25325 (N_25325,N_23022,N_22628);
xor U25326 (N_25326,N_23622,N_23477);
or U25327 (N_25327,N_22844,N_23865);
or U25328 (N_25328,N_23615,N_22862);
xnor U25329 (N_25329,N_22967,N_22842);
and U25330 (N_25330,N_22556,N_23560);
nor U25331 (N_25331,N_22999,N_23768);
or U25332 (N_25332,N_23872,N_23362);
or U25333 (N_25333,N_22954,N_22882);
or U25334 (N_25334,N_23212,N_23304);
nand U25335 (N_25335,N_22577,N_23525);
and U25336 (N_25336,N_22983,N_23342);
and U25337 (N_25337,N_23427,N_23154);
and U25338 (N_25338,N_22768,N_23603);
nand U25339 (N_25339,N_23406,N_22597);
and U25340 (N_25340,N_22613,N_23658);
nand U25341 (N_25341,N_23352,N_22901);
xor U25342 (N_25342,N_23943,N_22939);
nand U25343 (N_25343,N_23214,N_22646);
and U25344 (N_25344,N_23774,N_22647);
nor U25345 (N_25345,N_23314,N_23764);
xor U25346 (N_25346,N_23653,N_23453);
nor U25347 (N_25347,N_23852,N_22684);
or U25348 (N_25348,N_23429,N_22898);
xor U25349 (N_25349,N_23668,N_22859);
nor U25350 (N_25350,N_22675,N_23724);
nor U25351 (N_25351,N_22779,N_22503);
or U25352 (N_25352,N_23457,N_23602);
xor U25353 (N_25353,N_23549,N_23007);
nor U25354 (N_25354,N_22921,N_23843);
nand U25355 (N_25355,N_22516,N_23310);
or U25356 (N_25356,N_23753,N_22502);
xor U25357 (N_25357,N_22505,N_23271);
or U25358 (N_25358,N_22722,N_23495);
and U25359 (N_25359,N_23339,N_23713);
nor U25360 (N_25360,N_23705,N_23981);
xor U25361 (N_25361,N_23493,N_23420);
and U25362 (N_25362,N_23669,N_23215);
nand U25363 (N_25363,N_22732,N_22660);
nor U25364 (N_25364,N_23178,N_23771);
nand U25365 (N_25365,N_23334,N_22881);
or U25366 (N_25366,N_23384,N_22574);
and U25367 (N_25367,N_22865,N_23176);
and U25368 (N_25368,N_22640,N_23828);
nand U25369 (N_25369,N_23471,N_23814);
or U25370 (N_25370,N_22507,N_23769);
xnor U25371 (N_25371,N_23624,N_22786);
nor U25372 (N_25372,N_22578,N_23498);
nand U25373 (N_25373,N_22998,N_22542);
and U25374 (N_25374,N_23790,N_23063);
and U25375 (N_25375,N_22918,N_23613);
or U25376 (N_25376,N_22940,N_22843);
or U25377 (N_25377,N_23283,N_23150);
xor U25378 (N_25378,N_23536,N_23642);
and U25379 (N_25379,N_22807,N_22998);
nor U25380 (N_25380,N_23766,N_22549);
or U25381 (N_25381,N_23396,N_22981);
nand U25382 (N_25382,N_23442,N_23934);
nand U25383 (N_25383,N_23442,N_23333);
nor U25384 (N_25384,N_23074,N_23460);
and U25385 (N_25385,N_23190,N_23784);
xnor U25386 (N_25386,N_23452,N_23642);
nand U25387 (N_25387,N_23272,N_23474);
or U25388 (N_25388,N_23594,N_23039);
and U25389 (N_25389,N_23274,N_22862);
nor U25390 (N_25390,N_22735,N_23617);
nor U25391 (N_25391,N_23486,N_23325);
nand U25392 (N_25392,N_22504,N_23064);
xor U25393 (N_25393,N_22516,N_23755);
nand U25394 (N_25394,N_22930,N_22936);
nor U25395 (N_25395,N_23668,N_22679);
nor U25396 (N_25396,N_23761,N_23959);
xor U25397 (N_25397,N_23263,N_22725);
nor U25398 (N_25398,N_22830,N_23672);
nand U25399 (N_25399,N_23138,N_23307);
nand U25400 (N_25400,N_22632,N_23518);
nor U25401 (N_25401,N_23757,N_23991);
or U25402 (N_25402,N_23849,N_22941);
and U25403 (N_25403,N_23266,N_22967);
or U25404 (N_25404,N_23941,N_22863);
and U25405 (N_25405,N_23886,N_23791);
nor U25406 (N_25406,N_22685,N_23690);
xor U25407 (N_25407,N_22903,N_22747);
nor U25408 (N_25408,N_23564,N_22854);
or U25409 (N_25409,N_22720,N_22886);
nand U25410 (N_25410,N_22643,N_23844);
xnor U25411 (N_25411,N_23851,N_23132);
and U25412 (N_25412,N_23390,N_23961);
nand U25413 (N_25413,N_22632,N_22842);
nor U25414 (N_25414,N_22682,N_23429);
nand U25415 (N_25415,N_22545,N_22565);
and U25416 (N_25416,N_23534,N_23278);
nand U25417 (N_25417,N_23295,N_23034);
xor U25418 (N_25418,N_23070,N_23465);
nor U25419 (N_25419,N_23197,N_22946);
nor U25420 (N_25420,N_22741,N_22993);
nand U25421 (N_25421,N_23644,N_23765);
nor U25422 (N_25422,N_22683,N_23764);
and U25423 (N_25423,N_22587,N_22588);
or U25424 (N_25424,N_22711,N_23416);
xor U25425 (N_25425,N_23468,N_23628);
nand U25426 (N_25426,N_22917,N_23572);
xnor U25427 (N_25427,N_23787,N_23698);
nor U25428 (N_25428,N_23269,N_22540);
nand U25429 (N_25429,N_23379,N_22698);
or U25430 (N_25430,N_23366,N_23669);
and U25431 (N_25431,N_22565,N_23484);
nand U25432 (N_25432,N_23504,N_22894);
nor U25433 (N_25433,N_22717,N_22931);
xor U25434 (N_25434,N_23551,N_22903);
nand U25435 (N_25435,N_23561,N_23414);
nor U25436 (N_25436,N_23607,N_23385);
nor U25437 (N_25437,N_22938,N_23833);
or U25438 (N_25438,N_22898,N_22804);
nor U25439 (N_25439,N_23907,N_23028);
nor U25440 (N_25440,N_23666,N_23447);
xor U25441 (N_25441,N_23805,N_22746);
nand U25442 (N_25442,N_22904,N_23545);
or U25443 (N_25443,N_22636,N_23776);
and U25444 (N_25444,N_23945,N_23169);
xor U25445 (N_25445,N_23659,N_22579);
or U25446 (N_25446,N_23617,N_22925);
and U25447 (N_25447,N_23105,N_22531);
nand U25448 (N_25448,N_22950,N_22811);
and U25449 (N_25449,N_22507,N_23419);
and U25450 (N_25450,N_22580,N_23426);
and U25451 (N_25451,N_23241,N_23328);
xnor U25452 (N_25452,N_22954,N_22867);
nand U25453 (N_25453,N_23939,N_23523);
xnor U25454 (N_25454,N_23385,N_23714);
or U25455 (N_25455,N_23268,N_23918);
and U25456 (N_25456,N_23504,N_23509);
nor U25457 (N_25457,N_23410,N_22888);
nor U25458 (N_25458,N_23223,N_23813);
and U25459 (N_25459,N_23655,N_22909);
nor U25460 (N_25460,N_23560,N_23433);
and U25461 (N_25461,N_22932,N_23105);
nor U25462 (N_25462,N_22561,N_23614);
xnor U25463 (N_25463,N_23999,N_22742);
nand U25464 (N_25464,N_23901,N_23370);
and U25465 (N_25465,N_23658,N_23908);
nand U25466 (N_25466,N_23250,N_22869);
nor U25467 (N_25467,N_23852,N_23700);
or U25468 (N_25468,N_23748,N_23689);
and U25469 (N_25469,N_23413,N_23799);
nor U25470 (N_25470,N_23118,N_22996);
or U25471 (N_25471,N_22865,N_23635);
nand U25472 (N_25472,N_23520,N_23488);
nor U25473 (N_25473,N_23576,N_23531);
nand U25474 (N_25474,N_23905,N_23757);
nand U25475 (N_25475,N_22749,N_23570);
nand U25476 (N_25476,N_23758,N_23913);
or U25477 (N_25477,N_23032,N_22799);
and U25478 (N_25478,N_23124,N_23951);
nand U25479 (N_25479,N_23724,N_22835);
nand U25480 (N_25480,N_23339,N_23334);
xnor U25481 (N_25481,N_22608,N_23786);
nor U25482 (N_25482,N_23012,N_22983);
nand U25483 (N_25483,N_23506,N_23889);
and U25484 (N_25484,N_23244,N_22753);
nor U25485 (N_25485,N_23100,N_23214);
nand U25486 (N_25486,N_23337,N_23268);
xor U25487 (N_25487,N_22619,N_23901);
xor U25488 (N_25488,N_23354,N_23579);
nor U25489 (N_25489,N_22717,N_22712);
nor U25490 (N_25490,N_22908,N_23172);
xor U25491 (N_25491,N_23733,N_22841);
nor U25492 (N_25492,N_22613,N_22951);
nand U25493 (N_25493,N_23364,N_22969);
xnor U25494 (N_25494,N_23706,N_23629);
nand U25495 (N_25495,N_23677,N_23260);
and U25496 (N_25496,N_23913,N_22501);
nand U25497 (N_25497,N_22504,N_23759);
and U25498 (N_25498,N_23495,N_22779);
xnor U25499 (N_25499,N_23323,N_23236);
xor U25500 (N_25500,N_24902,N_24247);
or U25501 (N_25501,N_24613,N_25491);
nor U25502 (N_25502,N_24366,N_24005);
nand U25503 (N_25503,N_24768,N_24587);
nand U25504 (N_25504,N_24228,N_24173);
nand U25505 (N_25505,N_24614,N_24475);
or U25506 (N_25506,N_25441,N_24594);
or U25507 (N_25507,N_24822,N_24314);
nor U25508 (N_25508,N_24239,N_25149);
nor U25509 (N_25509,N_25367,N_24607);
or U25510 (N_25510,N_24726,N_25004);
or U25511 (N_25511,N_24604,N_25237);
or U25512 (N_25512,N_24263,N_24036);
nor U25513 (N_25513,N_25225,N_25317);
xnor U25514 (N_25514,N_24227,N_25482);
nand U25515 (N_25515,N_24689,N_24825);
nor U25516 (N_25516,N_25239,N_24723);
or U25517 (N_25517,N_25354,N_25002);
xnor U25518 (N_25518,N_24528,N_25226);
and U25519 (N_25519,N_25276,N_24801);
or U25520 (N_25520,N_25139,N_24894);
or U25521 (N_25521,N_24596,N_24017);
and U25522 (N_25522,N_24570,N_24013);
nor U25523 (N_25523,N_24750,N_24312);
nand U25524 (N_25524,N_24051,N_24905);
and U25525 (N_25525,N_24221,N_24123);
or U25526 (N_25526,N_25471,N_24110);
nand U25527 (N_25527,N_25403,N_24050);
nand U25528 (N_25528,N_24413,N_24521);
or U25529 (N_25529,N_24302,N_24915);
and U25530 (N_25530,N_24313,N_24569);
and U25531 (N_25531,N_24283,N_25171);
or U25532 (N_25532,N_24715,N_24298);
or U25533 (N_25533,N_24037,N_24149);
and U25534 (N_25534,N_25241,N_25425);
or U25535 (N_25535,N_24015,N_25386);
or U25536 (N_25536,N_24682,N_24972);
and U25537 (N_25537,N_24943,N_25447);
or U25538 (N_25538,N_24864,N_25153);
or U25539 (N_25539,N_24400,N_25359);
or U25540 (N_25540,N_24897,N_24002);
or U25541 (N_25541,N_24078,N_24277);
and U25542 (N_25542,N_24006,N_24291);
or U25543 (N_25543,N_25169,N_24875);
xor U25544 (N_25544,N_24793,N_24877);
nor U25545 (N_25545,N_24202,N_24821);
xnor U25546 (N_25546,N_25486,N_25434);
xnor U25547 (N_25547,N_24159,N_24270);
nor U25548 (N_25548,N_25093,N_24987);
nand U25549 (N_25549,N_24764,N_25026);
nor U25550 (N_25550,N_25019,N_24549);
xnor U25551 (N_25551,N_24395,N_25244);
nand U25552 (N_25552,N_24959,N_24072);
nor U25553 (N_25553,N_24354,N_24059);
nor U25554 (N_25554,N_24303,N_25389);
nand U25555 (N_25555,N_24345,N_24572);
nor U25556 (N_25556,N_25096,N_24847);
nor U25557 (N_25557,N_24486,N_25055);
nand U25558 (N_25558,N_24115,N_24082);
nor U25559 (N_25559,N_24522,N_24222);
or U25560 (N_25560,N_25206,N_25105);
xor U25561 (N_25561,N_25436,N_25017);
nor U25562 (N_25562,N_25191,N_25373);
and U25563 (N_25563,N_25208,N_24608);
nand U25564 (N_25564,N_24329,N_24212);
nand U25565 (N_25565,N_25051,N_24375);
nor U25566 (N_25566,N_25082,N_25448);
xor U25567 (N_25567,N_24249,N_25438);
and U25568 (N_25568,N_24139,N_24242);
nor U25569 (N_25569,N_25188,N_24049);
nor U25570 (N_25570,N_24069,N_24169);
nor U25571 (N_25571,N_24204,N_25463);
nand U25572 (N_25572,N_24516,N_24941);
nand U25573 (N_25573,N_24198,N_25047);
xnor U25574 (N_25574,N_25284,N_25492);
nand U25575 (N_25575,N_24033,N_25267);
or U25576 (N_25576,N_24349,N_24925);
xnor U25577 (N_25577,N_24372,N_24307);
xor U25578 (N_25578,N_24290,N_25398);
or U25579 (N_25579,N_24956,N_24097);
or U25580 (N_25580,N_24145,N_24885);
nor U25581 (N_25581,N_24863,N_24304);
nand U25582 (N_25582,N_24034,N_25077);
xnor U25583 (N_25583,N_25461,N_25134);
xnor U25584 (N_25584,N_25053,N_25074);
xor U25585 (N_25585,N_24610,N_24288);
xor U25586 (N_25586,N_24188,N_24416);
nor U25587 (N_25587,N_25102,N_24621);
and U25588 (N_25588,N_24189,N_25196);
nand U25589 (N_25589,N_24735,N_25407);
or U25590 (N_25590,N_25397,N_24510);
nor U25591 (N_25591,N_24359,N_24965);
or U25592 (N_25592,N_24612,N_24886);
and U25593 (N_25593,N_24519,N_25415);
and U25594 (N_25594,N_24167,N_24022);
xnor U25595 (N_25595,N_25370,N_25469);
and U25596 (N_25596,N_24710,N_25394);
and U25597 (N_25597,N_24357,N_25285);
and U25598 (N_25598,N_24857,N_25148);
or U25599 (N_25599,N_25100,N_24409);
or U25600 (N_25600,N_24784,N_24271);
and U25601 (N_25601,N_24624,N_25307);
or U25602 (N_25602,N_24152,N_25335);
xnor U25603 (N_25603,N_25057,N_24296);
or U25604 (N_25604,N_25104,N_24437);
nand U25605 (N_25605,N_24250,N_24999);
nand U25606 (N_25606,N_24282,N_24500);
xor U25607 (N_25607,N_24564,N_24674);
or U25608 (N_25608,N_25121,N_25003);
nor U25609 (N_25609,N_25301,N_24720);
and U25610 (N_25610,N_24812,N_25065);
and U25611 (N_25611,N_25315,N_25266);
nand U25612 (N_25612,N_25137,N_24356);
nand U25613 (N_25613,N_25443,N_24912);
nand U25614 (N_25614,N_24984,N_24490);
or U25615 (N_25615,N_25119,N_24224);
nor U25616 (N_25616,N_24402,N_24526);
nor U25617 (N_25617,N_24868,N_24969);
and U25618 (N_25618,N_24316,N_24178);
nand U25619 (N_25619,N_25323,N_25162);
and U25620 (N_25620,N_24806,N_24141);
xor U25621 (N_25621,N_24796,N_25110);
or U25622 (N_25622,N_24335,N_24245);
xnor U25623 (N_25623,N_24974,N_24916);
and U25624 (N_25624,N_24162,N_25193);
nand U25625 (N_25625,N_25311,N_25361);
nor U25626 (N_25626,N_25495,N_25336);
xnor U25627 (N_25627,N_24997,N_24117);
nor U25628 (N_25628,N_24603,N_24620);
xor U25629 (N_25629,N_24182,N_24834);
nand U25630 (N_25630,N_24636,N_24708);
xnor U25631 (N_25631,N_24071,N_24681);
and U25632 (N_25632,N_25108,N_25280);
nand U25633 (N_25633,N_24904,N_24127);
nor U25634 (N_25634,N_25473,N_25073);
nand U25635 (N_25635,N_24255,N_24087);
and U25636 (N_25636,N_24830,N_25001);
xnor U25637 (N_25637,N_24124,N_24991);
or U25638 (N_25638,N_25218,N_24370);
nor U25639 (N_25639,N_24581,N_25247);
or U25640 (N_25640,N_24794,N_24733);
nor U25641 (N_25641,N_25063,N_25458);
or U25642 (N_25642,N_25418,N_24090);
xnor U25643 (N_25643,N_25046,N_24898);
nand U25644 (N_25644,N_24404,N_25249);
xor U25645 (N_25645,N_24241,N_25221);
nand U25646 (N_25646,N_24927,N_24389);
xor U25647 (N_25647,N_24120,N_24958);
xor U25648 (N_25648,N_24839,N_25422);
nor U25649 (N_25649,N_24257,N_24197);
nand U25650 (N_25650,N_24836,N_24161);
nor U25651 (N_25651,N_24089,N_24718);
xnor U25652 (N_25652,N_24583,N_25352);
and U25653 (N_25653,N_24626,N_24252);
and U25654 (N_25654,N_24320,N_24448);
and U25655 (N_25655,N_24042,N_24088);
nor U25656 (N_25656,N_24405,N_24445);
xnor U25657 (N_25657,N_24333,N_24158);
nand U25658 (N_25658,N_24895,N_25168);
xor U25659 (N_25659,N_25433,N_24685);
or U25660 (N_25660,N_24632,N_24164);
and U25661 (N_25661,N_24003,N_24651);
nor U25662 (N_25662,N_24129,N_24163);
or U25663 (N_25663,N_24176,N_24440);
and U25664 (N_25664,N_25111,N_24668);
nor U25665 (N_25665,N_24630,N_24012);
nand U25666 (N_25666,N_25459,N_24929);
xor U25667 (N_25667,N_24766,N_24248);
xnor U25668 (N_25668,N_24433,N_25204);
or U25669 (N_25669,N_25303,N_25449);
xor U25670 (N_25670,N_24827,N_24695);
nand U25671 (N_25671,N_24213,N_24508);
and U25672 (N_25672,N_25405,N_24584);
or U25673 (N_25673,N_25031,N_25250);
nor U25674 (N_25674,N_24432,N_24231);
or U25675 (N_25675,N_24496,N_24253);
nand U25676 (N_25676,N_24175,N_25091);
xor U25677 (N_25677,N_24492,N_24442);
or U25678 (N_25678,N_24394,N_24845);
nor U25679 (N_25679,N_24443,N_25258);
nand U25680 (N_25680,N_25498,N_24215);
or U25681 (N_25681,N_24488,N_25291);
nand U25682 (N_25682,N_24779,N_24858);
nand U25683 (N_25683,N_24846,N_24172);
or U25684 (N_25684,N_25444,N_24007);
xnor U25685 (N_25685,N_24406,N_25076);
nor U25686 (N_25686,N_24616,N_25275);
nand U25687 (N_25687,N_24371,N_25480);
or U25688 (N_25688,N_25020,N_24048);
or U25689 (N_25689,N_24324,N_25177);
nor U25690 (N_25690,N_24435,N_24452);
and U25691 (N_25691,N_24226,N_24770);
xnor U25692 (N_25692,N_24073,N_24053);
nor U25693 (N_25693,N_25150,N_24949);
or U25694 (N_25694,N_24504,N_24571);
or U25695 (N_25695,N_24344,N_25342);
or U25696 (N_25696,N_24899,N_24415);
and U25697 (N_25697,N_24016,N_24111);
nor U25698 (N_25698,N_25279,N_24989);
or U25699 (N_25699,N_24837,N_25437);
nor U25700 (N_25700,N_24524,N_24514);
nor U25701 (N_25701,N_25287,N_24737);
nor U25702 (N_25702,N_24538,N_24031);
or U25703 (N_25703,N_24701,N_24852);
or U25704 (N_25704,N_24299,N_25489);
and U25705 (N_25705,N_25015,N_25261);
xnor U25706 (N_25706,N_25264,N_24932);
xnor U25707 (N_25707,N_24700,N_24833);
xnor U25708 (N_25708,N_25322,N_25494);
nand U25709 (N_25709,N_25138,N_24946);
nor U25710 (N_25710,N_24364,N_24600);
or U25711 (N_25711,N_24536,N_24154);
nand U25712 (N_25712,N_24489,N_24038);
xor U25713 (N_25713,N_24605,N_24382);
nor U25714 (N_25714,N_24166,N_24367);
nand U25715 (N_25715,N_24456,N_25045);
or U25716 (N_25716,N_24758,N_24635);
xnor U25717 (N_25717,N_24629,N_25292);
and U25718 (N_25718,N_24119,N_24975);
or U25719 (N_25719,N_25114,N_24434);
xor U25720 (N_25720,N_25120,N_24558);
nand U25721 (N_25721,N_24575,N_24933);
xnor U25722 (N_25722,N_25224,N_24641);
nand U25723 (N_25723,N_24799,N_25348);
or U25724 (N_25724,N_25088,N_24921);
and U25725 (N_25725,N_25470,N_24000);
nand U25726 (N_25726,N_25347,N_24196);
and U25727 (N_25727,N_24297,N_25211);
and U25728 (N_25728,N_25214,N_25205);
nand U25729 (N_25729,N_25126,N_24289);
and U25730 (N_25730,N_24191,N_24543);
nand U25731 (N_25731,N_24148,N_24655);
nor U25732 (N_25732,N_24118,N_24384);
nor U25733 (N_25733,N_24891,N_24961);
or U25734 (N_25734,N_24431,N_25079);
and U25735 (N_25735,N_25337,N_25421);
and U25736 (N_25736,N_24346,N_24547);
nor U25737 (N_25737,N_25351,N_25265);
and U25738 (N_25738,N_24754,N_25310);
and U25739 (N_25739,N_25064,N_24745);
nor U25740 (N_25740,N_24906,N_25253);
or U25741 (N_25741,N_24294,N_24983);
nand U25742 (N_25742,N_24803,N_24368);
nor U25743 (N_25743,N_24066,N_24043);
and U25744 (N_25744,N_25460,N_24676);
xor U25745 (N_25745,N_25339,N_24944);
nor U25746 (N_25746,N_25278,N_24537);
or U25747 (N_25747,N_25399,N_24950);
or U25748 (N_25748,N_24460,N_24646);
or U25749 (N_25749,N_24968,N_24347);
nor U25750 (N_25750,N_25081,N_24187);
and U25751 (N_25751,N_24499,N_24186);
xor U25752 (N_25752,N_24308,N_24782);
xnor U25753 (N_25753,N_24153,N_24407);
or U25754 (N_25754,N_25462,N_24512);
and U25755 (N_25755,N_24530,N_24267);
or U25756 (N_25756,N_24387,N_24062);
or U25757 (N_25757,N_24041,N_24540);
or U25758 (N_25758,N_24234,N_25029);
xnor U25759 (N_25759,N_25455,N_24840);
or U25760 (N_25760,N_25268,N_24218);
nand U25761 (N_25761,N_24468,N_24391);
nor U25762 (N_25762,N_24235,N_24731);
xnor U25763 (N_25763,N_25036,N_24686);
nor U25764 (N_25764,N_24890,N_25419);
nor U25765 (N_25765,N_24108,N_24986);
nor U25766 (N_25766,N_25487,N_24461);
and U25767 (N_25767,N_24467,N_24479);
and U25768 (N_25768,N_24619,N_24931);
xnor U25769 (N_25769,N_25199,N_25383);
or U25770 (N_25770,N_24820,N_24882);
xor U25771 (N_25771,N_24523,N_24692);
xor U25772 (N_25772,N_25230,N_25097);
and U25773 (N_25773,N_24714,N_24918);
or U25774 (N_25774,N_24278,N_24694);
nand U25775 (N_25775,N_24755,N_24075);
nor U25776 (N_25776,N_24014,N_24397);
nor U25777 (N_25777,N_25408,N_24470);
or U25778 (N_25778,N_24533,N_25167);
or U25779 (N_25779,N_24653,N_25028);
nand U25780 (N_25780,N_24137,N_24942);
or U25781 (N_25781,N_25228,N_24011);
and U25782 (N_25782,N_25067,N_24428);
or U25783 (N_25783,N_25166,N_25016);
nand U25784 (N_25784,N_24493,N_24903);
xnor U25785 (N_25785,N_24205,N_24896);
xor U25786 (N_25786,N_25009,N_24408);
xor U25787 (N_25787,N_24322,N_25164);
nor U25788 (N_25788,N_24763,N_25172);
nand U25789 (N_25789,N_24207,N_24615);
and U25790 (N_25790,N_24595,N_24552);
and U25791 (N_25791,N_25333,N_24502);
nand U25792 (N_25792,N_24273,N_24414);
and U25793 (N_25793,N_24562,N_24990);
nor U25794 (N_25794,N_24458,N_25037);
nor U25795 (N_25795,N_24705,N_24658);
xor U25796 (N_25796,N_25184,N_24568);
and U25797 (N_25797,N_24805,N_24759);
xor U25798 (N_25798,N_24819,N_24480);
or U25799 (N_25799,N_24647,N_24797);
xnor U25800 (N_25800,N_24995,N_25005);
nand U25801 (N_25801,N_24168,N_24450);
nand U25802 (N_25802,N_24696,N_25217);
and U25803 (N_25803,N_25018,N_25417);
or U25804 (N_25804,N_24369,N_25136);
or U25805 (N_25805,N_25158,N_24112);
and U25806 (N_25806,N_25227,N_25238);
xor U25807 (N_25807,N_24725,N_25042);
and U25808 (N_25808,N_24661,N_25198);
or U25809 (N_25809,N_25201,N_25320);
and U25810 (N_25810,N_24743,N_25318);
nand U25811 (N_25811,N_25451,N_24832);
and U25812 (N_25812,N_24665,N_24871);
or U25813 (N_25813,N_24085,N_24874);
xnor U25814 (N_25814,N_24240,N_25179);
nand U25815 (N_25815,N_25187,N_24441);
xor U25816 (N_25816,N_24976,N_25220);
nand U25817 (N_25817,N_24272,N_25393);
nor U25818 (N_25818,N_25127,N_24702);
nor U25819 (N_25819,N_24261,N_24876);
and U25820 (N_25820,N_24285,N_24854);
xor U25821 (N_25821,N_24515,N_24449);
and U25822 (N_25822,N_24068,N_24527);
nor U25823 (N_25823,N_24671,N_25334);
nand U25824 (N_25824,N_24749,N_25412);
and U25825 (N_25825,N_25061,N_24800);
xor U25826 (N_25826,N_25115,N_25445);
and U25827 (N_25827,N_24555,N_25007);
xnor U25828 (N_25828,N_24559,N_24849);
nor U25829 (N_25829,N_24951,N_24057);
nor U25830 (N_25830,N_24194,N_25066);
nor U25831 (N_25831,N_24778,N_24340);
or U25832 (N_25832,N_25080,N_24517);
or U25833 (N_25833,N_25474,N_24269);
or U25834 (N_25834,N_24791,N_24330);
xnor U25835 (N_25835,N_24459,N_24505);
nor U25836 (N_25836,N_24734,N_24520);
nand U25837 (N_25837,N_25014,N_24170);
and U25838 (N_25838,N_24473,N_24699);
or U25839 (N_25839,N_24729,N_24979);
nor U25840 (N_25840,N_25068,N_24396);
and U25841 (N_25841,N_24177,N_24327);
and U25842 (N_25842,N_24638,N_24730);
or U25843 (N_25843,N_25160,N_25295);
or U25844 (N_25844,N_25197,N_24548);
and U25845 (N_25845,N_25161,N_24421);
xor U25846 (N_25846,N_24645,N_24663);
or U25847 (N_25847,N_25476,N_24541);
and U25848 (N_25848,N_25453,N_24465);
xnor U25849 (N_25849,N_24598,N_24236);
nand U25850 (N_25850,N_24940,N_25212);
xor U25851 (N_25851,N_25475,N_24219);
nor U25852 (N_25852,N_24660,N_25270);
nor U25853 (N_25853,N_25147,N_25380);
xor U25854 (N_25854,N_24566,N_24055);
and U25855 (N_25855,N_24776,N_24666);
nand U25856 (N_25856,N_25376,N_24728);
nand U25857 (N_25857,N_24009,N_25098);
nand U25858 (N_25858,N_24321,N_25092);
or U25859 (N_25859,N_25194,N_24567);
nand U25860 (N_25860,N_25113,N_24029);
or U25861 (N_25861,N_25086,N_25173);
and U25862 (N_25862,N_24265,N_25229);
or U25863 (N_25863,N_24544,N_24982);
nand U25864 (N_25864,N_24310,N_25277);
nor U25865 (N_25865,N_25085,N_24266);
or U25866 (N_25866,N_25039,N_25331);
and U25867 (N_25867,N_24008,N_25499);
nand U25868 (N_25868,N_24004,N_24865);
or U25869 (N_25869,N_24789,N_25246);
nor U25870 (N_25870,N_24657,N_24293);
and U25871 (N_25871,N_24936,N_24040);
nor U25872 (N_25872,N_24080,N_24334);
or U25873 (N_25873,N_25360,N_24383);
nand U25874 (N_25874,N_25181,N_24351);
and U25875 (N_25875,N_24061,N_25000);
and U25876 (N_25876,N_25377,N_25349);
xor U25877 (N_25877,N_25297,N_24309);
or U25878 (N_25878,N_25006,N_24935);
xnor U25879 (N_25879,N_24039,N_24208);
nand U25880 (N_25880,N_24350,N_24948);
nor U25881 (N_25881,N_25248,N_25338);
xnor U25882 (N_25882,N_24455,N_24418);
and U25883 (N_25883,N_24697,N_24842);
nor U25884 (N_25884,N_24652,N_24996);
and U25885 (N_25885,N_24232,N_24977);
and U25886 (N_25886,N_25379,N_25456);
nand U25887 (N_25887,N_24602,N_24573);
nand U25888 (N_25888,N_24462,N_25165);
and U25889 (N_25889,N_24913,N_24962);
nor U25890 (N_25890,N_25210,N_24216);
or U25891 (N_25891,N_24973,N_25251);
nor U25892 (N_25892,N_24889,N_25056);
or U25893 (N_25893,N_24654,N_25305);
or U25894 (N_25894,N_24910,N_24870);
nor U25895 (N_25895,N_24147,N_24501);
nor U25896 (N_25896,N_25390,N_24992);
nor U25897 (N_25897,N_24126,N_24862);
or U25898 (N_25898,N_25344,N_24673);
and U25899 (N_25899,N_24268,N_25426);
nand U25900 (N_25900,N_24001,N_25054);
and U25901 (N_25901,N_24046,N_25371);
and U25902 (N_25902,N_24971,N_24811);
nor U25903 (N_25903,N_24554,N_24047);
nand U25904 (N_25904,N_24848,N_25343);
xor U25905 (N_25905,N_25234,N_24507);
and U25906 (N_25906,N_24027,N_25273);
nor U25907 (N_25907,N_25044,N_24683);
nor U25908 (N_25908,N_25013,N_24286);
nand U25909 (N_25909,N_24091,N_25298);
nor U25910 (N_25910,N_25116,N_24560);
xnor U25911 (N_25911,N_25384,N_24362);
and U25912 (N_25912,N_24884,N_24388);
nand U25913 (N_25913,N_24243,N_24179);
and U25914 (N_25914,N_24669,N_24199);
xnor U25915 (N_25915,N_25388,N_25151);
nor U25916 (N_25916,N_24880,N_24698);
nand U25917 (N_25917,N_24546,N_25428);
nor U25918 (N_25918,N_25385,N_25355);
and U25919 (N_25919,N_24417,N_25341);
and U25920 (N_25920,N_24058,N_24988);
and U25921 (N_25921,N_24648,N_24025);
and U25922 (N_25922,N_24130,N_24193);
nand U25923 (N_25923,N_24420,N_24643);
and U25924 (N_25924,N_24436,N_25254);
xor U25925 (N_25925,N_24023,N_24237);
nor U25926 (N_25926,N_25457,N_24967);
nor U25927 (N_25927,N_25022,N_25202);
nor U25928 (N_25928,N_24238,N_24352);
and U25929 (N_25929,N_25146,N_24143);
nand U25930 (N_25930,N_24945,N_24926);
nor U25931 (N_25931,N_24591,N_24074);
xor U25932 (N_25932,N_24229,N_24747);
nand U25933 (N_25933,N_24627,N_24095);
nor U25934 (N_25934,N_24305,N_24292);
xnor U25935 (N_25935,N_24438,N_25192);
nor U25936 (N_25936,N_24599,N_24336);
or U25937 (N_25937,N_24301,N_25252);
nand U25938 (N_25938,N_24879,N_25493);
and U25939 (N_25939,N_24326,N_24403);
nor U25940 (N_25940,N_25490,N_25402);
nand U25941 (N_25941,N_24860,N_24813);
nand U25942 (N_25942,N_24360,N_24328);
xnor U25943 (N_25943,N_25154,N_24952);
and U25944 (N_25944,N_24808,N_24065);
nand U25945 (N_25945,N_24279,N_24907);
or U25946 (N_25946,N_25152,N_24201);
and U25947 (N_25947,N_25157,N_24561);
nor U25948 (N_25948,N_24727,N_25306);
or U25949 (N_25949,N_24824,N_24831);
and U25950 (N_25950,N_24703,N_25364);
or U25951 (N_25951,N_24203,N_24223);
nand U25952 (N_25952,N_25118,N_24590);
or U25953 (N_25953,N_24760,N_24044);
nor U25954 (N_25954,N_24577,N_24772);
nand U25955 (N_25955,N_25262,N_24762);
xor U25956 (N_25956,N_24348,N_24556);
nor U25957 (N_25957,N_24195,N_25466);
nand U25958 (N_25958,N_25442,N_24746);
nand U25959 (N_25959,N_25083,N_24878);
nor U25960 (N_25960,N_24838,N_24183);
or U25961 (N_25961,N_24262,N_24707);
or U25962 (N_25962,N_25290,N_24787);
or U25963 (N_25963,N_25040,N_24659);
nand U25964 (N_25964,N_24780,N_24318);
nor U25965 (N_25965,N_24096,N_25101);
nand U25966 (N_25966,N_25274,N_24481);
nand U25967 (N_25967,N_24076,N_24717);
nand U25968 (N_25968,N_24276,N_25330);
or U25969 (N_25969,N_24244,N_24684);
and U25970 (N_25970,N_24260,N_24444);
or U25971 (N_25971,N_24476,N_24361);
or U25972 (N_25972,N_24251,N_24315);
nand U25973 (N_25973,N_24774,N_24019);
and U25974 (N_25974,N_24385,N_24274);
nor U25975 (N_25975,N_24872,N_24901);
nor U25976 (N_25976,N_25282,N_24939);
nor U25977 (N_25977,N_25484,N_25406);
nor U25978 (N_25978,N_24518,N_24398);
xnor U25979 (N_25979,N_24650,N_25123);
nor U25980 (N_25980,N_24919,N_25070);
xor U25981 (N_25981,N_25288,N_24736);
nand U25982 (N_25982,N_25219,N_25180);
nand U25983 (N_25983,N_24693,N_24841);
xor U25984 (N_25984,N_25131,N_24964);
or U25985 (N_25985,N_24116,N_24855);
or U25986 (N_25986,N_25145,N_24588);
nand U25987 (N_25987,N_24429,N_24633);
nand U25988 (N_25988,N_24200,N_25207);
or U25989 (N_25989,N_25060,N_24574);
nand U25990 (N_25990,N_25329,N_24484);
xnor U25991 (N_25991,N_24447,N_25382);
or U25992 (N_25992,N_24978,N_25050);
or U25993 (N_25993,N_24954,N_24190);
nor U25994 (N_25994,N_24181,N_24963);
or U25995 (N_25995,N_24063,N_25375);
nor U25996 (N_25996,N_24741,N_24677);
xnor U25997 (N_25997,N_25312,N_25358);
xor U25998 (N_25998,N_24716,N_24114);
or U25999 (N_25999,N_25087,N_24132);
and U26000 (N_26000,N_24498,N_24401);
nand U26001 (N_26001,N_25429,N_24103);
and U26002 (N_26002,N_24644,N_25189);
nor U26003 (N_26003,N_24815,N_24914);
xor U26004 (N_26004,N_24425,N_25129);
xor U26005 (N_26005,N_25034,N_24534);
xor U26006 (N_26006,N_24639,N_25141);
or U26007 (N_26007,N_24373,N_25481);
nand U26008 (N_26008,N_24081,N_24254);
nand U26009 (N_26009,N_25269,N_24144);
nand U26010 (N_26010,N_24711,N_24742);
xor U26011 (N_26011,N_24430,N_24210);
xnor U26012 (N_26012,N_24550,N_24474);
or U26013 (N_26013,N_25124,N_25195);
and U26014 (N_26014,N_24084,N_25125);
and U26015 (N_26015,N_24077,N_24920);
nor U26016 (N_26016,N_24032,N_25112);
or U26017 (N_26017,N_25027,N_24670);
xor U26018 (N_26018,N_25099,N_24482);
xnor U26019 (N_26019,N_24259,N_24125);
xor U26020 (N_26020,N_24998,N_24625);
or U26021 (N_26021,N_25272,N_24419);
or U26022 (N_26022,N_24341,N_24083);
nor U26023 (N_26023,N_25357,N_24592);
nor U26024 (N_26024,N_24390,N_24672);
or U26025 (N_26025,N_24970,N_25400);
nand U26026 (N_26026,N_25041,N_25378);
xnor U26027 (N_26027,N_24721,N_24628);
nand U26028 (N_26028,N_24753,N_24937);
nand U26029 (N_26029,N_25324,N_25430);
or U26030 (N_26030,N_24165,N_25143);
or U26031 (N_26031,N_25011,N_24994);
nand U26032 (N_26032,N_25156,N_25259);
and U26033 (N_26033,N_25058,N_24553);
and U26034 (N_26034,N_24911,N_25366);
xnor U26035 (N_26035,N_24873,N_24064);
nor U26036 (N_26036,N_24843,N_25133);
nand U26037 (N_26037,N_25052,N_25365);
or U26038 (N_26038,N_25049,N_25021);
nor U26039 (N_26039,N_24892,N_24740);
nand U26040 (N_26040,N_25369,N_25242);
and U26041 (N_26041,N_24769,N_24185);
or U26042 (N_26042,N_24640,N_25263);
and U26043 (N_26043,N_24930,N_24679);
nor U26044 (N_26044,N_24355,N_24586);
nand U26045 (N_26045,N_24680,N_25424);
nand U26046 (N_26046,N_24792,N_25023);
nand U26047 (N_26047,N_25103,N_24122);
and U26048 (N_26048,N_24133,N_25256);
or U26049 (N_26049,N_24513,N_24363);
nor U26050 (N_26050,N_25216,N_24411);
and U26051 (N_26051,N_24113,N_24532);
nor U26052 (N_26052,N_24102,N_25381);
xor U26053 (N_26053,N_25468,N_24757);
or U26054 (N_26054,N_25072,N_25240);
nor U26055 (N_26055,N_25440,N_24101);
xor U26056 (N_26056,N_25353,N_24258);
nor U26057 (N_26057,N_24284,N_25069);
xor U26058 (N_26058,N_24343,N_24576);
nor U26059 (N_26059,N_25467,N_25478);
xnor U26060 (N_26060,N_25095,N_24618);
nor U26061 (N_26061,N_25010,N_24211);
or U26062 (N_26062,N_24922,N_24823);
and U26063 (N_26063,N_24795,N_24331);
nor U26064 (N_26064,N_25175,N_24100);
nor U26065 (N_26065,N_24960,N_25107);
nand U26066 (N_26066,N_24788,N_25404);
or U26067 (N_26067,N_25483,N_24809);
nor U26068 (N_26068,N_25368,N_24192);
or U26069 (N_26069,N_24230,N_24423);
nor U26070 (N_26070,N_24160,N_24494);
or U26071 (N_26071,N_25130,N_24256);
and U26072 (N_26072,N_25372,N_24128);
nand U26073 (N_26073,N_25232,N_24451);
xor U26074 (N_26074,N_25321,N_25183);
or U26075 (N_26075,N_24589,N_25416);
nand U26076 (N_26076,N_24551,N_24802);
xor U26077 (N_26077,N_24601,N_25025);
xnor U26078 (N_26078,N_24887,N_24018);
xor U26079 (N_26079,N_24924,N_25465);
nor U26080 (N_26080,N_24928,N_24756);
and U26081 (N_26081,N_24478,N_24900);
xnor U26082 (N_26082,N_24739,N_24206);
nor U26083 (N_26083,N_25309,N_25304);
nand U26084 (N_26084,N_25243,N_25420);
or U26085 (N_26085,N_25485,N_24495);
or U26086 (N_26086,N_25132,N_24233);
nand U26087 (N_26087,N_25203,N_24798);
nand U26088 (N_26088,N_25413,N_25075);
nand U26089 (N_26089,N_24503,N_25326);
and U26090 (N_26090,N_24135,N_24511);
xnor U26091 (N_26091,N_25117,N_24867);
nand U26092 (N_26092,N_25427,N_24379);
nor U26093 (N_26093,N_24719,N_24980);
nand U26094 (N_26094,N_25163,N_24804);
or U26095 (N_26095,N_24487,N_25257);
or U26096 (N_26096,N_25308,N_25084);
and U26097 (N_26097,N_24985,N_24399);
or U26098 (N_26098,N_25078,N_24056);
and U26099 (N_26099,N_25496,N_24966);
xor U26100 (N_26100,N_25299,N_25283);
nand U26101 (N_26101,N_24280,N_25233);
nand U26102 (N_26102,N_24637,N_24631);
nand U26103 (N_26103,N_25038,N_25106);
xor U26104 (N_26104,N_24142,N_24332);
xor U26105 (N_26105,N_24107,N_25391);
and U26106 (N_26106,N_24535,N_24585);
nor U26107 (N_26107,N_24649,N_24374);
nand U26108 (N_26108,N_24859,N_25432);
or U26109 (N_26109,N_24761,N_24597);
nor U26110 (N_26110,N_24656,N_25008);
and U26111 (N_26111,N_25464,N_24623);
and U26112 (N_26112,N_24377,N_24751);
nand U26113 (N_26113,N_25294,N_25328);
nor U26114 (N_26114,N_24563,N_24771);
or U26115 (N_26115,N_24606,N_24180);
nand U26116 (N_26116,N_24953,N_25271);
and U26117 (N_26117,N_25236,N_24295);
xnor U26118 (N_26118,N_24509,N_24844);
xnor U26119 (N_26119,N_24317,N_24786);
and U26120 (N_26120,N_24045,N_25048);
nand U26121 (N_26121,N_24826,N_24439);
nor U26122 (N_26122,N_24579,N_24531);
xnor U26123 (N_26123,N_24225,N_24380);
nor U26124 (N_26124,N_24712,N_24908);
and U26125 (N_26125,N_24622,N_24079);
or U26126 (N_26126,N_25477,N_24020);
and U26127 (N_26127,N_24675,N_24093);
nand U26128 (N_26128,N_25223,N_25024);
nand U26129 (N_26129,N_24378,N_24104);
or U26130 (N_26130,N_24881,N_25409);
nand U26131 (N_26131,N_25452,N_24866);
nand U26132 (N_26132,N_25346,N_24325);
xor U26133 (N_26133,N_25327,N_24323);
or U26134 (N_26134,N_24578,N_24506);
xor U26135 (N_26135,N_24773,N_25374);
nor U26136 (N_26136,N_25245,N_24917);
or U26137 (N_26137,N_25286,N_25035);
nor U26138 (N_26138,N_25186,N_24790);
nand U26139 (N_26139,N_25043,N_24281);
xor U26140 (N_26140,N_24818,N_24957);
and U26141 (N_26141,N_24748,N_24311);
nand U26142 (N_26142,N_24817,N_24690);
and U26143 (N_26143,N_24171,N_25089);
nor U26144 (N_26144,N_24752,N_24883);
nor U26145 (N_26145,N_25159,N_25260);
or U26146 (N_26146,N_25431,N_24010);
and U26147 (N_26147,N_24381,N_24485);
xnor U26148 (N_26148,N_25356,N_25142);
or U26149 (N_26149,N_24021,N_25446);
nand U26150 (N_26150,N_24105,N_24816);
and U26151 (N_26151,N_24300,N_24030);
and U26152 (N_26152,N_24060,N_25316);
nor U26153 (N_26153,N_24457,N_24923);
nor U26154 (N_26154,N_24850,N_24497);
and U26155 (N_26155,N_24209,N_25300);
nand U26156 (N_26156,N_24156,N_25325);
xnor U26157 (N_26157,N_24464,N_24412);
nor U26158 (N_26158,N_25109,N_24611);
xor U26159 (N_26159,N_25170,N_24713);
nor U26160 (N_26160,N_24446,N_25012);
nand U26161 (N_26161,N_24454,N_24869);
and U26162 (N_26162,N_25289,N_24246);
xnor U26163 (N_26163,N_24642,N_24491);
nand U26164 (N_26164,N_24781,N_24828);
or U26165 (N_26165,N_25332,N_25182);
and U26166 (N_26166,N_24934,N_25435);
or U26167 (N_26167,N_25122,N_24427);
nand U26168 (N_26168,N_24483,N_25479);
nand U26169 (N_26169,N_24810,N_24342);
and U26170 (N_26170,N_24814,N_24909);
or U26171 (N_26171,N_24052,N_25176);
nor U26172 (N_26172,N_24938,N_25030);
or U26173 (N_26173,N_24358,N_24157);
or U26174 (N_26174,N_25313,N_24319);
nor U26175 (N_26175,N_25255,N_25450);
xor U26176 (N_26176,N_25033,N_24386);
xor U26177 (N_26177,N_24155,N_25302);
nor U26178 (N_26178,N_24136,N_24861);
or U26179 (N_26179,N_25395,N_24410);
nand U26180 (N_26180,N_24054,N_24593);
nand U26181 (N_26181,N_24807,N_24338);
xor U26182 (N_26182,N_25178,N_25094);
and U26183 (N_26183,N_24732,N_24220);
or U26184 (N_26184,N_24664,N_24092);
nand U26185 (N_26185,N_24529,N_24028);
nor U26186 (N_26186,N_25062,N_25144);
xor U26187 (N_26187,N_24086,N_24783);
and U26188 (N_26188,N_24856,N_25200);
nor U26189 (N_26189,N_24688,N_25423);
nand U26190 (N_26190,N_25414,N_24545);
or U26191 (N_26191,N_24138,N_24287);
nor U26192 (N_26192,N_25059,N_24453);
xnor U26193 (N_26193,N_24744,N_24106);
nor U26194 (N_26194,N_24477,N_24785);
xor U26195 (N_26195,N_25231,N_24617);
or U26196 (N_26196,N_24376,N_24131);
nand U26197 (N_26197,N_25350,N_25439);
or U26198 (N_26198,N_25340,N_25281);
or U26199 (N_26199,N_24609,N_24217);
nor U26200 (N_26200,N_25293,N_24121);
and U26201 (N_26201,N_24724,N_24634);
or U26202 (N_26202,N_24947,N_24067);
or U26203 (N_26203,N_25363,N_24704);
or U26204 (N_26204,N_24981,N_24678);
xor U26205 (N_26205,N_24888,N_24393);
or U26206 (N_26206,N_24662,N_24472);
xnor U26207 (N_26207,N_24851,N_24738);
and U26208 (N_26208,N_25472,N_25392);
nor U26209 (N_26209,N_25411,N_24098);
and U26210 (N_26210,N_24765,N_24109);
nor U26211 (N_26211,N_25140,N_24275);
nand U26212 (N_26212,N_25296,N_24463);
nand U26213 (N_26213,N_25362,N_25155);
xnor U26214 (N_26214,N_24893,N_24134);
nand U26215 (N_26215,N_25319,N_24070);
xnor U26216 (N_26216,N_24392,N_25174);
nand U26217 (N_26217,N_24424,N_24539);
or U26218 (N_26218,N_25387,N_24993);
xor U26219 (N_26219,N_25314,N_25185);
nand U26220 (N_26220,N_24094,N_24353);
xnor U26221 (N_26221,N_25128,N_25213);
and U26222 (N_26222,N_24955,N_25488);
nand U26223 (N_26223,N_25190,N_25401);
and U26224 (N_26224,N_24466,N_25235);
nand U26225 (N_26225,N_25497,N_25032);
and U26226 (N_26226,N_24767,N_25209);
xnor U26227 (N_26227,N_25071,N_24026);
and U26228 (N_26228,N_24667,N_25135);
nor U26229 (N_26229,N_24426,N_24184);
nand U26230 (N_26230,N_24024,N_24525);
xor U26231 (N_26231,N_24422,N_24099);
nor U26232 (N_26232,N_25222,N_24709);
xnor U26233 (N_26233,N_25090,N_24580);
and U26234 (N_26234,N_25215,N_24706);
nor U26235 (N_26235,N_24151,N_24146);
and U26236 (N_26236,N_24471,N_24150);
xor U26237 (N_26237,N_24365,N_24691);
and U26238 (N_26238,N_24035,N_24777);
xor U26239 (N_26239,N_25454,N_24306);
xnor U26240 (N_26240,N_25410,N_24214);
nor U26241 (N_26241,N_24835,N_24337);
xor U26242 (N_26242,N_24339,N_24542);
nor U26243 (N_26243,N_24140,N_24775);
or U26244 (N_26244,N_24829,N_24853);
xor U26245 (N_26245,N_24469,N_24557);
xor U26246 (N_26246,N_24687,N_25396);
nor U26247 (N_26247,N_24174,N_24565);
xor U26248 (N_26248,N_25345,N_24722);
or U26249 (N_26249,N_24582,N_24264);
or U26250 (N_26250,N_25326,N_24590);
nor U26251 (N_26251,N_24663,N_24393);
and U26252 (N_26252,N_24085,N_25283);
nor U26253 (N_26253,N_24798,N_25230);
and U26254 (N_26254,N_24251,N_25486);
or U26255 (N_26255,N_25160,N_24894);
xnor U26256 (N_26256,N_25250,N_24907);
or U26257 (N_26257,N_24988,N_24800);
nor U26258 (N_26258,N_25027,N_25141);
or U26259 (N_26259,N_24822,N_24090);
nor U26260 (N_26260,N_24318,N_24303);
or U26261 (N_26261,N_24536,N_25134);
xor U26262 (N_26262,N_24497,N_25382);
nor U26263 (N_26263,N_24344,N_24690);
or U26264 (N_26264,N_25464,N_25295);
nand U26265 (N_26265,N_25334,N_24073);
and U26266 (N_26266,N_24873,N_24702);
nand U26267 (N_26267,N_25298,N_24788);
and U26268 (N_26268,N_24999,N_24530);
nor U26269 (N_26269,N_24161,N_24365);
nand U26270 (N_26270,N_24923,N_24940);
and U26271 (N_26271,N_25291,N_24475);
nand U26272 (N_26272,N_24757,N_24926);
and U26273 (N_26273,N_24763,N_24152);
nor U26274 (N_26274,N_25029,N_24982);
and U26275 (N_26275,N_25497,N_24910);
nor U26276 (N_26276,N_24251,N_24811);
or U26277 (N_26277,N_24508,N_24482);
xor U26278 (N_26278,N_24911,N_24042);
xnor U26279 (N_26279,N_24132,N_25364);
and U26280 (N_26280,N_25103,N_25419);
xnor U26281 (N_26281,N_24570,N_24487);
or U26282 (N_26282,N_24610,N_24027);
or U26283 (N_26283,N_24148,N_24926);
xor U26284 (N_26284,N_24820,N_24180);
and U26285 (N_26285,N_24090,N_24597);
or U26286 (N_26286,N_24766,N_24944);
xnor U26287 (N_26287,N_24524,N_24241);
nand U26288 (N_26288,N_24741,N_24686);
nand U26289 (N_26289,N_25123,N_24283);
or U26290 (N_26290,N_25211,N_24103);
nor U26291 (N_26291,N_25058,N_24065);
nand U26292 (N_26292,N_24448,N_24479);
or U26293 (N_26293,N_25476,N_24037);
or U26294 (N_26294,N_24385,N_24793);
or U26295 (N_26295,N_24831,N_25315);
nand U26296 (N_26296,N_24834,N_24543);
nand U26297 (N_26297,N_25175,N_24013);
and U26298 (N_26298,N_24614,N_24211);
nand U26299 (N_26299,N_24706,N_24684);
xor U26300 (N_26300,N_24788,N_25393);
or U26301 (N_26301,N_25145,N_24273);
and U26302 (N_26302,N_25491,N_24238);
xnor U26303 (N_26303,N_24456,N_24592);
nor U26304 (N_26304,N_25064,N_25162);
or U26305 (N_26305,N_24873,N_24651);
nor U26306 (N_26306,N_24282,N_24701);
and U26307 (N_26307,N_25362,N_24255);
xnor U26308 (N_26308,N_25434,N_24227);
nor U26309 (N_26309,N_25148,N_25064);
nand U26310 (N_26310,N_25457,N_24263);
and U26311 (N_26311,N_24263,N_24450);
xnor U26312 (N_26312,N_24546,N_24742);
xor U26313 (N_26313,N_24614,N_24793);
xor U26314 (N_26314,N_24365,N_24286);
and U26315 (N_26315,N_25114,N_24097);
or U26316 (N_26316,N_24948,N_24973);
or U26317 (N_26317,N_24009,N_25492);
or U26318 (N_26318,N_24111,N_25470);
or U26319 (N_26319,N_24089,N_25354);
and U26320 (N_26320,N_24011,N_25265);
or U26321 (N_26321,N_24683,N_25405);
and U26322 (N_26322,N_24103,N_25152);
xor U26323 (N_26323,N_24798,N_25150);
nand U26324 (N_26324,N_24476,N_25216);
or U26325 (N_26325,N_24587,N_25019);
or U26326 (N_26326,N_24370,N_24133);
and U26327 (N_26327,N_24127,N_24656);
or U26328 (N_26328,N_25283,N_24281);
nand U26329 (N_26329,N_24615,N_24971);
and U26330 (N_26330,N_24266,N_25202);
and U26331 (N_26331,N_24296,N_24825);
or U26332 (N_26332,N_25295,N_25402);
or U26333 (N_26333,N_24191,N_24646);
nand U26334 (N_26334,N_24924,N_24061);
xnor U26335 (N_26335,N_25311,N_24882);
nand U26336 (N_26336,N_25463,N_25029);
xnor U26337 (N_26337,N_24347,N_25042);
nor U26338 (N_26338,N_24407,N_25332);
xnor U26339 (N_26339,N_24538,N_25250);
and U26340 (N_26340,N_24696,N_25066);
nand U26341 (N_26341,N_24029,N_25187);
or U26342 (N_26342,N_24873,N_24836);
nor U26343 (N_26343,N_25311,N_24512);
nand U26344 (N_26344,N_24427,N_24410);
xor U26345 (N_26345,N_24641,N_24504);
xnor U26346 (N_26346,N_25176,N_24940);
nand U26347 (N_26347,N_24071,N_24477);
nand U26348 (N_26348,N_24718,N_24927);
and U26349 (N_26349,N_24848,N_24738);
and U26350 (N_26350,N_25315,N_25393);
xor U26351 (N_26351,N_24080,N_24225);
nor U26352 (N_26352,N_24527,N_25412);
nor U26353 (N_26353,N_24992,N_25152);
xnor U26354 (N_26354,N_24494,N_24916);
and U26355 (N_26355,N_25478,N_25256);
nand U26356 (N_26356,N_25104,N_24024);
or U26357 (N_26357,N_24814,N_24673);
or U26358 (N_26358,N_24847,N_24645);
nor U26359 (N_26359,N_25464,N_24633);
or U26360 (N_26360,N_25326,N_25413);
nand U26361 (N_26361,N_24739,N_24536);
or U26362 (N_26362,N_25404,N_25397);
nor U26363 (N_26363,N_24671,N_24760);
nor U26364 (N_26364,N_24613,N_24078);
nor U26365 (N_26365,N_24508,N_24165);
or U26366 (N_26366,N_25320,N_25391);
or U26367 (N_26367,N_24128,N_25103);
nor U26368 (N_26368,N_24894,N_24423);
or U26369 (N_26369,N_24697,N_24198);
xnor U26370 (N_26370,N_25275,N_25030);
and U26371 (N_26371,N_25006,N_24575);
and U26372 (N_26372,N_24436,N_25062);
and U26373 (N_26373,N_24632,N_24778);
and U26374 (N_26374,N_24054,N_25096);
or U26375 (N_26375,N_24901,N_25210);
nor U26376 (N_26376,N_25363,N_24538);
nand U26377 (N_26377,N_25383,N_24445);
xor U26378 (N_26378,N_25295,N_24792);
xnor U26379 (N_26379,N_24194,N_24978);
xor U26380 (N_26380,N_24597,N_25174);
or U26381 (N_26381,N_24819,N_24679);
nand U26382 (N_26382,N_24257,N_24853);
and U26383 (N_26383,N_24465,N_24582);
nor U26384 (N_26384,N_25216,N_24180);
nor U26385 (N_26385,N_24735,N_24879);
or U26386 (N_26386,N_24495,N_25104);
xnor U26387 (N_26387,N_24645,N_24475);
and U26388 (N_26388,N_24333,N_24619);
nand U26389 (N_26389,N_25309,N_25091);
nor U26390 (N_26390,N_24135,N_24875);
or U26391 (N_26391,N_24326,N_24079);
xor U26392 (N_26392,N_24370,N_24595);
nand U26393 (N_26393,N_25025,N_25138);
nand U26394 (N_26394,N_24222,N_24829);
xor U26395 (N_26395,N_24582,N_24934);
xnor U26396 (N_26396,N_25020,N_24066);
nand U26397 (N_26397,N_24817,N_25106);
and U26398 (N_26398,N_24010,N_24482);
xnor U26399 (N_26399,N_24162,N_24074);
nor U26400 (N_26400,N_24785,N_25435);
and U26401 (N_26401,N_24885,N_24553);
xor U26402 (N_26402,N_24896,N_24824);
nor U26403 (N_26403,N_24358,N_24276);
and U26404 (N_26404,N_24401,N_24151);
nand U26405 (N_26405,N_24440,N_25342);
and U26406 (N_26406,N_25387,N_24212);
xnor U26407 (N_26407,N_24688,N_25053);
nor U26408 (N_26408,N_24224,N_24449);
and U26409 (N_26409,N_25320,N_25270);
nor U26410 (N_26410,N_24533,N_24756);
or U26411 (N_26411,N_24114,N_24891);
or U26412 (N_26412,N_24887,N_25385);
and U26413 (N_26413,N_24655,N_24963);
or U26414 (N_26414,N_24465,N_24466);
nand U26415 (N_26415,N_25298,N_25440);
or U26416 (N_26416,N_24894,N_24882);
xnor U26417 (N_26417,N_25407,N_25375);
xnor U26418 (N_26418,N_24824,N_24750);
nand U26419 (N_26419,N_25305,N_24779);
and U26420 (N_26420,N_25374,N_25159);
nand U26421 (N_26421,N_24290,N_24023);
xor U26422 (N_26422,N_24000,N_24075);
or U26423 (N_26423,N_24590,N_25147);
nand U26424 (N_26424,N_24943,N_25498);
xnor U26425 (N_26425,N_25469,N_24932);
nor U26426 (N_26426,N_25269,N_24670);
nand U26427 (N_26427,N_25191,N_24066);
and U26428 (N_26428,N_25362,N_24387);
nor U26429 (N_26429,N_25198,N_24201);
and U26430 (N_26430,N_24473,N_24462);
or U26431 (N_26431,N_25308,N_25326);
and U26432 (N_26432,N_25394,N_24080);
nor U26433 (N_26433,N_25391,N_24529);
nor U26434 (N_26434,N_25188,N_25126);
nand U26435 (N_26435,N_25043,N_24779);
nand U26436 (N_26436,N_24108,N_24317);
nor U26437 (N_26437,N_25049,N_25191);
nor U26438 (N_26438,N_24542,N_24496);
nor U26439 (N_26439,N_24728,N_25194);
or U26440 (N_26440,N_24696,N_24424);
xor U26441 (N_26441,N_24590,N_24663);
nand U26442 (N_26442,N_24663,N_24749);
xor U26443 (N_26443,N_24347,N_24664);
or U26444 (N_26444,N_24791,N_24904);
xnor U26445 (N_26445,N_24411,N_25065);
or U26446 (N_26446,N_24370,N_24221);
and U26447 (N_26447,N_24306,N_25468);
or U26448 (N_26448,N_24878,N_24431);
nand U26449 (N_26449,N_24474,N_25059);
nor U26450 (N_26450,N_24916,N_24277);
nand U26451 (N_26451,N_25035,N_24855);
or U26452 (N_26452,N_24251,N_24808);
or U26453 (N_26453,N_24322,N_25370);
or U26454 (N_26454,N_25378,N_24072);
and U26455 (N_26455,N_24647,N_24072);
and U26456 (N_26456,N_25226,N_24195);
and U26457 (N_26457,N_24848,N_24954);
xnor U26458 (N_26458,N_24379,N_24116);
or U26459 (N_26459,N_24881,N_24493);
and U26460 (N_26460,N_24415,N_25065);
or U26461 (N_26461,N_25113,N_25239);
nor U26462 (N_26462,N_25117,N_24353);
and U26463 (N_26463,N_24950,N_24868);
nor U26464 (N_26464,N_24090,N_24697);
nand U26465 (N_26465,N_24241,N_24087);
and U26466 (N_26466,N_25178,N_25186);
xor U26467 (N_26467,N_24224,N_25118);
nand U26468 (N_26468,N_24682,N_25444);
xor U26469 (N_26469,N_24276,N_24923);
and U26470 (N_26470,N_25349,N_24244);
nand U26471 (N_26471,N_25282,N_25117);
nand U26472 (N_26472,N_25122,N_24689);
xor U26473 (N_26473,N_25360,N_24366);
xor U26474 (N_26474,N_24686,N_25157);
xnor U26475 (N_26475,N_25477,N_24396);
or U26476 (N_26476,N_24545,N_24652);
nor U26477 (N_26477,N_24802,N_24247);
xor U26478 (N_26478,N_24663,N_24071);
or U26479 (N_26479,N_24204,N_24222);
and U26480 (N_26480,N_25308,N_25019);
and U26481 (N_26481,N_24953,N_25234);
xor U26482 (N_26482,N_24045,N_25416);
xor U26483 (N_26483,N_25095,N_24303);
nor U26484 (N_26484,N_24010,N_24931);
nand U26485 (N_26485,N_24942,N_24511);
xnor U26486 (N_26486,N_25270,N_25383);
xor U26487 (N_26487,N_24464,N_24823);
xnor U26488 (N_26488,N_24450,N_24145);
and U26489 (N_26489,N_24713,N_25338);
nand U26490 (N_26490,N_24571,N_25348);
or U26491 (N_26491,N_24819,N_24083);
and U26492 (N_26492,N_24990,N_25294);
nor U26493 (N_26493,N_24817,N_24715);
or U26494 (N_26494,N_24347,N_24213);
or U26495 (N_26495,N_24878,N_24561);
or U26496 (N_26496,N_24571,N_24735);
and U26497 (N_26497,N_24585,N_25332);
nor U26498 (N_26498,N_24069,N_24408);
or U26499 (N_26499,N_24034,N_25032);
nand U26500 (N_26500,N_24075,N_24948);
xor U26501 (N_26501,N_25185,N_24053);
nand U26502 (N_26502,N_24026,N_24162);
xor U26503 (N_26503,N_24540,N_24775);
or U26504 (N_26504,N_25183,N_24497);
nor U26505 (N_26505,N_24453,N_24909);
nor U26506 (N_26506,N_24085,N_24840);
or U26507 (N_26507,N_25145,N_24047);
and U26508 (N_26508,N_24833,N_25224);
nand U26509 (N_26509,N_24147,N_24703);
or U26510 (N_26510,N_24431,N_25013);
nand U26511 (N_26511,N_25179,N_24182);
or U26512 (N_26512,N_25055,N_24221);
xnor U26513 (N_26513,N_24983,N_24315);
nor U26514 (N_26514,N_24737,N_24083);
nand U26515 (N_26515,N_25026,N_24826);
or U26516 (N_26516,N_24460,N_25217);
xor U26517 (N_26517,N_24308,N_25198);
or U26518 (N_26518,N_25366,N_24813);
or U26519 (N_26519,N_24111,N_24779);
or U26520 (N_26520,N_24516,N_25277);
xnor U26521 (N_26521,N_25077,N_24109);
nand U26522 (N_26522,N_24569,N_25083);
xnor U26523 (N_26523,N_24529,N_24361);
and U26524 (N_26524,N_25320,N_24679);
xnor U26525 (N_26525,N_24797,N_25484);
xor U26526 (N_26526,N_24760,N_25185);
nand U26527 (N_26527,N_24404,N_25403);
or U26528 (N_26528,N_24928,N_25208);
or U26529 (N_26529,N_24201,N_25292);
and U26530 (N_26530,N_24924,N_24281);
xor U26531 (N_26531,N_24798,N_24459);
xor U26532 (N_26532,N_25448,N_24042);
nor U26533 (N_26533,N_24803,N_24609);
xor U26534 (N_26534,N_24756,N_25352);
xnor U26535 (N_26535,N_24150,N_25262);
nand U26536 (N_26536,N_24766,N_24319);
or U26537 (N_26537,N_24219,N_24472);
nor U26538 (N_26538,N_24410,N_24315);
xnor U26539 (N_26539,N_24297,N_24221);
xor U26540 (N_26540,N_24404,N_24989);
nor U26541 (N_26541,N_24774,N_24910);
xnor U26542 (N_26542,N_24150,N_24050);
and U26543 (N_26543,N_24916,N_24996);
xnor U26544 (N_26544,N_24754,N_24759);
nand U26545 (N_26545,N_25002,N_24515);
and U26546 (N_26546,N_25027,N_24759);
or U26547 (N_26547,N_25495,N_24955);
xor U26548 (N_26548,N_24085,N_24323);
nor U26549 (N_26549,N_24344,N_24623);
nor U26550 (N_26550,N_25378,N_24375);
xnor U26551 (N_26551,N_24457,N_24071);
and U26552 (N_26552,N_24293,N_24187);
or U26553 (N_26553,N_24517,N_24968);
and U26554 (N_26554,N_24174,N_24015);
and U26555 (N_26555,N_24802,N_24645);
xnor U26556 (N_26556,N_25329,N_24732);
nand U26557 (N_26557,N_24315,N_24019);
and U26558 (N_26558,N_25071,N_24158);
xnor U26559 (N_26559,N_24893,N_24958);
and U26560 (N_26560,N_24985,N_24965);
and U26561 (N_26561,N_25087,N_25057);
nand U26562 (N_26562,N_24870,N_25398);
nor U26563 (N_26563,N_25316,N_24893);
xnor U26564 (N_26564,N_24672,N_25467);
or U26565 (N_26565,N_24563,N_24257);
and U26566 (N_26566,N_25068,N_24071);
nand U26567 (N_26567,N_24781,N_24309);
nand U26568 (N_26568,N_25146,N_24282);
or U26569 (N_26569,N_25406,N_24714);
or U26570 (N_26570,N_25262,N_24151);
nand U26571 (N_26571,N_24583,N_25192);
nor U26572 (N_26572,N_24980,N_24078);
or U26573 (N_26573,N_24776,N_24156);
and U26574 (N_26574,N_24746,N_24156);
and U26575 (N_26575,N_25241,N_24215);
nor U26576 (N_26576,N_25081,N_25157);
nand U26577 (N_26577,N_24800,N_25174);
nand U26578 (N_26578,N_24605,N_24202);
nand U26579 (N_26579,N_24480,N_24503);
or U26580 (N_26580,N_24052,N_25367);
or U26581 (N_26581,N_25465,N_24309);
nor U26582 (N_26582,N_24167,N_24901);
xnor U26583 (N_26583,N_24857,N_25311);
nor U26584 (N_26584,N_24463,N_25238);
and U26585 (N_26585,N_24406,N_24652);
nor U26586 (N_26586,N_25295,N_24625);
or U26587 (N_26587,N_24843,N_24363);
nor U26588 (N_26588,N_24873,N_24759);
xor U26589 (N_26589,N_24693,N_24078);
or U26590 (N_26590,N_24794,N_25399);
or U26591 (N_26591,N_24273,N_25424);
nor U26592 (N_26592,N_24564,N_25209);
or U26593 (N_26593,N_25239,N_24240);
nand U26594 (N_26594,N_25188,N_24331);
nor U26595 (N_26595,N_24978,N_24896);
nor U26596 (N_26596,N_25326,N_25227);
nor U26597 (N_26597,N_24101,N_24477);
and U26598 (N_26598,N_24504,N_24940);
and U26599 (N_26599,N_24683,N_24616);
nand U26600 (N_26600,N_24841,N_24676);
nor U26601 (N_26601,N_24502,N_24468);
nor U26602 (N_26602,N_24524,N_24024);
nand U26603 (N_26603,N_24540,N_24369);
xnor U26604 (N_26604,N_24043,N_24545);
and U26605 (N_26605,N_24061,N_24383);
xor U26606 (N_26606,N_24143,N_24372);
nand U26607 (N_26607,N_25078,N_24442);
or U26608 (N_26608,N_24850,N_25119);
nor U26609 (N_26609,N_24209,N_24963);
nor U26610 (N_26610,N_24873,N_24634);
or U26611 (N_26611,N_25281,N_25153);
xor U26612 (N_26612,N_24756,N_25358);
and U26613 (N_26613,N_24215,N_25231);
xnor U26614 (N_26614,N_25227,N_25273);
or U26615 (N_26615,N_24083,N_24467);
or U26616 (N_26616,N_24497,N_25495);
and U26617 (N_26617,N_24047,N_24048);
nor U26618 (N_26618,N_24167,N_24003);
nor U26619 (N_26619,N_24394,N_24701);
and U26620 (N_26620,N_24911,N_24512);
and U26621 (N_26621,N_24253,N_25233);
nand U26622 (N_26622,N_24378,N_24338);
or U26623 (N_26623,N_25167,N_24133);
xnor U26624 (N_26624,N_24673,N_24067);
and U26625 (N_26625,N_25446,N_25287);
or U26626 (N_26626,N_25319,N_24378);
xor U26627 (N_26627,N_25220,N_25047);
nand U26628 (N_26628,N_25234,N_24436);
and U26629 (N_26629,N_25238,N_24467);
or U26630 (N_26630,N_25215,N_25453);
and U26631 (N_26631,N_25255,N_25430);
and U26632 (N_26632,N_25002,N_24604);
xnor U26633 (N_26633,N_24725,N_24106);
xnor U26634 (N_26634,N_24891,N_24758);
and U26635 (N_26635,N_24777,N_24962);
xor U26636 (N_26636,N_24636,N_24984);
or U26637 (N_26637,N_25173,N_25370);
nand U26638 (N_26638,N_24255,N_24911);
xnor U26639 (N_26639,N_24252,N_24306);
nor U26640 (N_26640,N_24568,N_24809);
and U26641 (N_26641,N_25461,N_24808);
nor U26642 (N_26642,N_24702,N_24280);
or U26643 (N_26643,N_24379,N_25155);
and U26644 (N_26644,N_24411,N_24110);
nand U26645 (N_26645,N_25280,N_24809);
or U26646 (N_26646,N_24359,N_24699);
or U26647 (N_26647,N_24174,N_24104);
nand U26648 (N_26648,N_24265,N_24217);
xor U26649 (N_26649,N_25119,N_25261);
and U26650 (N_26650,N_25102,N_25023);
xnor U26651 (N_26651,N_24150,N_24715);
nor U26652 (N_26652,N_24586,N_24881);
and U26653 (N_26653,N_24268,N_25179);
or U26654 (N_26654,N_24504,N_24648);
and U26655 (N_26655,N_25376,N_24710);
xor U26656 (N_26656,N_24228,N_24038);
nand U26657 (N_26657,N_24576,N_24191);
or U26658 (N_26658,N_25397,N_25243);
nand U26659 (N_26659,N_24664,N_25453);
nand U26660 (N_26660,N_24941,N_24207);
and U26661 (N_26661,N_25142,N_24887);
nand U26662 (N_26662,N_24239,N_24803);
nor U26663 (N_26663,N_24537,N_25392);
xor U26664 (N_26664,N_25438,N_24784);
or U26665 (N_26665,N_25426,N_24789);
or U26666 (N_26666,N_24242,N_24666);
or U26667 (N_26667,N_24192,N_24018);
nor U26668 (N_26668,N_25338,N_24419);
or U26669 (N_26669,N_25438,N_25081);
and U26670 (N_26670,N_24256,N_24015);
xnor U26671 (N_26671,N_24903,N_24847);
or U26672 (N_26672,N_24404,N_25035);
xnor U26673 (N_26673,N_24809,N_24662);
nor U26674 (N_26674,N_24169,N_25074);
nand U26675 (N_26675,N_24151,N_25123);
nor U26676 (N_26676,N_25173,N_25096);
xor U26677 (N_26677,N_24931,N_24828);
nand U26678 (N_26678,N_24628,N_25476);
nand U26679 (N_26679,N_24179,N_24358);
nor U26680 (N_26680,N_24606,N_24972);
or U26681 (N_26681,N_24490,N_25038);
nor U26682 (N_26682,N_24927,N_24234);
nand U26683 (N_26683,N_24370,N_24441);
and U26684 (N_26684,N_25100,N_24839);
nand U26685 (N_26685,N_24856,N_24885);
and U26686 (N_26686,N_25392,N_24010);
and U26687 (N_26687,N_24734,N_24650);
and U26688 (N_26688,N_25028,N_25131);
xnor U26689 (N_26689,N_24188,N_24364);
nand U26690 (N_26690,N_24235,N_25447);
and U26691 (N_26691,N_25247,N_25463);
nor U26692 (N_26692,N_25490,N_25226);
or U26693 (N_26693,N_24929,N_25416);
nor U26694 (N_26694,N_25403,N_25320);
nor U26695 (N_26695,N_24172,N_24756);
nand U26696 (N_26696,N_25054,N_24845);
xnor U26697 (N_26697,N_24625,N_24434);
or U26698 (N_26698,N_25358,N_24124);
nor U26699 (N_26699,N_24341,N_24594);
nand U26700 (N_26700,N_25007,N_25485);
nor U26701 (N_26701,N_24787,N_24015);
or U26702 (N_26702,N_24510,N_24630);
or U26703 (N_26703,N_25147,N_24995);
and U26704 (N_26704,N_24504,N_24148);
or U26705 (N_26705,N_25443,N_24285);
nor U26706 (N_26706,N_25128,N_24217);
or U26707 (N_26707,N_24027,N_25298);
xnor U26708 (N_26708,N_24095,N_24798);
xor U26709 (N_26709,N_24857,N_24462);
nor U26710 (N_26710,N_24047,N_25274);
xor U26711 (N_26711,N_25232,N_24262);
xor U26712 (N_26712,N_24200,N_25281);
xor U26713 (N_26713,N_24575,N_24648);
nor U26714 (N_26714,N_25341,N_24823);
nor U26715 (N_26715,N_24347,N_24110);
nor U26716 (N_26716,N_24910,N_24370);
xnor U26717 (N_26717,N_24345,N_25062);
nor U26718 (N_26718,N_24176,N_24642);
nand U26719 (N_26719,N_25187,N_25098);
and U26720 (N_26720,N_24002,N_24288);
nand U26721 (N_26721,N_25197,N_25040);
nand U26722 (N_26722,N_25116,N_24742);
and U26723 (N_26723,N_24775,N_24285);
and U26724 (N_26724,N_24361,N_24462);
or U26725 (N_26725,N_24258,N_25128);
nor U26726 (N_26726,N_24113,N_24905);
nor U26727 (N_26727,N_25481,N_25019);
nor U26728 (N_26728,N_24451,N_24212);
and U26729 (N_26729,N_25457,N_24874);
or U26730 (N_26730,N_24843,N_24459);
or U26731 (N_26731,N_24866,N_25408);
and U26732 (N_26732,N_25371,N_25029);
nand U26733 (N_26733,N_24538,N_24864);
nand U26734 (N_26734,N_25283,N_24042);
nand U26735 (N_26735,N_25313,N_24973);
or U26736 (N_26736,N_25481,N_24609);
nand U26737 (N_26737,N_25375,N_24503);
xnor U26738 (N_26738,N_25195,N_24599);
xnor U26739 (N_26739,N_24285,N_25332);
or U26740 (N_26740,N_24303,N_24892);
xnor U26741 (N_26741,N_24030,N_24650);
or U26742 (N_26742,N_24696,N_25395);
xnor U26743 (N_26743,N_24879,N_24564);
xor U26744 (N_26744,N_24675,N_25105);
or U26745 (N_26745,N_24541,N_25253);
and U26746 (N_26746,N_24725,N_24881);
nor U26747 (N_26747,N_24549,N_25491);
nor U26748 (N_26748,N_24909,N_24825);
nand U26749 (N_26749,N_24734,N_24489);
and U26750 (N_26750,N_24428,N_25280);
and U26751 (N_26751,N_24418,N_24990);
xor U26752 (N_26752,N_24053,N_25261);
nor U26753 (N_26753,N_24530,N_24763);
and U26754 (N_26754,N_24633,N_24657);
and U26755 (N_26755,N_24804,N_24653);
nor U26756 (N_26756,N_24936,N_24249);
and U26757 (N_26757,N_24557,N_24175);
nand U26758 (N_26758,N_24414,N_24606);
nand U26759 (N_26759,N_24564,N_24051);
or U26760 (N_26760,N_25297,N_25140);
and U26761 (N_26761,N_24521,N_24953);
nor U26762 (N_26762,N_24825,N_24042);
nand U26763 (N_26763,N_24369,N_24182);
xnor U26764 (N_26764,N_24343,N_24694);
or U26765 (N_26765,N_24177,N_25480);
or U26766 (N_26766,N_24655,N_25194);
and U26767 (N_26767,N_24245,N_25044);
xor U26768 (N_26768,N_25417,N_25189);
xor U26769 (N_26769,N_25037,N_25089);
xnor U26770 (N_26770,N_24100,N_24492);
and U26771 (N_26771,N_24081,N_25152);
nor U26772 (N_26772,N_24717,N_25353);
nand U26773 (N_26773,N_24306,N_24569);
xnor U26774 (N_26774,N_24996,N_25202);
or U26775 (N_26775,N_25499,N_24128);
nor U26776 (N_26776,N_24831,N_25214);
xor U26777 (N_26777,N_25367,N_24456);
nand U26778 (N_26778,N_25416,N_24795);
nor U26779 (N_26779,N_24479,N_25008);
and U26780 (N_26780,N_24853,N_24411);
or U26781 (N_26781,N_24822,N_24618);
nand U26782 (N_26782,N_24671,N_24628);
nor U26783 (N_26783,N_24046,N_25357);
nor U26784 (N_26784,N_25289,N_24873);
and U26785 (N_26785,N_24480,N_24502);
or U26786 (N_26786,N_24452,N_24472);
or U26787 (N_26787,N_24394,N_24186);
nand U26788 (N_26788,N_25048,N_24335);
nor U26789 (N_26789,N_25381,N_24541);
and U26790 (N_26790,N_24371,N_24204);
and U26791 (N_26791,N_24595,N_24867);
nor U26792 (N_26792,N_24311,N_25105);
nand U26793 (N_26793,N_24366,N_24991);
nand U26794 (N_26794,N_25072,N_25359);
nand U26795 (N_26795,N_24461,N_25006);
and U26796 (N_26796,N_24330,N_24228);
and U26797 (N_26797,N_24653,N_24692);
xor U26798 (N_26798,N_24128,N_24293);
and U26799 (N_26799,N_24569,N_25468);
nand U26800 (N_26800,N_25129,N_24417);
or U26801 (N_26801,N_25365,N_24716);
nor U26802 (N_26802,N_24577,N_24463);
xor U26803 (N_26803,N_24116,N_24250);
nand U26804 (N_26804,N_24137,N_24480);
nor U26805 (N_26805,N_24259,N_24128);
xor U26806 (N_26806,N_24882,N_24364);
xnor U26807 (N_26807,N_24232,N_25498);
and U26808 (N_26808,N_24946,N_25250);
nand U26809 (N_26809,N_25070,N_24147);
xor U26810 (N_26810,N_25467,N_24613);
or U26811 (N_26811,N_25451,N_24900);
and U26812 (N_26812,N_25148,N_24779);
nor U26813 (N_26813,N_25275,N_24947);
nand U26814 (N_26814,N_24544,N_24342);
or U26815 (N_26815,N_25314,N_24548);
and U26816 (N_26816,N_25416,N_24711);
and U26817 (N_26817,N_25274,N_24114);
nor U26818 (N_26818,N_24984,N_25228);
nor U26819 (N_26819,N_24521,N_24426);
and U26820 (N_26820,N_24732,N_24385);
and U26821 (N_26821,N_24711,N_24640);
xnor U26822 (N_26822,N_24732,N_24531);
nor U26823 (N_26823,N_24409,N_24289);
xor U26824 (N_26824,N_25355,N_24152);
nand U26825 (N_26825,N_24759,N_24618);
xnor U26826 (N_26826,N_24313,N_24291);
or U26827 (N_26827,N_24037,N_24744);
xnor U26828 (N_26828,N_25316,N_24222);
nor U26829 (N_26829,N_25148,N_25192);
xor U26830 (N_26830,N_25271,N_24603);
and U26831 (N_26831,N_24426,N_24357);
xnor U26832 (N_26832,N_24058,N_25021);
nor U26833 (N_26833,N_24753,N_24939);
and U26834 (N_26834,N_24197,N_24973);
xor U26835 (N_26835,N_25437,N_25174);
nand U26836 (N_26836,N_24760,N_25495);
nor U26837 (N_26837,N_25198,N_25176);
nand U26838 (N_26838,N_25177,N_24019);
nand U26839 (N_26839,N_25354,N_24775);
and U26840 (N_26840,N_24071,N_24116);
xnor U26841 (N_26841,N_24788,N_24584);
nor U26842 (N_26842,N_24014,N_24035);
nor U26843 (N_26843,N_25160,N_24056);
or U26844 (N_26844,N_24397,N_25471);
nor U26845 (N_26845,N_24958,N_24248);
nand U26846 (N_26846,N_25063,N_24411);
and U26847 (N_26847,N_24119,N_25268);
xor U26848 (N_26848,N_25114,N_24410);
and U26849 (N_26849,N_24003,N_24099);
nand U26850 (N_26850,N_24469,N_25035);
or U26851 (N_26851,N_25271,N_24629);
and U26852 (N_26852,N_24145,N_25375);
and U26853 (N_26853,N_25233,N_25150);
xor U26854 (N_26854,N_24841,N_24929);
nor U26855 (N_26855,N_25340,N_24116);
or U26856 (N_26856,N_25114,N_25414);
xnor U26857 (N_26857,N_24011,N_24438);
or U26858 (N_26858,N_24947,N_25475);
and U26859 (N_26859,N_24829,N_24444);
xor U26860 (N_26860,N_24190,N_25309);
and U26861 (N_26861,N_24386,N_24620);
or U26862 (N_26862,N_25470,N_24746);
and U26863 (N_26863,N_24286,N_24120);
and U26864 (N_26864,N_25407,N_24652);
xnor U26865 (N_26865,N_25088,N_24295);
nand U26866 (N_26866,N_24260,N_24135);
nor U26867 (N_26867,N_24321,N_24821);
nand U26868 (N_26868,N_25232,N_25012);
or U26869 (N_26869,N_24094,N_24115);
nand U26870 (N_26870,N_24538,N_24449);
and U26871 (N_26871,N_24817,N_25160);
and U26872 (N_26872,N_24490,N_24362);
xor U26873 (N_26873,N_25322,N_25283);
and U26874 (N_26874,N_25342,N_24857);
nand U26875 (N_26875,N_25200,N_25278);
and U26876 (N_26876,N_24380,N_24557);
xnor U26877 (N_26877,N_24911,N_24807);
and U26878 (N_26878,N_24152,N_24428);
nand U26879 (N_26879,N_25086,N_24505);
and U26880 (N_26880,N_24780,N_24055);
nor U26881 (N_26881,N_25468,N_24398);
xor U26882 (N_26882,N_25297,N_24045);
and U26883 (N_26883,N_24443,N_24564);
nor U26884 (N_26884,N_24656,N_24732);
or U26885 (N_26885,N_24268,N_25246);
xnor U26886 (N_26886,N_25160,N_25358);
nor U26887 (N_26887,N_24275,N_24003);
nor U26888 (N_26888,N_24635,N_24650);
xor U26889 (N_26889,N_24776,N_24417);
and U26890 (N_26890,N_25497,N_24653);
nand U26891 (N_26891,N_24286,N_24312);
xor U26892 (N_26892,N_24971,N_24840);
or U26893 (N_26893,N_25174,N_25306);
nand U26894 (N_26894,N_25415,N_24259);
and U26895 (N_26895,N_24168,N_24944);
nor U26896 (N_26896,N_25444,N_25350);
xnor U26897 (N_26897,N_24209,N_24398);
or U26898 (N_26898,N_25135,N_25242);
nand U26899 (N_26899,N_25141,N_24522);
nor U26900 (N_26900,N_24615,N_24451);
nor U26901 (N_26901,N_24716,N_24466);
nor U26902 (N_26902,N_25377,N_25101);
nand U26903 (N_26903,N_24647,N_24118);
nor U26904 (N_26904,N_24495,N_24388);
and U26905 (N_26905,N_24651,N_25103);
xnor U26906 (N_26906,N_24579,N_24607);
and U26907 (N_26907,N_25047,N_24675);
nor U26908 (N_26908,N_24363,N_24607);
nand U26909 (N_26909,N_25217,N_24982);
and U26910 (N_26910,N_25433,N_24248);
and U26911 (N_26911,N_24188,N_25192);
xor U26912 (N_26912,N_24936,N_25153);
xor U26913 (N_26913,N_25047,N_25137);
xor U26914 (N_26914,N_24668,N_24697);
xnor U26915 (N_26915,N_25004,N_25081);
or U26916 (N_26916,N_25241,N_25470);
xnor U26917 (N_26917,N_25430,N_25365);
xnor U26918 (N_26918,N_24708,N_24190);
and U26919 (N_26919,N_24740,N_25403);
nand U26920 (N_26920,N_25050,N_24824);
nand U26921 (N_26921,N_24119,N_24675);
and U26922 (N_26922,N_24532,N_24858);
xnor U26923 (N_26923,N_24164,N_24331);
nor U26924 (N_26924,N_24573,N_24144);
or U26925 (N_26925,N_24319,N_24156);
nand U26926 (N_26926,N_24009,N_25232);
xor U26927 (N_26927,N_25311,N_24050);
and U26928 (N_26928,N_24042,N_25354);
or U26929 (N_26929,N_25438,N_25317);
and U26930 (N_26930,N_24757,N_24759);
xnor U26931 (N_26931,N_24519,N_24835);
xnor U26932 (N_26932,N_25281,N_24664);
nand U26933 (N_26933,N_24620,N_25031);
nand U26934 (N_26934,N_25091,N_24894);
nor U26935 (N_26935,N_25328,N_24249);
and U26936 (N_26936,N_25114,N_24560);
or U26937 (N_26937,N_25155,N_24928);
nand U26938 (N_26938,N_24497,N_24655);
and U26939 (N_26939,N_24101,N_25088);
xor U26940 (N_26940,N_25208,N_25376);
and U26941 (N_26941,N_25186,N_25342);
or U26942 (N_26942,N_25291,N_25022);
nand U26943 (N_26943,N_24435,N_25132);
nand U26944 (N_26944,N_25255,N_24724);
xnor U26945 (N_26945,N_24150,N_25335);
and U26946 (N_26946,N_24822,N_24723);
and U26947 (N_26947,N_24404,N_24552);
nor U26948 (N_26948,N_25067,N_25037);
xor U26949 (N_26949,N_25040,N_25134);
xor U26950 (N_26950,N_25387,N_24939);
or U26951 (N_26951,N_24344,N_24159);
xor U26952 (N_26952,N_24087,N_24751);
or U26953 (N_26953,N_24206,N_24765);
or U26954 (N_26954,N_25072,N_24455);
xor U26955 (N_26955,N_24270,N_24806);
nand U26956 (N_26956,N_24847,N_24363);
or U26957 (N_26957,N_24396,N_24627);
or U26958 (N_26958,N_24629,N_25393);
nor U26959 (N_26959,N_25492,N_24973);
nand U26960 (N_26960,N_24090,N_25062);
and U26961 (N_26961,N_24207,N_24206);
xor U26962 (N_26962,N_24928,N_24697);
xnor U26963 (N_26963,N_25232,N_25331);
xnor U26964 (N_26964,N_24965,N_24234);
nand U26965 (N_26965,N_24869,N_25439);
nor U26966 (N_26966,N_24144,N_24833);
and U26967 (N_26967,N_24585,N_24645);
nand U26968 (N_26968,N_24579,N_25086);
or U26969 (N_26969,N_24593,N_25224);
nor U26970 (N_26970,N_24589,N_24193);
or U26971 (N_26971,N_24640,N_25327);
xnor U26972 (N_26972,N_25231,N_24402);
nor U26973 (N_26973,N_24750,N_24403);
nor U26974 (N_26974,N_24868,N_24686);
xor U26975 (N_26975,N_25059,N_25189);
and U26976 (N_26976,N_25425,N_24121);
nand U26977 (N_26977,N_25349,N_24366);
nor U26978 (N_26978,N_24584,N_24838);
xnor U26979 (N_26979,N_25332,N_25154);
xor U26980 (N_26980,N_24550,N_24215);
nor U26981 (N_26981,N_24744,N_24310);
xnor U26982 (N_26982,N_25084,N_24029);
or U26983 (N_26983,N_25103,N_24438);
and U26984 (N_26984,N_25484,N_25391);
xor U26985 (N_26985,N_24294,N_24097);
xor U26986 (N_26986,N_25109,N_24932);
nor U26987 (N_26987,N_25497,N_24473);
xnor U26988 (N_26988,N_24968,N_24454);
or U26989 (N_26989,N_24307,N_25389);
or U26990 (N_26990,N_25467,N_24631);
and U26991 (N_26991,N_25276,N_25490);
or U26992 (N_26992,N_24399,N_24662);
xnor U26993 (N_26993,N_25486,N_25346);
xnor U26994 (N_26994,N_24524,N_25098);
or U26995 (N_26995,N_24542,N_24201);
nand U26996 (N_26996,N_24547,N_24558);
xnor U26997 (N_26997,N_24021,N_25161);
nor U26998 (N_26998,N_24342,N_25342);
or U26999 (N_26999,N_24183,N_24144);
or U27000 (N_27000,N_26663,N_26617);
nor U27001 (N_27001,N_26272,N_26987);
nor U27002 (N_27002,N_25696,N_26571);
and U27003 (N_27003,N_26248,N_26463);
nand U27004 (N_27004,N_25551,N_26373);
or U27005 (N_27005,N_26243,N_25978);
nor U27006 (N_27006,N_26685,N_26730);
nand U27007 (N_27007,N_25744,N_25657);
and U27008 (N_27008,N_25732,N_25532);
and U27009 (N_27009,N_26060,N_26482);
or U27010 (N_27010,N_25623,N_26344);
xor U27011 (N_27011,N_26219,N_25812);
or U27012 (N_27012,N_26902,N_26061);
nor U27013 (N_27013,N_26895,N_26378);
or U27014 (N_27014,N_26704,N_25603);
nor U27015 (N_27015,N_26072,N_26599);
and U27016 (N_27016,N_26891,N_25935);
xor U27017 (N_27017,N_25593,N_26581);
nor U27018 (N_27018,N_25672,N_26129);
xor U27019 (N_27019,N_26466,N_25538);
nand U27020 (N_27020,N_25686,N_26973);
or U27021 (N_27021,N_26448,N_26346);
xor U27022 (N_27022,N_26552,N_25646);
nor U27023 (N_27023,N_26283,N_26253);
nand U27024 (N_27024,N_26406,N_26864);
xor U27025 (N_27025,N_26388,N_26351);
nand U27026 (N_27026,N_26369,N_26013);
and U27027 (N_27027,N_25618,N_26043);
xnor U27028 (N_27028,N_26083,N_25845);
and U27029 (N_27029,N_25960,N_25569);
and U27030 (N_27030,N_26657,N_25836);
nor U27031 (N_27031,N_25644,N_26554);
xor U27032 (N_27032,N_25826,N_26944);
nand U27033 (N_27033,N_25969,N_25785);
xor U27034 (N_27034,N_25681,N_26548);
nor U27035 (N_27035,N_26929,N_26458);
xnor U27036 (N_27036,N_26065,N_26208);
or U27037 (N_27037,N_25582,N_26792);
xor U27038 (N_27038,N_26303,N_26345);
xnor U27039 (N_27039,N_26665,N_26816);
nand U27040 (N_27040,N_25610,N_25757);
nor U27041 (N_27041,N_26756,N_26087);
and U27042 (N_27042,N_26031,N_25799);
nor U27043 (N_27043,N_26744,N_26880);
or U27044 (N_27044,N_26003,N_26115);
nor U27045 (N_27045,N_26680,N_25547);
or U27046 (N_27046,N_25819,N_25879);
or U27047 (N_27047,N_26338,N_25662);
and U27048 (N_27048,N_26920,N_26307);
nand U27049 (N_27049,N_26728,N_26370);
nand U27050 (N_27050,N_26313,N_25922);
xnor U27051 (N_27051,N_26337,N_26343);
xor U27052 (N_27052,N_25651,N_25703);
nor U27053 (N_27053,N_26385,N_25803);
nand U27054 (N_27054,N_26037,N_26726);
nor U27055 (N_27055,N_26504,N_26761);
xor U27056 (N_27056,N_26190,N_26855);
nand U27057 (N_27057,N_25984,N_26330);
xnor U27058 (N_27058,N_25876,N_26681);
nor U27059 (N_27059,N_26125,N_26171);
xor U27060 (N_27060,N_26032,N_25938);
nor U27061 (N_27061,N_25924,N_25509);
xnor U27062 (N_27062,N_26804,N_25758);
nand U27063 (N_27063,N_26425,N_26091);
or U27064 (N_27064,N_26052,N_26774);
and U27065 (N_27065,N_26019,N_26488);
nand U27066 (N_27066,N_26846,N_26305);
nand U27067 (N_27067,N_26831,N_26152);
and U27068 (N_27068,N_25998,N_26528);
xor U27069 (N_27069,N_25507,N_26834);
xor U27070 (N_27070,N_26945,N_26241);
and U27071 (N_27071,N_25863,N_26908);
xor U27072 (N_27072,N_25883,N_26637);
xor U27073 (N_27073,N_25846,N_26926);
and U27074 (N_27074,N_26712,N_25843);
nor U27075 (N_27075,N_25601,N_26602);
and U27076 (N_27076,N_26047,N_26240);
xnor U27077 (N_27077,N_26955,N_26517);
or U27078 (N_27078,N_26825,N_26262);
nor U27079 (N_27079,N_26718,N_25927);
nand U27080 (N_27080,N_26449,N_26661);
or U27081 (N_27081,N_26158,N_26021);
nor U27082 (N_27082,N_26470,N_26651);
and U27083 (N_27083,N_25536,N_25606);
and U27084 (N_27084,N_26779,N_25902);
nor U27085 (N_27085,N_25944,N_26906);
and U27086 (N_27086,N_26269,N_25660);
nand U27087 (N_27087,N_25663,N_26672);
nand U27088 (N_27088,N_26450,N_25760);
or U27089 (N_27089,N_25629,N_26803);
and U27090 (N_27090,N_25736,N_25788);
nor U27091 (N_27091,N_26411,N_26145);
or U27092 (N_27092,N_26819,N_26209);
or U27093 (N_27093,N_26678,N_26191);
and U27094 (N_27094,N_26278,N_25526);
nor U27095 (N_27095,N_25950,N_26772);
and U27096 (N_27096,N_26156,N_25945);
xor U27097 (N_27097,N_26359,N_26348);
and U27098 (N_27098,N_25572,N_26745);
or U27099 (N_27099,N_26592,N_25670);
xnor U27100 (N_27100,N_26192,N_25802);
and U27101 (N_27101,N_26994,N_25926);
or U27102 (N_27102,N_26312,N_26644);
nor U27103 (N_27103,N_26067,N_25896);
nor U27104 (N_27104,N_26384,N_25825);
nor U27105 (N_27105,N_26620,N_26252);
nor U27106 (N_27106,N_25971,N_26491);
and U27107 (N_27107,N_26120,N_26214);
and U27108 (N_27108,N_25913,N_26329);
nand U27109 (N_27109,N_26735,N_26877);
nor U27110 (N_27110,N_25999,N_26092);
nand U27111 (N_27111,N_26499,N_26341);
nand U27112 (N_27112,N_25828,N_25989);
nand U27113 (N_27113,N_25914,N_25722);
nor U27114 (N_27114,N_26520,N_26058);
nand U27115 (N_27115,N_25577,N_26628);
and U27116 (N_27116,N_26766,N_25514);
and U27117 (N_27117,N_25554,N_26597);
or U27118 (N_27118,N_26130,N_25553);
nor U27119 (N_27119,N_26195,N_26197);
nand U27120 (N_27120,N_26633,N_25980);
and U27121 (N_27121,N_26386,N_26234);
or U27122 (N_27122,N_25987,N_26818);
nand U27123 (N_27123,N_25833,N_26451);
and U27124 (N_27124,N_26161,N_26551);
nand U27125 (N_27125,N_25648,N_25979);
nor U27126 (N_27126,N_26703,N_26569);
and U27127 (N_27127,N_26649,N_25767);
nor U27128 (N_27128,N_26311,N_25740);
xnor U27129 (N_27129,N_25626,N_25977);
nor U27130 (N_27130,N_26280,N_25874);
and U27131 (N_27131,N_25542,N_25907);
nor U27132 (N_27132,N_26547,N_26453);
and U27133 (N_27133,N_26524,N_26939);
xor U27134 (N_27134,N_25659,N_25649);
nand U27135 (N_27135,N_26350,N_26108);
and U27136 (N_27136,N_26439,N_26423);
xor U27137 (N_27137,N_26276,N_25937);
or U27138 (N_27138,N_25993,N_26096);
and U27139 (N_27139,N_25673,N_26695);
nor U27140 (N_27140,N_25511,N_26967);
and U27141 (N_27141,N_26655,N_26498);
nand U27142 (N_27142,N_26110,N_26776);
nor U27143 (N_27143,N_26155,N_26900);
nand U27144 (N_27144,N_26437,N_26005);
nand U27145 (N_27145,N_26507,N_26268);
nor U27146 (N_27146,N_26500,N_25966);
xor U27147 (N_27147,N_26221,N_26188);
xor U27148 (N_27148,N_26217,N_26461);
nand U27149 (N_27149,N_25705,N_26583);
xor U27150 (N_27150,N_26873,N_26459);
and U27151 (N_27151,N_26057,N_26071);
nand U27152 (N_27152,N_26114,N_26187);
or U27153 (N_27153,N_26090,N_25591);
or U27154 (N_27154,N_25534,N_26297);
and U27155 (N_27155,N_25587,N_26296);
nor U27156 (N_27156,N_26646,N_26558);
nand U27157 (N_27157,N_26101,N_26505);
and U27158 (N_27158,N_26477,N_25602);
nor U27159 (N_27159,N_25682,N_25844);
xor U27160 (N_27160,N_26749,N_26412);
xor U27161 (N_27161,N_26164,N_25710);
or U27162 (N_27162,N_26143,N_26805);
or U27163 (N_27163,N_25640,N_26121);
nand U27164 (N_27164,N_26839,N_26431);
and U27165 (N_27165,N_26023,N_26142);
nor U27166 (N_27166,N_26426,N_25986);
xor U27167 (N_27167,N_26710,N_26075);
nor U27168 (N_27168,N_26850,N_26795);
nor U27169 (N_27169,N_26235,N_25574);
xor U27170 (N_27170,N_26227,N_25735);
nand U27171 (N_27171,N_26629,N_26686);
nand U27172 (N_27172,N_26225,N_26487);
nand U27173 (N_27173,N_26079,N_26490);
nand U27174 (N_27174,N_26591,N_26715);
nand U27175 (N_27175,N_25861,N_25747);
nand U27176 (N_27176,N_25880,N_26399);
xor U27177 (N_27177,N_25677,N_26961);
nor U27178 (N_27178,N_26882,N_26157);
nor U27179 (N_27179,N_26046,N_26977);
and U27180 (N_27180,N_26200,N_25668);
xor U27181 (N_27181,N_25680,N_25764);
or U27182 (N_27182,N_26347,N_26741);
and U27183 (N_27183,N_26403,N_26577);
nand U27184 (N_27184,N_25704,N_26748);
xnor U27185 (N_27185,N_26247,N_25755);
nand U27186 (N_27186,N_26204,N_26102);
nand U27187 (N_27187,N_25857,N_25807);
nand U27188 (N_27188,N_26522,N_25671);
xnor U27189 (N_27189,N_26233,N_25797);
nor U27190 (N_27190,N_26627,N_26027);
nand U27191 (N_27191,N_25991,N_25598);
nand U27192 (N_27192,N_25974,N_26683);
nand U27193 (N_27193,N_25564,N_26732);
or U27194 (N_27194,N_26717,N_25912);
xnor U27195 (N_27195,N_25639,N_25701);
and U27196 (N_27196,N_26053,N_25652);
and U27197 (N_27197,N_26495,N_26363);
nor U27198 (N_27198,N_25882,N_25821);
or U27199 (N_27199,N_25869,N_26940);
or U27200 (N_27200,N_25552,N_25988);
xnor U27201 (N_27201,N_26731,N_25820);
nor U27202 (N_27202,N_26335,N_25895);
xor U27203 (N_27203,N_26366,N_26184);
xnor U27204 (N_27204,N_25666,N_26324);
xnor U27205 (N_27205,N_26026,N_26327);
xor U27206 (N_27206,N_26572,N_26372);
and U27207 (N_27207,N_26068,N_26136);
nand U27208 (N_27208,N_25533,N_26601);
nor U27209 (N_27209,N_26632,N_25868);
or U27210 (N_27210,N_26625,N_25872);
nor U27211 (N_27211,N_25725,N_26442);
nand U27212 (N_27212,N_26754,N_26189);
xor U27213 (N_27213,N_25630,N_25523);
or U27214 (N_27214,N_25588,N_26829);
nand U27215 (N_27215,N_25516,N_26688);
nor U27216 (N_27216,N_26857,N_26727);
and U27217 (N_27217,N_25995,N_26802);
xnor U27218 (N_27218,N_26706,N_26094);
xor U27219 (N_27219,N_26010,N_26078);
xor U27220 (N_27220,N_26736,N_26393);
or U27221 (N_27221,N_26465,N_26475);
nand U27222 (N_27222,N_26070,N_26218);
xnor U27223 (N_27223,N_25904,N_26132);
and U27224 (N_27224,N_26245,N_26964);
and U27225 (N_27225,N_26401,N_26780);
or U27226 (N_27226,N_25724,N_26721);
or U27227 (N_27227,N_25518,N_26340);
nor U27228 (N_27228,N_26468,N_26045);
xor U27229 (N_27229,N_26796,N_26954);
and U27230 (N_27230,N_26974,N_26028);
nand U27231 (N_27231,N_25707,N_26516);
nor U27232 (N_27232,N_26981,N_26170);
or U27233 (N_27233,N_26525,N_26916);
and U27234 (N_27234,N_25555,N_26354);
and U27235 (N_27235,N_26968,N_26995);
nand U27236 (N_27236,N_25579,N_25996);
nor U27237 (N_27237,N_26565,N_26452);
and U27238 (N_27238,N_25787,N_26445);
nor U27239 (N_27239,N_25624,N_26871);
xnor U27240 (N_27240,N_26174,N_25834);
xnor U27241 (N_27241,N_26287,N_26733);
or U27242 (N_27242,N_26404,N_26224);
xor U27243 (N_27243,N_26652,N_25576);
nand U27244 (N_27244,N_25699,N_25911);
xnor U27245 (N_27245,N_26725,N_25645);
and U27246 (N_27246,N_26543,N_26951);
nor U27247 (N_27247,N_26589,N_26508);
or U27248 (N_27248,N_26865,N_25505);
xor U27249 (N_27249,N_26654,N_26687);
xor U27250 (N_27250,N_25730,N_25906);
xnor U27251 (N_27251,N_26063,N_26511);
and U27252 (N_27252,N_25708,N_25631);
and U27253 (N_27253,N_25885,N_26844);
or U27254 (N_27254,N_25992,N_26014);
and U27255 (N_27255,N_26642,N_25875);
and U27256 (N_27256,N_26367,N_26660);
or U27257 (N_27257,N_26462,N_26467);
or U27258 (N_27258,N_26407,N_25809);
and U27259 (N_27259,N_26986,N_26640);
nor U27260 (N_27260,N_25822,N_25786);
nand U27261 (N_27261,N_26938,N_26086);
xor U27262 (N_27262,N_26619,N_26910);
or U27263 (N_27263,N_25831,N_25625);
or U27264 (N_27264,N_26787,N_26390);
and U27265 (N_27265,N_26124,N_25908);
xnor U27266 (N_27266,N_26263,N_26700);
nand U27267 (N_27267,N_26009,N_26051);
or U27268 (N_27268,N_25897,N_25595);
and U27269 (N_27269,N_25684,N_26206);
nand U27270 (N_27270,N_25762,N_26867);
or U27271 (N_27271,N_26321,N_26635);
nand U27272 (N_27272,N_26118,N_25638);
nand U27273 (N_27273,N_26549,N_25801);
or U27274 (N_27274,N_26435,N_26203);
and U27275 (N_27275,N_25535,N_26755);
or U27276 (N_27276,N_26811,N_26285);
and U27277 (N_27277,N_26863,N_25756);
xnor U27278 (N_27278,N_26631,N_25866);
nand U27279 (N_27279,N_26006,N_26237);
xnor U27280 (N_27280,N_25530,N_25859);
and U27281 (N_27281,N_26116,N_26676);
nand U27282 (N_27282,N_26719,N_25543);
and U27283 (N_27283,N_26165,N_26395);
or U27284 (N_27284,N_26626,N_26705);
nand U27285 (N_27285,N_25774,N_25581);
nor U27286 (N_27286,N_26178,N_26007);
and U27287 (N_27287,N_25600,N_26849);
or U27288 (N_27288,N_26998,N_26778);
or U27289 (N_27289,N_26643,N_26220);
nand U27290 (N_27290,N_25900,N_25546);
nand U27291 (N_27291,N_26255,N_25550);
xnor U27292 (N_27292,N_26762,N_25584);
and U27293 (N_27293,N_25613,N_25818);
nand U27294 (N_27294,N_25813,N_26742);
and U27295 (N_27295,N_26653,N_26515);
nor U27296 (N_27296,N_26033,N_26941);
nand U27297 (N_27297,N_26133,N_26561);
or U27298 (N_27298,N_25743,N_25678);
or U27299 (N_27299,N_26568,N_26471);
and U27300 (N_27300,N_25622,N_26903);
xor U27301 (N_27301,N_26375,N_26647);
xnor U27302 (N_27302,N_25571,N_25531);
nor U27303 (N_27303,N_26207,N_25712);
nand U27304 (N_27304,N_25641,N_26966);
nand U27305 (N_27305,N_25519,N_26593);
or U27306 (N_27306,N_26257,N_25777);
nor U27307 (N_27307,N_26937,N_26925);
nor U27308 (N_27308,N_25715,N_25731);
or U27309 (N_27309,N_25634,N_26172);
nor U27310 (N_27310,N_26291,N_26914);
xor U27311 (N_27311,N_25515,N_26809);
nand U27312 (N_27312,N_25941,N_26794);
or U27313 (N_27313,N_26841,N_26290);
and U27314 (N_27314,N_26833,N_26506);
nand U27315 (N_27315,N_26519,N_26440);
and U27316 (N_27316,N_25964,N_26314);
or U27317 (N_27317,N_26334,N_25899);
xnor U27318 (N_27318,N_26739,N_25720);
and U27319 (N_27319,N_25847,N_25665);
and U27320 (N_27320,N_26239,N_26526);
nand U27321 (N_27321,N_26131,N_26898);
xor U27322 (N_27322,N_25607,N_25881);
and U27323 (N_27323,N_25842,N_26797);
or U27324 (N_27324,N_26163,N_26146);
and U27325 (N_27325,N_25617,N_25794);
nand U27326 (N_27326,N_26398,N_26952);
nand U27327 (N_27327,N_26302,N_26907);
nand U27328 (N_27328,N_26684,N_26746);
or U27329 (N_27329,N_26722,N_25967);
and U27330 (N_27330,N_25939,N_25916);
and U27331 (N_27331,N_25517,N_26881);
or U27332 (N_27332,N_26924,N_25942);
or U27333 (N_27333,N_25647,N_25580);
nand U27334 (N_27334,N_26082,N_26638);
nand U27335 (N_27335,N_26041,N_26383);
or U27336 (N_27336,N_25628,N_26605);
xnor U27337 (N_27337,N_25814,N_26623);
xor U27338 (N_27338,N_25537,N_26144);
nand U27339 (N_27339,N_26521,N_26897);
xor U27340 (N_27340,N_26325,N_26576);
nor U27341 (N_27341,N_26004,N_26402);
xnor U27342 (N_27342,N_26381,N_25775);
nand U27343 (N_27343,N_26409,N_26256);
xor U27344 (N_27344,N_26673,N_25653);
or U27345 (N_27345,N_26230,N_26799);
and U27346 (N_27346,N_26702,N_26523);
nand U27347 (N_27347,N_26064,N_26948);
or U27348 (N_27348,N_26358,N_26538);
xor U27349 (N_27349,N_26847,N_26711);
xnor U27350 (N_27350,N_25759,N_25763);
nand U27351 (N_27351,N_25697,N_26949);
and U27352 (N_27352,N_26899,N_26614);
xnor U27353 (N_27353,N_26969,N_26609);
nor U27354 (N_27354,N_25959,N_26943);
nand U27355 (N_27355,N_26109,N_26229);
nand U27356 (N_27356,N_26532,N_26339);
xnor U27357 (N_27357,N_25864,N_26213);
nor U27358 (N_27358,N_26387,N_26970);
xor U27359 (N_27359,N_26682,N_25521);
and U27360 (N_27360,N_26122,N_26277);
or U27361 (N_27361,N_26894,N_26408);
and U27362 (N_27362,N_26073,N_26616);
nor U27363 (N_27363,N_26273,N_26374);
nor U27364 (N_27364,N_26259,N_25962);
nand U27365 (N_27365,N_26852,N_26786);
xnor U27366 (N_27366,N_25621,N_26734);
xor U27367 (N_27367,N_26936,N_26472);
or U27368 (N_27368,N_25557,N_26615);
and U27369 (N_27369,N_26141,N_26985);
and U27370 (N_27370,N_25685,N_26555);
or U27371 (N_27371,N_26317,N_25510);
nand U27372 (N_27372,N_26413,N_26858);
and U27373 (N_27373,N_26333,N_26030);
nor U27374 (N_27374,N_25718,N_26231);
and U27375 (N_27375,N_26074,N_25965);
and U27376 (N_27376,N_26077,N_26062);
and U27377 (N_27377,N_26747,N_26024);
xnor U27378 (N_27378,N_25540,N_26604);
and U27379 (N_27379,N_25632,N_25958);
or U27380 (N_27380,N_26432,N_26832);
nor U27381 (N_27381,N_26757,N_26579);
and U27382 (N_27382,N_25816,N_25561);
or U27383 (N_27383,N_26677,N_26768);
xor U27384 (N_27384,N_26807,N_26137);
and U27385 (N_27385,N_26529,N_26199);
xnor U27386 (N_27386,N_26080,N_25596);
or U27387 (N_27387,N_25549,N_26275);
and U27388 (N_27388,N_26223,N_25727);
or U27389 (N_27389,N_26281,N_26999);
xnor U27390 (N_27390,N_26216,N_26148);
xor U27391 (N_27391,N_25956,N_26585);
or U27392 (N_27392,N_25806,N_25951);
and U27393 (N_27393,N_26845,N_25811);
nor U27394 (N_27394,N_26265,N_26460);
or U27395 (N_27395,N_25525,N_25943);
nor U27396 (N_27396,N_26098,N_26698);
nand U27397 (N_27397,N_26667,N_25709);
nor U27398 (N_27398,N_26194,N_26443);
nor U27399 (N_27399,N_26656,N_26574);
or U27400 (N_27400,N_26055,N_26671);
or U27401 (N_27401,N_26645,N_26915);
nand U27402 (N_27402,N_25862,N_26421);
and U27403 (N_27403,N_25506,N_26479);
and U27404 (N_27404,N_26557,N_25877);
and U27405 (N_27405,N_26536,N_26580);
nand U27406 (N_27406,N_26419,N_26455);
and U27407 (N_27407,N_26868,N_25783);
and U27408 (N_27408,N_25837,N_26489);
xnor U27409 (N_27409,N_25661,N_26621);
xor U27410 (N_27410,N_26160,N_25889);
xnor U27411 (N_27411,N_25545,N_26927);
and U27412 (N_27412,N_26493,N_26397);
or U27413 (N_27413,N_26691,N_26919);
xnor U27414 (N_27414,N_26389,N_26578);
and U27415 (N_27415,N_26696,N_26806);
or U27416 (N_27416,N_25560,N_26759);
xnor U27417 (N_27417,N_26128,N_25751);
xnor U27418 (N_27418,N_26167,N_26166);
xnor U27419 (N_27419,N_25856,N_26533);
nand U27420 (N_27420,N_26586,N_26016);
xor U27421 (N_27421,N_26959,N_26182);
nor U27422 (N_27422,N_26922,N_26872);
or U27423 (N_27423,N_26613,N_26228);
nand U27424 (N_27424,N_25796,N_26634);
or U27425 (N_27425,N_25815,N_26469);
xnor U27426 (N_27426,N_26510,N_26879);
nand U27427 (N_27427,N_25508,N_25589);
nand U27428 (N_27428,N_26991,N_26226);
xnor U27429 (N_27429,N_26662,N_26352);
xnor U27430 (N_27430,N_26149,N_26674);
and U27431 (N_27431,N_26035,N_26564);
xor U27432 (N_27432,N_25690,N_26414);
nand U27433 (N_27433,N_25539,N_26921);
xor U27434 (N_27434,N_26410,N_25575);
xnor U27435 (N_27435,N_26624,N_26002);
or U27436 (N_27436,N_25841,N_26556);
nor U27437 (N_27437,N_25592,N_26901);
or U27438 (N_27438,N_26485,N_26464);
or U27439 (N_27439,N_26048,N_25669);
nor U27440 (N_27440,N_26183,N_26288);
nor U27441 (N_27441,N_25749,N_26990);
nand U27442 (N_27442,N_26509,N_25698);
nor U27443 (N_27443,N_25655,N_26892);
and U27444 (N_27444,N_26567,N_25568);
nor U27445 (N_27445,N_25976,N_25700);
xnor U27446 (N_27446,N_26546,N_26689);
nor U27447 (N_27447,N_25766,N_26238);
and U27448 (N_27448,N_25983,N_26396);
or U27449 (N_27449,N_26843,N_25562);
nor U27450 (N_27450,N_25597,N_25910);
nor U27451 (N_27451,N_26758,N_25573);
nand U27452 (N_27452,N_26669,N_26293);
nand U27453 (N_27453,N_25503,N_25892);
nand U27454 (N_27454,N_25544,N_26198);
nor U27455 (N_27455,N_25702,N_26553);
or U27456 (N_27456,N_26284,N_25605);
xor U27457 (N_27457,N_26885,N_26417);
nand U27458 (N_27458,N_26588,N_25947);
nor U27459 (N_27459,N_25541,N_26416);
xnor U27460 (N_27460,N_26769,N_25693);
nand U27461 (N_27461,N_26049,N_26054);
and U27462 (N_27462,N_26315,N_25905);
and U27463 (N_27463,N_25848,N_25556);
nor U27464 (N_27464,N_26473,N_26600);
or U27465 (N_27465,N_26153,N_25878);
xnor U27466 (N_27466,N_26947,N_26486);
nor U27467 (N_27467,N_26205,N_25920);
xor U27468 (N_27468,N_26884,N_26518);
or U27469 (N_27469,N_25890,N_26169);
and U27470 (N_27470,N_26279,N_25716);
or U27471 (N_27471,N_25770,N_26050);
nor U27472 (N_27472,N_25734,N_26428);
xor U27473 (N_27473,N_25804,N_25524);
nor U27474 (N_27474,N_26988,N_25578);
nor U27475 (N_27475,N_26784,N_26760);
or U27476 (N_27476,N_25635,N_25620);
or U27477 (N_27477,N_26371,N_25952);
nand U27478 (N_27478,N_26851,N_26394);
nor U27479 (N_27479,N_26740,N_26770);
and U27480 (N_27480,N_26001,N_25955);
nand U27481 (N_27481,N_25817,N_25567);
nand U27482 (N_27482,N_26382,N_26095);
xor U27483 (N_27483,N_26815,N_26424);
or U27484 (N_27484,N_26038,N_25687);
nor U27485 (N_27485,N_26029,N_26353);
and U27486 (N_27486,N_26817,N_26971);
xor U27487 (N_27487,N_25838,N_26713);
nand U27488 (N_27488,N_26878,N_25745);
and U27489 (N_27489,N_26692,N_25683);
xnor U27490 (N_27490,N_25961,N_26789);
and U27491 (N_27491,N_26942,N_26232);
nand U27492 (N_27492,N_26022,N_25772);
nand U27493 (N_27493,N_26931,N_26295);
xor U27494 (N_27494,N_25870,N_25768);
and U27495 (N_27495,N_26008,N_25898);
and U27496 (N_27496,N_25765,N_25795);
and U27497 (N_27497,N_26222,N_26069);
nand U27498 (N_27498,N_26309,N_26151);
or U27499 (N_27499,N_26679,N_25840);
xor U27500 (N_27500,N_25789,N_26211);
or U27501 (N_27501,N_26636,N_26765);
or U27502 (N_27502,N_25750,N_25779);
nor U27503 (N_27503,N_26400,N_26310);
nor U27504 (N_27504,N_26059,N_25667);
or U27505 (N_27505,N_25798,N_25590);
and U27506 (N_27506,N_26377,N_25643);
nor U27507 (N_27507,N_26356,N_25917);
nand U27508 (N_27508,N_26360,N_25719);
and U27509 (N_27509,N_26590,N_26801);
or U27510 (N_27510,N_26446,N_25808);
nand U27511 (N_27511,N_26928,N_25865);
xnor U27512 (N_27512,N_26039,N_25504);
nor U27513 (N_27513,N_26853,N_26810);
or U27514 (N_27514,N_25746,N_26606);
and U27515 (N_27515,N_26162,N_25921);
nand U27516 (N_27516,N_25753,N_26821);
xor U27517 (N_27517,N_25949,N_26953);
nand U27518 (N_27518,N_26117,N_26773);
xor U27519 (N_27519,N_25994,N_26582);
nor U27520 (N_27520,N_26168,N_25741);
nor U27521 (N_27521,N_26011,N_26497);
and U27522 (N_27522,N_26201,N_25711);
nand U27523 (N_27523,N_26392,N_25559);
nand U27524 (N_27524,N_25527,N_25565);
and U27525 (N_27525,N_26550,N_25930);
nand U27526 (N_27526,N_26542,N_26539);
and U27527 (N_27527,N_26427,N_26598);
or U27528 (N_27528,N_26530,N_25891);
nand U27529 (N_27529,N_26368,N_26699);
and U27530 (N_27530,N_26134,N_26044);
xnor U27531 (N_27531,N_26319,N_26481);
and U27532 (N_27532,N_26537,N_26707);
and U27533 (N_27533,N_26242,N_26859);
or U27534 (N_27534,N_26862,N_25793);
xnor U27535 (N_27535,N_25805,N_26176);
nor U27536 (N_27536,N_25773,N_26015);
and U27537 (N_27537,N_26250,N_25776);
nand U27538 (N_27538,N_26668,N_26202);
nor U27539 (N_27539,N_26965,N_25835);
nand U27540 (N_27540,N_25501,N_25928);
or U27541 (N_27541,N_26186,N_26887);
nand U27542 (N_27542,N_25933,N_25633);
or U27543 (N_27543,N_26720,N_25609);
nor U27544 (N_27544,N_25827,N_26308);
or U27545 (N_27545,N_26418,N_26750);
xor U27546 (N_27546,N_26112,N_26336);
or U27547 (N_27547,N_26854,N_26531);
or U27548 (N_27548,N_26215,N_26105);
and U27549 (N_27549,N_26603,N_26000);
xnor U27550 (N_27550,N_25985,N_26886);
xnor U27551 (N_27551,N_25761,N_26982);
nand U27552 (N_27552,N_26181,N_26534);
nor U27553 (N_27553,N_26984,N_25970);
or U27554 (N_27554,N_25997,N_26081);
nor U27555 (N_27555,N_26540,N_26912);
nor U27556 (N_27556,N_25713,N_25782);
or U27557 (N_27557,N_26147,N_25679);
xnor U27558 (N_27558,N_26861,N_25901);
nor U27559 (N_27559,N_26956,N_26494);
nand U27560 (N_27560,N_26261,N_26650);
xor U27561 (N_27561,N_26788,N_25903);
and U27562 (N_27562,N_25717,N_25733);
nand U27563 (N_27563,N_26690,N_26512);
xnor U27564 (N_27564,N_26570,N_26249);
xnor U27565 (N_27565,N_26180,N_25729);
and U27566 (N_27566,N_26751,N_25873);
nand U27567 (N_27567,N_26298,N_26405);
nor U27568 (N_27568,N_26798,N_25723);
nand U27569 (N_27569,N_26017,N_26355);
nor U27570 (N_27570,N_25721,N_26874);
or U27571 (N_27571,N_26433,N_26391);
or U27572 (N_27572,N_26436,N_26274);
or U27573 (N_27573,N_25934,N_26830);
or U27574 (N_27574,N_26913,N_26210);
xor U27575 (N_27575,N_25594,N_26890);
or U27576 (N_27576,N_26342,N_26150);
nor U27577 (N_27577,N_26138,N_25931);
and U27578 (N_27578,N_26738,N_26267);
and U27579 (N_27579,N_26869,N_26587);
nand U27580 (N_27580,N_26483,N_25611);
or U27581 (N_27581,N_26379,N_25654);
or U27582 (N_27582,N_26103,N_26978);
nor U27583 (N_27583,N_26828,N_26575);
or U27584 (N_27584,N_25982,N_25918);
and U27585 (N_27585,N_26791,N_26905);
nor U27586 (N_27586,N_26478,N_26088);
xnor U27587 (N_27587,N_26270,N_26958);
and U27588 (N_27588,N_25851,N_26800);
nand U27589 (N_27589,N_26771,N_26454);
or U27590 (N_27590,N_26608,N_25692);
xor U27591 (N_27591,N_26827,N_26318);
xor U27592 (N_27592,N_25963,N_26502);
nand U27593 (N_27593,N_25919,N_26447);
nand U27594 (N_27594,N_26997,N_26610);
nand U27595 (N_27595,N_26848,N_25612);
or U27596 (N_27596,N_26664,N_25664);
nor U27597 (N_27597,N_26093,N_26697);
nand U27598 (N_27598,N_26976,N_26870);
nand U27599 (N_27599,N_25791,N_26056);
xor U27600 (N_27600,N_26630,N_26993);
or U27601 (N_27601,N_26618,N_26767);
and U27602 (N_27602,N_26709,N_26496);
nand U27603 (N_27603,N_25566,N_26896);
xnor U27604 (N_27604,N_26783,N_26962);
or U27605 (N_27605,N_25909,N_26289);
nor U27606 (N_27606,N_26782,N_25691);
nand U27607 (N_27607,N_25695,N_25867);
and U27608 (N_27608,N_26127,N_26266);
or U27609 (N_27609,N_26299,N_25855);
or U27610 (N_27610,N_26992,N_25599);
and U27611 (N_27611,N_26365,N_25925);
nand U27612 (N_27612,N_26573,N_26975);
or U27613 (N_27613,N_26701,N_25754);
xor U27614 (N_27614,N_26563,N_25946);
xor U27615 (N_27615,N_26753,N_26492);
nand U27616 (N_27616,N_26139,N_26126);
and U27617 (N_27617,N_26904,N_25502);
and U27618 (N_27618,N_26934,N_26775);
nand U27619 (N_27619,N_26434,N_26996);
xnor U27620 (N_27620,N_26380,N_25886);
nand U27621 (N_27621,N_26785,N_26244);
nor U27622 (N_27622,N_26527,N_26930);
nor U27623 (N_27623,N_26326,N_25784);
or U27624 (N_27624,N_25500,N_26935);
and U27625 (N_27625,N_26856,N_26097);
nor U27626 (N_27626,N_26866,N_26875);
and U27627 (N_27627,N_26193,N_26559);
and U27628 (N_27628,N_25706,N_25824);
or U27629 (N_27629,N_25688,N_26842);
and U27630 (N_27630,N_26781,N_26254);
and U27631 (N_27631,N_25830,N_25742);
xor U27632 (N_27632,N_26484,N_26876);
and U27633 (N_27633,N_25650,N_26331);
or U27634 (N_27634,N_25769,N_26271);
nor U27635 (N_27635,N_26979,N_26659);
or U27636 (N_27636,N_26476,N_26107);
nand U27637 (N_27637,N_26430,N_25570);
and U27638 (N_27638,N_26123,N_26541);
or U27639 (N_27639,N_25888,N_26076);
nor U27640 (N_27640,N_26179,N_26420);
xor U27641 (N_27641,N_26888,N_25860);
nand U27642 (N_27642,N_26544,N_26159);
or U27643 (N_27643,N_26584,N_26918);
xnor U27644 (N_27644,N_25975,N_26264);
nor U27645 (N_27645,N_25513,N_25829);
nor U27646 (N_27646,N_26514,N_26622);
nor U27647 (N_27647,N_26306,N_26972);
nand U27648 (N_27648,N_26826,N_26361);
nor U27649 (N_27649,N_26566,N_25675);
and U27650 (N_27650,N_25522,N_25953);
or U27651 (N_27651,N_26752,N_25957);
and U27652 (N_27652,N_25694,N_26670);
or U27653 (N_27653,N_26560,N_26596);
nand U27654 (N_27654,N_26456,N_26480);
and U27655 (N_27655,N_25585,N_25853);
nor U27656 (N_27656,N_26212,N_25627);
and U27657 (N_27657,N_26175,N_26813);
nor U27658 (N_27658,N_25832,N_25714);
and U27659 (N_27659,N_26362,N_26036);
xor U27660 (N_27660,N_25929,N_25923);
nor U27661 (N_27661,N_26562,N_26840);
and U27662 (N_27662,N_26357,N_26135);
and U27663 (N_27663,N_26814,N_26177);
xnor U27664 (N_27664,N_26763,N_26777);
xnor U27665 (N_27665,N_26724,N_25528);
nor U27666 (N_27666,N_25936,N_26950);
xnor U27667 (N_27667,N_25849,N_25940);
or U27668 (N_27668,N_26893,N_25968);
or U27669 (N_27669,N_25656,N_25800);
and U27670 (N_27670,N_26983,N_26328);
nor U27671 (N_27671,N_25615,N_26708);
nand U27672 (N_27672,N_25973,N_25674);
xnor U27673 (N_27673,N_25990,N_26932);
nor U27674 (N_27674,N_25894,N_25778);
and U27675 (N_27675,N_26611,N_25932);
and U27676 (N_27676,N_25728,N_25972);
xnor U27677 (N_27677,N_26364,N_25752);
or U27678 (N_27678,N_25676,N_26909);
xnor U27679 (N_27679,N_25529,N_26648);
xnor U27680 (N_27680,N_26104,N_26812);
nand U27681 (N_27681,N_26185,N_26594);
or U27682 (N_27682,N_26085,N_25852);
nor U27683 (N_27683,N_26764,N_26154);
nand U27684 (N_27684,N_26119,N_26089);
nor U27685 (N_27685,N_26444,N_26111);
nand U27686 (N_27686,N_26173,N_26933);
xnor U27687 (N_27687,N_26474,N_26911);
and U27688 (N_27688,N_26236,N_25636);
nor U27689 (N_27689,N_26883,N_26501);
nand U27690 (N_27690,N_26100,N_26376);
and U27691 (N_27691,N_26737,N_25748);
and U27692 (N_27692,N_26034,N_25823);
or U27693 (N_27693,N_25563,N_26980);
nand U27694 (N_27694,N_26860,N_26282);
xnor U27695 (N_27695,N_25790,N_26535);
and U27696 (N_27696,N_26332,N_26042);
nand U27697 (N_27697,N_26349,N_25548);
xnor U27698 (N_27698,N_26714,N_25780);
nand U27699 (N_27699,N_26675,N_26246);
nand U27700 (N_27700,N_26723,N_26820);
nand U27701 (N_27701,N_26106,N_25887);
and U27702 (N_27702,N_26066,N_25642);
or U27703 (N_27703,N_26196,N_26963);
xor U27704 (N_27704,N_26658,N_26304);
and U27705 (N_27705,N_25981,N_26457);
nand U27706 (N_27706,N_25614,N_25689);
or U27707 (N_27707,N_26793,N_26989);
nand U27708 (N_27708,N_26957,N_26837);
and U27709 (N_27709,N_26824,N_25839);
or U27710 (N_27710,N_25558,N_25739);
nor U27711 (N_27711,N_26020,N_26639);
xnor U27712 (N_27712,N_25637,N_26294);
nor U27713 (N_27713,N_25658,N_25954);
or U27714 (N_27714,N_25619,N_26323);
nand U27715 (N_27715,N_26040,N_26545);
xor U27716 (N_27716,N_26790,N_26838);
xor U27717 (N_27717,N_26258,N_25884);
or U27718 (N_27718,N_26836,N_26917);
and U27719 (N_27719,N_26641,N_25810);
nor U27720 (N_27720,N_26716,N_26018);
nor U27721 (N_27721,N_25858,N_26503);
nor U27722 (N_27722,N_26889,N_25738);
xor U27723 (N_27723,N_26595,N_25586);
and U27724 (N_27724,N_26415,N_25915);
xor U27725 (N_27725,N_25604,N_26251);
xnor U27726 (N_27726,N_26429,N_25520);
xnor U27727 (N_27727,N_26140,N_26025);
or U27728 (N_27728,N_25726,N_26693);
nand U27729 (N_27729,N_26822,N_26946);
xor U27730 (N_27730,N_26808,N_25583);
xor U27731 (N_27731,N_26099,N_26301);
and U27732 (N_27732,N_25948,N_25771);
nand U27733 (N_27733,N_25608,N_25616);
nand U27734 (N_27734,N_26084,N_25512);
nand U27735 (N_27735,N_26322,N_26666);
nand U27736 (N_27736,N_26286,N_26012);
nand U27737 (N_27737,N_26835,N_26729);
nand U27738 (N_27738,N_26438,N_26513);
or U27739 (N_27739,N_25850,N_26292);
xnor U27740 (N_27740,N_26694,N_25854);
or U27741 (N_27741,N_26923,N_26422);
nand U27742 (N_27742,N_26607,N_25737);
nor U27743 (N_27743,N_26960,N_26612);
or U27744 (N_27744,N_26823,N_26300);
and U27745 (N_27745,N_26441,N_25871);
and U27746 (N_27746,N_26113,N_25893);
xnor U27747 (N_27747,N_26320,N_26260);
xor U27748 (N_27748,N_25792,N_26743);
nand U27749 (N_27749,N_25781,N_26316);
or U27750 (N_27750,N_25649,N_26770);
nor U27751 (N_27751,N_26030,N_26015);
nor U27752 (N_27752,N_26188,N_26083);
or U27753 (N_27753,N_26933,N_26114);
xnor U27754 (N_27754,N_25588,N_26787);
or U27755 (N_27755,N_26538,N_26370);
nor U27756 (N_27756,N_26510,N_26305);
nand U27757 (N_27757,N_25519,N_25908);
xor U27758 (N_27758,N_26694,N_26679);
nand U27759 (N_27759,N_26829,N_25783);
or U27760 (N_27760,N_25665,N_25725);
nand U27761 (N_27761,N_26634,N_26566);
and U27762 (N_27762,N_26818,N_25684);
nor U27763 (N_27763,N_26948,N_25968);
nor U27764 (N_27764,N_26705,N_26119);
nand U27765 (N_27765,N_26857,N_26460);
and U27766 (N_27766,N_25775,N_26988);
nand U27767 (N_27767,N_26732,N_26002);
and U27768 (N_27768,N_26500,N_26691);
nor U27769 (N_27769,N_26077,N_25641);
nand U27770 (N_27770,N_25523,N_26578);
nand U27771 (N_27771,N_26466,N_25988);
xnor U27772 (N_27772,N_26241,N_26729);
xor U27773 (N_27773,N_25822,N_26341);
nand U27774 (N_27774,N_25600,N_26476);
xor U27775 (N_27775,N_26084,N_25923);
nor U27776 (N_27776,N_26076,N_25880);
or U27777 (N_27777,N_26294,N_26233);
nand U27778 (N_27778,N_26322,N_25573);
or U27779 (N_27779,N_25550,N_26446);
nand U27780 (N_27780,N_25516,N_26300);
or U27781 (N_27781,N_25587,N_26337);
nand U27782 (N_27782,N_26911,N_26579);
nor U27783 (N_27783,N_26564,N_25523);
nand U27784 (N_27784,N_26559,N_25557);
xor U27785 (N_27785,N_26495,N_26257);
and U27786 (N_27786,N_26490,N_26561);
or U27787 (N_27787,N_25597,N_26343);
or U27788 (N_27788,N_26598,N_25798);
xnor U27789 (N_27789,N_26041,N_26870);
or U27790 (N_27790,N_26052,N_25692);
nand U27791 (N_27791,N_25537,N_25839);
nor U27792 (N_27792,N_25589,N_26110);
nand U27793 (N_27793,N_25927,N_26870);
or U27794 (N_27794,N_25673,N_25872);
nor U27795 (N_27795,N_25701,N_26749);
xnor U27796 (N_27796,N_26776,N_25815);
and U27797 (N_27797,N_26243,N_26111);
xnor U27798 (N_27798,N_25986,N_25680);
and U27799 (N_27799,N_26449,N_26834);
nand U27800 (N_27800,N_26368,N_25683);
or U27801 (N_27801,N_25672,N_26986);
nand U27802 (N_27802,N_25817,N_25864);
or U27803 (N_27803,N_26885,N_25770);
and U27804 (N_27804,N_26352,N_26492);
and U27805 (N_27805,N_25807,N_26302);
xnor U27806 (N_27806,N_26903,N_26062);
or U27807 (N_27807,N_26897,N_26401);
and U27808 (N_27808,N_26294,N_26729);
or U27809 (N_27809,N_25812,N_25556);
nand U27810 (N_27810,N_26554,N_26692);
or U27811 (N_27811,N_25898,N_25816);
xnor U27812 (N_27812,N_26676,N_25669);
nor U27813 (N_27813,N_26768,N_26400);
or U27814 (N_27814,N_25589,N_26195);
nor U27815 (N_27815,N_26960,N_26672);
xor U27816 (N_27816,N_26368,N_26608);
and U27817 (N_27817,N_26716,N_26816);
nor U27818 (N_27818,N_25998,N_25988);
nor U27819 (N_27819,N_26139,N_26612);
xnor U27820 (N_27820,N_26914,N_26890);
nand U27821 (N_27821,N_25666,N_26813);
xor U27822 (N_27822,N_26379,N_26580);
nand U27823 (N_27823,N_26100,N_26185);
and U27824 (N_27824,N_26523,N_26999);
or U27825 (N_27825,N_26614,N_25936);
or U27826 (N_27826,N_25709,N_26422);
and U27827 (N_27827,N_26658,N_26927);
xnor U27828 (N_27828,N_25794,N_26108);
and U27829 (N_27829,N_25610,N_26590);
or U27830 (N_27830,N_26846,N_25513);
nor U27831 (N_27831,N_25636,N_25587);
or U27832 (N_27832,N_26232,N_26490);
xnor U27833 (N_27833,N_26092,N_26547);
or U27834 (N_27834,N_25711,N_25797);
nor U27835 (N_27835,N_26287,N_25566);
or U27836 (N_27836,N_25895,N_25627);
xor U27837 (N_27837,N_25524,N_25939);
and U27838 (N_27838,N_25731,N_25794);
nor U27839 (N_27839,N_26963,N_25894);
or U27840 (N_27840,N_26650,N_26330);
nor U27841 (N_27841,N_26359,N_25513);
xor U27842 (N_27842,N_26499,N_26202);
nor U27843 (N_27843,N_26727,N_26486);
xor U27844 (N_27844,N_25641,N_26547);
or U27845 (N_27845,N_26807,N_26456);
nor U27846 (N_27846,N_25933,N_26714);
and U27847 (N_27847,N_26800,N_26706);
or U27848 (N_27848,N_26977,N_26043);
xor U27849 (N_27849,N_26234,N_26421);
and U27850 (N_27850,N_26906,N_25929);
nand U27851 (N_27851,N_25931,N_26238);
and U27852 (N_27852,N_26789,N_26637);
xor U27853 (N_27853,N_26091,N_25575);
or U27854 (N_27854,N_26390,N_26508);
and U27855 (N_27855,N_26012,N_26483);
and U27856 (N_27856,N_26665,N_26917);
xor U27857 (N_27857,N_26346,N_26404);
nor U27858 (N_27858,N_25589,N_26466);
nand U27859 (N_27859,N_26170,N_26741);
nor U27860 (N_27860,N_25744,N_26137);
and U27861 (N_27861,N_26704,N_26463);
or U27862 (N_27862,N_26510,N_26457);
xor U27863 (N_27863,N_26830,N_25909);
or U27864 (N_27864,N_25665,N_26023);
and U27865 (N_27865,N_26582,N_25829);
xnor U27866 (N_27866,N_26035,N_26614);
nand U27867 (N_27867,N_26012,N_26713);
or U27868 (N_27868,N_26609,N_25825);
and U27869 (N_27869,N_25631,N_26289);
or U27870 (N_27870,N_25654,N_25836);
xnor U27871 (N_27871,N_26992,N_26176);
nand U27872 (N_27872,N_26406,N_26403);
xnor U27873 (N_27873,N_25780,N_25832);
nand U27874 (N_27874,N_25885,N_26858);
xnor U27875 (N_27875,N_26870,N_25962);
nand U27876 (N_27876,N_26783,N_26707);
and U27877 (N_27877,N_25587,N_26822);
or U27878 (N_27878,N_25944,N_25585);
nand U27879 (N_27879,N_25610,N_26211);
nand U27880 (N_27880,N_26771,N_26167);
or U27881 (N_27881,N_26224,N_26436);
and U27882 (N_27882,N_26790,N_26254);
xnor U27883 (N_27883,N_26570,N_25543);
and U27884 (N_27884,N_26217,N_26465);
xnor U27885 (N_27885,N_26863,N_25977);
nor U27886 (N_27886,N_26956,N_25978);
nand U27887 (N_27887,N_25771,N_25883);
and U27888 (N_27888,N_26580,N_26960);
and U27889 (N_27889,N_26001,N_25742);
and U27890 (N_27890,N_26283,N_26202);
nor U27891 (N_27891,N_26758,N_25772);
and U27892 (N_27892,N_26454,N_25828);
and U27893 (N_27893,N_25714,N_26079);
nor U27894 (N_27894,N_26112,N_26014);
nor U27895 (N_27895,N_26893,N_26607);
and U27896 (N_27896,N_25997,N_25884);
nand U27897 (N_27897,N_26618,N_25563);
nand U27898 (N_27898,N_26682,N_26550);
xnor U27899 (N_27899,N_25817,N_26436);
xnor U27900 (N_27900,N_26177,N_26607);
and U27901 (N_27901,N_26087,N_26674);
or U27902 (N_27902,N_26888,N_26391);
nand U27903 (N_27903,N_26483,N_26608);
xnor U27904 (N_27904,N_26247,N_25927);
nor U27905 (N_27905,N_26179,N_25858);
nor U27906 (N_27906,N_25827,N_25610);
or U27907 (N_27907,N_26937,N_26222);
and U27908 (N_27908,N_26416,N_25545);
nor U27909 (N_27909,N_25604,N_26980);
and U27910 (N_27910,N_26408,N_26983);
and U27911 (N_27911,N_25953,N_26948);
or U27912 (N_27912,N_26944,N_26744);
or U27913 (N_27913,N_26745,N_26257);
nand U27914 (N_27914,N_26142,N_26956);
nand U27915 (N_27915,N_26959,N_26245);
or U27916 (N_27916,N_26201,N_25697);
and U27917 (N_27917,N_25700,N_26623);
or U27918 (N_27918,N_26510,N_26143);
xor U27919 (N_27919,N_25785,N_26183);
or U27920 (N_27920,N_25561,N_26623);
nor U27921 (N_27921,N_26930,N_26338);
or U27922 (N_27922,N_26512,N_26064);
and U27923 (N_27923,N_26040,N_26015);
xor U27924 (N_27924,N_26171,N_26214);
nor U27925 (N_27925,N_25969,N_25985);
or U27926 (N_27926,N_26464,N_26284);
xor U27927 (N_27927,N_25537,N_26983);
and U27928 (N_27928,N_26344,N_26708);
nor U27929 (N_27929,N_26324,N_26862);
nand U27930 (N_27930,N_26315,N_26696);
nor U27931 (N_27931,N_26881,N_25898);
and U27932 (N_27932,N_25592,N_25830);
nand U27933 (N_27933,N_26222,N_25777);
or U27934 (N_27934,N_26341,N_26941);
and U27935 (N_27935,N_26948,N_26822);
nand U27936 (N_27936,N_26644,N_25516);
or U27937 (N_27937,N_26779,N_26523);
and U27938 (N_27938,N_26880,N_26416);
and U27939 (N_27939,N_26905,N_26302);
and U27940 (N_27940,N_25838,N_26471);
or U27941 (N_27941,N_25952,N_26701);
nor U27942 (N_27942,N_25733,N_25854);
nor U27943 (N_27943,N_26442,N_26807);
nor U27944 (N_27944,N_26459,N_25597);
or U27945 (N_27945,N_25793,N_25724);
nand U27946 (N_27946,N_26106,N_26501);
xnor U27947 (N_27947,N_26636,N_25949);
nand U27948 (N_27948,N_25763,N_26883);
xor U27949 (N_27949,N_26246,N_26696);
nand U27950 (N_27950,N_26147,N_25940);
xnor U27951 (N_27951,N_25844,N_26924);
nand U27952 (N_27952,N_26543,N_26120);
and U27953 (N_27953,N_26176,N_26475);
xnor U27954 (N_27954,N_26198,N_26599);
nor U27955 (N_27955,N_25524,N_26609);
and U27956 (N_27956,N_25581,N_25549);
xor U27957 (N_27957,N_26886,N_26803);
nor U27958 (N_27958,N_26968,N_26085);
xnor U27959 (N_27959,N_26382,N_26254);
nor U27960 (N_27960,N_26584,N_26546);
nor U27961 (N_27961,N_26806,N_26719);
or U27962 (N_27962,N_25806,N_25751);
xnor U27963 (N_27963,N_26723,N_26101);
and U27964 (N_27964,N_26951,N_26914);
and U27965 (N_27965,N_26268,N_26340);
or U27966 (N_27966,N_26681,N_25568);
nor U27967 (N_27967,N_26104,N_26944);
and U27968 (N_27968,N_26264,N_26482);
nor U27969 (N_27969,N_26720,N_25933);
xor U27970 (N_27970,N_25593,N_26385);
and U27971 (N_27971,N_25969,N_26563);
or U27972 (N_27972,N_26178,N_25861);
or U27973 (N_27973,N_26600,N_26548);
xor U27974 (N_27974,N_26970,N_26091);
nand U27975 (N_27975,N_26531,N_26106);
xnor U27976 (N_27976,N_25604,N_26017);
nor U27977 (N_27977,N_26540,N_26778);
nor U27978 (N_27978,N_26104,N_26824);
xnor U27979 (N_27979,N_25584,N_25630);
nand U27980 (N_27980,N_25561,N_26371);
and U27981 (N_27981,N_26462,N_25602);
nand U27982 (N_27982,N_25772,N_25715);
nand U27983 (N_27983,N_26139,N_26092);
nor U27984 (N_27984,N_25976,N_26541);
nor U27985 (N_27985,N_26702,N_26671);
nand U27986 (N_27986,N_25759,N_26457);
and U27987 (N_27987,N_26677,N_25722);
nor U27988 (N_27988,N_26860,N_26028);
or U27989 (N_27989,N_26050,N_26380);
nand U27990 (N_27990,N_26113,N_26039);
or U27991 (N_27991,N_26325,N_26109);
nor U27992 (N_27992,N_25504,N_26029);
nand U27993 (N_27993,N_26414,N_25573);
xnor U27994 (N_27994,N_26899,N_25968);
xor U27995 (N_27995,N_25631,N_25654);
nor U27996 (N_27996,N_25771,N_26343);
nor U27997 (N_27997,N_25686,N_25719);
and U27998 (N_27998,N_25821,N_25771);
nor U27999 (N_27999,N_26805,N_26904);
and U28000 (N_28000,N_25604,N_26776);
or U28001 (N_28001,N_26126,N_26280);
nand U28002 (N_28002,N_26841,N_26671);
nand U28003 (N_28003,N_25748,N_26885);
or U28004 (N_28004,N_26628,N_25869);
or U28005 (N_28005,N_26542,N_25857);
xor U28006 (N_28006,N_26058,N_26601);
and U28007 (N_28007,N_26090,N_26437);
and U28008 (N_28008,N_26829,N_26294);
nor U28009 (N_28009,N_26636,N_25655);
xnor U28010 (N_28010,N_26248,N_26326);
nand U28011 (N_28011,N_26261,N_26873);
and U28012 (N_28012,N_26793,N_25834);
or U28013 (N_28013,N_25984,N_25854);
nor U28014 (N_28014,N_25718,N_25886);
or U28015 (N_28015,N_25523,N_25797);
nor U28016 (N_28016,N_26059,N_26576);
nor U28017 (N_28017,N_26316,N_26688);
nor U28018 (N_28018,N_26516,N_26653);
or U28019 (N_28019,N_26624,N_25872);
or U28020 (N_28020,N_26686,N_26953);
nand U28021 (N_28021,N_26002,N_25988);
and U28022 (N_28022,N_26688,N_26919);
xor U28023 (N_28023,N_26317,N_25634);
nor U28024 (N_28024,N_25517,N_25586);
or U28025 (N_28025,N_25816,N_25598);
or U28026 (N_28026,N_25732,N_26349);
xor U28027 (N_28027,N_25757,N_26035);
or U28028 (N_28028,N_26637,N_25508);
xnor U28029 (N_28029,N_26374,N_25974);
and U28030 (N_28030,N_26497,N_26771);
nor U28031 (N_28031,N_26049,N_25794);
nand U28032 (N_28032,N_26363,N_25782);
xor U28033 (N_28033,N_25645,N_26464);
and U28034 (N_28034,N_26770,N_26199);
or U28035 (N_28035,N_26673,N_26153);
nand U28036 (N_28036,N_25910,N_25760);
and U28037 (N_28037,N_26841,N_25704);
xnor U28038 (N_28038,N_25563,N_26422);
nand U28039 (N_28039,N_26004,N_26009);
xor U28040 (N_28040,N_26311,N_25680);
and U28041 (N_28041,N_26479,N_26471);
xor U28042 (N_28042,N_25911,N_26176);
nand U28043 (N_28043,N_26403,N_25927);
xnor U28044 (N_28044,N_26477,N_26776);
and U28045 (N_28045,N_26069,N_26309);
xnor U28046 (N_28046,N_26234,N_26633);
xor U28047 (N_28047,N_26117,N_25710);
nand U28048 (N_28048,N_26807,N_26504);
and U28049 (N_28049,N_25521,N_26258);
xor U28050 (N_28050,N_26442,N_25616);
xor U28051 (N_28051,N_25851,N_26518);
or U28052 (N_28052,N_26325,N_26637);
and U28053 (N_28053,N_25660,N_26527);
xor U28054 (N_28054,N_25644,N_26267);
xor U28055 (N_28055,N_26348,N_25615);
nor U28056 (N_28056,N_26870,N_25701);
and U28057 (N_28057,N_25529,N_25711);
xor U28058 (N_28058,N_26129,N_26026);
nand U28059 (N_28059,N_25787,N_26974);
xor U28060 (N_28060,N_26017,N_26893);
nor U28061 (N_28061,N_26377,N_26029);
nand U28062 (N_28062,N_26698,N_26071);
nor U28063 (N_28063,N_26984,N_26030);
nand U28064 (N_28064,N_26078,N_26946);
or U28065 (N_28065,N_26010,N_25725);
nand U28066 (N_28066,N_25871,N_26832);
and U28067 (N_28067,N_26444,N_25917);
and U28068 (N_28068,N_26630,N_26859);
and U28069 (N_28069,N_25848,N_26347);
nand U28070 (N_28070,N_25778,N_26880);
or U28071 (N_28071,N_25570,N_26003);
nor U28072 (N_28072,N_25721,N_26211);
and U28073 (N_28073,N_26328,N_26447);
xor U28074 (N_28074,N_26195,N_25876);
xnor U28075 (N_28075,N_25674,N_26423);
and U28076 (N_28076,N_25606,N_26258);
or U28077 (N_28077,N_26055,N_25546);
xor U28078 (N_28078,N_25912,N_25503);
xor U28079 (N_28079,N_25863,N_26860);
or U28080 (N_28080,N_26827,N_26012);
nor U28081 (N_28081,N_25729,N_26914);
and U28082 (N_28082,N_25978,N_25526);
nor U28083 (N_28083,N_26751,N_26002);
xnor U28084 (N_28084,N_26006,N_26746);
nand U28085 (N_28085,N_26912,N_25955);
and U28086 (N_28086,N_26137,N_26214);
nor U28087 (N_28087,N_25855,N_26384);
xor U28088 (N_28088,N_26753,N_26590);
nor U28089 (N_28089,N_26770,N_25902);
xor U28090 (N_28090,N_25578,N_26633);
nor U28091 (N_28091,N_26410,N_26076);
nor U28092 (N_28092,N_26634,N_25648);
nand U28093 (N_28093,N_26036,N_25725);
and U28094 (N_28094,N_25702,N_26288);
or U28095 (N_28095,N_25865,N_26925);
and U28096 (N_28096,N_26461,N_26626);
nor U28097 (N_28097,N_25837,N_25948);
and U28098 (N_28098,N_25854,N_26862);
nand U28099 (N_28099,N_26492,N_25536);
xor U28100 (N_28100,N_26741,N_26893);
and U28101 (N_28101,N_26226,N_26849);
xnor U28102 (N_28102,N_26184,N_26235);
nor U28103 (N_28103,N_26479,N_26461);
nand U28104 (N_28104,N_25838,N_25982);
xnor U28105 (N_28105,N_26134,N_26744);
nor U28106 (N_28106,N_26716,N_26036);
or U28107 (N_28107,N_26810,N_25531);
and U28108 (N_28108,N_25502,N_25839);
nor U28109 (N_28109,N_26776,N_25784);
nor U28110 (N_28110,N_26051,N_26815);
or U28111 (N_28111,N_26490,N_26050);
or U28112 (N_28112,N_25999,N_26546);
xnor U28113 (N_28113,N_26476,N_26998);
or U28114 (N_28114,N_26582,N_25511);
and U28115 (N_28115,N_25844,N_26590);
xor U28116 (N_28116,N_26781,N_26636);
nand U28117 (N_28117,N_26070,N_26313);
and U28118 (N_28118,N_26977,N_26270);
nor U28119 (N_28119,N_25633,N_25635);
nor U28120 (N_28120,N_25571,N_26286);
or U28121 (N_28121,N_26078,N_26497);
or U28122 (N_28122,N_26046,N_26101);
or U28123 (N_28123,N_26262,N_26049);
nor U28124 (N_28124,N_26551,N_25607);
and U28125 (N_28125,N_26988,N_26843);
or U28126 (N_28126,N_26414,N_26617);
nand U28127 (N_28127,N_26760,N_26303);
and U28128 (N_28128,N_26239,N_26968);
nor U28129 (N_28129,N_25915,N_26996);
nand U28130 (N_28130,N_25977,N_26847);
nand U28131 (N_28131,N_26228,N_26505);
nand U28132 (N_28132,N_26241,N_25922);
or U28133 (N_28133,N_26468,N_26988);
nand U28134 (N_28134,N_26799,N_25733);
xnor U28135 (N_28135,N_25746,N_26383);
and U28136 (N_28136,N_25963,N_26172);
nand U28137 (N_28137,N_26510,N_25809);
nand U28138 (N_28138,N_25940,N_25511);
nor U28139 (N_28139,N_26234,N_26679);
and U28140 (N_28140,N_25560,N_25734);
nor U28141 (N_28141,N_26002,N_26813);
or U28142 (N_28142,N_26794,N_25741);
or U28143 (N_28143,N_26070,N_25880);
nor U28144 (N_28144,N_26169,N_26050);
or U28145 (N_28145,N_26895,N_25845);
or U28146 (N_28146,N_25553,N_26449);
or U28147 (N_28147,N_26823,N_26701);
and U28148 (N_28148,N_26641,N_25579);
xnor U28149 (N_28149,N_26144,N_25853);
nand U28150 (N_28150,N_25737,N_25735);
or U28151 (N_28151,N_26174,N_26168);
nand U28152 (N_28152,N_26450,N_26539);
nor U28153 (N_28153,N_25506,N_25755);
and U28154 (N_28154,N_26385,N_26819);
xor U28155 (N_28155,N_26845,N_26879);
and U28156 (N_28156,N_26433,N_26605);
xnor U28157 (N_28157,N_25812,N_26046);
nor U28158 (N_28158,N_26749,N_26536);
nand U28159 (N_28159,N_26722,N_26758);
and U28160 (N_28160,N_26469,N_26700);
nor U28161 (N_28161,N_26881,N_25703);
nor U28162 (N_28162,N_25694,N_26662);
and U28163 (N_28163,N_26691,N_26893);
and U28164 (N_28164,N_26678,N_25945);
nor U28165 (N_28165,N_26113,N_26124);
or U28166 (N_28166,N_26867,N_26249);
nand U28167 (N_28167,N_26100,N_26237);
nor U28168 (N_28168,N_25680,N_26755);
nor U28169 (N_28169,N_26240,N_26966);
nor U28170 (N_28170,N_25919,N_26578);
or U28171 (N_28171,N_25587,N_25980);
nor U28172 (N_28172,N_26705,N_25876);
nor U28173 (N_28173,N_26646,N_26285);
or U28174 (N_28174,N_26974,N_26849);
nand U28175 (N_28175,N_25799,N_26457);
or U28176 (N_28176,N_25987,N_26713);
nor U28177 (N_28177,N_26771,N_26943);
or U28178 (N_28178,N_26887,N_25653);
and U28179 (N_28179,N_26377,N_25698);
xnor U28180 (N_28180,N_26457,N_25587);
and U28181 (N_28181,N_25694,N_26949);
nor U28182 (N_28182,N_26711,N_25729);
or U28183 (N_28183,N_26538,N_26143);
nor U28184 (N_28184,N_26396,N_25961);
xnor U28185 (N_28185,N_26960,N_26838);
nand U28186 (N_28186,N_26393,N_26552);
nand U28187 (N_28187,N_25639,N_25687);
nor U28188 (N_28188,N_26069,N_25825);
xor U28189 (N_28189,N_25548,N_26491);
and U28190 (N_28190,N_26703,N_26364);
xor U28191 (N_28191,N_26539,N_26789);
and U28192 (N_28192,N_26095,N_25644);
and U28193 (N_28193,N_26311,N_25770);
and U28194 (N_28194,N_26084,N_26480);
nor U28195 (N_28195,N_25894,N_26531);
and U28196 (N_28196,N_26388,N_26416);
nor U28197 (N_28197,N_26318,N_25672);
nand U28198 (N_28198,N_25597,N_26331);
nand U28199 (N_28199,N_26665,N_26489);
xor U28200 (N_28200,N_26071,N_26533);
or U28201 (N_28201,N_26119,N_26159);
nand U28202 (N_28202,N_26170,N_25790);
nand U28203 (N_28203,N_25699,N_26138);
nand U28204 (N_28204,N_25590,N_25778);
nor U28205 (N_28205,N_26878,N_25934);
nand U28206 (N_28206,N_26582,N_25839);
nand U28207 (N_28207,N_26220,N_26114);
nor U28208 (N_28208,N_26496,N_26987);
nor U28209 (N_28209,N_25598,N_26493);
and U28210 (N_28210,N_26689,N_25715);
and U28211 (N_28211,N_26704,N_26970);
or U28212 (N_28212,N_26117,N_25635);
and U28213 (N_28213,N_26633,N_26869);
nand U28214 (N_28214,N_26251,N_25720);
nand U28215 (N_28215,N_26677,N_26190);
nand U28216 (N_28216,N_25765,N_25507);
or U28217 (N_28217,N_26514,N_25952);
and U28218 (N_28218,N_26807,N_25899);
nand U28219 (N_28219,N_25701,N_25826);
nor U28220 (N_28220,N_26001,N_26109);
and U28221 (N_28221,N_25780,N_26792);
nand U28222 (N_28222,N_26546,N_25572);
and U28223 (N_28223,N_25761,N_26011);
xor U28224 (N_28224,N_26719,N_25768);
and U28225 (N_28225,N_25937,N_26971);
or U28226 (N_28226,N_26678,N_25933);
nor U28227 (N_28227,N_26172,N_26213);
nand U28228 (N_28228,N_26148,N_26597);
nor U28229 (N_28229,N_25733,N_26573);
nor U28230 (N_28230,N_26491,N_25815);
nor U28231 (N_28231,N_25634,N_26512);
xor U28232 (N_28232,N_26958,N_26701);
and U28233 (N_28233,N_26742,N_26185);
xnor U28234 (N_28234,N_26231,N_26473);
nand U28235 (N_28235,N_26885,N_26526);
nor U28236 (N_28236,N_26220,N_25752);
nor U28237 (N_28237,N_26785,N_26089);
xnor U28238 (N_28238,N_25666,N_26081);
nor U28239 (N_28239,N_26444,N_26677);
and U28240 (N_28240,N_26145,N_26030);
xor U28241 (N_28241,N_25897,N_26219);
xnor U28242 (N_28242,N_25601,N_25527);
or U28243 (N_28243,N_26245,N_25716);
nand U28244 (N_28244,N_26794,N_25534);
nor U28245 (N_28245,N_26539,N_25681);
or U28246 (N_28246,N_25876,N_26446);
nand U28247 (N_28247,N_26773,N_25533);
nand U28248 (N_28248,N_26019,N_25868);
xnor U28249 (N_28249,N_26286,N_26538);
nand U28250 (N_28250,N_26294,N_25928);
nand U28251 (N_28251,N_25672,N_26010);
nand U28252 (N_28252,N_26887,N_26855);
and U28253 (N_28253,N_26090,N_26401);
nand U28254 (N_28254,N_26387,N_25525);
nor U28255 (N_28255,N_25634,N_26889);
nand U28256 (N_28256,N_25527,N_25524);
and U28257 (N_28257,N_26410,N_25978);
and U28258 (N_28258,N_26940,N_25886);
and U28259 (N_28259,N_26739,N_26163);
nor U28260 (N_28260,N_26645,N_25864);
and U28261 (N_28261,N_25811,N_26147);
nor U28262 (N_28262,N_26061,N_26125);
nor U28263 (N_28263,N_25533,N_26245);
or U28264 (N_28264,N_26317,N_26131);
nand U28265 (N_28265,N_26970,N_26024);
xor U28266 (N_28266,N_25762,N_26942);
and U28267 (N_28267,N_26283,N_26989);
nor U28268 (N_28268,N_26448,N_25694);
xnor U28269 (N_28269,N_26048,N_26951);
nand U28270 (N_28270,N_26561,N_26316);
or U28271 (N_28271,N_26616,N_26735);
and U28272 (N_28272,N_26302,N_26616);
nor U28273 (N_28273,N_26984,N_25842);
xnor U28274 (N_28274,N_26138,N_26201);
and U28275 (N_28275,N_26212,N_26875);
and U28276 (N_28276,N_25741,N_25760);
and U28277 (N_28277,N_25720,N_26995);
xnor U28278 (N_28278,N_26961,N_26315);
and U28279 (N_28279,N_25805,N_26676);
xnor U28280 (N_28280,N_25804,N_26982);
or U28281 (N_28281,N_25570,N_25532);
nor U28282 (N_28282,N_26956,N_25725);
xnor U28283 (N_28283,N_25936,N_26526);
nor U28284 (N_28284,N_25631,N_26240);
or U28285 (N_28285,N_26863,N_26137);
and U28286 (N_28286,N_26827,N_26775);
nand U28287 (N_28287,N_25664,N_26669);
or U28288 (N_28288,N_25739,N_25849);
xor U28289 (N_28289,N_25884,N_25554);
xnor U28290 (N_28290,N_26466,N_25510);
nand U28291 (N_28291,N_26519,N_25852);
xor U28292 (N_28292,N_26764,N_26375);
nand U28293 (N_28293,N_26656,N_26532);
and U28294 (N_28294,N_26516,N_25732);
nor U28295 (N_28295,N_26983,N_25635);
xnor U28296 (N_28296,N_26490,N_25951);
and U28297 (N_28297,N_26258,N_26528);
nand U28298 (N_28298,N_25898,N_26717);
and U28299 (N_28299,N_26735,N_26283);
nand U28300 (N_28300,N_26217,N_25677);
or U28301 (N_28301,N_26834,N_25686);
xor U28302 (N_28302,N_25541,N_26123);
and U28303 (N_28303,N_25682,N_25941);
and U28304 (N_28304,N_26995,N_26429);
nor U28305 (N_28305,N_25878,N_26338);
and U28306 (N_28306,N_26377,N_26619);
and U28307 (N_28307,N_26583,N_25692);
xor U28308 (N_28308,N_26517,N_26703);
xor U28309 (N_28309,N_26737,N_26105);
nor U28310 (N_28310,N_26036,N_25842);
xnor U28311 (N_28311,N_25541,N_25613);
nor U28312 (N_28312,N_26553,N_26850);
or U28313 (N_28313,N_25702,N_26332);
and U28314 (N_28314,N_26968,N_26522);
or U28315 (N_28315,N_26187,N_26958);
nand U28316 (N_28316,N_26288,N_26038);
and U28317 (N_28317,N_26950,N_26856);
xor U28318 (N_28318,N_26299,N_26244);
nand U28319 (N_28319,N_26840,N_25664);
nand U28320 (N_28320,N_26777,N_26504);
or U28321 (N_28321,N_26732,N_26524);
and U28322 (N_28322,N_26897,N_25898);
xor U28323 (N_28323,N_26324,N_26473);
xor U28324 (N_28324,N_26517,N_26975);
nor U28325 (N_28325,N_26338,N_26460);
nand U28326 (N_28326,N_25505,N_26801);
xnor U28327 (N_28327,N_25744,N_25809);
nand U28328 (N_28328,N_26344,N_25778);
nor U28329 (N_28329,N_26727,N_26583);
nand U28330 (N_28330,N_26490,N_25744);
xnor U28331 (N_28331,N_26866,N_26742);
or U28332 (N_28332,N_25583,N_26394);
nand U28333 (N_28333,N_26335,N_25690);
or U28334 (N_28334,N_26553,N_26109);
nand U28335 (N_28335,N_26682,N_26012);
nand U28336 (N_28336,N_26988,N_26092);
and U28337 (N_28337,N_26756,N_25630);
and U28338 (N_28338,N_25527,N_26953);
or U28339 (N_28339,N_26872,N_26740);
and U28340 (N_28340,N_26843,N_26013);
and U28341 (N_28341,N_26128,N_26562);
nand U28342 (N_28342,N_26278,N_25725);
and U28343 (N_28343,N_26880,N_26203);
xor U28344 (N_28344,N_25536,N_26577);
and U28345 (N_28345,N_26560,N_25852);
xor U28346 (N_28346,N_25540,N_26458);
nand U28347 (N_28347,N_26149,N_26303);
nor U28348 (N_28348,N_25524,N_25553);
nor U28349 (N_28349,N_26142,N_25755);
xnor U28350 (N_28350,N_26000,N_26932);
or U28351 (N_28351,N_25761,N_26786);
nand U28352 (N_28352,N_25786,N_26808);
nor U28353 (N_28353,N_25647,N_26910);
or U28354 (N_28354,N_25535,N_25702);
nand U28355 (N_28355,N_26339,N_25526);
xor U28356 (N_28356,N_25675,N_26258);
or U28357 (N_28357,N_25503,N_26987);
nand U28358 (N_28358,N_25701,N_26249);
xnor U28359 (N_28359,N_26139,N_26136);
xnor U28360 (N_28360,N_26295,N_25788);
and U28361 (N_28361,N_26235,N_26025);
or U28362 (N_28362,N_26651,N_26560);
and U28363 (N_28363,N_26125,N_25668);
nand U28364 (N_28364,N_25783,N_25834);
xnor U28365 (N_28365,N_26553,N_26832);
nor U28366 (N_28366,N_25565,N_26941);
nand U28367 (N_28367,N_26566,N_26554);
and U28368 (N_28368,N_25712,N_25598);
nor U28369 (N_28369,N_25534,N_25942);
nand U28370 (N_28370,N_25501,N_26768);
xor U28371 (N_28371,N_25908,N_26354);
and U28372 (N_28372,N_25918,N_26794);
xnor U28373 (N_28373,N_26583,N_26537);
nor U28374 (N_28374,N_26038,N_26504);
nor U28375 (N_28375,N_26205,N_26991);
nand U28376 (N_28376,N_26180,N_26391);
nand U28377 (N_28377,N_26162,N_26924);
nor U28378 (N_28378,N_26380,N_25584);
nor U28379 (N_28379,N_26906,N_26048);
and U28380 (N_28380,N_26474,N_26918);
nand U28381 (N_28381,N_26849,N_25834);
or U28382 (N_28382,N_26029,N_25657);
nor U28383 (N_28383,N_25898,N_25878);
nor U28384 (N_28384,N_25673,N_26967);
nand U28385 (N_28385,N_26029,N_25753);
xor U28386 (N_28386,N_25871,N_26300);
and U28387 (N_28387,N_25643,N_25564);
or U28388 (N_28388,N_26793,N_26976);
and U28389 (N_28389,N_25723,N_26873);
xor U28390 (N_28390,N_26036,N_26536);
nand U28391 (N_28391,N_26076,N_26879);
xor U28392 (N_28392,N_26261,N_26103);
and U28393 (N_28393,N_25549,N_26120);
nor U28394 (N_28394,N_25801,N_25939);
nand U28395 (N_28395,N_26777,N_26469);
or U28396 (N_28396,N_25894,N_25716);
and U28397 (N_28397,N_26109,N_25661);
and U28398 (N_28398,N_26058,N_26443);
xnor U28399 (N_28399,N_26165,N_25901);
nand U28400 (N_28400,N_25590,N_25845);
xnor U28401 (N_28401,N_26700,N_26300);
or U28402 (N_28402,N_26429,N_26708);
and U28403 (N_28403,N_26862,N_26480);
xor U28404 (N_28404,N_25685,N_25553);
and U28405 (N_28405,N_26786,N_26644);
or U28406 (N_28406,N_26295,N_26664);
nor U28407 (N_28407,N_26065,N_25809);
xor U28408 (N_28408,N_26147,N_25580);
nor U28409 (N_28409,N_25647,N_25659);
nor U28410 (N_28410,N_26483,N_26004);
nor U28411 (N_28411,N_26431,N_26430);
xnor U28412 (N_28412,N_26164,N_25850);
or U28413 (N_28413,N_26275,N_25622);
or U28414 (N_28414,N_26827,N_26761);
or U28415 (N_28415,N_25595,N_26306);
xnor U28416 (N_28416,N_26565,N_26841);
nand U28417 (N_28417,N_26251,N_26175);
nor U28418 (N_28418,N_25802,N_26816);
nand U28419 (N_28419,N_25563,N_26406);
and U28420 (N_28420,N_26553,N_26660);
nor U28421 (N_28421,N_26052,N_26905);
and U28422 (N_28422,N_26923,N_25889);
nor U28423 (N_28423,N_25510,N_25797);
or U28424 (N_28424,N_26690,N_25966);
xor U28425 (N_28425,N_26640,N_26983);
xor U28426 (N_28426,N_25618,N_26053);
and U28427 (N_28427,N_25867,N_25677);
xor U28428 (N_28428,N_26601,N_26344);
xor U28429 (N_28429,N_26177,N_26066);
xor U28430 (N_28430,N_26819,N_25767);
nand U28431 (N_28431,N_26341,N_25555);
nand U28432 (N_28432,N_26497,N_25854);
nor U28433 (N_28433,N_26978,N_26291);
nand U28434 (N_28434,N_25816,N_26351);
or U28435 (N_28435,N_26815,N_26785);
or U28436 (N_28436,N_25841,N_26822);
nand U28437 (N_28437,N_25783,N_25741);
nand U28438 (N_28438,N_26928,N_26554);
nor U28439 (N_28439,N_26756,N_25886);
and U28440 (N_28440,N_25525,N_26506);
and U28441 (N_28441,N_26641,N_26704);
and U28442 (N_28442,N_25794,N_26985);
nor U28443 (N_28443,N_26546,N_25721);
nand U28444 (N_28444,N_26618,N_26409);
or U28445 (N_28445,N_26432,N_25882);
nor U28446 (N_28446,N_25838,N_25763);
nor U28447 (N_28447,N_26694,N_25926);
xor U28448 (N_28448,N_25692,N_26051);
and U28449 (N_28449,N_26594,N_26549);
nand U28450 (N_28450,N_25646,N_26007);
or U28451 (N_28451,N_25799,N_25795);
xnor U28452 (N_28452,N_25825,N_26003);
nand U28453 (N_28453,N_26982,N_25734);
and U28454 (N_28454,N_26224,N_26487);
nor U28455 (N_28455,N_25795,N_26971);
and U28456 (N_28456,N_26817,N_25969);
or U28457 (N_28457,N_26179,N_26750);
xor U28458 (N_28458,N_26849,N_25761);
nor U28459 (N_28459,N_25506,N_26436);
xor U28460 (N_28460,N_26327,N_25985);
or U28461 (N_28461,N_26337,N_26396);
or U28462 (N_28462,N_26765,N_26867);
nand U28463 (N_28463,N_25990,N_26561);
or U28464 (N_28464,N_26716,N_25730);
xor U28465 (N_28465,N_25839,N_26390);
nand U28466 (N_28466,N_25885,N_26140);
or U28467 (N_28467,N_25896,N_25871);
xor U28468 (N_28468,N_26708,N_26407);
xor U28469 (N_28469,N_25813,N_26593);
nand U28470 (N_28470,N_25775,N_25668);
xor U28471 (N_28471,N_25504,N_25615);
nor U28472 (N_28472,N_25507,N_25795);
and U28473 (N_28473,N_26586,N_25820);
xor U28474 (N_28474,N_26075,N_25721);
or U28475 (N_28475,N_26977,N_26140);
xor U28476 (N_28476,N_26480,N_26546);
and U28477 (N_28477,N_25769,N_26993);
nor U28478 (N_28478,N_25538,N_26064);
or U28479 (N_28479,N_25701,N_26735);
nor U28480 (N_28480,N_26991,N_26022);
xnor U28481 (N_28481,N_26393,N_26602);
or U28482 (N_28482,N_25873,N_26428);
or U28483 (N_28483,N_25677,N_26553);
nand U28484 (N_28484,N_26318,N_25981);
nand U28485 (N_28485,N_25785,N_25673);
nor U28486 (N_28486,N_25795,N_25541);
or U28487 (N_28487,N_26312,N_26039);
or U28488 (N_28488,N_26532,N_26049);
xor U28489 (N_28489,N_25874,N_26207);
and U28490 (N_28490,N_26625,N_25871);
xnor U28491 (N_28491,N_26131,N_26380);
nor U28492 (N_28492,N_26261,N_25760);
and U28493 (N_28493,N_26747,N_26294);
xnor U28494 (N_28494,N_26601,N_26283);
nor U28495 (N_28495,N_26269,N_26998);
nor U28496 (N_28496,N_25784,N_26244);
or U28497 (N_28497,N_25608,N_25798);
or U28498 (N_28498,N_26295,N_25958);
or U28499 (N_28499,N_26734,N_25512);
or U28500 (N_28500,N_28048,N_28112);
or U28501 (N_28501,N_27903,N_28305);
and U28502 (N_28502,N_28252,N_27129);
xnor U28503 (N_28503,N_28096,N_27353);
or U28504 (N_28504,N_27762,N_27100);
xnor U28505 (N_28505,N_27653,N_27260);
xnor U28506 (N_28506,N_27450,N_28433);
and U28507 (N_28507,N_28205,N_28211);
or U28508 (N_28508,N_27757,N_27689);
or U28509 (N_28509,N_28282,N_27969);
or U28510 (N_28510,N_27044,N_28337);
xor U28511 (N_28511,N_27121,N_28271);
nand U28512 (N_28512,N_27791,N_27527);
and U28513 (N_28513,N_27273,N_27247);
xor U28514 (N_28514,N_27118,N_27367);
or U28515 (N_28515,N_27289,N_27190);
nor U28516 (N_28516,N_27440,N_28051);
or U28517 (N_28517,N_27461,N_27640);
nor U28518 (N_28518,N_27394,N_27886);
xnor U28519 (N_28519,N_28458,N_27449);
xor U28520 (N_28520,N_27560,N_27950);
nor U28521 (N_28521,N_27403,N_27995);
or U28522 (N_28522,N_28239,N_27153);
nor U28523 (N_28523,N_27170,N_27525);
and U28524 (N_28524,N_27931,N_28276);
or U28525 (N_28525,N_28439,N_28130);
and U28526 (N_28526,N_28092,N_28166);
xor U28527 (N_28527,N_27125,N_27441);
nand U28528 (N_28528,N_28331,N_27743);
xnor U28529 (N_28529,N_27774,N_27145);
and U28530 (N_28530,N_28097,N_27591);
nand U28531 (N_28531,N_27398,N_27928);
nand U28532 (N_28532,N_27466,N_27977);
nor U28533 (N_28533,N_28015,N_28493);
xnor U28534 (N_28534,N_28333,N_27671);
or U28535 (N_28535,N_27794,N_27956);
nor U28536 (N_28536,N_27152,N_28309);
xor U28537 (N_28537,N_27454,N_27068);
or U28538 (N_28538,N_27952,N_27694);
nand U28539 (N_28539,N_27104,N_27401);
xnor U28540 (N_28540,N_27963,N_28348);
nor U28541 (N_28541,N_27855,N_28310);
nor U28542 (N_28542,N_27438,N_28014);
nor U28543 (N_28543,N_27237,N_27057);
xor U28544 (N_28544,N_27526,N_27053);
and U28545 (N_28545,N_27204,N_27040);
nand U28546 (N_28546,N_28312,N_28264);
nor U28547 (N_28547,N_27410,N_27369);
or U28548 (N_28548,N_27140,N_27951);
nand U28549 (N_28549,N_28420,N_28406);
nor U28550 (N_28550,N_27524,N_28298);
and U28551 (N_28551,N_27662,N_27832);
nor U28552 (N_28552,N_27187,N_28029);
or U28553 (N_28553,N_27587,N_28040);
nor U28554 (N_28554,N_28449,N_28063);
nand U28555 (N_28555,N_27900,N_27275);
and U28556 (N_28556,N_27734,N_27637);
nand U28557 (N_28557,N_28463,N_27512);
and U28558 (N_28558,N_27491,N_27944);
nor U28559 (N_28559,N_28190,N_27478);
or U28560 (N_28560,N_27060,N_27785);
xor U28561 (N_28561,N_28451,N_27829);
xor U28562 (N_28562,N_27552,N_27983);
and U28563 (N_28563,N_27910,N_27284);
or U28564 (N_28564,N_27282,N_28056);
xnor U28565 (N_28565,N_27154,N_27501);
nor U28566 (N_28566,N_28383,N_27274);
xor U28567 (N_28567,N_28297,N_28440);
xnor U28568 (N_28568,N_27162,N_28293);
or U28569 (N_28569,N_27516,N_28146);
nand U28570 (N_28570,N_27146,N_27965);
or U28571 (N_28571,N_28000,N_27231);
nor U28572 (N_28572,N_27534,N_27608);
nor U28573 (N_28573,N_27864,N_27610);
nand U28574 (N_28574,N_27058,N_27473);
or U28575 (N_28575,N_28280,N_28486);
xnor U28576 (N_28576,N_27661,N_28374);
xor U28577 (N_28577,N_28295,N_27705);
or U28578 (N_28578,N_28428,N_27036);
or U28579 (N_28579,N_27188,N_27225);
and U28580 (N_28580,N_27913,N_27739);
or U28581 (N_28581,N_28425,N_28483);
nor U28582 (N_28582,N_27319,N_27167);
and U28583 (N_28583,N_28165,N_27322);
and U28584 (N_28584,N_27506,N_27737);
nor U28585 (N_28585,N_28140,N_28075);
nand U28586 (N_28586,N_27061,N_27250);
or U28587 (N_28587,N_27309,N_27173);
nor U28588 (N_28588,N_27198,N_27137);
nand U28589 (N_28589,N_27380,N_27652);
nor U28590 (N_28590,N_28119,N_27748);
or U28591 (N_28591,N_27769,N_27655);
nand U28592 (N_28592,N_27132,N_27136);
xnor U28593 (N_28593,N_28316,N_27625);
xnor U28594 (N_28594,N_27088,N_27984);
nor U28595 (N_28595,N_27479,N_27559);
nor U28596 (N_28596,N_27596,N_27782);
and U28597 (N_28597,N_27665,N_27642);
and U28598 (N_28598,N_27475,N_28371);
or U28599 (N_28599,N_27281,N_27432);
xnor U28600 (N_28600,N_27317,N_27311);
and U28601 (N_28601,N_27901,N_27701);
and U28602 (N_28602,N_27815,N_27487);
or U28603 (N_28603,N_27005,N_27863);
or U28604 (N_28604,N_28169,N_28033);
or U28605 (N_28605,N_28424,N_27464);
nor U28606 (N_28606,N_27488,N_28187);
nand U28607 (N_28607,N_28210,N_28030);
or U28608 (N_28608,N_28055,N_28226);
or U28609 (N_28609,N_27699,N_27019);
xnor U28610 (N_28610,N_27672,N_27481);
nand U28611 (N_28611,N_28275,N_27667);
nor U28612 (N_28612,N_27406,N_28490);
nand U28613 (N_28613,N_27008,N_28444);
and U28614 (N_28614,N_28317,N_27878);
nand U28615 (N_28615,N_27643,N_28034);
nor U28616 (N_28616,N_28343,N_28151);
xnor U28617 (N_28617,N_28476,N_27590);
nand U28618 (N_28618,N_28421,N_27230);
xor U28619 (N_28619,N_27426,N_27912);
and U28620 (N_28620,N_27312,N_28291);
or U28621 (N_28621,N_28286,N_27375);
nor U28622 (N_28622,N_28209,N_27666);
and U28623 (N_28623,N_28162,N_28240);
nand U28624 (N_28624,N_28397,N_27497);
nand U28625 (N_28625,N_27024,N_28437);
and U28626 (N_28626,N_27593,N_28141);
xor U28627 (N_28627,N_27766,N_27092);
and U28628 (N_28628,N_27072,N_28113);
nor U28629 (N_28629,N_27917,N_28289);
nor U28630 (N_28630,N_27081,N_28403);
or U28631 (N_28631,N_28179,N_27205);
or U28632 (N_28632,N_28136,N_28017);
or U28633 (N_28633,N_27255,N_27817);
nor U28634 (N_28634,N_27680,N_27644);
nor U28635 (N_28635,N_28147,N_28060);
nand U28636 (N_28636,N_27601,N_27707);
xnor U28637 (N_28637,N_27096,N_27548);
nor U28638 (N_28638,N_27651,N_27164);
xnor U28639 (N_28639,N_28314,N_27871);
and U28640 (N_28640,N_27206,N_28218);
nor U28641 (N_28641,N_27854,N_27895);
and U28642 (N_28642,N_27876,N_27254);
xnor U28643 (N_28643,N_28470,N_27731);
xor U28644 (N_28644,N_27872,N_27783);
xor U28645 (N_28645,N_28242,N_28247);
nor U28646 (N_28646,N_28329,N_28392);
xnor U28647 (N_28647,N_27557,N_27444);
nand U28648 (N_28648,N_27304,N_28159);
xnor U28649 (N_28649,N_27366,N_28244);
nand U28650 (N_28650,N_27489,N_27947);
and U28651 (N_28651,N_28079,N_27704);
nor U28652 (N_28652,N_27507,N_27603);
and U28653 (N_28653,N_27021,N_28487);
or U28654 (N_28654,N_27839,N_28038);
and U28655 (N_28655,N_27893,N_27733);
and U28656 (N_28656,N_27915,N_28241);
nand U28657 (N_28657,N_27113,N_27341);
nor U28658 (N_28658,N_27948,N_27509);
xnor U28659 (N_28659,N_27678,N_27307);
nor U28660 (N_28660,N_27267,N_28234);
and U28661 (N_28661,N_28059,N_27503);
or U28662 (N_28662,N_28465,N_28137);
xnor U28663 (N_28663,N_27883,N_27080);
nor U28664 (N_28664,N_28477,N_28229);
xnor U28665 (N_28665,N_28398,N_28422);
nor U28666 (N_28666,N_27709,N_28198);
and U28667 (N_28667,N_28028,N_27576);
nand U28668 (N_28668,N_27580,N_27921);
or U28669 (N_28669,N_27090,N_27636);
and U28670 (N_28670,N_27226,N_27124);
or U28671 (N_28671,N_27752,N_28116);
or U28672 (N_28672,N_27806,N_28388);
and U28673 (N_28673,N_28180,N_27758);
nor U28674 (N_28674,N_28126,N_27802);
xnor U28675 (N_28675,N_27433,N_27750);
nor U28676 (N_28676,N_27134,N_27435);
and U28677 (N_28677,N_28288,N_27617);
and U28678 (N_28678,N_27793,N_27979);
nand U28679 (N_28679,N_27741,N_27037);
nand U28680 (N_28680,N_27898,N_28199);
or U28681 (N_28681,N_27305,N_28156);
xor U28682 (N_28682,N_27561,N_27025);
and U28683 (N_28683,N_27386,N_27690);
nor U28684 (N_28684,N_28031,N_28294);
nor U28685 (N_28685,N_27214,N_27291);
nand U28686 (N_28686,N_27868,N_27174);
nor U28687 (N_28687,N_27097,N_27055);
and U28688 (N_28688,N_27959,N_28255);
and U28689 (N_28689,N_27911,N_28098);
nand U28690 (N_28690,N_28114,N_28266);
nand U28691 (N_28691,N_28182,N_28157);
xnor U28692 (N_28692,N_28010,N_28380);
and U28693 (N_28693,N_28323,N_28292);
nand U28694 (N_28694,N_28110,N_28217);
nor U28695 (N_28695,N_28172,N_27418);
and U28696 (N_28696,N_27339,N_28389);
or U28697 (N_28697,N_27451,N_27391);
nand U28698 (N_28698,N_27390,N_28132);
xor U28699 (N_28699,N_27896,N_27112);
xnor U28700 (N_28700,N_27881,N_28232);
nor U28701 (N_28701,N_27382,N_28274);
nor U28702 (N_28702,N_28448,N_27028);
nor U28703 (N_28703,N_27084,N_28251);
or U28704 (N_28704,N_28300,N_27935);
and U28705 (N_28705,N_27606,N_28134);
or U28706 (N_28706,N_27659,N_27941);
nand U28707 (N_28707,N_28479,N_28386);
nor U28708 (N_28708,N_27370,N_27141);
and U28709 (N_28709,N_28365,N_27348);
and U28710 (N_28710,N_27955,N_28296);
or U28711 (N_28711,N_27813,N_27934);
nand U28712 (N_28712,N_27455,N_27494);
or U28713 (N_28713,N_27909,N_27326);
nand U28714 (N_28714,N_27976,N_28003);
xor U28715 (N_28715,N_28046,N_28066);
xor U28716 (N_28716,N_28492,N_28131);
nand U28717 (N_28717,N_28102,N_28044);
nor U28718 (N_28718,N_27120,N_27978);
and U28719 (N_28719,N_27065,N_27003);
nor U28720 (N_28720,N_27975,N_27195);
and U28721 (N_28721,N_27685,N_27962);
or U28722 (N_28722,N_28468,N_28262);
xnor U28723 (N_28723,N_27632,N_27834);
or U28724 (N_28724,N_28069,N_27875);
and U28725 (N_28725,N_27123,N_27259);
nor U28726 (N_28726,N_28122,N_27344);
nand U28727 (N_28727,N_27788,N_27323);
nand U28728 (N_28728,N_27849,N_27980);
nor U28729 (N_28729,N_27692,N_28359);
nand U28730 (N_28730,N_28175,N_28236);
xor U28731 (N_28731,N_28108,N_28089);
or U28732 (N_28732,N_28260,N_27483);
and U28733 (N_28733,N_28285,N_27712);
and U28734 (N_28734,N_27989,N_27463);
nand U28735 (N_28735,N_28019,N_27159);
nor U28736 (N_28736,N_28171,N_28128);
nor U28737 (N_28737,N_28372,N_27658);
xor U28738 (N_28738,N_28133,N_27413);
nor U28739 (N_28739,N_27777,N_27837);
and U28740 (N_28740,N_27556,N_28407);
and U28741 (N_28741,N_27936,N_27575);
nor U28742 (N_28742,N_27789,N_27083);
or U28743 (N_28743,N_27365,N_27320);
xor U28744 (N_28744,N_28436,N_27098);
and U28745 (N_28745,N_27283,N_27286);
nand U28746 (N_28746,N_28191,N_27537);
xnor U28747 (N_28747,N_27315,N_27392);
nand U28748 (N_28748,N_28400,N_27867);
or U28749 (N_28749,N_28026,N_27328);
nand U28750 (N_28750,N_28022,N_28370);
or U28751 (N_28751,N_28154,N_27540);
nand U28752 (N_28752,N_27358,N_28036);
xor U28753 (N_28753,N_27990,N_27157);
xnor U28754 (N_28754,N_28461,N_27363);
or U28755 (N_28755,N_27039,N_27998);
or U28756 (N_28756,N_27856,N_28450);
xor U28757 (N_28757,N_27780,N_27285);
nand U28758 (N_28758,N_27352,N_28339);
nor U28759 (N_28759,N_28201,N_27108);
nand U28760 (N_28760,N_27045,N_27711);
and U28761 (N_28761,N_28409,N_28423);
nand U28762 (N_28762,N_28054,N_27754);
xnor U28763 (N_28763,N_27949,N_27439);
nor U28764 (N_28764,N_27811,N_27696);
nor U28765 (N_28765,N_28287,N_27840);
nor U28766 (N_28766,N_28302,N_27325);
nor U28767 (N_28767,N_27297,N_27932);
nor U28768 (N_28768,N_27776,N_27073);
or U28769 (N_28769,N_27833,N_28249);
nand U28770 (N_28770,N_28391,N_27589);
and U28771 (N_28771,N_28195,N_27654);
nand U28772 (N_28772,N_28043,N_28427);
or U28773 (N_28773,N_28341,N_28336);
or U28774 (N_28774,N_28369,N_27810);
xnor U28775 (N_28775,N_27614,N_27062);
and U28776 (N_28776,N_28250,N_28368);
nand U28777 (N_28777,N_27482,N_27574);
xor U28778 (N_28778,N_27182,N_27351);
nand U28779 (N_28779,N_27670,N_27818);
or U28780 (N_28780,N_27107,N_28441);
nor U28781 (N_28781,N_28315,N_27215);
or U28782 (N_28782,N_27469,N_28163);
nor U28783 (N_28783,N_28213,N_27229);
and U28784 (N_28784,N_28219,N_27533);
or U28785 (N_28785,N_28005,N_28037);
or U28786 (N_28786,N_27906,N_27517);
or U28787 (N_28787,N_27841,N_28068);
nor U28788 (N_28788,N_28485,N_28259);
and U28789 (N_28789,N_27476,N_27747);
xnor U28790 (N_28790,N_28321,N_28207);
nor U28791 (N_28791,N_28177,N_27316);
and U28792 (N_28792,N_28167,N_27877);
and U28793 (N_28793,N_27773,N_27046);
xor U28794 (N_28794,N_27076,N_27355);
or U28795 (N_28795,N_27436,N_27029);
xnor U28796 (N_28796,N_28047,N_27566);
and U28797 (N_28797,N_28404,N_27798);
nand U28798 (N_28798,N_27604,N_28138);
nand U28799 (N_28799,N_27649,N_28494);
or U28800 (N_28800,N_28174,N_27368);
nand U28801 (N_28801,N_27814,N_27117);
or U28802 (N_28802,N_27228,N_28283);
nor U28803 (N_28803,N_27718,N_28460);
or U28804 (N_28804,N_27781,N_27514);
nor U28805 (N_28805,N_27437,N_28127);
nor U28806 (N_28806,N_27716,N_27295);
and U28807 (N_28807,N_27656,N_28462);
xor U28808 (N_28808,N_28018,N_28100);
nor U28809 (N_28809,N_27966,N_27786);
or U28810 (N_28810,N_27714,N_27579);
and U28811 (N_28811,N_27735,N_28384);
or U28812 (N_28812,N_28189,N_27000);
and U28813 (N_28813,N_27795,N_27732);
and U28814 (N_28814,N_27144,N_27677);
xor U28815 (N_28815,N_27621,N_27349);
xor U28816 (N_28816,N_27627,N_28117);
and U28817 (N_28817,N_27521,N_28123);
nand U28818 (N_28818,N_27568,N_27477);
or U28819 (N_28819,N_27513,N_27333);
or U28820 (N_28820,N_27238,N_27940);
nand U28821 (N_28821,N_28105,N_27245);
xnor U28822 (N_28822,N_27462,N_27262);
nor U28823 (N_28823,N_27865,N_27414);
or U28824 (N_28824,N_27499,N_27650);
xnor U28825 (N_28825,N_27991,N_27329);
nand U28826 (N_28826,N_27495,N_27850);
xor U28827 (N_28827,N_27973,N_27095);
and U28828 (N_28828,N_27727,N_27530);
nand U28829 (N_28829,N_27122,N_27300);
nand U28830 (N_28830,N_27581,N_27419);
or U28831 (N_28831,N_28340,N_27862);
or U28832 (N_28832,N_27924,N_27302);
or U28833 (N_28833,N_27397,N_27018);
xnor U28834 (N_28834,N_27143,N_28115);
or U28835 (N_28835,N_27184,N_28202);
nor U28836 (N_28836,N_27324,N_27171);
xnor U28837 (N_28837,N_28322,N_27888);
and U28838 (N_28838,N_28385,N_27359);
and U28839 (N_28839,N_27086,N_27584);
and U28840 (N_28840,N_28222,N_28027);
nand U28841 (N_28841,N_28489,N_27056);
or U28842 (N_28842,N_27256,N_27142);
nor U28843 (N_28843,N_28058,N_27429);
xnor U28844 (N_28844,N_27101,N_28067);
or U28845 (N_28845,N_28469,N_27772);
nand U28846 (N_28846,N_27937,N_28290);
xnor U28847 (N_28847,N_28072,N_27816);
and U28848 (N_28848,N_28254,N_28184);
xnor U28849 (N_28849,N_27961,N_27918);
xor U28850 (N_28850,N_27387,N_27356);
nor U28851 (N_28851,N_27942,N_28246);
nand U28852 (N_28852,N_28367,N_27916);
xnor U28853 (N_28853,N_27720,N_27586);
nor U28854 (N_28854,N_27180,N_27052);
and U28855 (N_28855,N_27823,N_28170);
nor U28856 (N_28856,N_28438,N_27460);
nand U28857 (N_28857,N_27892,N_27729);
nand U28858 (N_28858,N_28065,N_27957);
nor U28859 (N_28859,N_27303,N_28495);
or U28860 (N_28860,N_27964,N_28429);
nand U28861 (N_28861,N_27595,N_27089);
and U28862 (N_28862,N_27031,N_27510);
nand U28863 (N_28863,N_27110,N_27508);
xor U28864 (N_28864,N_28042,N_27549);
xor U28865 (N_28865,N_28349,N_27175);
xor U28866 (N_28866,N_27266,N_27213);
or U28867 (N_28867,N_27828,N_28362);
or U28868 (N_28868,N_28445,N_28381);
xnor U28869 (N_28869,N_28197,N_27087);
nand U28870 (N_28870,N_27257,N_28376);
nand U28871 (N_28871,N_28273,N_27759);
nand U28872 (N_28872,N_27801,N_28363);
xor U28873 (N_28873,N_27193,N_28311);
or U28874 (N_28874,N_27336,N_27023);
nand U28875 (N_28875,N_27445,N_27074);
nand U28876 (N_28876,N_28328,N_28330);
and U28877 (N_28877,N_27075,N_28334);
or U28878 (N_28878,N_27562,N_28164);
or U28879 (N_28879,N_27456,N_28093);
nor U28880 (N_28880,N_28077,N_27428);
or U28881 (N_28881,N_27538,N_27035);
nor U28882 (N_28882,N_27771,N_27105);
and U28883 (N_28883,N_28107,N_27264);
or U28884 (N_28884,N_28272,N_28415);
or U28885 (N_28885,N_27417,N_27411);
nand U28886 (N_28886,N_28011,N_27176);
xor U28887 (N_28887,N_27033,N_27668);
or U28888 (N_28888,N_27623,N_27400);
and U28889 (N_28889,N_27519,N_27156);
xnor U28890 (N_28890,N_27845,N_27384);
nand U28891 (N_28891,N_27372,N_28347);
and U28892 (N_28892,N_27093,N_27130);
nand U28893 (N_28893,N_27778,N_28039);
or U28894 (N_28894,N_28150,N_27611);
nor U28895 (N_28895,N_27700,N_27395);
and U28896 (N_28896,N_27314,N_28121);
xnor U28897 (N_28897,N_28106,N_27020);
nor U28898 (N_28898,N_27027,N_28326);
or U28899 (N_28899,N_28045,N_28263);
xnor U28900 (N_28900,N_28431,N_27605);
and U28901 (N_28901,N_27049,N_27004);
nor U28902 (N_28902,N_27127,N_28214);
xor U28903 (N_28903,N_28355,N_27091);
nand U28904 (N_28904,N_27465,N_27629);
nor U28905 (N_28905,N_27313,N_27337);
xor U28906 (N_28906,N_27338,N_27012);
and U28907 (N_28907,N_27181,N_27493);
nand U28908 (N_28908,N_27128,N_28480);
nand U28909 (N_28909,N_28012,N_28084);
and U28910 (N_28910,N_27034,N_27927);
xnor U28911 (N_28911,N_27981,N_27899);
nand U28912 (N_28912,N_27242,N_27362);
or U28913 (N_28913,N_27796,N_27111);
or U28914 (N_28914,N_28307,N_27343);
or U28915 (N_28915,N_27770,N_27588);
xnor U28916 (N_28916,N_27929,N_27999);
nand U28917 (N_28917,N_27119,N_28256);
xnor U28918 (N_28918,N_27103,N_28426);
xnor U28919 (N_28919,N_27288,N_27660);
and U28920 (N_28920,N_28332,N_27066);
xor U28921 (N_28921,N_27787,N_28281);
xnor U28922 (N_28922,N_27330,N_27115);
nor U28923 (N_28923,N_27669,N_28443);
and U28924 (N_28924,N_27224,N_28008);
nand U28925 (N_28925,N_28418,N_27933);
or U28926 (N_28926,N_28491,N_28088);
or U28927 (N_28927,N_27749,N_28153);
xnor U28928 (N_28928,N_27236,N_27613);
xor U28929 (N_28929,N_27189,N_28109);
nand U28930 (N_28930,N_27011,N_27663);
xnor U28931 (N_28931,N_27631,N_28020);
or U28932 (N_28932,N_27048,N_27249);
or U28933 (N_28933,N_27270,N_27523);
or U28934 (N_28934,N_27471,N_27407);
and U28935 (N_28935,N_27434,N_27197);
or U28936 (N_28936,N_28204,N_27563);
or U28937 (N_28937,N_27708,N_27717);
and U28938 (N_28938,N_27378,N_28373);
nor U28939 (N_28939,N_27821,N_27582);
or U28940 (N_28940,N_27502,N_27290);
nor U28941 (N_28941,N_28181,N_27930);
or U28942 (N_28942,N_27972,N_27554);
xor U28943 (N_28943,N_28073,N_27939);
xnor U28944 (N_28944,N_28454,N_28432);
nor U28945 (N_28945,N_28399,N_27904);
xnor U28946 (N_28946,N_27607,N_27001);
nand U28947 (N_28947,N_27222,N_27425);
nor U28948 (N_28948,N_27292,N_27172);
nand U28949 (N_28949,N_27470,N_27819);
nor U28950 (N_28950,N_27071,N_28095);
nor U28951 (N_28951,N_27880,N_27693);
or U28952 (N_28952,N_27234,N_27109);
xnor U28953 (N_28953,N_27698,N_27015);
xor U28954 (N_28954,N_27296,N_27721);
xor U28955 (N_28955,N_27616,N_27169);
or U28956 (N_28956,N_27064,N_28346);
nand U28957 (N_28957,N_28375,N_27272);
or U28958 (N_28958,N_27728,N_27017);
nand U28959 (N_28959,N_27293,N_27006);
xnor U28960 (N_28960,N_27997,N_27306);
and U28961 (N_28961,N_27836,N_27177);
xnor U28962 (N_28962,N_27278,N_27340);
xor U28963 (N_28963,N_27106,N_28344);
or U28964 (N_28964,N_28243,N_28324);
nor U28965 (N_28965,N_27207,N_27452);
nand U28966 (N_28966,N_27412,N_27622);
nand U28967 (N_28967,N_27925,N_28083);
nor U28968 (N_28968,N_27539,N_28475);
or U28969 (N_28969,N_28090,N_27953);
xor U28970 (N_28970,N_27615,N_28230);
and U28971 (N_28971,N_27824,N_27800);
or U28972 (N_28972,N_27646,N_27252);
and U28973 (N_28973,N_27674,N_28253);
or U28974 (N_28974,N_27371,N_27457);
nand U28975 (N_28975,N_27740,N_27321);
nand U28976 (N_28976,N_27504,N_27423);
nor U28977 (N_28977,N_27847,N_28208);
xnor U28978 (N_28978,N_27612,N_27396);
xor U28979 (N_28979,N_28456,N_27009);
nand U28980 (N_28980,N_27299,N_28087);
nor U28981 (N_28981,N_27446,N_27681);
or U28982 (N_28982,N_27389,N_27243);
or U28983 (N_28983,N_28455,N_27047);
or U28984 (N_28984,N_27767,N_28142);
xor U28985 (N_28985,N_27738,N_27448);
xor U28986 (N_28986,N_28396,N_27138);
or U28987 (N_28987,N_27746,N_27726);
nor U28988 (N_28988,N_27719,N_27258);
xnor U28989 (N_28989,N_27094,N_27196);
nor U28990 (N_28990,N_27069,N_28158);
and U28991 (N_28991,N_28016,N_28358);
and U28992 (N_28992,N_28284,N_27848);
nand U28993 (N_28993,N_27235,N_27424);
and U28994 (N_28994,N_27203,N_28278);
or U28995 (N_28995,N_28301,N_27161);
xor U28996 (N_28996,N_27459,N_27553);
and U28997 (N_28997,N_27542,N_27240);
nand U28998 (N_28998,N_27807,N_27223);
nor U28999 (N_28999,N_27342,N_27042);
or U29000 (N_29000,N_27051,N_27280);
or U29001 (N_29001,N_27715,N_27151);
and U29002 (N_29002,N_28412,N_27163);
nor U29003 (N_29003,N_27870,N_28318);
nand U29004 (N_29004,N_27480,N_28129);
and U29005 (N_29005,N_27985,N_28024);
xnor U29006 (N_29006,N_27713,N_28231);
nand U29007 (N_29007,N_28228,N_27695);
or U29008 (N_29008,N_27179,N_27954);
and U29009 (N_29009,N_27421,N_27573);
or U29010 (N_29010,N_27986,N_27753);
or U29011 (N_29011,N_27706,N_27710);
xor U29012 (N_29012,N_28173,N_28120);
nand U29013 (N_29013,N_27191,N_27531);
or U29014 (N_29014,N_27914,N_27216);
and U29015 (N_29015,N_27803,N_27102);
and U29016 (N_29016,N_28086,N_27388);
or U29017 (N_29017,N_27239,N_28013);
xor U29018 (N_29018,N_27013,N_28101);
and U29019 (N_29019,N_27768,N_27026);
nor U29020 (N_29020,N_28378,N_27458);
nand U29021 (N_29021,N_28099,N_27415);
nand U29022 (N_29022,N_27691,N_27808);
or U29023 (N_29023,N_28482,N_27014);
xnor U29024 (N_29024,N_27158,N_27345);
nor U29025 (N_29025,N_28419,N_28447);
nand U29026 (N_29026,N_27682,N_28413);
xnor U29027 (N_29027,N_27185,N_28248);
xor U29028 (N_29028,N_27873,N_28216);
and U29029 (N_29029,N_28354,N_27844);
nor U29030 (N_29030,N_27133,N_27567);
nor U29031 (N_29031,N_27126,N_27890);
and U29032 (N_29032,N_27529,N_27041);
and U29033 (N_29033,N_27385,N_28269);
and U29034 (N_29034,N_28227,N_27070);
nor U29035 (N_29035,N_27967,N_28453);
xor U29036 (N_29036,N_27861,N_27838);
and U29037 (N_29037,N_27879,N_27298);
or U29038 (N_29038,N_27244,N_28382);
xnor U29039 (N_29039,N_27360,N_28416);
or U29040 (N_29040,N_27261,N_27569);
or U29041 (N_29041,N_27373,N_27201);
nor U29042 (N_29042,N_27377,N_27246);
or U29043 (N_29043,N_28076,N_27988);
nand U29044 (N_29044,N_28002,N_27702);
nor U29045 (N_29045,N_27558,N_27843);
xnor U29046 (N_29046,N_27265,N_27301);
or U29047 (N_29047,N_28471,N_28484);
or U29048 (N_29048,N_27761,N_27869);
xor U29049 (N_29049,N_27790,N_27598);
nor U29050 (N_29050,N_28057,N_27500);
nand U29051 (N_29051,N_27381,N_27550);
and U29052 (N_29052,N_27742,N_27926);
and U29053 (N_29053,N_27647,N_28446);
and U29054 (N_29054,N_27736,N_27050);
xnor U29055 (N_29055,N_27943,N_28081);
xnor U29056 (N_29056,N_27679,N_27541);
nand U29057 (N_29057,N_27592,N_28221);
and U29058 (N_29058,N_28356,N_27379);
xnor U29059 (N_29059,N_28325,N_28304);
nor U29060 (N_29060,N_27149,N_28473);
xor U29061 (N_29061,N_28145,N_28496);
nor U29062 (N_29062,N_27993,N_28041);
or U29063 (N_29063,N_28335,N_27346);
or U29064 (N_29064,N_28435,N_27453);
xor U29065 (N_29065,N_27805,N_28303);
xnor U29066 (N_29066,N_27422,N_27082);
nor U29067 (N_29067,N_28499,N_28035);
or U29068 (N_29068,N_28139,N_27420);
nand U29069 (N_29069,N_28327,N_27891);
or U29070 (N_29070,N_27308,N_27186);
and U29071 (N_29071,N_28320,N_27114);
nor U29072 (N_29072,N_27007,N_28111);
nor U29073 (N_29073,N_27155,N_27211);
nand U29074 (N_29074,N_28160,N_27724);
nor U29075 (N_29075,N_27490,N_27431);
or U29076 (N_29076,N_28258,N_27889);
nor U29077 (N_29077,N_28094,N_27335);
or U29078 (N_29078,N_28408,N_27897);
nor U29079 (N_29079,N_27248,N_27987);
and U29080 (N_29080,N_27826,N_27851);
and U29081 (N_29081,N_28103,N_28203);
nor U29082 (N_29082,N_28009,N_27251);
nor U29083 (N_29083,N_27619,N_28080);
nand U29084 (N_29084,N_27287,N_27907);
nor U29085 (N_29085,N_27996,N_28004);
or U29086 (N_29086,N_27131,N_28053);
or U29087 (N_29087,N_28161,N_28238);
and U29088 (N_29088,N_27218,N_27408);
nor U29089 (N_29089,N_27528,N_28459);
and U29090 (N_29090,N_27994,N_28268);
nand U29091 (N_29091,N_28342,N_27820);
xor U29092 (N_29092,N_28434,N_28245);
nand U29093 (N_29093,N_27555,N_28149);
or U29094 (N_29094,N_27217,N_27269);
nand U29095 (N_29095,N_27697,N_27532);
xor U29096 (N_29096,N_28313,N_27192);
nor U29097 (N_29097,N_27809,N_28078);
or U29098 (N_29098,N_28417,N_27657);
or U29099 (N_29099,N_28194,N_28070);
or U29100 (N_29100,N_27347,N_27884);
xnor U29101 (N_29101,N_28125,N_27609);
or U29102 (N_29102,N_27799,N_28082);
and U29103 (N_29103,N_28366,N_27038);
and U29104 (N_29104,N_28402,N_27830);
or U29105 (N_29105,N_27253,N_27639);
nor U29106 (N_29106,N_27673,N_28006);
xnor U29107 (N_29107,N_27354,N_28267);
nand U29108 (N_29108,N_27467,N_27812);
and U29109 (N_29109,N_27565,N_27725);
or U29110 (N_29110,N_27970,N_28064);
nand U29111 (N_29111,N_27536,N_27232);
xor U29112 (N_29112,N_27905,N_28442);
xor U29113 (N_29113,N_27486,N_27294);
or U29114 (N_29114,N_27010,N_28497);
xnor U29115 (N_29115,N_27498,N_28466);
nand U29116 (N_29116,N_28176,N_27402);
and U29117 (N_29117,N_27518,N_28379);
or U29118 (N_29118,N_27472,N_27350);
nor U29119 (N_29119,N_27210,N_27427);
and U29120 (N_29120,N_27332,N_27022);
nor U29121 (N_29121,N_28353,N_28411);
xnor U29122 (N_29122,N_27597,N_28498);
and U29123 (N_29123,N_28049,N_27277);
and U29124 (N_29124,N_27675,N_27543);
nand U29125 (N_29125,N_27168,N_27178);
and U29126 (N_29126,N_27765,N_27945);
nor U29127 (N_29127,N_28261,N_27764);
nand U29128 (N_29128,N_27825,N_27219);
or U29129 (N_29129,N_27887,N_27443);
and U29130 (N_29130,N_28481,N_27946);
and U29131 (N_29131,N_27902,N_27971);
xnor U29132 (N_29132,N_27515,N_27416);
nor U29133 (N_29133,N_28193,N_27522);
and U29134 (N_29134,N_27393,N_27846);
nand U29135 (N_29135,N_27067,N_28085);
nor U29136 (N_29136,N_28308,N_28212);
and U29137 (N_29137,N_28001,N_28061);
nor U29138 (N_29138,N_28233,N_28104);
nand U29139 (N_29139,N_28350,N_28395);
or U29140 (N_29140,N_27775,N_27860);
nand U29141 (N_29141,N_27628,N_28393);
nor U29142 (N_29142,N_27135,N_28074);
and U29143 (N_29143,N_27688,N_27165);
nor U29144 (N_29144,N_27468,N_28360);
and U29145 (N_29145,N_27722,N_27572);
nor U29146 (N_29146,N_27634,N_27212);
xnor U29147 (N_29147,N_27938,N_28224);
and U29148 (N_29148,N_28192,N_27002);
nor U29149 (N_29149,N_27723,N_27919);
or U29150 (N_29150,N_28124,N_27200);
or U29151 (N_29151,N_27835,N_28299);
xnor U29152 (N_29152,N_28200,N_28270);
xor U29153 (N_29153,N_27227,N_27570);
xnor U29154 (N_29154,N_27279,N_27032);
or U29155 (N_29155,N_27147,N_27208);
nand U29156 (N_29156,N_28361,N_28357);
nor U29157 (N_29157,N_27600,N_27547);
xnor U29158 (N_29158,N_27202,N_27318);
or U29159 (N_29159,N_27908,N_28279);
xnor U29160 (N_29160,N_27703,N_27645);
nand U29161 (N_29161,N_27505,N_27078);
and U29162 (N_29162,N_27276,N_27376);
xnor U29163 (N_29163,N_27882,N_28377);
or U29164 (N_29164,N_27492,N_28215);
nor U29165 (N_29165,N_28050,N_28338);
or U29166 (N_29166,N_27511,N_28364);
or U29167 (N_29167,N_27842,N_27920);
and U29168 (N_29168,N_28352,N_28467);
nor U29169 (N_29169,N_28021,N_27043);
nand U29170 (N_29170,N_27077,N_27139);
and U29171 (N_29171,N_27241,N_27804);
nand U29172 (N_29172,N_27676,N_27564);
nor U29173 (N_29173,N_27831,N_27116);
nand U29174 (N_29174,N_27641,N_27751);
xnor U29175 (N_29175,N_28265,N_27404);
or U29176 (N_29176,N_28186,N_28351);
or U29177 (N_29177,N_27474,N_27442);
nor U29178 (N_29178,N_28472,N_28118);
or U29179 (N_29179,N_27648,N_27520);
nor U29180 (N_29180,N_27763,N_28319);
or U29181 (N_29181,N_27744,N_27827);
nand U29182 (N_29182,N_27885,N_27585);
nand U29183 (N_29183,N_28223,N_27779);
nor U29184 (N_29184,N_27544,N_28390);
nand U29185 (N_29185,N_27405,N_27221);
nand U29186 (N_29186,N_27664,N_28394);
and U29187 (N_29187,N_28032,N_27430);
or U29188 (N_29188,N_27583,N_27797);
xnor U29189 (N_29189,N_28148,N_27485);
nor U29190 (N_29190,N_27577,N_28387);
or U29191 (N_29191,N_27310,N_27399);
xor U29192 (N_29192,N_27361,N_27496);
or U29193 (N_29193,N_27571,N_27974);
nor U29194 (N_29194,N_27857,N_27633);
and U29195 (N_29195,N_27209,N_28052);
nand U29196 (N_29196,N_28188,N_28183);
or U29197 (N_29197,N_27374,N_27858);
and U29198 (N_29198,N_27099,N_27409);
nor U29199 (N_29199,N_27866,N_28401);
and U29200 (N_29200,N_27822,N_27484);
and U29201 (N_29201,N_27853,N_28091);
nor U29202 (N_29202,N_27859,N_27578);
xor U29203 (N_29203,N_27079,N_27992);
nor U29204 (N_29204,N_27327,N_27626);
xor U29205 (N_29205,N_28405,N_27635);
and U29206 (N_29206,N_28457,N_28071);
nor U29207 (N_29207,N_28206,N_27160);
nor U29208 (N_29208,N_27199,N_28025);
nor U29209 (N_29209,N_28414,N_27599);
nand U29210 (N_29210,N_28023,N_28345);
and U29211 (N_29211,N_28474,N_27016);
xnor U29212 (N_29212,N_27268,N_28478);
nor U29213 (N_29213,N_27233,N_27745);
and U29214 (N_29214,N_27271,N_27958);
and U29215 (N_29215,N_28196,N_27684);
nor U29216 (N_29216,N_27535,N_28306);
and U29217 (N_29217,N_28135,N_27683);
xnor U29218 (N_29218,N_28144,N_28152);
xor U29219 (N_29219,N_27594,N_28062);
nor U29220 (N_29220,N_27755,N_27852);
xor U29221 (N_29221,N_28257,N_27968);
and U29222 (N_29222,N_27602,N_27150);
nand U29223 (N_29223,N_27334,N_27982);
and U29224 (N_29224,N_27263,N_28007);
nand U29225 (N_29225,N_28237,N_28168);
nand U29226 (N_29226,N_28220,N_28185);
xor U29227 (N_29227,N_28235,N_28410);
and U29228 (N_29228,N_28143,N_27054);
or U29229 (N_29229,N_27063,N_27630);
xor U29230 (N_29230,N_27894,N_28277);
xnor U29231 (N_29231,N_27364,N_27085);
and U29232 (N_29232,N_27447,N_27792);
xor U29233 (N_29233,N_28464,N_27620);
nor U29234 (N_29234,N_27756,N_27148);
nand U29235 (N_29235,N_27357,N_27551);
and U29236 (N_29236,N_27383,N_27874);
and U29237 (N_29237,N_27059,N_27618);
or U29238 (N_29238,N_28488,N_27686);
nor U29239 (N_29239,N_27220,N_27030);
nand U29240 (N_29240,N_27331,N_27960);
or U29241 (N_29241,N_27922,N_27784);
or U29242 (N_29242,N_27730,N_28225);
and U29243 (N_29243,N_27546,N_27194);
xor U29244 (N_29244,N_27624,N_27545);
and U29245 (N_29245,N_27166,N_28452);
and U29246 (N_29246,N_27183,N_27638);
and U29247 (N_29247,N_27687,N_27923);
nand U29248 (N_29248,N_28155,N_27760);
nand U29249 (N_29249,N_28430,N_28178);
or U29250 (N_29250,N_27784,N_27379);
or U29251 (N_29251,N_27756,N_27887);
and U29252 (N_29252,N_28318,N_27537);
nor U29253 (N_29253,N_27053,N_27345);
nor U29254 (N_29254,N_27130,N_27807);
xor U29255 (N_29255,N_27358,N_28138);
and U29256 (N_29256,N_27819,N_27700);
and U29257 (N_29257,N_28222,N_28158);
or U29258 (N_29258,N_28417,N_28304);
xor U29259 (N_29259,N_27930,N_27890);
nor U29260 (N_29260,N_27853,N_27473);
and U29261 (N_29261,N_28292,N_27576);
and U29262 (N_29262,N_27803,N_27401);
xnor U29263 (N_29263,N_28208,N_27523);
or U29264 (N_29264,N_27827,N_28152);
nor U29265 (N_29265,N_27868,N_27086);
xnor U29266 (N_29266,N_27369,N_27933);
nor U29267 (N_29267,N_27953,N_27990);
or U29268 (N_29268,N_28078,N_27472);
and U29269 (N_29269,N_27881,N_28047);
xor U29270 (N_29270,N_27603,N_28277);
and U29271 (N_29271,N_27797,N_27280);
and U29272 (N_29272,N_27035,N_27973);
nor U29273 (N_29273,N_28108,N_28193);
nand U29274 (N_29274,N_27526,N_27405);
nor U29275 (N_29275,N_27606,N_27226);
and U29276 (N_29276,N_27187,N_28435);
and U29277 (N_29277,N_27117,N_28097);
and U29278 (N_29278,N_28061,N_28088);
xnor U29279 (N_29279,N_27978,N_27799);
nor U29280 (N_29280,N_27751,N_27964);
or U29281 (N_29281,N_27469,N_28181);
xnor U29282 (N_29282,N_27601,N_28480);
or U29283 (N_29283,N_27431,N_28185);
xnor U29284 (N_29284,N_27680,N_27408);
nand U29285 (N_29285,N_28072,N_27582);
nand U29286 (N_29286,N_27007,N_28355);
nand U29287 (N_29287,N_28483,N_28442);
or U29288 (N_29288,N_27228,N_27470);
xor U29289 (N_29289,N_27044,N_27926);
and U29290 (N_29290,N_27145,N_28141);
nand U29291 (N_29291,N_28082,N_27663);
nor U29292 (N_29292,N_27618,N_27715);
nor U29293 (N_29293,N_27034,N_27265);
and U29294 (N_29294,N_27230,N_27051);
or U29295 (N_29295,N_27467,N_27520);
xor U29296 (N_29296,N_27492,N_27567);
xor U29297 (N_29297,N_27708,N_28126);
nor U29298 (N_29298,N_27114,N_27350);
and U29299 (N_29299,N_27163,N_27379);
and U29300 (N_29300,N_28141,N_27892);
and U29301 (N_29301,N_27675,N_28084);
and U29302 (N_29302,N_27330,N_27574);
nor U29303 (N_29303,N_27206,N_27037);
nand U29304 (N_29304,N_28487,N_27039);
nor U29305 (N_29305,N_27077,N_28376);
or U29306 (N_29306,N_27104,N_27037);
nand U29307 (N_29307,N_27273,N_27971);
and U29308 (N_29308,N_28408,N_28386);
xnor U29309 (N_29309,N_27612,N_27670);
or U29310 (N_29310,N_28226,N_27091);
nor U29311 (N_29311,N_28051,N_27721);
or U29312 (N_29312,N_27464,N_27864);
xor U29313 (N_29313,N_27914,N_27860);
nor U29314 (N_29314,N_27930,N_28288);
nand U29315 (N_29315,N_28078,N_27656);
nand U29316 (N_29316,N_27153,N_28408);
or U29317 (N_29317,N_27333,N_27086);
xnor U29318 (N_29318,N_27689,N_28023);
nor U29319 (N_29319,N_28416,N_27502);
xor U29320 (N_29320,N_27600,N_27805);
and U29321 (N_29321,N_28329,N_28235);
or U29322 (N_29322,N_27197,N_28227);
xor U29323 (N_29323,N_28110,N_28170);
or U29324 (N_29324,N_28381,N_28279);
and U29325 (N_29325,N_27290,N_27678);
and U29326 (N_29326,N_27979,N_27723);
nor U29327 (N_29327,N_28298,N_27720);
xnor U29328 (N_29328,N_27677,N_27304);
xnor U29329 (N_29329,N_27755,N_28064);
xor U29330 (N_29330,N_28485,N_27954);
nand U29331 (N_29331,N_27651,N_28156);
xnor U29332 (N_29332,N_27036,N_27257);
nor U29333 (N_29333,N_27067,N_27547);
nand U29334 (N_29334,N_27780,N_27758);
and U29335 (N_29335,N_27750,N_28217);
nor U29336 (N_29336,N_27075,N_27716);
or U29337 (N_29337,N_27647,N_27388);
xor U29338 (N_29338,N_27874,N_28149);
xnor U29339 (N_29339,N_27087,N_28207);
nand U29340 (N_29340,N_27386,N_27359);
nor U29341 (N_29341,N_27497,N_28153);
nor U29342 (N_29342,N_27178,N_27551);
nand U29343 (N_29343,N_27529,N_28167);
nor U29344 (N_29344,N_27344,N_27863);
nand U29345 (N_29345,N_28173,N_28283);
nor U29346 (N_29346,N_27982,N_27143);
nand U29347 (N_29347,N_27162,N_28371);
xnor U29348 (N_29348,N_27603,N_27242);
and U29349 (N_29349,N_27327,N_27242);
or U29350 (N_29350,N_27499,N_27004);
and U29351 (N_29351,N_27599,N_27464);
nand U29352 (N_29352,N_27800,N_27026);
xor U29353 (N_29353,N_27256,N_28313);
or U29354 (N_29354,N_27356,N_27535);
nand U29355 (N_29355,N_27849,N_27898);
nand U29356 (N_29356,N_28225,N_27996);
nand U29357 (N_29357,N_27061,N_27823);
xnor U29358 (N_29358,N_27132,N_28006);
and U29359 (N_29359,N_27591,N_27015);
nor U29360 (N_29360,N_28041,N_27100);
and U29361 (N_29361,N_27746,N_27897);
xor U29362 (N_29362,N_27745,N_28354);
xor U29363 (N_29363,N_27352,N_27608);
nor U29364 (N_29364,N_27735,N_27536);
xor U29365 (N_29365,N_27559,N_27489);
nand U29366 (N_29366,N_27083,N_27142);
nor U29367 (N_29367,N_27358,N_28153);
nor U29368 (N_29368,N_28445,N_27950);
xor U29369 (N_29369,N_28304,N_27615);
and U29370 (N_29370,N_27062,N_27730);
or U29371 (N_29371,N_27327,N_28491);
nor U29372 (N_29372,N_27787,N_27676);
or U29373 (N_29373,N_28320,N_28130);
or U29374 (N_29374,N_28045,N_27653);
nand U29375 (N_29375,N_27245,N_27267);
xnor U29376 (N_29376,N_28003,N_27127);
nor U29377 (N_29377,N_28236,N_27105);
or U29378 (N_29378,N_27638,N_27319);
and U29379 (N_29379,N_27347,N_28146);
nand U29380 (N_29380,N_27492,N_27902);
xnor U29381 (N_29381,N_28467,N_27147);
xnor U29382 (N_29382,N_28416,N_27395);
xor U29383 (N_29383,N_27847,N_28479);
nand U29384 (N_29384,N_28496,N_27918);
nand U29385 (N_29385,N_28213,N_27568);
xnor U29386 (N_29386,N_27847,N_27132);
nand U29387 (N_29387,N_27888,N_27335);
nand U29388 (N_29388,N_27247,N_28368);
or U29389 (N_29389,N_27517,N_27034);
and U29390 (N_29390,N_27777,N_27845);
or U29391 (N_29391,N_28168,N_27757);
or U29392 (N_29392,N_27548,N_28001);
or U29393 (N_29393,N_27281,N_27083);
and U29394 (N_29394,N_27672,N_27108);
nor U29395 (N_29395,N_28483,N_27420);
and U29396 (N_29396,N_28067,N_28077);
nor U29397 (N_29397,N_28083,N_27070);
xnor U29398 (N_29398,N_27414,N_28301);
and U29399 (N_29399,N_27674,N_27534);
nor U29400 (N_29400,N_28066,N_27705);
xnor U29401 (N_29401,N_28111,N_27992);
nor U29402 (N_29402,N_27910,N_27206);
and U29403 (N_29403,N_27163,N_28028);
xor U29404 (N_29404,N_27578,N_28264);
and U29405 (N_29405,N_27991,N_27972);
and U29406 (N_29406,N_28281,N_27771);
or U29407 (N_29407,N_27425,N_27550);
and U29408 (N_29408,N_27917,N_27321);
and U29409 (N_29409,N_28169,N_27668);
nor U29410 (N_29410,N_28113,N_27671);
nand U29411 (N_29411,N_27995,N_27476);
xnor U29412 (N_29412,N_28116,N_27766);
or U29413 (N_29413,N_28008,N_28192);
nand U29414 (N_29414,N_27974,N_27815);
nor U29415 (N_29415,N_28259,N_28195);
nand U29416 (N_29416,N_27498,N_28091);
xor U29417 (N_29417,N_27526,N_27913);
and U29418 (N_29418,N_28370,N_28187);
xor U29419 (N_29419,N_27773,N_27731);
nor U29420 (N_29420,N_27679,N_28305);
and U29421 (N_29421,N_27649,N_27638);
and U29422 (N_29422,N_27612,N_27700);
xor U29423 (N_29423,N_27507,N_27628);
and U29424 (N_29424,N_27290,N_27473);
nand U29425 (N_29425,N_27722,N_27187);
or U29426 (N_29426,N_27274,N_28291);
xnor U29427 (N_29427,N_27585,N_27940);
and U29428 (N_29428,N_28395,N_27322);
or U29429 (N_29429,N_27235,N_27842);
and U29430 (N_29430,N_27841,N_27058);
or U29431 (N_29431,N_28300,N_27012);
and U29432 (N_29432,N_27724,N_27011);
or U29433 (N_29433,N_27976,N_28354);
and U29434 (N_29434,N_27228,N_27216);
nor U29435 (N_29435,N_27409,N_28470);
xnor U29436 (N_29436,N_27925,N_27008);
nand U29437 (N_29437,N_27317,N_27539);
nand U29438 (N_29438,N_27427,N_27742);
xnor U29439 (N_29439,N_28442,N_27484);
and U29440 (N_29440,N_28369,N_27502);
xnor U29441 (N_29441,N_27711,N_27445);
nand U29442 (N_29442,N_27019,N_27969);
or U29443 (N_29443,N_27055,N_28248);
xnor U29444 (N_29444,N_28131,N_27151);
or U29445 (N_29445,N_27683,N_27202);
nand U29446 (N_29446,N_27447,N_27925);
and U29447 (N_29447,N_27349,N_28329);
and U29448 (N_29448,N_27577,N_27763);
or U29449 (N_29449,N_28291,N_27328);
xnor U29450 (N_29450,N_27295,N_27636);
nand U29451 (N_29451,N_28346,N_27801);
and U29452 (N_29452,N_27171,N_27614);
nand U29453 (N_29453,N_28344,N_27653);
and U29454 (N_29454,N_28296,N_27237);
nor U29455 (N_29455,N_28139,N_27045);
nor U29456 (N_29456,N_28039,N_27823);
xor U29457 (N_29457,N_27075,N_27178);
or U29458 (N_29458,N_27546,N_27774);
and U29459 (N_29459,N_28465,N_28107);
nor U29460 (N_29460,N_27433,N_28088);
or U29461 (N_29461,N_27084,N_28175);
xnor U29462 (N_29462,N_28216,N_28099);
or U29463 (N_29463,N_28435,N_28396);
nor U29464 (N_29464,N_28169,N_28419);
xor U29465 (N_29465,N_28103,N_27692);
nand U29466 (N_29466,N_28445,N_27058);
or U29467 (N_29467,N_27225,N_27960);
xnor U29468 (N_29468,N_27562,N_28390);
and U29469 (N_29469,N_27791,N_27924);
xnor U29470 (N_29470,N_28272,N_27912);
and U29471 (N_29471,N_28499,N_27747);
or U29472 (N_29472,N_27480,N_28356);
nand U29473 (N_29473,N_27623,N_28239);
nor U29474 (N_29474,N_27247,N_27891);
or U29475 (N_29475,N_28452,N_27053);
nor U29476 (N_29476,N_28337,N_27765);
nand U29477 (N_29477,N_28375,N_27262);
nand U29478 (N_29478,N_28222,N_27205);
nand U29479 (N_29479,N_28181,N_27683);
xor U29480 (N_29480,N_28296,N_27416);
nand U29481 (N_29481,N_28490,N_27537);
or U29482 (N_29482,N_27551,N_28296);
or U29483 (N_29483,N_28375,N_27500);
xnor U29484 (N_29484,N_27038,N_28095);
nor U29485 (N_29485,N_27495,N_27500);
xor U29486 (N_29486,N_28382,N_27071);
xnor U29487 (N_29487,N_28486,N_27003);
or U29488 (N_29488,N_27275,N_28263);
nor U29489 (N_29489,N_28347,N_28075);
and U29490 (N_29490,N_27998,N_28420);
nand U29491 (N_29491,N_27543,N_27622);
xnor U29492 (N_29492,N_27352,N_28130);
xor U29493 (N_29493,N_27450,N_27414);
xnor U29494 (N_29494,N_27045,N_27850);
or U29495 (N_29495,N_27537,N_28483);
or U29496 (N_29496,N_27670,N_28142);
and U29497 (N_29497,N_28440,N_27558);
and U29498 (N_29498,N_27920,N_27593);
nand U29499 (N_29499,N_27486,N_28335);
or U29500 (N_29500,N_27401,N_28315);
nor U29501 (N_29501,N_27885,N_27074);
nor U29502 (N_29502,N_27691,N_27188);
xor U29503 (N_29503,N_28042,N_27931);
nor U29504 (N_29504,N_28332,N_27608);
nor U29505 (N_29505,N_27972,N_27339);
or U29506 (N_29506,N_28219,N_27519);
nand U29507 (N_29507,N_28214,N_27970);
or U29508 (N_29508,N_28428,N_28109);
nor U29509 (N_29509,N_28072,N_27768);
or U29510 (N_29510,N_27016,N_27075);
nand U29511 (N_29511,N_27288,N_27503);
xnor U29512 (N_29512,N_27338,N_27890);
nor U29513 (N_29513,N_27649,N_27417);
or U29514 (N_29514,N_27327,N_27530);
or U29515 (N_29515,N_27494,N_27926);
and U29516 (N_29516,N_27547,N_27695);
nand U29517 (N_29517,N_27230,N_27552);
nand U29518 (N_29518,N_28104,N_28150);
nand U29519 (N_29519,N_27133,N_27604);
xnor U29520 (N_29520,N_28078,N_27939);
or U29521 (N_29521,N_27439,N_27908);
or U29522 (N_29522,N_27202,N_27256);
nand U29523 (N_29523,N_27632,N_28243);
nand U29524 (N_29524,N_27010,N_27471);
xor U29525 (N_29525,N_27306,N_28301);
and U29526 (N_29526,N_27973,N_27042);
or U29527 (N_29527,N_27457,N_28099);
nor U29528 (N_29528,N_28307,N_27515);
or U29529 (N_29529,N_28343,N_28403);
or U29530 (N_29530,N_27476,N_27443);
nor U29531 (N_29531,N_28353,N_27889);
xnor U29532 (N_29532,N_27856,N_27114);
or U29533 (N_29533,N_27890,N_28473);
nand U29534 (N_29534,N_27840,N_27419);
and U29535 (N_29535,N_27430,N_28440);
xnor U29536 (N_29536,N_27154,N_27173);
or U29537 (N_29537,N_27073,N_27731);
nand U29538 (N_29538,N_28248,N_28125);
xnor U29539 (N_29539,N_27289,N_27320);
and U29540 (N_29540,N_28176,N_27332);
xnor U29541 (N_29541,N_28158,N_27850);
and U29542 (N_29542,N_27060,N_28009);
nand U29543 (N_29543,N_27225,N_27419);
nand U29544 (N_29544,N_27687,N_27870);
and U29545 (N_29545,N_28304,N_27677);
or U29546 (N_29546,N_27368,N_27906);
xnor U29547 (N_29547,N_27938,N_27399);
or U29548 (N_29548,N_27975,N_28239);
and U29549 (N_29549,N_28313,N_28073);
xnor U29550 (N_29550,N_28021,N_27604);
xor U29551 (N_29551,N_27909,N_27789);
nor U29552 (N_29552,N_27558,N_27447);
and U29553 (N_29553,N_27957,N_27578);
and U29554 (N_29554,N_28469,N_27131);
xnor U29555 (N_29555,N_27638,N_28307);
and U29556 (N_29556,N_28219,N_27188);
xnor U29557 (N_29557,N_27868,N_28271);
and U29558 (N_29558,N_28218,N_27340);
nor U29559 (N_29559,N_27025,N_28069);
and U29560 (N_29560,N_27158,N_27165);
and U29561 (N_29561,N_28139,N_27314);
or U29562 (N_29562,N_27393,N_27592);
xnor U29563 (N_29563,N_28265,N_27707);
and U29564 (N_29564,N_27432,N_27667);
nor U29565 (N_29565,N_27968,N_27671);
nand U29566 (N_29566,N_27585,N_27164);
and U29567 (N_29567,N_27214,N_27841);
and U29568 (N_29568,N_27708,N_27762);
or U29569 (N_29569,N_27205,N_27518);
nor U29570 (N_29570,N_28115,N_28349);
nand U29571 (N_29571,N_27643,N_27362);
nor U29572 (N_29572,N_27797,N_27033);
or U29573 (N_29573,N_28447,N_27168);
nand U29574 (N_29574,N_28473,N_27564);
xnor U29575 (N_29575,N_27257,N_27334);
or U29576 (N_29576,N_27211,N_27316);
or U29577 (N_29577,N_27390,N_28362);
xor U29578 (N_29578,N_28440,N_28407);
xnor U29579 (N_29579,N_28395,N_27637);
or U29580 (N_29580,N_27561,N_27183);
or U29581 (N_29581,N_27934,N_28375);
and U29582 (N_29582,N_28093,N_28013);
and U29583 (N_29583,N_28291,N_27860);
and U29584 (N_29584,N_28045,N_27347);
nand U29585 (N_29585,N_28318,N_27648);
nand U29586 (N_29586,N_27991,N_28233);
and U29587 (N_29587,N_27614,N_27719);
nor U29588 (N_29588,N_28419,N_27111);
xor U29589 (N_29589,N_27908,N_28223);
or U29590 (N_29590,N_28161,N_27916);
xor U29591 (N_29591,N_27778,N_27133);
or U29592 (N_29592,N_27089,N_28346);
and U29593 (N_29593,N_27060,N_28064);
nor U29594 (N_29594,N_28397,N_28162);
xor U29595 (N_29595,N_27211,N_27152);
nand U29596 (N_29596,N_28177,N_27870);
nor U29597 (N_29597,N_27044,N_27872);
xnor U29598 (N_29598,N_27206,N_28066);
and U29599 (N_29599,N_27398,N_28337);
nand U29600 (N_29600,N_28069,N_27318);
and U29601 (N_29601,N_27264,N_27024);
or U29602 (N_29602,N_27784,N_28432);
nand U29603 (N_29603,N_27151,N_28180);
xor U29604 (N_29604,N_27596,N_27347);
nand U29605 (N_29605,N_28442,N_27322);
nand U29606 (N_29606,N_27399,N_27447);
nor U29607 (N_29607,N_27778,N_27338);
nand U29608 (N_29608,N_27521,N_28462);
xor U29609 (N_29609,N_28164,N_27125);
and U29610 (N_29610,N_28366,N_27509);
xor U29611 (N_29611,N_28136,N_27142);
or U29612 (N_29612,N_27418,N_27925);
and U29613 (N_29613,N_27695,N_28253);
or U29614 (N_29614,N_27554,N_28194);
xnor U29615 (N_29615,N_27398,N_27746);
and U29616 (N_29616,N_28153,N_27837);
nor U29617 (N_29617,N_27540,N_28149);
nand U29618 (N_29618,N_27445,N_27706);
and U29619 (N_29619,N_28098,N_27199);
nand U29620 (N_29620,N_28251,N_27068);
nand U29621 (N_29621,N_27063,N_27395);
and U29622 (N_29622,N_27600,N_27061);
or U29623 (N_29623,N_28102,N_27744);
and U29624 (N_29624,N_27823,N_28203);
or U29625 (N_29625,N_27422,N_27531);
nand U29626 (N_29626,N_27510,N_28051);
or U29627 (N_29627,N_27387,N_27143);
nor U29628 (N_29628,N_28245,N_27139);
or U29629 (N_29629,N_28375,N_28395);
or U29630 (N_29630,N_28126,N_27983);
nand U29631 (N_29631,N_28411,N_27121);
nor U29632 (N_29632,N_27962,N_27341);
nor U29633 (N_29633,N_28100,N_27401);
nand U29634 (N_29634,N_27293,N_28413);
nand U29635 (N_29635,N_28134,N_28321);
nor U29636 (N_29636,N_28115,N_27972);
and U29637 (N_29637,N_27110,N_27952);
nor U29638 (N_29638,N_27375,N_27175);
nand U29639 (N_29639,N_28192,N_27384);
nor U29640 (N_29640,N_28029,N_28161);
nand U29641 (N_29641,N_27480,N_27248);
nand U29642 (N_29642,N_27552,N_28253);
or U29643 (N_29643,N_27666,N_27085);
nand U29644 (N_29644,N_27261,N_27352);
nand U29645 (N_29645,N_27127,N_27099);
and U29646 (N_29646,N_28497,N_27335);
and U29647 (N_29647,N_27739,N_28464);
or U29648 (N_29648,N_27193,N_28263);
xor U29649 (N_29649,N_27893,N_28459);
or U29650 (N_29650,N_27592,N_27624);
xnor U29651 (N_29651,N_27032,N_27631);
nand U29652 (N_29652,N_27178,N_28356);
and U29653 (N_29653,N_27456,N_27567);
or U29654 (N_29654,N_28068,N_28260);
xnor U29655 (N_29655,N_27158,N_28209);
xnor U29656 (N_29656,N_27263,N_28466);
xnor U29657 (N_29657,N_27447,N_28357);
nand U29658 (N_29658,N_28255,N_27393);
nand U29659 (N_29659,N_28486,N_27832);
or U29660 (N_29660,N_28008,N_27864);
nand U29661 (N_29661,N_27665,N_27066);
nand U29662 (N_29662,N_28038,N_28092);
and U29663 (N_29663,N_27964,N_28135);
and U29664 (N_29664,N_28375,N_28052);
nand U29665 (N_29665,N_27989,N_27713);
nand U29666 (N_29666,N_27269,N_28390);
nor U29667 (N_29667,N_27875,N_27734);
or U29668 (N_29668,N_27116,N_27778);
xor U29669 (N_29669,N_28043,N_27769);
nor U29670 (N_29670,N_27490,N_27274);
or U29671 (N_29671,N_27590,N_27964);
xor U29672 (N_29672,N_28197,N_27715);
xor U29673 (N_29673,N_27958,N_27976);
or U29674 (N_29674,N_27388,N_27899);
xnor U29675 (N_29675,N_27001,N_27032);
and U29676 (N_29676,N_27944,N_27235);
nand U29677 (N_29677,N_28400,N_28289);
nor U29678 (N_29678,N_27464,N_27474);
and U29679 (N_29679,N_27650,N_27062);
or U29680 (N_29680,N_27532,N_28428);
nand U29681 (N_29681,N_28455,N_27325);
nand U29682 (N_29682,N_27841,N_28383);
nand U29683 (N_29683,N_27645,N_27303);
xor U29684 (N_29684,N_27772,N_28474);
nor U29685 (N_29685,N_27186,N_27214);
xnor U29686 (N_29686,N_27609,N_27841);
and U29687 (N_29687,N_27641,N_27169);
and U29688 (N_29688,N_28170,N_27595);
nor U29689 (N_29689,N_27175,N_27294);
nand U29690 (N_29690,N_28265,N_27825);
nand U29691 (N_29691,N_27742,N_27931);
nand U29692 (N_29692,N_27569,N_28405);
nor U29693 (N_29693,N_27878,N_28391);
xor U29694 (N_29694,N_27741,N_28195);
and U29695 (N_29695,N_27579,N_27756);
or U29696 (N_29696,N_28415,N_27458);
or U29697 (N_29697,N_27028,N_28131);
nor U29698 (N_29698,N_27187,N_27881);
nand U29699 (N_29699,N_27068,N_28226);
nand U29700 (N_29700,N_27435,N_28305);
nor U29701 (N_29701,N_27704,N_28048);
or U29702 (N_29702,N_27350,N_27771);
or U29703 (N_29703,N_27192,N_28053);
nor U29704 (N_29704,N_28287,N_27067);
xnor U29705 (N_29705,N_27121,N_27696);
xnor U29706 (N_29706,N_27359,N_27987);
nor U29707 (N_29707,N_27354,N_27036);
or U29708 (N_29708,N_28482,N_27768);
and U29709 (N_29709,N_27599,N_28477);
or U29710 (N_29710,N_28179,N_27395);
nor U29711 (N_29711,N_28272,N_27532);
xnor U29712 (N_29712,N_27555,N_27060);
and U29713 (N_29713,N_28263,N_28103);
xor U29714 (N_29714,N_27430,N_28111);
or U29715 (N_29715,N_27178,N_27367);
and U29716 (N_29716,N_27625,N_28117);
xnor U29717 (N_29717,N_27192,N_28361);
nand U29718 (N_29718,N_27687,N_27668);
and U29719 (N_29719,N_27262,N_27200);
and U29720 (N_29720,N_28417,N_28471);
and U29721 (N_29721,N_28342,N_27291);
xor U29722 (N_29722,N_28260,N_28182);
xnor U29723 (N_29723,N_27165,N_27236);
xor U29724 (N_29724,N_28345,N_27783);
or U29725 (N_29725,N_27284,N_27295);
xnor U29726 (N_29726,N_28239,N_27378);
nor U29727 (N_29727,N_28037,N_27150);
nor U29728 (N_29728,N_28094,N_27048);
and U29729 (N_29729,N_27200,N_27797);
and U29730 (N_29730,N_27801,N_27375);
and U29731 (N_29731,N_27229,N_27810);
and U29732 (N_29732,N_27713,N_27095);
or U29733 (N_29733,N_28058,N_28423);
or U29734 (N_29734,N_27834,N_28256);
nor U29735 (N_29735,N_28260,N_28221);
nor U29736 (N_29736,N_27915,N_27729);
nor U29737 (N_29737,N_27338,N_27265);
nor U29738 (N_29738,N_27248,N_27271);
or U29739 (N_29739,N_28151,N_27809);
nor U29740 (N_29740,N_27370,N_28102);
xnor U29741 (N_29741,N_27722,N_28137);
or U29742 (N_29742,N_27098,N_27862);
xor U29743 (N_29743,N_27659,N_27856);
nand U29744 (N_29744,N_27956,N_28363);
or U29745 (N_29745,N_27942,N_28495);
nand U29746 (N_29746,N_27894,N_28458);
nor U29747 (N_29747,N_28022,N_27941);
nand U29748 (N_29748,N_28220,N_27825);
or U29749 (N_29749,N_27436,N_27399);
xnor U29750 (N_29750,N_28143,N_27880);
or U29751 (N_29751,N_27258,N_27604);
and U29752 (N_29752,N_27744,N_28266);
xor U29753 (N_29753,N_27223,N_27713);
and U29754 (N_29754,N_27013,N_27246);
or U29755 (N_29755,N_27849,N_27766);
xnor U29756 (N_29756,N_27260,N_27008);
xnor U29757 (N_29757,N_27564,N_27029);
xnor U29758 (N_29758,N_28440,N_28141);
nand U29759 (N_29759,N_28418,N_27983);
or U29760 (N_29760,N_27424,N_27114);
or U29761 (N_29761,N_28466,N_28446);
xnor U29762 (N_29762,N_28095,N_27150);
nor U29763 (N_29763,N_28322,N_28126);
xor U29764 (N_29764,N_27132,N_27167);
nor U29765 (N_29765,N_27015,N_27714);
nor U29766 (N_29766,N_27158,N_27929);
or U29767 (N_29767,N_28031,N_27590);
nand U29768 (N_29768,N_27979,N_28157);
or U29769 (N_29769,N_28053,N_27254);
nor U29770 (N_29770,N_27209,N_27777);
and U29771 (N_29771,N_27890,N_27695);
nor U29772 (N_29772,N_27774,N_27364);
and U29773 (N_29773,N_27848,N_27501);
nand U29774 (N_29774,N_28311,N_28054);
and U29775 (N_29775,N_27873,N_27134);
and U29776 (N_29776,N_27235,N_27652);
and U29777 (N_29777,N_27115,N_28230);
nand U29778 (N_29778,N_28287,N_28017);
nor U29779 (N_29779,N_28259,N_27303);
and U29780 (N_29780,N_27553,N_28202);
and U29781 (N_29781,N_27588,N_27093);
nor U29782 (N_29782,N_27606,N_27868);
xnor U29783 (N_29783,N_28224,N_28319);
xnor U29784 (N_29784,N_27067,N_28480);
nor U29785 (N_29785,N_27089,N_27723);
xor U29786 (N_29786,N_27746,N_27262);
nand U29787 (N_29787,N_28340,N_28248);
nor U29788 (N_29788,N_27668,N_27491);
nor U29789 (N_29789,N_27439,N_28269);
or U29790 (N_29790,N_28002,N_27660);
xor U29791 (N_29791,N_27329,N_27813);
and U29792 (N_29792,N_28369,N_28429);
nand U29793 (N_29793,N_27429,N_27659);
nand U29794 (N_29794,N_27365,N_27755);
xnor U29795 (N_29795,N_28146,N_27627);
xnor U29796 (N_29796,N_27324,N_28275);
or U29797 (N_29797,N_27143,N_27084);
xor U29798 (N_29798,N_27506,N_27478);
nor U29799 (N_29799,N_27178,N_27379);
and U29800 (N_29800,N_27382,N_27754);
and U29801 (N_29801,N_27854,N_27570);
nand U29802 (N_29802,N_27446,N_28238);
or U29803 (N_29803,N_27375,N_27966);
and U29804 (N_29804,N_28268,N_27041);
xor U29805 (N_29805,N_27349,N_27892);
and U29806 (N_29806,N_28356,N_27172);
and U29807 (N_29807,N_28061,N_27593);
and U29808 (N_29808,N_27685,N_27478);
nor U29809 (N_29809,N_27794,N_28247);
nor U29810 (N_29810,N_28063,N_28013);
nand U29811 (N_29811,N_27515,N_28042);
and U29812 (N_29812,N_27866,N_27070);
or U29813 (N_29813,N_28387,N_28194);
xnor U29814 (N_29814,N_28115,N_27236);
xnor U29815 (N_29815,N_27820,N_27887);
nand U29816 (N_29816,N_28125,N_28262);
nor U29817 (N_29817,N_27104,N_27218);
nand U29818 (N_29818,N_27612,N_28392);
and U29819 (N_29819,N_27593,N_27086);
or U29820 (N_29820,N_27727,N_27047);
xnor U29821 (N_29821,N_27252,N_28299);
xor U29822 (N_29822,N_27179,N_27062);
nand U29823 (N_29823,N_27607,N_27701);
nand U29824 (N_29824,N_28482,N_27809);
nor U29825 (N_29825,N_27620,N_27544);
xor U29826 (N_29826,N_28211,N_27945);
nor U29827 (N_29827,N_27626,N_28270);
nand U29828 (N_29828,N_27832,N_27245);
nor U29829 (N_29829,N_27069,N_28127);
xor U29830 (N_29830,N_27577,N_27738);
nor U29831 (N_29831,N_27626,N_27768);
nor U29832 (N_29832,N_27100,N_28069);
xnor U29833 (N_29833,N_28473,N_28255);
nand U29834 (N_29834,N_27011,N_27149);
xor U29835 (N_29835,N_27767,N_27624);
nand U29836 (N_29836,N_27330,N_27303);
and U29837 (N_29837,N_28061,N_27123);
and U29838 (N_29838,N_28434,N_27901);
nand U29839 (N_29839,N_28205,N_28239);
nand U29840 (N_29840,N_27206,N_27561);
nor U29841 (N_29841,N_27330,N_27475);
and U29842 (N_29842,N_28179,N_27715);
xnor U29843 (N_29843,N_28395,N_28438);
nor U29844 (N_29844,N_28446,N_28499);
and U29845 (N_29845,N_28031,N_27046);
xor U29846 (N_29846,N_27787,N_27891);
or U29847 (N_29847,N_27519,N_27359);
nand U29848 (N_29848,N_27378,N_27037);
and U29849 (N_29849,N_27756,N_27050);
and U29850 (N_29850,N_27909,N_27011);
and U29851 (N_29851,N_27051,N_27417);
nor U29852 (N_29852,N_28413,N_27971);
nor U29853 (N_29853,N_27824,N_27310);
xnor U29854 (N_29854,N_27205,N_27372);
and U29855 (N_29855,N_28150,N_27619);
and U29856 (N_29856,N_27342,N_28476);
nor U29857 (N_29857,N_27717,N_28495);
or U29858 (N_29858,N_28423,N_27537);
nand U29859 (N_29859,N_28363,N_28322);
xnor U29860 (N_29860,N_28425,N_28277);
nand U29861 (N_29861,N_27869,N_27920);
nand U29862 (N_29862,N_28484,N_28015);
nor U29863 (N_29863,N_28208,N_27114);
nand U29864 (N_29864,N_27269,N_27010);
or U29865 (N_29865,N_27658,N_27741);
nand U29866 (N_29866,N_27163,N_27717);
nand U29867 (N_29867,N_28332,N_27981);
or U29868 (N_29868,N_27547,N_27532);
or U29869 (N_29869,N_27520,N_28092);
xor U29870 (N_29870,N_28087,N_27650);
xor U29871 (N_29871,N_28455,N_28158);
nor U29872 (N_29872,N_28129,N_27683);
or U29873 (N_29873,N_27484,N_28064);
xnor U29874 (N_29874,N_28302,N_27960);
xor U29875 (N_29875,N_28447,N_28198);
xor U29876 (N_29876,N_28185,N_27583);
nand U29877 (N_29877,N_28177,N_28014);
nand U29878 (N_29878,N_27147,N_27591);
nand U29879 (N_29879,N_27534,N_27058);
nand U29880 (N_29880,N_27283,N_28495);
nand U29881 (N_29881,N_27774,N_27895);
nor U29882 (N_29882,N_28061,N_27423);
xor U29883 (N_29883,N_28403,N_27334);
xor U29884 (N_29884,N_27906,N_27660);
nand U29885 (N_29885,N_27936,N_28422);
nand U29886 (N_29886,N_27326,N_27608);
xor U29887 (N_29887,N_27011,N_27726);
nor U29888 (N_29888,N_28128,N_28062);
xnor U29889 (N_29889,N_28393,N_28204);
nand U29890 (N_29890,N_27143,N_28383);
or U29891 (N_29891,N_27853,N_28306);
nor U29892 (N_29892,N_28005,N_27632);
nand U29893 (N_29893,N_28266,N_27209);
nand U29894 (N_29894,N_28194,N_27712);
or U29895 (N_29895,N_28079,N_28234);
nor U29896 (N_29896,N_28434,N_28048);
nand U29897 (N_29897,N_28339,N_27929);
xor U29898 (N_29898,N_28272,N_28130);
or U29899 (N_29899,N_27468,N_27297);
and U29900 (N_29900,N_27753,N_27352);
or U29901 (N_29901,N_28027,N_28371);
nor U29902 (N_29902,N_27243,N_27737);
xnor U29903 (N_29903,N_27511,N_27971);
nor U29904 (N_29904,N_27784,N_27549);
nand U29905 (N_29905,N_28344,N_28406);
xor U29906 (N_29906,N_27759,N_27483);
xnor U29907 (N_29907,N_27688,N_27530);
nand U29908 (N_29908,N_28316,N_27020);
nand U29909 (N_29909,N_27439,N_27537);
or U29910 (N_29910,N_27315,N_28406);
and U29911 (N_29911,N_27986,N_27899);
nor U29912 (N_29912,N_27234,N_27123);
and U29913 (N_29913,N_27095,N_27732);
nand U29914 (N_29914,N_27015,N_27908);
and U29915 (N_29915,N_27545,N_28204);
xnor U29916 (N_29916,N_28098,N_28344);
and U29917 (N_29917,N_28205,N_27749);
or U29918 (N_29918,N_27295,N_27043);
or U29919 (N_29919,N_28418,N_28002);
nor U29920 (N_29920,N_27492,N_28187);
xor U29921 (N_29921,N_27180,N_28286);
and U29922 (N_29922,N_28362,N_27840);
nand U29923 (N_29923,N_27707,N_27991);
xnor U29924 (N_29924,N_27405,N_28122);
nand U29925 (N_29925,N_27623,N_27086);
nor U29926 (N_29926,N_27029,N_27087);
or U29927 (N_29927,N_28201,N_28425);
nand U29928 (N_29928,N_27445,N_27515);
nand U29929 (N_29929,N_28164,N_27003);
or U29930 (N_29930,N_28281,N_27182);
and U29931 (N_29931,N_27781,N_27612);
and U29932 (N_29932,N_27184,N_27369);
and U29933 (N_29933,N_28444,N_27787);
and U29934 (N_29934,N_28382,N_28412);
xor U29935 (N_29935,N_27347,N_28298);
nand U29936 (N_29936,N_27390,N_27651);
nor U29937 (N_29937,N_27444,N_27977);
and U29938 (N_29938,N_27702,N_28373);
xor U29939 (N_29939,N_28442,N_28272);
nand U29940 (N_29940,N_28476,N_28478);
nand U29941 (N_29941,N_28181,N_27183);
or U29942 (N_29942,N_27134,N_27652);
or U29943 (N_29943,N_28231,N_28401);
and U29944 (N_29944,N_28154,N_28085);
or U29945 (N_29945,N_27019,N_27551);
and U29946 (N_29946,N_28130,N_27737);
and U29947 (N_29947,N_27976,N_27921);
and U29948 (N_29948,N_27309,N_27969);
and U29949 (N_29949,N_27550,N_27735);
xor U29950 (N_29950,N_27996,N_27414);
or U29951 (N_29951,N_27214,N_27369);
and U29952 (N_29952,N_28303,N_27954);
nor U29953 (N_29953,N_27410,N_27275);
nor U29954 (N_29954,N_28249,N_28136);
or U29955 (N_29955,N_28076,N_28327);
or U29956 (N_29956,N_28200,N_28140);
nand U29957 (N_29957,N_27993,N_28427);
and U29958 (N_29958,N_27444,N_28395);
nor U29959 (N_29959,N_27698,N_28220);
nand U29960 (N_29960,N_27262,N_27996);
and U29961 (N_29961,N_27904,N_27373);
nand U29962 (N_29962,N_28348,N_28290);
and U29963 (N_29963,N_27040,N_27938);
xor U29964 (N_29964,N_27165,N_27468);
and U29965 (N_29965,N_28432,N_27984);
nor U29966 (N_29966,N_28205,N_27352);
and U29967 (N_29967,N_27850,N_28042);
nor U29968 (N_29968,N_27362,N_27388);
and U29969 (N_29969,N_28305,N_27548);
and U29970 (N_29970,N_27609,N_28095);
nand U29971 (N_29971,N_27300,N_28411);
xor U29972 (N_29972,N_27016,N_27143);
nand U29973 (N_29973,N_27566,N_28428);
and U29974 (N_29974,N_27806,N_28300);
xnor U29975 (N_29975,N_27022,N_27033);
or U29976 (N_29976,N_27122,N_27538);
or U29977 (N_29977,N_27929,N_27023);
xor U29978 (N_29978,N_28419,N_28191);
nor U29979 (N_29979,N_27910,N_28339);
nand U29980 (N_29980,N_28137,N_27347);
nor U29981 (N_29981,N_27149,N_28207);
nor U29982 (N_29982,N_27098,N_28063);
nand U29983 (N_29983,N_27899,N_27785);
or U29984 (N_29984,N_27855,N_27456);
nor U29985 (N_29985,N_27176,N_27577);
and U29986 (N_29986,N_28393,N_28121);
or U29987 (N_29987,N_27927,N_27951);
and U29988 (N_29988,N_27522,N_27937);
nor U29989 (N_29989,N_28256,N_28277);
or U29990 (N_29990,N_28021,N_27858);
xor U29991 (N_29991,N_27525,N_27399);
and U29992 (N_29992,N_27701,N_27179);
nand U29993 (N_29993,N_27980,N_27162);
or U29994 (N_29994,N_27752,N_27075);
or U29995 (N_29995,N_28212,N_27296);
nor U29996 (N_29996,N_27202,N_27417);
nand U29997 (N_29997,N_27846,N_28121);
or U29998 (N_29998,N_27873,N_27071);
nand U29999 (N_29999,N_27120,N_27625);
nand UO_0 (O_0,N_29909,N_29523);
or UO_1 (O_1,N_28960,N_29275);
nor UO_2 (O_2,N_28830,N_29607);
nor UO_3 (O_3,N_29305,N_29257);
and UO_4 (O_4,N_29724,N_29211);
xnor UO_5 (O_5,N_29098,N_28521);
xor UO_6 (O_6,N_28745,N_29524);
xnor UO_7 (O_7,N_29267,N_28528);
nor UO_8 (O_8,N_29792,N_28545);
nor UO_9 (O_9,N_28571,N_28657);
or UO_10 (O_10,N_28766,N_28635);
nor UO_11 (O_11,N_29033,N_28692);
xor UO_12 (O_12,N_29201,N_29738);
nand UO_13 (O_13,N_29761,N_29590);
and UO_14 (O_14,N_29494,N_29695);
xnor UO_15 (O_15,N_29625,N_29018);
nand UO_16 (O_16,N_29003,N_29131);
and UO_17 (O_17,N_28877,N_29775);
or UO_18 (O_18,N_29173,N_29939);
and UO_19 (O_19,N_28770,N_29468);
and UO_20 (O_20,N_29973,N_28733);
or UO_21 (O_21,N_29671,N_29778);
and UO_22 (O_22,N_28682,N_28974);
nor UO_23 (O_23,N_28547,N_29285);
xnor UO_24 (O_24,N_29500,N_28985);
nor UO_25 (O_25,N_29965,N_29370);
and UO_26 (O_26,N_29447,N_29953);
nand UO_27 (O_27,N_29216,N_29774);
nand UO_28 (O_28,N_28947,N_28829);
xor UO_29 (O_29,N_29197,N_29437);
and UO_30 (O_30,N_29956,N_28640);
and UO_31 (O_31,N_29776,N_29927);
and UO_32 (O_32,N_29502,N_29052);
nor UO_33 (O_33,N_29470,N_29672);
nor UO_34 (O_34,N_29054,N_28567);
and UO_35 (O_35,N_29731,N_29568);
and UO_36 (O_36,N_29151,N_29519);
nor UO_37 (O_37,N_28645,N_29821);
nor UO_38 (O_38,N_28796,N_29260);
and UO_39 (O_39,N_28826,N_29846);
and UO_40 (O_40,N_29797,N_28563);
nand UO_41 (O_41,N_29988,N_28566);
xor UO_42 (O_42,N_29908,N_28973);
nand UO_43 (O_43,N_29628,N_28643);
xor UO_44 (O_44,N_28557,N_29357);
nor UO_45 (O_45,N_29273,N_28772);
xor UO_46 (O_46,N_29212,N_28734);
nand UO_47 (O_47,N_29990,N_29402);
xor UO_48 (O_48,N_28593,N_28506);
nand UO_49 (O_49,N_29472,N_29079);
and UO_50 (O_50,N_28831,N_29620);
or UO_51 (O_51,N_28648,N_28976);
and UO_52 (O_52,N_29220,N_29382);
nand UO_53 (O_53,N_28542,N_29691);
and UO_54 (O_54,N_28763,N_29159);
and UO_55 (O_55,N_29100,N_29160);
or UO_56 (O_56,N_28790,N_29594);
or UO_57 (O_57,N_29486,N_29873);
or UO_58 (O_58,N_29284,N_28711);
nand UO_59 (O_59,N_29036,N_29076);
and UO_60 (O_60,N_28505,N_29348);
nand UO_61 (O_61,N_29515,N_29541);
xnor UO_62 (O_62,N_28875,N_29898);
xnor UO_63 (O_63,N_29705,N_29204);
xor UO_64 (O_64,N_28750,N_29001);
nand UO_65 (O_65,N_29042,N_29392);
or UO_66 (O_66,N_29613,N_29750);
and UO_67 (O_67,N_29399,N_29442);
and UO_68 (O_68,N_29851,N_29393);
nand UO_69 (O_69,N_29600,N_29106);
xnor UO_70 (O_70,N_29194,N_28997);
and UO_71 (O_71,N_28760,N_28696);
or UO_72 (O_72,N_28769,N_29592);
xnor UO_73 (O_73,N_29896,N_29794);
nor UO_74 (O_74,N_29069,N_29654);
and UO_75 (O_75,N_28833,N_28848);
nor UO_76 (O_76,N_29129,N_29218);
nand UO_77 (O_77,N_29945,N_29187);
or UO_78 (O_78,N_29017,N_29553);
or UO_79 (O_79,N_29640,N_29058);
and UO_80 (O_80,N_29756,N_28922);
nand UO_81 (O_81,N_29090,N_29875);
nor UO_82 (O_82,N_28579,N_29698);
nand UO_83 (O_83,N_29149,N_29814);
or UO_84 (O_84,N_28749,N_28503);
nor UO_85 (O_85,N_29192,N_29591);
nand UO_86 (O_86,N_28511,N_29509);
nor UO_87 (O_87,N_29865,N_29274);
or UO_88 (O_88,N_28585,N_28556);
and UO_89 (O_89,N_29715,N_29006);
xnor UO_90 (O_90,N_29381,N_29292);
or UO_91 (O_91,N_29180,N_28927);
and UO_92 (O_92,N_28930,N_29475);
nand UO_93 (O_93,N_29632,N_29025);
or UO_94 (O_94,N_29853,N_28880);
xor UO_95 (O_95,N_29708,N_29164);
nand UO_96 (O_96,N_29200,N_28683);
or UO_97 (O_97,N_29935,N_28785);
and UO_98 (O_98,N_28607,N_29063);
xnor UO_99 (O_99,N_29765,N_29354);
xnor UO_100 (O_100,N_29810,N_28610);
xor UO_101 (O_101,N_28553,N_28820);
nor UO_102 (O_102,N_28951,N_28688);
nor UO_103 (O_103,N_29855,N_29035);
nor UO_104 (O_104,N_29377,N_28741);
and UO_105 (O_105,N_29168,N_29453);
or UO_106 (O_106,N_29233,N_29314);
xnor UO_107 (O_107,N_29718,N_29389);
or UO_108 (O_108,N_29940,N_29852);
nor UO_109 (O_109,N_29493,N_28946);
and UO_110 (O_110,N_29167,N_29499);
nand UO_111 (O_111,N_29330,N_29764);
or UO_112 (O_112,N_29638,N_29564);
nand UO_113 (O_113,N_29996,N_29007);
nand UO_114 (O_114,N_29914,N_28799);
or UO_115 (O_115,N_29078,N_28989);
nand UO_116 (O_116,N_29970,N_29126);
nand UO_117 (O_117,N_29408,N_28809);
or UO_118 (O_118,N_29240,N_28810);
nor UO_119 (O_119,N_28846,N_28726);
nor UO_120 (O_120,N_28834,N_29783);
or UO_121 (O_121,N_29202,N_28580);
nor UO_122 (O_122,N_29981,N_29758);
nand UO_123 (O_123,N_28982,N_29315);
nand UO_124 (O_124,N_28981,N_29045);
and UO_125 (O_125,N_28941,N_29575);
and UO_126 (O_126,N_29862,N_29527);
xor UO_127 (O_127,N_29107,N_28923);
and UO_128 (O_128,N_29642,N_29024);
nand UO_129 (O_129,N_29955,N_28870);
nor UO_130 (O_130,N_29977,N_28658);
or UO_131 (O_131,N_29184,N_29546);
xor UO_132 (O_132,N_29436,N_29863);
or UO_133 (O_133,N_29234,N_29390);
xnor UO_134 (O_134,N_29712,N_28709);
xor UO_135 (O_135,N_29349,N_28616);
and UO_136 (O_136,N_28937,N_29146);
nand UO_137 (O_137,N_29352,N_28746);
and UO_138 (O_138,N_29333,N_29105);
xnor UO_139 (O_139,N_29697,N_29368);
nor UO_140 (O_140,N_29322,N_29929);
nand UO_141 (O_141,N_28501,N_29605);
or UO_142 (O_142,N_29367,N_28592);
xor UO_143 (O_143,N_29872,N_29931);
nor UO_144 (O_144,N_28847,N_28597);
and UO_145 (O_145,N_29243,N_28878);
or UO_146 (O_146,N_29162,N_28732);
xnor UO_147 (O_147,N_29815,N_29842);
nand UO_148 (O_148,N_29729,N_29175);
and UO_149 (O_149,N_29646,N_29771);
and UO_150 (O_150,N_29089,N_29518);
and UO_151 (O_151,N_29190,N_29849);
or UO_152 (O_152,N_29743,N_29316);
xnor UO_153 (O_153,N_28980,N_28523);
nand UO_154 (O_154,N_28869,N_29210);
and UO_155 (O_155,N_29811,N_28715);
nand UO_156 (O_156,N_29868,N_28577);
or UO_157 (O_157,N_29356,N_29414);
or UO_158 (O_158,N_29166,N_29823);
nand UO_159 (O_159,N_29425,N_29951);
xnor UO_160 (O_160,N_29488,N_29959);
or UO_161 (O_161,N_28605,N_28817);
and UO_162 (O_162,N_29699,N_29336);
or UO_163 (O_163,N_29912,N_29982);
or UO_164 (O_164,N_29361,N_29533);
nand UO_165 (O_165,N_28558,N_29497);
nor UO_166 (O_166,N_28797,N_28686);
or UO_167 (O_167,N_29769,N_29287);
and UO_168 (O_168,N_29484,N_29682);
nand UO_169 (O_169,N_28704,N_28918);
nor UO_170 (O_170,N_29396,N_29338);
or UO_171 (O_171,N_29938,N_28589);
and UO_172 (O_172,N_29351,N_29680);
nor UO_173 (O_173,N_29154,N_28794);
and UO_174 (O_174,N_28910,N_29318);
and UO_175 (O_175,N_29727,N_29850);
and UO_176 (O_176,N_29586,N_29827);
xor UO_177 (O_177,N_28583,N_29644);
xnor UO_178 (O_178,N_29936,N_29504);
xor UO_179 (O_179,N_28990,N_29547);
nand UO_180 (O_180,N_28907,N_28689);
nand UO_181 (O_181,N_29016,N_29373);
xor UO_182 (O_182,N_29911,N_29817);
xor UO_183 (O_183,N_28572,N_29968);
nand UO_184 (O_184,N_29127,N_29961);
or UO_185 (O_185,N_28838,N_29398);
or UO_186 (O_186,N_28536,N_29165);
xor UO_187 (O_187,N_28892,N_29614);
or UO_188 (O_188,N_29177,N_29550);
or UO_189 (O_189,N_29919,N_29585);
xor UO_190 (O_190,N_29884,N_29269);
xor UO_191 (O_191,N_29302,N_29334);
xnor UO_192 (O_192,N_28762,N_29716);
nand UO_193 (O_193,N_29458,N_29156);
and UO_194 (O_194,N_29785,N_28620);
xnor UO_195 (O_195,N_29490,N_29920);
nand UO_196 (O_196,N_29601,N_29571);
nor UO_197 (O_197,N_28590,N_28828);
and UO_198 (O_198,N_29128,N_29508);
or UO_199 (O_199,N_29290,N_29678);
nand UO_200 (O_200,N_29028,N_29788);
nand UO_201 (O_201,N_29294,N_28791);
and UO_202 (O_202,N_29531,N_29023);
xnor UO_203 (O_203,N_29121,N_28768);
nor UO_204 (O_204,N_29557,N_29264);
or UO_205 (O_205,N_28964,N_29395);
and UO_206 (O_206,N_28986,N_29662);
xor UO_207 (O_207,N_29144,N_29913);
nor UO_208 (O_208,N_28897,N_29700);
nor UO_209 (O_209,N_29812,N_29748);
nor UO_210 (O_210,N_29781,N_28913);
nor UO_211 (O_211,N_28876,N_29065);
xor UO_212 (O_212,N_28613,N_28803);
and UO_213 (O_213,N_28824,N_29195);
xnor UO_214 (O_214,N_29083,N_29782);
or UO_215 (O_215,N_29015,N_28646);
and UO_216 (O_216,N_28578,N_29230);
or UO_217 (O_217,N_28518,N_28653);
nand UO_218 (O_218,N_29483,N_28871);
nor UO_219 (O_219,N_29856,N_28510);
and UO_220 (O_220,N_29498,N_29434);
nand UO_221 (O_221,N_29448,N_28759);
or UO_222 (O_222,N_29391,N_29692);
and UO_223 (O_223,N_29934,N_28984);
nand UO_224 (O_224,N_29635,N_28576);
xnor UO_225 (O_225,N_29525,N_29661);
or UO_226 (O_226,N_28669,N_28717);
xnor UO_227 (O_227,N_28540,N_29477);
or UO_228 (O_228,N_29561,N_28866);
nand UO_229 (O_229,N_28618,N_29304);
nor UO_230 (O_230,N_28912,N_28938);
nand UO_231 (O_231,N_29476,N_29784);
xor UO_232 (O_232,N_29344,N_29530);
xor UO_233 (O_233,N_29053,N_29343);
or UO_234 (O_234,N_29949,N_28595);
or UO_235 (O_235,N_29182,N_29994);
nor UO_236 (O_236,N_29624,N_29582);
nor UO_237 (O_237,N_29516,N_29051);
nand UO_238 (O_238,N_28958,N_29403);
nor UO_239 (O_239,N_29584,N_29118);
or UO_240 (O_240,N_29094,N_29169);
or UO_241 (O_241,N_28935,N_29213);
or UO_242 (O_242,N_29971,N_29907);
and UO_243 (O_243,N_29186,N_29379);
xor UO_244 (O_244,N_29219,N_28701);
xnor UO_245 (O_245,N_29378,N_29577);
and UO_246 (O_246,N_28743,N_28944);
xor UO_247 (O_247,N_28779,N_29835);
or UO_248 (O_248,N_28719,N_29365);
nor UO_249 (O_249,N_28537,N_28802);
or UO_250 (O_250,N_29313,N_28666);
and UO_251 (O_251,N_29746,N_28917);
and UO_252 (O_252,N_29460,N_29854);
nand UO_253 (O_253,N_29960,N_28647);
and UO_254 (O_254,N_29545,N_29183);
or UO_255 (O_255,N_29086,N_28783);
nand UO_256 (O_256,N_29627,N_28978);
or UO_257 (O_257,N_29658,N_29072);
nand UO_258 (O_258,N_28899,N_29848);
nor UO_259 (O_259,N_29215,N_29780);
nor UO_260 (O_260,N_29109,N_29890);
nand UO_261 (O_261,N_29371,N_29193);
or UO_262 (O_262,N_29095,N_29634);
or UO_263 (O_263,N_28955,N_28823);
and UO_264 (O_264,N_29674,N_29163);
nor UO_265 (O_265,N_29214,N_29196);
nand UO_266 (O_266,N_28681,N_29113);
xnor UO_267 (O_267,N_29623,N_28539);
nor UO_268 (O_268,N_28967,N_29300);
nor UO_269 (O_269,N_29103,N_28656);
nand UO_270 (O_270,N_28934,N_29013);
nand UO_271 (O_271,N_29085,N_29239);
and UO_272 (O_272,N_28994,N_28529);
or UO_273 (O_273,N_29102,N_29353);
nand UO_274 (O_274,N_29725,N_29535);
nand UO_275 (O_275,N_29819,N_29445);
or UO_276 (O_276,N_29657,N_29153);
xor UO_277 (O_277,N_29123,N_29521);
xnor UO_278 (O_278,N_29228,N_29917);
and UO_279 (O_279,N_28601,N_29062);
nand UO_280 (O_280,N_28588,N_28811);
nor UO_281 (O_281,N_29581,N_29655);
nor UO_282 (O_282,N_28806,N_28835);
and UO_283 (O_283,N_29122,N_28623);
xnor UO_284 (O_284,N_29070,N_29900);
and UO_285 (O_285,N_29363,N_29097);
and UO_286 (O_286,N_29728,N_29610);
and UO_287 (O_287,N_28805,N_28581);
and UO_288 (O_288,N_29717,N_28814);
nor UO_289 (O_289,N_29301,N_29805);
xnor UO_290 (O_290,N_29793,N_29384);
nand UO_291 (O_291,N_28965,N_28513);
or UO_292 (O_292,N_28586,N_28929);
or UO_293 (O_293,N_29005,N_28881);
and UO_294 (O_294,N_29226,N_28534);
xnor UO_295 (O_295,N_29950,N_28676);
nor UO_296 (O_296,N_29713,N_28840);
xnor UO_297 (O_297,N_29837,N_29155);
or UO_298 (O_298,N_29439,N_28628);
nand UO_299 (O_299,N_29060,N_28919);
nor UO_300 (O_300,N_29878,N_28856);
and UO_301 (O_301,N_29707,N_29622);
xnor UO_302 (O_302,N_29732,N_28611);
xnor UO_303 (O_303,N_28614,N_29432);
xnor UO_304 (O_304,N_28776,N_29138);
nor UO_305 (O_305,N_28694,N_29387);
or UO_306 (O_306,N_28707,N_29386);
and UO_307 (O_307,N_28854,N_29451);
and UO_308 (O_308,N_28525,N_29651);
nor UO_309 (O_309,N_29995,N_29847);
nand UO_310 (O_310,N_29752,N_29135);
xnor UO_311 (O_311,N_28924,N_28564);
xnor UO_312 (O_312,N_28544,N_29150);
or UO_313 (O_313,N_28861,N_29014);
or UO_314 (O_314,N_29510,N_29987);
or UO_315 (O_315,N_28873,N_29492);
and UO_316 (O_316,N_29174,N_29539);
nor UO_317 (O_317,N_29383,N_29282);
xnor UO_318 (O_318,N_29191,N_29004);
nand UO_319 (O_319,N_29760,N_29027);
xnor UO_320 (O_320,N_28690,N_29690);
xor UO_321 (O_321,N_29507,N_29554);
nand UO_322 (O_322,N_28863,N_28740);
or UO_323 (O_323,N_29091,N_29822);
and UO_324 (O_324,N_29059,N_28987);
xor UO_325 (O_325,N_28738,N_29721);
nor UO_326 (O_326,N_29286,N_29309);
nor UO_327 (O_327,N_29420,N_29572);
nand UO_328 (O_328,N_28526,N_28890);
nor UO_329 (O_329,N_29740,N_29522);
nand UO_330 (O_330,N_29719,N_29667);
xnor UO_331 (O_331,N_29972,N_29242);
and UO_332 (O_332,N_28889,N_29019);
nor UO_333 (O_333,N_29465,N_29400);
nand UO_334 (O_334,N_28971,N_29943);
xor UO_335 (O_335,N_29040,N_28995);
or UO_336 (O_336,N_29474,N_28520);
xnor UO_337 (O_337,N_28668,N_29566);
nand UO_338 (O_338,N_29710,N_29653);
and UO_339 (O_339,N_29388,N_28655);
and UO_340 (O_340,N_28731,N_29340);
xnor UO_341 (O_341,N_29558,N_29983);
nor UO_342 (O_342,N_29355,N_29733);
and UO_343 (O_343,N_29735,N_29992);
or UO_344 (O_344,N_29997,N_28742);
nand UO_345 (O_345,N_29247,N_29830);
and UO_346 (O_346,N_29542,N_29906);
nand UO_347 (O_347,N_29406,N_29171);
nand UO_348 (O_348,N_29636,N_28651);
nor UO_349 (O_349,N_29328,N_28781);
nor UO_350 (O_350,N_29454,N_29469);
or UO_351 (O_351,N_29009,N_29012);
and UO_352 (O_352,N_29142,N_29485);
nand UO_353 (O_353,N_29583,N_29362);
or UO_354 (O_354,N_29463,N_29626);
and UO_355 (O_355,N_29404,N_28954);
or UO_356 (O_356,N_29459,N_29844);
or UO_357 (O_357,N_28562,N_29329);
xnor UO_358 (O_358,N_29332,N_28702);
or UO_359 (O_359,N_29963,N_29528);
or UO_360 (O_360,N_29739,N_28902);
and UO_361 (O_361,N_29134,N_29081);
nor UO_362 (O_362,N_29573,N_28722);
or UO_363 (O_363,N_29244,N_29092);
nor UO_364 (O_364,N_28568,N_28737);
xnor UO_365 (O_365,N_29958,N_29181);
nor UO_366 (O_366,N_29962,N_28561);
or UO_367 (O_367,N_29172,N_29857);
or UO_368 (O_368,N_29077,N_28975);
and UO_369 (O_369,N_28793,N_29471);
nor UO_370 (O_370,N_29580,N_29669);
nor UO_371 (O_371,N_28718,N_28920);
nand UO_372 (O_372,N_29231,N_29339);
nand UO_373 (O_373,N_29777,N_28514);
and UO_374 (O_374,N_29238,N_28667);
and UO_375 (O_375,N_28533,N_28724);
and UO_376 (O_376,N_28691,N_29495);
and UO_377 (O_377,N_29446,N_28560);
nor UO_378 (O_378,N_29041,N_28721);
xor UO_379 (O_379,N_29262,N_29986);
and UO_380 (O_380,N_28596,N_28940);
nand UO_381 (O_381,N_29899,N_28860);
xnor UO_382 (O_382,N_29256,N_29457);
and UO_383 (O_383,N_28789,N_28903);
or UO_384 (O_384,N_29029,N_29616);
and UO_385 (O_385,N_28661,N_29800);
and UO_386 (O_386,N_28700,N_29589);
and UO_387 (O_387,N_29125,N_28550);
xor UO_388 (O_388,N_29540,N_28801);
and UO_389 (O_389,N_29306,N_28538);
nor UO_390 (O_390,N_28959,N_29737);
nor UO_391 (O_391,N_29241,N_29845);
xor UO_392 (O_392,N_29124,N_29071);
nor UO_393 (O_393,N_29902,N_29688);
or UO_394 (O_394,N_29544,N_29073);
or UO_395 (O_395,N_28798,N_29574);
xnor UO_396 (O_396,N_29277,N_29517);
xnor UO_397 (O_397,N_28808,N_29503);
nor UO_398 (O_398,N_29158,N_28603);
nand UO_399 (O_399,N_29754,N_29803);
or UO_400 (O_400,N_29350,N_28756);
or UO_401 (O_401,N_29619,N_29770);
xor UO_402 (O_402,N_29461,N_29422);
nand UO_403 (O_403,N_28604,N_28627);
nor UO_404 (O_404,N_29871,N_29978);
nor UO_405 (O_405,N_28859,N_28736);
xor UO_406 (O_406,N_28852,N_29345);
or UO_407 (O_407,N_28758,N_28939);
and UO_408 (O_408,N_28548,N_29789);
xnor UO_409 (O_409,N_29966,N_28530);
xor UO_410 (O_410,N_29321,N_28509);
or UO_411 (O_411,N_29551,N_29002);
nor UO_412 (O_412,N_29813,N_29921);
nor UO_413 (O_413,N_29888,N_29762);
or UO_414 (O_414,N_28842,N_29555);
and UO_415 (O_415,N_29820,N_29272);
or UO_416 (O_416,N_29808,N_29993);
nor UO_417 (O_417,N_28624,N_29643);
nand UO_418 (O_418,N_29787,N_29511);
nand UO_419 (O_419,N_29745,N_29675);
or UO_420 (O_420,N_29254,N_29520);
or UO_421 (O_421,N_28712,N_29679);
nand UO_422 (O_422,N_29417,N_29380);
xor UO_423 (O_423,N_29056,N_29877);
nand UO_424 (O_424,N_28839,N_28699);
and UO_425 (O_425,N_29137,N_29189);
or UO_426 (O_426,N_29407,N_29008);
and UO_427 (O_427,N_29630,N_28952);
and UO_428 (O_428,N_29341,N_29308);
nand UO_429 (O_429,N_29376,N_28804);
and UO_430 (O_430,N_28950,N_29617);
and UO_431 (O_431,N_28754,N_29609);
xor UO_432 (O_432,N_29816,N_29409);
and UO_433 (O_433,N_29714,N_29491);
xnor UO_434 (O_434,N_29998,N_29549);
nand UO_435 (O_435,N_29882,N_28629);
or UO_436 (O_436,N_29067,N_29093);
or UO_437 (O_437,N_29299,N_29394);
and UO_438 (O_438,N_29905,N_28713);
nor UO_439 (O_439,N_29763,N_29869);
nor UO_440 (O_440,N_28502,N_28851);
xnor UO_441 (O_441,N_28551,N_28874);
and UO_442 (O_442,N_29602,N_29178);
nor UO_443 (O_443,N_29964,N_29369);
or UO_444 (O_444,N_28634,N_29289);
and UO_445 (O_445,N_28723,N_29536);
nand UO_446 (O_446,N_28757,N_28504);
xnor UO_447 (O_447,N_28761,N_29225);
nand UO_448 (O_448,N_28541,N_29578);
nor UO_449 (O_449,N_29032,N_29064);
nor UO_450 (O_450,N_29119,N_28784);
and UO_451 (O_451,N_29832,N_28915);
xnor UO_452 (O_452,N_28821,N_29147);
xor UO_453 (O_453,N_29587,N_29283);
nor UO_454 (O_454,N_29298,N_29188);
xnor UO_455 (O_455,N_28896,N_28948);
nand UO_456 (O_456,N_28708,N_29450);
or UO_457 (O_457,N_29615,N_29276);
xor UO_458 (O_458,N_28966,N_29412);
xnor UO_459 (O_459,N_28853,N_29595);
nand UO_460 (O_460,N_28895,N_29596);
nor UO_461 (O_461,N_29824,N_29883);
xnor UO_462 (O_462,N_28633,N_29799);
xnor UO_463 (O_463,N_29199,N_29747);
xnor UO_464 (O_464,N_29798,N_28570);
xor UO_465 (O_465,N_29428,N_29433);
and UO_466 (O_466,N_29604,N_28705);
or UO_467 (O_467,N_29980,N_29924);
and UO_468 (O_468,N_28687,N_28664);
or UO_469 (O_469,N_28972,N_28926);
and UO_470 (O_470,N_29834,N_29757);
and UO_471 (O_471,N_28632,N_29647);
nor UO_472 (O_472,N_29809,N_28788);
nand UO_473 (O_473,N_28622,N_29804);
or UO_474 (O_474,N_29829,N_28963);
and UO_475 (O_475,N_29741,N_29796);
xnor UO_476 (O_476,N_28698,N_29424);
or UO_477 (O_477,N_28898,N_29826);
nor UO_478 (O_478,N_29038,N_28884);
xor UO_479 (O_479,N_29423,N_29297);
and UO_480 (O_480,N_29744,N_28559);
and UO_481 (O_481,N_29429,N_28663);
or UO_482 (O_482,N_28706,N_29320);
nor UO_483 (O_483,N_28642,N_29359);
nand UO_484 (O_484,N_29020,N_29331);
xnor UO_485 (O_485,N_28816,N_28905);
nor UO_486 (O_486,N_29880,N_28775);
or UO_487 (O_487,N_29117,N_29974);
and UO_488 (O_488,N_28591,N_28879);
xnor UO_489 (O_489,N_29133,N_29891);
xor UO_490 (O_490,N_29327,N_29270);
and UO_491 (O_491,N_29694,N_28906);
or UO_492 (O_492,N_28693,N_28991);
or UO_493 (O_493,N_29224,N_29656);
or UO_494 (O_494,N_28836,N_29456);
xor UO_495 (O_495,N_29579,N_28729);
nor UO_496 (O_496,N_28673,N_28925);
or UO_497 (O_497,N_29157,N_28956);
xor UO_498 (O_498,N_28787,N_29074);
nor UO_499 (O_499,N_29670,N_29496);
nor UO_500 (O_500,N_29532,N_29206);
and UO_501 (O_501,N_29026,N_29588);
nor UO_502 (O_502,N_29802,N_29405);
nor UO_503 (O_503,N_29879,N_29480);
nor UO_504 (O_504,N_29537,N_29481);
nand UO_505 (O_505,N_29258,N_28858);
or UO_506 (O_506,N_28600,N_29598);
and UO_507 (O_507,N_28630,N_29702);
or UO_508 (O_508,N_29082,N_29538);
or UO_509 (O_509,N_29176,N_29841);
nor UO_510 (O_510,N_28644,N_29985);
or UO_511 (O_511,N_28886,N_29720);
nor UO_512 (O_512,N_28771,N_28680);
or UO_513 (O_513,N_28998,N_28818);
nand UO_514 (O_514,N_29110,N_29952);
nand UO_515 (O_515,N_29031,N_29099);
and UO_516 (O_516,N_28662,N_29111);
xor UO_517 (O_517,N_28710,N_29999);
nand UO_518 (O_518,N_28827,N_29291);
and UO_519 (O_519,N_29790,N_29957);
nand UO_520 (O_520,N_28774,N_29932);
or UO_521 (O_521,N_29366,N_28594);
or UO_522 (O_522,N_29360,N_28739);
nor UO_523 (O_523,N_29043,N_29597);
nand UO_524 (O_524,N_29565,N_29413);
or UO_525 (O_525,N_28862,N_29203);
xor UO_526 (O_526,N_29385,N_29317);
nor UO_527 (O_527,N_29441,N_28598);
and UO_528 (O_528,N_29037,N_29892);
xnor UO_529 (O_529,N_29818,N_28507);
or UO_530 (O_530,N_29222,N_28650);
and UO_531 (O_531,N_28638,N_28641);
nor UO_532 (O_532,N_29839,N_29969);
nand UO_533 (O_533,N_28850,N_29021);
or UO_534 (O_534,N_29648,N_28970);
xor UO_535 (O_535,N_28532,N_28867);
or UO_536 (O_536,N_29645,N_28639);
and UO_537 (O_537,N_29411,N_29288);
xor UO_538 (O_538,N_29268,N_29055);
xor UO_539 (O_539,N_28602,N_29666);
or UO_540 (O_540,N_28744,N_29438);
or UO_541 (O_541,N_29979,N_29556);
and UO_542 (O_542,N_29473,N_29759);
nor UO_543 (O_543,N_28637,N_29926);
xnor UO_544 (O_544,N_28909,N_29681);
xor UO_545 (O_545,N_29044,N_29342);
nand UO_546 (O_546,N_29548,N_29120);
nand UO_547 (O_547,N_29736,N_29944);
and UO_548 (O_548,N_29910,N_29140);
xnor UO_549 (O_549,N_29840,N_28730);
and UO_550 (O_550,N_29335,N_29132);
xnor UO_551 (O_551,N_29751,N_28543);
or UO_552 (O_552,N_28697,N_28936);
nand UO_553 (O_553,N_29726,N_28845);
nor UO_554 (O_554,N_29066,N_28765);
xor UO_555 (O_555,N_29410,N_29552);
or UO_556 (O_556,N_28883,N_29255);
nand UO_557 (O_557,N_29312,N_29375);
and UO_558 (O_558,N_28949,N_29593);
nand UO_559 (O_559,N_29084,N_29989);
nor UO_560 (O_560,N_28764,N_29916);
xor UO_561 (O_561,N_29723,N_28996);
nor UO_562 (O_562,N_29806,N_28555);
nor UO_563 (O_563,N_28901,N_29709);
and UO_564 (O_564,N_29543,N_29440);
and UO_565 (O_565,N_28928,N_29534);
nor UO_566 (O_566,N_28612,N_28515);
and UO_567 (O_567,N_28961,N_29684);
or UO_568 (O_568,N_28968,N_29374);
nor UO_569 (O_569,N_29325,N_29876);
or UO_570 (O_570,N_29941,N_29416);
and UO_571 (O_571,N_29722,N_28777);
nor UO_572 (O_572,N_29567,N_28979);
or UO_573 (O_573,N_29000,N_28795);
nor UO_574 (O_574,N_29612,N_28815);
nand UO_575 (O_575,N_28606,N_28773);
xor UO_576 (O_576,N_29034,N_28625);
nor UO_577 (O_577,N_29418,N_29833);
xnor UO_578 (O_578,N_28675,N_28512);
and UO_579 (O_579,N_29659,N_29886);
or UO_580 (O_580,N_29462,N_28685);
xnor UO_581 (O_581,N_29665,N_29807);
and UO_582 (O_582,N_28660,N_29749);
and UO_583 (O_583,N_28582,N_28868);
xor UO_584 (O_584,N_29734,N_28516);
and UO_585 (O_585,N_29112,N_29148);
nor UO_586 (O_586,N_29831,N_29265);
nand UO_587 (O_587,N_29650,N_29246);
or UO_588 (O_588,N_29867,N_28931);
xnor UO_589 (O_589,N_29161,N_29293);
nand UO_590 (O_590,N_28751,N_29562);
or UO_591 (O_591,N_29772,N_28969);
and UO_592 (O_592,N_28665,N_28865);
and UO_593 (O_593,N_28916,N_29467);
nand UO_594 (O_594,N_29621,N_28893);
and UO_595 (O_595,N_29271,N_28755);
xor UO_596 (O_596,N_29307,N_29928);
nor UO_597 (O_597,N_28945,N_28843);
nor UO_598 (O_598,N_29514,N_29633);
or UO_599 (O_599,N_28908,N_29208);
or UO_600 (O_600,N_29742,N_28631);
xor UO_601 (O_601,N_29311,N_29050);
or UO_602 (O_602,N_29179,N_29730);
nand UO_603 (O_603,N_29889,N_29608);
or UO_604 (O_604,N_29116,N_28911);
nand UO_605 (O_605,N_29337,N_29221);
nand UO_606 (O_606,N_28569,N_29046);
xnor UO_607 (O_607,N_29431,N_29925);
nor UO_608 (O_608,N_28747,N_29048);
nand UO_609 (O_609,N_29791,N_28584);
nand UO_610 (O_610,N_28609,N_29894);
and UO_611 (O_611,N_29237,N_28753);
or UO_612 (O_612,N_29205,N_28999);
or UO_613 (O_613,N_29114,N_29143);
nand UO_614 (O_614,N_28531,N_29703);
or UO_615 (O_615,N_29505,N_28554);
or UO_616 (O_616,N_28894,N_28678);
or UO_617 (O_617,N_28857,N_28933);
or UO_618 (O_618,N_29825,N_28552);
nand UO_619 (O_619,N_29030,N_28962);
nand UO_620 (O_620,N_29755,N_28573);
nand UO_621 (O_621,N_29087,N_29130);
nand UO_622 (O_622,N_29115,N_29660);
and UO_623 (O_623,N_28695,N_29874);
and UO_624 (O_624,N_29415,N_29047);
nor UO_625 (O_625,N_28812,N_29466);
and UO_626 (O_626,N_29088,N_28619);
nor UO_627 (O_627,N_28659,N_29435);
or UO_628 (O_628,N_29768,N_29506);
nor UO_629 (O_629,N_28508,N_28546);
xnor UO_630 (O_630,N_28636,N_29096);
or UO_631 (O_631,N_29893,N_28983);
nand UO_632 (O_632,N_29198,N_29022);
nand UO_633 (O_633,N_28932,N_28716);
nor UO_634 (O_634,N_29346,N_28957);
or UO_635 (O_635,N_29637,N_28674);
and UO_636 (O_636,N_28587,N_29010);
nor UO_637 (O_637,N_29049,N_28778);
xor UO_638 (O_638,N_29559,N_28837);
nor UO_639 (O_639,N_29947,N_28819);
xnor UO_640 (O_640,N_28807,N_29364);
or UO_641 (O_641,N_29779,N_29946);
xnor UO_642 (O_642,N_29248,N_28519);
nor UO_643 (O_643,N_28615,N_28864);
nor UO_644 (O_644,N_29828,N_29421);
or UO_645 (O_645,N_28844,N_29933);
nor UO_646 (O_646,N_29280,N_29786);
and UO_647 (O_647,N_29209,N_29245);
and UO_648 (O_648,N_29901,N_29080);
or UO_649 (O_649,N_29039,N_28599);
and UO_650 (O_650,N_28621,N_29139);
xor UO_651 (O_651,N_28992,N_28677);
xor UO_652 (O_652,N_29217,N_29185);
xnor UO_653 (O_653,N_28822,N_29766);
nor UO_654 (O_654,N_28574,N_29108);
nand UO_655 (O_655,N_29948,N_29075);
or UO_656 (O_656,N_28953,N_28780);
nand UO_657 (O_657,N_29296,N_29903);
or UO_658 (O_658,N_29859,N_28703);
and UO_659 (O_659,N_28841,N_29685);
nor UO_660 (O_660,N_29881,N_29937);
or UO_661 (O_661,N_29991,N_29278);
and UO_662 (O_662,N_29897,N_29836);
or UO_663 (O_663,N_29606,N_29560);
and UO_664 (O_664,N_29136,N_28832);
nand UO_665 (O_665,N_29649,N_29922);
and UO_666 (O_666,N_29870,N_29864);
nor UO_667 (O_667,N_28943,N_28671);
xor UO_668 (O_668,N_29455,N_28527);
nor UO_669 (O_669,N_29487,N_29529);
nand UO_670 (O_670,N_28522,N_29310);
nand UO_671 (O_671,N_29673,N_29235);
or UO_672 (O_672,N_29773,N_29860);
nand UO_673 (O_673,N_29478,N_29319);
or UO_674 (O_674,N_28670,N_29279);
or UO_675 (O_675,N_29693,N_28900);
nor UO_676 (O_676,N_28988,N_29639);
and UO_677 (O_677,N_29430,N_29101);
or UO_678 (O_678,N_28565,N_28649);
or UO_679 (O_679,N_29141,N_29942);
or UO_680 (O_680,N_28748,N_29753);
and UO_681 (O_681,N_29570,N_29683);
xnor UO_682 (O_682,N_29858,N_28575);
or UO_683 (O_683,N_28887,N_29664);
xor UO_684 (O_684,N_28714,N_29631);
and UO_685 (O_685,N_29887,N_29569);
nand UO_686 (O_686,N_29687,N_28767);
nor UO_687 (O_687,N_29207,N_28725);
or UO_688 (O_688,N_29426,N_29711);
nand UO_689 (O_689,N_28617,N_29427);
nand UO_690 (O_690,N_29249,N_29295);
xor UO_691 (O_691,N_29629,N_29904);
or UO_692 (O_692,N_28720,N_29915);
nor UO_693 (O_693,N_29689,N_28849);
xnor UO_694 (O_694,N_29263,N_29686);
and UO_695 (O_695,N_28728,N_28825);
nand UO_696 (O_696,N_29861,N_29261);
nor UO_697 (O_697,N_29838,N_28855);
nand UO_698 (O_698,N_29252,N_29251);
xor UO_699 (O_699,N_28684,N_29061);
and UO_700 (O_700,N_29324,N_29843);
xnor UO_701 (O_701,N_28921,N_29223);
nor UO_702 (O_702,N_29401,N_28727);
and UO_703 (O_703,N_28993,N_28608);
or UO_704 (O_704,N_29145,N_29975);
nand UO_705 (O_705,N_29885,N_29563);
and UO_706 (O_706,N_29236,N_29419);
or UO_707 (O_707,N_29967,N_29652);
nor UO_708 (O_708,N_29326,N_29676);
nand UO_709 (O_709,N_29266,N_28672);
nor UO_710 (O_710,N_29923,N_29347);
or UO_711 (O_711,N_29011,N_29866);
nor UO_712 (O_712,N_28652,N_29303);
nand UO_713 (O_713,N_29229,N_29663);
and UO_714 (O_714,N_29930,N_29057);
or UO_715 (O_715,N_29767,N_29512);
or UO_716 (O_716,N_28914,N_28813);
nand UO_717 (O_717,N_28782,N_28679);
or UO_718 (O_718,N_29599,N_29618);
nand UO_719 (O_719,N_29281,N_29801);
xnor UO_720 (O_720,N_28800,N_28891);
nor UO_721 (O_721,N_28524,N_28626);
or UO_722 (O_722,N_29976,N_29501);
nor UO_723 (O_723,N_29443,N_28904);
nor UO_724 (O_724,N_28792,N_28882);
and UO_725 (O_725,N_29152,N_29397);
nor UO_726 (O_726,N_29668,N_29232);
nor UO_727 (O_727,N_28500,N_29677);
and UO_728 (O_728,N_29464,N_29449);
and UO_729 (O_729,N_29170,N_29513);
nor UO_730 (O_730,N_29372,N_29704);
xor UO_731 (O_731,N_29253,N_29641);
and UO_732 (O_732,N_29954,N_29250);
and UO_733 (O_733,N_29984,N_29259);
or UO_734 (O_734,N_29482,N_28872);
nor UO_735 (O_735,N_29489,N_28535);
xor UO_736 (O_736,N_28942,N_29104);
nor UO_737 (O_737,N_28977,N_29526);
nand UO_738 (O_738,N_28888,N_29706);
and UO_739 (O_739,N_28885,N_28654);
xnor UO_740 (O_740,N_29068,N_29323);
nand UO_741 (O_741,N_29696,N_28735);
and UO_742 (O_742,N_29895,N_28517);
nor UO_743 (O_743,N_29795,N_29227);
nor UO_744 (O_744,N_29918,N_29358);
or UO_745 (O_745,N_29479,N_29452);
nand UO_746 (O_746,N_29701,N_28549);
nor UO_747 (O_747,N_28786,N_29611);
or UO_748 (O_748,N_29603,N_28752);
and UO_749 (O_749,N_29444,N_29576);
xnor UO_750 (O_750,N_29102,N_29075);
nand UO_751 (O_751,N_29723,N_28819);
or UO_752 (O_752,N_29514,N_28798);
and UO_753 (O_753,N_29304,N_28638);
xor UO_754 (O_754,N_29686,N_29669);
and UO_755 (O_755,N_29004,N_29214);
xor UO_756 (O_756,N_28542,N_28755);
nand UO_757 (O_757,N_29187,N_29912);
or UO_758 (O_758,N_28755,N_28992);
xor UO_759 (O_759,N_28797,N_29050);
nand UO_760 (O_760,N_29028,N_28747);
nor UO_761 (O_761,N_29654,N_28593);
xnor UO_762 (O_762,N_29027,N_29855);
nand UO_763 (O_763,N_29656,N_28928);
or UO_764 (O_764,N_29923,N_29022);
or UO_765 (O_765,N_28776,N_29784);
nor UO_766 (O_766,N_28516,N_29338);
or UO_767 (O_767,N_29887,N_29106);
and UO_768 (O_768,N_29228,N_28808);
nand UO_769 (O_769,N_28879,N_29817);
xnor UO_770 (O_770,N_29156,N_29462);
nand UO_771 (O_771,N_28800,N_29361);
and UO_772 (O_772,N_28988,N_29704);
nand UO_773 (O_773,N_29982,N_28642);
or UO_774 (O_774,N_28529,N_28586);
nand UO_775 (O_775,N_29932,N_29195);
nand UO_776 (O_776,N_28936,N_29523);
nor UO_777 (O_777,N_28593,N_29504);
and UO_778 (O_778,N_29264,N_28543);
and UO_779 (O_779,N_28905,N_28989);
xnor UO_780 (O_780,N_29167,N_29836);
nor UO_781 (O_781,N_28921,N_29233);
nand UO_782 (O_782,N_29504,N_29040);
nor UO_783 (O_783,N_29329,N_29438);
nor UO_784 (O_784,N_29682,N_29077);
nor UO_785 (O_785,N_29569,N_28950);
or UO_786 (O_786,N_28751,N_28589);
or UO_787 (O_787,N_29462,N_29526);
or UO_788 (O_788,N_29408,N_29007);
or UO_789 (O_789,N_29282,N_29955);
nand UO_790 (O_790,N_28939,N_28776);
or UO_791 (O_791,N_28560,N_29587);
nand UO_792 (O_792,N_28841,N_29053);
xor UO_793 (O_793,N_29707,N_29355);
nor UO_794 (O_794,N_28608,N_29405);
and UO_795 (O_795,N_29077,N_29944);
nand UO_796 (O_796,N_28905,N_29519);
nand UO_797 (O_797,N_29674,N_28606);
and UO_798 (O_798,N_29963,N_29365);
nand UO_799 (O_799,N_28553,N_29713);
nand UO_800 (O_800,N_28903,N_29773);
nand UO_801 (O_801,N_28519,N_29022);
and UO_802 (O_802,N_28704,N_29251);
nor UO_803 (O_803,N_29479,N_28746);
or UO_804 (O_804,N_28682,N_29828);
xnor UO_805 (O_805,N_29683,N_29851);
and UO_806 (O_806,N_28566,N_28998);
nand UO_807 (O_807,N_29769,N_29303);
or UO_808 (O_808,N_28765,N_29663);
xor UO_809 (O_809,N_29701,N_29151);
xnor UO_810 (O_810,N_28665,N_29157);
nand UO_811 (O_811,N_29306,N_29591);
and UO_812 (O_812,N_28752,N_29428);
xnor UO_813 (O_813,N_28662,N_29708);
nand UO_814 (O_814,N_29281,N_29474);
nor UO_815 (O_815,N_29573,N_28508);
xor UO_816 (O_816,N_29387,N_28572);
or UO_817 (O_817,N_29178,N_29886);
nor UO_818 (O_818,N_29340,N_28606);
nand UO_819 (O_819,N_29858,N_29705);
and UO_820 (O_820,N_28709,N_29523);
and UO_821 (O_821,N_29220,N_29080);
xor UO_822 (O_822,N_28939,N_29890);
and UO_823 (O_823,N_28624,N_29578);
nand UO_824 (O_824,N_29218,N_29236);
xnor UO_825 (O_825,N_29846,N_29911);
nand UO_826 (O_826,N_28618,N_28681);
xnor UO_827 (O_827,N_29340,N_29140);
nand UO_828 (O_828,N_28566,N_29885);
and UO_829 (O_829,N_29753,N_28693);
nand UO_830 (O_830,N_29554,N_29643);
nor UO_831 (O_831,N_29594,N_28622);
or UO_832 (O_832,N_29237,N_29927);
nand UO_833 (O_833,N_28538,N_29272);
or UO_834 (O_834,N_29034,N_28946);
nand UO_835 (O_835,N_29152,N_28523);
nor UO_836 (O_836,N_28789,N_29332);
xor UO_837 (O_837,N_28696,N_29239);
or UO_838 (O_838,N_28622,N_28973);
nand UO_839 (O_839,N_28677,N_29923);
or UO_840 (O_840,N_28697,N_29001);
nor UO_841 (O_841,N_29194,N_29212);
nor UO_842 (O_842,N_29254,N_28999);
xnor UO_843 (O_843,N_29011,N_29650);
xnor UO_844 (O_844,N_29278,N_29545);
and UO_845 (O_845,N_29221,N_29223);
nor UO_846 (O_846,N_28731,N_29938);
nor UO_847 (O_847,N_29748,N_29959);
nor UO_848 (O_848,N_28755,N_28715);
or UO_849 (O_849,N_28675,N_29057);
nand UO_850 (O_850,N_29838,N_28739);
nand UO_851 (O_851,N_29456,N_29431);
nand UO_852 (O_852,N_29181,N_28669);
and UO_853 (O_853,N_28713,N_29249);
or UO_854 (O_854,N_29501,N_29582);
nor UO_855 (O_855,N_28789,N_29305);
and UO_856 (O_856,N_28934,N_29951);
xnor UO_857 (O_857,N_29184,N_29882);
xnor UO_858 (O_858,N_29932,N_28608);
and UO_859 (O_859,N_29493,N_28595);
nand UO_860 (O_860,N_28889,N_29529);
or UO_861 (O_861,N_29004,N_28594);
or UO_862 (O_862,N_29957,N_28797);
xor UO_863 (O_863,N_29234,N_28663);
xnor UO_864 (O_864,N_29637,N_29493);
nor UO_865 (O_865,N_29216,N_29265);
nor UO_866 (O_866,N_29873,N_28574);
or UO_867 (O_867,N_28801,N_28766);
xnor UO_868 (O_868,N_29662,N_28882);
nand UO_869 (O_869,N_29268,N_29749);
nand UO_870 (O_870,N_29264,N_29580);
xnor UO_871 (O_871,N_28557,N_29912);
xor UO_872 (O_872,N_29350,N_28844);
and UO_873 (O_873,N_29953,N_29673);
or UO_874 (O_874,N_28599,N_29850);
xor UO_875 (O_875,N_29969,N_29173);
nand UO_876 (O_876,N_29744,N_29854);
xor UO_877 (O_877,N_28630,N_28679);
nor UO_878 (O_878,N_28593,N_29028);
nor UO_879 (O_879,N_28582,N_29273);
xnor UO_880 (O_880,N_29716,N_28649);
xor UO_881 (O_881,N_28743,N_29576);
and UO_882 (O_882,N_29626,N_29112);
xor UO_883 (O_883,N_28961,N_28927);
xnor UO_884 (O_884,N_29619,N_29791);
nor UO_885 (O_885,N_29883,N_29553);
nand UO_886 (O_886,N_29619,N_28957);
or UO_887 (O_887,N_29190,N_28956);
nand UO_888 (O_888,N_28841,N_29984);
nand UO_889 (O_889,N_29586,N_28612);
xor UO_890 (O_890,N_28856,N_29639);
or UO_891 (O_891,N_29631,N_29142);
xor UO_892 (O_892,N_29651,N_29667);
and UO_893 (O_893,N_29926,N_29881);
nor UO_894 (O_894,N_29898,N_29058);
or UO_895 (O_895,N_29351,N_28758);
nor UO_896 (O_896,N_29072,N_28653);
nor UO_897 (O_897,N_28537,N_29293);
xor UO_898 (O_898,N_29032,N_29149);
xor UO_899 (O_899,N_29069,N_29820);
and UO_900 (O_900,N_29094,N_28683);
xnor UO_901 (O_901,N_29390,N_29253);
and UO_902 (O_902,N_29544,N_29137);
nand UO_903 (O_903,N_28616,N_28765);
and UO_904 (O_904,N_29572,N_29180);
xor UO_905 (O_905,N_29055,N_28914);
xor UO_906 (O_906,N_28740,N_29323);
nor UO_907 (O_907,N_28707,N_29541);
nor UO_908 (O_908,N_29973,N_29794);
nor UO_909 (O_909,N_29130,N_29006);
or UO_910 (O_910,N_29350,N_29386);
xor UO_911 (O_911,N_29121,N_29630);
or UO_912 (O_912,N_29598,N_29959);
or UO_913 (O_913,N_29062,N_28682);
or UO_914 (O_914,N_29295,N_29141);
nor UO_915 (O_915,N_29062,N_29771);
or UO_916 (O_916,N_29218,N_28515);
or UO_917 (O_917,N_29683,N_28503);
or UO_918 (O_918,N_28646,N_29018);
and UO_919 (O_919,N_29242,N_28685);
nor UO_920 (O_920,N_28586,N_29641);
xor UO_921 (O_921,N_28855,N_29680);
and UO_922 (O_922,N_28655,N_29512);
and UO_923 (O_923,N_29284,N_29007);
xor UO_924 (O_924,N_28523,N_28936);
nand UO_925 (O_925,N_28841,N_28697);
and UO_926 (O_926,N_29151,N_29363);
nor UO_927 (O_927,N_29832,N_28855);
and UO_928 (O_928,N_29944,N_29161);
nand UO_929 (O_929,N_28994,N_29944);
and UO_930 (O_930,N_28714,N_29915);
or UO_931 (O_931,N_28749,N_29835);
xnor UO_932 (O_932,N_29732,N_28944);
nor UO_933 (O_933,N_29124,N_28571);
nor UO_934 (O_934,N_28949,N_28826);
or UO_935 (O_935,N_28952,N_28807);
or UO_936 (O_936,N_29930,N_29527);
xor UO_937 (O_937,N_28514,N_29466);
nor UO_938 (O_938,N_28764,N_29300);
nor UO_939 (O_939,N_29216,N_29304);
xor UO_940 (O_940,N_29148,N_29193);
nand UO_941 (O_941,N_28667,N_29956);
or UO_942 (O_942,N_28540,N_28860);
nor UO_943 (O_943,N_29444,N_29309);
or UO_944 (O_944,N_28645,N_29812);
nand UO_945 (O_945,N_29651,N_29622);
or UO_946 (O_946,N_29939,N_29550);
nand UO_947 (O_947,N_29953,N_29244);
nand UO_948 (O_948,N_28781,N_29823);
nand UO_949 (O_949,N_29051,N_28969);
xor UO_950 (O_950,N_28853,N_29218);
nand UO_951 (O_951,N_29853,N_29598);
or UO_952 (O_952,N_29636,N_29956);
nand UO_953 (O_953,N_28704,N_29701);
xnor UO_954 (O_954,N_28811,N_28658);
xor UO_955 (O_955,N_29475,N_28566);
and UO_956 (O_956,N_28979,N_29458);
xnor UO_957 (O_957,N_28728,N_29073);
nand UO_958 (O_958,N_29064,N_28603);
xnor UO_959 (O_959,N_28979,N_29351);
and UO_960 (O_960,N_29836,N_28562);
xor UO_961 (O_961,N_28631,N_29128);
or UO_962 (O_962,N_29764,N_28979);
nor UO_963 (O_963,N_28861,N_29880);
or UO_964 (O_964,N_29060,N_28657);
nor UO_965 (O_965,N_29726,N_28688);
nand UO_966 (O_966,N_28971,N_28611);
or UO_967 (O_967,N_29953,N_29162);
nor UO_968 (O_968,N_28870,N_29627);
or UO_969 (O_969,N_28749,N_29066);
nand UO_970 (O_970,N_29891,N_29695);
nand UO_971 (O_971,N_28831,N_29277);
nand UO_972 (O_972,N_29879,N_29083);
nor UO_973 (O_973,N_28778,N_29700);
nand UO_974 (O_974,N_29085,N_29506);
xor UO_975 (O_975,N_28546,N_29549);
or UO_976 (O_976,N_29432,N_29075);
and UO_977 (O_977,N_29721,N_29208);
or UO_978 (O_978,N_29513,N_28759);
xnor UO_979 (O_979,N_28564,N_29842);
nand UO_980 (O_980,N_28663,N_28841);
xnor UO_981 (O_981,N_29624,N_28678);
and UO_982 (O_982,N_29109,N_29023);
nor UO_983 (O_983,N_29523,N_28966);
and UO_984 (O_984,N_29548,N_28643);
nand UO_985 (O_985,N_29340,N_29774);
or UO_986 (O_986,N_28987,N_28695);
xor UO_987 (O_987,N_29331,N_29218);
nand UO_988 (O_988,N_29700,N_28961);
xnor UO_989 (O_989,N_28764,N_29930);
and UO_990 (O_990,N_29226,N_28557);
and UO_991 (O_991,N_29950,N_29493);
and UO_992 (O_992,N_29535,N_29860);
and UO_993 (O_993,N_29760,N_29482);
nand UO_994 (O_994,N_28541,N_28548);
and UO_995 (O_995,N_29778,N_29765);
and UO_996 (O_996,N_29749,N_29083);
nor UO_997 (O_997,N_29125,N_29900);
or UO_998 (O_998,N_29586,N_29018);
nor UO_999 (O_999,N_28578,N_28581);
nand UO_1000 (O_1000,N_29781,N_29830);
or UO_1001 (O_1001,N_29510,N_29005);
or UO_1002 (O_1002,N_29618,N_28783);
nand UO_1003 (O_1003,N_29150,N_28905);
nand UO_1004 (O_1004,N_29053,N_28686);
or UO_1005 (O_1005,N_29306,N_28509);
xor UO_1006 (O_1006,N_29677,N_29768);
nor UO_1007 (O_1007,N_28744,N_29455);
xnor UO_1008 (O_1008,N_29159,N_29643);
nand UO_1009 (O_1009,N_28503,N_29687);
xor UO_1010 (O_1010,N_29583,N_28658);
xnor UO_1011 (O_1011,N_29820,N_28585);
nor UO_1012 (O_1012,N_28828,N_29507);
and UO_1013 (O_1013,N_28665,N_29556);
xor UO_1014 (O_1014,N_29231,N_29814);
nand UO_1015 (O_1015,N_28974,N_28849);
nor UO_1016 (O_1016,N_28979,N_29031);
and UO_1017 (O_1017,N_29122,N_29264);
nor UO_1018 (O_1018,N_29415,N_29312);
nand UO_1019 (O_1019,N_29623,N_29639);
nand UO_1020 (O_1020,N_28627,N_29271);
nor UO_1021 (O_1021,N_28707,N_29835);
and UO_1022 (O_1022,N_29988,N_29404);
or UO_1023 (O_1023,N_29706,N_28539);
xnor UO_1024 (O_1024,N_29059,N_29995);
nand UO_1025 (O_1025,N_29299,N_28794);
nand UO_1026 (O_1026,N_29433,N_29498);
nor UO_1027 (O_1027,N_29508,N_29715);
xor UO_1028 (O_1028,N_28825,N_29874);
nand UO_1029 (O_1029,N_28536,N_29336);
nor UO_1030 (O_1030,N_29830,N_29881);
or UO_1031 (O_1031,N_28629,N_29507);
nor UO_1032 (O_1032,N_29092,N_29875);
or UO_1033 (O_1033,N_28956,N_28589);
nor UO_1034 (O_1034,N_29619,N_28838);
xor UO_1035 (O_1035,N_29752,N_29320);
xnor UO_1036 (O_1036,N_29486,N_29884);
or UO_1037 (O_1037,N_28943,N_28923);
and UO_1038 (O_1038,N_28531,N_29875);
nand UO_1039 (O_1039,N_29433,N_29806);
or UO_1040 (O_1040,N_29416,N_29240);
nor UO_1041 (O_1041,N_29488,N_28935);
and UO_1042 (O_1042,N_28673,N_28765);
nand UO_1043 (O_1043,N_29365,N_28906);
xnor UO_1044 (O_1044,N_29085,N_28916);
nand UO_1045 (O_1045,N_28514,N_29046);
nand UO_1046 (O_1046,N_29427,N_29477);
and UO_1047 (O_1047,N_29780,N_29845);
nand UO_1048 (O_1048,N_29410,N_28865);
xor UO_1049 (O_1049,N_29504,N_29462);
xnor UO_1050 (O_1050,N_29867,N_29566);
and UO_1051 (O_1051,N_28514,N_28925);
nand UO_1052 (O_1052,N_29664,N_29435);
nand UO_1053 (O_1053,N_29718,N_28968);
or UO_1054 (O_1054,N_28610,N_29344);
or UO_1055 (O_1055,N_28906,N_29631);
or UO_1056 (O_1056,N_29031,N_28680);
xnor UO_1057 (O_1057,N_29648,N_29275);
nand UO_1058 (O_1058,N_28685,N_28570);
xor UO_1059 (O_1059,N_29397,N_28829);
nand UO_1060 (O_1060,N_28701,N_29034);
and UO_1061 (O_1061,N_29749,N_29734);
nor UO_1062 (O_1062,N_29439,N_29792);
or UO_1063 (O_1063,N_29434,N_29633);
nand UO_1064 (O_1064,N_28722,N_28676);
nand UO_1065 (O_1065,N_29402,N_29397);
nand UO_1066 (O_1066,N_29736,N_29475);
and UO_1067 (O_1067,N_28869,N_29299);
nand UO_1068 (O_1068,N_29887,N_28820);
xor UO_1069 (O_1069,N_29702,N_29768);
nor UO_1070 (O_1070,N_28712,N_28976);
nand UO_1071 (O_1071,N_29027,N_28528);
xnor UO_1072 (O_1072,N_29652,N_29274);
nor UO_1073 (O_1073,N_29922,N_28730);
nand UO_1074 (O_1074,N_29151,N_29689);
nor UO_1075 (O_1075,N_29699,N_28763);
or UO_1076 (O_1076,N_29069,N_28886);
nand UO_1077 (O_1077,N_28801,N_29001);
nor UO_1078 (O_1078,N_28555,N_29165);
or UO_1079 (O_1079,N_29360,N_29277);
nor UO_1080 (O_1080,N_29749,N_28657);
nor UO_1081 (O_1081,N_29102,N_29781);
nor UO_1082 (O_1082,N_29363,N_29411);
xnor UO_1083 (O_1083,N_29795,N_29760);
or UO_1084 (O_1084,N_29966,N_29111);
nand UO_1085 (O_1085,N_28525,N_28554);
and UO_1086 (O_1086,N_29384,N_28842);
or UO_1087 (O_1087,N_29815,N_28942);
nand UO_1088 (O_1088,N_29825,N_29667);
or UO_1089 (O_1089,N_28651,N_29865);
or UO_1090 (O_1090,N_28602,N_28705);
xnor UO_1091 (O_1091,N_29212,N_29803);
nor UO_1092 (O_1092,N_29340,N_29263);
and UO_1093 (O_1093,N_29433,N_28581);
or UO_1094 (O_1094,N_28995,N_28629);
nand UO_1095 (O_1095,N_29611,N_29467);
nor UO_1096 (O_1096,N_29865,N_28762);
or UO_1097 (O_1097,N_29624,N_29691);
nand UO_1098 (O_1098,N_29568,N_29141);
and UO_1099 (O_1099,N_29470,N_28554);
and UO_1100 (O_1100,N_28766,N_28940);
xnor UO_1101 (O_1101,N_29334,N_29949);
or UO_1102 (O_1102,N_28848,N_29124);
or UO_1103 (O_1103,N_29432,N_28962);
nand UO_1104 (O_1104,N_28748,N_28782);
or UO_1105 (O_1105,N_29894,N_28804);
nand UO_1106 (O_1106,N_29779,N_29759);
xor UO_1107 (O_1107,N_29379,N_29843);
or UO_1108 (O_1108,N_29266,N_29771);
nand UO_1109 (O_1109,N_28720,N_29920);
xor UO_1110 (O_1110,N_29080,N_29087);
or UO_1111 (O_1111,N_29069,N_29013);
xor UO_1112 (O_1112,N_29213,N_28787);
xor UO_1113 (O_1113,N_29726,N_28981);
and UO_1114 (O_1114,N_29810,N_29220);
or UO_1115 (O_1115,N_29896,N_28968);
nand UO_1116 (O_1116,N_29741,N_29272);
and UO_1117 (O_1117,N_28621,N_28605);
xnor UO_1118 (O_1118,N_29512,N_28667);
and UO_1119 (O_1119,N_29617,N_29937);
and UO_1120 (O_1120,N_28756,N_29037);
nand UO_1121 (O_1121,N_29664,N_29959);
xnor UO_1122 (O_1122,N_28949,N_29000);
nor UO_1123 (O_1123,N_28527,N_28733);
nor UO_1124 (O_1124,N_29807,N_29057);
and UO_1125 (O_1125,N_29151,N_29774);
and UO_1126 (O_1126,N_29164,N_28959);
or UO_1127 (O_1127,N_28674,N_29109);
and UO_1128 (O_1128,N_28556,N_29727);
xnor UO_1129 (O_1129,N_29735,N_29378);
nor UO_1130 (O_1130,N_28545,N_28585);
xnor UO_1131 (O_1131,N_29948,N_28785);
nor UO_1132 (O_1132,N_29175,N_29520);
or UO_1133 (O_1133,N_28969,N_29711);
and UO_1134 (O_1134,N_29466,N_29849);
xor UO_1135 (O_1135,N_28963,N_28828);
or UO_1136 (O_1136,N_28633,N_28739);
or UO_1137 (O_1137,N_29294,N_29989);
or UO_1138 (O_1138,N_29992,N_28780);
and UO_1139 (O_1139,N_28822,N_29944);
nand UO_1140 (O_1140,N_29341,N_28662);
and UO_1141 (O_1141,N_29232,N_29868);
nand UO_1142 (O_1142,N_29350,N_29244);
and UO_1143 (O_1143,N_29100,N_29009);
xor UO_1144 (O_1144,N_28846,N_29162);
nand UO_1145 (O_1145,N_29479,N_29781);
nand UO_1146 (O_1146,N_29690,N_29710);
xor UO_1147 (O_1147,N_29350,N_29801);
and UO_1148 (O_1148,N_28922,N_29610);
xor UO_1149 (O_1149,N_28880,N_28579);
xor UO_1150 (O_1150,N_29906,N_28727);
nand UO_1151 (O_1151,N_29447,N_28551);
and UO_1152 (O_1152,N_29947,N_29961);
nand UO_1153 (O_1153,N_28587,N_28618);
or UO_1154 (O_1154,N_29235,N_28634);
and UO_1155 (O_1155,N_29257,N_28784);
nand UO_1156 (O_1156,N_28685,N_28504);
xnor UO_1157 (O_1157,N_29978,N_28936);
nand UO_1158 (O_1158,N_29853,N_29566);
or UO_1159 (O_1159,N_29262,N_28987);
and UO_1160 (O_1160,N_29851,N_29534);
or UO_1161 (O_1161,N_29225,N_29175);
nor UO_1162 (O_1162,N_29183,N_29863);
or UO_1163 (O_1163,N_28549,N_29200);
xnor UO_1164 (O_1164,N_29937,N_29269);
and UO_1165 (O_1165,N_29344,N_29010);
and UO_1166 (O_1166,N_29387,N_28685);
or UO_1167 (O_1167,N_28584,N_29045);
nor UO_1168 (O_1168,N_29927,N_29247);
and UO_1169 (O_1169,N_29060,N_28583);
xnor UO_1170 (O_1170,N_29084,N_28624);
and UO_1171 (O_1171,N_29336,N_29062);
nand UO_1172 (O_1172,N_28588,N_28596);
and UO_1173 (O_1173,N_28829,N_29655);
and UO_1174 (O_1174,N_29296,N_28952);
xor UO_1175 (O_1175,N_29352,N_28571);
nor UO_1176 (O_1176,N_29660,N_29489);
nor UO_1177 (O_1177,N_29534,N_28816);
and UO_1178 (O_1178,N_28798,N_29312);
xnor UO_1179 (O_1179,N_29914,N_29335);
xnor UO_1180 (O_1180,N_29860,N_29972);
xnor UO_1181 (O_1181,N_29645,N_29963);
nand UO_1182 (O_1182,N_29411,N_29050);
xor UO_1183 (O_1183,N_29294,N_28866);
or UO_1184 (O_1184,N_28863,N_28747);
nor UO_1185 (O_1185,N_29060,N_29187);
nand UO_1186 (O_1186,N_28795,N_29685);
or UO_1187 (O_1187,N_29713,N_28996);
nor UO_1188 (O_1188,N_28709,N_29100);
nand UO_1189 (O_1189,N_28759,N_29333);
nor UO_1190 (O_1190,N_29539,N_29588);
xor UO_1191 (O_1191,N_29577,N_28873);
nor UO_1192 (O_1192,N_29592,N_28644);
nor UO_1193 (O_1193,N_29908,N_28620);
and UO_1194 (O_1194,N_28857,N_28767);
and UO_1195 (O_1195,N_28682,N_29429);
nor UO_1196 (O_1196,N_29404,N_29614);
nand UO_1197 (O_1197,N_28554,N_29337);
and UO_1198 (O_1198,N_28685,N_28828);
nor UO_1199 (O_1199,N_28930,N_29021);
and UO_1200 (O_1200,N_28969,N_29085);
xnor UO_1201 (O_1201,N_28605,N_29578);
nor UO_1202 (O_1202,N_29948,N_29008);
xnor UO_1203 (O_1203,N_28761,N_28959);
nor UO_1204 (O_1204,N_28548,N_29672);
xnor UO_1205 (O_1205,N_28570,N_29850);
nand UO_1206 (O_1206,N_28784,N_29521);
nand UO_1207 (O_1207,N_29244,N_29973);
nor UO_1208 (O_1208,N_28971,N_28902);
or UO_1209 (O_1209,N_28797,N_29902);
nand UO_1210 (O_1210,N_29210,N_29499);
or UO_1211 (O_1211,N_29530,N_29086);
nor UO_1212 (O_1212,N_28799,N_28601);
or UO_1213 (O_1213,N_29269,N_29157);
or UO_1214 (O_1214,N_28844,N_29792);
nor UO_1215 (O_1215,N_29326,N_29746);
or UO_1216 (O_1216,N_28827,N_28881);
and UO_1217 (O_1217,N_29803,N_29266);
xor UO_1218 (O_1218,N_29753,N_28749);
nand UO_1219 (O_1219,N_29400,N_28856);
nand UO_1220 (O_1220,N_29400,N_29421);
or UO_1221 (O_1221,N_28566,N_29086);
or UO_1222 (O_1222,N_28718,N_29224);
nand UO_1223 (O_1223,N_29990,N_28668);
and UO_1224 (O_1224,N_29374,N_29416);
or UO_1225 (O_1225,N_29222,N_29865);
xnor UO_1226 (O_1226,N_28695,N_28773);
xor UO_1227 (O_1227,N_29139,N_28555);
nor UO_1228 (O_1228,N_28705,N_29112);
nand UO_1229 (O_1229,N_29320,N_29078);
or UO_1230 (O_1230,N_29561,N_28602);
xnor UO_1231 (O_1231,N_29076,N_29348);
nor UO_1232 (O_1232,N_29708,N_29599);
or UO_1233 (O_1233,N_29335,N_28575);
and UO_1234 (O_1234,N_29298,N_29320);
or UO_1235 (O_1235,N_29464,N_28642);
nor UO_1236 (O_1236,N_29268,N_28969);
and UO_1237 (O_1237,N_29514,N_29713);
xor UO_1238 (O_1238,N_29713,N_29417);
xnor UO_1239 (O_1239,N_29518,N_29443);
nand UO_1240 (O_1240,N_29730,N_29534);
and UO_1241 (O_1241,N_29464,N_28683);
xor UO_1242 (O_1242,N_29536,N_28631);
and UO_1243 (O_1243,N_29256,N_28689);
or UO_1244 (O_1244,N_28803,N_29888);
and UO_1245 (O_1245,N_29084,N_28849);
and UO_1246 (O_1246,N_29489,N_28987);
or UO_1247 (O_1247,N_29136,N_28950);
or UO_1248 (O_1248,N_28949,N_29156);
and UO_1249 (O_1249,N_29950,N_29420);
nor UO_1250 (O_1250,N_28541,N_28868);
or UO_1251 (O_1251,N_29794,N_29575);
nand UO_1252 (O_1252,N_28607,N_29503);
and UO_1253 (O_1253,N_28539,N_28516);
xor UO_1254 (O_1254,N_28543,N_29483);
nand UO_1255 (O_1255,N_28778,N_29403);
nor UO_1256 (O_1256,N_29417,N_29839);
nand UO_1257 (O_1257,N_28952,N_29014);
xor UO_1258 (O_1258,N_29900,N_29467);
xnor UO_1259 (O_1259,N_28513,N_29634);
nand UO_1260 (O_1260,N_29046,N_29556);
nand UO_1261 (O_1261,N_29324,N_28587);
or UO_1262 (O_1262,N_29135,N_29042);
nand UO_1263 (O_1263,N_29666,N_29296);
and UO_1264 (O_1264,N_29712,N_29485);
or UO_1265 (O_1265,N_28967,N_29648);
xor UO_1266 (O_1266,N_28607,N_29091);
nand UO_1267 (O_1267,N_29388,N_28993);
nor UO_1268 (O_1268,N_29474,N_29396);
nor UO_1269 (O_1269,N_29910,N_29700);
xnor UO_1270 (O_1270,N_29116,N_29907);
or UO_1271 (O_1271,N_28635,N_29715);
or UO_1272 (O_1272,N_28991,N_28716);
and UO_1273 (O_1273,N_29574,N_29669);
nand UO_1274 (O_1274,N_29696,N_29558);
nand UO_1275 (O_1275,N_29982,N_29762);
xor UO_1276 (O_1276,N_28734,N_29457);
and UO_1277 (O_1277,N_29145,N_28647);
nor UO_1278 (O_1278,N_29012,N_29183);
or UO_1279 (O_1279,N_28539,N_29772);
nand UO_1280 (O_1280,N_29607,N_28772);
nor UO_1281 (O_1281,N_29512,N_28962);
and UO_1282 (O_1282,N_29672,N_29816);
or UO_1283 (O_1283,N_29162,N_29675);
xnor UO_1284 (O_1284,N_29550,N_29136);
and UO_1285 (O_1285,N_29253,N_29098);
or UO_1286 (O_1286,N_28603,N_29215);
nand UO_1287 (O_1287,N_29575,N_29048);
nand UO_1288 (O_1288,N_28682,N_29838);
or UO_1289 (O_1289,N_29521,N_29806);
nor UO_1290 (O_1290,N_28923,N_28648);
nor UO_1291 (O_1291,N_29630,N_29042);
nor UO_1292 (O_1292,N_28611,N_28746);
nor UO_1293 (O_1293,N_29179,N_29058);
or UO_1294 (O_1294,N_28592,N_28990);
xor UO_1295 (O_1295,N_29914,N_28721);
nor UO_1296 (O_1296,N_29368,N_29761);
and UO_1297 (O_1297,N_28574,N_28752);
nor UO_1298 (O_1298,N_29648,N_28517);
xnor UO_1299 (O_1299,N_28682,N_28522);
or UO_1300 (O_1300,N_29782,N_28830);
and UO_1301 (O_1301,N_29235,N_29246);
nor UO_1302 (O_1302,N_29043,N_28536);
nand UO_1303 (O_1303,N_29890,N_28614);
and UO_1304 (O_1304,N_29287,N_29952);
or UO_1305 (O_1305,N_29819,N_29937);
and UO_1306 (O_1306,N_29225,N_29641);
or UO_1307 (O_1307,N_29529,N_29646);
xor UO_1308 (O_1308,N_29399,N_29300);
xnor UO_1309 (O_1309,N_29842,N_29686);
nor UO_1310 (O_1310,N_28990,N_28856);
nand UO_1311 (O_1311,N_29658,N_28915);
nor UO_1312 (O_1312,N_29752,N_29960);
nand UO_1313 (O_1313,N_28544,N_28745);
nand UO_1314 (O_1314,N_29713,N_29820);
nor UO_1315 (O_1315,N_28550,N_29888);
nand UO_1316 (O_1316,N_29234,N_28961);
or UO_1317 (O_1317,N_28688,N_28718);
and UO_1318 (O_1318,N_29893,N_29743);
nor UO_1319 (O_1319,N_28998,N_29555);
xnor UO_1320 (O_1320,N_29258,N_28897);
nor UO_1321 (O_1321,N_29517,N_28656);
nor UO_1322 (O_1322,N_28562,N_29692);
and UO_1323 (O_1323,N_29342,N_28900);
xor UO_1324 (O_1324,N_28980,N_29746);
nand UO_1325 (O_1325,N_29934,N_29541);
xnor UO_1326 (O_1326,N_29569,N_29934);
or UO_1327 (O_1327,N_28666,N_28981);
nor UO_1328 (O_1328,N_29870,N_29276);
or UO_1329 (O_1329,N_29050,N_29974);
nor UO_1330 (O_1330,N_29955,N_29078);
and UO_1331 (O_1331,N_28896,N_28958);
nor UO_1332 (O_1332,N_28995,N_29361);
or UO_1333 (O_1333,N_29305,N_28792);
xnor UO_1334 (O_1334,N_28963,N_29815);
xnor UO_1335 (O_1335,N_28996,N_29704);
and UO_1336 (O_1336,N_29009,N_28744);
or UO_1337 (O_1337,N_29057,N_29549);
or UO_1338 (O_1338,N_29399,N_28809);
nand UO_1339 (O_1339,N_29030,N_29871);
or UO_1340 (O_1340,N_28665,N_29421);
nand UO_1341 (O_1341,N_28820,N_28942);
nand UO_1342 (O_1342,N_29122,N_29705);
xnor UO_1343 (O_1343,N_29165,N_28545);
and UO_1344 (O_1344,N_29438,N_29374);
xor UO_1345 (O_1345,N_29209,N_29668);
nand UO_1346 (O_1346,N_29014,N_29998);
nand UO_1347 (O_1347,N_29389,N_29993);
xnor UO_1348 (O_1348,N_29432,N_29552);
xnor UO_1349 (O_1349,N_29177,N_29610);
nor UO_1350 (O_1350,N_29448,N_29630);
nor UO_1351 (O_1351,N_29780,N_29118);
or UO_1352 (O_1352,N_28854,N_29309);
xor UO_1353 (O_1353,N_29904,N_28717);
nor UO_1354 (O_1354,N_29996,N_28781);
and UO_1355 (O_1355,N_28952,N_29236);
nor UO_1356 (O_1356,N_29387,N_29704);
nor UO_1357 (O_1357,N_28808,N_28633);
or UO_1358 (O_1358,N_29469,N_29289);
nand UO_1359 (O_1359,N_28924,N_29918);
and UO_1360 (O_1360,N_28894,N_29213);
nand UO_1361 (O_1361,N_29394,N_28558);
nand UO_1362 (O_1362,N_29130,N_29591);
and UO_1363 (O_1363,N_29052,N_28893);
and UO_1364 (O_1364,N_29418,N_28897);
xor UO_1365 (O_1365,N_29719,N_29288);
and UO_1366 (O_1366,N_29097,N_29354);
xor UO_1367 (O_1367,N_29325,N_28853);
or UO_1368 (O_1368,N_29016,N_29082);
nor UO_1369 (O_1369,N_29962,N_28740);
or UO_1370 (O_1370,N_28818,N_28821);
or UO_1371 (O_1371,N_29428,N_29189);
or UO_1372 (O_1372,N_29887,N_29359);
nor UO_1373 (O_1373,N_29343,N_28823);
and UO_1374 (O_1374,N_29671,N_29708);
nand UO_1375 (O_1375,N_29775,N_29203);
nor UO_1376 (O_1376,N_29963,N_29862);
nand UO_1377 (O_1377,N_29318,N_29520);
nand UO_1378 (O_1378,N_29398,N_29626);
or UO_1379 (O_1379,N_28625,N_28997);
nand UO_1380 (O_1380,N_28719,N_28798);
or UO_1381 (O_1381,N_29478,N_29102);
nor UO_1382 (O_1382,N_29476,N_29226);
or UO_1383 (O_1383,N_29888,N_28798);
xnor UO_1384 (O_1384,N_28722,N_28732);
and UO_1385 (O_1385,N_28805,N_29026);
nor UO_1386 (O_1386,N_29136,N_29656);
nand UO_1387 (O_1387,N_29993,N_29202);
xor UO_1388 (O_1388,N_28913,N_28524);
nand UO_1389 (O_1389,N_28505,N_28948);
or UO_1390 (O_1390,N_29875,N_28810);
and UO_1391 (O_1391,N_29058,N_29733);
xor UO_1392 (O_1392,N_29059,N_29280);
or UO_1393 (O_1393,N_29782,N_29063);
nor UO_1394 (O_1394,N_29418,N_28738);
nor UO_1395 (O_1395,N_29967,N_29541);
nand UO_1396 (O_1396,N_28519,N_29695);
xor UO_1397 (O_1397,N_29223,N_29258);
and UO_1398 (O_1398,N_29918,N_28563);
nor UO_1399 (O_1399,N_29002,N_29063);
and UO_1400 (O_1400,N_28663,N_29512);
nor UO_1401 (O_1401,N_29975,N_29299);
and UO_1402 (O_1402,N_29177,N_29950);
xor UO_1403 (O_1403,N_29806,N_28543);
nand UO_1404 (O_1404,N_29043,N_29100);
and UO_1405 (O_1405,N_28878,N_29442);
xnor UO_1406 (O_1406,N_28577,N_29886);
or UO_1407 (O_1407,N_29243,N_29228);
nor UO_1408 (O_1408,N_29780,N_29161);
nor UO_1409 (O_1409,N_28976,N_29626);
or UO_1410 (O_1410,N_28981,N_28619);
or UO_1411 (O_1411,N_28599,N_28733);
or UO_1412 (O_1412,N_28941,N_29765);
nor UO_1413 (O_1413,N_29513,N_28934);
nor UO_1414 (O_1414,N_29464,N_28836);
nor UO_1415 (O_1415,N_28588,N_29137);
and UO_1416 (O_1416,N_28943,N_29961);
or UO_1417 (O_1417,N_29083,N_29956);
and UO_1418 (O_1418,N_29793,N_29513);
nand UO_1419 (O_1419,N_29612,N_29010);
or UO_1420 (O_1420,N_28517,N_28812);
nand UO_1421 (O_1421,N_29807,N_29602);
and UO_1422 (O_1422,N_28853,N_28711);
nor UO_1423 (O_1423,N_29370,N_28802);
or UO_1424 (O_1424,N_29524,N_29230);
nor UO_1425 (O_1425,N_29780,N_29732);
nand UO_1426 (O_1426,N_29948,N_28857);
or UO_1427 (O_1427,N_29805,N_29763);
nand UO_1428 (O_1428,N_29938,N_29227);
and UO_1429 (O_1429,N_29021,N_29430);
xor UO_1430 (O_1430,N_29833,N_29010);
nand UO_1431 (O_1431,N_29441,N_28628);
xnor UO_1432 (O_1432,N_29483,N_29745);
nand UO_1433 (O_1433,N_29067,N_28707);
and UO_1434 (O_1434,N_29735,N_29335);
or UO_1435 (O_1435,N_29305,N_28685);
nand UO_1436 (O_1436,N_28914,N_28521);
xor UO_1437 (O_1437,N_28731,N_29651);
or UO_1438 (O_1438,N_29455,N_29280);
xnor UO_1439 (O_1439,N_28777,N_29529);
xor UO_1440 (O_1440,N_29395,N_29701);
nand UO_1441 (O_1441,N_28752,N_28622);
nor UO_1442 (O_1442,N_29751,N_28927);
or UO_1443 (O_1443,N_29363,N_28500);
xor UO_1444 (O_1444,N_29277,N_28970);
nor UO_1445 (O_1445,N_28631,N_28893);
nor UO_1446 (O_1446,N_29275,N_28758);
xnor UO_1447 (O_1447,N_28585,N_29433);
xnor UO_1448 (O_1448,N_28823,N_28538);
nand UO_1449 (O_1449,N_29248,N_29226);
and UO_1450 (O_1450,N_29333,N_29420);
and UO_1451 (O_1451,N_28983,N_29828);
xnor UO_1452 (O_1452,N_29971,N_29452);
nor UO_1453 (O_1453,N_29903,N_29928);
or UO_1454 (O_1454,N_28651,N_29049);
xnor UO_1455 (O_1455,N_29948,N_28563);
nor UO_1456 (O_1456,N_29736,N_29202);
and UO_1457 (O_1457,N_28886,N_29061);
nand UO_1458 (O_1458,N_29865,N_29760);
or UO_1459 (O_1459,N_29751,N_28800);
nand UO_1460 (O_1460,N_29782,N_28784);
nand UO_1461 (O_1461,N_29736,N_29148);
and UO_1462 (O_1462,N_29080,N_29199);
nor UO_1463 (O_1463,N_29396,N_28533);
nor UO_1464 (O_1464,N_29796,N_28788);
xnor UO_1465 (O_1465,N_28526,N_29357);
or UO_1466 (O_1466,N_29663,N_29641);
nand UO_1467 (O_1467,N_29325,N_29931);
xor UO_1468 (O_1468,N_29487,N_28665);
xnor UO_1469 (O_1469,N_28736,N_28997);
and UO_1470 (O_1470,N_29652,N_29068);
nor UO_1471 (O_1471,N_28839,N_29589);
nor UO_1472 (O_1472,N_29993,N_28941);
nand UO_1473 (O_1473,N_29338,N_28744);
nand UO_1474 (O_1474,N_29102,N_28782);
xor UO_1475 (O_1475,N_28510,N_29101);
or UO_1476 (O_1476,N_28694,N_29015);
xor UO_1477 (O_1477,N_29779,N_29993);
nor UO_1478 (O_1478,N_29410,N_29823);
xor UO_1479 (O_1479,N_28925,N_29104);
and UO_1480 (O_1480,N_29630,N_29827);
xnor UO_1481 (O_1481,N_29713,N_29793);
and UO_1482 (O_1482,N_29016,N_28996);
nand UO_1483 (O_1483,N_29370,N_28904);
nor UO_1484 (O_1484,N_29799,N_29299);
xor UO_1485 (O_1485,N_29612,N_29676);
and UO_1486 (O_1486,N_29859,N_28991);
xnor UO_1487 (O_1487,N_29802,N_28723);
nand UO_1488 (O_1488,N_29186,N_28736);
nand UO_1489 (O_1489,N_28855,N_29180);
xor UO_1490 (O_1490,N_28851,N_28801);
or UO_1491 (O_1491,N_28934,N_29194);
xnor UO_1492 (O_1492,N_29670,N_29855);
or UO_1493 (O_1493,N_29511,N_29533);
nand UO_1494 (O_1494,N_29965,N_29432);
xor UO_1495 (O_1495,N_29252,N_29536);
nor UO_1496 (O_1496,N_29128,N_28551);
or UO_1497 (O_1497,N_29806,N_29745);
or UO_1498 (O_1498,N_29965,N_29960);
nor UO_1499 (O_1499,N_29535,N_28754);
or UO_1500 (O_1500,N_29550,N_29522);
or UO_1501 (O_1501,N_29195,N_28507);
nand UO_1502 (O_1502,N_29617,N_29780);
nand UO_1503 (O_1503,N_28840,N_28649);
nand UO_1504 (O_1504,N_28817,N_28714);
or UO_1505 (O_1505,N_28677,N_29190);
and UO_1506 (O_1506,N_29667,N_29610);
or UO_1507 (O_1507,N_29623,N_29131);
or UO_1508 (O_1508,N_29260,N_28868);
and UO_1509 (O_1509,N_28626,N_29679);
nand UO_1510 (O_1510,N_28955,N_29324);
nand UO_1511 (O_1511,N_29415,N_29601);
or UO_1512 (O_1512,N_29165,N_29135);
xnor UO_1513 (O_1513,N_29517,N_28800);
xnor UO_1514 (O_1514,N_29744,N_28934);
xnor UO_1515 (O_1515,N_29852,N_29427);
nor UO_1516 (O_1516,N_28756,N_29223);
nand UO_1517 (O_1517,N_29329,N_28508);
nand UO_1518 (O_1518,N_28580,N_29648);
or UO_1519 (O_1519,N_29442,N_29902);
xnor UO_1520 (O_1520,N_28745,N_29437);
xor UO_1521 (O_1521,N_28961,N_29997);
xnor UO_1522 (O_1522,N_28668,N_28527);
or UO_1523 (O_1523,N_28779,N_29002);
and UO_1524 (O_1524,N_28514,N_29118);
and UO_1525 (O_1525,N_29733,N_28629);
nor UO_1526 (O_1526,N_28816,N_28899);
or UO_1527 (O_1527,N_29521,N_29934);
nor UO_1528 (O_1528,N_28572,N_29231);
nor UO_1529 (O_1529,N_29476,N_28852);
nor UO_1530 (O_1530,N_29076,N_29653);
and UO_1531 (O_1531,N_29667,N_29542);
xnor UO_1532 (O_1532,N_29661,N_28520);
or UO_1533 (O_1533,N_29376,N_29417);
xnor UO_1534 (O_1534,N_28735,N_29276);
nand UO_1535 (O_1535,N_29252,N_28677);
xnor UO_1536 (O_1536,N_28625,N_29474);
nand UO_1537 (O_1537,N_29486,N_29695);
nand UO_1538 (O_1538,N_29295,N_29941);
and UO_1539 (O_1539,N_29061,N_28948);
nor UO_1540 (O_1540,N_29674,N_29420);
and UO_1541 (O_1541,N_29517,N_29489);
and UO_1542 (O_1542,N_28831,N_28666);
or UO_1543 (O_1543,N_29945,N_29019);
nand UO_1544 (O_1544,N_29532,N_29368);
xnor UO_1545 (O_1545,N_28661,N_29748);
nand UO_1546 (O_1546,N_28988,N_29274);
and UO_1547 (O_1547,N_29453,N_28871);
nor UO_1548 (O_1548,N_29525,N_29599);
xor UO_1549 (O_1549,N_29429,N_28778);
nand UO_1550 (O_1550,N_29796,N_29975);
xor UO_1551 (O_1551,N_29072,N_29534);
nand UO_1552 (O_1552,N_29922,N_28824);
nand UO_1553 (O_1553,N_29957,N_29693);
and UO_1554 (O_1554,N_28673,N_29336);
xor UO_1555 (O_1555,N_29667,N_29401);
xor UO_1556 (O_1556,N_29011,N_29751);
nor UO_1557 (O_1557,N_29070,N_29669);
and UO_1558 (O_1558,N_29485,N_29475);
and UO_1559 (O_1559,N_29868,N_29989);
xor UO_1560 (O_1560,N_29439,N_29575);
or UO_1561 (O_1561,N_29530,N_29212);
nand UO_1562 (O_1562,N_29116,N_29070);
nand UO_1563 (O_1563,N_29174,N_29310);
and UO_1564 (O_1564,N_28710,N_28675);
nor UO_1565 (O_1565,N_28782,N_28775);
nor UO_1566 (O_1566,N_29736,N_29452);
nor UO_1567 (O_1567,N_28555,N_29556);
nor UO_1568 (O_1568,N_28504,N_28841);
and UO_1569 (O_1569,N_29411,N_29216);
and UO_1570 (O_1570,N_29604,N_28894);
and UO_1571 (O_1571,N_29587,N_28624);
and UO_1572 (O_1572,N_28739,N_29190);
nand UO_1573 (O_1573,N_28885,N_29742);
nand UO_1574 (O_1574,N_29361,N_29124);
xnor UO_1575 (O_1575,N_29035,N_29496);
nand UO_1576 (O_1576,N_29748,N_28867);
or UO_1577 (O_1577,N_28555,N_28951);
or UO_1578 (O_1578,N_29484,N_29422);
and UO_1579 (O_1579,N_29970,N_28728);
nand UO_1580 (O_1580,N_28533,N_29143);
nor UO_1581 (O_1581,N_29246,N_29853);
xnor UO_1582 (O_1582,N_29239,N_29177);
nor UO_1583 (O_1583,N_28979,N_29812);
or UO_1584 (O_1584,N_29495,N_29671);
nor UO_1585 (O_1585,N_29019,N_29195);
or UO_1586 (O_1586,N_28862,N_29571);
or UO_1587 (O_1587,N_29165,N_29316);
nor UO_1588 (O_1588,N_29973,N_28956);
and UO_1589 (O_1589,N_29259,N_28951);
xor UO_1590 (O_1590,N_28781,N_29708);
and UO_1591 (O_1591,N_29431,N_28912);
nand UO_1592 (O_1592,N_29504,N_29024);
nand UO_1593 (O_1593,N_29061,N_29368);
nor UO_1594 (O_1594,N_28634,N_29703);
and UO_1595 (O_1595,N_28867,N_29635);
or UO_1596 (O_1596,N_28849,N_29466);
nand UO_1597 (O_1597,N_28620,N_28665);
or UO_1598 (O_1598,N_29282,N_29837);
xnor UO_1599 (O_1599,N_28636,N_29621);
nor UO_1600 (O_1600,N_29165,N_28693);
xor UO_1601 (O_1601,N_28571,N_28667);
and UO_1602 (O_1602,N_29791,N_29033);
and UO_1603 (O_1603,N_29555,N_29086);
nand UO_1604 (O_1604,N_28579,N_29556);
nor UO_1605 (O_1605,N_29447,N_28918);
nor UO_1606 (O_1606,N_28891,N_29067);
nand UO_1607 (O_1607,N_29628,N_29427);
nand UO_1608 (O_1608,N_28559,N_29597);
or UO_1609 (O_1609,N_28728,N_28585);
nor UO_1610 (O_1610,N_29858,N_29088);
nand UO_1611 (O_1611,N_28617,N_29018);
nand UO_1612 (O_1612,N_29443,N_29982);
and UO_1613 (O_1613,N_28629,N_29449);
nor UO_1614 (O_1614,N_29227,N_28549);
or UO_1615 (O_1615,N_28912,N_28824);
and UO_1616 (O_1616,N_29186,N_29158);
or UO_1617 (O_1617,N_29809,N_29914);
or UO_1618 (O_1618,N_29870,N_28799);
or UO_1619 (O_1619,N_28794,N_29900);
and UO_1620 (O_1620,N_29155,N_29933);
and UO_1621 (O_1621,N_29926,N_29980);
nor UO_1622 (O_1622,N_29688,N_28872);
or UO_1623 (O_1623,N_28696,N_29876);
nor UO_1624 (O_1624,N_28779,N_29434);
and UO_1625 (O_1625,N_29283,N_29648);
nor UO_1626 (O_1626,N_29406,N_29185);
nor UO_1627 (O_1627,N_28895,N_28556);
nor UO_1628 (O_1628,N_29779,N_28531);
nor UO_1629 (O_1629,N_29018,N_29125);
xor UO_1630 (O_1630,N_29248,N_29567);
xor UO_1631 (O_1631,N_29411,N_29012);
nand UO_1632 (O_1632,N_28917,N_29870);
nor UO_1633 (O_1633,N_28872,N_29028);
nor UO_1634 (O_1634,N_29532,N_28619);
xor UO_1635 (O_1635,N_29786,N_29514);
nand UO_1636 (O_1636,N_28921,N_28863);
and UO_1637 (O_1637,N_29698,N_28707);
and UO_1638 (O_1638,N_28815,N_29758);
and UO_1639 (O_1639,N_28872,N_28682);
or UO_1640 (O_1640,N_28545,N_29745);
xnor UO_1641 (O_1641,N_28681,N_29742);
nand UO_1642 (O_1642,N_28973,N_28955);
xnor UO_1643 (O_1643,N_28642,N_29888);
nor UO_1644 (O_1644,N_29930,N_28555);
or UO_1645 (O_1645,N_28856,N_29182);
or UO_1646 (O_1646,N_29892,N_28698);
nand UO_1647 (O_1647,N_29894,N_29848);
xor UO_1648 (O_1648,N_29921,N_29121);
nand UO_1649 (O_1649,N_28882,N_29475);
xnor UO_1650 (O_1650,N_28842,N_29780);
xnor UO_1651 (O_1651,N_29077,N_29811);
or UO_1652 (O_1652,N_28602,N_29950);
nor UO_1653 (O_1653,N_28559,N_29720);
xor UO_1654 (O_1654,N_29787,N_28816);
nor UO_1655 (O_1655,N_28694,N_28784);
xor UO_1656 (O_1656,N_29038,N_28993);
xor UO_1657 (O_1657,N_29695,N_29645);
and UO_1658 (O_1658,N_29922,N_29559);
xnor UO_1659 (O_1659,N_28595,N_28952);
or UO_1660 (O_1660,N_29239,N_29276);
nor UO_1661 (O_1661,N_28644,N_29777);
xnor UO_1662 (O_1662,N_29710,N_29382);
and UO_1663 (O_1663,N_29543,N_28913);
nand UO_1664 (O_1664,N_29430,N_29716);
and UO_1665 (O_1665,N_28501,N_28818);
nor UO_1666 (O_1666,N_28710,N_28942);
nor UO_1667 (O_1667,N_28815,N_29021);
nand UO_1668 (O_1668,N_29167,N_29237);
or UO_1669 (O_1669,N_29640,N_29168);
nor UO_1670 (O_1670,N_28610,N_28773);
xor UO_1671 (O_1671,N_29036,N_29526);
and UO_1672 (O_1672,N_28617,N_29739);
nand UO_1673 (O_1673,N_29816,N_29658);
xnor UO_1674 (O_1674,N_28738,N_29896);
and UO_1675 (O_1675,N_29698,N_29276);
or UO_1676 (O_1676,N_28770,N_29047);
nor UO_1677 (O_1677,N_28668,N_29779);
or UO_1678 (O_1678,N_29956,N_29223);
nand UO_1679 (O_1679,N_29876,N_29494);
or UO_1680 (O_1680,N_28814,N_29687);
nor UO_1681 (O_1681,N_29093,N_29853);
nor UO_1682 (O_1682,N_29569,N_29801);
or UO_1683 (O_1683,N_28677,N_28865);
nand UO_1684 (O_1684,N_28655,N_29438);
nor UO_1685 (O_1685,N_29747,N_28832);
and UO_1686 (O_1686,N_29354,N_29294);
or UO_1687 (O_1687,N_29048,N_29192);
xor UO_1688 (O_1688,N_29717,N_28934);
or UO_1689 (O_1689,N_29591,N_29880);
nor UO_1690 (O_1690,N_29604,N_28943);
nor UO_1691 (O_1691,N_28919,N_29522);
or UO_1692 (O_1692,N_29380,N_29103);
nor UO_1693 (O_1693,N_29143,N_28958);
or UO_1694 (O_1694,N_29583,N_29021);
or UO_1695 (O_1695,N_28763,N_29216);
nand UO_1696 (O_1696,N_29345,N_29216);
and UO_1697 (O_1697,N_29329,N_29809);
nand UO_1698 (O_1698,N_29366,N_29548);
xor UO_1699 (O_1699,N_28588,N_29277);
xor UO_1700 (O_1700,N_29771,N_29779);
and UO_1701 (O_1701,N_28910,N_29910);
and UO_1702 (O_1702,N_29343,N_28642);
xor UO_1703 (O_1703,N_29125,N_29448);
nor UO_1704 (O_1704,N_29786,N_29757);
and UO_1705 (O_1705,N_29627,N_28843);
or UO_1706 (O_1706,N_29082,N_28644);
xnor UO_1707 (O_1707,N_28578,N_28664);
nand UO_1708 (O_1708,N_29641,N_29950);
and UO_1709 (O_1709,N_29781,N_28863);
or UO_1710 (O_1710,N_28836,N_28993);
xor UO_1711 (O_1711,N_29439,N_28620);
nand UO_1712 (O_1712,N_29439,N_29688);
or UO_1713 (O_1713,N_28520,N_29713);
or UO_1714 (O_1714,N_29067,N_29710);
or UO_1715 (O_1715,N_28590,N_28670);
xor UO_1716 (O_1716,N_29103,N_28946);
and UO_1717 (O_1717,N_29289,N_29707);
nor UO_1718 (O_1718,N_29812,N_28910);
nand UO_1719 (O_1719,N_29535,N_29146);
nor UO_1720 (O_1720,N_28616,N_29468);
xor UO_1721 (O_1721,N_29247,N_29526);
and UO_1722 (O_1722,N_29968,N_29663);
or UO_1723 (O_1723,N_29025,N_29382);
nor UO_1724 (O_1724,N_29740,N_29707);
and UO_1725 (O_1725,N_29302,N_29410);
or UO_1726 (O_1726,N_29650,N_28732);
nand UO_1727 (O_1727,N_28538,N_29687);
or UO_1728 (O_1728,N_29721,N_28791);
nand UO_1729 (O_1729,N_29181,N_28715);
nor UO_1730 (O_1730,N_29191,N_29186);
nor UO_1731 (O_1731,N_29142,N_28552);
or UO_1732 (O_1732,N_29212,N_29521);
nor UO_1733 (O_1733,N_29363,N_28939);
nor UO_1734 (O_1734,N_28585,N_29773);
nand UO_1735 (O_1735,N_28907,N_29099);
nor UO_1736 (O_1736,N_29919,N_28558);
or UO_1737 (O_1737,N_28947,N_29314);
nand UO_1738 (O_1738,N_29443,N_29363);
nor UO_1739 (O_1739,N_29667,N_29956);
xor UO_1740 (O_1740,N_28923,N_29060);
and UO_1741 (O_1741,N_29542,N_28663);
nand UO_1742 (O_1742,N_28826,N_28709);
xor UO_1743 (O_1743,N_29761,N_28856);
nand UO_1744 (O_1744,N_29144,N_29731);
nor UO_1745 (O_1745,N_29775,N_29878);
or UO_1746 (O_1746,N_28538,N_29144);
nand UO_1747 (O_1747,N_29600,N_29963);
and UO_1748 (O_1748,N_29961,N_28670);
or UO_1749 (O_1749,N_29058,N_29137);
xnor UO_1750 (O_1750,N_29546,N_29960);
nand UO_1751 (O_1751,N_29556,N_29405);
xor UO_1752 (O_1752,N_29978,N_29889);
or UO_1753 (O_1753,N_29693,N_28899);
nor UO_1754 (O_1754,N_28918,N_29769);
xor UO_1755 (O_1755,N_29702,N_29529);
nand UO_1756 (O_1756,N_29867,N_29296);
nor UO_1757 (O_1757,N_29101,N_28585);
and UO_1758 (O_1758,N_29422,N_29978);
xor UO_1759 (O_1759,N_29509,N_29461);
nand UO_1760 (O_1760,N_29431,N_29827);
nand UO_1761 (O_1761,N_29578,N_28705);
nor UO_1762 (O_1762,N_29436,N_28876);
and UO_1763 (O_1763,N_29098,N_29005);
or UO_1764 (O_1764,N_28541,N_29340);
and UO_1765 (O_1765,N_29796,N_28650);
nor UO_1766 (O_1766,N_28902,N_28638);
nor UO_1767 (O_1767,N_29426,N_29739);
nor UO_1768 (O_1768,N_29755,N_29180);
or UO_1769 (O_1769,N_29687,N_29592);
or UO_1770 (O_1770,N_28706,N_29807);
nand UO_1771 (O_1771,N_28726,N_28994);
xor UO_1772 (O_1772,N_28915,N_29122);
nor UO_1773 (O_1773,N_29784,N_29877);
nor UO_1774 (O_1774,N_28533,N_28572);
xor UO_1775 (O_1775,N_28976,N_29023);
xor UO_1776 (O_1776,N_29099,N_29353);
nand UO_1777 (O_1777,N_29147,N_29398);
and UO_1778 (O_1778,N_29152,N_28538);
and UO_1779 (O_1779,N_28579,N_29237);
nor UO_1780 (O_1780,N_28735,N_29813);
and UO_1781 (O_1781,N_29403,N_29815);
xor UO_1782 (O_1782,N_29442,N_29764);
nor UO_1783 (O_1783,N_29995,N_29946);
nor UO_1784 (O_1784,N_29489,N_28669);
nor UO_1785 (O_1785,N_29665,N_28726);
nand UO_1786 (O_1786,N_29809,N_28859);
or UO_1787 (O_1787,N_28826,N_28637);
or UO_1788 (O_1788,N_29973,N_29815);
xnor UO_1789 (O_1789,N_28840,N_28872);
nand UO_1790 (O_1790,N_28738,N_28526);
and UO_1791 (O_1791,N_29135,N_28742);
or UO_1792 (O_1792,N_28915,N_29088);
or UO_1793 (O_1793,N_29677,N_29969);
xnor UO_1794 (O_1794,N_29650,N_28658);
nand UO_1795 (O_1795,N_29194,N_28658);
nand UO_1796 (O_1796,N_29481,N_28627);
nor UO_1797 (O_1797,N_29792,N_29634);
nand UO_1798 (O_1798,N_29634,N_29567);
or UO_1799 (O_1799,N_28761,N_29086);
xor UO_1800 (O_1800,N_29021,N_29346);
xnor UO_1801 (O_1801,N_29919,N_29122);
nand UO_1802 (O_1802,N_28783,N_29428);
xnor UO_1803 (O_1803,N_28665,N_28761);
xnor UO_1804 (O_1804,N_29095,N_28811);
nor UO_1805 (O_1805,N_29356,N_28971);
or UO_1806 (O_1806,N_28669,N_29211);
nor UO_1807 (O_1807,N_28720,N_29304);
and UO_1808 (O_1808,N_29353,N_28917);
nor UO_1809 (O_1809,N_28665,N_29481);
nand UO_1810 (O_1810,N_29121,N_29603);
or UO_1811 (O_1811,N_29624,N_29255);
nor UO_1812 (O_1812,N_29668,N_29741);
xor UO_1813 (O_1813,N_28803,N_29346);
or UO_1814 (O_1814,N_29873,N_29020);
nand UO_1815 (O_1815,N_29634,N_28778);
and UO_1816 (O_1816,N_29925,N_29824);
and UO_1817 (O_1817,N_29271,N_29533);
nand UO_1818 (O_1818,N_28876,N_29191);
or UO_1819 (O_1819,N_29860,N_29756);
nand UO_1820 (O_1820,N_29127,N_29719);
nand UO_1821 (O_1821,N_28703,N_29877);
nor UO_1822 (O_1822,N_28876,N_29131);
nor UO_1823 (O_1823,N_29147,N_28921);
xnor UO_1824 (O_1824,N_29621,N_28687);
and UO_1825 (O_1825,N_29941,N_28638);
nand UO_1826 (O_1826,N_29781,N_29497);
xnor UO_1827 (O_1827,N_29922,N_29643);
or UO_1828 (O_1828,N_29896,N_29058);
nand UO_1829 (O_1829,N_29942,N_29428);
nand UO_1830 (O_1830,N_29147,N_28593);
xor UO_1831 (O_1831,N_28923,N_28685);
and UO_1832 (O_1832,N_28633,N_29815);
or UO_1833 (O_1833,N_28875,N_29045);
nor UO_1834 (O_1834,N_29028,N_29321);
xnor UO_1835 (O_1835,N_29863,N_29655);
nand UO_1836 (O_1836,N_28830,N_28661);
nor UO_1837 (O_1837,N_29340,N_28571);
nand UO_1838 (O_1838,N_29531,N_29691);
or UO_1839 (O_1839,N_29013,N_28967);
and UO_1840 (O_1840,N_28915,N_29164);
or UO_1841 (O_1841,N_29876,N_29290);
or UO_1842 (O_1842,N_28869,N_29076);
nor UO_1843 (O_1843,N_28968,N_29358);
or UO_1844 (O_1844,N_29343,N_28962);
or UO_1845 (O_1845,N_29207,N_29264);
nand UO_1846 (O_1846,N_29216,N_29598);
nand UO_1847 (O_1847,N_29103,N_28748);
or UO_1848 (O_1848,N_28788,N_28902);
and UO_1849 (O_1849,N_29099,N_29993);
nor UO_1850 (O_1850,N_29936,N_29226);
nor UO_1851 (O_1851,N_28620,N_29231);
or UO_1852 (O_1852,N_28708,N_28775);
or UO_1853 (O_1853,N_28531,N_29938);
and UO_1854 (O_1854,N_28653,N_29533);
and UO_1855 (O_1855,N_29186,N_28835);
nand UO_1856 (O_1856,N_29351,N_28834);
or UO_1857 (O_1857,N_29775,N_29393);
xor UO_1858 (O_1858,N_29981,N_29799);
and UO_1859 (O_1859,N_29677,N_29370);
and UO_1860 (O_1860,N_29858,N_29093);
xnor UO_1861 (O_1861,N_29091,N_29613);
nor UO_1862 (O_1862,N_29430,N_29784);
and UO_1863 (O_1863,N_29643,N_28760);
nand UO_1864 (O_1864,N_29662,N_28790);
nand UO_1865 (O_1865,N_29597,N_28975);
xnor UO_1866 (O_1866,N_28769,N_29898);
or UO_1867 (O_1867,N_29323,N_29214);
xnor UO_1868 (O_1868,N_28869,N_29852);
nor UO_1869 (O_1869,N_29283,N_28626);
xnor UO_1870 (O_1870,N_29532,N_29424);
nor UO_1871 (O_1871,N_29231,N_28911);
and UO_1872 (O_1872,N_29375,N_29988);
or UO_1873 (O_1873,N_29053,N_29682);
and UO_1874 (O_1874,N_29094,N_28744);
nand UO_1875 (O_1875,N_29710,N_29907);
nand UO_1876 (O_1876,N_29413,N_29528);
and UO_1877 (O_1877,N_28599,N_29411);
and UO_1878 (O_1878,N_28912,N_28949);
xor UO_1879 (O_1879,N_29473,N_29896);
nand UO_1880 (O_1880,N_28848,N_29008);
nand UO_1881 (O_1881,N_29713,N_29734);
or UO_1882 (O_1882,N_29800,N_28834);
nand UO_1883 (O_1883,N_29321,N_28684);
xor UO_1884 (O_1884,N_29037,N_29056);
nand UO_1885 (O_1885,N_29700,N_29032);
or UO_1886 (O_1886,N_29275,N_28769);
or UO_1887 (O_1887,N_28625,N_28604);
nor UO_1888 (O_1888,N_28638,N_29428);
or UO_1889 (O_1889,N_29910,N_29182);
nand UO_1890 (O_1890,N_29486,N_29438);
xnor UO_1891 (O_1891,N_28896,N_28738);
and UO_1892 (O_1892,N_29880,N_28732);
nor UO_1893 (O_1893,N_29995,N_29224);
xnor UO_1894 (O_1894,N_28826,N_29942);
nor UO_1895 (O_1895,N_29237,N_29644);
nor UO_1896 (O_1896,N_29675,N_29001);
nand UO_1897 (O_1897,N_29490,N_28976);
nand UO_1898 (O_1898,N_29694,N_29592);
or UO_1899 (O_1899,N_28900,N_29446);
nor UO_1900 (O_1900,N_29953,N_29999);
and UO_1901 (O_1901,N_28541,N_28679);
nor UO_1902 (O_1902,N_29621,N_29706);
and UO_1903 (O_1903,N_29396,N_29195);
nand UO_1904 (O_1904,N_29202,N_29643);
and UO_1905 (O_1905,N_28541,N_29821);
nand UO_1906 (O_1906,N_29280,N_29062);
nor UO_1907 (O_1907,N_28636,N_29535);
xor UO_1908 (O_1908,N_28867,N_29094);
xor UO_1909 (O_1909,N_28718,N_29847);
and UO_1910 (O_1910,N_29351,N_29992);
nand UO_1911 (O_1911,N_28573,N_28653);
nand UO_1912 (O_1912,N_29045,N_28770);
nand UO_1913 (O_1913,N_29073,N_28971);
nand UO_1914 (O_1914,N_28823,N_29375);
nand UO_1915 (O_1915,N_29831,N_29872);
or UO_1916 (O_1916,N_29012,N_29093);
xor UO_1917 (O_1917,N_28685,N_28918);
nand UO_1918 (O_1918,N_29370,N_28528);
or UO_1919 (O_1919,N_29717,N_29261);
nand UO_1920 (O_1920,N_29693,N_28742);
or UO_1921 (O_1921,N_28778,N_28974);
nor UO_1922 (O_1922,N_28701,N_28731);
nor UO_1923 (O_1923,N_29439,N_29789);
nand UO_1924 (O_1924,N_29363,N_29883);
nand UO_1925 (O_1925,N_29363,N_29461);
nand UO_1926 (O_1926,N_28714,N_29513);
nand UO_1927 (O_1927,N_28848,N_29098);
xnor UO_1928 (O_1928,N_28702,N_29048);
xor UO_1929 (O_1929,N_29792,N_28608);
and UO_1930 (O_1930,N_29547,N_28536);
and UO_1931 (O_1931,N_29867,N_28838);
and UO_1932 (O_1932,N_28775,N_28609);
or UO_1933 (O_1933,N_29988,N_29536);
nand UO_1934 (O_1934,N_28550,N_28588);
or UO_1935 (O_1935,N_29637,N_29816);
nor UO_1936 (O_1936,N_29268,N_28601);
nor UO_1937 (O_1937,N_29814,N_28952);
nand UO_1938 (O_1938,N_29400,N_28989);
nor UO_1939 (O_1939,N_29917,N_29063);
nand UO_1940 (O_1940,N_29077,N_29800);
xor UO_1941 (O_1941,N_29548,N_29505);
xor UO_1942 (O_1942,N_29415,N_29033);
and UO_1943 (O_1943,N_28938,N_29211);
nand UO_1944 (O_1944,N_28834,N_28504);
and UO_1945 (O_1945,N_28930,N_29338);
and UO_1946 (O_1946,N_29218,N_28792);
xor UO_1947 (O_1947,N_29269,N_29016);
or UO_1948 (O_1948,N_28577,N_28778);
or UO_1949 (O_1949,N_29282,N_29263);
and UO_1950 (O_1950,N_29645,N_29460);
xnor UO_1951 (O_1951,N_28981,N_28858);
nand UO_1952 (O_1952,N_29901,N_28563);
and UO_1953 (O_1953,N_29107,N_29074);
nand UO_1954 (O_1954,N_28823,N_29174);
nand UO_1955 (O_1955,N_29641,N_29572);
xor UO_1956 (O_1956,N_29203,N_29617);
and UO_1957 (O_1957,N_29145,N_29519);
or UO_1958 (O_1958,N_29507,N_29461);
nor UO_1959 (O_1959,N_29975,N_28742);
nand UO_1960 (O_1960,N_29981,N_28771);
and UO_1961 (O_1961,N_29719,N_29786);
xnor UO_1962 (O_1962,N_29171,N_29535);
and UO_1963 (O_1963,N_28932,N_29906);
nand UO_1964 (O_1964,N_28668,N_29333);
and UO_1965 (O_1965,N_29668,N_28841);
nand UO_1966 (O_1966,N_29225,N_28700);
or UO_1967 (O_1967,N_29341,N_29963);
nor UO_1968 (O_1968,N_29722,N_29417);
or UO_1969 (O_1969,N_28698,N_28625);
or UO_1970 (O_1970,N_29862,N_29059);
nor UO_1971 (O_1971,N_28787,N_28509);
and UO_1972 (O_1972,N_28522,N_29900);
nand UO_1973 (O_1973,N_29167,N_28663);
xor UO_1974 (O_1974,N_29977,N_28514);
nor UO_1975 (O_1975,N_29823,N_28663);
nor UO_1976 (O_1976,N_28808,N_29013);
or UO_1977 (O_1977,N_29854,N_28570);
or UO_1978 (O_1978,N_28926,N_29966);
and UO_1979 (O_1979,N_28549,N_29206);
xnor UO_1980 (O_1980,N_28888,N_28783);
xor UO_1981 (O_1981,N_28950,N_29805);
nor UO_1982 (O_1982,N_29127,N_29059);
nand UO_1983 (O_1983,N_29889,N_29520);
nor UO_1984 (O_1984,N_29796,N_29773);
nand UO_1985 (O_1985,N_29625,N_29373);
nor UO_1986 (O_1986,N_29554,N_28560);
or UO_1987 (O_1987,N_28899,N_29832);
or UO_1988 (O_1988,N_29266,N_29794);
or UO_1989 (O_1989,N_28678,N_29235);
or UO_1990 (O_1990,N_29495,N_28715);
nor UO_1991 (O_1991,N_28639,N_29014);
nor UO_1992 (O_1992,N_28932,N_29452);
and UO_1993 (O_1993,N_29093,N_28592);
nor UO_1994 (O_1994,N_29876,N_29633);
xnor UO_1995 (O_1995,N_28858,N_29871);
nand UO_1996 (O_1996,N_28556,N_28833);
nor UO_1997 (O_1997,N_29249,N_29588);
and UO_1998 (O_1998,N_29570,N_28725);
nand UO_1999 (O_1999,N_29078,N_29789);
nand UO_2000 (O_2000,N_28618,N_28561);
nand UO_2001 (O_2001,N_29566,N_29948);
nor UO_2002 (O_2002,N_29353,N_29357);
nand UO_2003 (O_2003,N_28973,N_29073);
xnor UO_2004 (O_2004,N_29751,N_29844);
or UO_2005 (O_2005,N_29496,N_28510);
and UO_2006 (O_2006,N_29738,N_29616);
or UO_2007 (O_2007,N_29656,N_28877);
xnor UO_2008 (O_2008,N_29473,N_29521);
or UO_2009 (O_2009,N_29057,N_29723);
nand UO_2010 (O_2010,N_29494,N_28628);
and UO_2011 (O_2011,N_28524,N_28963);
and UO_2012 (O_2012,N_29935,N_28500);
or UO_2013 (O_2013,N_29150,N_29375);
xor UO_2014 (O_2014,N_29337,N_29309);
nand UO_2015 (O_2015,N_28716,N_29779);
nor UO_2016 (O_2016,N_28557,N_29864);
xor UO_2017 (O_2017,N_28617,N_29655);
and UO_2018 (O_2018,N_29349,N_29454);
or UO_2019 (O_2019,N_29422,N_29510);
nor UO_2020 (O_2020,N_29051,N_29637);
xnor UO_2021 (O_2021,N_29338,N_28920);
xor UO_2022 (O_2022,N_29815,N_28877);
nand UO_2023 (O_2023,N_29133,N_29745);
or UO_2024 (O_2024,N_29314,N_29797);
nor UO_2025 (O_2025,N_28840,N_29564);
nor UO_2026 (O_2026,N_29820,N_29522);
or UO_2027 (O_2027,N_29477,N_28863);
or UO_2028 (O_2028,N_29469,N_29364);
nor UO_2029 (O_2029,N_29793,N_29700);
xnor UO_2030 (O_2030,N_29329,N_29664);
xnor UO_2031 (O_2031,N_29838,N_29606);
nand UO_2032 (O_2032,N_28863,N_29722);
and UO_2033 (O_2033,N_29143,N_28889);
nor UO_2034 (O_2034,N_28994,N_29891);
and UO_2035 (O_2035,N_28798,N_29476);
nor UO_2036 (O_2036,N_29299,N_28722);
and UO_2037 (O_2037,N_29815,N_29208);
xnor UO_2038 (O_2038,N_28898,N_29704);
xor UO_2039 (O_2039,N_28770,N_29530);
nor UO_2040 (O_2040,N_29231,N_29021);
and UO_2041 (O_2041,N_28896,N_29313);
xor UO_2042 (O_2042,N_28764,N_29416);
nand UO_2043 (O_2043,N_29927,N_29503);
xnor UO_2044 (O_2044,N_29004,N_28857);
nor UO_2045 (O_2045,N_28945,N_29394);
nand UO_2046 (O_2046,N_28898,N_29490);
nand UO_2047 (O_2047,N_28886,N_29606);
xor UO_2048 (O_2048,N_29993,N_28758);
nor UO_2049 (O_2049,N_29010,N_29954);
nor UO_2050 (O_2050,N_28526,N_28972);
nor UO_2051 (O_2051,N_28951,N_29759);
or UO_2052 (O_2052,N_29438,N_28692);
xnor UO_2053 (O_2053,N_28553,N_29473);
xor UO_2054 (O_2054,N_29251,N_28884);
nor UO_2055 (O_2055,N_28626,N_29754);
or UO_2056 (O_2056,N_29978,N_29094);
nand UO_2057 (O_2057,N_28859,N_28783);
or UO_2058 (O_2058,N_29819,N_29016);
or UO_2059 (O_2059,N_29422,N_28535);
or UO_2060 (O_2060,N_29284,N_28762);
nor UO_2061 (O_2061,N_29534,N_29385);
and UO_2062 (O_2062,N_29207,N_29629);
or UO_2063 (O_2063,N_28765,N_28987);
and UO_2064 (O_2064,N_29928,N_29550);
or UO_2065 (O_2065,N_29300,N_29755);
xnor UO_2066 (O_2066,N_28522,N_28756);
and UO_2067 (O_2067,N_29229,N_29985);
and UO_2068 (O_2068,N_28734,N_29608);
nand UO_2069 (O_2069,N_29207,N_29784);
and UO_2070 (O_2070,N_28879,N_29170);
xor UO_2071 (O_2071,N_29152,N_29262);
xor UO_2072 (O_2072,N_28844,N_29295);
nand UO_2073 (O_2073,N_29046,N_29672);
xor UO_2074 (O_2074,N_29883,N_28849);
nand UO_2075 (O_2075,N_28717,N_28991);
xor UO_2076 (O_2076,N_28938,N_28826);
nor UO_2077 (O_2077,N_29747,N_28807);
and UO_2078 (O_2078,N_29598,N_28523);
and UO_2079 (O_2079,N_29537,N_29294);
and UO_2080 (O_2080,N_28664,N_29747);
and UO_2081 (O_2081,N_29757,N_29188);
xnor UO_2082 (O_2082,N_29341,N_29749);
nor UO_2083 (O_2083,N_28972,N_29098);
or UO_2084 (O_2084,N_29979,N_29064);
nor UO_2085 (O_2085,N_28779,N_29706);
xnor UO_2086 (O_2086,N_29520,N_29702);
and UO_2087 (O_2087,N_29423,N_29035);
xnor UO_2088 (O_2088,N_29223,N_28926);
xor UO_2089 (O_2089,N_28502,N_29835);
and UO_2090 (O_2090,N_28596,N_29637);
nand UO_2091 (O_2091,N_29603,N_29484);
and UO_2092 (O_2092,N_28676,N_29017);
or UO_2093 (O_2093,N_29322,N_28581);
nor UO_2094 (O_2094,N_28887,N_29315);
or UO_2095 (O_2095,N_29577,N_29529);
or UO_2096 (O_2096,N_29385,N_29286);
and UO_2097 (O_2097,N_28546,N_28549);
nor UO_2098 (O_2098,N_29698,N_29459);
and UO_2099 (O_2099,N_28946,N_28916);
or UO_2100 (O_2100,N_29822,N_29562);
xnor UO_2101 (O_2101,N_29023,N_29467);
nand UO_2102 (O_2102,N_28977,N_29661);
or UO_2103 (O_2103,N_29439,N_29925);
or UO_2104 (O_2104,N_29843,N_29856);
nand UO_2105 (O_2105,N_29754,N_29351);
nand UO_2106 (O_2106,N_29142,N_29844);
or UO_2107 (O_2107,N_29465,N_28962);
nand UO_2108 (O_2108,N_29528,N_29751);
xnor UO_2109 (O_2109,N_29744,N_29400);
or UO_2110 (O_2110,N_28719,N_29287);
and UO_2111 (O_2111,N_28712,N_28651);
xor UO_2112 (O_2112,N_28841,N_29308);
xor UO_2113 (O_2113,N_29910,N_29970);
nor UO_2114 (O_2114,N_28611,N_29608);
or UO_2115 (O_2115,N_28562,N_29699);
xor UO_2116 (O_2116,N_29077,N_29134);
nand UO_2117 (O_2117,N_29696,N_28591);
nand UO_2118 (O_2118,N_29315,N_28918);
and UO_2119 (O_2119,N_28933,N_29967);
and UO_2120 (O_2120,N_29886,N_29223);
or UO_2121 (O_2121,N_29969,N_28596);
or UO_2122 (O_2122,N_29713,N_28504);
or UO_2123 (O_2123,N_29009,N_28630);
xor UO_2124 (O_2124,N_29481,N_29107);
nor UO_2125 (O_2125,N_29365,N_29872);
xnor UO_2126 (O_2126,N_28579,N_28511);
nor UO_2127 (O_2127,N_29840,N_29566);
nand UO_2128 (O_2128,N_29441,N_29410);
xnor UO_2129 (O_2129,N_29521,N_29816);
nor UO_2130 (O_2130,N_29863,N_28577);
and UO_2131 (O_2131,N_29455,N_28868);
xnor UO_2132 (O_2132,N_28585,N_29539);
nand UO_2133 (O_2133,N_28661,N_29913);
and UO_2134 (O_2134,N_29274,N_29972);
nor UO_2135 (O_2135,N_28910,N_28531);
and UO_2136 (O_2136,N_29287,N_29539);
or UO_2137 (O_2137,N_28606,N_28983);
or UO_2138 (O_2138,N_28669,N_29307);
xor UO_2139 (O_2139,N_29288,N_29029);
xor UO_2140 (O_2140,N_29166,N_29694);
and UO_2141 (O_2141,N_28565,N_29108);
nor UO_2142 (O_2142,N_29678,N_29059);
xnor UO_2143 (O_2143,N_29311,N_28565);
xor UO_2144 (O_2144,N_28804,N_29372);
and UO_2145 (O_2145,N_28853,N_29994);
nor UO_2146 (O_2146,N_28799,N_29941);
nand UO_2147 (O_2147,N_29056,N_28969);
nand UO_2148 (O_2148,N_28513,N_29195);
xnor UO_2149 (O_2149,N_28913,N_29383);
nand UO_2150 (O_2150,N_29912,N_28821);
xnor UO_2151 (O_2151,N_29200,N_29930);
nor UO_2152 (O_2152,N_28714,N_29011);
and UO_2153 (O_2153,N_29120,N_28626);
nor UO_2154 (O_2154,N_28875,N_29529);
or UO_2155 (O_2155,N_29292,N_29749);
xor UO_2156 (O_2156,N_29243,N_29317);
nor UO_2157 (O_2157,N_28577,N_29778);
and UO_2158 (O_2158,N_28519,N_29595);
xor UO_2159 (O_2159,N_29410,N_28826);
nand UO_2160 (O_2160,N_28592,N_29621);
nor UO_2161 (O_2161,N_28657,N_29669);
nand UO_2162 (O_2162,N_29543,N_28923);
nor UO_2163 (O_2163,N_29048,N_29136);
and UO_2164 (O_2164,N_28742,N_29841);
nand UO_2165 (O_2165,N_28611,N_29439);
nor UO_2166 (O_2166,N_29066,N_29813);
nor UO_2167 (O_2167,N_28519,N_29992);
nand UO_2168 (O_2168,N_29435,N_29663);
nand UO_2169 (O_2169,N_29766,N_28725);
or UO_2170 (O_2170,N_29290,N_29416);
nand UO_2171 (O_2171,N_29352,N_28684);
and UO_2172 (O_2172,N_29874,N_29087);
or UO_2173 (O_2173,N_29669,N_28666);
xor UO_2174 (O_2174,N_28535,N_29144);
nor UO_2175 (O_2175,N_28893,N_28598);
and UO_2176 (O_2176,N_28940,N_29917);
nor UO_2177 (O_2177,N_29712,N_28783);
xor UO_2178 (O_2178,N_29117,N_28546);
nor UO_2179 (O_2179,N_28684,N_28893);
nor UO_2180 (O_2180,N_28525,N_29193);
nor UO_2181 (O_2181,N_29140,N_29855);
nand UO_2182 (O_2182,N_28905,N_29974);
or UO_2183 (O_2183,N_29498,N_29802);
xor UO_2184 (O_2184,N_29792,N_28833);
xor UO_2185 (O_2185,N_28687,N_29286);
xnor UO_2186 (O_2186,N_28865,N_29835);
nand UO_2187 (O_2187,N_29236,N_28550);
nand UO_2188 (O_2188,N_29218,N_29131);
or UO_2189 (O_2189,N_29413,N_29959);
or UO_2190 (O_2190,N_29775,N_28759);
nand UO_2191 (O_2191,N_28763,N_28830);
and UO_2192 (O_2192,N_29253,N_28571);
and UO_2193 (O_2193,N_28875,N_28973);
xnor UO_2194 (O_2194,N_29648,N_29836);
nand UO_2195 (O_2195,N_29173,N_28600);
nand UO_2196 (O_2196,N_29599,N_29352);
nor UO_2197 (O_2197,N_29773,N_29595);
xor UO_2198 (O_2198,N_29517,N_29555);
nor UO_2199 (O_2199,N_29414,N_29913);
xnor UO_2200 (O_2200,N_29600,N_29313);
xnor UO_2201 (O_2201,N_29754,N_29406);
or UO_2202 (O_2202,N_29255,N_29792);
and UO_2203 (O_2203,N_29307,N_29769);
nand UO_2204 (O_2204,N_29186,N_29208);
and UO_2205 (O_2205,N_29236,N_29597);
nor UO_2206 (O_2206,N_29213,N_29394);
and UO_2207 (O_2207,N_29709,N_28638);
and UO_2208 (O_2208,N_28508,N_29389);
xnor UO_2209 (O_2209,N_28787,N_29728);
and UO_2210 (O_2210,N_28766,N_29050);
nand UO_2211 (O_2211,N_28641,N_28812);
xor UO_2212 (O_2212,N_28673,N_29501);
xnor UO_2213 (O_2213,N_29586,N_29014);
nand UO_2214 (O_2214,N_29681,N_29411);
and UO_2215 (O_2215,N_29897,N_29945);
xnor UO_2216 (O_2216,N_29988,N_28717);
nor UO_2217 (O_2217,N_29299,N_29886);
nor UO_2218 (O_2218,N_28830,N_28913);
nor UO_2219 (O_2219,N_28802,N_29008);
or UO_2220 (O_2220,N_28745,N_29576);
nor UO_2221 (O_2221,N_29018,N_28668);
nand UO_2222 (O_2222,N_28501,N_29349);
xnor UO_2223 (O_2223,N_29431,N_29804);
and UO_2224 (O_2224,N_29779,N_29261);
nand UO_2225 (O_2225,N_28791,N_29547);
or UO_2226 (O_2226,N_28745,N_29161);
nand UO_2227 (O_2227,N_29843,N_28763);
and UO_2228 (O_2228,N_28630,N_29029);
or UO_2229 (O_2229,N_28547,N_29989);
xor UO_2230 (O_2230,N_29443,N_29926);
and UO_2231 (O_2231,N_29108,N_29319);
xnor UO_2232 (O_2232,N_28675,N_29569);
xor UO_2233 (O_2233,N_29895,N_28685);
or UO_2234 (O_2234,N_29785,N_28796);
nor UO_2235 (O_2235,N_28658,N_28505);
and UO_2236 (O_2236,N_29336,N_29250);
nor UO_2237 (O_2237,N_29676,N_29046);
and UO_2238 (O_2238,N_28764,N_28739);
nor UO_2239 (O_2239,N_28879,N_29449);
xor UO_2240 (O_2240,N_28770,N_28778);
nor UO_2241 (O_2241,N_28908,N_29275);
xnor UO_2242 (O_2242,N_28961,N_29544);
xnor UO_2243 (O_2243,N_29472,N_28801);
or UO_2244 (O_2244,N_28811,N_29076);
xnor UO_2245 (O_2245,N_28583,N_29524);
or UO_2246 (O_2246,N_29914,N_29204);
xnor UO_2247 (O_2247,N_29710,N_29760);
xnor UO_2248 (O_2248,N_28537,N_29741);
or UO_2249 (O_2249,N_29047,N_29052);
or UO_2250 (O_2250,N_29621,N_29265);
nor UO_2251 (O_2251,N_29172,N_28521);
nand UO_2252 (O_2252,N_29035,N_29750);
and UO_2253 (O_2253,N_29458,N_28810);
xor UO_2254 (O_2254,N_29662,N_29185);
or UO_2255 (O_2255,N_29174,N_28513);
xnor UO_2256 (O_2256,N_29501,N_29407);
nor UO_2257 (O_2257,N_29144,N_29852);
nor UO_2258 (O_2258,N_29297,N_29429);
xnor UO_2259 (O_2259,N_29095,N_29368);
xor UO_2260 (O_2260,N_28595,N_28728);
nand UO_2261 (O_2261,N_28619,N_28940);
nor UO_2262 (O_2262,N_29644,N_29478);
nand UO_2263 (O_2263,N_29361,N_29976);
and UO_2264 (O_2264,N_29324,N_29148);
xor UO_2265 (O_2265,N_29264,N_29494);
xnor UO_2266 (O_2266,N_29746,N_28848);
nor UO_2267 (O_2267,N_29598,N_29380);
nor UO_2268 (O_2268,N_29351,N_29152);
xnor UO_2269 (O_2269,N_28638,N_29672);
nor UO_2270 (O_2270,N_28952,N_29673);
or UO_2271 (O_2271,N_29961,N_29529);
and UO_2272 (O_2272,N_28921,N_29816);
nand UO_2273 (O_2273,N_28851,N_29160);
xor UO_2274 (O_2274,N_28541,N_28650);
nor UO_2275 (O_2275,N_29623,N_29421);
nand UO_2276 (O_2276,N_29315,N_29711);
nor UO_2277 (O_2277,N_29106,N_28589);
xor UO_2278 (O_2278,N_28597,N_29208);
and UO_2279 (O_2279,N_29651,N_29638);
nor UO_2280 (O_2280,N_29363,N_28808);
nor UO_2281 (O_2281,N_29176,N_28630);
and UO_2282 (O_2282,N_29395,N_28944);
or UO_2283 (O_2283,N_29916,N_29351);
nor UO_2284 (O_2284,N_29009,N_29423);
or UO_2285 (O_2285,N_29642,N_29554);
xnor UO_2286 (O_2286,N_29810,N_29011);
nor UO_2287 (O_2287,N_29899,N_29417);
xor UO_2288 (O_2288,N_29352,N_29694);
nand UO_2289 (O_2289,N_29446,N_28712);
xnor UO_2290 (O_2290,N_29518,N_28830);
and UO_2291 (O_2291,N_29106,N_29972);
xnor UO_2292 (O_2292,N_28952,N_29441);
nand UO_2293 (O_2293,N_28503,N_29227);
nor UO_2294 (O_2294,N_29298,N_29458);
xnor UO_2295 (O_2295,N_29800,N_29194);
and UO_2296 (O_2296,N_28820,N_29227);
xnor UO_2297 (O_2297,N_29719,N_29611);
nand UO_2298 (O_2298,N_28541,N_29936);
xnor UO_2299 (O_2299,N_28702,N_29032);
nor UO_2300 (O_2300,N_29001,N_29059);
and UO_2301 (O_2301,N_28575,N_28939);
nand UO_2302 (O_2302,N_28746,N_29509);
nand UO_2303 (O_2303,N_29822,N_28812);
nor UO_2304 (O_2304,N_29102,N_29219);
nor UO_2305 (O_2305,N_29145,N_29346);
and UO_2306 (O_2306,N_29710,N_29507);
or UO_2307 (O_2307,N_28826,N_28591);
xnor UO_2308 (O_2308,N_29025,N_29267);
or UO_2309 (O_2309,N_29959,N_29242);
or UO_2310 (O_2310,N_29349,N_29296);
and UO_2311 (O_2311,N_29425,N_29365);
nor UO_2312 (O_2312,N_29964,N_29487);
nor UO_2313 (O_2313,N_29629,N_29258);
nor UO_2314 (O_2314,N_29853,N_28632);
nand UO_2315 (O_2315,N_29616,N_28560);
xor UO_2316 (O_2316,N_29606,N_28862);
xor UO_2317 (O_2317,N_28990,N_29730);
nor UO_2318 (O_2318,N_29350,N_29779);
or UO_2319 (O_2319,N_29878,N_29716);
or UO_2320 (O_2320,N_29996,N_29658);
and UO_2321 (O_2321,N_29499,N_29740);
and UO_2322 (O_2322,N_28601,N_29148);
nor UO_2323 (O_2323,N_29778,N_29494);
nor UO_2324 (O_2324,N_29714,N_29628);
nand UO_2325 (O_2325,N_29189,N_28950);
nand UO_2326 (O_2326,N_28935,N_28538);
nand UO_2327 (O_2327,N_28550,N_28674);
xnor UO_2328 (O_2328,N_29611,N_29629);
xor UO_2329 (O_2329,N_29356,N_29195);
or UO_2330 (O_2330,N_28709,N_28576);
nor UO_2331 (O_2331,N_28554,N_28911);
and UO_2332 (O_2332,N_28512,N_29013);
xor UO_2333 (O_2333,N_29010,N_28746);
nand UO_2334 (O_2334,N_29168,N_28569);
and UO_2335 (O_2335,N_29741,N_28626);
nor UO_2336 (O_2336,N_28653,N_28520);
and UO_2337 (O_2337,N_29959,N_29873);
nor UO_2338 (O_2338,N_29570,N_28568);
nor UO_2339 (O_2339,N_29461,N_29277);
xnor UO_2340 (O_2340,N_29161,N_28910);
and UO_2341 (O_2341,N_28998,N_29649);
xor UO_2342 (O_2342,N_29816,N_29633);
or UO_2343 (O_2343,N_29362,N_28633);
nor UO_2344 (O_2344,N_29738,N_29555);
or UO_2345 (O_2345,N_29158,N_29695);
nor UO_2346 (O_2346,N_28579,N_29398);
xnor UO_2347 (O_2347,N_28609,N_28557);
xnor UO_2348 (O_2348,N_28695,N_28510);
nor UO_2349 (O_2349,N_28618,N_29236);
nand UO_2350 (O_2350,N_29523,N_28863);
nor UO_2351 (O_2351,N_28750,N_29338);
nor UO_2352 (O_2352,N_29420,N_29877);
or UO_2353 (O_2353,N_28622,N_29219);
nor UO_2354 (O_2354,N_28794,N_29696);
xnor UO_2355 (O_2355,N_29694,N_29681);
and UO_2356 (O_2356,N_29452,N_29902);
nand UO_2357 (O_2357,N_28865,N_29779);
and UO_2358 (O_2358,N_29649,N_29243);
nor UO_2359 (O_2359,N_29916,N_28618);
xnor UO_2360 (O_2360,N_29076,N_28529);
and UO_2361 (O_2361,N_29465,N_29383);
and UO_2362 (O_2362,N_29293,N_29204);
and UO_2363 (O_2363,N_28560,N_29992);
xnor UO_2364 (O_2364,N_29755,N_29900);
nor UO_2365 (O_2365,N_28601,N_29997);
nor UO_2366 (O_2366,N_29869,N_29876);
nor UO_2367 (O_2367,N_29398,N_29301);
and UO_2368 (O_2368,N_29942,N_29499);
xnor UO_2369 (O_2369,N_28892,N_29871);
or UO_2370 (O_2370,N_28933,N_29143);
xnor UO_2371 (O_2371,N_29625,N_28745);
and UO_2372 (O_2372,N_29959,N_29397);
nand UO_2373 (O_2373,N_29566,N_28898);
xnor UO_2374 (O_2374,N_28715,N_29845);
or UO_2375 (O_2375,N_28789,N_28973);
nand UO_2376 (O_2376,N_28526,N_28791);
xnor UO_2377 (O_2377,N_28590,N_29700);
and UO_2378 (O_2378,N_29271,N_29906);
nand UO_2379 (O_2379,N_28517,N_29805);
nand UO_2380 (O_2380,N_29171,N_29681);
and UO_2381 (O_2381,N_29458,N_29158);
xor UO_2382 (O_2382,N_28977,N_29979);
xor UO_2383 (O_2383,N_29201,N_28904);
xor UO_2384 (O_2384,N_28896,N_29578);
or UO_2385 (O_2385,N_29254,N_28577);
nor UO_2386 (O_2386,N_29631,N_28618);
xor UO_2387 (O_2387,N_28762,N_29729);
and UO_2388 (O_2388,N_28788,N_29030);
nor UO_2389 (O_2389,N_29469,N_29397);
and UO_2390 (O_2390,N_29230,N_29418);
or UO_2391 (O_2391,N_29312,N_29511);
nor UO_2392 (O_2392,N_29497,N_29830);
or UO_2393 (O_2393,N_28790,N_29943);
nand UO_2394 (O_2394,N_29416,N_29403);
and UO_2395 (O_2395,N_28897,N_29397);
or UO_2396 (O_2396,N_28650,N_29778);
nand UO_2397 (O_2397,N_29931,N_28843);
nor UO_2398 (O_2398,N_29279,N_29345);
and UO_2399 (O_2399,N_29791,N_28896);
nor UO_2400 (O_2400,N_29226,N_28526);
or UO_2401 (O_2401,N_29975,N_29486);
nor UO_2402 (O_2402,N_28768,N_28937);
and UO_2403 (O_2403,N_29197,N_29561);
xnor UO_2404 (O_2404,N_29751,N_29091);
xor UO_2405 (O_2405,N_28661,N_29404);
nand UO_2406 (O_2406,N_29513,N_29519);
xor UO_2407 (O_2407,N_29196,N_28897);
nor UO_2408 (O_2408,N_29684,N_28531);
xor UO_2409 (O_2409,N_29965,N_28800);
xor UO_2410 (O_2410,N_28550,N_29328);
or UO_2411 (O_2411,N_29174,N_29189);
and UO_2412 (O_2412,N_28558,N_28930);
or UO_2413 (O_2413,N_29221,N_29252);
and UO_2414 (O_2414,N_29108,N_29956);
nor UO_2415 (O_2415,N_28522,N_28662);
nor UO_2416 (O_2416,N_28932,N_29742);
nand UO_2417 (O_2417,N_29214,N_28739);
or UO_2418 (O_2418,N_29677,N_29803);
nand UO_2419 (O_2419,N_28992,N_29605);
or UO_2420 (O_2420,N_29833,N_28875);
nor UO_2421 (O_2421,N_28782,N_28988);
or UO_2422 (O_2422,N_29529,N_29850);
nor UO_2423 (O_2423,N_28913,N_28829);
nor UO_2424 (O_2424,N_29752,N_29610);
xor UO_2425 (O_2425,N_29904,N_29715);
and UO_2426 (O_2426,N_29494,N_29156);
nand UO_2427 (O_2427,N_28742,N_29102);
nor UO_2428 (O_2428,N_29935,N_29389);
nor UO_2429 (O_2429,N_29856,N_28713);
xnor UO_2430 (O_2430,N_29312,N_28523);
and UO_2431 (O_2431,N_28509,N_29869);
or UO_2432 (O_2432,N_29994,N_29930);
and UO_2433 (O_2433,N_29345,N_28553);
and UO_2434 (O_2434,N_28786,N_29349);
xor UO_2435 (O_2435,N_29752,N_29390);
nand UO_2436 (O_2436,N_29530,N_28934);
nor UO_2437 (O_2437,N_29118,N_29879);
xnor UO_2438 (O_2438,N_29165,N_29828);
xnor UO_2439 (O_2439,N_29388,N_29899);
or UO_2440 (O_2440,N_28558,N_28738);
xor UO_2441 (O_2441,N_29209,N_29942);
nand UO_2442 (O_2442,N_28794,N_29651);
nor UO_2443 (O_2443,N_29200,N_29222);
xor UO_2444 (O_2444,N_29452,N_29944);
nor UO_2445 (O_2445,N_28984,N_28588);
or UO_2446 (O_2446,N_29707,N_29937);
and UO_2447 (O_2447,N_28874,N_28929);
nand UO_2448 (O_2448,N_28992,N_28927);
nand UO_2449 (O_2449,N_29504,N_29412);
nor UO_2450 (O_2450,N_29790,N_29846);
nand UO_2451 (O_2451,N_28655,N_29616);
and UO_2452 (O_2452,N_29022,N_28830);
xnor UO_2453 (O_2453,N_29626,N_29691);
nand UO_2454 (O_2454,N_29715,N_29059);
nor UO_2455 (O_2455,N_29631,N_28820);
nand UO_2456 (O_2456,N_29836,N_29397);
and UO_2457 (O_2457,N_29388,N_28537);
nor UO_2458 (O_2458,N_28900,N_29353);
and UO_2459 (O_2459,N_28622,N_28860);
xnor UO_2460 (O_2460,N_29623,N_28501);
or UO_2461 (O_2461,N_29034,N_29874);
nand UO_2462 (O_2462,N_28847,N_29892);
nor UO_2463 (O_2463,N_29995,N_29502);
nor UO_2464 (O_2464,N_28517,N_28888);
or UO_2465 (O_2465,N_28561,N_29484);
or UO_2466 (O_2466,N_28767,N_29091);
nand UO_2467 (O_2467,N_29341,N_29797);
and UO_2468 (O_2468,N_28848,N_29294);
nand UO_2469 (O_2469,N_29672,N_29799);
xor UO_2470 (O_2470,N_29319,N_28526);
xor UO_2471 (O_2471,N_28814,N_28880);
nor UO_2472 (O_2472,N_29887,N_29699);
and UO_2473 (O_2473,N_29472,N_29497);
xnor UO_2474 (O_2474,N_29981,N_29561);
nand UO_2475 (O_2475,N_29667,N_29633);
nand UO_2476 (O_2476,N_29387,N_29860);
xnor UO_2477 (O_2477,N_28846,N_29183);
xor UO_2478 (O_2478,N_29524,N_29562);
or UO_2479 (O_2479,N_28599,N_29663);
and UO_2480 (O_2480,N_29506,N_29704);
or UO_2481 (O_2481,N_29961,N_29851);
nand UO_2482 (O_2482,N_29276,N_29123);
xnor UO_2483 (O_2483,N_29821,N_29638);
and UO_2484 (O_2484,N_29047,N_28957);
nand UO_2485 (O_2485,N_29474,N_29785);
or UO_2486 (O_2486,N_29451,N_29000);
or UO_2487 (O_2487,N_28861,N_29493);
xor UO_2488 (O_2488,N_28956,N_29720);
nand UO_2489 (O_2489,N_28867,N_28605);
or UO_2490 (O_2490,N_29734,N_28555);
or UO_2491 (O_2491,N_29710,N_29202);
xnor UO_2492 (O_2492,N_28559,N_28915);
xnor UO_2493 (O_2493,N_29566,N_29475);
nand UO_2494 (O_2494,N_29485,N_29087);
nand UO_2495 (O_2495,N_28954,N_29242);
xnor UO_2496 (O_2496,N_29717,N_29747);
nor UO_2497 (O_2497,N_29264,N_29242);
nand UO_2498 (O_2498,N_28641,N_29635);
nand UO_2499 (O_2499,N_28659,N_29100);
nor UO_2500 (O_2500,N_29990,N_28969);
nand UO_2501 (O_2501,N_28512,N_29390);
nor UO_2502 (O_2502,N_28963,N_29120);
nor UO_2503 (O_2503,N_28678,N_29168);
or UO_2504 (O_2504,N_29041,N_29234);
and UO_2505 (O_2505,N_28965,N_28896);
nand UO_2506 (O_2506,N_28711,N_29894);
and UO_2507 (O_2507,N_29337,N_29090);
and UO_2508 (O_2508,N_28886,N_29149);
nand UO_2509 (O_2509,N_29698,N_28668);
xor UO_2510 (O_2510,N_29620,N_28582);
nand UO_2511 (O_2511,N_28776,N_29718);
nand UO_2512 (O_2512,N_28904,N_29561);
nand UO_2513 (O_2513,N_28718,N_29886);
nand UO_2514 (O_2514,N_28922,N_28559);
nor UO_2515 (O_2515,N_29817,N_28515);
or UO_2516 (O_2516,N_29006,N_29830);
nor UO_2517 (O_2517,N_29421,N_29715);
or UO_2518 (O_2518,N_29609,N_29056);
nor UO_2519 (O_2519,N_29177,N_29740);
and UO_2520 (O_2520,N_29374,N_28977);
or UO_2521 (O_2521,N_29978,N_29890);
or UO_2522 (O_2522,N_29997,N_29277);
or UO_2523 (O_2523,N_29187,N_29017);
xor UO_2524 (O_2524,N_29640,N_29139);
nand UO_2525 (O_2525,N_29772,N_29557);
nor UO_2526 (O_2526,N_29418,N_28977);
and UO_2527 (O_2527,N_29379,N_29192);
or UO_2528 (O_2528,N_29757,N_29155);
nand UO_2529 (O_2529,N_29301,N_29396);
or UO_2530 (O_2530,N_28519,N_29280);
or UO_2531 (O_2531,N_29434,N_28678);
xor UO_2532 (O_2532,N_29800,N_28878);
nor UO_2533 (O_2533,N_29327,N_28679);
or UO_2534 (O_2534,N_29871,N_29163);
nor UO_2535 (O_2535,N_28736,N_28509);
and UO_2536 (O_2536,N_29422,N_28930);
and UO_2537 (O_2537,N_29628,N_29313);
nand UO_2538 (O_2538,N_28715,N_29821);
nor UO_2539 (O_2539,N_29497,N_29994);
nor UO_2540 (O_2540,N_28854,N_29198);
nand UO_2541 (O_2541,N_29394,N_29285);
and UO_2542 (O_2542,N_29861,N_29556);
nor UO_2543 (O_2543,N_28568,N_29612);
and UO_2544 (O_2544,N_29281,N_28690);
or UO_2545 (O_2545,N_29284,N_29765);
nor UO_2546 (O_2546,N_28725,N_29442);
xor UO_2547 (O_2547,N_29831,N_29421);
and UO_2548 (O_2548,N_28506,N_29834);
and UO_2549 (O_2549,N_28946,N_29075);
and UO_2550 (O_2550,N_28862,N_28999);
xnor UO_2551 (O_2551,N_29142,N_29394);
or UO_2552 (O_2552,N_29026,N_29259);
and UO_2553 (O_2553,N_29798,N_29489);
or UO_2554 (O_2554,N_28763,N_29877);
nor UO_2555 (O_2555,N_29644,N_28782);
or UO_2556 (O_2556,N_29693,N_28877);
xor UO_2557 (O_2557,N_29248,N_29093);
and UO_2558 (O_2558,N_29525,N_28672);
and UO_2559 (O_2559,N_29538,N_29673);
xor UO_2560 (O_2560,N_29626,N_29677);
and UO_2561 (O_2561,N_28520,N_29097);
or UO_2562 (O_2562,N_28937,N_29945);
and UO_2563 (O_2563,N_29153,N_29555);
xnor UO_2564 (O_2564,N_29301,N_29272);
nor UO_2565 (O_2565,N_29618,N_28811);
and UO_2566 (O_2566,N_29706,N_29046);
or UO_2567 (O_2567,N_29076,N_28822);
xor UO_2568 (O_2568,N_28880,N_28687);
nand UO_2569 (O_2569,N_29500,N_29872);
nor UO_2570 (O_2570,N_29250,N_28707);
xor UO_2571 (O_2571,N_29692,N_29445);
nor UO_2572 (O_2572,N_29635,N_29941);
xnor UO_2573 (O_2573,N_29673,N_29504);
or UO_2574 (O_2574,N_29229,N_28949);
nand UO_2575 (O_2575,N_29785,N_28849);
or UO_2576 (O_2576,N_29393,N_29222);
xor UO_2577 (O_2577,N_29595,N_29463);
nor UO_2578 (O_2578,N_29755,N_29453);
nand UO_2579 (O_2579,N_28653,N_29835);
and UO_2580 (O_2580,N_28648,N_29216);
nor UO_2581 (O_2581,N_29825,N_29718);
or UO_2582 (O_2582,N_29904,N_29091);
nand UO_2583 (O_2583,N_29985,N_29467);
and UO_2584 (O_2584,N_29077,N_29810);
nand UO_2585 (O_2585,N_28995,N_28592);
nand UO_2586 (O_2586,N_28516,N_28822);
and UO_2587 (O_2587,N_29454,N_29650);
nand UO_2588 (O_2588,N_29014,N_29779);
nand UO_2589 (O_2589,N_29161,N_29450);
nor UO_2590 (O_2590,N_29111,N_29185);
or UO_2591 (O_2591,N_29420,N_28882);
and UO_2592 (O_2592,N_29105,N_29611);
and UO_2593 (O_2593,N_29957,N_29439);
nand UO_2594 (O_2594,N_29635,N_28822);
nand UO_2595 (O_2595,N_28542,N_28674);
xnor UO_2596 (O_2596,N_29476,N_28699);
nand UO_2597 (O_2597,N_29195,N_29865);
nor UO_2598 (O_2598,N_29094,N_29216);
nor UO_2599 (O_2599,N_28755,N_28905);
or UO_2600 (O_2600,N_29603,N_29964);
xnor UO_2601 (O_2601,N_28973,N_29470);
nand UO_2602 (O_2602,N_28801,N_29237);
or UO_2603 (O_2603,N_29828,N_29606);
or UO_2604 (O_2604,N_28503,N_29952);
and UO_2605 (O_2605,N_29082,N_29502);
and UO_2606 (O_2606,N_28770,N_28547);
xnor UO_2607 (O_2607,N_29417,N_28715);
xnor UO_2608 (O_2608,N_29096,N_29728);
xnor UO_2609 (O_2609,N_29863,N_28584);
or UO_2610 (O_2610,N_29463,N_29134);
xnor UO_2611 (O_2611,N_29429,N_29798);
nand UO_2612 (O_2612,N_29818,N_29502);
nand UO_2613 (O_2613,N_29996,N_29470);
or UO_2614 (O_2614,N_28668,N_28652);
or UO_2615 (O_2615,N_29213,N_28920);
or UO_2616 (O_2616,N_29248,N_29111);
and UO_2617 (O_2617,N_29989,N_29269);
or UO_2618 (O_2618,N_28886,N_29187);
and UO_2619 (O_2619,N_29341,N_29687);
or UO_2620 (O_2620,N_29806,N_29969);
or UO_2621 (O_2621,N_29910,N_28691);
xor UO_2622 (O_2622,N_29476,N_29963);
and UO_2623 (O_2623,N_28909,N_29896);
nand UO_2624 (O_2624,N_29766,N_29465);
nor UO_2625 (O_2625,N_29014,N_28780);
xnor UO_2626 (O_2626,N_28808,N_29653);
nor UO_2627 (O_2627,N_28646,N_29020);
xnor UO_2628 (O_2628,N_29931,N_29703);
and UO_2629 (O_2629,N_29933,N_29539);
nand UO_2630 (O_2630,N_29408,N_28876);
xnor UO_2631 (O_2631,N_29583,N_29793);
and UO_2632 (O_2632,N_29556,N_29150);
xnor UO_2633 (O_2633,N_29499,N_29986);
nor UO_2634 (O_2634,N_29145,N_28680);
and UO_2635 (O_2635,N_29507,N_29504);
or UO_2636 (O_2636,N_29861,N_29596);
xnor UO_2637 (O_2637,N_28992,N_28900);
or UO_2638 (O_2638,N_28737,N_29361);
and UO_2639 (O_2639,N_28725,N_28962);
xnor UO_2640 (O_2640,N_29451,N_28758);
nor UO_2641 (O_2641,N_29360,N_29002);
nand UO_2642 (O_2642,N_28800,N_29936);
or UO_2643 (O_2643,N_28835,N_29820);
nand UO_2644 (O_2644,N_29461,N_29379);
or UO_2645 (O_2645,N_29725,N_28595);
or UO_2646 (O_2646,N_29424,N_29247);
xor UO_2647 (O_2647,N_29916,N_28721);
and UO_2648 (O_2648,N_29724,N_28880);
nor UO_2649 (O_2649,N_29262,N_28678);
and UO_2650 (O_2650,N_28935,N_28600);
nor UO_2651 (O_2651,N_28958,N_28699);
or UO_2652 (O_2652,N_29981,N_29745);
xor UO_2653 (O_2653,N_28673,N_29782);
xnor UO_2654 (O_2654,N_29840,N_29017);
nand UO_2655 (O_2655,N_29441,N_29191);
xor UO_2656 (O_2656,N_28815,N_28836);
nand UO_2657 (O_2657,N_29036,N_29400);
xor UO_2658 (O_2658,N_29798,N_28945);
nor UO_2659 (O_2659,N_28572,N_29353);
or UO_2660 (O_2660,N_29287,N_29062);
nand UO_2661 (O_2661,N_29904,N_28553);
or UO_2662 (O_2662,N_29346,N_29936);
and UO_2663 (O_2663,N_28920,N_28942);
nor UO_2664 (O_2664,N_28771,N_29873);
nand UO_2665 (O_2665,N_29945,N_29204);
nand UO_2666 (O_2666,N_29279,N_28673);
nand UO_2667 (O_2667,N_29921,N_29725);
nor UO_2668 (O_2668,N_29764,N_28844);
nor UO_2669 (O_2669,N_29045,N_29842);
xor UO_2670 (O_2670,N_29817,N_28731);
xor UO_2671 (O_2671,N_29038,N_29868);
and UO_2672 (O_2672,N_29505,N_29616);
and UO_2673 (O_2673,N_28654,N_29682);
and UO_2674 (O_2674,N_29856,N_29571);
nand UO_2675 (O_2675,N_29051,N_29291);
or UO_2676 (O_2676,N_29492,N_29035);
nor UO_2677 (O_2677,N_29030,N_28766);
nor UO_2678 (O_2678,N_28581,N_29667);
xor UO_2679 (O_2679,N_29899,N_29522);
nor UO_2680 (O_2680,N_29227,N_29727);
nor UO_2681 (O_2681,N_28764,N_28628);
and UO_2682 (O_2682,N_28822,N_29572);
nor UO_2683 (O_2683,N_29550,N_29521);
or UO_2684 (O_2684,N_29758,N_28919);
or UO_2685 (O_2685,N_28812,N_28796);
nor UO_2686 (O_2686,N_29804,N_28883);
or UO_2687 (O_2687,N_29314,N_28603);
or UO_2688 (O_2688,N_29956,N_29666);
nor UO_2689 (O_2689,N_28847,N_29511);
xnor UO_2690 (O_2690,N_29181,N_29658);
nand UO_2691 (O_2691,N_29319,N_29972);
nor UO_2692 (O_2692,N_29734,N_29526);
xor UO_2693 (O_2693,N_28978,N_28979);
nand UO_2694 (O_2694,N_29357,N_29723);
nor UO_2695 (O_2695,N_28938,N_29096);
or UO_2696 (O_2696,N_28948,N_29899);
xor UO_2697 (O_2697,N_28520,N_29399);
nand UO_2698 (O_2698,N_28991,N_29123);
nand UO_2699 (O_2699,N_29170,N_28794);
or UO_2700 (O_2700,N_29005,N_29519);
nor UO_2701 (O_2701,N_28964,N_28743);
nand UO_2702 (O_2702,N_29431,N_29049);
nor UO_2703 (O_2703,N_29550,N_29892);
nand UO_2704 (O_2704,N_29871,N_29214);
xor UO_2705 (O_2705,N_29068,N_29939);
xor UO_2706 (O_2706,N_29770,N_29869);
or UO_2707 (O_2707,N_29883,N_29172);
and UO_2708 (O_2708,N_28912,N_29887);
nor UO_2709 (O_2709,N_29269,N_29391);
and UO_2710 (O_2710,N_29402,N_29399);
nand UO_2711 (O_2711,N_28693,N_29403);
nand UO_2712 (O_2712,N_29880,N_29291);
nor UO_2713 (O_2713,N_29311,N_28506);
xnor UO_2714 (O_2714,N_28719,N_28901);
and UO_2715 (O_2715,N_28774,N_29288);
nor UO_2716 (O_2716,N_29911,N_28689);
nor UO_2717 (O_2717,N_28924,N_28997);
nor UO_2718 (O_2718,N_29149,N_28718);
nand UO_2719 (O_2719,N_29900,N_29715);
and UO_2720 (O_2720,N_28779,N_28945);
nand UO_2721 (O_2721,N_29291,N_29660);
or UO_2722 (O_2722,N_29910,N_29349);
xnor UO_2723 (O_2723,N_29432,N_29300);
xor UO_2724 (O_2724,N_29701,N_29978);
and UO_2725 (O_2725,N_28619,N_29829);
or UO_2726 (O_2726,N_28973,N_29432);
or UO_2727 (O_2727,N_29472,N_29932);
and UO_2728 (O_2728,N_28965,N_28703);
xor UO_2729 (O_2729,N_28728,N_29328);
nor UO_2730 (O_2730,N_28661,N_29553);
nor UO_2731 (O_2731,N_29959,N_28708);
nor UO_2732 (O_2732,N_29491,N_29824);
or UO_2733 (O_2733,N_29536,N_29619);
nand UO_2734 (O_2734,N_29431,N_29720);
and UO_2735 (O_2735,N_29100,N_29824);
nor UO_2736 (O_2736,N_29936,N_29015);
xor UO_2737 (O_2737,N_29657,N_28893);
and UO_2738 (O_2738,N_29065,N_29525);
nor UO_2739 (O_2739,N_29770,N_29528);
nand UO_2740 (O_2740,N_28556,N_29609);
nand UO_2741 (O_2741,N_29888,N_28626);
nor UO_2742 (O_2742,N_28933,N_29184);
or UO_2743 (O_2743,N_29966,N_29572);
nand UO_2744 (O_2744,N_28605,N_29438);
or UO_2745 (O_2745,N_29134,N_29770);
nand UO_2746 (O_2746,N_29338,N_28523);
and UO_2747 (O_2747,N_29743,N_29845);
xor UO_2748 (O_2748,N_29739,N_28657);
and UO_2749 (O_2749,N_29970,N_28676);
and UO_2750 (O_2750,N_28639,N_28847);
nor UO_2751 (O_2751,N_28840,N_29804);
and UO_2752 (O_2752,N_29487,N_29317);
nor UO_2753 (O_2753,N_28692,N_29243);
xnor UO_2754 (O_2754,N_29412,N_29565);
nor UO_2755 (O_2755,N_29076,N_28840);
xor UO_2756 (O_2756,N_28845,N_29254);
or UO_2757 (O_2757,N_28999,N_29132);
xnor UO_2758 (O_2758,N_29690,N_28630);
xnor UO_2759 (O_2759,N_29558,N_28856);
nand UO_2760 (O_2760,N_29383,N_29819);
nand UO_2761 (O_2761,N_28734,N_29422);
and UO_2762 (O_2762,N_29208,N_28664);
and UO_2763 (O_2763,N_29131,N_28821);
or UO_2764 (O_2764,N_28967,N_29370);
and UO_2765 (O_2765,N_29278,N_28985);
or UO_2766 (O_2766,N_28802,N_28925);
and UO_2767 (O_2767,N_28805,N_29184);
xor UO_2768 (O_2768,N_28697,N_29986);
nand UO_2769 (O_2769,N_29586,N_29509);
nand UO_2770 (O_2770,N_28755,N_29215);
xor UO_2771 (O_2771,N_29458,N_29054);
xnor UO_2772 (O_2772,N_29638,N_28905);
nand UO_2773 (O_2773,N_29580,N_29296);
or UO_2774 (O_2774,N_29899,N_29878);
and UO_2775 (O_2775,N_29327,N_29005);
or UO_2776 (O_2776,N_29046,N_29331);
nor UO_2777 (O_2777,N_29264,N_28627);
xor UO_2778 (O_2778,N_29793,N_28579);
xnor UO_2779 (O_2779,N_29259,N_28914);
xnor UO_2780 (O_2780,N_29908,N_29638);
and UO_2781 (O_2781,N_29237,N_28965);
nor UO_2782 (O_2782,N_29131,N_29289);
nand UO_2783 (O_2783,N_29353,N_29055);
nand UO_2784 (O_2784,N_29000,N_29868);
xnor UO_2785 (O_2785,N_29497,N_29408);
xnor UO_2786 (O_2786,N_28712,N_28974);
xnor UO_2787 (O_2787,N_29946,N_29174);
xnor UO_2788 (O_2788,N_28629,N_29448);
or UO_2789 (O_2789,N_28638,N_29541);
and UO_2790 (O_2790,N_28855,N_29604);
nand UO_2791 (O_2791,N_29656,N_29891);
or UO_2792 (O_2792,N_28567,N_29459);
xor UO_2793 (O_2793,N_29039,N_29633);
and UO_2794 (O_2794,N_28537,N_29630);
nand UO_2795 (O_2795,N_29458,N_29934);
nand UO_2796 (O_2796,N_29837,N_29168);
nand UO_2797 (O_2797,N_28762,N_29002);
or UO_2798 (O_2798,N_29405,N_29058);
nand UO_2799 (O_2799,N_28851,N_28986);
or UO_2800 (O_2800,N_29405,N_29374);
xor UO_2801 (O_2801,N_28666,N_29295);
or UO_2802 (O_2802,N_29551,N_29990);
xnor UO_2803 (O_2803,N_29773,N_29517);
nor UO_2804 (O_2804,N_29716,N_29975);
nand UO_2805 (O_2805,N_29202,N_29054);
or UO_2806 (O_2806,N_29434,N_29150);
nor UO_2807 (O_2807,N_29602,N_29851);
xnor UO_2808 (O_2808,N_29824,N_29007);
nor UO_2809 (O_2809,N_29627,N_29487);
nor UO_2810 (O_2810,N_29118,N_28706);
xor UO_2811 (O_2811,N_28971,N_29719);
or UO_2812 (O_2812,N_28669,N_28690);
or UO_2813 (O_2813,N_29334,N_29005);
nor UO_2814 (O_2814,N_29038,N_29621);
and UO_2815 (O_2815,N_29300,N_28544);
or UO_2816 (O_2816,N_29520,N_28960);
xnor UO_2817 (O_2817,N_29604,N_29430);
or UO_2818 (O_2818,N_28610,N_29656);
or UO_2819 (O_2819,N_29221,N_28748);
and UO_2820 (O_2820,N_29882,N_29635);
nand UO_2821 (O_2821,N_29954,N_29520);
or UO_2822 (O_2822,N_28856,N_29457);
and UO_2823 (O_2823,N_29256,N_29251);
and UO_2824 (O_2824,N_29708,N_29114);
and UO_2825 (O_2825,N_28952,N_29419);
nor UO_2826 (O_2826,N_29748,N_29186);
xor UO_2827 (O_2827,N_29201,N_28580);
xnor UO_2828 (O_2828,N_29089,N_29749);
nor UO_2829 (O_2829,N_29678,N_28673);
or UO_2830 (O_2830,N_29668,N_28789);
or UO_2831 (O_2831,N_29437,N_29947);
nand UO_2832 (O_2832,N_29890,N_29757);
xnor UO_2833 (O_2833,N_29190,N_29515);
xor UO_2834 (O_2834,N_29719,N_29977);
xor UO_2835 (O_2835,N_28755,N_29613);
nand UO_2836 (O_2836,N_28646,N_29213);
or UO_2837 (O_2837,N_29423,N_29927);
nor UO_2838 (O_2838,N_29833,N_29829);
nand UO_2839 (O_2839,N_28669,N_29116);
nand UO_2840 (O_2840,N_29808,N_28571);
nand UO_2841 (O_2841,N_29767,N_28693);
nor UO_2842 (O_2842,N_28653,N_29431);
and UO_2843 (O_2843,N_29257,N_28529);
nand UO_2844 (O_2844,N_28520,N_28990);
nor UO_2845 (O_2845,N_29955,N_29316);
xor UO_2846 (O_2846,N_29999,N_28913);
and UO_2847 (O_2847,N_29580,N_29435);
xnor UO_2848 (O_2848,N_29236,N_28837);
nor UO_2849 (O_2849,N_28990,N_29614);
and UO_2850 (O_2850,N_28700,N_29038);
or UO_2851 (O_2851,N_29668,N_29261);
nand UO_2852 (O_2852,N_29910,N_28764);
nand UO_2853 (O_2853,N_28805,N_29694);
xor UO_2854 (O_2854,N_29473,N_29684);
nor UO_2855 (O_2855,N_29004,N_28682);
xor UO_2856 (O_2856,N_29794,N_29480);
xor UO_2857 (O_2857,N_29908,N_28645);
nand UO_2858 (O_2858,N_28584,N_28903);
nor UO_2859 (O_2859,N_29415,N_29366);
or UO_2860 (O_2860,N_28887,N_29357);
xor UO_2861 (O_2861,N_28670,N_28688);
or UO_2862 (O_2862,N_29812,N_28955);
xnor UO_2863 (O_2863,N_29954,N_29730);
xor UO_2864 (O_2864,N_29783,N_29008);
xor UO_2865 (O_2865,N_29538,N_29032);
and UO_2866 (O_2866,N_28976,N_29452);
or UO_2867 (O_2867,N_28985,N_29519);
xnor UO_2868 (O_2868,N_29213,N_29360);
and UO_2869 (O_2869,N_29116,N_28626);
or UO_2870 (O_2870,N_29851,N_29496);
nand UO_2871 (O_2871,N_29402,N_29071);
or UO_2872 (O_2872,N_29802,N_29220);
nor UO_2873 (O_2873,N_29554,N_28646);
and UO_2874 (O_2874,N_29080,N_28966);
nor UO_2875 (O_2875,N_29913,N_29945);
or UO_2876 (O_2876,N_28711,N_29902);
xor UO_2877 (O_2877,N_29440,N_28918);
and UO_2878 (O_2878,N_29737,N_29018);
or UO_2879 (O_2879,N_29329,N_28523);
nand UO_2880 (O_2880,N_29820,N_29246);
nand UO_2881 (O_2881,N_29534,N_28633);
or UO_2882 (O_2882,N_28807,N_29077);
nor UO_2883 (O_2883,N_29026,N_29335);
or UO_2884 (O_2884,N_28961,N_29117);
nand UO_2885 (O_2885,N_29736,N_29456);
and UO_2886 (O_2886,N_28625,N_29284);
xor UO_2887 (O_2887,N_29016,N_29604);
xnor UO_2888 (O_2888,N_29637,N_28704);
nand UO_2889 (O_2889,N_28594,N_28982);
and UO_2890 (O_2890,N_29886,N_29075);
and UO_2891 (O_2891,N_29375,N_29161);
nor UO_2892 (O_2892,N_28727,N_29482);
and UO_2893 (O_2893,N_29308,N_29438);
and UO_2894 (O_2894,N_28928,N_28778);
xnor UO_2895 (O_2895,N_29000,N_29277);
xnor UO_2896 (O_2896,N_28990,N_29115);
or UO_2897 (O_2897,N_28653,N_29300);
nor UO_2898 (O_2898,N_29417,N_29222);
nand UO_2899 (O_2899,N_28941,N_29011);
and UO_2900 (O_2900,N_29220,N_28579);
and UO_2901 (O_2901,N_29914,N_28666);
and UO_2902 (O_2902,N_29633,N_29623);
nor UO_2903 (O_2903,N_29035,N_28542);
and UO_2904 (O_2904,N_28760,N_28652);
xor UO_2905 (O_2905,N_28730,N_29445);
xnor UO_2906 (O_2906,N_29074,N_29159);
nor UO_2907 (O_2907,N_29662,N_29778);
nand UO_2908 (O_2908,N_29894,N_29712);
and UO_2909 (O_2909,N_29681,N_29176);
nand UO_2910 (O_2910,N_28974,N_29275);
and UO_2911 (O_2911,N_29520,N_28917);
nand UO_2912 (O_2912,N_28720,N_28672);
xor UO_2913 (O_2913,N_28624,N_29592);
xor UO_2914 (O_2914,N_29615,N_29863);
nand UO_2915 (O_2915,N_29790,N_29582);
or UO_2916 (O_2916,N_28514,N_28930);
and UO_2917 (O_2917,N_28891,N_29651);
xor UO_2918 (O_2918,N_29427,N_29805);
xor UO_2919 (O_2919,N_29887,N_29764);
xor UO_2920 (O_2920,N_29939,N_29127);
and UO_2921 (O_2921,N_28873,N_29185);
or UO_2922 (O_2922,N_29149,N_29682);
and UO_2923 (O_2923,N_28693,N_29762);
nor UO_2924 (O_2924,N_29763,N_28889);
or UO_2925 (O_2925,N_29861,N_29463);
xor UO_2926 (O_2926,N_29945,N_29625);
xor UO_2927 (O_2927,N_28902,N_29803);
or UO_2928 (O_2928,N_28909,N_29146);
and UO_2929 (O_2929,N_28829,N_28936);
and UO_2930 (O_2930,N_28510,N_29155);
and UO_2931 (O_2931,N_29990,N_29583);
or UO_2932 (O_2932,N_29655,N_29500);
nor UO_2933 (O_2933,N_29199,N_28786);
nand UO_2934 (O_2934,N_28645,N_29670);
nor UO_2935 (O_2935,N_28936,N_29113);
and UO_2936 (O_2936,N_29753,N_28901);
nand UO_2937 (O_2937,N_29141,N_29145);
and UO_2938 (O_2938,N_29634,N_29768);
or UO_2939 (O_2939,N_29114,N_29734);
and UO_2940 (O_2940,N_29187,N_29497);
nor UO_2941 (O_2941,N_29714,N_29245);
or UO_2942 (O_2942,N_29297,N_28704);
and UO_2943 (O_2943,N_29109,N_29074);
nand UO_2944 (O_2944,N_29402,N_28757);
nand UO_2945 (O_2945,N_29934,N_28817);
nor UO_2946 (O_2946,N_28883,N_29159);
or UO_2947 (O_2947,N_28935,N_28548);
nand UO_2948 (O_2948,N_29925,N_29212);
nand UO_2949 (O_2949,N_29537,N_28918);
xnor UO_2950 (O_2950,N_28808,N_29894);
or UO_2951 (O_2951,N_29609,N_28782);
or UO_2952 (O_2952,N_28748,N_28928);
or UO_2953 (O_2953,N_28806,N_29026);
nor UO_2954 (O_2954,N_29363,N_28554);
nor UO_2955 (O_2955,N_29859,N_29069);
xnor UO_2956 (O_2956,N_29749,N_29319);
nor UO_2957 (O_2957,N_29523,N_29965);
or UO_2958 (O_2958,N_29286,N_29659);
or UO_2959 (O_2959,N_29259,N_29406);
nor UO_2960 (O_2960,N_29864,N_29066);
nand UO_2961 (O_2961,N_29500,N_28503);
nand UO_2962 (O_2962,N_28950,N_29432);
nand UO_2963 (O_2963,N_28514,N_28979);
xor UO_2964 (O_2964,N_28858,N_28855);
nor UO_2965 (O_2965,N_29036,N_28734);
and UO_2966 (O_2966,N_29038,N_28595);
or UO_2967 (O_2967,N_28831,N_28815);
xor UO_2968 (O_2968,N_29806,N_28694);
nand UO_2969 (O_2969,N_29061,N_28853);
and UO_2970 (O_2970,N_29508,N_29477);
and UO_2971 (O_2971,N_29462,N_29485);
nand UO_2972 (O_2972,N_29143,N_28720);
and UO_2973 (O_2973,N_29555,N_29010);
and UO_2974 (O_2974,N_29126,N_29647);
or UO_2975 (O_2975,N_29823,N_29401);
and UO_2976 (O_2976,N_29651,N_29364);
and UO_2977 (O_2977,N_28813,N_29505);
nor UO_2978 (O_2978,N_29238,N_29704);
nor UO_2979 (O_2979,N_28693,N_28818);
and UO_2980 (O_2980,N_29200,N_29334);
or UO_2981 (O_2981,N_29260,N_29064);
nor UO_2982 (O_2982,N_28886,N_29998);
nor UO_2983 (O_2983,N_29693,N_29034);
xnor UO_2984 (O_2984,N_29615,N_29770);
or UO_2985 (O_2985,N_28648,N_29074);
nand UO_2986 (O_2986,N_28692,N_29972);
or UO_2987 (O_2987,N_29073,N_29133);
and UO_2988 (O_2988,N_28971,N_29090);
and UO_2989 (O_2989,N_29519,N_29515);
nor UO_2990 (O_2990,N_29345,N_29791);
and UO_2991 (O_2991,N_29737,N_28669);
or UO_2992 (O_2992,N_29322,N_29254);
nand UO_2993 (O_2993,N_29198,N_29612);
and UO_2994 (O_2994,N_29469,N_29639);
nor UO_2995 (O_2995,N_28716,N_29597);
and UO_2996 (O_2996,N_28559,N_28833);
and UO_2997 (O_2997,N_28801,N_28813);
and UO_2998 (O_2998,N_29637,N_29232);
and UO_2999 (O_2999,N_29765,N_29388);
xor UO_3000 (O_3000,N_28729,N_28758);
or UO_3001 (O_3001,N_28624,N_29805);
or UO_3002 (O_3002,N_29517,N_28803);
nor UO_3003 (O_3003,N_28962,N_29629);
nor UO_3004 (O_3004,N_29785,N_29620);
xor UO_3005 (O_3005,N_28894,N_29001);
nor UO_3006 (O_3006,N_29338,N_28893);
or UO_3007 (O_3007,N_29889,N_29461);
xnor UO_3008 (O_3008,N_28830,N_29319);
nor UO_3009 (O_3009,N_29536,N_29333);
xnor UO_3010 (O_3010,N_29167,N_29324);
xor UO_3011 (O_3011,N_29045,N_29449);
nand UO_3012 (O_3012,N_29025,N_28668);
nor UO_3013 (O_3013,N_28525,N_29433);
nand UO_3014 (O_3014,N_29731,N_28709);
xnor UO_3015 (O_3015,N_29259,N_29866);
or UO_3016 (O_3016,N_29734,N_29249);
nand UO_3017 (O_3017,N_29123,N_29015);
nand UO_3018 (O_3018,N_28580,N_29241);
or UO_3019 (O_3019,N_29546,N_28787);
nor UO_3020 (O_3020,N_29816,N_29670);
nand UO_3021 (O_3021,N_28623,N_28773);
xnor UO_3022 (O_3022,N_29153,N_28573);
nor UO_3023 (O_3023,N_29660,N_29824);
nor UO_3024 (O_3024,N_29762,N_29976);
xnor UO_3025 (O_3025,N_29203,N_28818);
or UO_3026 (O_3026,N_29575,N_29730);
nand UO_3027 (O_3027,N_28517,N_28571);
or UO_3028 (O_3028,N_29432,N_29061);
nand UO_3029 (O_3029,N_28712,N_29040);
nand UO_3030 (O_3030,N_29446,N_29321);
nor UO_3031 (O_3031,N_29993,N_28794);
and UO_3032 (O_3032,N_28568,N_29251);
nand UO_3033 (O_3033,N_29672,N_28844);
nor UO_3034 (O_3034,N_29078,N_29378);
xor UO_3035 (O_3035,N_29063,N_28831);
or UO_3036 (O_3036,N_29412,N_29670);
xnor UO_3037 (O_3037,N_29893,N_29058);
nand UO_3038 (O_3038,N_29262,N_28807);
and UO_3039 (O_3039,N_28515,N_29457);
or UO_3040 (O_3040,N_28613,N_29020);
xor UO_3041 (O_3041,N_29794,N_29027);
nand UO_3042 (O_3042,N_29511,N_28912);
or UO_3043 (O_3043,N_29689,N_29743);
nand UO_3044 (O_3044,N_29829,N_28657);
xnor UO_3045 (O_3045,N_29147,N_29569);
or UO_3046 (O_3046,N_29377,N_29485);
nand UO_3047 (O_3047,N_29396,N_28771);
or UO_3048 (O_3048,N_29563,N_28759);
nor UO_3049 (O_3049,N_29239,N_28973);
xor UO_3050 (O_3050,N_29405,N_29298);
and UO_3051 (O_3051,N_29369,N_29400);
or UO_3052 (O_3052,N_28794,N_29441);
xnor UO_3053 (O_3053,N_28505,N_29623);
or UO_3054 (O_3054,N_29468,N_28517);
nor UO_3055 (O_3055,N_29236,N_29121);
nand UO_3056 (O_3056,N_29605,N_29074);
nor UO_3057 (O_3057,N_29410,N_29727);
nor UO_3058 (O_3058,N_29683,N_28529);
or UO_3059 (O_3059,N_28893,N_29955);
and UO_3060 (O_3060,N_28648,N_29924);
or UO_3061 (O_3061,N_29802,N_29125);
xor UO_3062 (O_3062,N_29501,N_29595);
nor UO_3063 (O_3063,N_29954,N_28906);
nor UO_3064 (O_3064,N_28643,N_29363);
nand UO_3065 (O_3065,N_28609,N_28800);
nand UO_3066 (O_3066,N_29546,N_29039);
nand UO_3067 (O_3067,N_28972,N_28699);
nor UO_3068 (O_3068,N_28571,N_28520);
xnor UO_3069 (O_3069,N_28635,N_29771);
nor UO_3070 (O_3070,N_29656,N_29374);
nor UO_3071 (O_3071,N_29747,N_29292);
xnor UO_3072 (O_3072,N_29743,N_28501);
and UO_3073 (O_3073,N_28716,N_29729);
nor UO_3074 (O_3074,N_28723,N_29901);
and UO_3075 (O_3075,N_28574,N_29419);
nand UO_3076 (O_3076,N_28586,N_29065);
xor UO_3077 (O_3077,N_29720,N_29677);
xor UO_3078 (O_3078,N_29401,N_29951);
nor UO_3079 (O_3079,N_29130,N_29978);
and UO_3080 (O_3080,N_28781,N_28854);
and UO_3081 (O_3081,N_28519,N_29159);
or UO_3082 (O_3082,N_29437,N_29494);
or UO_3083 (O_3083,N_29306,N_29531);
xnor UO_3084 (O_3084,N_29317,N_29625);
nor UO_3085 (O_3085,N_29404,N_29336);
and UO_3086 (O_3086,N_29970,N_29324);
nand UO_3087 (O_3087,N_29738,N_28515);
nor UO_3088 (O_3088,N_29480,N_29729);
xnor UO_3089 (O_3089,N_28654,N_28799);
nor UO_3090 (O_3090,N_29945,N_29571);
or UO_3091 (O_3091,N_29674,N_29767);
nand UO_3092 (O_3092,N_29856,N_29273);
or UO_3093 (O_3093,N_29765,N_29977);
or UO_3094 (O_3094,N_29812,N_29661);
or UO_3095 (O_3095,N_29757,N_29595);
or UO_3096 (O_3096,N_29291,N_28555);
and UO_3097 (O_3097,N_29420,N_28912);
and UO_3098 (O_3098,N_29882,N_28824);
nor UO_3099 (O_3099,N_29549,N_29201);
and UO_3100 (O_3100,N_29782,N_29842);
and UO_3101 (O_3101,N_28908,N_28877);
or UO_3102 (O_3102,N_29258,N_29769);
and UO_3103 (O_3103,N_29339,N_29909);
and UO_3104 (O_3104,N_29569,N_28500);
nor UO_3105 (O_3105,N_28980,N_29821);
nor UO_3106 (O_3106,N_28588,N_28591);
and UO_3107 (O_3107,N_28879,N_28677);
nor UO_3108 (O_3108,N_29246,N_29666);
or UO_3109 (O_3109,N_28547,N_28565);
nand UO_3110 (O_3110,N_29876,N_29180);
nor UO_3111 (O_3111,N_29361,N_29804);
nor UO_3112 (O_3112,N_29424,N_29502);
nor UO_3113 (O_3113,N_29507,N_29877);
nand UO_3114 (O_3114,N_29455,N_28807);
nor UO_3115 (O_3115,N_29216,N_28817);
nor UO_3116 (O_3116,N_28519,N_28848);
or UO_3117 (O_3117,N_29074,N_28819);
xor UO_3118 (O_3118,N_28603,N_28785);
nand UO_3119 (O_3119,N_28659,N_28526);
xnor UO_3120 (O_3120,N_29779,N_29155);
and UO_3121 (O_3121,N_29508,N_28971);
xor UO_3122 (O_3122,N_29033,N_29814);
or UO_3123 (O_3123,N_29514,N_29745);
nand UO_3124 (O_3124,N_28674,N_29497);
nand UO_3125 (O_3125,N_29629,N_29909);
xor UO_3126 (O_3126,N_28911,N_29519);
or UO_3127 (O_3127,N_28569,N_29323);
or UO_3128 (O_3128,N_28672,N_29650);
or UO_3129 (O_3129,N_28623,N_29924);
nand UO_3130 (O_3130,N_29395,N_29430);
nor UO_3131 (O_3131,N_28710,N_29400);
nand UO_3132 (O_3132,N_29983,N_29791);
nand UO_3133 (O_3133,N_29355,N_29138);
nand UO_3134 (O_3134,N_28587,N_29355);
nand UO_3135 (O_3135,N_29453,N_29309);
and UO_3136 (O_3136,N_29418,N_28680);
xor UO_3137 (O_3137,N_29564,N_29309);
xnor UO_3138 (O_3138,N_28915,N_29578);
nor UO_3139 (O_3139,N_29894,N_29384);
and UO_3140 (O_3140,N_29679,N_29641);
nand UO_3141 (O_3141,N_29138,N_29430);
nor UO_3142 (O_3142,N_29995,N_28787);
nand UO_3143 (O_3143,N_29033,N_28569);
xor UO_3144 (O_3144,N_29177,N_29903);
or UO_3145 (O_3145,N_29009,N_28680);
nand UO_3146 (O_3146,N_29728,N_29479);
xor UO_3147 (O_3147,N_28657,N_28842);
nor UO_3148 (O_3148,N_29699,N_28714);
xnor UO_3149 (O_3149,N_29891,N_28637);
or UO_3150 (O_3150,N_28857,N_28949);
and UO_3151 (O_3151,N_29120,N_29738);
nor UO_3152 (O_3152,N_29194,N_29560);
xnor UO_3153 (O_3153,N_29141,N_29062);
nand UO_3154 (O_3154,N_29521,N_29715);
xor UO_3155 (O_3155,N_29819,N_28647);
nor UO_3156 (O_3156,N_28652,N_29025);
or UO_3157 (O_3157,N_28550,N_29253);
and UO_3158 (O_3158,N_29593,N_29702);
or UO_3159 (O_3159,N_29680,N_29297);
and UO_3160 (O_3160,N_29957,N_29892);
xor UO_3161 (O_3161,N_29180,N_29881);
nand UO_3162 (O_3162,N_29273,N_28519);
and UO_3163 (O_3163,N_29137,N_29387);
nor UO_3164 (O_3164,N_29426,N_29052);
and UO_3165 (O_3165,N_29536,N_29361);
nor UO_3166 (O_3166,N_29425,N_28895);
and UO_3167 (O_3167,N_29120,N_28545);
or UO_3168 (O_3168,N_29693,N_29464);
and UO_3169 (O_3169,N_29428,N_29250);
nor UO_3170 (O_3170,N_29029,N_29713);
nor UO_3171 (O_3171,N_28569,N_29812);
nand UO_3172 (O_3172,N_28891,N_28809);
or UO_3173 (O_3173,N_29619,N_28876);
nand UO_3174 (O_3174,N_29359,N_28765);
or UO_3175 (O_3175,N_29182,N_29128);
and UO_3176 (O_3176,N_28704,N_29609);
or UO_3177 (O_3177,N_29854,N_29709);
nand UO_3178 (O_3178,N_28974,N_29071);
nand UO_3179 (O_3179,N_29688,N_29986);
nand UO_3180 (O_3180,N_29943,N_28525);
or UO_3181 (O_3181,N_29830,N_29486);
nand UO_3182 (O_3182,N_29254,N_28762);
nor UO_3183 (O_3183,N_28833,N_28808);
nor UO_3184 (O_3184,N_29881,N_29349);
xnor UO_3185 (O_3185,N_29293,N_29104);
or UO_3186 (O_3186,N_29271,N_29334);
xnor UO_3187 (O_3187,N_29954,N_29754);
xnor UO_3188 (O_3188,N_29368,N_29225);
nand UO_3189 (O_3189,N_28516,N_28965);
or UO_3190 (O_3190,N_29579,N_28806);
nand UO_3191 (O_3191,N_28551,N_29450);
nand UO_3192 (O_3192,N_28743,N_28856);
and UO_3193 (O_3193,N_29894,N_29486);
nor UO_3194 (O_3194,N_29293,N_29560);
and UO_3195 (O_3195,N_29117,N_29655);
xnor UO_3196 (O_3196,N_28907,N_29120);
nand UO_3197 (O_3197,N_28603,N_29906);
nor UO_3198 (O_3198,N_28544,N_29353);
or UO_3199 (O_3199,N_29782,N_28619);
nand UO_3200 (O_3200,N_28953,N_28886);
nand UO_3201 (O_3201,N_29244,N_28720);
or UO_3202 (O_3202,N_29975,N_29933);
nand UO_3203 (O_3203,N_28915,N_29172);
and UO_3204 (O_3204,N_29570,N_29944);
or UO_3205 (O_3205,N_28539,N_28715);
or UO_3206 (O_3206,N_29693,N_29729);
nor UO_3207 (O_3207,N_28522,N_29066);
and UO_3208 (O_3208,N_29789,N_28859);
and UO_3209 (O_3209,N_28553,N_29876);
nand UO_3210 (O_3210,N_29440,N_29982);
xnor UO_3211 (O_3211,N_28581,N_29278);
xor UO_3212 (O_3212,N_28851,N_29487);
nor UO_3213 (O_3213,N_28550,N_28721);
xnor UO_3214 (O_3214,N_28969,N_29045);
or UO_3215 (O_3215,N_29390,N_29202);
nor UO_3216 (O_3216,N_28636,N_29378);
nor UO_3217 (O_3217,N_28722,N_29392);
nand UO_3218 (O_3218,N_29912,N_29979);
and UO_3219 (O_3219,N_29201,N_28797);
and UO_3220 (O_3220,N_29560,N_29978);
or UO_3221 (O_3221,N_29873,N_28629);
nor UO_3222 (O_3222,N_29044,N_28716);
xor UO_3223 (O_3223,N_29631,N_28688);
or UO_3224 (O_3224,N_29953,N_29455);
xor UO_3225 (O_3225,N_29478,N_28890);
and UO_3226 (O_3226,N_28567,N_29184);
or UO_3227 (O_3227,N_28688,N_29254);
and UO_3228 (O_3228,N_29345,N_29338);
xnor UO_3229 (O_3229,N_29799,N_29656);
nor UO_3230 (O_3230,N_29089,N_28941);
or UO_3231 (O_3231,N_29103,N_28531);
or UO_3232 (O_3232,N_28559,N_29945);
nor UO_3233 (O_3233,N_28722,N_29875);
or UO_3234 (O_3234,N_29479,N_29511);
nand UO_3235 (O_3235,N_29558,N_29812);
nand UO_3236 (O_3236,N_29279,N_29394);
or UO_3237 (O_3237,N_29066,N_29365);
or UO_3238 (O_3238,N_29615,N_29614);
and UO_3239 (O_3239,N_28932,N_28523);
xnor UO_3240 (O_3240,N_29932,N_29567);
nand UO_3241 (O_3241,N_28932,N_28622);
nand UO_3242 (O_3242,N_29720,N_29949);
nand UO_3243 (O_3243,N_28652,N_29795);
nand UO_3244 (O_3244,N_29542,N_29861);
or UO_3245 (O_3245,N_29227,N_28997);
nand UO_3246 (O_3246,N_29631,N_29229);
nand UO_3247 (O_3247,N_29387,N_29805);
and UO_3248 (O_3248,N_29670,N_29550);
or UO_3249 (O_3249,N_28603,N_29022);
nor UO_3250 (O_3250,N_28707,N_29968);
nand UO_3251 (O_3251,N_29726,N_29021);
nand UO_3252 (O_3252,N_28617,N_28745);
or UO_3253 (O_3253,N_29283,N_29363);
nor UO_3254 (O_3254,N_29949,N_28619);
nand UO_3255 (O_3255,N_29589,N_29633);
nor UO_3256 (O_3256,N_29060,N_28725);
nand UO_3257 (O_3257,N_29398,N_29039);
nor UO_3258 (O_3258,N_29271,N_28652);
nand UO_3259 (O_3259,N_29236,N_29565);
or UO_3260 (O_3260,N_29541,N_28681);
xnor UO_3261 (O_3261,N_29881,N_28646);
and UO_3262 (O_3262,N_28603,N_29522);
or UO_3263 (O_3263,N_29696,N_29463);
and UO_3264 (O_3264,N_28557,N_28704);
nand UO_3265 (O_3265,N_28993,N_29921);
nand UO_3266 (O_3266,N_28605,N_28954);
and UO_3267 (O_3267,N_29730,N_29378);
xnor UO_3268 (O_3268,N_29115,N_28773);
and UO_3269 (O_3269,N_29649,N_29469);
nand UO_3270 (O_3270,N_29978,N_29598);
xor UO_3271 (O_3271,N_29221,N_29799);
nand UO_3272 (O_3272,N_29405,N_29110);
and UO_3273 (O_3273,N_29032,N_29829);
xor UO_3274 (O_3274,N_29790,N_29437);
and UO_3275 (O_3275,N_29331,N_29904);
nor UO_3276 (O_3276,N_28807,N_28540);
xor UO_3277 (O_3277,N_28692,N_28597);
or UO_3278 (O_3278,N_28572,N_28889);
nand UO_3279 (O_3279,N_29934,N_29595);
and UO_3280 (O_3280,N_28685,N_29049);
nor UO_3281 (O_3281,N_28717,N_29247);
nor UO_3282 (O_3282,N_29276,N_29424);
or UO_3283 (O_3283,N_29827,N_29454);
xor UO_3284 (O_3284,N_28980,N_29642);
nand UO_3285 (O_3285,N_28770,N_29261);
or UO_3286 (O_3286,N_29820,N_29830);
or UO_3287 (O_3287,N_28898,N_28561);
nor UO_3288 (O_3288,N_29789,N_28828);
and UO_3289 (O_3289,N_28686,N_29416);
nor UO_3290 (O_3290,N_28566,N_29382);
nand UO_3291 (O_3291,N_29759,N_29182);
or UO_3292 (O_3292,N_29077,N_28867);
or UO_3293 (O_3293,N_29715,N_28575);
nand UO_3294 (O_3294,N_29984,N_29425);
xor UO_3295 (O_3295,N_28894,N_28507);
and UO_3296 (O_3296,N_29872,N_29091);
nor UO_3297 (O_3297,N_29301,N_28514);
nand UO_3298 (O_3298,N_28889,N_29978);
or UO_3299 (O_3299,N_29410,N_29955);
or UO_3300 (O_3300,N_28728,N_29520);
and UO_3301 (O_3301,N_29315,N_29837);
or UO_3302 (O_3302,N_29449,N_29074);
nor UO_3303 (O_3303,N_29764,N_29885);
nand UO_3304 (O_3304,N_28841,N_29969);
nor UO_3305 (O_3305,N_29761,N_29910);
and UO_3306 (O_3306,N_28803,N_29974);
xnor UO_3307 (O_3307,N_28782,N_29257);
and UO_3308 (O_3308,N_29731,N_29388);
and UO_3309 (O_3309,N_29172,N_29023);
or UO_3310 (O_3310,N_29782,N_29667);
nor UO_3311 (O_3311,N_28577,N_29091);
nor UO_3312 (O_3312,N_28729,N_29869);
or UO_3313 (O_3313,N_29634,N_29642);
or UO_3314 (O_3314,N_28745,N_29139);
xnor UO_3315 (O_3315,N_29194,N_28954);
xor UO_3316 (O_3316,N_29327,N_29958);
xnor UO_3317 (O_3317,N_29746,N_28755);
nor UO_3318 (O_3318,N_29545,N_28594);
nor UO_3319 (O_3319,N_28947,N_29586);
nor UO_3320 (O_3320,N_28615,N_29477);
or UO_3321 (O_3321,N_29728,N_28582);
and UO_3322 (O_3322,N_29305,N_29565);
and UO_3323 (O_3323,N_28965,N_28624);
or UO_3324 (O_3324,N_29416,N_29351);
nand UO_3325 (O_3325,N_29749,N_29553);
or UO_3326 (O_3326,N_28600,N_28655);
xor UO_3327 (O_3327,N_29333,N_28601);
nor UO_3328 (O_3328,N_28652,N_29399);
or UO_3329 (O_3329,N_28509,N_28945);
nand UO_3330 (O_3330,N_29931,N_29502);
nor UO_3331 (O_3331,N_29675,N_28998);
nor UO_3332 (O_3332,N_29463,N_28571);
and UO_3333 (O_3333,N_29483,N_28907);
xnor UO_3334 (O_3334,N_29115,N_29928);
or UO_3335 (O_3335,N_28552,N_29000);
nor UO_3336 (O_3336,N_29171,N_29643);
nor UO_3337 (O_3337,N_28810,N_28969);
xnor UO_3338 (O_3338,N_29072,N_29164);
or UO_3339 (O_3339,N_28856,N_28835);
or UO_3340 (O_3340,N_28857,N_29127);
nand UO_3341 (O_3341,N_28524,N_29077);
nand UO_3342 (O_3342,N_29277,N_28690);
nor UO_3343 (O_3343,N_29155,N_29253);
and UO_3344 (O_3344,N_29111,N_28911);
xnor UO_3345 (O_3345,N_29952,N_28826);
or UO_3346 (O_3346,N_28895,N_29043);
or UO_3347 (O_3347,N_28507,N_29377);
xor UO_3348 (O_3348,N_29171,N_29722);
xor UO_3349 (O_3349,N_29233,N_29414);
and UO_3350 (O_3350,N_29424,N_28613);
and UO_3351 (O_3351,N_28655,N_29491);
nand UO_3352 (O_3352,N_28654,N_28818);
nor UO_3353 (O_3353,N_28821,N_29499);
nand UO_3354 (O_3354,N_29644,N_28955);
nor UO_3355 (O_3355,N_28697,N_28910);
or UO_3356 (O_3356,N_29001,N_29922);
nand UO_3357 (O_3357,N_29900,N_29564);
and UO_3358 (O_3358,N_29574,N_28635);
nor UO_3359 (O_3359,N_29519,N_29438);
or UO_3360 (O_3360,N_29075,N_28799);
nand UO_3361 (O_3361,N_29211,N_28896);
and UO_3362 (O_3362,N_29601,N_29140);
or UO_3363 (O_3363,N_29704,N_29960);
and UO_3364 (O_3364,N_28839,N_29015);
and UO_3365 (O_3365,N_28851,N_28861);
xor UO_3366 (O_3366,N_28765,N_29040);
or UO_3367 (O_3367,N_29721,N_29915);
nand UO_3368 (O_3368,N_29112,N_29360);
and UO_3369 (O_3369,N_28729,N_28627);
nand UO_3370 (O_3370,N_29327,N_28745);
nor UO_3371 (O_3371,N_28527,N_29727);
nand UO_3372 (O_3372,N_28969,N_29654);
and UO_3373 (O_3373,N_29355,N_28799);
xor UO_3374 (O_3374,N_29464,N_29399);
nand UO_3375 (O_3375,N_29984,N_29545);
nor UO_3376 (O_3376,N_28802,N_29288);
or UO_3377 (O_3377,N_29215,N_28809);
or UO_3378 (O_3378,N_28542,N_29743);
nor UO_3379 (O_3379,N_29153,N_28624);
or UO_3380 (O_3380,N_29832,N_29152);
or UO_3381 (O_3381,N_29913,N_28626);
and UO_3382 (O_3382,N_29804,N_28527);
or UO_3383 (O_3383,N_29764,N_28755);
xor UO_3384 (O_3384,N_28528,N_29597);
and UO_3385 (O_3385,N_29476,N_28577);
nor UO_3386 (O_3386,N_29518,N_29689);
nand UO_3387 (O_3387,N_29959,N_29494);
nor UO_3388 (O_3388,N_28864,N_29762);
nand UO_3389 (O_3389,N_29390,N_28814);
and UO_3390 (O_3390,N_28618,N_28995);
nor UO_3391 (O_3391,N_29188,N_29551);
nand UO_3392 (O_3392,N_28579,N_29771);
nor UO_3393 (O_3393,N_28629,N_28706);
and UO_3394 (O_3394,N_29549,N_29647);
nor UO_3395 (O_3395,N_29774,N_29316);
nor UO_3396 (O_3396,N_29353,N_28998);
nor UO_3397 (O_3397,N_28850,N_29099);
and UO_3398 (O_3398,N_29268,N_28566);
or UO_3399 (O_3399,N_29268,N_29411);
nor UO_3400 (O_3400,N_29371,N_29937);
nand UO_3401 (O_3401,N_28975,N_29998);
nand UO_3402 (O_3402,N_28823,N_28552);
nor UO_3403 (O_3403,N_28840,N_29640);
or UO_3404 (O_3404,N_29994,N_29251);
xnor UO_3405 (O_3405,N_29443,N_29848);
nand UO_3406 (O_3406,N_29496,N_29383);
or UO_3407 (O_3407,N_29991,N_28776);
or UO_3408 (O_3408,N_29162,N_29657);
xnor UO_3409 (O_3409,N_28834,N_29285);
xor UO_3410 (O_3410,N_29278,N_28924);
nor UO_3411 (O_3411,N_29243,N_29104);
nor UO_3412 (O_3412,N_29736,N_29300);
nor UO_3413 (O_3413,N_28716,N_28628);
nor UO_3414 (O_3414,N_28679,N_29928);
or UO_3415 (O_3415,N_28818,N_28876);
or UO_3416 (O_3416,N_29945,N_29148);
xor UO_3417 (O_3417,N_29848,N_29705);
and UO_3418 (O_3418,N_29564,N_29795);
nand UO_3419 (O_3419,N_28836,N_28692);
nor UO_3420 (O_3420,N_28843,N_29530);
xor UO_3421 (O_3421,N_28714,N_29592);
and UO_3422 (O_3422,N_29122,N_29158);
nand UO_3423 (O_3423,N_29912,N_29598);
nor UO_3424 (O_3424,N_29421,N_29234);
xor UO_3425 (O_3425,N_29495,N_28678);
xnor UO_3426 (O_3426,N_29735,N_29950);
nand UO_3427 (O_3427,N_29931,N_29151);
nor UO_3428 (O_3428,N_29242,N_29962);
xor UO_3429 (O_3429,N_29941,N_29312);
nor UO_3430 (O_3430,N_28847,N_28925);
nor UO_3431 (O_3431,N_29797,N_29763);
xor UO_3432 (O_3432,N_29532,N_28662);
xor UO_3433 (O_3433,N_28625,N_28831);
or UO_3434 (O_3434,N_28890,N_29998);
or UO_3435 (O_3435,N_29463,N_29552);
nor UO_3436 (O_3436,N_28707,N_28859);
xnor UO_3437 (O_3437,N_28513,N_29686);
nand UO_3438 (O_3438,N_28668,N_28623);
nor UO_3439 (O_3439,N_29310,N_29399);
nor UO_3440 (O_3440,N_29032,N_29222);
and UO_3441 (O_3441,N_29669,N_29955);
nor UO_3442 (O_3442,N_29483,N_28968);
or UO_3443 (O_3443,N_29235,N_29843);
and UO_3444 (O_3444,N_28713,N_29100);
xnor UO_3445 (O_3445,N_29236,N_28576);
and UO_3446 (O_3446,N_28829,N_28891);
nor UO_3447 (O_3447,N_28673,N_29493);
xnor UO_3448 (O_3448,N_28925,N_28942);
nor UO_3449 (O_3449,N_28633,N_28649);
nand UO_3450 (O_3450,N_29480,N_28517);
or UO_3451 (O_3451,N_29993,N_29138);
and UO_3452 (O_3452,N_28867,N_29262);
xor UO_3453 (O_3453,N_29040,N_29785);
xor UO_3454 (O_3454,N_28644,N_29391);
nand UO_3455 (O_3455,N_28562,N_29183);
nand UO_3456 (O_3456,N_28983,N_29346);
and UO_3457 (O_3457,N_29982,N_29996);
xnor UO_3458 (O_3458,N_28977,N_29682);
and UO_3459 (O_3459,N_28761,N_29799);
or UO_3460 (O_3460,N_29066,N_28672);
nor UO_3461 (O_3461,N_29938,N_29443);
and UO_3462 (O_3462,N_29400,N_29734);
and UO_3463 (O_3463,N_29668,N_29878);
and UO_3464 (O_3464,N_29418,N_29964);
and UO_3465 (O_3465,N_28558,N_28913);
xor UO_3466 (O_3466,N_29785,N_29432);
nand UO_3467 (O_3467,N_29484,N_29855);
nand UO_3468 (O_3468,N_29097,N_28959);
nor UO_3469 (O_3469,N_28846,N_28989);
xnor UO_3470 (O_3470,N_29308,N_29706);
nand UO_3471 (O_3471,N_28874,N_29875);
nor UO_3472 (O_3472,N_29918,N_29134);
xor UO_3473 (O_3473,N_28521,N_29726);
and UO_3474 (O_3474,N_29714,N_29340);
nor UO_3475 (O_3475,N_28834,N_28706);
or UO_3476 (O_3476,N_29528,N_29511);
nor UO_3477 (O_3477,N_28649,N_29921);
or UO_3478 (O_3478,N_28929,N_29912);
and UO_3479 (O_3479,N_29418,N_29749);
or UO_3480 (O_3480,N_29488,N_29306);
xor UO_3481 (O_3481,N_29518,N_29935);
xnor UO_3482 (O_3482,N_29935,N_28767);
xor UO_3483 (O_3483,N_28601,N_28932);
and UO_3484 (O_3484,N_29678,N_28985);
nand UO_3485 (O_3485,N_29194,N_28648);
nor UO_3486 (O_3486,N_28891,N_28835);
or UO_3487 (O_3487,N_29558,N_28883);
xor UO_3488 (O_3488,N_29054,N_29495);
nand UO_3489 (O_3489,N_28625,N_29944);
and UO_3490 (O_3490,N_29003,N_29989);
xnor UO_3491 (O_3491,N_29085,N_29972);
or UO_3492 (O_3492,N_29848,N_29548);
nand UO_3493 (O_3493,N_28891,N_28638);
or UO_3494 (O_3494,N_29623,N_29554);
nor UO_3495 (O_3495,N_29438,N_29286);
nor UO_3496 (O_3496,N_29393,N_29281);
nor UO_3497 (O_3497,N_29075,N_29191);
or UO_3498 (O_3498,N_29250,N_29471);
nor UO_3499 (O_3499,N_28804,N_29711);
endmodule