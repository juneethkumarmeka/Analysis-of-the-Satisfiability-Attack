module basic_1000_10000_1500_4_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_71,In_64);
nand U1 (N_1,In_382,In_67);
xnor U2 (N_2,In_190,In_209);
nand U3 (N_3,In_758,In_844);
nand U4 (N_4,In_569,In_250);
xnor U5 (N_5,In_474,In_286);
nand U6 (N_6,In_980,In_682);
nand U7 (N_7,In_867,In_994);
nand U8 (N_8,In_764,In_621);
xor U9 (N_9,In_352,In_907);
and U10 (N_10,In_429,In_582);
and U11 (N_11,In_350,In_399);
xor U12 (N_12,In_44,In_896);
nand U13 (N_13,In_273,In_483);
nor U14 (N_14,In_534,In_501);
nor U15 (N_15,In_365,In_949);
xor U16 (N_16,In_46,In_699);
and U17 (N_17,In_704,In_132);
xnor U18 (N_18,In_99,In_683);
nand U19 (N_19,In_532,In_998);
nand U20 (N_20,In_767,In_301);
or U21 (N_21,In_206,In_517);
nor U22 (N_22,In_351,In_601);
and U23 (N_23,In_289,In_234);
xor U24 (N_24,In_218,In_282);
and U25 (N_25,In_367,In_735);
and U26 (N_26,In_540,In_107);
nor U27 (N_27,In_886,In_82);
or U28 (N_28,In_225,In_748);
and U29 (N_29,In_554,In_463);
nand U30 (N_30,In_586,In_491);
or U31 (N_31,In_130,In_871);
nand U32 (N_32,In_29,In_864);
nand U33 (N_33,In_914,In_470);
nand U34 (N_34,In_556,In_295);
nor U35 (N_35,In_703,In_828);
nand U36 (N_36,In_435,In_428);
xor U37 (N_37,In_387,In_523);
nor U38 (N_38,In_305,In_434);
or U39 (N_39,In_233,In_24);
nor U40 (N_40,In_665,In_698);
xnor U41 (N_41,In_149,In_482);
xor U42 (N_42,In_162,In_159);
or U43 (N_43,In_872,In_814);
and U44 (N_44,In_673,In_507);
xor U45 (N_45,In_430,In_707);
or U46 (N_46,In_50,In_737);
and U47 (N_47,In_216,In_792);
nor U48 (N_48,In_204,In_17);
and U49 (N_49,In_759,In_10);
nor U50 (N_50,In_560,In_808);
and U51 (N_51,In_466,In_404);
or U52 (N_52,In_43,In_617);
and U53 (N_53,In_720,In_300);
xor U54 (N_54,In_761,In_395);
nor U55 (N_55,In_181,In_302);
or U56 (N_56,In_402,In_854);
and U57 (N_57,In_215,In_409);
or U58 (N_58,In_819,In_13);
and U59 (N_59,In_440,In_34);
nand U60 (N_60,In_203,In_857);
and U61 (N_61,In_178,In_228);
nand U62 (N_62,In_311,In_691);
nand U63 (N_63,In_48,In_347);
and U64 (N_64,In_354,In_275);
nor U65 (N_65,In_106,In_661);
xor U66 (N_66,In_655,In_499);
nor U67 (N_67,In_171,In_199);
and U68 (N_68,In_198,In_620);
nand U69 (N_69,In_985,In_238);
or U70 (N_70,In_160,In_913);
xnor U71 (N_71,In_585,In_213);
nand U72 (N_72,In_977,In_739);
xnor U73 (N_73,In_425,In_336);
nor U74 (N_74,In_133,In_342);
xnor U75 (N_75,In_740,In_320);
and U76 (N_76,In_955,In_923);
or U77 (N_77,In_142,In_257);
xnor U78 (N_78,In_32,In_26);
nor U79 (N_79,In_448,In_385);
nand U80 (N_80,In_324,In_960);
or U81 (N_81,In_86,In_235);
or U82 (N_82,In_416,In_115);
and U83 (N_83,In_276,In_578);
xor U84 (N_84,In_627,In_245);
xnor U85 (N_85,In_239,In_150);
and U86 (N_86,In_625,In_990);
or U87 (N_87,In_774,In_91);
xnor U88 (N_88,In_194,In_76);
or U89 (N_89,In_475,In_900);
nand U90 (N_90,In_151,In_653);
xor U91 (N_91,In_614,In_120);
and U92 (N_92,In_974,In_754);
and U93 (N_93,In_542,In_833);
xnor U94 (N_94,In_403,In_810);
or U95 (N_95,In_779,In_495);
nand U96 (N_96,In_35,In_606);
nand U97 (N_97,In_368,In_39);
nor U98 (N_98,In_284,In_340);
nand U99 (N_99,In_846,In_196);
nand U100 (N_100,In_423,In_591);
nand U101 (N_101,In_825,In_244);
xnor U102 (N_102,In_695,In_906);
nor U103 (N_103,In_894,In_714);
and U104 (N_104,In_656,In_877);
nor U105 (N_105,In_467,In_552);
nand U106 (N_106,In_797,In_323);
nand U107 (N_107,In_805,In_161);
and U108 (N_108,In_769,In_663);
and U109 (N_109,In_636,In_826);
and U110 (N_110,In_790,In_885);
nand U111 (N_111,In_644,In_935);
nand U112 (N_112,In_873,In_270);
or U113 (N_113,In_904,In_47);
xor U114 (N_114,In_730,In_392);
xor U115 (N_115,In_638,In_464);
nor U116 (N_116,In_979,In_749);
nor U117 (N_117,In_890,In_148);
and U118 (N_118,In_820,In_381);
or U119 (N_119,In_845,In_796);
nor U120 (N_120,In_237,In_711);
xnor U121 (N_121,In_271,In_917);
nand U122 (N_122,In_94,In_118);
and U123 (N_123,In_415,In_191);
and U124 (N_124,In_874,In_5);
and U125 (N_125,In_603,In_3);
and U126 (N_126,In_478,In_202);
xor U127 (N_127,In_798,In_911);
and U128 (N_128,In_959,In_146);
nand U129 (N_129,In_297,In_229);
or U130 (N_130,In_255,In_861);
xnor U131 (N_131,In_346,In_581);
nand U132 (N_132,In_223,In_593);
and U133 (N_133,In_427,In_398);
and U134 (N_134,In_135,In_875);
xor U135 (N_135,In_200,In_973);
and U136 (N_136,In_667,In_42);
nor U137 (N_137,In_611,In_953);
nor U138 (N_138,In_752,In_948);
and U139 (N_139,In_377,In_530);
nand U140 (N_140,In_144,In_348);
nor U141 (N_141,In_253,In_622);
nor U142 (N_142,In_310,In_224);
and U143 (N_143,In_211,In_545);
and U144 (N_144,In_602,In_38);
or U145 (N_145,In_176,In_131);
nor U146 (N_146,In_480,In_111);
or U147 (N_147,In_139,In_188);
nor U148 (N_148,In_391,In_45);
nand U149 (N_149,In_962,In_443);
or U150 (N_150,In_509,In_81);
and U151 (N_151,In_78,In_956);
and U152 (N_152,In_788,In_497);
or U153 (N_153,In_265,In_127);
and U154 (N_154,In_226,In_88);
nand U155 (N_155,In_950,In_744);
nor U156 (N_156,In_193,In_791);
nand U157 (N_157,In_241,In_596);
or U158 (N_158,In_681,In_256);
and U159 (N_159,In_468,In_794);
xnor U160 (N_160,In_869,In_549);
or U161 (N_161,In_164,In_53);
or U162 (N_162,In_174,In_671);
nand U163 (N_163,In_712,In_353);
or U164 (N_164,In_658,In_941);
and U165 (N_165,In_511,In_702);
xnor U166 (N_166,In_726,In_745);
or U167 (N_167,In_49,In_997);
nand U168 (N_168,In_30,In_325);
nand U169 (N_169,In_855,In_801);
or U170 (N_170,In_701,In_125);
nor U171 (N_171,In_477,In_778);
nand U172 (N_172,In_571,In_982);
xnor U173 (N_173,In_918,In_338);
and U174 (N_174,In_664,In_442);
or U175 (N_175,In_362,In_122);
or U176 (N_176,In_921,In_668);
xor U177 (N_177,In_16,In_274);
or U178 (N_178,In_341,In_946);
or U179 (N_179,In_772,In_167);
xnor U180 (N_180,In_361,In_37);
nand U181 (N_181,In_283,In_709);
nand U182 (N_182,In_232,In_266);
xnor U183 (N_183,In_966,In_77);
and U184 (N_184,In_500,In_597);
and U185 (N_185,In_592,In_938);
or U186 (N_186,In_700,In_628);
nand U187 (N_187,In_105,In_564);
nor U188 (N_188,In_902,In_830);
or U189 (N_189,In_121,In_768);
nand U190 (N_190,In_600,In_944);
nor U191 (N_191,In_880,In_41);
or U192 (N_192,In_901,In_390);
or U193 (N_193,In_568,In_996);
nand U194 (N_194,In_449,In_618);
nor U195 (N_195,In_492,In_780);
nand U196 (N_196,In_108,In_616);
nor U197 (N_197,In_248,In_660);
and U198 (N_198,In_565,In_981);
nor U199 (N_199,In_876,In_74);
nor U200 (N_200,In_456,In_588);
or U201 (N_201,In_531,In_134);
xor U202 (N_202,In_639,In_690);
or U203 (N_203,In_420,In_836);
nand U204 (N_204,In_328,In_558);
nand U205 (N_205,In_623,In_9);
nand U206 (N_206,In_192,In_97);
nand U207 (N_207,In_450,In_84);
nor U208 (N_208,In_786,In_298);
nand U209 (N_209,In_490,In_760);
nand U210 (N_210,In_363,In_789);
or U211 (N_211,In_424,In_782);
and U212 (N_212,In_376,In_612);
nor U213 (N_213,In_165,In_799);
or U214 (N_214,In_129,In_576);
nor U215 (N_215,In_605,In_267);
nor U216 (N_216,In_494,In_73);
nor U217 (N_217,In_718,In_455);
nor U218 (N_218,In_433,In_963);
and U219 (N_219,In_14,In_411);
or U220 (N_220,In_487,In_356);
xor U221 (N_221,In_66,In_460);
xor U222 (N_222,In_680,In_344);
nand U223 (N_223,In_153,In_599);
and U224 (N_224,In_369,In_22);
nand U225 (N_225,In_821,In_303);
or U226 (N_226,In_113,In_169);
xnor U227 (N_227,In_393,In_738);
nor U228 (N_228,In_657,In_197);
and U229 (N_229,In_843,In_945);
nand U230 (N_230,In_514,In_291);
nor U231 (N_231,In_931,In_888);
and U232 (N_232,In_75,In_573);
and U233 (N_233,In_919,In_168);
or U234 (N_234,In_575,In_476);
nor U235 (N_235,In_848,In_230);
or U236 (N_236,In_33,In_781);
xnor U237 (N_237,In_498,In_154);
nor U238 (N_238,In_924,In_529);
xnor U239 (N_239,In_645,In_916);
and U240 (N_240,In_678,In_68);
xnor U241 (N_241,In_526,In_584);
and U242 (N_242,In_555,In_319);
xnor U243 (N_243,In_374,In_227);
and U244 (N_244,In_635,In_626);
and U245 (N_245,In_504,In_992);
xnor U246 (N_246,In_217,In_615);
or U247 (N_247,In_640,In_572);
nand U248 (N_248,In_109,In_832);
xnor U249 (N_249,In_987,In_254);
nor U250 (N_250,In_807,In_776);
xnor U251 (N_251,In_69,In_834);
xnor U252 (N_252,In_418,In_290);
or U253 (N_253,In_307,In_851);
and U254 (N_254,In_706,In_803);
nand U255 (N_255,In_823,In_590);
nand U256 (N_256,In_25,In_243);
nor U257 (N_257,In_662,In_447);
and U258 (N_258,In_63,In_784);
xor U259 (N_259,In_878,In_858);
xnor U260 (N_260,In_991,In_879);
or U261 (N_261,In_143,In_70);
or U262 (N_262,In_141,In_335);
xor U263 (N_263,In_396,In_967);
and U264 (N_264,In_570,In_454);
nor U265 (N_265,In_859,In_471);
and U266 (N_266,In_692,In_686);
nand U267 (N_267,In_54,In_446);
nor U268 (N_268,In_897,In_795);
xor U269 (N_269,In_371,In_370);
nor U270 (N_270,In_158,In_563);
and U271 (N_271,In_296,In_670);
nor U272 (N_272,In_21,In_515);
xor U273 (N_273,In_189,In_536);
nor U274 (N_274,In_895,In_334);
nand U275 (N_275,In_642,In_743);
and U276 (N_276,In_400,In_57);
xor U277 (N_277,In_419,In_750);
or U278 (N_278,In_262,In_426);
nor U279 (N_279,In_976,In_332);
nor U280 (N_280,In_212,In_58);
xor U281 (N_281,In_716,In_461);
nor U282 (N_282,In_98,In_0);
nor U283 (N_283,In_594,In_908);
nand U284 (N_284,In_770,In_157);
nor U285 (N_285,In_451,In_751);
or U286 (N_286,In_688,In_827);
and U287 (N_287,In_983,In_553);
and U288 (N_288,In_550,In_824);
xnor U289 (N_289,In_2,In_465);
nor U290 (N_290,In_771,In_696);
nor U291 (N_291,In_723,In_231);
xnor U292 (N_292,In_183,In_378);
and U293 (N_293,In_986,In_8);
or U294 (N_294,In_533,In_163);
or U295 (N_295,In_28,In_708);
nand U296 (N_296,In_689,In_502);
nand U297 (N_297,In_731,In_258);
nand U298 (N_298,In_925,In_863);
nor U299 (N_299,In_236,In_337);
and U300 (N_300,In_889,In_62);
nor U301 (N_301,In_722,In_518);
xor U302 (N_302,In_800,In_201);
nor U303 (N_303,In_505,In_866);
xor U304 (N_304,In_422,In_804);
nand U305 (N_305,In_488,In_818);
xnor U306 (N_306,In_380,In_123);
or U307 (N_307,In_733,In_138);
or U308 (N_308,In_437,In_186);
nand U309 (N_309,In_421,In_112);
nor U310 (N_310,In_506,In_898);
nand U311 (N_311,In_309,In_83);
nor U312 (N_312,In_372,In_417);
xnor U313 (N_313,In_145,In_961);
xor U314 (N_314,In_485,In_103);
nand U315 (N_315,In_479,In_452);
or U316 (N_316,In_631,In_912);
and U317 (N_317,In_710,In_321);
xnor U318 (N_318,In_715,In_903);
nand U319 (N_319,In_412,In_59);
xor U320 (N_320,In_175,In_459);
nor U321 (N_321,In_727,In_734);
nor U322 (N_322,In_666,In_694);
nor U323 (N_323,In_436,In_728);
and U324 (N_324,In_242,In_170);
or U325 (N_325,In_56,In_978);
or U326 (N_326,In_732,In_849);
nor U327 (N_327,In_383,In_920);
nand U328 (N_328,In_389,In_357);
nor U329 (N_329,In_968,In_85);
nor U330 (N_330,In_51,In_802);
xnor U331 (N_331,In_535,In_995);
or U332 (N_332,In_445,In_742);
xnor U333 (N_333,In_339,In_318);
and U334 (N_334,In_100,In_128);
or U335 (N_335,In_314,In_287);
xor U336 (N_336,In_184,In_755);
and U337 (N_337,In_4,In_355);
xnor U338 (N_338,In_179,In_31);
xnor U339 (N_339,In_652,In_541);
or U340 (N_340,In_272,In_187);
nor U341 (N_341,In_503,In_577);
and U342 (N_342,In_763,In_595);
and U343 (N_343,In_364,In_156);
and U344 (N_344,In_589,In_566);
and U345 (N_345,In_528,In_608);
xor U346 (N_346,In_126,In_954);
xnor U347 (N_347,In_835,In_697);
nand U348 (N_348,In_842,In_326);
and U349 (N_349,In_773,In_19);
nor U350 (N_350,In_246,In_538);
xnor U351 (N_351,In_312,In_705);
and U352 (N_352,In_721,In_330);
nand U353 (N_353,In_910,In_777);
nand U354 (N_354,In_294,In_604);
and U355 (N_355,In_288,In_331);
and U356 (N_356,In_27,In_643);
nor U357 (N_357,In_358,In_785);
and U358 (N_358,In_349,In_12);
or U359 (N_359,In_493,In_841);
nand U360 (N_360,In_23,In_95);
and U361 (N_361,In_971,In_439);
or U362 (N_362,In_943,In_96);
or U363 (N_363,In_951,In_20);
xor U364 (N_364,In_579,In_928);
nand U365 (N_365,In_343,In_268);
or U366 (N_366,In_308,In_6);
and U367 (N_367,In_887,In_117);
or U368 (N_368,In_512,In_373);
or U369 (N_369,In_304,In_583);
xnor U370 (N_370,In_546,In_852);
xor U371 (N_371,In_972,In_685);
xor U372 (N_372,In_155,In_394);
nor U373 (N_373,In_522,In_259);
and U374 (N_374,In_386,In_926);
nand U375 (N_375,In_87,In_940);
and U376 (N_376,In_279,In_927);
or U377 (N_377,In_934,In_313);
xor U378 (N_378,In_587,In_672);
nand U379 (N_379,In_654,In_18);
and U380 (N_380,In_195,In_952);
nor U381 (N_381,In_840,In_783);
nand U382 (N_382,In_219,In_317);
and U383 (N_383,In_89,In_741);
xor U384 (N_384,In_865,In_205);
and U385 (N_385,In_676,In_646);
and U386 (N_386,In_838,In_185);
xnor U387 (N_387,In_140,In_489);
nor U388 (N_388,In_173,In_881);
nor U389 (N_389,In_958,In_999);
nor U390 (N_390,In_110,In_260);
or U391 (N_391,In_101,In_736);
and U392 (N_392,In_481,In_562);
nor U393 (N_393,In_947,In_136);
or U394 (N_394,In_251,In_856);
nand U395 (N_395,In_609,In_850);
or U396 (N_396,In_360,In_299);
nand U397 (N_397,In_641,In_915);
xor U398 (N_398,In_669,In_438);
xor U399 (N_399,In_397,In_757);
or U400 (N_400,In_79,In_388);
xor U401 (N_401,In_379,In_527);
nor U402 (N_402,In_306,In_269);
or U403 (N_403,In_551,In_484);
or U404 (N_404,In_264,In_933);
or U405 (N_405,In_384,In_932);
and U406 (N_406,In_793,In_717);
nand U407 (N_407,In_375,In_166);
xnor U408 (N_408,In_102,In_674);
nand U409 (N_409,In_675,In_648);
or U410 (N_410,In_182,In_93);
nor U411 (N_411,In_431,In_853);
and U412 (N_412,In_208,In_942);
nand U413 (N_413,In_905,In_548);
and U414 (N_414,In_345,In_172);
xnor U415 (N_415,In_847,In_327);
and U416 (N_416,In_634,In_809);
or U417 (N_417,In_247,In_557);
nand U418 (N_418,In_293,In_180);
and U419 (N_419,In_893,In_839);
nand U420 (N_420,In_870,In_936);
xnor U421 (N_421,In_278,In_650);
nand U422 (N_422,In_177,In_862);
and U423 (N_423,In_72,In_831);
nand U424 (N_424,In_537,In_762);
or U425 (N_425,In_322,In_598);
nor U426 (N_426,In_55,In_909);
nor U427 (N_427,In_787,In_519);
xnor U428 (N_428,In_984,In_679);
and U429 (N_429,In_413,In_263);
or U430 (N_430,In_547,In_472);
and U431 (N_431,In_969,In_883);
or U432 (N_432,In_316,In_210);
and U433 (N_433,In_817,In_92);
nand U434 (N_434,In_104,In_405);
and U435 (N_435,In_610,In_252);
and U436 (N_436,In_937,In_975);
or U437 (N_437,In_989,In_486);
xnor U438 (N_438,In_806,In_221);
xnor U439 (N_439,In_410,In_329);
nand U440 (N_440,In_543,In_988);
or U441 (N_441,In_457,In_453);
or U442 (N_442,In_765,In_152);
or U443 (N_443,In_747,In_651);
and U444 (N_444,In_406,In_899);
xnor U445 (N_445,In_469,In_524);
and U446 (N_446,In_359,In_965);
or U447 (N_447,In_822,In_607);
xor U448 (N_448,In_366,In_473);
nand U449 (N_449,In_525,In_892);
xnor U450 (N_450,In_713,In_633);
nand U451 (N_451,In_408,In_7);
nand U452 (N_452,In_401,In_891);
nand U453 (N_453,In_684,In_285);
nand U454 (N_454,In_414,In_929);
or U455 (N_455,In_147,In_816);
xnor U456 (N_456,In_207,In_214);
nor U457 (N_457,In_333,In_629);
nor U458 (N_458,In_725,In_970);
or U459 (N_459,In_724,In_15);
nor U460 (N_460,In_613,In_630);
or U461 (N_461,In_508,In_137);
or U462 (N_462,In_249,In_90);
or U463 (N_463,In_521,In_1);
or U464 (N_464,In_65,In_561);
and U465 (N_465,In_659,In_567);
nor U466 (N_466,In_619,In_119);
or U467 (N_467,In_922,In_281);
nand U468 (N_468,In_80,In_222);
nor U469 (N_469,In_407,In_957);
xor U470 (N_470,In_632,In_580);
xor U471 (N_471,In_496,In_277);
or U472 (N_472,In_766,In_292);
nor U473 (N_473,In_939,In_813);
nand U474 (N_474,In_513,In_868);
and U475 (N_475,In_458,In_964);
nand U476 (N_476,In_649,In_432);
and U477 (N_477,In_860,In_315);
xor U478 (N_478,In_753,In_775);
nor U479 (N_479,In_637,In_544);
xor U480 (N_480,In_729,In_40);
and U481 (N_481,In_884,In_837);
or U482 (N_482,In_60,In_811);
and U483 (N_483,In_261,In_687);
nand U484 (N_484,In_815,In_52);
nand U485 (N_485,In_114,In_11);
and U486 (N_486,In_539,In_559);
nand U487 (N_487,In_520,In_624);
xor U488 (N_488,In_993,In_220);
nor U489 (N_489,In_462,In_61);
or U490 (N_490,In_882,In_746);
nor U491 (N_491,In_516,In_36);
nand U492 (N_492,In_930,In_510);
and U493 (N_493,In_441,In_444);
nand U494 (N_494,In_124,In_647);
nand U495 (N_495,In_677,In_240);
or U496 (N_496,In_756,In_116);
or U497 (N_497,In_812,In_280);
or U498 (N_498,In_693,In_719);
and U499 (N_499,In_574,In_829);
nand U500 (N_500,In_124,In_894);
and U501 (N_501,In_891,In_582);
nand U502 (N_502,In_471,In_831);
and U503 (N_503,In_267,In_13);
or U504 (N_504,In_43,In_647);
or U505 (N_505,In_912,In_517);
and U506 (N_506,In_741,In_821);
or U507 (N_507,In_922,In_761);
and U508 (N_508,In_272,In_364);
nand U509 (N_509,In_265,In_509);
xor U510 (N_510,In_146,In_5);
or U511 (N_511,In_483,In_351);
nor U512 (N_512,In_341,In_405);
nor U513 (N_513,In_643,In_632);
and U514 (N_514,In_896,In_559);
nand U515 (N_515,In_271,In_460);
xnor U516 (N_516,In_38,In_15);
and U517 (N_517,In_534,In_756);
nor U518 (N_518,In_519,In_852);
nand U519 (N_519,In_264,In_969);
nor U520 (N_520,In_654,In_235);
xnor U521 (N_521,In_290,In_694);
and U522 (N_522,In_779,In_712);
or U523 (N_523,In_329,In_188);
nor U524 (N_524,In_875,In_416);
nand U525 (N_525,In_364,In_43);
nor U526 (N_526,In_272,In_323);
xnor U527 (N_527,In_2,In_434);
nand U528 (N_528,In_147,In_564);
nand U529 (N_529,In_141,In_727);
nor U530 (N_530,In_357,In_806);
nor U531 (N_531,In_900,In_152);
nand U532 (N_532,In_202,In_409);
or U533 (N_533,In_419,In_148);
xor U534 (N_534,In_233,In_863);
xor U535 (N_535,In_80,In_136);
and U536 (N_536,In_60,In_471);
and U537 (N_537,In_893,In_422);
or U538 (N_538,In_474,In_393);
nand U539 (N_539,In_632,In_965);
xnor U540 (N_540,In_279,In_199);
xnor U541 (N_541,In_95,In_187);
and U542 (N_542,In_808,In_515);
nand U543 (N_543,In_99,In_733);
or U544 (N_544,In_57,In_240);
and U545 (N_545,In_543,In_903);
xor U546 (N_546,In_132,In_512);
or U547 (N_547,In_937,In_816);
xnor U548 (N_548,In_680,In_144);
xnor U549 (N_549,In_36,In_222);
nor U550 (N_550,In_113,In_724);
xnor U551 (N_551,In_727,In_182);
or U552 (N_552,In_51,In_453);
nor U553 (N_553,In_554,In_971);
nor U554 (N_554,In_150,In_440);
nand U555 (N_555,In_687,In_737);
xnor U556 (N_556,In_266,In_611);
xor U557 (N_557,In_561,In_570);
and U558 (N_558,In_873,In_446);
nor U559 (N_559,In_462,In_443);
xnor U560 (N_560,In_538,In_995);
and U561 (N_561,In_747,In_739);
nor U562 (N_562,In_634,In_469);
or U563 (N_563,In_935,In_826);
xnor U564 (N_564,In_105,In_403);
or U565 (N_565,In_615,In_153);
nor U566 (N_566,In_445,In_164);
and U567 (N_567,In_478,In_686);
and U568 (N_568,In_477,In_826);
or U569 (N_569,In_873,In_681);
or U570 (N_570,In_112,In_262);
xnor U571 (N_571,In_172,In_837);
xor U572 (N_572,In_522,In_647);
or U573 (N_573,In_250,In_424);
and U574 (N_574,In_985,In_696);
and U575 (N_575,In_920,In_97);
or U576 (N_576,In_118,In_343);
or U577 (N_577,In_886,In_258);
nor U578 (N_578,In_895,In_973);
and U579 (N_579,In_820,In_438);
or U580 (N_580,In_443,In_174);
xor U581 (N_581,In_662,In_971);
xnor U582 (N_582,In_627,In_55);
xor U583 (N_583,In_530,In_603);
or U584 (N_584,In_546,In_678);
xor U585 (N_585,In_6,In_286);
nor U586 (N_586,In_653,In_932);
nand U587 (N_587,In_360,In_494);
or U588 (N_588,In_380,In_157);
xnor U589 (N_589,In_979,In_427);
xor U590 (N_590,In_702,In_413);
xor U591 (N_591,In_664,In_592);
xor U592 (N_592,In_816,In_817);
and U593 (N_593,In_178,In_697);
xnor U594 (N_594,In_840,In_981);
nand U595 (N_595,In_418,In_711);
nor U596 (N_596,In_317,In_772);
xnor U597 (N_597,In_53,In_239);
nor U598 (N_598,In_229,In_985);
xnor U599 (N_599,In_145,In_460);
or U600 (N_600,In_217,In_517);
nor U601 (N_601,In_227,In_454);
nor U602 (N_602,In_982,In_666);
or U603 (N_603,In_748,In_6);
or U604 (N_604,In_403,In_702);
nor U605 (N_605,In_419,In_418);
xor U606 (N_606,In_841,In_875);
nor U607 (N_607,In_475,In_142);
and U608 (N_608,In_746,In_879);
xnor U609 (N_609,In_140,In_5);
xor U610 (N_610,In_98,In_332);
xor U611 (N_611,In_900,In_467);
or U612 (N_612,In_229,In_414);
and U613 (N_613,In_649,In_759);
nor U614 (N_614,In_450,In_324);
or U615 (N_615,In_828,In_764);
or U616 (N_616,In_72,In_5);
or U617 (N_617,In_260,In_318);
and U618 (N_618,In_61,In_558);
or U619 (N_619,In_546,In_921);
xor U620 (N_620,In_304,In_614);
xor U621 (N_621,In_10,In_60);
or U622 (N_622,In_702,In_787);
nor U623 (N_623,In_190,In_738);
nand U624 (N_624,In_260,In_816);
xnor U625 (N_625,In_752,In_724);
or U626 (N_626,In_382,In_711);
and U627 (N_627,In_669,In_648);
or U628 (N_628,In_953,In_732);
xnor U629 (N_629,In_718,In_128);
nor U630 (N_630,In_456,In_127);
nor U631 (N_631,In_251,In_214);
and U632 (N_632,In_217,In_583);
nand U633 (N_633,In_177,In_578);
xor U634 (N_634,In_703,In_222);
nor U635 (N_635,In_176,In_806);
and U636 (N_636,In_676,In_725);
nor U637 (N_637,In_328,In_758);
nand U638 (N_638,In_391,In_865);
and U639 (N_639,In_224,In_486);
xnor U640 (N_640,In_261,In_10);
or U641 (N_641,In_156,In_434);
and U642 (N_642,In_219,In_491);
xnor U643 (N_643,In_678,In_852);
or U644 (N_644,In_738,In_226);
nor U645 (N_645,In_539,In_63);
xor U646 (N_646,In_995,In_545);
xor U647 (N_647,In_135,In_554);
or U648 (N_648,In_50,In_564);
or U649 (N_649,In_781,In_193);
nor U650 (N_650,In_691,In_492);
nor U651 (N_651,In_971,In_881);
nor U652 (N_652,In_641,In_774);
xor U653 (N_653,In_303,In_768);
or U654 (N_654,In_389,In_517);
or U655 (N_655,In_938,In_281);
and U656 (N_656,In_264,In_682);
nor U657 (N_657,In_415,In_217);
nand U658 (N_658,In_620,In_768);
and U659 (N_659,In_606,In_821);
xnor U660 (N_660,In_376,In_511);
and U661 (N_661,In_285,In_820);
and U662 (N_662,In_93,In_883);
nand U663 (N_663,In_489,In_335);
and U664 (N_664,In_350,In_32);
nor U665 (N_665,In_323,In_79);
nand U666 (N_666,In_344,In_435);
xnor U667 (N_667,In_193,In_452);
nand U668 (N_668,In_900,In_438);
nor U669 (N_669,In_204,In_833);
and U670 (N_670,In_877,In_206);
xnor U671 (N_671,In_595,In_17);
and U672 (N_672,In_467,In_38);
nor U673 (N_673,In_532,In_402);
nor U674 (N_674,In_334,In_961);
nand U675 (N_675,In_699,In_705);
nor U676 (N_676,In_24,In_871);
xor U677 (N_677,In_81,In_31);
xor U678 (N_678,In_805,In_346);
xnor U679 (N_679,In_133,In_327);
and U680 (N_680,In_808,In_645);
or U681 (N_681,In_406,In_689);
nor U682 (N_682,In_621,In_830);
and U683 (N_683,In_993,In_507);
xor U684 (N_684,In_391,In_583);
and U685 (N_685,In_239,In_371);
nand U686 (N_686,In_874,In_324);
or U687 (N_687,In_611,In_296);
or U688 (N_688,In_927,In_76);
nor U689 (N_689,In_78,In_116);
and U690 (N_690,In_225,In_137);
nand U691 (N_691,In_59,In_943);
xor U692 (N_692,In_50,In_895);
nor U693 (N_693,In_261,In_564);
nor U694 (N_694,In_842,In_691);
nor U695 (N_695,In_756,In_458);
xnor U696 (N_696,In_629,In_321);
nor U697 (N_697,In_829,In_702);
or U698 (N_698,In_326,In_688);
or U699 (N_699,In_40,In_81);
or U700 (N_700,In_650,In_846);
nor U701 (N_701,In_346,In_965);
xor U702 (N_702,In_250,In_219);
nand U703 (N_703,In_215,In_796);
or U704 (N_704,In_972,In_385);
nand U705 (N_705,In_828,In_876);
and U706 (N_706,In_978,In_476);
nand U707 (N_707,In_314,In_639);
nand U708 (N_708,In_283,In_803);
nor U709 (N_709,In_927,In_644);
and U710 (N_710,In_682,In_150);
xor U711 (N_711,In_333,In_961);
nor U712 (N_712,In_94,In_986);
and U713 (N_713,In_71,In_250);
nor U714 (N_714,In_636,In_162);
nor U715 (N_715,In_182,In_675);
or U716 (N_716,In_808,In_250);
and U717 (N_717,In_222,In_170);
nor U718 (N_718,In_944,In_247);
nor U719 (N_719,In_661,In_672);
nor U720 (N_720,In_931,In_908);
nand U721 (N_721,In_536,In_635);
and U722 (N_722,In_782,In_206);
and U723 (N_723,In_816,In_176);
nand U724 (N_724,In_488,In_614);
or U725 (N_725,In_821,In_644);
nand U726 (N_726,In_689,In_463);
nor U727 (N_727,In_435,In_18);
or U728 (N_728,In_42,In_730);
nor U729 (N_729,In_908,In_530);
nand U730 (N_730,In_300,In_130);
or U731 (N_731,In_64,In_29);
nand U732 (N_732,In_885,In_405);
xnor U733 (N_733,In_520,In_766);
xor U734 (N_734,In_229,In_102);
or U735 (N_735,In_820,In_813);
xor U736 (N_736,In_158,In_630);
nand U737 (N_737,In_384,In_632);
or U738 (N_738,In_483,In_578);
or U739 (N_739,In_619,In_80);
or U740 (N_740,In_760,In_705);
nand U741 (N_741,In_12,In_303);
and U742 (N_742,In_974,In_885);
nor U743 (N_743,In_326,In_931);
nand U744 (N_744,In_883,In_433);
nor U745 (N_745,In_462,In_569);
xnor U746 (N_746,In_614,In_775);
nor U747 (N_747,In_821,In_623);
and U748 (N_748,In_675,In_211);
or U749 (N_749,In_670,In_464);
nor U750 (N_750,In_345,In_0);
and U751 (N_751,In_500,In_713);
xor U752 (N_752,In_847,In_488);
xnor U753 (N_753,In_322,In_463);
and U754 (N_754,In_21,In_24);
xor U755 (N_755,In_521,In_473);
nor U756 (N_756,In_970,In_269);
nand U757 (N_757,In_354,In_558);
and U758 (N_758,In_645,In_766);
nor U759 (N_759,In_205,In_606);
xnor U760 (N_760,In_338,In_601);
and U761 (N_761,In_660,In_683);
or U762 (N_762,In_920,In_679);
or U763 (N_763,In_3,In_829);
xnor U764 (N_764,In_689,In_865);
xnor U765 (N_765,In_725,In_69);
xor U766 (N_766,In_456,In_436);
nor U767 (N_767,In_123,In_873);
or U768 (N_768,In_473,In_325);
or U769 (N_769,In_950,In_532);
nand U770 (N_770,In_494,In_630);
nand U771 (N_771,In_375,In_661);
xnor U772 (N_772,In_836,In_503);
xor U773 (N_773,In_992,In_908);
or U774 (N_774,In_117,In_677);
and U775 (N_775,In_454,In_368);
and U776 (N_776,In_966,In_944);
and U777 (N_777,In_307,In_729);
or U778 (N_778,In_946,In_988);
and U779 (N_779,In_638,In_255);
and U780 (N_780,In_974,In_23);
and U781 (N_781,In_666,In_103);
nor U782 (N_782,In_707,In_804);
or U783 (N_783,In_291,In_719);
nand U784 (N_784,In_848,In_839);
or U785 (N_785,In_124,In_411);
or U786 (N_786,In_600,In_900);
nand U787 (N_787,In_418,In_605);
or U788 (N_788,In_958,In_87);
and U789 (N_789,In_42,In_451);
or U790 (N_790,In_266,In_623);
and U791 (N_791,In_650,In_909);
or U792 (N_792,In_855,In_414);
nand U793 (N_793,In_130,In_467);
and U794 (N_794,In_282,In_726);
nand U795 (N_795,In_493,In_149);
xnor U796 (N_796,In_278,In_384);
nand U797 (N_797,In_357,In_431);
xor U798 (N_798,In_267,In_143);
and U799 (N_799,In_458,In_939);
nor U800 (N_800,In_233,In_455);
nor U801 (N_801,In_210,In_36);
and U802 (N_802,In_781,In_792);
nand U803 (N_803,In_25,In_796);
nand U804 (N_804,In_399,In_636);
nand U805 (N_805,In_755,In_382);
xnor U806 (N_806,In_863,In_933);
nand U807 (N_807,In_958,In_940);
and U808 (N_808,In_615,In_862);
and U809 (N_809,In_660,In_175);
and U810 (N_810,In_38,In_854);
nand U811 (N_811,In_486,In_553);
nand U812 (N_812,In_185,In_820);
nor U813 (N_813,In_485,In_734);
nor U814 (N_814,In_653,In_171);
or U815 (N_815,In_846,In_567);
or U816 (N_816,In_428,In_967);
nor U817 (N_817,In_653,In_937);
or U818 (N_818,In_29,In_514);
nand U819 (N_819,In_873,In_486);
and U820 (N_820,In_472,In_136);
or U821 (N_821,In_481,In_321);
and U822 (N_822,In_985,In_659);
and U823 (N_823,In_61,In_891);
nor U824 (N_824,In_56,In_64);
or U825 (N_825,In_320,In_133);
xor U826 (N_826,In_880,In_186);
and U827 (N_827,In_960,In_559);
xor U828 (N_828,In_284,In_936);
or U829 (N_829,In_45,In_191);
or U830 (N_830,In_325,In_551);
xnor U831 (N_831,In_773,In_784);
and U832 (N_832,In_149,In_697);
nor U833 (N_833,In_109,In_423);
nor U834 (N_834,In_505,In_464);
nand U835 (N_835,In_851,In_283);
or U836 (N_836,In_326,In_641);
and U837 (N_837,In_805,In_947);
nor U838 (N_838,In_435,In_700);
xnor U839 (N_839,In_834,In_67);
nand U840 (N_840,In_332,In_308);
or U841 (N_841,In_382,In_786);
and U842 (N_842,In_251,In_297);
and U843 (N_843,In_725,In_968);
xor U844 (N_844,In_412,In_370);
nor U845 (N_845,In_246,In_744);
and U846 (N_846,In_960,In_541);
xnor U847 (N_847,In_127,In_332);
xor U848 (N_848,In_481,In_470);
xor U849 (N_849,In_452,In_928);
or U850 (N_850,In_611,In_888);
nor U851 (N_851,In_311,In_717);
and U852 (N_852,In_241,In_203);
and U853 (N_853,In_535,In_3);
or U854 (N_854,In_405,In_476);
or U855 (N_855,In_391,In_255);
or U856 (N_856,In_642,In_253);
or U857 (N_857,In_963,In_328);
nor U858 (N_858,In_61,In_280);
nor U859 (N_859,In_460,In_978);
nor U860 (N_860,In_312,In_227);
and U861 (N_861,In_682,In_449);
and U862 (N_862,In_15,In_764);
xor U863 (N_863,In_268,In_866);
nand U864 (N_864,In_308,In_687);
xor U865 (N_865,In_947,In_397);
nor U866 (N_866,In_101,In_497);
or U867 (N_867,In_174,In_753);
nor U868 (N_868,In_447,In_799);
xor U869 (N_869,In_674,In_784);
nand U870 (N_870,In_697,In_968);
and U871 (N_871,In_782,In_523);
or U872 (N_872,In_836,In_706);
or U873 (N_873,In_43,In_687);
nor U874 (N_874,In_421,In_545);
or U875 (N_875,In_761,In_297);
or U876 (N_876,In_37,In_642);
or U877 (N_877,In_154,In_186);
nand U878 (N_878,In_726,In_830);
and U879 (N_879,In_960,In_95);
nor U880 (N_880,In_955,In_603);
nand U881 (N_881,In_744,In_128);
and U882 (N_882,In_455,In_366);
xor U883 (N_883,In_589,In_493);
xor U884 (N_884,In_464,In_764);
or U885 (N_885,In_770,In_8);
or U886 (N_886,In_187,In_496);
xnor U887 (N_887,In_836,In_439);
xnor U888 (N_888,In_770,In_853);
xnor U889 (N_889,In_12,In_69);
nor U890 (N_890,In_735,In_383);
and U891 (N_891,In_670,In_747);
nor U892 (N_892,In_947,In_305);
and U893 (N_893,In_176,In_213);
and U894 (N_894,In_219,In_851);
and U895 (N_895,In_502,In_808);
or U896 (N_896,In_370,In_944);
nand U897 (N_897,In_631,In_768);
and U898 (N_898,In_989,In_280);
nor U899 (N_899,In_154,In_840);
nor U900 (N_900,In_779,In_330);
and U901 (N_901,In_917,In_790);
nand U902 (N_902,In_125,In_580);
xnor U903 (N_903,In_845,In_440);
nor U904 (N_904,In_239,In_720);
nor U905 (N_905,In_550,In_679);
or U906 (N_906,In_82,In_344);
nor U907 (N_907,In_784,In_391);
nor U908 (N_908,In_972,In_978);
xor U909 (N_909,In_402,In_649);
nand U910 (N_910,In_257,In_228);
nand U911 (N_911,In_668,In_764);
nand U912 (N_912,In_679,In_662);
nand U913 (N_913,In_860,In_560);
nor U914 (N_914,In_287,In_689);
and U915 (N_915,In_223,In_842);
nand U916 (N_916,In_840,In_825);
nor U917 (N_917,In_949,In_147);
xnor U918 (N_918,In_376,In_360);
nand U919 (N_919,In_254,In_505);
nand U920 (N_920,In_414,In_513);
nand U921 (N_921,In_715,In_768);
and U922 (N_922,In_175,In_479);
nor U923 (N_923,In_59,In_315);
nor U924 (N_924,In_375,In_480);
and U925 (N_925,In_35,In_776);
nor U926 (N_926,In_402,In_505);
xnor U927 (N_927,In_836,In_829);
nand U928 (N_928,In_772,In_927);
xor U929 (N_929,In_602,In_976);
nor U930 (N_930,In_133,In_973);
and U931 (N_931,In_333,In_574);
or U932 (N_932,In_805,In_80);
nor U933 (N_933,In_698,In_988);
and U934 (N_934,In_414,In_924);
xor U935 (N_935,In_777,In_684);
and U936 (N_936,In_123,In_323);
and U937 (N_937,In_570,In_728);
nor U938 (N_938,In_542,In_897);
xor U939 (N_939,In_261,In_881);
and U940 (N_940,In_900,In_502);
xor U941 (N_941,In_370,In_778);
nand U942 (N_942,In_575,In_944);
or U943 (N_943,In_601,In_207);
nand U944 (N_944,In_10,In_898);
xor U945 (N_945,In_568,In_127);
xnor U946 (N_946,In_585,In_558);
nand U947 (N_947,In_934,In_153);
and U948 (N_948,In_562,In_583);
nor U949 (N_949,In_60,In_669);
nand U950 (N_950,In_647,In_159);
nand U951 (N_951,In_104,In_409);
nor U952 (N_952,In_731,In_222);
nand U953 (N_953,In_655,In_451);
nor U954 (N_954,In_116,In_44);
xnor U955 (N_955,In_963,In_700);
or U956 (N_956,In_703,In_768);
or U957 (N_957,In_683,In_533);
and U958 (N_958,In_181,In_765);
nand U959 (N_959,In_217,In_128);
and U960 (N_960,In_872,In_272);
nor U961 (N_961,In_916,In_877);
or U962 (N_962,In_385,In_503);
xnor U963 (N_963,In_453,In_243);
nand U964 (N_964,In_513,In_166);
xnor U965 (N_965,In_648,In_752);
nand U966 (N_966,In_61,In_948);
nor U967 (N_967,In_109,In_786);
and U968 (N_968,In_905,In_282);
nor U969 (N_969,In_911,In_442);
xor U970 (N_970,In_935,In_193);
and U971 (N_971,In_743,In_10);
nor U972 (N_972,In_198,In_534);
or U973 (N_973,In_136,In_226);
nand U974 (N_974,In_597,In_871);
or U975 (N_975,In_139,In_475);
and U976 (N_976,In_186,In_76);
or U977 (N_977,In_193,In_37);
and U978 (N_978,In_963,In_894);
nor U979 (N_979,In_868,In_282);
or U980 (N_980,In_865,In_495);
and U981 (N_981,In_739,In_278);
or U982 (N_982,In_341,In_632);
nand U983 (N_983,In_974,In_718);
xor U984 (N_984,In_972,In_242);
or U985 (N_985,In_345,In_641);
nand U986 (N_986,In_559,In_920);
and U987 (N_987,In_774,In_441);
nor U988 (N_988,In_834,In_510);
or U989 (N_989,In_491,In_538);
nor U990 (N_990,In_391,In_786);
nor U991 (N_991,In_311,In_637);
and U992 (N_992,In_606,In_622);
or U993 (N_993,In_448,In_617);
nor U994 (N_994,In_573,In_25);
xor U995 (N_995,In_583,In_477);
and U996 (N_996,In_245,In_391);
nand U997 (N_997,In_627,In_108);
or U998 (N_998,In_496,In_426);
nor U999 (N_999,In_726,In_487);
nand U1000 (N_1000,In_399,In_915);
nand U1001 (N_1001,In_670,In_868);
nand U1002 (N_1002,In_641,In_393);
or U1003 (N_1003,In_415,In_259);
xor U1004 (N_1004,In_495,In_408);
or U1005 (N_1005,In_745,In_468);
and U1006 (N_1006,In_792,In_899);
xor U1007 (N_1007,In_832,In_393);
or U1008 (N_1008,In_666,In_417);
or U1009 (N_1009,In_980,In_160);
and U1010 (N_1010,In_409,In_577);
or U1011 (N_1011,In_731,In_337);
xnor U1012 (N_1012,In_633,In_671);
nand U1013 (N_1013,In_602,In_451);
nand U1014 (N_1014,In_891,In_463);
nor U1015 (N_1015,In_970,In_91);
nor U1016 (N_1016,In_466,In_418);
nor U1017 (N_1017,In_313,In_289);
or U1018 (N_1018,In_428,In_235);
nor U1019 (N_1019,In_933,In_428);
nor U1020 (N_1020,In_211,In_191);
nor U1021 (N_1021,In_19,In_417);
xor U1022 (N_1022,In_474,In_713);
nor U1023 (N_1023,In_330,In_75);
or U1024 (N_1024,In_287,In_445);
and U1025 (N_1025,In_597,In_826);
or U1026 (N_1026,In_898,In_164);
and U1027 (N_1027,In_185,In_445);
xnor U1028 (N_1028,In_198,In_836);
xor U1029 (N_1029,In_28,In_515);
and U1030 (N_1030,In_705,In_723);
nor U1031 (N_1031,In_291,In_717);
nor U1032 (N_1032,In_558,In_105);
and U1033 (N_1033,In_193,In_467);
or U1034 (N_1034,In_862,In_842);
nand U1035 (N_1035,In_52,In_22);
and U1036 (N_1036,In_547,In_897);
or U1037 (N_1037,In_742,In_309);
or U1038 (N_1038,In_685,In_425);
xnor U1039 (N_1039,In_817,In_762);
nor U1040 (N_1040,In_461,In_872);
xnor U1041 (N_1041,In_686,In_991);
or U1042 (N_1042,In_777,In_671);
xnor U1043 (N_1043,In_57,In_229);
and U1044 (N_1044,In_469,In_560);
or U1045 (N_1045,In_397,In_881);
and U1046 (N_1046,In_380,In_524);
and U1047 (N_1047,In_268,In_810);
or U1048 (N_1048,In_17,In_680);
nor U1049 (N_1049,In_626,In_428);
and U1050 (N_1050,In_273,In_269);
nor U1051 (N_1051,In_854,In_586);
nand U1052 (N_1052,In_715,In_331);
nand U1053 (N_1053,In_1,In_738);
xor U1054 (N_1054,In_704,In_100);
nand U1055 (N_1055,In_436,In_383);
or U1056 (N_1056,In_903,In_725);
xor U1057 (N_1057,In_760,In_184);
nand U1058 (N_1058,In_332,In_820);
nor U1059 (N_1059,In_539,In_246);
and U1060 (N_1060,In_928,In_653);
nor U1061 (N_1061,In_421,In_146);
nand U1062 (N_1062,In_576,In_486);
nor U1063 (N_1063,In_572,In_127);
or U1064 (N_1064,In_976,In_301);
nor U1065 (N_1065,In_715,In_187);
xnor U1066 (N_1066,In_47,In_90);
nor U1067 (N_1067,In_602,In_907);
xor U1068 (N_1068,In_778,In_118);
or U1069 (N_1069,In_38,In_486);
nor U1070 (N_1070,In_462,In_785);
nor U1071 (N_1071,In_806,In_463);
nand U1072 (N_1072,In_568,In_343);
and U1073 (N_1073,In_136,In_456);
or U1074 (N_1074,In_38,In_223);
and U1075 (N_1075,In_160,In_921);
nor U1076 (N_1076,In_123,In_667);
xnor U1077 (N_1077,In_755,In_941);
xnor U1078 (N_1078,In_50,In_373);
nor U1079 (N_1079,In_972,In_898);
xor U1080 (N_1080,In_791,In_555);
or U1081 (N_1081,In_887,In_835);
or U1082 (N_1082,In_88,In_403);
nor U1083 (N_1083,In_460,In_561);
and U1084 (N_1084,In_113,In_355);
nand U1085 (N_1085,In_194,In_241);
nand U1086 (N_1086,In_306,In_109);
xor U1087 (N_1087,In_216,In_254);
xnor U1088 (N_1088,In_198,In_241);
and U1089 (N_1089,In_544,In_193);
nand U1090 (N_1090,In_706,In_989);
or U1091 (N_1091,In_24,In_121);
xor U1092 (N_1092,In_813,In_462);
and U1093 (N_1093,In_255,In_225);
nand U1094 (N_1094,In_469,In_51);
and U1095 (N_1095,In_786,In_511);
or U1096 (N_1096,In_430,In_983);
nand U1097 (N_1097,In_709,In_949);
nor U1098 (N_1098,In_18,In_606);
xor U1099 (N_1099,In_900,In_886);
and U1100 (N_1100,In_520,In_361);
or U1101 (N_1101,In_86,In_949);
nor U1102 (N_1102,In_218,In_139);
xnor U1103 (N_1103,In_322,In_756);
nor U1104 (N_1104,In_470,In_665);
nand U1105 (N_1105,In_109,In_719);
nor U1106 (N_1106,In_289,In_940);
or U1107 (N_1107,In_804,In_853);
nand U1108 (N_1108,In_414,In_810);
nor U1109 (N_1109,In_480,In_430);
or U1110 (N_1110,In_574,In_19);
nand U1111 (N_1111,In_581,In_724);
or U1112 (N_1112,In_73,In_947);
or U1113 (N_1113,In_315,In_817);
nor U1114 (N_1114,In_254,In_107);
nor U1115 (N_1115,In_740,In_98);
or U1116 (N_1116,In_501,In_522);
or U1117 (N_1117,In_42,In_376);
nand U1118 (N_1118,In_491,In_113);
nand U1119 (N_1119,In_433,In_581);
nor U1120 (N_1120,In_434,In_750);
nor U1121 (N_1121,In_288,In_703);
and U1122 (N_1122,In_918,In_711);
nor U1123 (N_1123,In_782,In_656);
and U1124 (N_1124,In_387,In_506);
and U1125 (N_1125,In_184,In_99);
xnor U1126 (N_1126,In_820,In_762);
nand U1127 (N_1127,In_686,In_720);
xor U1128 (N_1128,In_485,In_239);
and U1129 (N_1129,In_371,In_222);
xor U1130 (N_1130,In_621,In_52);
nor U1131 (N_1131,In_674,In_613);
xnor U1132 (N_1132,In_594,In_441);
or U1133 (N_1133,In_89,In_983);
and U1134 (N_1134,In_826,In_996);
nor U1135 (N_1135,In_523,In_238);
nor U1136 (N_1136,In_467,In_401);
xor U1137 (N_1137,In_597,In_406);
nand U1138 (N_1138,In_690,In_909);
or U1139 (N_1139,In_212,In_177);
nand U1140 (N_1140,In_202,In_448);
nand U1141 (N_1141,In_587,In_348);
nand U1142 (N_1142,In_839,In_319);
or U1143 (N_1143,In_437,In_193);
nor U1144 (N_1144,In_461,In_361);
or U1145 (N_1145,In_73,In_963);
xnor U1146 (N_1146,In_600,In_619);
and U1147 (N_1147,In_16,In_540);
or U1148 (N_1148,In_765,In_539);
nand U1149 (N_1149,In_487,In_339);
and U1150 (N_1150,In_16,In_910);
xnor U1151 (N_1151,In_821,In_483);
or U1152 (N_1152,In_920,In_987);
nand U1153 (N_1153,In_328,In_44);
nor U1154 (N_1154,In_826,In_716);
or U1155 (N_1155,In_717,In_899);
xor U1156 (N_1156,In_290,In_175);
and U1157 (N_1157,In_867,In_690);
nor U1158 (N_1158,In_251,In_720);
nand U1159 (N_1159,In_982,In_195);
nor U1160 (N_1160,In_813,In_835);
and U1161 (N_1161,In_576,In_406);
xor U1162 (N_1162,In_2,In_95);
nor U1163 (N_1163,In_373,In_545);
nand U1164 (N_1164,In_47,In_256);
or U1165 (N_1165,In_197,In_722);
or U1166 (N_1166,In_46,In_908);
xnor U1167 (N_1167,In_879,In_573);
xnor U1168 (N_1168,In_504,In_643);
or U1169 (N_1169,In_385,In_129);
or U1170 (N_1170,In_76,In_841);
xnor U1171 (N_1171,In_237,In_770);
xor U1172 (N_1172,In_354,In_129);
xor U1173 (N_1173,In_540,In_273);
nand U1174 (N_1174,In_116,In_52);
and U1175 (N_1175,In_582,In_809);
nor U1176 (N_1176,In_246,In_184);
or U1177 (N_1177,In_365,In_134);
or U1178 (N_1178,In_841,In_632);
nor U1179 (N_1179,In_290,In_654);
and U1180 (N_1180,In_771,In_822);
xnor U1181 (N_1181,In_540,In_594);
xor U1182 (N_1182,In_4,In_519);
or U1183 (N_1183,In_687,In_602);
nor U1184 (N_1184,In_444,In_678);
nor U1185 (N_1185,In_868,In_66);
or U1186 (N_1186,In_760,In_112);
nor U1187 (N_1187,In_560,In_573);
nor U1188 (N_1188,In_920,In_628);
nor U1189 (N_1189,In_247,In_4);
nand U1190 (N_1190,In_587,In_253);
nor U1191 (N_1191,In_134,In_743);
nor U1192 (N_1192,In_964,In_724);
xnor U1193 (N_1193,In_879,In_774);
nand U1194 (N_1194,In_128,In_192);
nor U1195 (N_1195,In_774,In_678);
xnor U1196 (N_1196,In_724,In_83);
or U1197 (N_1197,In_462,In_193);
nor U1198 (N_1198,In_782,In_920);
xor U1199 (N_1199,In_957,In_716);
and U1200 (N_1200,In_964,In_746);
or U1201 (N_1201,In_575,In_863);
nand U1202 (N_1202,In_733,In_791);
nor U1203 (N_1203,In_40,In_741);
nor U1204 (N_1204,In_472,In_969);
and U1205 (N_1205,In_71,In_855);
xor U1206 (N_1206,In_144,In_507);
nor U1207 (N_1207,In_306,In_782);
nand U1208 (N_1208,In_8,In_386);
or U1209 (N_1209,In_973,In_166);
xnor U1210 (N_1210,In_216,In_417);
and U1211 (N_1211,In_801,In_217);
nand U1212 (N_1212,In_404,In_943);
or U1213 (N_1213,In_581,In_855);
nor U1214 (N_1214,In_817,In_574);
or U1215 (N_1215,In_105,In_98);
nand U1216 (N_1216,In_380,In_187);
nand U1217 (N_1217,In_279,In_460);
nor U1218 (N_1218,In_913,In_839);
or U1219 (N_1219,In_792,In_892);
and U1220 (N_1220,In_824,In_168);
nand U1221 (N_1221,In_590,In_912);
and U1222 (N_1222,In_825,In_19);
nor U1223 (N_1223,In_454,In_524);
or U1224 (N_1224,In_300,In_855);
and U1225 (N_1225,In_707,In_101);
or U1226 (N_1226,In_6,In_679);
or U1227 (N_1227,In_598,In_435);
xnor U1228 (N_1228,In_945,In_760);
nand U1229 (N_1229,In_613,In_728);
xnor U1230 (N_1230,In_90,In_267);
nor U1231 (N_1231,In_876,In_441);
and U1232 (N_1232,In_765,In_526);
nand U1233 (N_1233,In_948,In_187);
nor U1234 (N_1234,In_431,In_324);
and U1235 (N_1235,In_219,In_901);
xor U1236 (N_1236,In_472,In_687);
nand U1237 (N_1237,In_542,In_288);
or U1238 (N_1238,In_439,In_464);
nor U1239 (N_1239,In_225,In_838);
or U1240 (N_1240,In_240,In_909);
and U1241 (N_1241,In_697,In_951);
and U1242 (N_1242,In_973,In_706);
and U1243 (N_1243,In_168,In_926);
nand U1244 (N_1244,In_560,In_206);
and U1245 (N_1245,In_3,In_14);
or U1246 (N_1246,In_886,In_245);
xor U1247 (N_1247,In_191,In_311);
or U1248 (N_1248,In_491,In_308);
and U1249 (N_1249,In_513,In_225);
xnor U1250 (N_1250,In_405,In_717);
xor U1251 (N_1251,In_531,In_819);
and U1252 (N_1252,In_892,In_877);
or U1253 (N_1253,In_254,In_894);
and U1254 (N_1254,In_121,In_120);
or U1255 (N_1255,In_750,In_4);
or U1256 (N_1256,In_5,In_812);
nor U1257 (N_1257,In_74,In_194);
or U1258 (N_1258,In_341,In_137);
nand U1259 (N_1259,In_192,In_731);
xnor U1260 (N_1260,In_594,In_259);
and U1261 (N_1261,In_645,In_355);
nand U1262 (N_1262,In_150,In_395);
nand U1263 (N_1263,In_993,In_946);
and U1264 (N_1264,In_240,In_921);
nor U1265 (N_1265,In_281,In_847);
and U1266 (N_1266,In_591,In_901);
or U1267 (N_1267,In_919,In_953);
nand U1268 (N_1268,In_891,In_299);
xnor U1269 (N_1269,In_176,In_138);
and U1270 (N_1270,In_645,In_493);
and U1271 (N_1271,In_480,In_147);
nor U1272 (N_1272,In_349,In_651);
or U1273 (N_1273,In_985,In_172);
nor U1274 (N_1274,In_520,In_92);
or U1275 (N_1275,In_276,In_284);
xor U1276 (N_1276,In_943,In_814);
or U1277 (N_1277,In_551,In_584);
or U1278 (N_1278,In_414,In_500);
xnor U1279 (N_1279,In_365,In_856);
and U1280 (N_1280,In_312,In_339);
or U1281 (N_1281,In_132,In_27);
xnor U1282 (N_1282,In_961,In_994);
and U1283 (N_1283,In_220,In_506);
and U1284 (N_1284,In_560,In_444);
and U1285 (N_1285,In_8,In_368);
or U1286 (N_1286,In_727,In_832);
and U1287 (N_1287,In_473,In_650);
nor U1288 (N_1288,In_991,In_933);
nor U1289 (N_1289,In_295,In_71);
nor U1290 (N_1290,In_541,In_258);
or U1291 (N_1291,In_639,In_56);
nand U1292 (N_1292,In_858,In_841);
xor U1293 (N_1293,In_677,In_600);
nor U1294 (N_1294,In_775,In_77);
and U1295 (N_1295,In_818,In_288);
and U1296 (N_1296,In_650,In_306);
nand U1297 (N_1297,In_514,In_362);
or U1298 (N_1298,In_338,In_116);
and U1299 (N_1299,In_940,In_52);
xor U1300 (N_1300,In_371,In_493);
and U1301 (N_1301,In_275,In_208);
nor U1302 (N_1302,In_663,In_307);
xor U1303 (N_1303,In_21,In_252);
and U1304 (N_1304,In_478,In_77);
nor U1305 (N_1305,In_93,In_59);
xor U1306 (N_1306,In_306,In_167);
nor U1307 (N_1307,In_472,In_949);
nor U1308 (N_1308,In_660,In_897);
or U1309 (N_1309,In_237,In_460);
xnor U1310 (N_1310,In_434,In_598);
xor U1311 (N_1311,In_708,In_78);
and U1312 (N_1312,In_976,In_267);
and U1313 (N_1313,In_97,In_314);
nand U1314 (N_1314,In_44,In_169);
and U1315 (N_1315,In_477,In_462);
nor U1316 (N_1316,In_730,In_48);
or U1317 (N_1317,In_661,In_274);
xor U1318 (N_1318,In_753,In_470);
or U1319 (N_1319,In_610,In_21);
xor U1320 (N_1320,In_153,In_970);
nor U1321 (N_1321,In_374,In_80);
and U1322 (N_1322,In_968,In_749);
and U1323 (N_1323,In_398,In_736);
nand U1324 (N_1324,In_577,In_324);
nand U1325 (N_1325,In_416,In_160);
or U1326 (N_1326,In_226,In_76);
nand U1327 (N_1327,In_757,In_295);
xnor U1328 (N_1328,In_88,In_416);
nand U1329 (N_1329,In_947,In_535);
and U1330 (N_1330,In_274,In_896);
and U1331 (N_1331,In_215,In_433);
xnor U1332 (N_1332,In_717,In_172);
xor U1333 (N_1333,In_229,In_895);
or U1334 (N_1334,In_227,In_576);
and U1335 (N_1335,In_959,In_43);
and U1336 (N_1336,In_533,In_291);
nor U1337 (N_1337,In_79,In_306);
xnor U1338 (N_1338,In_277,In_202);
and U1339 (N_1339,In_213,In_964);
or U1340 (N_1340,In_109,In_795);
nor U1341 (N_1341,In_299,In_753);
nor U1342 (N_1342,In_520,In_850);
nor U1343 (N_1343,In_756,In_984);
nand U1344 (N_1344,In_182,In_576);
nor U1345 (N_1345,In_442,In_332);
nand U1346 (N_1346,In_721,In_937);
nand U1347 (N_1347,In_317,In_30);
or U1348 (N_1348,In_719,In_584);
nand U1349 (N_1349,In_237,In_276);
nand U1350 (N_1350,In_263,In_325);
or U1351 (N_1351,In_499,In_919);
nor U1352 (N_1352,In_420,In_442);
nand U1353 (N_1353,In_618,In_103);
or U1354 (N_1354,In_185,In_329);
and U1355 (N_1355,In_508,In_449);
xor U1356 (N_1356,In_462,In_829);
nor U1357 (N_1357,In_163,In_554);
xnor U1358 (N_1358,In_228,In_615);
or U1359 (N_1359,In_253,In_485);
nor U1360 (N_1360,In_44,In_556);
xnor U1361 (N_1361,In_899,In_982);
and U1362 (N_1362,In_554,In_920);
xnor U1363 (N_1363,In_124,In_696);
nand U1364 (N_1364,In_67,In_736);
nand U1365 (N_1365,In_508,In_644);
nand U1366 (N_1366,In_954,In_54);
nand U1367 (N_1367,In_219,In_433);
nand U1368 (N_1368,In_450,In_503);
nand U1369 (N_1369,In_415,In_764);
or U1370 (N_1370,In_746,In_214);
nor U1371 (N_1371,In_137,In_990);
xor U1372 (N_1372,In_39,In_865);
nand U1373 (N_1373,In_189,In_586);
nor U1374 (N_1374,In_377,In_211);
nand U1375 (N_1375,In_412,In_213);
nor U1376 (N_1376,In_54,In_332);
and U1377 (N_1377,In_657,In_597);
or U1378 (N_1378,In_839,In_456);
or U1379 (N_1379,In_979,In_760);
xor U1380 (N_1380,In_440,In_594);
nand U1381 (N_1381,In_184,In_478);
nor U1382 (N_1382,In_620,In_635);
nor U1383 (N_1383,In_193,In_482);
nor U1384 (N_1384,In_826,In_773);
or U1385 (N_1385,In_238,In_510);
nand U1386 (N_1386,In_511,In_74);
xor U1387 (N_1387,In_381,In_868);
xnor U1388 (N_1388,In_804,In_81);
xor U1389 (N_1389,In_154,In_915);
or U1390 (N_1390,In_343,In_559);
and U1391 (N_1391,In_402,In_642);
and U1392 (N_1392,In_47,In_720);
nand U1393 (N_1393,In_592,In_318);
nor U1394 (N_1394,In_386,In_974);
xor U1395 (N_1395,In_112,In_934);
and U1396 (N_1396,In_126,In_65);
xor U1397 (N_1397,In_18,In_863);
and U1398 (N_1398,In_302,In_702);
xor U1399 (N_1399,In_549,In_552);
and U1400 (N_1400,In_82,In_349);
nor U1401 (N_1401,In_9,In_607);
or U1402 (N_1402,In_634,In_838);
nor U1403 (N_1403,In_126,In_318);
nand U1404 (N_1404,In_36,In_368);
xnor U1405 (N_1405,In_670,In_595);
or U1406 (N_1406,In_329,In_68);
xor U1407 (N_1407,In_713,In_963);
xnor U1408 (N_1408,In_878,In_678);
or U1409 (N_1409,In_696,In_624);
nand U1410 (N_1410,In_246,In_487);
and U1411 (N_1411,In_519,In_29);
nand U1412 (N_1412,In_38,In_136);
nor U1413 (N_1413,In_951,In_100);
and U1414 (N_1414,In_904,In_656);
and U1415 (N_1415,In_772,In_303);
xor U1416 (N_1416,In_123,In_641);
and U1417 (N_1417,In_300,In_238);
and U1418 (N_1418,In_399,In_80);
nand U1419 (N_1419,In_866,In_879);
or U1420 (N_1420,In_863,In_151);
and U1421 (N_1421,In_817,In_600);
nor U1422 (N_1422,In_220,In_677);
and U1423 (N_1423,In_462,In_988);
and U1424 (N_1424,In_728,In_973);
nor U1425 (N_1425,In_403,In_936);
nand U1426 (N_1426,In_425,In_853);
xor U1427 (N_1427,In_7,In_949);
nand U1428 (N_1428,In_970,In_219);
and U1429 (N_1429,In_482,In_650);
nor U1430 (N_1430,In_847,In_573);
and U1431 (N_1431,In_847,In_167);
or U1432 (N_1432,In_616,In_567);
nand U1433 (N_1433,In_934,In_443);
xor U1434 (N_1434,In_449,In_995);
xnor U1435 (N_1435,In_67,In_693);
nor U1436 (N_1436,In_282,In_12);
nor U1437 (N_1437,In_41,In_835);
xnor U1438 (N_1438,In_91,In_313);
nor U1439 (N_1439,In_933,In_654);
or U1440 (N_1440,In_754,In_516);
and U1441 (N_1441,In_662,In_555);
or U1442 (N_1442,In_6,In_998);
xor U1443 (N_1443,In_386,In_765);
nand U1444 (N_1444,In_984,In_17);
nand U1445 (N_1445,In_320,In_834);
nor U1446 (N_1446,In_634,In_803);
nor U1447 (N_1447,In_785,In_828);
nor U1448 (N_1448,In_746,In_189);
or U1449 (N_1449,In_518,In_322);
xnor U1450 (N_1450,In_417,In_126);
xnor U1451 (N_1451,In_218,In_948);
or U1452 (N_1452,In_260,In_156);
and U1453 (N_1453,In_354,In_800);
and U1454 (N_1454,In_380,In_894);
nor U1455 (N_1455,In_923,In_637);
nor U1456 (N_1456,In_543,In_468);
xnor U1457 (N_1457,In_399,In_605);
xnor U1458 (N_1458,In_789,In_559);
nor U1459 (N_1459,In_671,In_743);
or U1460 (N_1460,In_975,In_752);
or U1461 (N_1461,In_929,In_711);
nor U1462 (N_1462,In_835,In_160);
and U1463 (N_1463,In_355,In_922);
and U1464 (N_1464,In_7,In_574);
nand U1465 (N_1465,In_878,In_185);
nand U1466 (N_1466,In_344,In_156);
nand U1467 (N_1467,In_192,In_101);
or U1468 (N_1468,In_136,In_775);
or U1469 (N_1469,In_710,In_655);
xnor U1470 (N_1470,In_415,In_744);
nand U1471 (N_1471,In_294,In_162);
nor U1472 (N_1472,In_763,In_447);
nor U1473 (N_1473,In_657,In_170);
nand U1474 (N_1474,In_116,In_760);
nor U1475 (N_1475,In_97,In_380);
or U1476 (N_1476,In_179,In_213);
nand U1477 (N_1477,In_72,In_969);
xnor U1478 (N_1478,In_856,In_244);
or U1479 (N_1479,In_394,In_689);
xnor U1480 (N_1480,In_822,In_487);
nor U1481 (N_1481,In_252,In_424);
xnor U1482 (N_1482,In_333,In_543);
or U1483 (N_1483,In_936,In_345);
nor U1484 (N_1484,In_391,In_345);
or U1485 (N_1485,In_860,In_925);
and U1486 (N_1486,In_592,In_355);
xnor U1487 (N_1487,In_667,In_181);
nand U1488 (N_1488,In_567,In_876);
or U1489 (N_1489,In_987,In_547);
and U1490 (N_1490,In_29,In_375);
or U1491 (N_1491,In_516,In_912);
nand U1492 (N_1492,In_667,In_804);
nand U1493 (N_1493,In_869,In_767);
nor U1494 (N_1494,In_788,In_423);
nor U1495 (N_1495,In_989,In_55);
nand U1496 (N_1496,In_921,In_705);
or U1497 (N_1497,In_229,In_602);
xnor U1498 (N_1498,In_407,In_796);
xor U1499 (N_1499,In_254,In_939);
or U1500 (N_1500,In_408,In_506);
xnor U1501 (N_1501,In_999,In_641);
nor U1502 (N_1502,In_626,In_382);
xnor U1503 (N_1503,In_183,In_6);
or U1504 (N_1504,In_43,In_254);
and U1505 (N_1505,In_331,In_387);
or U1506 (N_1506,In_885,In_459);
and U1507 (N_1507,In_748,In_168);
nor U1508 (N_1508,In_11,In_373);
nor U1509 (N_1509,In_851,In_935);
nand U1510 (N_1510,In_864,In_789);
nand U1511 (N_1511,In_545,In_46);
and U1512 (N_1512,In_938,In_4);
nor U1513 (N_1513,In_313,In_940);
and U1514 (N_1514,In_745,In_9);
or U1515 (N_1515,In_104,In_815);
nand U1516 (N_1516,In_792,In_48);
or U1517 (N_1517,In_638,In_275);
or U1518 (N_1518,In_0,In_363);
and U1519 (N_1519,In_295,In_607);
nand U1520 (N_1520,In_362,In_202);
and U1521 (N_1521,In_335,In_294);
nor U1522 (N_1522,In_585,In_98);
nand U1523 (N_1523,In_60,In_104);
nor U1524 (N_1524,In_67,In_924);
or U1525 (N_1525,In_305,In_986);
or U1526 (N_1526,In_835,In_705);
xnor U1527 (N_1527,In_674,In_233);
nor U1528 (N_1528,In_264,In_19);
nand U1529 (N_1529,In_346,In_869);
or U1530 (N_1530,In_929,In_113);
or U1531 (N_1531,In_37,In_50);
or U1532 (N_1532,In_590,In_579);
and U1533 (N_1533,In_230,In_80);
nand U1534 (N_1534,In_39,In_390);
xnor U1535 (N_1535,In_299,In_874);
nand U1536 (N_1536,In_182,In_283);
and U1537 (N_1537,In_332,In_783);
xnor U1538 (N_1538,In_193,In_295);
or U1539 (N_1539,In_252,In_460);
nand U1540 (N_1540,In_499,In_808);
xnor U1541 (N_1541,In_463,In_956);
or U1542 (N_1542,In_637,In_438);
nand U1543 (N_1543,In_102,In_576);
nand U1544 (N_1544,In_420,In_598);
nand U1545 (N_1545,In_449,In_203);
xnor U1546 (N_1546,In_86,In_750);
nand U1547 (N_1547,In_237,In_792);
or U1548 (N_1548,In_642,In_894);
xnor U1549 (N_1549,In_175,In_455);
nand U1550 (N_1550,In_948,In_19);
nor U1551 (N_1551,In_556,In_808);
nand U1552 (N_1552,In_820,In_888);
or U1553 (N_1553,In_72,In_57);
or U1554 (N_1554,In_558,In_306);
nor U1555 (N_1555,In_233,In_28);
and U1556 (N_1556,In_403,In_705);
nor U1557 (N_1557,In_637,In_449);
nor U1558 (N_1558,In_188,In_634);
xnor U1559 (N_1559,In_328,In_787);
xnor U1560 (N_1560,In_13,In_438);
and U1561 (N_1561,In_713,In_344);
nor U1562 (N_1562,In_587,In_197);
or U1563 (N_1563,In_272,In_816);
and U1564 (N_1564,In_353,In_960);
or U1565 (N_1565,In_202,In_626);
and U1566 (N_1566,In_275,In_733);
nand U1567 (N_1567,In_201,In_702);
or U1568 (N_1568,In_234,In_531);
nor U1569 (N_1569,In_790,In_311);
nand U1570 (N_1570,In_810,In_68);
nand U1571 (N_1571,In_568,In_112);
nand U1572 (N_1572,In_207,In_110);
and U1573 (N_1573,In_768,In_896);
or U1574 (N_1574,In_171,In_873);
nor U1575 (N_1575,In_135,In_826);
and U1576 (N_1576,In_897,In_509);
or U1577 (N_1577,In_513,In_181);
nand U1578 (N_1578,In_804,In_603);
nand U1579 (N_1579,In_121,In_496);
nand U1580 (N_1580,In_344,In_34);
nand U1581 (N_1581,In_899,In_810);
and U1582 (N_1582,In_915,In_448);
or U1583 (N_1583,In_600,In_856);
xnor U1584 (N_1584,In_925,In_732);
and U1585 (N_1585,In_345,In_591);
xor U1586 (N_1586,In_942,In_974);
or U1587 (N_1587,In_613,In_125);
nand U1588 (N_1588,In_648,In_380);
and U1589 (N_1589,In_852,In_868);
nand U1590 (N_1590,In_589,In_708);
or U1591 (N_1591,In_46,In_244);
nor U1592 (N_1592,In_585,In_293);
and U1593 (N_1593,In_525,In_718);
xnor U1594 (N_1594,In_243,In_972);
nor U1595 (N_1595,In_291,In_932);
or U1596 (N_1596,In_782,In_197);
and U1597 (N_1597,In_613,In_352);
nor U1598 (N_1598,In_682,In_89);
and U1599 (N_1599,In_283,In_92);
nor U1600 (N_1600,In_987,In_258);
xnor U1601 (N_1601,In_174,In_34);
xor U1602 (N_1602,In_353,In_90);
xor U1603 (N_1603,In_933,In_117);
nor U1604 (N_1604,In_585,In_695);
xor U1605 (N_1605,In_715,In_604);
nor U1606 (N_1606,In_743,In_305);
or U1607 (N_1607,In_326,In_350);
and U1608 (N_1608,In_820,In_721);
or U1609 (N_1609,In_648,In_717);
or U1610 (N_1610,In_542,In_247);
nor U1611 (N_1611,In_889,In_717);
nand U1612 (N_1612,In_653,In_552);
and U1613 (N_1613,In_33,In_355);
and U1614 (N_1614,In_563,In_923);
and U1615 (N_1615,In_580,In_367);
and U1616 (N_1616,In_347,In_808);
nor U1617 (N_1617,In_692,In_416);
and U1618 (N_1618,In_320,In_504);
xor U1619 (N_1619,In_496,In_771);
xnor U1620 (N_1620,In_691,In_425);
and U1621 (N_1621,In_778,In_867);
or U1622 (N_1622,In_581,In_877);
or U1623 (N_1623,In_198,In_760);
nor U1624 (N_1624,In_762,In_452);
nand U1625 (N_1625,In_25,In_425);
xnor U1626 (N_1626,In_391,In_18);
or U1627 (N_1627,In_19,In_26);
and U1628 (N_1628,In_473,In_637);
nor U1629 (N_1629,In_685,In_272);
and U1630 (N_1630,In_79,In_330);
nor U1631 (N_1631,In_262,In_994);
and U1632 (N_1632,In_262,In_104);
xor U1633 (N_1633,In_371,In_658);
and U1634 (N_1634,In_705,In_583);
or U1635 (N_1635,In_435,In_95);
xor U1636 (N_1636,In_203,In_865);
or U1637 (N_1637,In_218,In_200);
or U1638 (N_1638,In_889,In_644);
nand U1639 (N_1639,In_311,In_283);
or U1640 (N_1640,In_43,In_686);
or U1641 (N_1641,In_137,In_821);
and U1642 (N_1642,In_13,In_883);
or U1643 (N_1643,In_204,In_101);
or U1644 (N_1644,In_185,In_78);
or U1645 (N_1645,In_893,In_662);
or U1646 (N_1646,In_366,In_650);
or U1647 (N_1647,In_918,In_314);
nor U1648 (N_1648,In_553,In_138);
nand U1649 (N_1649,In_51,In_884);
xor U1650 (N_1650,In_246,In_652);
or U1651 (N_1651,In_954,In_960);
xor U1652 (N_1652,In_297,In_600);
and U1653 (N_1653,In_828,In_136);
and U1654 (N_1654,In_348,In_987);
nor U1655 (N_1655,In_983,In_488);
or U1656 (N_1656,In_970,In_291);
nor U1657 (N_1657,In_528,In_13);
nor U1658 (N_1658,In_800,In_91);
nand U1659 (N_1659,In_148,In_709);
and U1660 (N_1660,In_667,In_565);
or U1661 (N_1661,In_338,In_458);
nor U1662 (N_1662,In_575,In_315);
xor U1663 (N_1663,In_807,In_783);
nand U1664 (N_1664,In_742,In_598);
or U1665 (N_1665,In_745,In_977);
xnor U1666 (N_1666,In_994,In_325);
or U1667 (N_1667,In_538,In_77);
nand U1668 (N_1668,In_486,In_893);
and U1669 (N_1669,In_215,In_837);
nor U1670 (N_1670,In_884,In_636);
or U1671 (N_1671,In_418,In_437);
nand U1672 (N_1672,In_476,In_330);
nand U1673 (N_1673,In_856,In_112);
and U1674 (N_1674,In_909,In_90);
nor U1675 (N_1675,In_936,In_915);
or U1676 (N_1676,In_3,In_664);
and U1677 (N_1677,In_784,In_829);
nor U1678 (N_1678,In_288,In_867);
or U1679 (N_1679,In_690,In_37);
nor U1680 (N_1680,In_627,In_931);
xor U1681 (N_1681,In_58,In_810);
nand U1682 (N_1682,In_14,In_558);
nand U1683 (N_1683,In_127,In_365);
and U1684 (N_1684,In_128,In_94);
nor U1685 (N_1685,In_683,In_103);
nor U1686 (N_1686,In_405,In_664);
nand U1687 (N_1687,In_828,In_568);
and U1688 (N_1688,In_994,In_270);
nor U1689 (N_1689,In_817,In_257);
xnor U1690 (N_1690,In_823,In_829);
nor U1691 (N_1691,In_680,In_908);
or U1692 (N_1692,In_406,In_36);
xor U1693 (N_1693,In_945,In_433);
xor U1694 (N_1694,In_146,In_230);
nand U1695 (N_1695,In_523,In_525);
and U1696 (N_1696,In_230,In_314);
or U1697 (N_1697,In_901,In_321);
xnor U1698 (N_1698,In_384,In_433);
and U1699 (N_1699,In_818,In_585);
and U1700 (N_1700,In_104,In_332);
xor U1701 (N_1701,In_77,In_610);
nand U1702 (N_1702,In_431,In_832);
or U1703 (N_1703,In_379,In_131);
nor U1704 (N_1704,In_358,In_254);
nand U1705 (N_1705,In_490,In_870);
and U1706 (N_1706,In_484,In_851);
nand U1707 (N_1707,In_871,In_244);
and U1708 (N_1708,In_745,In_18);
and U1709 (N_1709,In_254,In_667);
xor U1710 (N_1710,In_216,In_412);
nor U1711 (N_1711,In_454,In_857);
or U1712 (N_1712,In_684,In_276);
and U1713 (N_1713,In_931,In_758);
and U1714 (N_1714,In_252,In_713);
nand U1715 (N_1715,In_541,In_473);
nor U1716 (N_1716,In_973,In_717);
nor U1717 (N_1717,In_913,In_91);
nor U1718 (N_1718,In_141,In_734);
xnor U1719 (N_1719,In_841,In_787);
and U1720 (N_1720,In_287,In_925);
xor U1721 (N_1721,In_562,In_323);
nand U1722 (N_1722,In_444,In_370);
or U1723 (N_1723,In_706,In_945);
nand U1724 (N_1724,In_851,In_940);
nor U1725 (N_1725,In_706,In_152);
and U1726 (N_1726,In_128,In_421);
or U1727 (N_1727,In_223,In_719);
or U1728 (N_1728,In_65,In_93);
xor U1729 (N_1729,In_985,In_433);
or U1730 (N_1730,In_390,In_104);
nand U1731 (N_1731,In_418,In_783);
and U1732 (N_1732,In_984,In_181);
nor U1733 (N_1733,In_244,In_319);
or U1734 (N_1734,In_721,In_945);
xnor U1735 (N_1735,In_732,In_505);
nor U1736 (N_1736,In_883,In_736);
and U1737 (N_1737,In_380,In_600);
or U1738 (N_1738,In_471,In_985);
nand U1739 (N_1739,In_3,In_737);
and U1740 (N_1740,In_564,In_400);
nor U1741 (N_1741,In_213,In_923);
nand U1742 (N_1742,In_982,In_763);
nand U1743 (N_1743,In_614,In_357);
nor U1744 (N_1744,In_76,In_787);
xnor U1745 (N_1745,In_718,In_22);
nor U1746 (N_1746,In_824,In_490);
or U1747 (N_1747,In_907,In_393);
or U1748 (N_1748,In_749,In_384);
nor U1749 (N_1749,In_143,In_75);
or U1750 (N_1750,In_70,In_676);
nand U1751 (N_1751,In_121,In_467);
xor U1752 (N_1752,In_488,In_51);
and U1753 (N_1753,In_457,In_770);
and U1754 (N_1754,In_545,In_908);
or U1755 (N_1755,In_172,In_229);
or U1756 (N_1756,In_286,In_232);
nor U1757 (N_1757,In_531,In_67);
or U1758 (N_1758,In_15,In_918);
xnor U1759 (N_1759,In_235,In_441);
nand U1760 (N_1760,In_539,In_78);
or U1761 (N_1761,In_847,In_406);
and U1762 (N_1762,In_393,In_310);
xor U1763 (N_1763,In_629,In_370);
or U1764 (N_1764,In_925,In_895);
xnor U1765 (N_1765,In_132,In_407);
nor U1766 (N_1766,In_526,In_808);
nor U1767 (N_1767,In_800,In_339);
nand U1768 (N_1768,In_73,In_257);
nand U1769 (N_1769,In_106,In_349);
nor U1770 (N_1770,In_83,In_285);
or U1771 (N_1771,In_753,In_966);
or U1772 (N_1772,In_59,In_51);
nand U1773 (N_1773,In_278,In_237);
nor U1774 (N_1774,In_921,In_517);
xnor U1775 (N_1775,In_112,In_308);
and U1776 (N_1776,In_60,In_487);
and U1777 (N_1777,In_506,In_627);
nor U1778 (N_1778,In_557,In_197);
nor U1779 (N_1779,In_663,In_62);
or U1780 (N_1780,In_164,In_770);
nor U1781 (N_1781,In_356,In_632);
and U1782 (N_1782,In_556,In_453);
nor U1783 (N_1783,In_520,In_525);
or U1784 (N_1784,In_290,In_934);
or U1785 (N_1785,In_913,In_768);
and U1786 (N_1786,In_777,In_629);
or U1787 (N_1787,In_686,In_767);
nor U1788 (N_1788,In_762,In_722);
nor U1789 (N_1789,In_772,In_862);
or U1790 (N_1790,In_386,In_586);
nand U1791 (N_1791,In_830,In_6);
and U1792 (N_1792,In_83,In_677);
or U1793 (N_1793,In_170,In_145);
nor U1794 (N_1794,In_480,In_878);
nand U1795 (N_1795,In_561,In_864);
nand U1796 (N_1796,In_41,In_908);
nor U1797 (N_1797,In_784,In_795);
and U1798 (N_1798,In_784,In_725);
nor U1799 (N_1799,In_61,In_763);
nor U1800 (N_1800,In_534,In_265);
xnor U1801 (N_1801,In_613,In_696);
or U1802 (N_1802,In_186,In_715);
or U1803 (N_1803,In_884,In_325);
xnor U1804 (N_1804,In_303,In_992);
nor U1805 (N_1805,In_758,In_972);
nand U1806 (N_1806,In_166,In_733);
or U1807 (N_1807,In_535,In_794);
xor U1808 (N_1808,In_80,In_772);
nor U1809 (N_1809,In_957,In_3);
xnor U1810 (N_1810,In_956,In_8);
nand U1811 (N_1811,In_589,In_738);
xnor U1812 (N_1812,In_339,In_392);
nor U1813 (N_1813,In_94,In_880);
nor U1814 (N_1814,In_315,In_327);
nand U1815 (N_1815,In_814,In_448);
nor U1816 (N_1816,In_609,In_280);
xnor U1817 (N_1817,In_616,In_39);
and U1818 (N_1818,In_926,In_14);
xnor U1819 (N_1819,In_604,In_136);
or U1820 (N_1820,In_289,In_235);
xor U1821 (N_1821,In_101,In_723);
and U1822 (N_1822,In_822,In_884);
nand U1823 (N_1823,In_128,In_677);
xnor U1824 (N_1824,In_316,In_698);
or U1825 (N_1825,In_937,In_397);
nand U1826 (N_1826,In_579,In_249);
nand U1827 (N_1827,In_361,In_791);
or U1828 (N_1828,In_894,In_623);
nor U1829 (N_1829,In_166,In_937);
or U1830 (N_1830,In_618,In_236);
and U1831 (N_1831,In_674,In_461);
xnor U1832 (N_1832,In_481,In_226);
xor U1833 (N_1833,In_282,In_299);
nor U1834 (N_1834,In_32,In_116);
and U1835 (N_1835,In_424,In_62);
xnor U1836 (N_1836,In_404,In_610);
nor U1837 (N_1837,In_718,In_551);
and U1838 (N_1838,In_844,In_878);
nand U1839 (N_1839,In_669,In_626);
and U1840 (N_1840,In_59,In_797);
xor U1841 (N_1841,In_548,In_77);
and U1842 (N_1842,In_914,In_687);
nor U1843 (N_1843,In_755,In_696);
nand U1844 (N_1844,In_4,In_32);
nor U1845 (N_1845,In_40,In_872);
xor U1846 (N_1846,In_21,In_654);
or U1847 (N_1847,In_830,In_787);
xor U1848 (N_1848,In_681,In_792);
nand U1849 (N_1849,In_98,In_193);
or U1850 (N_1850,In_642,In_882);
nor U1851 (N_1851,In_514,In_565);
nand U1852 (N_1852,In_977,In_753);
xnor U1853 (N_1853,In_686,In_143);
and U1854 (N_1854,In_391,In_970);
nor U1855 (N_1855,In_955,In_132);
nor U1856 (N_1856,In_300,In_77);
xnor U1857 (N_1857,In_69,In_284);
xnor U1858 (N_1858,In_228,In_871);
or U1859 (N_1859,In_209,In_470);
xnor U1860 (N_1860,In_861,In_385);
nand U1861 (N_1861,In_458,In_520);
nand U1862 (N_1862,In_233,In_478);
xnor U1863 (N_1863,In_427,In_771);
nand U1864 (N_1864,In_33,In_252);
nand U1865 (N_1865,In_248,In_811);
and U1866 (N_1866,In_127,In_819);
and U1867 (N_1867,In_763,In_824);
xor U1868 (N_1868,In_717,In_208);
nor U1869 (N_1869,In_598,In_113);
xnor U1870 (N_1870,In_648,In_148);
nor U1871 (N_1871,In_752,In_18);
nor U1872 (N_1872,In_474,In_710);
nor U1873 (N_1873,In_686,In_208);
nor U1874 (N_1874,In_99,In_330);
nor U1875 (N_1875,In_754,In_638);
nand U1876 (N_1876,In_109,In_23);
and U1877 (N_1877,In_361,In_450);
nor U1878 (N_1878,In_961,In_496);
nand U1879 (N_1879,In_386,In_27);
or U1880 (N_1880,In_869,In_463);
nand U1881 (N_1881,In_963,In_660);
nand U1882 (N_1882,In_618,In_128);
nand U1883 (N_1883,In_708,In_744);
nand U1884 (N_1884,In_61,In_211);
or U1885 (N_1885,In_85,In_245);
xnor U1886 (N_1886,In_211,In_186);
nor U1887 (N_1887,In_975,In_507);
xor U1888 (N_1888,In_497,In_862);
nand U1889 (N_1889,In_501,In_629);
nand U1890 (N_1890,In_499,In_798);
or U1891 (N_1891,In_864,In_595);
nor U1892 (N_1892,In_501,In_401);
and U1893 (N_1893,In_865,In_224);
and U1894 (N_1894,In_614,In_66);
xnor U1895 (N_1895,In_307,In_559);
or U1896 (N_1896,In_987,In_766);
nor U1897 (N_1897,In_150,In_607);
nor U1898 (N_1898,In_166,In_731);
nor U1899 (N_1899,In_699,In_357);
nor U1900 (N_1900,In_799,In_326);
nand U1901 (N_1901,In_183,In_973);
xnor U1902 (N_1902,In_374,In_154);
and U1903 (N_1903,In_890,In_258);
xnor U1904 (N_1904,In_947,In_794);
nor U1905 (N_1905,In_305,In_56);
nor U1906 (N_1906,In_370,In_939);
and U1907 (N_1907,In_336,In_76);
xor U1908 (N_1908,In_677,In_32);
and U1909 (N_1909,In_518,In_73);
or U1910 (N_1910,In_308,In_472);
xor U1911 (N_1911,In_559,In_548);
or U1912 (N_1912,In_407,In_700);
nor U1913 (N_1913,In_446,In_727);
or U1914 (N_1914,In_137,In_480);
and U1915 (N_1915,In_546,In_513);
xnor U1916 (N_1916,In_838,In_925);
nand U1917 (N_1917,In_801,In_120);
xnor U1918 (N_1918,In_357,In_403);
nor U1919 (N_1919,In_917,In_324);
nand U1920 (N_1920,In_678,In_531);
xor U1921 (N_1921,In_146,In_799);
nand U1922 (N_1922,In_465,In_993);
or U1923 (N_1923,In_922,In_282);
xor U1924 (N_1924,In_755,In_82);
xor U1925 (N_1925,In_295,In_968);
nor U1926 (N_1926,In_206,In_3);
nand U1927 (N_1927,In_174,In_888);
xor U1928 (N_1928,In_26,In_864);
nor U1929 (N_1929,In_919,In_740);
nor U1930 (N_1930,In_638,In_862);
nand U1931 (N_1931,In_942,In_665);
nand U1932 (N_1932,In_346,In_394);
and U1933 (N_1933,In_702,In_620);
nor U1934 (N_1934,In_423,In_123);
nand U1935 (N_1935,In_521,In_50);
or U1936 (N_1936,In_721,In_124);
xnor U1937 (N_1937,In_183,In_125);
and U1938 (N_1938,In_384,In_185);
nor U1939 (N_1939,In_26,In_487);
xor U1940 (N_1940,In_533,In_102);
and U1941 (N_1941,In_540,In_42);
xor U1942 (N_1942,In_845,In_800);
or U1943 (N_1943,In_89,In_498);
nor U1944 (N_1944,In_337,In_609);
and U1945 (N_1945,In_951,In_338);
xor U1946 (N_1946,In_495,In_811);
xnor U1947 (N_1947,In_462,In_920);
or U1948 (N_1948,In_94,In_672);
nor U1949 (N_1949,In_783,In_469);
nor U1950 (N_1950,In_603,In_264);
and U1951 (N_1951,In_632,In_816);
and U1952 (N_1952,In_949,In_615);
nor U1953 (N_1953,In_523,In_867);
or U1954 (N_1954,In_451,In_474);
xnor U1955 (N_1955,In_385,In_894);
nand U1956 (N_1956,In_700,In_515);
or U1957 (N_1957,In_771,In_683);
nand U1958 (N_1958,In_712,In_512);
nand U1959 (N_1959,In_36,In_868);
and U1960 (N_1960,In_761,In_900);
xnor U1961 (N_1961,In_598,In_367);
nor U1962 (N_1962,In_742,In_779);
xor U1963 (N_1963,In_414,In_910);
and U1964 (N_1964,In_965,In_863);
xnor U1965 (N_1965,In_858,In_703);
xor U1966 (N_1966,In_687,In_608);
or U1967 (N_1967,In_383,In_597);
or U1968 (N_1968,In_951,In_754);
and U1969 (N_1969,In_655,In_759);
and U1970 (N_1970,In_862,In_336);
nor U1971 (N_1971,In_602,In_841);
nand U1972 (N_1972,In_965,In_575);
nor U1973 (N_1973,In_163,In_125);
nand U1974 (N_1974,In_721,In_32);
and U1975 (N_1975,In_662,In_909);
xnor U1976 (N_1976,In_685,In_976);
and U1977 (N_1977,In_825,In_955);
and U1978 (N_1978,In_618,In_640);
or U1979 (N_1979,In_656,In_973);
xnor U1980 (N_1980,In_672,In_973);
and U1981 (N_1981,In_87,In_821);
and U1982 (N_1982,In_844,In_122);
nor U1983 (N_1983,In_63,In_337);
xor U1984 (N_1984,In_782,In_219);
nand U1985 (N_1985,In_766,In_442);
nand U1986 (N_1986,In_463,In_9);
xnor U1987 (N_1987,In_884,In_6);
or U1988 (N_1988,In_136,In_610);
or U1989 (N_1989,In_139,In_33);
nand U1990 (N_1990,In_576,In_230);
xnor U1991 (N_1991,In_343,In_71);
or U1992 (N_1992,In_512,In_826);
nor U1993 (N_1993,In_463,In_549);
and U1994 (N_1994,In_792,In_813);
nor U1995 (N_1995,In_383,In_185);
and U1996 (N_1996,In_123,In_221);
nor U1997 (N_1997,In_255,In_65);
xnor U1998 (N_1998,In_37,In_149);
or U1999 (N_1999,In_614,In_752);
or U2000 (N_2000,In_253,In_475);
xnor U2001 (N_2001,In_542,In_455);
nor U2002 (N_2002,In_663,In_948);
xnor U2003 (N_2003,In_538,In_887);
and U2004 (N_2004,In_267,In_571);
or U2005 (N_2005,In_840,In_47);
and U2006 (N_2006,In_8,In_302);
xnor U2007 (N_2007,In_180,In_109);
and U2008 (N_2008,In_376,In_279);
nor U2009 (N_2009,In_595,In_904);
nor U2010 (N_2010,In_543,In_410);
or U2011 (N_2011,In_845,In_756);
and U2012 (N_2012,In_805,In_65);
xor U2013 (N_2013,In_350,In_836);
nand U2014 (N_2014,In_365,In_116);
nor U2015 (N_2015,In_443,In_461);
xnor U2016 (N_2016,In_136,In_501);
nor U2017 (N_2017,In_441,In_238);
nor U2018 (N_2018,In_718,In_565);
or U2019 (N_2019,In_746,In_838);
or U2020 (N_2020,In_643,In_500);
nor U2021 (N_2021,In_151,In_470);
nor U2022 (N_2022,In_523,In_620);
and U2023 (N_2023,In_987,In_593);
and U2024 (N_2024,In_149,In_196);
nand U2025 (N_2025,In_685,In_43);
xnor U2026 (N_2026,In_391,In_957);
xor U2027 (N_2027,In_827,In_103);
and U2028 (N_2028,In_195,In_130);
nor U2029 (N_2029,In_389,In_627);
nor U2030 (N_2030,In_957,In_914);
nor U2031 (N_2031,In_460,In_376);
or U2032 (N_2032,In_919,In_229);
nand U2033 (N_2033,In_661,In_276);
nand U2034 (N_2034,In_111,In_560);
nand U2035 (N_2035,In_221,In_353);
nand U2036 (N_2036,In_555,In_905);
and U2037 (N_2037,In_394,In_605);
nand U2038 (N_2038,In_427,In_881);
and U2039 (N_2039,In_571,In_93);
nand U2040 (N_2040,In_521,In_990);
or U2041 (N_2041,In_444,In_122);
or U2042 (N_2042,In_330,In_861);
or U2043 (N_2043,In_150,In_400);
xor U2044 (N_2044,In_99,In_412);
or U2045 (N_2045,In_127,In_493);
nand U2046 (N_2046,In_479,In_143);
or U2047 (N_2047,In_560,In_182);
xor U2048 (N_2048,In_273,In_565);
xor U2049 (N_2049,In_19,In_673);
xor U2050 (N_2050,In_906,In_348);
nor U2051 (N_2051,In_774,In_452);
nand U2052 (N_2052,In_840,In_669);
nor U2053 (N_2053,In_294,In_375);
or U2054 (N_2054,In_356,In_690);
and U2055 (N_2055,In_599,In_629);
xor U2056 (N_2056,In_140,In_776);
nor U2057 (N_2057,In_340,In_589);
or U2058 (N_2058,In_857,In_937);
xor U2059 (N_2059,In_404,In_792);
or U2060 (N_2060,In_80,In_598);
xor U2061 (N_2061,In_415,In_535);
and U2062 (N_2062,In_248,In_361);
nor U2063 (N_2063,In_387,In_561);
nand U2064 (N_2064,In_410,In_703);
and U2065 (N_2065,In_399,In_787);
nor U2066 (N_2066,In_936,In_230);
nand U2067 (N_2067,In_553,In_210);
or U2068 (N_2068,In_616,In_509);
and U2069 (N_2069,In_589,In_477);
nand U2070 (N_2070,In_436,In_668);
or U2071 (N_2071,In_195,In_441);
nor U2072 (N_2072,In_488,In_431);
or U2073 (N_2073,In_600,In_635);
xnor U2074 (N_2074,In_376,In_621);
or U2075 (N_2075,In_184,In_880);
or U2076 (N_2076,In_248,In_313);
or U2077 (N_2077,In_434,In_72);
and U2078 (N_2078,In_549,In_482);
and U2079 (N_2079,In_192,In_21);
or U2080 (N_2080,In_656,In_690);
or U2081 (N_2081,In_424,In_32);
nor U2082 (N_2082,In_203,In_883);
xor U2083 (N_2083,In_327,In_116);
xnor U2084 (N_2084,In_672,In_827);
nand U2085 (N_2085,In_91,In_435);
nand U2086 (N_2086,In_768,In_229);
or U2087 (N_2087,In_377,In_578);
or U2088 (N_2088,In_717,In_726);
and U2089 (N_2089,In_906,In_229);
xor U2090 (N_2090,In_782,In_758);
or U2091 (N_2091,In_922,In_807);
nand U2092 (N_2092,In_324,In_345);
xor U2093 (N_2093,In_108,In_26);
xor U2094 (N_2094,In_697,In_915);
or U2095 (N_2095,In_192,In_135);
and U2096 (N_2096,In_639,In_724);
nand U2097 (N_2097,In_492,In_322);
and U2098 (N_2098,In_367,In_913);
or U2099 (N_2099,In_403,In_58);
or U2100 (N_2100,In_743,In_419);
or U2101 (N_2101,In_525,In_492);
xnor U2102 (N_2102,In_288,In_1);
nor U2103 (N_2103,In_978,In_906);
nand U2104 (N_2104,In_132,In_557);
or U2105 (N_2105,In_385,In_899);
xor U2106 (N_2106,In_334,In_159);
and U2107 (N_2107,In_900,In_313);
or U2108 (N_2108,In_622,In_537);
nor U2109 (N_2109,In_347,In_490);
nor U2110 (N_2110,In_689,In_795);
and U2111 (N_2111,In_354,In_857);
nand U2112 (N_2112,In_759,In_875);
nor U2113 (N_2113,In_74,In_393);
xor U2114 (N_2114,In_766,In_722);
nand U2115 (N_2115,In_415,In_794);
and U2116 (N_2116,In_485,In_89);
or U2117 (N_2117,In_814,In_398);
xnor U2118 (N_2118,In_884,In_707);
and U2119 (N_2119,In_577,In_202);
and U2120 (N_2120,In_10,In_773);
nor U2121 (N_2121,In_599,In_568);
and U2122 (N_2122,In_317,In_265);
nand U2123 (N_2123,In_510,In_474);
nand U2124 (N_2124,In_231,In_617);
nor U2125 (N_2125,In_920,In_741);
nor U2126 (N_2126,In_806,In_603);
nand U2127 (N_2127,In_441,In_481);
xor U2128 (N_2128,In_124,In_313);
xor U2129 (N_2129,In_909,In_258);
nor U2130 (N_2130,In_811,In_846);
xnor U2131 (N_2131,In_402,In_987);
nor U2132 (N_2132,In_483,In_908);
xor U2133 (N_2133,In_104,In_278);
nor U2134 (N_2134,In_652,In_552);
or U2135 (N_2135,In_618,In_609);
nand U2136 (N_2136,In_578,In_328);
or U2137 (N_2137,In_288,In_797);
and U2138 (N_2138,In_972,In_440);
xor U2139 (N_2139,In_922,In_507);
and U2140 (N_2140,In_172,In_815);
and U2141 (N_2141,In_108,In_435);
or U2142 (N_2142,In_796,In_75);
nor U2143 (N_2143,In_579,In_168);
nor U2144 (N_2144,In_682,In_7);
nand U2145 (N_2145,In_506,In_499);
or U2146 (N_2146,In_493,In_259);
nor U2147 (N_2147,In_132,In_229);
nor U2148 (N_2148,In_755,In_797);
nor U2149 (N_2149,In_422,In_941);
and U2150 (N_2150,In_467,In_266);
or U2151 (N_2151,In_825,In_777);
or U2152 (N_2152,In_790,In_216);
or U2153 (N_2153,In_377,In_658);
or U2154 (N_2154,In_744,In_641);
xnor U2155 (N_2155,In_966,In_908);
and U2156 (N_2156,In_979,In_118);
nor U2157 (N_2157,In_798,In_577);
and U2158 (N_2158,In_84,In_331);
and U2159 (N_2159,In_74,In_235);
or U2160 (N_2160,In_761,In_343);
nor U2161 (N_2161,In_951,In_668);
or U2162 (N_2162,In_959,In_398);
or U2163 (N_2163,In_757,In_412);
nand U2164 (N_2164,In_223,In_591);
xnor U2165 (N_2165,In_95,In_85);
and U2166 (N_2166,In_734,In_245);
and U2167 (N_2167,In_922,In_259);
nand U2168 (N_2168,In_281,In_395);
nor U2169 (N_2169,In_705,In_548);
or U2170 (N_2170,In_373,In_110);
or U2171 (N_2171,In_770,In_303);
and U2172 (N_2172,In_21,In_940);
nor U2173 (N_2173,In_802,In_972);
nand U2174 (N_2174,In_441,In_259);
nor U2175 (N_2175,In_703,In_581);
nor U2176 (N_2176,In_365,In_831);
xor U2177 (N_2177,In_617,In_423);
nor U2178 (N_2178,In_730,In_354);
and U2179 (N_2179,In_653,In_663);
nand U2180 (N_2180,In_486,In_400);
nor U2181 (N_2181,In_853,In_669);
and U2182 (N_2182,In_648,In_283);
nor U2183 (N_2183,In_422,In_872);
nor U2184 (N_2184,In_185,In_490);
and U2185 (N_2185,In_702,In_865);
nor U2186 (N_2186,In_856,In_698);
nor U2187 (N_2187,In_943,In_66);
xnor U2188 (N_2188,In_508,In_150);
nor U2189 (N_2189,In_848,In_416);
or U2190 (N_2190,In_455,In_861);
and U2191 (N_2191,In_884,In_355);
nor U2192 (N_2192,In_337,In_891);
or U2193 (N_2193,In_341,In_450);
or U2194 (N_2194,In_621,In_89);
and U2195 (N_2195,In_842,In_224);
nor U2196 (N_2196,In_296,In_919);
and U2197 (N_2197,In_514,In_228);
nand U2198 (N_2198,In_220,In_451);
and U2199 (N_2199,In_999,In_228);
nor U2200 (N_2200,In_296,In_710);
nand U2201 (N_2201,In_558,In_691);
nor U2202 (N_2202,In_32,In_113);
xnor U2203 (N_2203,In_301,In_108);
and U2204 (N_2204,In_86,In_580);
nand U2205 (N_2205,In_635,In_17);
nor U2206 (N_2206,In_713,In_182);
or U2207 (N_2207,In_335,In_558);
xor U2208 (N_2208,In_286,In_604);
xnor U2209 (N_2209,In_869,In_195);
nand U2210 (N_2210,In_264,In_851);
nand U2211 (N_2211,In_319,In_153);
nand U2212 (N_2212,In_258,In_549);
and U2213 (N_2213,In_323,In_184);
nand U2214 (N_2214,In_215,In_306);
nor U2215 (N_2215,In_481,In_308);
and U2216 (N_2216,In_528,In_6);
nor U2217 (N_2217,In_14,In_44);
and U2218 (N_2218,In_238,In_560);
or U2219 (N_2219,In_995,In_621);
or U2220 (N_2220,In_36,In_197);
or U2221 (N_2221,In_48,In_421);
nand U2222 (N_2222,In_855,In_379);
nand U2223 (N_2223,In_65,In_10);
nand U2224 (N_2224,In_986,In_257);
or U2225 (N_2225,In_576,In_871);
and U2226 (N_2226,In_975,In_967);
xnor U2227 (N_2227,In_322,In_504);
xor U2228 (N_2228,In_13,In_56);
or U2229 (N_2229,In_611,In_248);
nor U2230 (N_2230,In_331,In_966);
xnor U2231 (N_2231,In_352,In_468);
nor U2232 (N_2232,In_796,In_781);
xnor U2233 (N_2233,In_411,In_808);
nand U2234 (N_2234,In_168,In_578);
nor U2235 (N_2235,In_894,In_574);
or U2236 (N_2236,In_531,In_945);
or U2237 (N_2237,In_294,In_3);
and U2238 (N_2238,In_222,In_844);
nand U2239 (N_2239,In_278,In_276);
and U2240 (N_2240,In_368,In_32);
nand U2241 (N_2241,In_338,In_922);
nor U2242 (N_2242,In_592,In_151);
xnor U2243 (N_2243,In_42,In_520);
nor U2244 (N_2244,In_802,In_585);
or U2245 (N_2245,In_138,In_552);
xor U2246 (N_2246,In_208,In_850);
and U2247 (N_2247,In_497,In_127);
xor U2248 (N_2248,In_795,In_173);
nor U2249 (N_2249,In_35,In_319);
nor U2250 (N_2250,In_988,In_728);
or U2251 (N_2251,In_367,In_914);
nand U2252 (N_2252,In_374,In_658);
nand U2253 (N_2253,In_14,In_770);
or U2254 (N_2254,In_774,In_442);
and U2255 (N_2255,In_491,In_270);
or U2256 (N_2256,In_763,In_979);
and U2257 (N_2257,In_35,In_955);
nand U2258 (N_2258,In_301,In_329);
nand U2259 (N_2259,In_819,In_502);
or U2260 (N_2260,In_782,In_657);
nor U2261 (N_2261,In_650,In_101);
or U2262 (N_2262,In_614,In_650);
and U2263 (N_2263,In_432,In_239);
nand U2264 (N_2264,In_833,In_866);
and U2265 (N_2265,In_666,In_254);
nor U2266 (N_2266,In_12,In_101);
xnor U2267 (N_2267,In_371,In_152);
xor U2268 (N_2268,In_75,In_98);
or U2269 (N_2269,In_2,In_773);
nand U2270 (N_2270,In_669,In_87);
and U2271 (N_2271,In_197,In_373);
xnor U2272 (N_2272,In_777,In_618);
or U2273 (N_2273,In_145,In_73);
and U2274 (N_2274,In_501,In_614);
nor U2275 (N_2275,In_288,In_904);
or U2276 (N_2276,In_339,In_511);
nor U2277 (N_2277,In_528,In_248);
or U2278 (N_2278,In_139,In_549);
nor U2279 (N_2279,In_389,In_15);
nor U2280 (N_2280,In_75,In_978);
nor U2281 (N_2281,In_877,In_527);
or U2282 (N_2282,In_216,In_441);
and U2283 (N_2283,In_242,In_446);
xor U2284 (N_2284,In_911,In_156);
nor U2285 (N_2285,In_706,In_412);
nand U2286 (N_2286,In_900,In_52);
or U2287 (N_2287,In_794,In_784);
nor U2288 (N_2288,In_738,In_721);
nand U2289 (N_2289,In_758,In_428);
and U2290 (N_2290,In_996,In_515);
xor U2291 (N_2291,In_701,In_774);
nand U2292 (N_2292,In_325,In_909);
xnor U2293 (N_2293,In_425,In_66);
nand U2294 (N_2294,In_198,In_926);
or U2295 (N_2295,In_150,In_573);
and U2296 (N_2296,In_969,In_445);
nor U2297 (N_2297,In_908,In_821);
xnor U2298 (N_2298,In_470,In_992);
nor U2299 (N_2299,In_556,In_766);
nor U2300 (N_2300,In_670,In_351);
or U2301 (N_2301,In_140,In_569);
nor U2302 (N_2302,In_368,In_638);
nand U2303 (N_2303,In_559,In_682);
nor U2304 (N_2304,In_315,In_711);
xor U2305 (N_2305,In_784,In_311);
nand U2306 (N_2306,In_338,In_881);
and U2307 (N_2307,In_54,In_904);
and U2308 (N_2308,In_632,In_188);
xor U2309 (N_2309,In_706,In_558);
xnor U2310 (N_2310,In_373,In_651);
and U2311 (N_2311,In_359,In_936);
nand U2312 (N_2312,In_188,In_234);
nor U2313 (N_2313,In_601,In_166);
nor U2314 (N_2314,In_112,In_61);
and U2315 (N_2315,In_305,In_303);
or U2316 (N_2316,In_706,In_505);
or U2317 (N_2317,In_956,In_259);
nand U2318 (N_2318,In_160,In_354);
nor U2319 (N_2319,In_971,In_322);
nand U2320 (N_2320,In_657,In_523);
or U2321 (N_2321,In_399,In_97);
nand U2322 (N_2322,In_735,In_414);
or U2323 (N_2323,In_157,In_563);
or U2324 (N_2324,In_61,In_726);
and U2325 (N_2325,In_255,In_897);
or U2326 (N_2326,In_965,In_267);
or U2327 (N_2327,In_372,In_578);
nor U2328 (N_2328,In_480,In_359);
or U2329 (N_2329,In_987,In_231);
nor U2330 (N_2330,In_813,In_828);
nand U2331 (N_2331,In_996,In_567);
or U2332 (N_2332,In_172,In_378);
or U2333 (N_2333,In_136,In_781);
or U2334 (N_2334,In_384,In_199);
nor U2335 (N_2335,In_728,In_640);
nor U2336 (N_2336,In_968,In_468);
or U2337 (N_2337,In_418,In_326);
or U2338 (N_2338,In_575,In_678);
and U2339 (N_2339,In_686,In_806);
xnor U2340 (N_2340,In_891,In_896);
or U2341 (N_2341,In_107,In_665);
and U2342 (N_2342,In_592,In_994);
or U2343 (N_2343,In_197,In_886);
nor U2344 (N_2344,In_159,In_88);
xnor U2345 (N_2345,In_551,In_431);
nand U2346 (N_2346,In_457,In_390);
or U2347 (N_2347,In_307,In_428);
xor U2348 (N_2348,In_990,In_886);
nand U2349 (N_2349,In_288,In_250);
and U2350 (N_2350,In_250,In_811);
xnor U2351 (N_2351,In_415,In_841);
or U2352 (N_2352,In_385,In_461);
or U2353 (N_2353,In_64,In_93);
or U2354 (N_2354,In_847,In_856);
nor U2355 (N_2355,In_332,In_160);
or U2356 (N_2356,In_760,In_518);
or U2357 (N_2357,In_289,In_191);
nand U2358 (N_2358,In_77,In_992);
or U2359 (N_2359,In_210,In_321);
or U2360 (N_2360,In_835,In_428);
or U2361 (N_2361,In_421,In_356);
or U2362 (N_2362,In_846,In_70);
nand U2363 (N_2363,In_739,In_94);
xnor U2364 (N_2364,In_672,In_780);
or U2365 (N_2365,In_168,In_556);
xor U2366 (N_2366,In_816,In_418);
and U2367 (N_2367,In_782,In_819);
and U2368 (N_2368,In_926,In_510);
and U2369 (N_2369,In_46,In_918);
nand U2370 (N_2370,In_696,In_918);
nand U2371 (N_2371,In_34,In_120);
or U2372 (N_2372,In_724,In_132);
nor U2373 (N_2373,In_348,In_563);
xnor U2374 (N_2374,In_46,In_246);
xor U2375 (N_2375,In_283,In_898);
nand U2376 (N_2376,In_174,In_117);
and U2377 (N_2377,In_870,In_781);
nand U2378 (N_2378,In_386,In_867);
nor U2379 (N_2379,In_467,In_940);
or U2380 (N_2380,In_998,In_624);
nand U2381 (N_2381,In_175,In_879);
or U2382 (N_2382,In_787,In_282);
or U2383 (N_2383,In_19,In_169);
or U2384 (N_2384,In_585,In_87);
xor U2385 (N_2385,In_384,In_512);
xnor U2386 (N_2386,In_218,In_466);
or U2387 (N_2387,In_913,In_200);
or U2388 (N_2388,In_589,In_173);
nand U2389 (N_2389,In_120,In_713);
and U2390 (N_2390,In_560,In_128);
and U2391 (N_2391,In_342,In_971);
and U2392 (N_2392,In_702,In_337);
nor U2393 (N_2393,In_40,In_401);
and U2394 (N_2394,In_118,In_260);
xnor U2395 (N_2395,In_113,In_116);
or U2396 (N_2396,In_642,In_483);
nand U2397 (N_2397,In_921,In_232);
and U2398 (N_2398,In_875,In_302);
xnor U2399 (N_2399,In_180,In_389);
nor U2400 (N_2400,In_57,In_650);
xor U2401 (N_2401,In_68,In_637);
xor U2402 (N_2402,In_682,In_315);
nor U2403 (N_2403,In_781,In_530);
and U2404 (N_2404,In_774,In_647);
or U2405 (N_2405,In_43,In_183);
xnor U2406 (N_2406,In_546,In_750);
nand U2407 (N_2407,In_967,In_401);
nand U2408 (N_2408,In_322,In_108);
xor U2409 (N_2409,In_620,In_634);
xnor U2410 (N_2410,In_968,In_989);
xnor U2411 (N_2411,In_547,In_768);
or U2412 (N_2412,In_165,In_213);
or U2413 (N_2413,In_138,In_969);
xor U2414 (N_2414,In_122,In_961);
or U2415 (N_2415,In_415,In_226);
nor U2416 (N_2416,In_511,In_617);
nor U2417 (N_2417,In_304,In_220);
xnor U2418 (N_2418,In_35,In_527);
nor U2419 (N_2419,In_948,In_784);
or U2420 (N_2420,In_276,In_158);
and U2421 (N_2421,In_403,In_391);
or U2422 (N_2422,In_146,In_355);
nor U2423 (N_2423,In_979,In_219);
nand U2424 (N_2424,In_701,In_339);
nand U2425 (N_2425,In_286,In_963);
or U2426 (N_2426,In_574,In_163);
nor U2427 (N_2427,In_865,In_234);
and U2428 (N_2428,In_178,In_138);
nand U2429 (N_2429,In_979,In_336);
xnor U2430 (N_2430,In_311,In_148);
and U2431 (N_2431,In_483,In_455);
nand U2432 (N_2432,In_612,In_518);
nor U2433 (N_2433,In_978,In_392);
nor U2434 (N_2434,In_407,In_824);
xor U2435 (N_2435,In_829,In_848);
nand U2436 (N_2436,In_468,In_994);
nor U2437 (N_2437,In_704,In_523);
nand U2438 (N_2438,In_999,In_676);
nor U2439 (N_2439,In_296,In_352);
or U2440 (N_2440,In_906,In_35);
xor U2441 (N_2441,In_775,In_652);
and U2442 (N_2442,In_281,In_136);
or U2443 (N_2443,In_366,In_270);
nor U2444 (N_2444,In_790,In_531);
nor U2445 (N_2445,In_831,In_639);
xor U2446 (N_2446,In_234,In_999);
nor U2447 (N_2447,In_118,In_464);
or U2448 (N_2448,In_313,In_195);
nor U2449 (N_2449,In_474,In_92);
xnor U2450 (N_2450,In_952,In_770);
xnor U2451 (N_2451,In_345,In_627);
nand U2452 (N_2452,In_537,In_807);
xnor U2453 (N_2453,In_628,In_325);
xnor U2454 (N_2454,In_355,In_468);
xor U2455 (N_2455,In_807,In_824);
or U2456 (N_2456,In_191,In_456);
nor U2457 (N_2457,In_613,In_574);
nand U2458 (N_2458,In_695,In_990);
and U2459 (N_2459,In_913,In_530);
or U2460 (N_2460,In_616,In_638);
or U2461 (N_2461,In_294,In_572);
nand U2462 (N_2462,In_521,In_76);
or U2463 (N_2463,In_436,In_753);
nor U2464 (N_2464,In_850,In_731);
and U2465 (N_2465,In_438,In_537);
or U2466 (N_2466,In_556,In_243);
xnor U2467 (N_2467,In_342,In_497);
xnor U2468 (N_2468,In_401,In_119);
or U2469 (N_2469,In_392,In_212);
nor U2470 (N_2470,In_608,In_557);
or U2471 (N_2471,In_785,In_80);
and U2472 (N_2472,In_469,In_162);
nor U2473 (N_2473,In_566,In_190);
or U2474 (N_2474,In_899,In_534);
and U2475 (N_2475,In_16,In_190);
nor U2476 (N_2476,In_539,In_903);
nand U2477 (N_2477,In_317,In_653);
nor U2478 (N_2478,In_167,In_129);
xor U2479 (N_2479,In_19,In_722);
xnor U2480 (N_2480,In_437,In_597);
nand U2481 (N_2481,In_829,In_591);
xnor U2482 (N_2482,In_563,In_899);
and U2483 (N_2483,In_650,In_726);
and U2484 (N_2484,In_360,In_976);
and U2485 (N_2485,In_825,In_163);
or U2486 (N_2486,In_687,In_666);
nand U2487 (N_2487,In_895,In_203);
xnor U2488 (N_2488,In_216,In_383);
nor U2489 (N_2489,In_917,In_96);
xor U2490 (N_2490,In_732,In_431);
nand U2491 (N_2491,In_362,In_816);
nand U2492 (N_2492,In_609,In_51);
nand U2493 (N_2493,In_589,In_59);
or U2494 (N_2494,In_875,In_457);
nand U2495 (N_2495,In_297,In_673);
and U2496 (N_2496,In_227,In_119);
xor U2497 (N_2497,In_254,In_311);
xnor U2498 (N_2498,In_743,In_816);
nor U2499 (N_2499,In_677,In_68);
nor U2500 (N_2500,N_1563,N_2187);
xor U2501 (N_2501,N_91,N_1378);
nor U2502 (N_2502,N_1309,N_1230);
nand U2503 (N_2503,N_539,N_877);
nand U2504 (N_2504,N_2053,N_1333);
nand U2505 (N_2505,N_1623,N_685);
nor U2506 (N_2506,N_1229,N_2371);
and U2507 (N_2507,N_311,N_383);
and U2508 (N_2508,N_2112,N_887);
xor U2509 (N_2509,N_1792,N_785);
and U2510 (N_2510,N_2195,N_917);
nor U2511 (N_2511,N_1139,N_899);
or U2512 (N_2512,N_2246,N_628);
nand U2513 (N_2513,N_218,N_697);
nand U2514 (N_2514,N_1868,N_2449);
and U2515 (N_2515,N_1736,N_734);
nand U2516 (N_2516,N_2135,N_563);
xnor U2517 (N_2517,N_1488,N_446);
xor U2518 (N_2518,N_2236,N_2490);
xnor U2519 (N_2519,N_2274,N_2466);
or U2520 (N_2520,N_1216,N_1547);
xnor U2521 (N_2521,N_1747,N_1249);
xnor U2522 (N_2522,N_1227,N_12);
or U2523 (N_2523,N_2029,N_935);
nor U2524 (N_2524,N_1921,N_1844);
nand U2525 (N_2525,N_1087,N_864);
xnor U2526 (N_2526,N_469,N_566);
nand U2527 (N_2527,N_773,N_98);
nand U2528 (N_2528,N_2482,N_307);
nand U2529 (N_2529,N_1538,N_1281);
nand U2530 (N_2530,N_950,N_1449);
nand U2531 (N_2531,N_447,N_819);
and U2532 (N_2532,N_1337,N_1317);
nor U2533 (N_2533,N_528,N_989);
xnor U2534 (N_2534,N_1793,N_932);
and U2535 (N_2535,N_1905,N_385);
and U2536 (N_2536,N_1257,N_597);
or U2537 (N_2537,N_1806,N_1602);
and U2538 (N_2538,N_2244,N_1698);
nor U2539 (N_2539,N_1511,N_410);
nor U2540 (N_2540,N_1832,N_2492);
nand U2541 (N_2541,N_1886,N_20);
nor U2542 (N_2542,N_669,N_262);
and U2543 (N_2543,N_2400,N_1579);
nand U2544 (N_2544,N_2476,N_1245);
nor U2545 (N_2545,N_2253,N_127);
nand U2546 (N_2546,N_1759,N_1517);
nand U2547 (N_2547,N_1816,N_1874);
xor U2548 (N_2548,N_1489,N_209);
nand U2549 (N_2549,N_114,N_2457);
or U2550 (N_2550,N_1676,N_1325);
or U2551 (N_2551,N_1758,N_1487);
and U2552 (N_2552,N_776,N_1408);
or U2553 (N_2553,N_691,N_1068);
and U2554 (N_2554,N_2252,N_1721);
nand U2555 (N_2555,N_492,N_1091);
nand U2556 (N_2556,N_987,N_1479);
nand U2557 (N_2557,N_1589,N_329);
or U2558 (N_2558,N_1770,N_1541);
nor U2559 (N_2559,N_1282,N_1319);
xnor U2560 (N_2560,N_1077,N_71);
or U2561 (N_2561,N_1404,N_242);
nor U2562 (N_2562,N_2369,N_0);
nand U2563 (N_2563,N_716,N_2199);
or U2564 (N_2564,N_1653,N_1316);
xnor U2565 (N_2565,N_487,N_2356);
nor U2566 (N_2566,N_2198,N_614);
nand U2567 (N_2567,N_670,N_1671);
or U2568 (N_2568,N_2307,N_738);
nand U2569 (N_2569,N_914,N_1312);
nand U2570 (N_2570,N_580,N_644);
and U2571 (N_2571,N_2342,N_373);
nor U2572 (N_2572,N_1716,N_1358);
xor U2573 (N_2573,N_948,N_2247);
and U2574 (N_2574,N_2407,N_1925);
and U2575 (N_2575,N_1730,N_253);
and U2576 (N_2576,N_1196,N_1284);
nand U2577 (N_2577,N_1145,N_2170);
or U2578 (N_2578,N_207,N_646);
or U2579 (N_2579,N_2145,N_954);
nor U2580 (N_2580,N_305,N_2139);
nand U2581 (N_2581,N_518,N_783);
xnor U2582 (N_2582,N_2264,N_238);
nor U2583 (N_2583,N_2161,N_1565);
nor U2584 (N_2584,N_2041,N_717);
nand U2585 (N_2585,N_1968,N_2431);
nand U2586 (N_2586,N_321,N_757);
nand U2587 (N_2587,N_2385,N_1117);
xor U2588 (N_2588,N_273,N_2470);
or U2589 (N_2589,N_1748,N_46);
or U2590 (N_2590,N_1395,N_1696);
or U2591 (N_2591,N_156,N_1536);
nor U2592 (N_2592,N_713,N_274);
or U2593 (N_2593,N_366,N_549);
and U2594 (N_2594,N_1507,N_266);
nor U2595 (N_2595,N_101,N_2167);
or U2596 (N_2596,N_1013,N_1784);
and U2597 (N_2597,N_2005,N_892);
or U2598 (N_2598,N_1928,N_1867);
or U2599 (N_2599,N_472,N_1761);
xnor U2600 (N_2600,N_2281,N_2233);
and U2601 (N_2601,N_1749,N_1024);
or U2602 (N_2602,N_573,N_1382);
and U2603 (N_2603,N_1750,N_1687);
nor U2604 (N_2604,N_821,N_559);
nand U2605 (N_2605,N_2220,N_1067);
xor U2606 (N_2606,N_22,N_665);
and U2607 (N_2607,N_2339,N_2353);
xor U2608 (N_2608,N_845,N_2294);
or U2609 (N_2609,N_1324,N_1858);
nor U2610 (N_2610,N_2308,N_1185);
and U2611 (N_2611,N_2463,N_17);
or U2612 (N_2612,N_1214,N_1393);
nor U2613 (N_2613,N_2438,N_533);
and U2614 (N_2614,N_379,N_2206);
nor U2615 (N_2615,N_916,N_1963);
nor U2616 (N_2616,N_2079,N_1423);
xor U2617 (N_2617,N_1104,N_416);
and U2618 (N_2618,N_1113,N_289);
xor U2619 (N_2619,N_2212,N_1987);
or U2620 (N_2620,N_687,N_1109);
nor U2621 (N_2621,N_692,N_648);
nand U2622 (N_2622,N_1140,N_286);
nor U2623 (N_2623,N_317,N_949);
nand U2624 (N_2624,N_927,N_1420);
nand U2625 (N_2625,N_89,N_2081);
and U2626 (N_2626,N_1344,N_2332);
and U2627 (N_2627,N_582,N_1752);
and U2628 (N_2628,N_1418,N_1595);
nor U2629 (N_2629,N_2266,N_451);
nand U2630 (N_2630,N_1900,N_116);
or U2631 (N_2631,N_2424,N_1743);
nand U2632 (N_2632,N_1634,N_724);
and U2633 (N_2633,N_1590,N_806);
nor U2634 (N_2634,N_980,N_513);
and U2635 (N_2635,N_995,N_173);
nand U2636 (N_2636,N_2087,N_583);
nor U2637 (N_2637,N_909,N_283);
nand U2638 (N_2638,N_2034,N_88);
and U2639 (N_2639,N_29,N_2372);
xnor U2640 (N_2640,N_831,N_464);
nand U2641 (N_2641,N_1485,N_937);
nor U2642 (N_2642,N_1756,N_777);
xnor U2643 (N_2643,N_1754,N_118);
or U2644 (N_2644,N_970,N_42);
or U2645 (N_2645,N_2046,N_296);
xor U2646 (N_2646,N_394,N_1371);
or U2647 (N_2647,N_710,N_2391);
xnor U2648 (N_2648,N_2306,N_1656);
and U2649 (N_2649,N_2050,N_2100);
or U2650 (N_2650,N_702,N_222);
or U2651 (N_2651,N_2191,N_246);
and U2652 (N_2652,N_1034,N_217);
nor U2653 (N_2653,N_2062,N_1674);
and U2654 (N_2654,N_1052,N_835);
nor U2655 (N_2655,N_371,N_143);
or U2656 (N_2656,N_780,N_2322);
xnor U2657 (N_2657,N_1797,N_43);
and U2658 (N_2658,N_2134,N_141);
xor U2659 (N_2659,N_395,N_468);
and U2660 (N_2660,N_784,N_1992);
nor U2661 (N_2661,N_60,N_1151);
xor U2662 (N_2662,N_1880,N_1470);
xnor U2663 (N_2663,N_766,N_965);
and U2664 (N_2664,N_2288,N_2373);
and U2665 (N_2665,N_1259,N_737);
nand U2666 (N_2666,N_616,N_195);
nor U2667 (N_2667,N_868,N_1913);
nand U2668 (N_2668,N_1019,N_2259);
nand U2669 (N_2669,N_730,N_2317);
nand U2670 (N_2670,N_2418,N_695);
nand U2671 (N_2671,N_2107,N_2299);
nand U2672 (N_2672,N_499,N_2343);
nand U2673 (N_2673,N_2027,N_402);
nand U2674 (N_2674,N_2155,N_789);
nor U2675 (N_2675,N_2061,N_1815);
xnor U2676 (N_2676,N_3,N_2360);
xnor U2677 (N_2677,N_538,N_1801);
nor U2678 (N_2678,N_1247,N_258);
nor U2679 (N_2679,N_2172,N_2284);
xor U2680 (N_2680,N_1457,N_904);
nor U2681 (N_2681,N_2475,N_803);
or U2682 (N_2682,N_1958,N_2464);
or U2683 (N_2683,N_1430,N_1057);
and U2684 (N_2684,N_1646,N_675);
or U2685 (N_2685,N_134,N_1606);
nor U2686 (N_2686,N_558,N_2359);
nand U2687 (N_2687,N_225,N_1296);
xnor U2688 (N_2688,N_1668,N_554);
nor U2689 (N_2689,N_1889,N_928);
and U2690 (N_2690,N_2440,N_1628);
nor U2691 (N_2691,N_983,N_1362);
or U2692 (N_2692,N_1454,N_1381);
and U2693 (N_2693,N_1755,N_1512);
nor U2694 (N_2694,N_411,N_654);
nand U2695 (N_2695,N_1795,N_2309);
xnor U2696 (N_2696,N_363,N_1854);
xnor U2697 (N_2697,N_221,N_1875);
or U2698 (N_2698,N_2150,N_1798);
xnor U2699 (N_2699,N_2403,N_1156);
xnor U2700 (N_2700,N_1675,N_1767);
and U2701 (N_2701,N_991,N_1187);
nor U2702 (N_2702,N_815,N_2228);
nor U2703 (N_2703,N_1008,N_1805);
or U2704 (N_2704,N_753,N_2349);
nand U2705 (N_2705,N_421,N_38);
nand U2706 (N_2706,N_2337,N_1659);
nor U2707 (N_2707,N_1890,N_2311);
and U2708 (N_2708,N_105,N_126);
xnor U2709 (N_2709,N_2346,N_1966);
nand U2710 (N_2710,N_1411,N_1389);
or U2711 (N_2711,N_1321,N_1814);
xor U2712 (N_2712,N_1825,N_1424);
nor U2713 (N_2713,N_2076,N_805);
xor U2714 (N_2714,N_1531,N_2003);
or U2715 (N_2715,N_1225,N_153);
nor U2716 (N_2716,N_512,N_609);
or U2717 (N_2717,N_861,N_1573);
and U2718 (N_2718,N_1335,N_893);
nand U2719 (N_2719,N_1728,N_715);
or U2720 (N_2720,N_546,N_2180);
nand U2721 (N_2721,N_2310,N_1197);
nor U2722 (N_2722,N_1753,N_629);
or U2723 (N_2723,N_2248,N_2009);
xnor U2724 (N_2724,N_1211,N_1283);
nor U2725 (N_2725,N_964,N_1455);
or U2726 (N_2726,N_1045,N_1189);
and U2727 (N_2727,N_1887,N_1345);
and U2728 (N_2728,N_1038,N_684);
xor U2729 (N_2729,N_1846,N_461);
nor U2730 (N_2730,N_1322,N_2217);
xor U2731 (N_2731,N_2125,N_445);
and U2732 (N_2732,N_1932,N_586);
nor U2733 (N_2733,N_519,N_2397);
and U2734 (N_2734,N_723,N_1453);
and U2735 (N_2735,N_1710,N_1069);
xnor U2736 (N_2736,N_2188,N_293);
or U2737 (N_2737,N_921,N_774);
nor U2738 (N_2738,N_2143,N_223);
and U2739 (N_2739,N_701,N_1516);
or U2740 (N_2740,N_2160,N_2133);
nor U2741 (N_2741,N_650,N_393);
xnor U2742 (N_2742,N_2085,N_1560);
nand U2743 (N_2743,N_1372,N_2065);
or U2744 (N_2744,N_457,N_206);
nor U2745 (N_2745,N_1224,N_2096);
nor U2746 (N_2746,N_604,N_1603);
and U2747 (N_2747,N_1501,N_2405);
nand U2748 (N_2748,N_1441,N_2108);
or U2749 (N_2749,N_1678,N_1587);
nand U2750 (N_2750,N_1093,N_210);
and U2751 (N_2751,N_79,N_325);
xnor U2752 (N_2752,N_568,N_10);
nand U2753 (N_2753,N_930,N_2486);
nand U2754 (N_2754,N_1436,N_97);
and U2755 (N_2755,N_352,N_982);
and U2756 (N_2756,N_2347,N_1975);
nor U2757 (N_2757,N_1799,N_2408);
nand U2758 (N_2758,N_889,N_1871);
or U2759 (N_2759,N_709,N_944);
xnor U2760 (N_2760,N_2280,N_1170);
xor U2761 (N_2761,N_2493,N_213);
nor U2762 (N_2762,N_339,N_1592);
and U2763 (N_2763,N_2434,N_1385);
and U2764 (N_2764,N_1359,N_993);
and U2765 (N_2765,N_1369,N_2442);
nand U2766 (N_2766,N_902,N_2304);
nor U2767 (N_2767,N_1964,N_2415);
nand U2768 (N_2768,N_2465,N_1996);
nand U2769 (N_2769,N_1163,N_1570);
nand U2770 (N_2770,N_1435,N_1315);
and U2771 (N_2771,N_1114,N_1202);
and U2772 (N_2772,N_1919,N_2256);
nor U2773 (N_2773,N_2197,N_1561);
or U2774 (N_2774,N_2024,N_618);
nor U2775 (N_2775,N_560,N_2473);
and U2776 (N_2776,N_291,N_1190);
and U2777 (N_2777,N_132,N_1360);
or U2778 (N_2778,N_504,N_2481);
or U2779 (N_2779,N_1556,N_2251);
and U2780 (N_2780,N_630,N_1231);
or U2781 (N_2781,N_1645,N_2093);
nand U2782 (N_2782,N_356,N_2156);
and U2783 (N_2783,N_1270,N_1515);
nand U2784 (N_2784,N_550,N_429);
or U2785 (N_2785,N_163,N_2084);
nand U2786 (N_2786,N_525,N_2377);
or U2787 (N_2787,N_1011,N_1161);
xnor U2788 (N_2788,N_1861,N_1047);
or U2789 (N_2789,N_475,N_340);
xnor U2790 (N_2790,N_219,N_833);
xnor U2791 (N_2791,N_2474,N_1703);
nand U2792 (N_2792,N_256,N_2042);
xnor U2793 (N_2793,N_862,N_1959);
or U2794 (N_2794,N_1251,N_497);
or U2795 (N_2795,N_1707,N_1402);
or U2796 (N_2796,N_1502,N_1461);
and U2797 (N_2797,N_1751,N_1621);
nor U2798 (N_2798,N_1988,N_72);
nor U2799 (N_2799,N_2394,N_2417);
and U2800 (N_2800,N_2268,N_11);
xnor U2801 (N_2801,N_615,N_2092);
nand U2802 (N_2802,N_740,N_400);
and U2803 (N_2803,N_162,N_1734);
nor U2804 (N_2804,N_2401,N_2363);
xnor U2805 (N_2805,N_1810,N_635);
and U2806 (N_2806,N_51,N_1400);
xor U2807 (N_2807,N_761,N_2026);
or U2808 (N_2808,N_590,N_2190);
nand U2809 (N_2809,N_1416,N_1833);
and U2810 (N_2810,N_1374,N_1642);
and U2811 (N_2811,N_2478,N_1285);
or U2812 (N_2812,N_1210,N_1397);
xnor U2813 (N_2813,N_1809,N_1108);
or U2814 (N_2814,N_1204,N_1514);
xnor U2815 (N_2815,N_2113,N_728);
and U2816 (N_2816,N_463,N_1783);
xor U2817 (N_2817,N_1972,N_617);
xor U2818 (N_2818,N_678,N_2293);
xnor U2819 (N_2819,N_631,N_1070);
xnor U2820 (N_2820,N_1533,N_1569);
xor U2821 (N_2821,N_1171,N_1528);
nand U2822 (N_2822,N_1279,N_1119);
or U2823 (N_2823,N_767,N_302);
nand U2824 (N_2824,N_2048,N_413);
xor U2825 (N_2825,N_138,N_2276);
nand U2826 (N_2826,N_460,N_751);
and U2827 (N_2827,N_1226,N_924);
nand U2828 (N_2828,N_2056,N_1931);
nor U2829 (N_2829,N_417,N_2104);
or U2830 (N_2830,N_2402,N_2469);
nand U2831 (N_2831,N_1179,N_1843);
and U2832 (N_2832,N_2144,N_828);
or U2833 (N_2833,N_31,N_945);
xnor U2834 (N_2834,N_1971,N_2207);
xnor U2835 (N_2835,N_1760,N_199);
and U2836 (N_2836,N_287,N_1203);
nand U2837 (N_2837,N_507,N_848);
nand U2838 (N_2838,N_1001,N_1271);
and U2839 (N_2839,N_1215,N_1380);
or U2840 (N_2840,N_1101,N_1513);
and U2841 (N_2841,N_1619,N_1191);
nand U2842 (N_2842,N_1158,N_2324);
or U2843 (N_2843,N_1604,N_735);
and U2844 (N_2844,N_1873,N_365);
nor U2845 (N_2845,N_2498,N_387);
or U2846 (N_2846,N_522,N_2265);
or U2847 (N_2847,N_1437,N_279);
or U2848 (N_2848,N_1732,N_398);
nand U2849 (N_2849,N_659,N_1029);
nand U2850 (N_2850,N_1015,N_432);
nor U2851 (N_2851,N_2215,N_575);
or U2852 (N_2852,N_2254,N_2350);
xnor U2853 (N_2853,N_1403,N_2455);
nand U2854 (N_2854,N_1166,N_64);
nand U2855 (N_2855,N_348,N_2318);
and U2856 (N_2856,N_1276,N_1127);
and U2857 (N_2857,N_235,N_407);
nor U2858 (N_2858,N_1559,N_284);
or U2859 (N_2859,N_375,N_78);
nand U2860 (N_2860,N_2030,N_2389);
or U2861 (N_2861,N_778,N_891);
and U2862 (N_2862,N_1432,N_1320);
xnor U2863 (N_2863,N_1912,N_939);
xnor U2864 (N_2864,N_1148,N_178);
and U2865 (N_2865,N_1291,N_2014);
nor U2866 (N_2866,N_2430,N_2319);
nor U2867 (N_2867,N_39,N_1265);
or U2868 (N_2868,N_2361,N_1818);
nand U2869 (N_2869,N_1834,N_613);
xnor U2870 (N_2870,N_459,N_1338);
nand U2871 (N_2871,N_633,N_61);
nor U2872 (N_2872,N_547,N_869);
xnor U2873 (N_2873,N_1848,N_32);
nor U2874 (N_2874,N_1711,N_2270);
or U2875 (N_2875,N_344,N_190);
or U2876 (N_2876,N_956,N_986);
or U2877 (N_2877,N_1419,N_2448);
xnor U2878 (N_2878,N_1005,N_2095);
nand U2879 (N_2879,N_216,N_294);
and U2880 (N_2880,N_579,N_1938);
nor U2881 (N_2881,N_380,N_2429);
xnor U2882 (N_2882,N_2345,N_1107);
nand U2883 (N_2883,N_1980,N_2458);
nand U2884 (N_2884,N_1597,N_2379);
nor U2885 (N_2885,N_722,N_1121);
nor U2886 (N_2886,N_409,N_224);
nand U2887 (N_2887,N_557,N_1865);
nand U2888 (N_2888,N_1655,N_1280);
nor U2889 (N_2889,N_2086,N_938);
or U2890 (N_2890,N_1268,N_489);
nand U2891 (N_2891,N_2239,N_170);
nor U2892 (N_2892,N_739,N_1260);
xor U2893 (N_2893,N_1327,N_482);
xor U2894 (N_2894,N_233,N_1762);
nor U2895 (N_2895,N_2398,N_1521);
or U2896 (N_2896,N_1974,N_1578);
nand U2897 (N_2897,N_124,N_58);
or U2898 (N_2898,N_1930,N_2058);
nor U2899 (N_2899,N_656,N_50);
and U2900 (N_2900,N_103,N_1099);
nand U2901 (N_2901,N_74,N_2189);
xnor U2902 (N_2902,N_2312,N_414);
nand U2903 (N_2903,N_354,N_2269);
and U2904 (N_2904,N_2219,N_825);
xnor U2905 (N_2905,N_1841,N_2015);
xor U2906 (N_2906,N_943,N_2105);
nand U2907 (N_2907,N_1465,N_106);
and U2908 (N_2908,N_1510,N_164);
or U2909 (N_2909,N_1663,N_1388);
and U2910 (N_2910,N_1680,N_1499);
nor U2911 (N_2911,N_1056,N_2427);
nand U2912 (N_2912,N_2146,N_2016);
nand U2913 (N_2913,N_527,N_1852);
xnor U2914 (N_2914,N_2295,N_683);
or U2915 (N_2915,N_189,N_1774);
or U2916 (N_2916,N_676,N_2071);
or U2917 (N_2917,N_529,N_240);
nand U2918 (N_2918,N_1986,N_186);
nor U2919 (N_2919,N_448,N_2428);
xnor U2920 (N_2920,N_1433,N_1855);
and U2921 (N_2921,N_746,N_1526);
nand U2922 (N_2922,N_688,N_667);
and U2923 (N_2923,N_2049,N_350);
or U2924 (N_2924,N_1136,N_318);
and U2925 (N_2925,N_2376,N_2255);
or U2926 (N_2926,N_2366,N_1950);
or U2927 (N_2927,N_673,N_330);
xnor U2928 (N_2928,N_1994,N_272);
and U2929 (N_2929,N_1049,N_1414);
nor U2930 (N_2930,N_639,N_2227);
or U2931 (N_2931,N_1830,N_435);
or U2932 (N_2932,N_1647,N_1648);
or U2933 (N_2933,N_1851,N_2224);
nor U2934 (N_2934,N_483,N_2432);
xor U2935 (N_2935,N_406,N_800);
and U2936 (N_2936,N_433,N_467);
xor U2937 (N_2937,N_2290,N_1062);
and U2938 (N_2938,N_44,N_1287);
and U2939 (N_2939,N_1175,N_1731);
or U2940 (N_2940,N_1576,N_1879);
or U2941 (N_2941,N_270,N_1450);
nor U2942 (N_2942,N_1105,N_655);
nor U2943 (N_2943,N_1473,N_725);
and U2944 (N_2944,N_1310,N_1791);
nor U2945 (N_2945,N_205,N_841);
nand U2946 (N_2946,N_1872,N_2127);
and U2947 (N_2947,N_2314,N_1115);
xor U2948 (N_2948,N_2173,N_1464);
nand U2949 (N_2949,N_193,N_1033);
nand U2950 (N_2950,N_1920,N_1278);
nor U2951 (N_2951,N_2148,N_1857);
and U2952 (N_2952,N_686,N_1976);
or U2953 (N_2953,N_1244,N_2211);
and U2954 (N_2954,N_896,N_920);
nand U2955 (N_2955,N_1012,N_2454);
xor U2956 (N_2956,N_1662,N_929);
nor U2957 (N_2957,N_1134,N_1486);
or U2958 (N_2958,N_1869,N_754);
nor U2959 (N_2959,N_1209,N_1532);
nand U2960 (N_2960,N_80,N_49);
nand U2961 (N_2961,N_2320,N_601);
nor U2962 (N_2962,N_2203,N_2077);
nand U2963 (N_2963,N_2140,N_1817);
nand U2964 (N_2964,N_1347,N_727);
and U2965 (N_2965,N_622,N_1688);
xor U2966 (N_2966,N_1295,N_2262);
nor U2967 (N_2967,N_337,N_1631);
nor U2968 (N_2968,N_1535,N_1629);
nor U2969 (N_2969,N_2232,N_2132);
xnor U2970 (N_2970,N_1933,N_1723);
nand U2971 (N_2971,N_1415,N_1443);
xor U2972 (N_2972,N_2285,N_741);
xor U2973 (N_2973,N_359,N_1738);
xor U2974 (N_2974,N_2040,N_1496);
nand U2975 (N_2975,N_1735,N_82);
and U2976 (N_2976,N_775,N_1159);
nor U2977 (N_2977,N_1949,N_2151);
nand U2978 (N_2978,N_1907,N_1220);
nand U2979 (N_2979,N_45,N_649);
xor U2980 (N_2980,N_1083,N_1222);
nor U2981 (N_2981,N_588,N_1406);
xnor U2982 (N_2982,N_1088,N_1788);
nand U2983 (N_2983,N_752,N_719);
or U2984 (N_2984,N_1258,N_1670);
nor U2985 (N_2985,N_1639,N_1314);
xor U2986 (N_2986,N_281,N_1304);
xnor U2987 (N_2987,N_158,N_1553);
nand U2988 (N_2988,N_1059,N_47);
nor U2989 (N_2989,N_2047,N_2450);
and U2990 (N_2990,N_133,N_2396);
nand U2991 (N_2991,N_574,N_436);
nand U2992 (N_2992,N_595,N_2018);
nor U2993 (N_2993,N_690,N_56);
xor U2994 (N_2994,N_1583,N_768);
or U2995 (N_2995,N_802,N_962);
xnor U2996 (N_2996,N_992,N_931);
xnor U2997 (N_2997,N_641,N_30);
nor U2998 (N_2998,N_1456,N_257);
nand U2999 (N_2999,N_677,N_1769);
nor U3000 (N_3000,N_1383,N_8);
nor U3001 (N_3001,N_1348,N_1041);
nand U3002 (N_3002,N_376,N_1914);
and U3003 (N_3003,N_1956,N_1891);
xor U3004 (N_3004,N_1878,N_2485);
nand U3005 (N_3005,N_555,N_2334);
xor U3006 (N_3006,N_1635,N_96);
xnor U3007 (N_3007,N_1174,N_420);
xnor U3008 (N_3008,N_1010,N_374);
and U3009 (N_3009,N_922,N_144);
and U3010 (N_3010,N_1458,N_2067);
xnor U3011 (N_3011,N_1398,N_494);
nor U3012 (N_3012,N_1819,N_1842);
or U3013 (N_3013,N_2447,N_506);
nor U3014 (N_3014,N_2181,N_2064);
and U3015 (N_3015,N_1060,N_2202);
or U3016 (N_3016,N_215,N_439);
xor U3017 (N_3017,N_2157,N_1706);
or U3018 (N_3018,N_336,N_2163);
xor U3019 (N_3019,N_1079,N_2002);
or U3020 (N_3020,N_48,N_1352);
nand U3021 (N_3021,N_1684,N_1394);
xnor U3022 (N_3022,N_2165,N_1906);
nand U3023 (N_3023,N_227,N_661);
or U3024 (N_3024,N_894,N_427);
nor U3025 (N_3025,N_820,N_1413);
xnor U3026 (N_3026,N_1575,N_229);
xor U3027 (N_3027,N_90,N_1445);
nor U3028 (N_3028,N_1452,N_1474);
nor U3029 (N_3029,N_2273,N_171);
xor U3030 (N_3030,N_1981,N_817);
and U3031 (N_3031,N_2193,N_794);
and U3032 (N_3032,N_1048,N_1255);
or U3033 (N_3033,N_2439,N_2278);
xor U3034 (N_3034,N_2487,N_16);
nor U3035 (N_3035,N_157,N_1772);
and U3036 (N_3036,N_1742,N_634);
nand U3037 (N_3037,N_540,N_1290);
and U3038 (N_3038,N_57,N_1591);
or U3039 (N_3039,N_1129,N_1112);
xnor U3040 (N_3040,N_23,N_107);
nand U3041 (N_3041,N_1026,N_578);
nor U3042 (N_3042,N_2326,N_2028);
xnor U3043 (N_3043,N_1942,N_2351);
xor U3044 (N_3044,N_424,N_2072);
and U3045 (N_3045,N_7,N_1982);
nor U3046 (N_3046,N_405,N_589);
and U3047 (N_3047,N_2433,N_338);
and U3048 (N_3048,N_501,N_1692);
nor U3049 (N_3049,N_760,N_1686);
nand U3050 (N_3050,N_1935,N_382);
nor U3051 (N_3051,N_859,N_1522);
or U3052 (N_3052,N_838,N_357);
or U3053 (N_3053,N_2336,N_750);
xnor U3054 (N_3054,N_1776,N_1241);
or U3055 (N_3055,N_315,N_372);
xor U3056 (N_3056,N_389,N_1529);
xor U3057 (N_3057,N_1167,N_796);
or U3058 (N_3058,N_2245,N_2499);
and U3059 (N_3059,N_997,N_1654);
xnor U3060 (N_3060,N_1835,N_179);
nand U3061 (N_3061,N_2162,N_470);
nor U3062 (N_3062,N_1697,N_1796);
nand U3063 (N_3063,N_154,N_312);
xnor U3064 (N_3064,N_1340,N_1970);
and U3065 (N_3065,N_147,N_152);
nand U3066 (N_3066,N_25,N_1000);
nand U3067 (N_3067,N_689,N_810);
nand U3068 (N_3068,N_985,N_769);
nand U3069 (N_3069,N_812,N_292);
nand U3070 (N_3070,N_941,N_1745);
and U3071 (N_3071,N_28,N_181);
nor U3072 (N_3072,N_721,N_1803);
xnor U3073 (N_3073,N_816,N_886);
and U3074 (N_3074,N_1401,N_2277);
xnor U3075 (N_3075,N_425,N_975);
nand U3076 (N_3076,N_1995,N_1076);
and U3077 (N_3077,N_1650,N_882);
and U3078 (N_3078,N_493,N_1409);
nand U3079 (N_3079,N_75,N_1263);
nor U3080 (N_3080,N_2069,N_392);
nor U3081 (N_3081,N_1807,N_779);
xor U3082 (N_3082,N_1331,N_984);
or U3083 (N_3083,N_860,N_1286);
and U3084 (N_3084,N_2364,N_1585);
nor U3085 (N_3085,N_241,N_624);
or U3086 (N_3086,N_1120,N_129);
nand U3087 (N_3087,N_2213,N_2395);
or U3088 (N_3088,N_718,N_309);
nand U3089 (N_3089,N_703,N_883);
or U3090 (N_3090,N_1657,N_2289);
xor U3091 (N_3091,N_936,N_1699);
xor U3092 (N_3092,N_341,N_2249);
and U3093 (N_3093,N_1375,N_1192);
and U3094 (N_3094,N_1491,N_818);
and U3095 (N_3095,N_905,N_1839);
or U3096 (N_3096,N_2001,N_1882);
nor U3097 (N_3097,N_1941,N_155);
xnor U3098 (N_3098,N_1272,N_2461);
nand U3099 (N_3099,N_1665,N_553);
or U3100 (N_3100,N_1440,N_150);
nor U3101 (N_3101,N_1789,N_1468);
xnor U3102 (N_3102,N_1764,N_576);
nor U3103 (N_3103,N_1078,N_1178);
nor U3104 (N_3104,N_1106,N_2216);
or U3105 (N_3105,N_1664,N_581);
or U3106 (N_3106,N_303,N_1638);
or U3107 (N_3107,N_1143,N_1035);
nand U3108 (N_3108,N_93,N_790);
or U3109 (N_3109,N_264,N_2128);
nand U3110 (N_3110,N_2021,N_2226);
nand U3111 (N_3111,N_1630,N_131);
nor U3112 (N_3112,N_960,N_1110);
nor U3113 (N_3113,N_822,N_1864);
or U3114 (N_3114,N_1626,N_1460);
nand U3115 (N_3115,N_636,N_708);
or U3116 (N_3116,N_1918,N_254);
and U3117 (N_3117,N_732,N_2025);
nor U3118 (N_3118,N_537,N_571);
nor U3119 (N_3119,N_214,N_1572);
or U3120 (N_3120,N_895,N_1594);
xor U3121 (N_3121,N_367,N_807);
nor U3122 (N_3122,N_1566,N_1096);
and U3123 (N_3123,N_1346,N_19);
xor U3124 (N_3124,N_1885,N_2238);
nand U3125 (N_3125,N_2411,N_1896);
xor U3126 (N_3126,N_1182,N_1787);
xor U3127 (N_3127,N_749,N_62);
nand U3128 (N_3128,N_1548,N_251);
nand U3129 (N_3129,N_73,N_1219);
nor U3130 (N_3130,N_1082,N_396);
nor U3131 (N_3131,N_663,N_1823);
and U3132 (N_3132,N_165,N_2240);
and U3133 (N_3133,N_1677,N_349);
xnor U3134 (N_3134,N_1781,N_2036);
nor U3135 (N_3135,N_1739,N_1527);
nand U3136 (N_3136,N_2393,N_236);
nand U3137 (N_3137,N_2111,N_1520);
nor U3138 (N_3138,N_2102,N_592);
nand U3139 (N_3139,N_2088,N_1102);
and U3140 (N_3140,N_1275,N_1624);
xnor U3141 (N_3141,N_2422,N_1138);
and U3142 (N_3142,N_953,N_569);
or U3143 (N_3143,N_1307,N_110);
or U3144 (N_3144,N_1016,N_1269);
nor U3145 (N_3145,N_2459,N_1826);
nand U3146 (N_3146,N_2222,N_1644);
nand U3147 (N_3147,N_1357,N_364);
xor U3148 (N_3148,N_1612,N_174);
nand U3149 (N_3149,N_1558,N_2115);
and U3150 (N_3150,N_1303,N_450);
or U3151 (N_3151,N_878,N_1822);
and U3152 (N_3152,N_1695,N_188);
nor U3153 (N_3153,N_1355,N_1926);
nor U3154 (N_3154,N_1252,N_1961);
nand U3155 (N_3155,N_68,N_473);
or U3156 (N_3156,N_484,N_2022);
nand U3157 (N_3157,N_377,N_2164);
xnor U3158 (N_3158,N_515,N_598);
xor U3159 (N_3159,N_1944,N_2119);
and U3160 (N_3160,N_2054,N_1407);
and U3161 (N_3161,N_204,N_1977);
xnor U3162 (N_3162,N_747,N_2380);
nand U3163 (N_3163,N_857,N_1899);
xnor U3164 (N_3164,N_2443,N_671);
and U3165 (N_3165,N_1552,N_1218);
and U3166 (N_3166,N_1044,N_1555);
or U3167 (N_3167,N_607,N_95);
nor U3168 (N_3168,N_840,N_632);
or U3169 (N_3169,N_2169,N_2330);
and U3170 (N_3170,N_1543,N_1534);
and U3171 (N_3171,N_187,N_1051);
nor U3172 (N_3172,N_1238,N_541);
and U3173 (N_3173,N_517,N_2384);
nor U3174 (N_3174,N_220,N_1600);
nand U3175 (N_3175,N_781,N_2044);
xor U3176 (N_3176,N_1153,N_1997);
nand U3177 (N_3177,N_2329,N_1386);
nor U3178 (N_3178,N_1608,N_1652);
xor U3179 (N_3179,N_606,N_552);
and U3180 (N_3180,N_422,N_263);
xor U3181 (N_3181,N_1545,N_1160);
xnor U3182 (N_3182,N_486,N_1953);
nand U3183 (N_3183,N_1392,N_1544);
nor U3184 (N_3184,N_1475,N_37);
and U3185 (N_3185,N_2416,N_477);
or U3186 (N_3186,N_925,N_465);
xor U3187 (N_3187,N_1042,N_2365);
and U3188 (N_3188,N_2007,N_942);
nor U3189 (N_3189,N_1353,N_798);
or U3190 (N_3190,N_2419,N_957);
or U3191 (N_3191,N_508,N_770);
nand U3192 (N_3192,N_743,N_1651);
and U3193 (N_3193,N_1037,N_345);
xnor U3194 (N_3194,N_626,N_971);
and U3195 (N_3195,N_1361,N_100);
nand U3196 (N_3196,N_1633,N_1632);
xnor U3197 (N_3197,N_1162,N_1326);
and U3198 (N_3198,N_1999,N_121);
and U3199 (N_3199,N_587,N_125);
or U3200 (N_3200,N_1080,N_1828);
nor U3201 (N_3201,N_1240,N_196);
and U3202 (N_3202,N_1542,N_2328);
and U3203 (N_3203,N_681,N_182);
and U3204 (N_3204,N_764,N_961);
and U3205 (N_3205,N_1298,N_444);
or U3206 (N_3206,N_1990,N_1838);
nor U3207 (N_3207,N_1622,N_1757);
nand U3208 (N_3208,N_1794,N_652);
nor U3209 (N_3209,N_1292,N_787);
xor U3210 (N_3210,N_197,N_1863);
and U3211 (N_3211,N_478,N_1773);
or U3212 (N_3212,N_551,N_1613);
xnor U3213 (N_3213,N_2413,N_314);
nand U3214 (N_3214,N_1934,N_1264);
nand U3215 (N_3215,N_1733,N_1494);
nor U3216 (N_3216,N_384,N_854);
xor U3217 (N_3217,N_832,N_63);
xor U3218 (N_3218,N_1682,N_1718);
and U3219 (N_3219,N_2286,N_1596);
or U3220 (N_3220,N_842,N_1130);
nor U3221 (N_3221,N_245,N_2296);
nand U3222 (N_3222,N_612,N_608);
xnor U3223 (N_3223,N_353,N_1387);
nor U3224 (N_3224,N_912,N_645);
nand U3225 (N_3225,N_1336,N_521);
and U3226 (N_3226,N_998,N_1500);
and U3227 (N_3227,N_947,N_280);
or U3228 (N_3228,N_2176,N_1615);
and U3229 (N_3229,N_1176,N_449);
nand U3230 (N_3230,N_1169,N_1993);
xor U3231 (N_3231,N_27,N_175);
or U3232 (N_3232,N_177,N_1658);
nor U3233 (N_3233,N_865,N_1356);
nor U3234 (N_3234,N_86,N_1800);
xnor U3235 (N_3235,N_1379,N_584);
or U3236 (N_3236,N_919,N_1448);
nor U3237 (N_3237,N_355,N_275);
xnor U3238 (N_3238,N_875,N_423);
and U3239 (N_3239,N_874,N_1582);
nand U3240 (N_3240,N_1039,N_1952);
nor U3241 (N_3241,N_53,N_2472);
or U3242 (N_3242,N_2467,N_2420);
and U3243 (N_3243,N_347,N_1277);
xor U3244 (N_3244,N_55,N_167);
nand U3245 (N_3245,N_672,N_35);
or U3246 (N_3246,N_610,N_1288);
and U3247 (N_3247,N_2260,N_999);
or U3248 (N_3248,N_706,N_2099);
and U3249 (N_3249,N_1827,N_208);
nand U3250 (N_3250,N_327,N_1701);
xnor U3251 (N_3251,N_1683,N_334);
or U3252 (N_3252,N_638,N_1998);
nand U3253 (N_3253,N_1313,N_1421);
xor U3254 (N_3254,N_2231,N_1601);
xnor U3255 (N_3255,N_866,N_2019);
nor U3256 (N_3256,N_978,N_694);
nand U3257 (N_3257,N_443,N_1365);
xor U3258 (N_3258,N_1717,N_1232);
nor U3259 (N_3259,N_250,N_1482);
or U3260 (N_3260,N_2272,N_2074);
and U3261 (N_3261,N_1812,N_969);
xor U3262 (N_3262,N_362,N_1866);
xnor U3263 (N_3263,N_1412,N_1574);
xor U3264 (N_3264,N_2083,N_1343);
xor U3265 (N_3265,N_1539,N_2315);
nor U3266 (N_3266,N_1128,N_159);
nand U3267 (N_3267,N_282,N_1962);
or U3268 (N_3268,N_2243,N_627);
and U3269 (N_3269,N_13,N_748);
xor U3270 (N_3270,N_109,N_83);
nand U3271 (N_3271,N_1154,N_603);
xnor U3272 (N_3272,N_1431,N_591);
and U3273 (N_3273,N_1092,N_94);
or U3274 (N_3274,N_698,N_1031);
nor U3275 (N_3275,N_903,N_853);
nor U3276 (N_3276,N_370,N_1205);
or U3277 (N_3277,N_788,N_813);
nor U3278 (N_3278,N_850,N_834);
xor U3279 (N_3279,N_531,N_1261);
and U3280 (N_3280,N_1235,N_1085);
and U3281 (N_3281,N_2441,N_2103);
nand U3282 (N_3282,N_2383,N_452);
xnor U3283 (N_3283,N_2109,N_2031);
and U3284 (N_3284,N_2382,N_705);
xnor U3285 (N_3285,N_1895,N_2480);
nor U3286 (N_3286,N_602,N_731);
xnor U3287 (N_3287,N_2409,N_1332);
nor U3288 (N_3288,N_1061,N_399);
xor U3289 (N_3289,N_1116,N_1493);
or U3290 (N_3290,N_2000,N_804);
or U3291 (N_3291,N_434,N_1429);
or U3292 (N_3292,N_111,N_1133);
xor U3293 (N_3293,N_1540,N_1122);
or U3294 (N_3294,N_1929,N_2179);
nand U3295 (N_3295,N_1877,N_168);
xnor U3296 (N_3296,N_1323,N_756);
and U3297 (N_3297,N_2267,N_1765);
nor U3298 (N_3298,N_879,N_1065);
and U3299 (N_3299,N_801,N_276);
and U3300 (N_3300,N_1146,N_136);
xor U3301 (N_3301,N_1447,N_139);
nand U3302 (N_3302,N_2341,N_2237);
or U3303 (N_3303,N_623,N_4);
nor U3304 (N_3304,N_933,N_1367);
and U3305 (N_3305,N_990,N_298);
nand U3306 (N_3306,N_117,N_268);
nand U3307 (N_3307,N_1020,N_1704);
xnor U3308 (N_3308,N_403,N_401);
xor U3309 (N_3309,N_194,N_1168);
and U3310 (N_3310,N_1442,N_973);
nand U3311 (N_3311,N_1551,N_1318);
nor U3312 (N_3312,N_1937,N_1186);
nand U3313 (N_3313,N_1266,N_476);
nand U3314 (N_3314,N_169,N_1207);
or U3315 (N_3315,N_918,N_2182);
nor U3316 (N_3316,N_66,N_923);
nor U3317 (N_3317,N_2070,N_1973);
and U3318 (N_3318,N_1439,N_2392);
nor U3319 (N_3319,N_1546,N_77);
nor U3320 (N_3320,N_2292,N_1965);
or U3321 (N_3321,N_34,N_243);
nor U3322 (N_3322,N_1308,N_2234);
nor U3323 (N_3323,N_898,N_1046);
nand U3324 (N_3324,N_1236,N_261);
and U3325 (N_3325,N_1405,N_509);
and U3326 (N_3326,N_271,N_824);
and U3327 (N_3327,N_1273,N_959);
nor U3328 (N_3328,N_113,N_2137);
and U3329 (N_3329,N_1009,N_2123);
xor U3330 (N_3330,N_765,N_2208);
and U3331 (N_3331,N_54,N_1525);
nor U3332 (N_3332,N_1428,N_323);
nor U3333 (N_3333,N_2357,N_977);
and U3334 (N_3334,N_1094,N_277);
or U3335 (N_3335,N_1021,N_2352);
nor U3336 (N_3336,N_981,N_85);
or U3337 (N_3337,N_1208,N_510);
nor U3338 (N_3338,N_1804,N_530);
and U3339 (N_3339,N_1125,N_1763);
nor U3340 (N_3340,N_585,N_2147);
nand U3341 (N_3341,N_2090,N_1084);
and U3342 (N_3342,N_1672,N_1893);
xnor U3343 (N_3343,N_2124,N_1685);
or U3344 (N_3344,N_1911,N_1666);
and U3345 (N_3345,N_2425,N_397);
or U3346 (N_3346,N_2287,N_570);
xor U3347 (N_3347,N_1715,N_593);
and U3348 (N_3348,N_596,N_260);
xnor U3349 (N_3349,N_21,N_1840);
and U3350 (N_3350,N_1847,N_711);
and U3351 (N_3351,N_658,N_1775);
nand U3352 (N_3352,N_1860,N_430);
xnor U3353 (N_3353,N_2479,N_1228);
or U3354 (N_3354,N_1599,N_1778);
nand U3355 (N_3355,N_2210,N_1845);
nor U3356 (N_3356,N_1302,N_232);
nand U3357 (N_3357,N_1713,N_1097);
or U3358 (N_3358,N_33,N_481);
nor U3359 (N_3359,N_1299,N_1649);
nand U3360 (N_3360,N_1616,N_870);
or U3361 (N_3361,N_926,N_2120);
or U3362 (N_3362,N_1262,N_599);
nand U3363 (N_3363,N_316,N_619);
or U3364 (N_3364,N_852,N_1055);
xnor U3365 (N_3365,N_1495,N_346);
nand U3366 (N_3366,N_542,N_2488);
or U3367 (N_3367,N_1329,N_1853);
nand U3368 (N_3368,N_881,N_600);
xor U3369 (N_3369,N_1714,N_908);
nand U3370 (N_3370,N_474,N_1267);
nand U3371 (N_3371,N_1377,N_1476);
and U3372 (N_3372,N_1425,N_1892);
or U3373 (N_3373,N_647,N_637);
and U3374 (N_3374,N_1484,N_1111);
nor U3375 (N_3375,N_498,N_1184);
nor U3376 (N_3376,N_2325,N_906);
nand U3377 (N_3377,N_1777,N_958);
and U3378 (N_3378,N_2126,N_826);
nor U3379 (N_3379,N_1193,N_556);
nand U3380 (N_3380,N_2153,N_1720);
or U3381 (N_3381,N_368,N_2250);
nor U3382 (N_3382,N_2032,N_733);
or U3383 (N_3383,N_799,N_1519);
nor U3384 (N_3384,N_1050,N_331);
xnor U3385 (N_3385,N_1562,N_76);
nor U3386 (N_3386,N_288,N_1581);
or U3387 (N_3387,N_1350,N_332);
nand U3388 (N_3388,N_2390,N_1472);
nor U3389 (N_3389,N_1177,N_145);
xnor U3390 (N_3390,N_1915,N_122);
xor U3391 (N_3391,N_2279,N_811);
nor U3392 (N_3392,N_2241,N_1691);
or U3393 (N_3393,N_762,N_1144);
nor U3394 (N_3394,N_543,N_2039);
and U3395 (N_3395,N_836,N_668);
nor U3396 (N_3396,N_2406,N_1212);
nor U3397 (N_3397,N_2313,N_161);
or U3398 (N_3398,N_2175,N_172);
and U3399 (N_3399,N_1233,N_1480);
or U3400 (N_3400,N_2082,N_437);
nor U3401 (N_3401,N_1640,N_577);
nand U3402 (N_3402,N_2381,N_1422);
xor U3403 (N_3403,N_87,N_2075);
nand U3404 (N_3404,N_809,N_2333);
nand U3405 (N_3405,N_1923,N_736);
or U3406 (N_3406,N_1984,N_795);
and U3407 (N_3407,N_2423,N_2462);
xnor U3408 (N_3408,N_2444,N_1478);
and U3409 (N_3409,N_901,N_1983);
nand U3410 (N_3410,N_712,N_505);
nand U3411 (N_3411,N_2271,N_1341);
and U3412 (N_3412,N_491,N_1253);
and U3413 (N_3413,N_128,N_1064);
nand U3414 (N_3414,N_1618,N_200);
and U3415 (N_3415,N_1242,N_1213);
nor U3416 (N_3416,N_1836,N_2331);
and U3417 (N_3417,N_2141,N_2106);
nor U3418 (N_3418,N_2177,N_1504);
xnor U3419 (N_3419,N_2037,N_1368);
xor U3420 (N_3420,N_1066,N_15);
xor U3421 (N_3421,N_1780,N_1802);
and U3422 (N_3422,N_462,N_1030);
or U3423 (N_3423,N_1201,N_2205);
nor U3424 (N_3424,N_1311,N_666);
nor U3425 (N_3425,N_69,N_704);
xor U3426 (N_3426,N_976,N_640);
xor U3427 (N_3427,N_745,N_1903);
xnor U3428 (N_3428,N_2185,N_707);
nand U3429 (N_3429,N_2184,N_2235);
xnor U3430 (N_3430,N_115,N_2321);
nor U3431 (N_3431,N_1702,N_782);
nand U3432 (N_3432,N_1681,N_2158);
and U3433 (N_3433,N_1689,N_1927);
and U3434 (N_3434,N_404,N_1342);
or U3435 (N_3435,N_680,N_1779);
or U3436 (N_3436,N_1924,N_351);
xnor U3437 (N_3437,N_2004,N_1813);
xnor U3438 (N_3438,N_166,N_142);
xnor U3439 (N_3439,N_2221,N_2223);
nor U3440 (N_3440,N_2456,N_1550);
or U3441 (N_3441,N_1014,N_202);
nand U3442 (N_3442,N_1741,N_2043);
nor U3443 (N_3443,N_440,N_2121);
xor U3444 (N_3444,N_471,N_2200);
or U3445 (N_3445,N_1506,N_1364);
xor U3446 (N_3446,N_108,N_26);
xnor U3447 (N_3447,N_1712,N_791);
nor U3448 (N_3448,N_534,N_532);
and U3449 (N_3449,N_2283,N_2011);
nand U3450 (N_3450,N_1945,N_228);
nor U3451 (N_3451,N_2495,N_319);
nand U3452 (N_3452,N_1947,N_1894);
nor U3453 (N_3453,N_1137,N_290);
nand U3454 (N_3454,N_1157,N_310);
nor U3455 (N_3455,N_562,N_548);
xnor U3456 (N_3456,N_1274,N_24);
and U3457 (N_3457,N_1881,N_1571);
nand U3458 (N_3458,N_2477,N_304);
nand U3459 (N_3459,N_285,N_2300);
nor U3460 (N_3460,N_1523,N_70);
or U3461 (N_3461,N_1549,N_180);
nor U3462 (N_3462,N_1577,N_1444);
and U3463 (N_3463,N_1090,N_1567);
and U3464 (N_3464,N_40,N_1217);
and U3465 (N_3465,N_726,N_1916);
and U3466 (N_3466,N_1849,N_2152);
or U3467 (N_3467,N_2225,N_1305);
xor U3468 (N_3468,N_2305,N_1611);
nor U3469 (N_3469,N_843,N_2275);
or U3470 (N_3470,N_979,N_1370);
nor U3471 (N_3471,N_1605,N_1301);
or U3472 (N_3472,N_2006,N_2483);
nor U3473 (N_3473,N_1991,N_2362);
or U3474 (N_3474,N_2435,N_2412);
and U3475 (N_3475,N_1985,N_2129);
or U3476 (N_3476,N_849,N_2059);
or U3477 (N_3477,N_2340,N_84);
or U3478 (N_3478,N_104,N_2387);
xnor U3479 (N_3479,N_1198,N_2209);
xor U3480 (N_3480,N_342,N_1607);
nand U3481 (N_3481,N_381,N_36);
or U3482 (N_3482,N_758,N_1584);
xor U3483 (N_3483,N_2370,N_1248);
or U3484 (N_3484,N_5,N_565);
nand U3485 (N_3485,N_1859,N_1155);
xor U3486 (N_3486,N_2055,N_2078);
or U3487 (N_3487,N_847,N_1625);
nor U3488 (N_3488,N_1366,N_1498);
and U3489 (N_3489,N_1123,N_1328);
nand U3490 (N_3490,N_2117,N_1223);
nor U3491 (N_3491,N_940,N_1363);
nor U3492 (N_3492,N_490,N_1306);
nand U3493 (N_3493,N_611,N_880);
nand U3494 (N_3494,N_1183,N_755);
or U3495 (N_3495,N_2008,N_1790);
xnor U3496 (N_3496,N_65,N_184);
xnor U3497 (N_3497,N_1524,N_1737);
nand U3498 (N_3498,N_278,N_2496);
nor U3499 (N_3499,N_1194,N_2327);
nor U3500 (N_3500,N_2038,N_660);
and U3501 (N_3501,N_2316,N_700);
xor U3502 (N_3502,N_1462,N_1820);
and U3503 (N_3503,N_1373,N_523);
nor U3504 (N_3504,N_2174,N_2194);
and U3505 (N_3505,N_2196,N_1246);
nor U3506 (N_3506,N_651,N_479);
nor U3507 (N_3507,N_2229,N_234);
or U3508 (N_3508,N_2142,N_1554);
xor U3509 (N_3509,N_458,N_1391);
nand U3510 (N_3510,N_1951,N_1740);
or U3511 (N_3511,N_2192,N_211);
and U3512 (N_3512,N_431,N_2068);
or U3513 (N_3513,N_1126,N_1376);
xnor U3514 (N_3514,N_2471,N_2302);
xnor U3515 (N_3515,N_2051,N_1726);
nor U3516 (N_3516,N_313,N_1427);
nand U3517 (N_3517,N_2214,N_2122);
nor U3518 (N_3518,N_1694,N_1936);
nor U3519 (N_3519,N_2374,N_2110);
or U3520 (N_3520,N_729,N_1300);
nor U3521 (N_3521,N_1917,N_1294);
xor U3522 (N_3522,N_1446,N_1131);
nor U3523 (N_3523,N_14,N_1614);
nand U3524 (N_3524,N_1568,N_496);
nor U3525 (N_3525,N_1063,N_1609);
and U3526 (N_3526,N_511,N_1426);
nor U3527 (N_3527,N_814,N_1492);
xor U3528 (N_3528,N_2386,N_149);
nand U3529 (N_3529,N_322,N_1195);
and U3530 (N_3530,N_2484,N_2012);
nor U3531 (N_3531,N_441,N_488);
or U3532 (N_3532,N_1679,N_974);
nand U3533 (N_3533,N_662,N_388);
nor U3534 (N_3534,N_176,N_267);
xnor U3535 (N_3535,N_1497,N_306);
nor U3536 (N_3536,N_2094,N_955);
nor U3537 (N_3537,N_1610,N_1149);
nand U3538 (N_3538,N_524,N_1434);
or U3539 (N_3539,N_1481,N_391);
or U3540 (N_3540,N_1467,N_269);
or U3541 (N_3541,N_1641,N_237);
and U3542 (N_3542,N_855,N_771);
nand U3543 (N_3543,N_1339,N_453);
xor U3544 (N_3544,N_572,N_1199);
xnor U3545 (N_3545,N_1254,N_1884);
nor U3546 (N_3546,N_1297,N_827);
xnor U3547 (N_3547,N_418,N_839);
and U3548 (N_3548,N_1943,N_520);
or U3549 (N_3549,N_120,N_2297);
nand U3550 (N_3550,N_1508,N_2291);
nand U3551 (N_3551,N_1946,N_1598);
nand U3552 (N_3552,N_1459,N_1673);
xor U3553 (N_3553,N_485,N_642);
nor U3554 (N_3554,N_2282,N_390);
and U3555 (N_3555,N_2426,N_112);
nor U3556 (N_3556,N_1243,N_1172);
nor U3557 (N_3557,N_1384,N_1940);
nor U3558 (N_3558,N_876,N_2159);
nor U3559 (N_3559,N_1708,N_742);
or U3560 (N_3560,N_2118,N_907);
and U3561 (N_3561,N_2136,N_911);
and U3562 (N_3562,N_1660,N_1831);
and U3563 (N_3563,N_2057,N_130);
and U3564 (N_3564,N_1960,N_2303);
or U3565 (N_3565,N_41,N_1221);
nor U3566 (N_3566,N_1719,N_714);
nand U3567 (N_3567,N_2367,N_230);
nor U3568 (N_3568,N_442,N_2218);
nand U3569 (N_3569,N_1636,N_1725);
or U3570 (N_3570,N_249,N_900);
xnor U3571 (N_3571,N_871,N_500);
nor U3572 (N_3572,N_2168,N_858);
and U3573 (N_3573,N_808,N_867);
nor U3574 (N_3574,N_328,N_1032);
xor U3575 (N_3575,N_2,N_378);
xnor U3576 (N_3576,N_1580,N_140);
or U3577 (N_3577,N_1053,N_191);
xor U3578 (N_3578,N_333,N_2335);
and U3579 (N_3579,N_1768,N_137);
and U3580 (N_3580,N_934,N_1181);
or U3581 (N_3581,N_1399,N_1593);
xor U3582 (N_3582,N_1902,N_1883);
and U3583 (N_3583,N_1811,N_1729);
or U3584 (N_3584,N_2130,N_2399);
or U3585 (N_3585,N_1081,N_2494);
nor U3586 (N_3586,N_1709,N_1006);
and U3587 (N_3587,N_1898,N_1180);
or U3588 (N_3588,N_1390,N_1693);
xor U3589 (N_3589,N_1237,N_119);
nand U3590 (N_3590,N_1821,N_2414);
nand U3591 (N_3591,N_1098,N_1888);
xor U3592 (N_3592,N_2052,N_913);
and U3593 (N_3593,N_369,N_1862);
or U3594 (N_3594,N_564,N_2171);
and U3595 (N_3595,N_657,N_2258);
and U3596 (N_3596,N_1417,N_203);
nor U3597 (N_3597,N_2388,N_59);
xnor U3598 (N_3598,N_1142,N_454);
and U3599 (N_3599,N_1617,N_1856);
nand U3600 (N_3600,N_844,N_872);
or U3601 (N_3601,N_968,N_1808);
nand U3602 (N_3602,N_2033,N_873);
and U3603 (N_3603,N_160,N_1954);
and U3604 (N_3604,N_2368,N_212);
nor U3605 (N_3605,N_1330,N_1451);
or U3606 (N_3606,N_885,N_2186);
nor U3607 (N_3607,N_252,N_1922);
xnor U3608 (N_3608,N_516,N_772);
or U3609 (N_3609,N_52,N_2298);
xnor U3610 (N_3610,N_415,N_664);
nor U3611 (N_3611,N_1256,N_299);
or U3612 (N_3612,N_1028,N_1948);
and U3613 (N_3613,N_653,N_151);
and U3614 (N_3614,N_185,N_2451);
or U3615 (N_3615,N_1043,N_1349);
or U3616 (N_3616,N_1469,N_1910);
or U3617 (N_3617,N_1054,N_1289);
and U3618 (N_3618,N_966,N_308);
xor U3619 (N_3619,N_1661,N_295);
nand U3620 (N_3620,N_2445,N_2404);
nor U3621 (N_3621,N_1744,N_1908);
nand U3622 (N_3622,N_456,N_699);
nor U3623 (N_3623,N_1705,N_2491);
nor U3624 (N_3624,N_226,N_915);
and U3625 (N_3625,N_2338,N_1025);
xnor U3626 (N_3626,N_2421,N_301);
nand U3627 (N_3627,N_1643,N_544);
or U3628 (N_3628,N_183,N_786);
xor U3629 (N_3629,N_343,N_335);
nor U3630 (N_3630,N_1957,N_1072);
or U3631 (N_3631,N_248,N_297);
or U3632 (N_3632,N_720,N_1537);
and U3633 (N_3633,N_1850,N_6);
nor U3634 (N_3634,N_1206,N_102);
or U3635 (N_3635,N_605,N_2045);
nor U3636 (N_3636,N_1438,N_2242);
nand U3637 (N_3637,N_1466,N_265);
nand U3638 (N_3638,N_1007,N_2453);
and U3639 (N_3639,N_851,N_2301);
or U3640 (N_3640,N_1017,N_2063);
or U3641 (N_3641,N_1089,N_994);
or U3642 (N_3642,N_148,N_1766);
and U3643 (N_3643,N_2101,N_1901);
nor U3644 (N_3644,N_1124,N_1410);
xor U3645 (N_3645,N_890,N_2166);
nor U3646 (N_3646,N_1904,N_884);
and U3647 (N_3647,N_1477,N_1786);
nand U3648 (N_3648,N_2080,N_438);
nand U3649 (N_3649,N_1073,N_2089);
nor U3650 (N_3650,N_2060,N_2201);
and U3651 (N_3651,N_1354,N_763);
or U3652 (N_3652,N_1471,N_1164);
and U3653 (N_3653,N_2116,N_1967);
xnor U3654 (N_3654,N_1979,N_1505);
or U3655 (N_3655,N_2035,N_1141);
xor U3656 (N_3656,N_988,N_621);
xor U3657 (N_3657,N_495,N_594);
nor U3658 (N_3658,N_1200,N_793);
xnor U3659 (N_3659,N_1086,N_1782);
or U3660 (N_3660,N_2323,N_1518);
nor U3661 (N_3661,N_1989,N_135);
nor U3662 (N_3662,N_201,N_2446);
nand U3663 (N_3663,N_693,N_320);
or U3664 (N_3664,N_996,N_1188);
or U3665 (N_3665,N_1100,N_231);
nor U3666 (N_3666,N_1118,N_679);
xnor U3667 (N_3667,N_2098,N_1396);
or U3668 (N_3668,N_2073,N_1103);
and U3669 (N_3669,N_1564,N_837);
xnor U3670 (N_3670,N_1071,N_620);
xor U3671 (N_3671,N_1250,N_2131);
nor U3672 (N_3672,N_1040,N_792);
nand U3673 (N_3673,N_386,N_567);
and U3674 (N_3674,N_952,N_946);
xnor U3675 (N_3675,N_696,N_643);
xor U3676 (N_3676,N_2154,N_1509);
or U3677 (N_3677,N_2066,N_1058);
and U3678 (N_3678,N_1135,N_1530);
nand U3679 (N_3679,N_1727,N_2149);
and U3680 (N_3680,N_536,N_2378);
nand U3681 (N_3681,N_1620,N_2138);
or U3682 (N_3682,N_239,N_2261);
or U3683 (N_3683,N_1829,N_1690);
nand U3684 (N_3684,N_1023,N_1724);
and U3685 (N_3685,N_67,N_2410);
xor U3686 (N_3686,N_1490,N_1667);
or U3687 (N_3687,N_1669,N_1234);
and U3688 (N_3688,N_503,N_2348);
and U3689 (N_3689,N_759,N_1785);
nor U3690 (N_3690,N_2023,N_2497);
xnor U3691 (N_3691,N_545,N_830);
or U3692 (N_3692,N_1027,N_2460);
and U3693 (N_3693,N_1,N_744);
or U3694 (N_3694,N_2437,N_797);
and U3695 (N_3695,N_1239,N_255);
xnor U3696 (N_3696,N_2257,N_1637);
and U3697 (N_3697,N_324,N_1036);
or U3698 (N_3698,N_1909,N_535);
or U3699 (N_3699,N_1018,N_1876);
and U3700 (N_3700,N_1939,N_2091);
nor U3701 (N_3701,N_1173,N_1627);
and U3702 (N_3702,N_1588,N_863);
nor U3703 (N_3703,N_1147,N_408);
xor U3704 (N_3704,N_1483,N_2178);
nor U3705 (N_3705,N_244,N_2263);
or U3706 (N_3706,N_823,N_2452);
nand U3707 (N_3707,N_526,N_2114);
nand U3708 (N_3708,N_682,N_428);
nand U3709 (N_3709,N_1557,N_1022);
xor U3710 (N_3710,N_1700,N_99);
nand U3711 (N_3711,N_412,N_426);
nand U3712 (N_3712,N_18,N_198);
nor U3713 (N_3713,N_2097,N_1293);
nand U3714 (N_3714,N_951,N_2355);
nand U3715 (N_3715,N_2183,N_910);
nand U3716 (N_3716,N_2013,N_561);
and U3717 (N_3717,N_9,N_1351);
nand U3718 (N_3718,N_1132,N_480);
nor U3719 (N_3719,N_1004,N_1837);
nor U3720 (N_3720,N_1503,N_1003);
nor U3721 (N_3721,N_2358,N_326);
xor U3722 (N_3722,N_846,N_897);
and U3723 (N_3723,N_963,N_1463);
xnor U3724 (N_3724,N_502,N_829);
nor U3725 (N_3725,N_2354,N_92);
xnor U3726 (N_3726,N_247,N_419);
nor U3727 (N_3727,N_1150,N_514);
xnor U3728 (N_3728,N_1586,N_625);
nand U3729 (N_3729,N_1334,N_2468);
and U3730 (N_3730,N_674,N_2204);
xor U3731 (N_3731,N_146,N_1824);
or U3732 (N_3732,N_1722,N_1002);
xnor U3733 (N_3733,N_1978,N_1771);
nand U3734 (N_3734,N_972,N_259);
nand U3735 (N_3735,N_1897,N_888);
nand U3736 (N_3736,N_360,N_2020);
nor U3737 (N_3737,N_1969,N_2436);
and U3738 (N_3738,N_361,N_856);
nand U3739 (N_3739,N_1074,N_2017);
nor U3740 (N_3740,N_455,N_81);
xnor U3741 (N_3741,N_2344,N_1095);
or U3742 (N_3742,N_1955,N_123);
xnor U3743 (N_3743,N_967,N_2010);
or U3744 (N_3744,N_466,N_1165);
or U3745 (N_3745,N_192,N_2375);
and U3746 (N_3746,N_1075,N_2489);
nand U3747 (N_3747,N_1746,N_2230);
and U3748 (N_3748,N_1870,N_300);
xnor U3749 (N_3749,N_358,N_1152);
and U3750 (N_3750,N_82,N_1745);
or U3751 (N_3751,N_2355,N_2025);
nor U3752 (N_3752,N_2092,N_320);
nand U3753 (N_3753,N_427,N_1830);
xnor U3754 (N_3754,N_1320,N_2058);
nor U3755 (N_3755,N_1346,N_1681);
nand U3756 (N_3756,N_2345,N_982);
xor U3757 (N_3757,N_516,N_1470);
nand U3758 (N_3758,N_1940,N_1034);
and U3759 (N_3759,N_1026,N_1097);
or U3760 (N_3760,N_1780,N_1249);
nor U3761 (N_3761,N_763,N_588);
or U3762 (N_3762,N_2297,N_2386);
or U3763 (N_3763,N_1805,N_613);
or U3764 (N_3764,N_741,N_312);
nand U3765 (N_3765,N_2146,N_315);
and U3766 (N_3766,N_965,N_1834);
or U3767 (N_3767,N_1181,N_1532);
and U3768 (N_3768,N_2383,N_860);
or U3769 (N_3769,N_890,N_1935);
and U3770 (N_3770,N_1029,N_180);
xnor U3771 (N_3771,N_2183,N_2408);
or U3772 (N_3772,N_2368,N_272);
xor U3773 (N_3773,N_1938,N_2131);
xnor U3774 (N_3774,N_771,N_568);
nor U3775 (N_3775,N_1917,N_944);
xor U3776 (N_3776,N_1409,N_2116);
nor U3777 (N_3777,N_1842,N_2217);
nand U3778 (N_3778,N_179,N_1531);
or U3779 (N_3779,N_387,N_2436);
xor U3780 (N_3780,N_644,N_1637);
nand U3781 (N_3781,N_1280,N_998);
nor U3782 (N_3782,N_1868,N_2313);
or U3783 (N_3783,N_1016,N_831);
or U3784 (N_3784,N_2254,N_665);
xnor U3785 (N_3785,N_1660,N_544);
or U3786 (N_3786,N_1616,N_1315);
nor U3787 (N_3787,N_1552,N_978);
nand U3788 (N_3788,N_1861,N_851);
nand U3789 (N_3789,N_803,N_1441);
xor U3790 (N_3790,N_236,N_286);
or U3791 (N_3791,N_813,N_1532);
nor U3792 (N_3792,N_2248,N_942);
nor U3793 (N_3793,N_1056,N_1482);
or U3794 (N_3794,N_1793,N_191);
xnor U3795 (N_3795,N_484,N_1661);
nand U3796 (N_3796,N_2352,N_420);
and U3797 (N_3797,N_2298,N_339);
nand U3798 (N_3798,N_78,N_299);
xor U3799 (N_3799,N_606,N_384);
nand U3800 (N_3800,N_85,N_2137);
and U3801 (N_3801,N_580,N_2049);
nor U3802 (N_3802,N_1443,N_1874);
xnor U3803 (N_3803,N_3,N_2356);
xor U3804 (N_3804,N_1496,N_1378);
and U3805 (N_3805,N_1366,N_1623);
or U3806 (N_3806,N_384,N_537);
and U3807 (N_3807,N_520,N_2476);
xnor U3808 (N_3808,N_109,N_1211);
nand U3809 (N_3809,N_510,N_484);
nand U3810 (N_3810,N_852,N_895);
or U3811 (N_3811,N_1748,N_1007);
nor U3812 (N_3812,N_70,N_2155);
or U3813 (N_3813,N_1537,N_1397);
and U3814 (N_3814,N_568,N_669);
or U3815 (N_3815,N_1639,N_1984);
nor U3816 (N_3816,N_467,N_830);
xnor U3817 (N_3817,N_1388,N_2097);
nor U3818 (N_3818,N_2256,N_505);
nor U3819 (N_3819,N_1309,N_574);
or U3820 (N_3820,N_2186,N_711);
nand U3821 (N_3821,N_2471,N_2072);
and U3822 (N_3822,N_1923,N_1125);
and U3823 (N_3823,N_1061,N_970);
nor U3824 (N_3824,N_68,N_1943);
nor U3825 (N_3825,N_1851,N_1873);
and U3826 (N_3826,N_1867,N_2350);
nand U3827 (N_3827,N_2392,N_249);
nand U3828 (N_3828,N_1404,N_604);
or U3829 (N_3829,N_2195,N_1983);
nor U3830 (N_3830,N_1635,N_1632);
xor U3831 (N_3831,N_2267,N_2350);
nor U3832 (N_3832,N_2064,N_2153);
xor U3833 (N_3833,N_167,N_1163);
xnor U3834 (N_3834,N_1210,N_7);
nand U3835 (N_3835,N_161,N_1353);
xnor U3836 (N_3836,N_747,N_616);
nand U3837 (N_3837,N_810,N_1167);
nor U3838 (N_3838,N_749,N_1704);
xor U3839 (N_3839,N_2377,N_2496);
nand U3840 (N_3840,N_433,N_600);
xor U3841 (N_3841,N_552,N_272);
or U3842 (N_3842,N_1435,N_1230);
or U3843 (N_3843,N_1248,N_2472);
nand U3844 (N_3844,N_927,N_1767);
nand U3845 (N_3845,N_1162,N_1858);
and U3846 (N_3846,N_45,N_2117);
xor U3847 (N_3847,N_925,N_1128);
nor U3848 (N_3848,N_58,N_519);
nor U3849 (N_3849,N_1554,N_622);
xnor U3850 (N_3850,N_858,N_999);
nor U3851 (N_3851,N_709,N_1757);
nand U3852 (N_3852,N_895,N_1451);
xor U3853 (N_3853,N_1977,N_609);
and U3854 (N_3854,N_1435,N_2139);
and U3855 (N_3855,N_2214,N_1515);
nand U3856 (N_3856,N_2136,N_868);
or U3857 (N_3857,N_2163,N_721);
xor U3858 (N_3858,N_2464,N_455);
or U3859 (N_3859,N_1715,N_2172);
xor U3860 (N_3860,N_1378,N_1484);
xor U3861 (N_3861,N_1604,N_896);
nor U3862 (N_3862,N_653,N_2405);
nand U3863 (N_3863,N_1568,N_2402);
xnor U3864 (N_3864,N_514,N_1381);
xor U3865 (N_3865,N_1328,N_697);
nand U3866 (N_3866,N_2141,N_2420);
and U3867 (N_3867,N_190,N_2270);
xor U3868 (N_3868,N_899,N_575);
or U3869 (N_3869,N_229,N_387);
nand U3870 (N_3870,N_890,N_7);
xor U3871 (N_3871,N_1541,N_724);
xor U3872 (N_3872,N_1793,N_749);
and U3873 (N_3873,N_1752,N_832);
xnor U3874 (N_3874,N_670,N_1202);
xor U3875 (N_3875,N_2113,N_871);
or U3876 (N_3876,N_1850,N_2408);
nand U3877 (N_3877,N_978,N_1322);
and U3878 (N_3878,N_1019,N_1052);
and U3879 (N_3879,N_2438,N_2046);
nand U3880 (N_3880,N_1827,N_845);
or U3881 (N_3881,N_2498,N_1854);
and U3882 (N_3882,N_2437,N_1801);
or U3883 (N_3883,N_482,N_1319);
or U3884 (N_3884,N_995,N_654);
nand U3885 (N_3885,N_2455,N_97);
and U3886 (N_3886,N_2089,N_2423);
and U3887 (N_3887,N_123,N_1948);
or U3888 (N_3888,N_2236,N_415);
and U3889 (N_3889,N_962,N_1601);
nor U3890 (N_3890,N_232,N_1146);
nor U3891 (N_3891,N_520,N_259);
xor U3892 (N_3892,N_2274,N_1294);
nand U3893 (N_3893,N_1283,N_414);
nor U3894 (N_3894,N_1495,N_947);
nand U3895 (N_3895,N_1754,N_1432);
xor U3896 (N_3896,N_2389,N_996);
and U3897 (N_3897,N_2004,N_262);
or U3898 (N_3898,N_2012,N_2279);
xor U3899 (N_3899,N_1723,N_1052);
nor U3900 (N_3900,N_654,N_2326);
and U3901 (N_3901,N_1764,N_1224);
or U3902 (N_3902,N_513,N_804);
nand U3903 (N_3903,N_2038,N_2466);
xnor U3904 (N_3904,N_2329,N_948);
nor U3905 (N_3905,N_877,N_769);
and U3906 (N_3906,N_1021,N_396);
xor U3907 (N_3907,N_1950,N_1004);
nor U3908 (N_3908,N_1726,N_2231);
or U3909 (N_3909,N_1072,N_1749);
and U3910 (N_3910,N_305,N_2489);
nand U3911 (N_3911,N_110,N_437);
xor U3912 (N_3912,N_1943,N_1325);
xnor U3913 (N_3913,N_336,N_498);
xnor U3914 (N_3914,N_2228,N_1326);
xor U3915 (N_3915,N_1361,N_786);
nand U3916 (N_3916,N_1686,N_1439);
nor U3917 (N_3917,N_2079,N_1637);
xnor U3918 (N_3918,N_1248,N_329);
xnor U3919 (N_3919,N_5,N_1245);
and U3920 (N_3920,N_2411,N_2434);
nor U3921 (N_3921,N_1331,N_919);
nor U3922 (N_3922,N_1600,N_894);
nor U3923 (N_3923,N_781,N_1164);
xnor U3924 (N_3924,N_874,N_2102);
or U3925 (N_3925,N_691,N_1826);
nand U3926 (N_3926,N_2490,N_127);
nand U3927 (N_3927,N_1252,N_2131);
and U3928 (N_3928,N_868,N_1519);
nand U3929 (N_3929,N_1791,N_1097);
xnor U3930 (N_3930,N_147,N_1678);
nand U3931 (N_3931,N_234,N_745);
nor U3932 (N_3932,N_418,N_176);
xor U3933 (N_3933,N_2325,N_1133);
nand U3934 (N_3934,N_183,N_1948);
and U3935 (N_3935,N_884,N_2134);
nand U3936 (N_3936,N_1730,N_783);
nor U3937 (N_3937,N_2169,N_212);
or U3938 (N_3938,N_1208,N_261);
nor U3939 (N_3939,N_1932,N_1625);
nor U3940 (N_3940,N_1036,N_4);
nand U3941 (N_3941,N_891,N_1187);
nand U3942 (N_3942,N_2025,N_1354);
xor U3943 (N_3943,N_1551,N_151);
or U3944 (N_3944,N_1109,N_1877);
and U3945 (N_3945,N_1834,N_2406);
or U3946 (N_3946,N_1621,N_1501);
nor U3947 (N_3947,N_1634,N_2017);
nand U3948 (N_3948,N_446,N_883);
nand U3949 (N_3949,N_1642,N_1802);
and U3950 (N_3950,N_498,N_2485);
xnor U3951 (N_3951,N_887,N_1703);
nand U3952 (N_3952,N_2332,N_309);
and U3953 (N_3953,N_72,N_646);
xor U3954 (N_3954,N_2492,N_541);
nand U3955 (N_3955,N_2073,N_1683);
or U3956 (N_3956,N_335,N_905);
or U3957 (N_3957,N_373,N_636);
xnor U3958 (N_3958,N_902,N_767);
xnor U3959 (N_3959,N_79,N_884);
nand U3960 (N_3960,N_1630,N_1450);
nand U3961 (N_3961,N_598,N_975);
nor U3962 (N_3962,N_224,N_2165);
xor U3963 (N_3963,N_459,N_2234);
or U3964 (N_3964,N_1553,N_845);
xnor U3965 (N_3965,N_1534,N_1810);
xnor U3966 (N_3966,N_1952,N_2368);
or U3967 (N_3967,N_2085,N_531);
nand U3968 (N_3968,N_1337,N_952);
nor U3969 (N_3969,N_2283,N_1634);
nor U3970 (N_3970,N_408,N_692);
and U3971 (N_3971,N_2362,N_1845);
nand U3972 (N_3972,N_1220,N_415);
or U3973 (N_3973,N_2026,N_433);
nand U3974 (N_3974,N_2211,N_1677);
and U3975 (N_3975,N_1829,N_1647);
and U3976 (N_3976,N_2142,N_961);
and U3977 (N_3977,N_1782,N_745);
or U3978 (N_3978,N_533,N_1012);
xnor U3979 (N_3979,N_2115,N_1662);
and U3980 (N_3980,N_1380,N_732);
nor U3981 (N_3981,N_663,N_976);
xnor U3982 (N_3982,N_930,N_1997);
and U3983 (N_3983,N_968,N_2014);
nand U3984 (N_3984,N_1332,N_2234);
and U3985 (N_3985,N_2285,N_2218);
nor U3986 (N_3986,N_177,N_1578);
nand U3987 (N_3987,N_1002,N_1334);
or U3988 (N_3988,N_207,N_928);
and U3989 (N_3989,N_108,N_899);
nand U3990 (N_3990,N_1042,N_1493);
and U3991 (N_3991,N_2259,N_1601);
and U3992 (N_3992,N_2187,N_2190);
or U3993 (N_3993,N_2094,N_1808);
nor U3994 (N_3994,N_583,N_613);
or U3995 (N_3995,N_645,N_1982);
or U3996 (N_3996,N_108,N_2222);
xor U3997 (N_3997,N_2215,N_1754);
xor U3998 (N_3998,N_1633,N_1268);
or U3999 (N_3999,N_1322,N_239);
or U4000 (N_4000,N_728,N_2402);
or U4001 (N_4001,N_1906,N_175);
xor U4002 (N_4002,N_2298,N_2109);
nor U4003 (N_4003,N_2358,N_370);
nor U4004 (N_4004,N_2248,N_2404);
xor U4005 (N_4005,N_399,N_1729);
xor U4006 (N_4006,N_2058,N_395);
nor U4007 (N_4007,N_1674,N_2376);
or U4008 (N_4008,N_1150,N_532);
or U4009 (N_4009,N_398,N_1373);
nor U4010 (N_4010,N_2494,N_2240);
and U4011 (N_4011,N_1692,N_1690);
nand U4012 (N_4012,N_567,N_2312);
and U4013 (N_4013,N_2329,N_922);
nor U4014 (N_4014,N_1809,N_1200);
and U4015 (N_4015,N_1104,N_1525);
nand U4016 (N_4016,N_1529,N_1317);
or U4017 (N_4017,N_1251,N_1774);
nand U4018 (N_4018,N_2097,N_1214);
nor U4019 (N_4019,N_417,N_1748);
xnor U4020 (N_4020,N_459,N_1614);
nand U4021 (N_4021,N_2355,N_1000);
nand U4022 (N_4022,N_1371,N_2072);
xor U4023 (N_4023,N_1115,N_1221);
nor U4024 (N_4024,N_1632,N_856);
nor U4025 (N_4025,N_907,N_961);
nand U4026 (N_4026,N_1735,N_1284);
nor U4027 (N_4027,N_102,N_2291);
or U4028 (N_4028,N_1747,N_1620);
nor U4029 (N_4029,N_2400,N_463);
xor U4030 (N_4030,N_1792,N_2134);
xnor U4031 (N_4031,N_428,N_239);
and U4032 (N_4032,N_1127,N_508);
and U4033 (N_4033,N_690,N_1654);
nand U4034 (N_4034,N_2308,N_1959);
and U4035 (N_4035,N_297,N_1890);
nor U4036 (N_4036,N_1507,N_1615);
or U4037 (N_4037,N_2246,N_2408);
nor U4038 (N_4038,N_2050,N_1862);
xnor U4039 (N_4039,N_2380,N_76);
nor U4040 (N_4040,N_2113,N_256);
or U4041 (N_4041,N_888,N_2268);
and U4042 (N_4042,N_1435,N_709);
and U4043 (N_4043,N_663,N_147);
or U4044 (N_4044,N_777,N_1407);
nand U4045 (N_4045,N_1778,N_68);
nor U4046 (N_4046,N_1433,N_1478);
or U4047 (N_4047,N_1965,N_1605);
xnor U4048 (N_4048,N_2180,N_1591);
or U4049 (N_4049,N_526,N_830);
nand U4050 (N_4050,N_513,N_1593);
nand U4051 (N_4051,N_1017,N_1639);
xor U4052 (N_4052,N_869,N_2297);
xor U4053 (N_4053,N_642,N_257);
xnor U4054 (N_4054,N_445,N_528);
or U4055 (N_4055,N_2052,N_1190);
xnor U4056 (N_4056,N_1478,N_1818);
xnor U4057 (N_4057,N_2291,N_2385);
and U4058 (N_4058,N_42,N_572);
or U4059 (N_4059,N_1580,N_561);
xnor U4060 (N_4060,N_1788,N_139);
nand U4061 (N_4061,N_2360,N_644);
nand U4062 (N_4062,N_2320,N_2330);
nand U4063 (N_4063,N_527,N_1545);
nand U4064 (N_4064,N_789,N_1786);
nand U4065 (N_4065,N_917,N_1167);
and U4066 (N_4066,N_946,N_331);
nor U4067 (N_4067,N_312,N_1438);
nand U4068 (N_4068,N_1786,N_2072);
or U4069 (N_4069,N_39,N_316);
nor U4070 (N_4070,N_2294,N_1793);
and U4071 (N_4071,N_1416,N_204);
xor U4072 (N_4072,N_2489,N_1278);
or U4073 (N_4073,N_1771,N_1387);
xor U4074 (N_4074,N_1923,N_850);
nand U4075 (N_4075,N_818,N_972);
or U4076 (N_4076,N_152,N_1919);
nor U4077 (N_4077,N_402,N_702);
or U4078 (N_4078,N_80,N_326);
nand U4079 (N_4079,N_1823,N_831);
xnor U4080 (N_4080,N_2455,N_910);
and U4081 (N_4081,N_1142,N_135);
or U4082 (N_4082,N_2336,N_1510);
and U4083 (N_4083,N_77,N_1996);
xnor U4084 (N_4084,N_1154,N_1029);
and U4085 (N_4085,N_2448,N_1457);
or U4086 (N_4086,N_481,N_2282);
nand U4087 (N_4087,N_1024,N_492);
or U4088 (N_4088,N_2369,N_2460);
or U4089 (N_4089,N_1792,N_633);
nor U4090 (N_4090,N_1175,N_1447);
or U4091 (N_4091,N_694,N_121);
xor U4092 (N_4092,N_1589,N_975);
or U4093 (N_4093,N_476,N_2147);
nand U4094 (N_4094,N_463,N_2112);
or U4095 (N_4095,N_323,N_2025);
or U4096 (N_4096,N_421,N_1802);
nor U4097 (N_4097,N_1641,N_72);
or U4098 (N_4098,N_890,N_1334);
xnor U4099 (N_4099,N_2409,N_1743);
nand U4100 (N_4100,N_2271,N_2301);
nand U4101 (N_4101,N_449,N_1302);
and U4102 (N_4102,N_2392,N_1971);
and U4103 (N_4103,N_203,N_2047);
nand U4104 (N_4104,N_1734,N_2423);
or U4105 (N_4105,N_1613,N_1741);
and U4106 (N_4106,N_2034,N_725);
nor U4107 (N_4107,N_598,N_372);
and U4108 (N_4108,N_1610,N_2294);
xor U4109 (N_4109,N_618,N_168);
nor U4110 (N_4110,N_2274,N_2069);
or U4111 (N_4111,N_1679,N_2205);
or U4112 (N_4112,N_1591,N_457);
and U4113 (N_4113,N_385,N_1637);
nand U4114 (N_4114,N_401,N_1924);
nand U4115 (N_4115,N_45,N_1613);
and U4116 (N_4116,N_104,N_724);
nor U4117 (N_4117,N_2128,N_2332);
nand U4118 (N_4118,N_1463,N_157);
or U4119 (N_4119,N_391,N_1202);
xor U4120 (N_4120,N_2205,N_1844);
and U4121 (N_4121,N_1608,N_837);
xnor U4122 (N_4122,N_283,N_210);
xor U4123 (N_4123,N_1532,N_2312);
nor U4124 (N_4124,N_853,N_1617);
nor U4125 (N_4125,N_767,N_270);
nor U4126 (N_4126,N_1955,N_1422);
and U4127 (N_4127,N_1377,N_1871);
xor U4128 (N_4128,N_2109,N_938);
xnor U4129 (N_4129,N_1852,N_768);
xnor U4130 (N_4130,N_738,N_2198);
or U4131 (N_4131,N_2268,N_2174);
or U4132 (N_4132,N_2031,N_1633);
nor U4133 (N_4133,N_676,N_337);
and U4134 (N_4134,N_1582,N_822);
and U4135 (N_4135,N_1130,N_1534);
nand U4136 (N_4136,N_2068,N_2367);
nand U4137 (N_4137,N_638,N_2084);
nand U4138 (N_4138,N_1108,N_853);
xor U4139 (N_4139,N_730,N_1958);
or U4140 (N_4140,N_1189,N_2391);
or U4141 (N_4141,N_2096,N_58);
nand U4142 (N_4142,N_93,N_2128);
nand U4143 (N_4143,N_197,N_826);
or U4144 (N_4144,N_1676,N_683);
or U4145 (N_4145,N_1809,N_2009);
or U4146 (N_4146,N_2310,N_404);
nand U4147 (N_4147,N_2400,N_2173);
nor U4148 (N_4148,N_1769,N_814);
and U4149 (N_4149,N_1812,N_33);
and U4150 (N_4150,N_336,N_846);
or U4151 (N_4151,N_1766,N_15);
nor U4152 (N_4152,N_1192,N_231);
xnor U4153 (N_4153,N_2271,N_980);
nand U4154 (N_4154,N_443,N_1076);
or U4155 (N_4155,N_389,N_1160);
nor U4156 (N_4156,N_1015,N_2029);
and U4157 (N_4157,N_215,N_2156);
xnor U4158 (N_4158,N_333,N_2394);
nand U4159 (N_4159,N_791,N_2231);
nor U4160 (N_4160,N_885,N_1234);
or U4161 (N_4161,N_1833,N_1905);
nand U4162 (N_4162,N_1694,N_1956);
nand U4163 (N_4163,N_2011,N_2277);
and U4164 (N_4164,N_1369,N_846);
xor U4165 (N_4165,N_1670,N_812);
nand U4166 (N_4166,N_321,N_644);
nand U4167 (N_4167,N_1181,N_408);
xnor U4168 (N_4168,N_1764,N_504);
nor U4169 (N_4169,N_665,N_1348);
nor U4170 (N_4170,N_968,N_1726);
and U4171 (N_4171,N_1756,N_2479);
and U4172 (N_4172,N_2388,N_1342);
nor U4173 (N_4173,N_1257,N_2480);
or U4174 (N_4174,N_1637,N_1638);
and U4175 (N_4175,N_1843,N_2178);
and U4176 (N_4176,N_2490,N_38);
nor U4177 (N_4177,N_436,N_1713);
xor U4178 (N_4178,N_2177,N_1127);
and U4179 (N_4179,N_1797,N_840);
and U4180 (N_4180,N_773,N_1383);
nor U4181 (N_4181,N_554,N_669);
nand U4182 (N_4182,N_66,N_1312);
or U4183 (N_4183,N_2209,N_15);
nand U4184 (N_4184,N_1296,N_625);
and U4185 (N_4185,N_1454,N_1666);
or U4186 (N_4186,N_1702,N_1374);
nor U4187 (N_4187,N_1288,N_43);
or U4188 (N_4188,N_1312,N_2169);
or U4189 (N_4189,N_1977,N_461);
nor U4190 (N_4190,N_1371,N_218);
and U4191 (N_4191,N_2162,N_2180);
and U4192 (N_4192,N_383,N_960);
nand U4193 (N_4193,N_1901,N_1852);
nand U4194 (N_4194,N_2136,N_407);
and U4195 (N_4195,N_1875,N_1719);
nand U4196 (N_4196,N_59,N_1942);
xor U4197 (N_4197,N_865,N_575);
and U4198 (N_4198,N_1942,N_601);
xnor U4199 (N_4199,N_1925,N_392);
nand U4200 (N_4200,N_1247,N_2412);
and U4201 (N_4201,N_1173,N_1354);
nand U4202 (N_4202,N_578,N_1135);
xnor U4203 (N_4203,N_1238,N_2242);
nor U4204 (N_4204,N_1229,N_1473);
nor U4205 (N_4205,N_376,N_66);
and U4206 (N_4206,N_2493,N_2075);
nor U4207 (N_4207,N_1362,N_412);
and U4208 (N_4208,N_1484,N_1373);
and U4209 (N_4209,N_193,N_2311);
and U4210 (N_4210,N_2091,N_217);
nor U4211 (N_4211,N_1925,N_76);
xnor U4212 (N_4212,N_1952,N_47);
nor U4213 (N_4213,N_1268,N_2222);
xor U4214 (N_4214,N_2200,N_1340);
nor U4215 (N_4215,N_2236,N_2379);
xor U4216 (N_4216,N_226,N_1252);
and U4217 (N_4217,N_1130,N_722);
nor U4218 (N_4218,N_2184,N_1475);
or U4219 (N_4219,N_625,N_1819);
or U4220 (N_4220,N_192,N_1764);
xor U4221 (N_4221,N_1617,N_1964);
nor U4222 (N_4222,N_1742,N_1453);
nor U4223 (N_4223,N_54,N_1962);
and U4224 (N_4224,N_1589,N_897);
xnor U4225 (N_4225,N_992,N_756);
xnor U4226 (N_4226,N_86,N_2000);
xnor U4227 (N_4227,N_261,N_1417);
nand U4228 (N_4228,N_1279,N_1754);
xnor U4229 (N_4229,N_560,N_19);
xor U4230 (N_4230,N_1276,N_1153);
and U4231 (N_4231,N_1401,N_2402);
or U4232 (N_4232,N_1893,N_1164);
and U4233 (N_4233,N_503,N_1256);
nand U4234 (N_4234,N_2472,N_847);
or U4235 (N_4235,N_1744,N_2444);
or U4236 (N_4236,N_1999,N_1615);
nand U4237 (N_4237,N_1439,N_617);
nor U4238 (N_4238,N_1015,N_1617);
xor U4239 (N_4239,N_56,N_349);
xnor U4240 (N_4240,N_819,N_1729);
nand U4241 (N_4241,N_515,N_581);
xnor U4242 (N_4242,N_2258,N_1604);
nand U4243 (N_4243,N_1065,N_1330);
or U4244 (N_4244,N_733,N_989);
nor U4245 (N_4245,N_493,N_1162);
or U4246 (N_4246,N_341,N_168);
xor U4247 (N_4247,N_1208,N_1321);
and U4248 (N_4248,N_1654,N_1924);
nand U4249 (N_4249,N_944,N_985);
xnor U4250 (N_4250,N_1227,N_36);
nand U4251 (N_4251,N_1522,N_1061);
nand U4252 (N_4252,N_474,N_2101);
or U4253 (N_4253,N_707,N_2078);
nand U4254 (N_4254,N_409,N_1181);
nor U4255 (N_4255,N_10,N_658);
nand U4256 (N_4256,N_2098,N_733);
xor U4257 (N_4257,N_2161,N_2110);
or U4258 (N_4258,N_2129,N_675);
nor U4259 (N_4259,N_186,N_1778);
or U4260 (N_4260,N_621,N_64);
or U4261 (N_4261,N_1475,N_2497);
and U4262 (N_4262,N_101,N_1414);
or U4263 (N_4263,N_252,N_489);
or U4264 (N_4264,N_1664,N_2372);
or U4265 (N_4265,N_1743,N_1280);
nor U4266 (N_4266,N_990,N_1042);
nor U4267 (N_4267,N_2113,N_522);
xor U4268 (N_4268,N_396,N_926);
nand U4269 (N_4269,N_476,N_576);
nor U4270 (N_4270,N_2074,N_42);
nand U4271 (N_4271,N_1012,N_1041);
nor U4272 (N_4272,N_61,N_1424);
nor U4273 (N_4273,N_2169,N_2);
nor U4274 (N_4274,N_1951,N_527);
xnor U4275 (N_4275,N_101,N_1469);
xor U4276 (N_4276,N_471,N_1325);
xnor U4277 (N_4277,N_207,N_2412);
and U4278 (N_4278,N_2164,N_1960);
nor U4279 (N_4279,N_636,N_324);
nand U4280 (N_4280,N_1025,N_735);
and U4281 (N_4281,N_2459,N_260);
nor U4282 (N_4282,N_965,N_724);
and U4283 (N_4283,N_1223,N_452);
nand U4284 (N_4284,N_179,N_127);
and U4285 (N_4285,N_350,N_1298);
xnor U4286 (N_4286,N_2171,N_1336);
xnor U4287 (N_4287,N_1213,N_1450);
nand U4288 (N_4288,N_299,N_1624);
or U4289 (N_4289,N_975,N_97);
xor U4290 (N_4290,N_2350,N_2059);
nor U4291 (N_4291,N_1322,N_2426);
nor U4292 (N_4292,N_1175,N_2093);
nor U4293 (N_4293,N_59,N_1448);
nand U4294 (N_4294,N_1225,N_1961);
or U4295 (N_4295,N_1400,N_885);
xnor U4296 (N_4296,N_1848,N_404);
or U4297 (N_4297,N_119,N_1818);
or U4298 (N_4298,N_927,N_270);
or U4299 (N_4299,N_1928,N_406);
nand U4300 (N_4300,N_1671,N_27);
or U4301 (N_4301,N_981,N_389);
nand U4302 (N_4302,N_2027,N_87);
xnor U4303 (N_4303,N_762,N_2428);
xor U4304 (N_4304,N_210,N_2318);
nand U4305 (N_4305,N_200,N_495);
xnor U4306 (N_4306,N_561,N_858);
nor U4307 (N_4307,N_474,N_2122);
nor U4308 (N_4308,N_1290,N_900);
and U4309 (N_4309,N_54,N_1015);
nand U4310 (N_4310,N_2460,N_2420);
and U4311 (N_4311,N_901,N_1695);
and U4312 (N_4312,N_1430,N_168);
xor U4313 (N_4313,N_2132,N_1456);
or U4314 (N_4314,N_2026,N_41);
xor U4315 (N_4315,N_1445,N_2262);
xor U4316 (N_4316,N_832,N_258);
xnor U4317 (N_4317,N_499,N_105);
nand U4318 (N_4318,N_255,N_511);
nand U4319 (N_4319,N_922,N_691);
xnor U4320 (N_4320,N_2325,N_985);
nand U4321 (N_4321,N_1540,N_9);
and U4322 (N_4322,N_2155,N_150);
or U4323 (N_4323,N_2328,N_820);
nand U4324 (N_4324,N_1781,N_157);
nand U4325 (N_4325,N_45,N_1316);
or U4326 (N_4326,N_520,N_1609);
nand U4327 (N_4327,N_928,N_758);
and U4328 (N_4328,N_489,N_591);
nor U4329 (N_4329,N_1583,N_1636);
and U4330 (N_4330,N_511,N_2237);
nand U4331 (N_4331,N_258,N_2089);
nor U4332 (N_4332,N_2241,N_1403);
and U4333 (N_4333,N_2219,N_2442);
xor U4334 (N_4334,N_1110,N_236);
nand U4335 (N_4335,N_1408,N_1495);
nand U4336 (N_4336,N_1499,N_603);
xor U4337 (N_4337,N_871,N_1574);
and U4338 (N_4338,N_188,N_1760);
nor U4339 (N_4339,N_359,N_356);
or U4340 (N_4340,N_979,N_1342);
and U4341 (N_4341,N_647,N_441);
or U4342 (N_4342,N_1467,N_225);
nor U4343 (N_4343,N_2057,N_2272);
nand U4344 (N_4344,N_1485,N_1843);
nand U4345 (N_4345,N_850,N_630);
and U4346 (N_4346,N_1242,N_342);
and U4347 (N_4347,N_2361,N_1805);
nor U4348 (N_4348,N_1208,N_1461);
or U4349 (N_4349,N_1768,N_1787);
or U4350 (N_4350,N_1635,N_2274);
and U4351 (N_4351,N_143,N_51);
nor U4352 (N_4352,N_1012,N_979);
and U4353 (N_4353,N_1028,N_1848);
or U4354 (N_4354,N_1320,N_387);
nand U4355 (N_4355,N_2049,N_608);
nor U4356 (N_4356,N_1007,N_1658);
and U4357 (N_4357,N_474,N_1238);
or U4358 (N_4358,N_410,N_1811);
nor U4359 (N_4359,N_488,N_314);
and U4360 (N_4360,N_1981,N_2016);
nor U4361 (N_4361,N_918,N_1391);
xnor U4362 (N_4362,N_1214,N_1564);
xnor U4363 (N_4363,N_2086,N_2129);
nand U4364 (N_4364,N_1725,N_1401);
nand U4365 (N_4365,N_846,N_1020);
xor U4366 (N_4366,N_1117,N_472);
nor U4367 (N_4367,N_1535,N_113);
or U4368 (N_4368,N_1840,N_1924);
xnor U4369 (N_4369,N_1035,N_148);
xnor U4370 (N_4370,N_1735,N_2449);
and U4371 (N_4371,N_1059,N_1023);
nand U4372 (N_4372,N_1273,N_1189);
and U4373 (N_4373,N_795,N_970);
or U4374 (N_4374,N_232,N_2220);
and U4375 (N_4375,N_1769,N_262);
and U4376 (N_4376,N_1035,N_2067);
nor U4377 (N_4377,N_2317,N_1564);
or U4378 (N_4378,N_2383,N_1071);
and U4379 (N_4379,N_929,N_1342);
nor U4380 (N_4380,N_1060,N_2238);
nand U4381 (N_4381,N_1607,N_1975);
and U4382 (N_4382,N_37,N_1614);
nand U4383 (N_4383,N_2291,N_962);
xor U4384 (N_4384,N_1185,N_1238);
nor U4385 (N_4385,N_1727,N_2489);
and U4386 (N_4386,N_2492,N_2222);
nor U4387 (N_4387,N_1589,N_2049);
xnor U4388 (N_4388,N_1113,N_1769);
nor U4389 (N_4389,N_736,N_681);
nand U4390 (N_4390,N_809,N_634);
nor U4391 (N_4391,N_1217,N_345);
xnor U4392 (N_4392,N_2426,N_998);
or U4393 (N_4393,N_1966,N_122);
and U4394 (N_4394,N_1517,N_2445);
xor U4395 (N_4395,N_2335,N_2402);
nor U4396 (N_4396,N_1669,N_895);
or U4397 (N_4397,N_2458,N_997);
and U4398 (N_4398,N_21,N_892);
or U4399 (N_4399,N_2478,N_1303);
nor U4400 (N_4400,N_1352,N_1014);
xnor U4401 (N_4401,N_2360,N_2175);
and U4402 (N_4402,N_189,N_143);
xor U4403 (N_4403,N_499,N_612);
or U4404 (N_4404,N_629,N_2012);
xor U4405 (N_4405,N_736,N_402);
or U4406 (N_4406,N_2195,N_589);
nor U4407 (N_4407,N_499,N_2149);
nor U4408 (N_4408,N_1742,N_1085);
and U4409 (N_4409,N_1068,N_2210);
nand U4410 (N_4410,N_2061,N_201);
nor U4411 (N_4411,N_565,N_597);
nand U4412 (N_4412,N_1245,N_1894);
xnor U4413 (N_4413,N_2133,N_1338);
and U4414 (N_4414,N_550,N_1061);
and U4415 (N_4415,N_2281,N_2341);
xnor U4416 (N_4416,N_496,N_779);
nand U4417 (N_4417,N_2257,N_1234);
or U4418 (N_4418,N_1859,N_2125);
xor U4419 (N_4419,N_2343,N_967);
xor U4420 (N_4420,N_1937,N_580);
xnor U4421 (N_4421,N_2066,N_1610);
and U4422 (N_4422,N_1527,N_2082);
or U4423 (N_4423,N_743,N_659);
and U4424 (N_4424,N_1353,N_1905);
xnor U4425 (N_4425,N_448,N_1669);
nand U4426 (N_4426,N_1880,N_115);
nand U4427 (N_4427,N_1598,N_833);
and U4428 (N_4428,N_819,N_1938);
xor U4429 (N_4429,N_529,N_298);
xnor U4430 (N_4430,N_138,N_142);
nor U4431 (N_4431,N_1394,N_2385);
xor U4432 (N_4432,N_1244,N_1298);
nor U4433 (N_4433,N_993,N_367);
or U4434 (N_4434,N_836,N_1685);
nand U4435 (N_4435,N_2260,N_519);
xnor U4436 (N_4436,N_829,N_313);
or U4437 (N_4437,N_2036,N_2292);
nand U4438 (N_4438,N_294,N_2235);
and U4439 (N_4439,N_1788,N_738);
or U4440 (N_4440,N_1215,N_1481);
or U4441 (N_4441,N_1693,N_1926);
nand U4442 (N_4442,N_2085,N_986);
xnor U4443 (N_4443,N_1639,N_2408);
xnor U4444 (N_4444,N_2222,N_640);
and U4445 (N_4445,N_11,N_445);
xnor U4446 (N_4446,N_2054,N_858);
nor U4447 (N_4447,N_1608,N_1182);
nor U4448 (N_4448,N_1513,N_1179);
and U4449 (N_4449,N_395,N_919);
nor U4450 (N_4450,N_1502,N_453);
xnor U4451 (N_4451,N_143,N_520);
nor U4452 (N_4452,N_2032,N_151);
xnor U4453 (N_4453,N_2084,N_1177);
and U4454 (N_4454,N_2246,N_1598);
and U4455 (N_4455,N_2176,N_1012);
or U4456 (N_4456,N_2241,N_1149);
nor U4457 (N_4457,N_339,N_111);
and U4458 (N_4458,N_2011,N_3);
xor U4459 (N_4459,N_2364,N_904);
or U4460 (N_4460,N_267,N_1375);
or U4461 (N_4461,N_1825,N_670);
nor U4462 (N_4462,N_169,N_7);
xor U4463 (N_4463,N_2246,N_553);
nor U4464 (N_4464,N_2219,N_762);
nor U4465 (N_4465,N_1263,N_1166);
and U4466 (N_4466,N_514,N_2006);
or U4467 (N_4467,N_602,N_1600);
nand U4468 (N_4468,N_2432,N_2101);
or U4469 (N_4469,N_1264,N_1759);
xnor U4470 (N_4470,N_980,N_1973);
or U4471 (N_4471,N_1466,N_1821);
and U4472 (N_4472,N_2073,N_418);
and U4473 (N_4473,N_2231,N_941);
and U4474 (N_4474,N_465,N_37);
xnor U4475 (N_4475,N_2434,N_1758);
or U4476 (N_4476,N_1765,N_775);
or U4477 (N_4477,N_2293,N_2422);
nand U4478 (N_4478,N_2499,N_2204);
xnor U4479 (N_4479,N_1078,N_1224);
or U4480 (N_4480,N_402,N_2076);
or U4481 (N_4481,N_1401,N_205);
or U4482 (N_4482,N_1649,N_1531);
or U4483 (N_4483,N_60,N_2292);
or U4484 (N_4484,N_2076,N_525);
xor U4485 (N_4485,N_542,N_346);
and U4486 (N_4486,N_1234,N_236);
or U4487 (N_4487,N_144,N_997);
nor U4488 (N_4488,N_133,N_2346);
and U4489 (N_4489,N_1394,N_1711);
or U4490 (N_4490,N_1251,N_129);
or U4491 (N_4491,N_1392,N_2468);
nand U4492 (N_4492,N_240,N_2187);
nand U4493 (N_4493,N_2096,N_2244);
xnor U4494 (N_4494,N_1572,N_63);
or U4495 (N_4495,N_1067,N_66);
and U4496 (N_4496,N_313,N_1563);
nand U4497 (N_4497,N_2127,N_2278);
nand U4498 (N_4498,N_201,N_2407);
and U4499 (N_4499,N_2283,N_993);
nand U4500 (N_4500,N_1322,N_1185);
nor U4501 (N_4501,N_424,N_600);
nand U4502 (N_4502,N_819,N_603);
and U4503 (N_4503,N_516,N_2364);
xnor U4504 (N_4504,N_1710,N_2062);
and U4505 (N_4505,N_2089,N_795);
or U4506 (N_4506,N_1402,N_1311);
and U4507 (N_4507,N_1745,N_1122);
xnor U4508 (N_4508,N_1773,N_683);
nor U4509 (N_4509,N_2424,N_578);
nor U4510 (N_4510,N_1408,N_372);
or U4511 (N_4511,N_1230,N_2388);
nor U4512 (N_4512,N_937,N_1534);
nor U4513 (N_4513,N_447,N_2193);
and U4514 (N_4514,N_1403,N_845);
xor U4515 (N_4515,N_180,N_1076);
xnor U4516 (N_4516,N_1929,N_169);
or U4517 (N_4517,N_2214,N_1977);
nor U4518 (N_4518,N_7,N_1277);
xnor U4519 (N_4519,N_1272,N_2387);
and U4520 (N_4520,N_292,N_856);
and U4521 (N_4521,N_1300,N_1319);
nor U4522 (N_4522,N_1871,N_943);
or U4523 (N_4523,N_1636,N_1213);
and U4524 (N_4524,N_217,N_1629);
nor U4525 (N_4525,N_2301,N_964);
xnor U4526 (N_4526,N_979,N_1259);
xnor U4527 (N_4527,N_438,N_362);
nor U4528 (N_4528,N_2007,N_729);
or U4529 (N_4529,N_903,N_841);
nor U4530 (N_4530,N_1000,N_690);
xor U4531 (N_4531,N_1586,N_508);
or U4532 (N_4532,N_220,N_629);
or U4533 (N_4533,N_1183,N_2220);
xnor U4534 (N_4534,N_1773,N_727);
nor U4535 (N_4535,N_1470,N_1216);
xor U4536 (N_4536,N_1081,N_2334);
nor U4537 (N_4537,N_1682,N_435);
or U4538 (N_4538,N_112,N_818);
nor U4539 (N_4539,N_2154,N_2318);
nor U4540 (N_4540,N_25,N_1133);
nand U4541 (N_4541,N_2324,N_2410);
nand U4542 (N_4542,N_1213,N_978);
and U4543 (N_4543,N_1778,N_484);
nor U4544 (N_4544,N_257,N_2411);
nand U4545 (N_4545,N_1147,N_1330);
xor U4546 (N_4546,N_522,N_1499);
and U4547 (N_4547,N_2178,N_839);
or U4548 (N_4548,N_258,N_769);
xor U4549 (N_4549,N_2185,N_581);
or U4550 (N_4550,N_1760,N_245);
xor U4551 (N_4551,N_113,N_2082);
xnor U4552 (N_4552,N_271,N_908);
xnor U4553 (N_4553,N_915,N_2250);
nor U4554 (N_4554,N_1253,N_2015);
xor U4555 (N_4555,N_221,N_1362);
nand U4556 (N_4556,N_2426,N_1633);
nor U4557 (N_4557,N_947,N_1437);
nand U4558 (N_4558,N_448,N_1754);
nor U4559 (N_4559,N_179,N_1226);
or U4560 (N_4560,N_104,N_2096);
or U4561 (N_4561,N_845,N_638);
nor U4562 (N_4562,N_437,N_1691);
and U4563 (N_4563,N_667,N_393);
xnor U4564 (N_4564,N_408,N_1596);
nand U4565 (N_4565,N_214,N_540);
or U4566 (N_4566,N_38,N_160);
xor U4567 (N_4567,N_692,N_1474);
nand U4568 (N_4568,N_826,N_1151);
or U4569 (N_4569,N_314,N_303);
and U4570 (N_4570,N_854,N_1946);
xor U4571 (N_4571,N_638,N_1169);
nor U4572 (N_4572,N_76,N_131);
and U4573 (N_4573,N_1474,N_445);
nand U4574 (N_4574,N_368,N_58);
nor U4575 (N_4575,N_811,N_2119);
nor U4576 (N_4576,N_425,N_2312);
and U4577 (N_4577,N_1550,N_206);
nor U4578 (N_4578,N_954,N_229);
xnor U4579 (N_4579,N_1365,N_488);
and U4580 (N_4580,N_378,N_879);
and U4581 (N_4581,N_1331,N_1955);
and U4582 (N_4582,N_1179,N_1468);
xor U4583 (N_4583,N_1846,N_79);
or U4584 (N_4584,N_1760,N_2232);
nand U4585 (N_4585,N_1678,N_1828);
and U4586 (N_4586,N_1334,N_928);
nor U4587 (N_4587,N_353,N_1716);
nand U4588 (N_4588,N_1147,N_288);
or U4589 (N_4589,N_569,N_1294);
or U4590 (N_4590,N_1747,N_486);
nand U4591 (N_4591,N_722,N_2436);
nor U4592 (N_4592,N_1269,N_773);
nand U4593 (N_4593,N_1750,N_1166);
and U4594 (N_4594,N_1828,N_2044);
nand U4595 (N_4595,N_1260,N_258);
xnor U4596 (N_4596,N_1569,N_990);
nand U4597 (N_4597,N_1147,N_309);
nand U4598 (N_4598,N_1345,N_195);
nor U4599 (N_4599,N_2415,N_1100);
or U4600 (N_4600,N_598,N_502);
and U4601 (N_4601,N_1171,N_1459);
nor U4602 (N_4602,N_1592,N_713);
and U4603 (N_4603,N_183,N_1507);
or U4604 (N_4604,N_944,N_677);
xor U4605 (N_4605,N_417,N_239);
nor U4606 (N_4606,N_2066,N_234);
xnor U4607 (N_4607,N_1721,N_1058);
nand U4608 (N_4608,N_239,N_1205);
and U4609 (N_4609,N_1365,N_2040);
xnor U4610 (N_4610,N_1376,N_499);
xor U4611 (N_4611,N_615,N_161);
xor U4612 (N_4612,N_513,N_2202);
and U4613 (N_4613,N_1095,N_884);
nor U4614 (N_4614,N_2010,N_1156);
or U4615 (N_4615,N_266,N_1580);
xnor U4616 (N_4616,N_237,N_1823);
nand U4617 (N_4617,N_2489,N_776);
xnor U4618 (N_4618,N_13,N_890);
xor U4619 (N_4619,N_2376,N_1835);
and U4620 (N_4620,N_1287,N_124);
and U4621 (N_4621,N_2110,N_1152);
or U4622 (N_4622,N_1875,N_1614);
and U4623 (N_4623,N_997,N_1549);
or U4624 (N_4624,N_296,N_1923);
or U4625 (N_4625,N_2094,N_1249);
or U4626 (N_4626,N_69,N_1649);
nand U4627 (N_4627,N_1128,N_734);
xnor U4628 (N_4628,N_1474,N_2145);
nor U4629 (N_4629,N_52,N_332);
nor U4630 (N_4630,N_2039,N_2150);
or U4631 (N_4631,N_560,N_1054);
nand U4632 (N_4632,N_1503,N_2109);
or U4633 (N_4633,N_1639,N_338);
xor U4634 (N_4634,N_1464,N_1222);
or U4635 (N_4635,N_1552,N_188);
nor U4636 (N_4636,N_891,N_1532);
nand U4637 (N_4637,N_1877,N_62);
nor U4638 (N_4638,N_1344,N_1146);
nor U4639 (N_4639,N_815,N_1037);
nand U4640 (N_4640,N_1216,N_1262);
xor U4641 (N_4641,N_195,N_1580);
nor U4642 (N_4642,N_2479,N_1849);
xor U4643 (N_4643,N_2062,N_873);
nor U4644 (N_4644,N_1263,N_1457);
xor U4645 (N_4645,N_2224,N_943);
and U4646 (N_4646,N_2000,N_745);
and U4647 (N_4647,N_283,N_965);
nand U4648 (N_4648,N_866,N_1620);
xnor U4649 (N_4649,N_745,N_1724);
nor U4650 (N_4650,N_2453,N_1311);
nand U4651 (N_4651,N_2176,N_915);
or U4652 (N_4652,N_2149,N_595);
nand U4653 (N_4653,N_1439,N_15);
and U4654 (N_4654,N_1041,N_1233);
nand U4655 (N_4655,N_1290,N_586);
nand U4656 (N_4656,N_1130,N_1062);
nor U4657 (N_4657,N_995,N_783);
and U4658 (N_4658,N_1846,N_308);
nor U4659 (N_4659,N_606,N_888);
xnor U4660 (N_4660,N_1000,N_1713);
and U4661 (N_4661,N_624,N_578);
nor U4662 (N_4662,N_602,N_2303);
nand U4663 (N_4663,N_351,N_341);
nor U4664 (N_4664,N_2274,N_1307);
xor U4665 (N_4665,N_78,N_2048);
nand U4666 (N_4666,N_2075,N_1041);
xnor U4667 (N_4667,N_521,N_714);
nand U4668 (N_4668,N_226,N_529);
nand U4669 (N_4669,N_791,N_696);
nand U4670 (N_4670,N_1315,N_965);
or U4671 (N_4671,N_774,N_2148);
nor U4672 (N_4672,N_1678,N_1322);
nand U4673 (N_4673,N_2183,N_313);
or U4674 (N_4674,N_1328,N_1943);
xnor U4675 (N_4675,N_442,N_1720);
nand U4676 (N_4676,N_1228,N_890);
nor U4677 (N_4677,N_2319,N_805);
nor U4678 (N_4678,N_2308,N_980);
and U4679 (N_4679,N_86,N_1624);
nand U4680 (N_4680,N_1134,N_906);
or U4681 (N_4681,N_2013,N_692);
nor U4682 (N_4682,N_652,N_290);
or U4683 (N_4683,N_1867,N_948);
nor U4684 (N_4684,N_514,N_300);
nand U4685 (N_4685,N_1566,N_724);
or U4686 (N_4686,N_458,N_292);
and U4687 (N_4687,N_1097,N_1882);
nand U4688 (N_4688,N_876,N_1458);
nor U4689 (N_4689,N_2026,N_1833);
and U4690 (N_4690,N_1776,N_1418);
nor U4691 (N_4691,N_1617,N_2381);
xnor U4692 (N_4692,N_303,N_2436);
or U4693 (N_4693,N_1767,N_2431);
nand U4694 (N_4694,N_159,N_58);
and U4695 (N_4695,N_2057,N_2069);
nand U4696 (N_4696,N_1430,N_1728);
xnor U4697 (N_4697,N_1981,N_2068);
or U4698 (N_4698,N_2131,N_1573);
nor U4699 (N_4699,N_2283,N_1016);
nor U4700 (N_4700,N_1609,N_93);
and U4701 (N_4701,N_1007,N_211);
and U4702 (N_4702,N_391,N_1813);
nand U4703 (N_4703,N_673,N_502);
nor U4704 (N_4704,N_665,N_516);
nand U4705 (N_4705,N_1997,N_294);
nand U4706 (N_4706,N_1124,N_363);
xor U4707 (N_4707,N_1375,N_1532);
or U4708 (N_4708,N_1717,N_2458);
xnor U4709 (N_4709,N_711,N_1033);
xnor U4710 (N_4710,N_1993,N_2457);
nor U4711 (N_4711,N_1628,N_595);
and U4712 (N_4712,N_1840,N_2466);
xor U4713 (N_4713,N_1118,N_2297);
and U4714 (N_4714,N_1812,N_353);
xnor U4715 (N_4715,N_781,N_1681);
nor U4716 (N_4716,N_1959,N_2388);
and U4717 (N_4717,N_1231,N_114);
nand U4718 (N_4718,N_2244,N_1829);
or U4719 (N_4719,N_1407,N_1816);
or U4720 (N_4720,N_1787,N_1922);
nand U4721 (N_4721,N_110,N_1160);
and U4722 (N_4722,N_644,N_2263);
and U4723 (N_4723,N_573,N_1934);
nor U4724 (N_4724,N_1292,N_334);
nand U4725 (N_4725,N_768,N_704);
xnor U4726 (N_4726,N_2108,N_1382);
and U4727 (N_4727,N_629,N_690);
nor U4728 (N_4728,N_1854,N_2215);
nor U4729 (N_4729,N_340,N_1724);
and U4730 (N_4730,N_1979,N_711);
or U4731 (N_4731,N_1962,N_922);
nand U4732 (N_4732,N_1762,N_1764);
nand U4733 (N_4733,N_2287,N_951);
and U4734 (N_4734,N_26,N_1403);
nand U4735 (N_4735,N_10,N_2320);
or U4736 (N_4736,N_701,N_475);
nand U4737 (N_4737,N_1725,N_2368);
and U4738 (N_4738,N_566,N_1179);
and U4739 (N_4739,N_135,N_423);
or U4740 (N_4740,N_740,N_1187);
or U4741 (N_4741,N_1894,N_2053);
nor U4742 (N_4742,N_2403,N_2158);
nand U4743 (N_4743,N_2168,N_1964);
nand U4744 (N_4744,N_1425,N_506);
and U4745 (N_4745,N_708,N_934);
and U4746 (N_4746,N_301,N_1100);
or U4747 (N_4747,N_1845,N_589);
or U4748 (N_4748,N_923,N_2192);
and U4749 (N_4749,N_498,N_1223);
nand U4750 (N_4750,N_856,N_264);
or U4751 (N_4751,N_16,N_1615);
or U4752 (N_4752,N_57,N_1201);
xnor U4753 (N_4753,N_2182,N_1515);
nor U4754 (N_4754,N_2144,N_423);
or U4755 (N_4755,N_1171,N_854);
nor U4756 (N_4756,N_1727,N_1960);
xor U4757 (N_4757,N_2190,N_2159);
xor U4758 (N_4758,N_448,N_874);
xnor U4759 (N_4759,N_925,N_1789);
or U4760 (N_4760,N_769,N_2049);
nor U4761 (N_4761,N_1192,N_2008);
nand U4762 (N_4762,N_699,N_863);
or U4763 (N_4763,N_2103,N_1720);
xnor U4764 (N_4764,N_1194,N_1681);
and U4765 (N_4765,N_2201,N_1371);
nand U4766 (N_4766,N_1715,N_1322);
nand U4767 (N_4767,N_911,N_1436);
xnor U4768 (N_4768,N_187,N_486);
xnor U4769 (N_4769,N_2448,N_658);
or U4770 (N_4770,N_2150,N_1025);
or U4771 (N_4771,N_22,N_1314);
nand U4772 (N_4772,N_949,N_953);
xnor U4773 (N_4773,N_2360,N_1425);
or U4774 (N_4774,N_615,N_1125);
nand U4775 (N_4775,N_1322,N_1447);
or U4776 (N_4776,N_1214,N_1277);
and U4777 (N_4777,N_330,N_1024);
xnor U4778 (N_4778,N_835,N_2031);
nor U4779 (N_4779,N_316,N_2234);
and U4780 (N_4780,N_1949,N_1260);
xnor U4781 (N_4781,N_2218,N_1704);
nor U4782 (N_4782,N_943,N_1248);
or U4783 (N_4783,N_1383,N_530);
nand U4784 (N_4784,N_317,N_2132);
nor U4785 (N_4785,N_326,N_2455);
nor U4786 (N_4786,N_2104,N_1778);
nor U4787 (N_4787,N_1867,N_2050);
or U4788 (N_4788,N_2411,N_1730);
or U4789 (N_4789,N_179,N_606);
or U4790 (N_4790,N_1143,N_471);
nor U4791 (N_4791,N_709,N_694);
xnor U4792 (N_4792,N_1664,N_97);
or U4793 (N_4793,N_1315,N_758);
nand U4794 (N_4794,N_2126,N_1998);
or U4795 (N_4795,N_1952,N_138);
nor U4796 (N_4796,N_2466,N_456);
and U4797 (N_4797,N_107,N_498);
xor U4798 (N_4798,N_1032,N_1009);
nand U4799 (N_4799,N_760,N_1585);
nor U4800 (N_4800,N_456,N_1489);
nor U4801 (N_4801,N_2147,N_382);
and U4802 (N_4802,N_2139,N_1733);
nand U4803 (N_4803,N_844,N_804);
and U4804 (N_4804,N_406,N_915);
xnor U4805 (N_4805,N_575,N_554);
or U4806 (N_4806,N_994,N_51);
xor U4807 (N_4807,N_2013,N_1361);
or U4808 (N_4808,N_2463,N_2143);
nand U4809 (N_4809,N_1702,N_716);
and U4810 (N_4810,N_57,N_1349);
and U4811 (N_4811,N_1976,N_1149);
xor U4812 (N_4812,N_364,N_1548);
nor U4813 (N_4813,N_1958,N_930);
xor U4814 (N_4814,N_188,N_1901);
xnor U4815 (N_4815,N_839,N_2472);
nand U4816 (N_4816,N_2080,N_150);
xnor U4817 (N_4817,N_2412,N_785);
nand U4818 (N_4818,N_922,N_1551);
xor U4819 (N_4819,N_197,N_236);
or U4820 (N_4820,N_73,N_1966);
xnor U4821 (N_4821,N_572,N_2112);
or U4822 (N_4822,N_2455,N_2165);
nor U4823 (N_4823,N_687,N_1539);
and U4824 (N_4824,N_2467,N_1838);
xnor U4825 (N_4825,N_2426,N_2278);
and U4826 (N_4826,N_70,N_493);
nor U4827 (N_4827,N_1747,N_432);
nand U4828 (N_4828,N_212,N_31);
and U4829 (N_4829,N_1294,N_144);
or U4830 (N_4830,N_656,N_648);
nand U4831 (N_4831,N_659,N_1563);
nor U4832 (N_4832,N_1731,N_1771);
and U4833 (N_4833,N_2152,N_1730);
xor U4834 (N_4834,N_627,N_1974);
and U4835 (N_4835,N_998,N_474);
and U4836 (N_4836,N_1034,N_1469);
or U4837 (N_4837,N_1955,N_842);
and U4838 (N_4838,N_1492,N_1442);
or U4839 (N_4839,N_1447,N_34);
nand U4840 (N_4840,N_873,N_1455);
or U4841 (N_4841,N_2465,N_1430);
and U4842 (N_4842,N_636,N_982);
nor U4843 (N_4843,N_1242,N_1743);
xor U4844 (N_4844,N_1857,N_205);
nand U4845 (N_4845,N_1686,N_2432);
nand U4846 (N_4846,N_569,N_1060);
or U4847 (N_4847,N_910,N_2168);
nor U4848 (N_4848,N_311,N_2372);
nand U4849 (N_4849,N_857,N_1988);
nor U4850 (N_4850,N_421,N_1680);
nor U4851 (N_4851,N_431,N_323);
nand U4852 (N_4852,N_671,N_2459);
nor U4853 (N_4853,N_1413,N_2232);
and U4854 (N_4854,N_11,N_381);
xnor U4855 (N_4855,N_2016,N_2397);
xor U4856 (N_4856,N_2052,N_1776);
nand U4857 (N_4857,N_709,N_1146);
xor U4858 (N_4858,N_1745,N_2447);
nor U4859 (N_4859,N_685,N_240);
xnor U4860 (N_4860,N_901,N_1718);
nand U4861 (N_4861,N_1228,N_1019);
and U4862 (N_4862,N_762,N_1275);
and U4863 (N_4863,N_707,N_429);
xor U4864 (N_4864,N_562,N_884);
nand U4865 (N_4865,N_485,N_2037);
nand U4866 (N_4866,N_724,N_1753);
xnor U4867 (N_4867,N_1605,N_478);
nand U4868 (N_4868,N_1158,N_994);
or U4869 (N_4869,N_2090,N_1892);
nor U4870 (N_4870,N_1878,N_1629);
nor U4871 (N_4871,N_128,N_1397);
xnor U4872 (N_4872,N_1215,N_1174);
nor U4873 (N_4873,N_331,N_1301);
or U4874 (N_4874,N_353,N_2150);
nand U4875 (N_4875,N_1604,N_1072);
nand U4876 (N_4876,N_610,N_2093);
or U4877 (N_4877,N_1280,N_2480);
or U4878 (N_4878,N_1882,N_2277);
and U4879 (N_4879,N_1228,N_2323);
nand U4880 (N_4880,N_1373,N_1534);
or U4881 (N_4881,N_306,N_1024);
nor U4882 (N_4882,N_192,N_1296);
nand U4883 (N_4883,N_1194,N_494);
and U4884 (N_4884,N_2484,N_1113);
or U4885 (N_4885,N_1191,N_2291);
nor U4886 (N_4886,N_121,N_1373);
and U4887 (N_4887,N_1195,N_1799);
xnor U4888 (N_4888,N_47,N_177);
nor U4889 (N_4889,N_1025,N_1316);
nor U4890 (N_4890,N_1945,N_2171);
nand U4891 (N_4891,N_1363,N_2215);
nor U4892 (N_4892,N_87,N_1032);
nor U4893 (N_4893,N_943,N_1291);
nor U4894 (N_4894,N_1005,N_962);
or U4895 (N_4895,N_918,N_391);
xnor U4896 (N_4896,N_1824,N_1644);
or U4897 (N_4897,N_1140,N_1337);
nor U4898 (N_4898,N_1435,N_2273);
nand U4899 (N_4899,N_2457,N_10);
nand U4900 (N_4900,N_2107,N_1146);
and U4901 (N_4901,N_1707,N_618);
xnor U4902 (N_4902,N_1291,N_1935);
nand U4903 (N_4903,N_1099,N_287);
nand U4904 (N_4904,N_1429,N_2254);
nor U4905 (N_4905,N_646,N_1889);
or U4906 (N_4906,N_2024,N_270);
or U4907 (N_4907,N_291,N_354);
xor U4908 (N_4908,N_1843,N_793);
and U4909 (N_4909,N_1944,N_2142);
nand U4910 (N_4910,N_1398,N_685);
xnor U4911 (N_4911,N_422,N_2216);
nor U4912 (N_4912,N_1491,N_1074);
and U4913 (N_4913,N_475,N_1952);
nor U4914 (N_4914,N_54,N_425);
nor U4915 (N_4915,N_999,N_1804);
and U4916 (N_4916,N_2459,N_362);
or U4917 (N_4917,N_1578,N_2474);
xnor U4918 (N_4918,N_237,N_1204);
nand U4919 (N_4919,N_675,N_2330);
xnor U4920 (N_4920,N_1981,N_42);
xnor U4921 (N_4921,N_2490,N_69);
or U4922 (N_4922,N_1308,N_1707);
xor U4923 (N_4923,N_2072,N_1910);
and U4924 (N_4924,N_2098,N_105);
or U4925 (N_4925,N_263,N_935);
xor U4926 (N_4926,N_2314,N_1213);
or U4927 (N_4927,N_1365,N_2048);
or U4928 (N_4928,N_695,N_1133);
and U4929 (N_4929,N_1479,N_1533);
xor U4930 (N_4930,N_1608,N_1298);
and U4931 (N_4931,N_1351,N_356);
nor U4932 (N_4932,N_483,N_1628);
or U4933 (N_4933,N_970,N_417);
and U4934 (N_4934,N_1133,N_834);
xnor U4935 (N_4935,N_2291,N_1069);
or U4936 (N_4936,N_1857,N_1336);
nor U4937 (N_4937,N_910,N_221);
nand U4938 (N_4938,N_2133,N_1646);
xor U4939 (N_4939,N_1361,N_1043);
nand U4940 (N_4940,N_1577,N_8);
nand U4941 (N_4941,N_730,N_1678);
or U4942 (N_4942,N_602,N_1974);
and U4943 (N_4943,N_2137,N_382);
or U4944 (N_4944,N_1866,N_2328);
or U4945 (N_4945,N_2010,N_1866);
or U4946 (N_4946,N_1264,N_1772);
nor U4947 (N_4947,N_1233,N_1410);
and U4948 (N_4948,N_334,N_2338);
nand U4949 (N_4949,N_911,N_1528);
nand U4950 (N_4950,N_969,N_2075);
nor U4951 (N_4951,N_1130,N_1501);
xor U4952 (N_4952,N_801,N_1348);
nand U4953 (N_4953,N_206,N_167);
xnor U4954 (N_4954,N_2,N_1098);
or U4955 (N_4955,N_348,N_1156);
xor U4956 (N_4956,N_305,N_2284);
or U4957 (N_4957,N_727,N_147);
and U4958 (N_4958,N_435,N_1487);
nor U4959 (N_4959,N_1844,N_1739);
xor U4960 (N_4960,N_882,N_1923);
nand U4961 (N_4961,N_1762,N_2081);
or U4962 (N_4962,N_2455,N_2412);
or U4963 (N_4963,N_2065,N_2037);
and U4964 (N_4964,N_1848,N_2180);
xnor U4965 (N_4965,N_1555,N_496);
and U4966 (N_4966,N_1307,N_1675);
or U4967 (N_4967,N_1540,N_774);
nor U4968 (N_4968,N_234,N_2004);
xor U4969 (N_4969,N_1533,N_377);
nand U4970 (N_4970,N_846,N_2101);
nand U4971 (N_4971,N_2048,N_1312);
and U4972 (N_4972,N_522,N_2159);
nor U4973 (N_4973,N_1694,N_556);
and U4974 (N_4974,N_1761,N_431);
nor U4975 (N_4975,N_1814,N_64);
nand U4976 (N_4976,N_1573,N_265);
nand U4977 (N_4977,N_354,N_2430);
xnor U4978 (N_4978,N_1000,N_186);
and U4979 (N_4979,N_441,N_2467);
or U4980 (N_4980,N_1158,N_2427);
or U4981 (N_4981,N_1686,N_1906);
xor U4982 (N_4982,N_772,N_90);
nand U4983 (N_4983,N_2437,N_551);
and U4984 (N_4984,N_1495,N_852);
nand U4985 (N_4985,N_1861,N_2115);
xnor U4986 (N_4986,N_396,N_200);
and U4987 (N_4987,N_1428,N_382);
nor U4988 (N_4988,N_99,N_1061);
and U4989 (N_4989,N_2301,N_793);
and U4990 (N_4990,N_1938,N_1791);
or U4991 (N_4991,N_939,N_843);
or U4992 (N_4992,N_769,N_832);
nand U4993 (N_4993,N_337,N_1468);
and U4994 (N_4994,N_342,N_2290);
or U4995 (N_4995,N_1600,N_237);
nor U4996 (N_4996,N_1934,N_1438);
and U4997 (N_4997,N_1322,N_884);
nand U4998 (N_4998,N_1921,N_2130);
xnor U4999 (N_4999,N_1584,N_1974);
or U5000 (N_5000,N_4028,N_4702);
or U5001 (N_5001,N_2950,N_4160);
xor U5002 (N_5002,N_4378,N_4249);
nand U5003 (N_5003,N_4223,N_2962);
xnor U5004 (N_5004,N_4693,N_4845);
nand U5005 (N_5005,N_3478,N_3281);
or U5006 (N_5006,N_3545,N_3671);
nand U5007 (N_5007,N_4295,N_3130);
nand U5008 (N_5008,N_4641,N_4260);
nand U5009 (N_5009,N_3474,N_3405);
nor U5010 (N_5010,N_4317,N_3160);
nor U5011 (N_5011,N_4143,N_2589);
or U5012 (N_5012,N_2599,N_3053);
xor U5013 (N_5013,N_4785,N_3084);
and U5014 (N_5014,N_4145,N_3429);
or U5015 (N_5015,N_4895,N_2554);
or U5016 (N_5016,N_4154,N_3414);
xnor U5017 (N_5017,N_4089,N_4023);
nor U5018 (N_5018,N_4902,N_3180);
and U5019 (N_5019,N_4423,N_3852);
nand U5020 (N_5020,N_3468,N_3347);
xor U5021 (N_5021,N_3781,N_4220);
nand U5022 (N_5022,N_3629,N_3119);
nand U5023 (N_5023,N_3096,N_4933);
and U5024 (N_5024,N_2657,N_3584);
xnor U5025 (N_5025,N_2618,N_2863);
or U5026 (N_5026,N_3200,N_4903);
or U5027 (N_5027,N_4653,N_4024);
or U5028 (N_5028,N_4130,N_4180);
and U5029 (N_5029,N_3595,N_4385);
xor U5030 (N_5030,N_3668,N_4993);
and U5031 (N_5031,N_3390,N_4448);
nor U5032 (N_5032,N_3935,N_4603);
and U5033 (N_5033,N_4711,N_3460);
nand U5034 (N_5034,N_3503,N_4809);
nand U5035 (N_5035,N_3989,N_3889);
nor U5036 (N_5036,N_4998,N_3607);
and U5037 (N_5037,N_2829,N_4971);
xor U5038 (N_5038,N_2516,N_4112);
and U5039 (N_5039,N_3520,N_3375);
and U5040 (N_5040,N_3866,N_2854);
or U5041 (N_5041,N_3363,N_2750);
nor U5042 (N_5042,N_2563,N_4060);
and U5043 (N_5043,N_4324,N_3477);
nor U5044 (N_5044,N_4549,N_2893);
xor U5045 (N_5045,N_2576,N_4818);
and U5046 (N_5046,N_4339,N_3135);
or U5047 (N_5047,N_2556,N_3123);
nand U5048 (N_5048,N_2934,N_2600);
nand U5049 (N_5049,N_4616,N_3402);
and U5050 (N_5050,N_3634,N_3336);
and U5051 (N_5051,N_3069,N_3580);
and U5052 (N_5052,N_4842,N_4777);
xor U5053 (N_5053,N_2942,N_4128);
or U5054 (N_5054,N_2896,N_3490);
xnor U5055 (N_5055,N_2721,N_4783);
and U5056 (N_5056,N_2525,N_4577);
and U5057 (N_5057,N_4639,N_3100);
nor U5058 (N_5058,N_4999,N_4330);
xor U5059 (N_5059,N_3761,N_4623);
and U5060 (N_5060,N_3001,N_4586);
nor U5061 (N_5061,N_3941,N_3922);
nor U5062 (N_5062,N_3211,N_4564);
nor U5063 (N_5063,N_3071,N_3717);
or U5064 (N_5064,N_4765,N_4788);
xnor U5065 (N_5065,N_3996,N_2875);
nand U5066 (N_5066,N_4228,N_2695);
or U5067 (N_5067,N_3558,N_4259);
or U5068 (N_5068,N_4408,N_3527);
nor U5069 (N_5069,N_2637,N_4253);
nand U5070 (N_5070,N_2931,N_4874);
or U5071 (N_5071,N_3698,N_3563);
xnor U5072 (N_5072,N_4437,N_3279);
or U5073 (N_5073,N_4728,N_3877);
and U5074 (N_5074,N_4012,N_3117);
and U5075 (N_5075,N_4410,N_3859);
or U5076 (N_5076,N_4663,N_3846);
nand U5077 (N_5077,N_3099,N_4994);
or U5078 (N_5078,N_3713,N_2597);
xnor U5079 (N_5079,N_2763,N_3173);
or U5080 (N_5080,N_4900,N_3514);
and U5081 (N_5081,N_3658,N_4397);
and U5082 (N_5082,N_2997,N_2892);
and U5083 (N_5083,N_3313,N_2545);
nor U5084 (N_5084,N_3526,N_4794);
or U5085 (N_5085,N_3222,N_3716);
nor U5086 (N_5086,N_4735,N_2538);
xor U5087 (N_5087,N_3942,N_4951);
nor U5088 (N_5088,N_3861,N_2617);
xnor U5089 (N_5089,N_4924,N_4161);
nor U5090 (N_5090,N_3983,N_3087);
xnor U5091 (N_5091,N_4395,N_3155);
xor U5092 (N_5092,N_3720,N_4801);
or U5093 (N_5093,N_3554,N_2921);
nor U5094 (N_5094,N_3733,N_3725);
nand U5095 (N_5095,N_4747,N_3093);
or U5096 (N_5096,N_4309,N_2676);
and U5097 (N_5097,N_4310,N_4950);
and U5098 (N_5098,N_4977,N_3268);
nor U5099 (N_5099,N_4347,N_4188);
xnor U5100 (N_5100,N_4399,N_4019);
nor U5101 (N_5101,N_4961,N_2666);
or U5102 (N_5102,N_4480,N_3938);
xnor U5103 (N_5103,N_4512,N_4943);
xor U5104 (N_5104,N_4468,N_4532);
nor U5105 (N_5105,N_4667,N_4001);
nand U5106 (N_5106,N_2838,N_4888);
and U5107 (N_5107,N_3463,N_4827);
nor U5108 (N_5108,N_2552,N_4167);
nor U5109 (N_5109,N_3351,N_4569);
nor U5110 (N_5110,N_3420,N_2996);
nor U5111 (N_5111,N_2639,N_3752);
xor U5112 (N_5112,N_2782,N_2543);
xnor U5113 (N_5113,N_3924,N_4633);
nor U5114 (N_5114,N_3748,N_3743);
xnor U5115 (N_5115,N_4715,N_2794);
nor U5116 (N_5116,N_3749,N_2880);
and U5117 (N_5117,N_3711,N_3524);
nor U5118 (N_5118,N_3505,N_4732);
xor U5119 (N_5119,N_3359,N_3872);
nor U5120 (N_5120,N_4445,N_3699);
or U5121 (N_5121,N_3328,N_4414);
and U5122 (N_5122,N_3926,N_3642);
nor U5123 (N_5123,N_3059,N_3330);
nor U5124 (N_5124,N_3814,N_3194);
and U5125 (N_5125,N_3774,N_4617);
and U5126 (N_5126,N_3339,N_4336);
or U5127 (N_5127,N_3611,N_4053);
or U5128 (N_5128,N_3113,N_3101);
nor U5129 (N_5129,N_4748,N_4926);
or U5130 (N_5130,N_2603,N_2746);
nand U5131 (N_5131,N_4579,N_2566);
or U5132 (N_5132,N_2923,N_4505);
nor U5133 (N_5133,N_4450,N_3192);
and U5134 (N_5134,N_4604,N_4707);
nand U5135 (N_5135,N_2963,N_4521);
nand U5136 (N_5136,N_3236,N_4609);
nor U5137 (N_5137,N_3254,N_2990);
xnor U5138 (N_5138,N_4102,N_4153);
or U5139 (N_5139,N_4919,N_3483);
nor U5140 (N_5140,N_3432,N_4029);
nor U5141 (N_5141,N_3754,N_4236);
xor U5142 (N_5142,N_3032,N_2508);
nor U5143 (N_5143,N_3435,N_4830);
nand U5144 (N_5144,N_4773,N_4768);
and U5145 (N_5145,N_4490,N_4529);
or U5146 (N_5146,N_3147,N_3516);
nor U5147 (N_5147,N_2752,N_4911);
and U5148 (N_5148,N_3309,N_3930);
or U5149 (N_5149,N_4590,N_3450);
nand U5150 (N_5150,N_2675,N_3470);
nand U5151 (N_5151,N_4956,N_2581);
nor U5152 (N_5152,N_3849,N_4120);
nand U5153 (N_5153,N_4519,N_2672);
nor U5154 (N_5154,N_3887,N_4074);
and U5155 (N_5155,N_3971,N_2805);
nand U5156 (N_5156,N_3455,N_4214);
and U5157 (N_5157,N_2674,N_4033);
xnor U5158 (N_5158,N_3547,N_4449);
xor U5159 (N_5159,N_2661,N_3571);
xnor U5160 (N_5160,N_3240,N_2653);
nand U5161 (N_5161,N_2799,N_4257);
nor U5162 (N_5162,N_4816,N_4698);
and U5163 (N_5163,N_3341,N_3002);
or U5164 (N_5164,N_3488,N_4456);
or U5165 (N_5165,N_3204,N_3386);
nor U5166 (N_5166,N_2646,N_4864);
or U5167 (N_5167,N_2774,N_4492);
nand U5168 (N_5168,N_4857,N_3462);
and U5169 (N_5169,N_3756,N_2885);
and U5170 (N_5170,N_3045,N_4756);
nand U5171 (N_5171,N_3937,N_4200);
and U5172 (N_5172,N_3835,N_3810);
or U5173 (N_5173,N_4158,N_4557);
or U5174 (N_5174,N_4051,N_2640);
nand U5175 (N_5175,N_4184,N_3539);
nor U5176 (N_5176,N_4194,N_3424);
nand U5177 (N_5177,N_3140,N_4493);
xor U5178 (N_5178,N_4806,N_4644);
or U5179 (N_5179,N_3449,N_3657);
or U5180 (N_5180,N_2770,N_4871);
nor U5181 (N_5181,N_2976,N_3706);
and U5182 (N_5182,N_4566,N_3290);
or U5183 (N_5183,N_3316,N_4418);
and U5184 (N_5184,N_4186,N_3479);
and U5185 (N_5185,N_3320,N_3112);
xnor U5186 (N_5186,N_3688,N_3573);
xnor U5187 (N_5187,N_4246,N_2729);
nand U5188 (N_5188,N_3158,N_4042);
xor U5189 (N_5189,N_4093,N_4988);
and U5190 (N_5190,N_2788,N_4299);
nand U5191 (N_5191,N_3960,N_4750);
and U5192 (N_5192,N_4782,N_2908);
xor U5193 (N_5193,N_4542,N_2687);
nand U5194 (N_5194,N_4137,N_2680);
xor U5195 (N_5195,N_4099,N_4591);
or U5196 (N_5196,N_2755,N_3104);
nor U5197 (N_5197,N_3667,N_3932);
xor U5198 (N_5198,N_2502,N_4851);
or U5199 (N_5199,N_2699,N_3624);
nor U5200 (N_5200,N_3065,N_4491);
and U5201 (N_5201,N_3610,N_4092);
and U5202 (N_5202,N_3355,N_2647);
and U5203 (N_5203,N_2866,N_3023);
xor U5204 (N_5204,N_2784,N_4925);
and U5205 (N_5205,N_3793,N_2801);
and U5206 (N_5206,N_3257,N_4537);
or U5207 (N_5207,N_3900,N_4858);
and U5208 (N_5208,N_4442,N_3251);
nand U5209 (N_5209,N_3874,N_3530);
and U5210 (N_5210,N_3466,N_3740);
nor U5211 (N_5211,N_2883,N_4247);
xor U5212 (N_5212,N_4831,N_4985);
and U5213 (N_5213,N_3929,N_4095);
nor U5214 (N_5214,N_2772,N_4274);
and U5215 (N_5215,N_2771,N_4032);
xnor U5216 (N_5216,N_2937,N_2621);
xnor U5217 (N_5217,N_2605,N_4912);
nor U5218 (N_5218,N_2590,N_4034);
and U5219 (N_5219,N_3256,N_4567);
or U5220 (N_5220,N_4196,N_3796);
and U5221 (N_5221,N_3805,N_3606);
and U5222 (N_5222,N_2822,N_2503);
and U5223 (N_5223,N_4428,N_3788);
and U5224 (N_5224,N_2722,N_3430);
or U5225 (N_5225,N_4381,N_4780);
nand U5226 (N_5226,N_4968,N_4435);
or U5227 (N_5227,N_3618,N_2871);
and U5228 (N_5228,N_2933,N_4642);
and U5229 (N_5229,N_4499,N_4561);
xnor U5230 (N_5230,N_4386,N_4531);
or U5231 (N_5231,N_2660,N_3213);
or U5232 (N_5232,N_4689,N_4893);
nand U5233 (N_5233,N_2751,N_4573);
nor U5234 (N_5234,N_3304,N_4524);
nand U5235 (N_5235,N_3364,N_3982);
xor U5236 (N_5236,N_4256,N_2724);
nand U5237 (N_5237,N_4219,N_2717);
nor U5238 (N_5238,N_3288,N_2807);
xor U5239 (N_5239,N_3311,N_4345);
and U5240 (N_5240,N_4975,N_4664);
nand U5241 (N_5241,N_2993,N_3225);
and U5242 (N_5242,N_3380,N_4387);
nand U5243 (N_5243,N_2733,N_4122);
xnor U5244 (N_5244,N_3409,N_4821);
and U5245 (N_5245,N_2864,N_2865);
nor U5246 (N_5246,N_4085,N_2671);
xnor U5247 (N_5247,N_4458,N_3764);
xnor U5248 (N_5248,N_3946,N_4477);
xnor U5249 (N_5249,N_2927,N_4930);
or U5250 (N_5250,N_3569,N_3063);
nor U5251 (N_5251,N_3763,N_2626);
or U5252 (N_5252,N_3722,N_3917);
nand U5253 (N_5253,N_3145,N_3831);
nor U5254 (N_5254,N_3593,N_4904);
nand U5255 (N_5255,N_2564,N_3437);
xor U5256 (N_5256,N_4587,N_3510);
nor U5257 (N_5257,N_4036,N_2814);
nand U5258 (N_5258,N_4181,N_2796);
and U5259 (N_5259,N_4856,N_2941);
nor U5260 (N_5260,N_4212,N_4031);
nor U5261 (N_5261,N_3552,N_3305);
xor U5262 (N_5262,N_3597,N_3999);
xor U5263 (N_5263,N_3948,N_4726);
xor U5264 (N_5264,N_3915,N_2940);
and U5265 (N_5265,N_4280,N_3438);
or U5266 (N_5266,N_3888,N_2585);
xor U5267 (N_5267,N_2586,N_4126);
and U5268 (N_5268,N_3858,N_4147);
xor U5269 (N_5269,N_4133,N_3659);
nand U5270 (N_5270,N_3945,N_3739);
xnor U5271 (N_5271,N_4081,N_4610);
nor U5272 (N_5272,N_4100,N_3841);
or U5273 (N_5273,N_2810,N_3442);
xnor U5274 (N_5274,N_4357,N_4189);
or U5275 (N_5275,N_3548,N_4670);
nor U5276 (N_5276,N_3675,N_4709);
nand U5277 (N_5277,N_3321,N_4880);
or U5278 (N_5278,N_2766,N_3689);
xnor U5279 (N_5279,N_4771,N_2943);
nor U5280 (N_5280,N_4276,N_4284);
or U5281 (N_5281,N_3684,N_2749);
nand U5282 (N_5282,N_3406,N_4764);
and U5283 (N_5283,N_3780,N_3031);
and U5284 (N_5284,N_3056,N_3966);
and U5285 (N_5285,N_4578,N_4742);
or U5286 (N_5286,N_3102,N_3700);
nor U5287 (N_5287,N_3994,N_3857);
and U5288 (N_5288,N_3324,N_4142);
xnor U5289 (N_5289,N_4839,N_4621);
or U5290 (N_5290,N_4206,N_4679);
and U5291 (N_5291,N_3591,N_2951);
nand U5292 (N_5292,N_4749,N_4662);
or U5293 (N_5293,N_4101,N_2759);
nand U5294 (N_5294,N_3010,N_3656);
nand U5295 (N_5295,N_4465,N_4854);
nor U5296 (N_5296,N_4928,N_4955);
nand U5297 (N_5297,N_3775,N_4453);
xnor U5298 (N_5298,N_4175,N_2999);
nand U5299 (N_5299,N_4834,N_2507);
nor U5300 (N_5300,N_4164,N_3559);
xnor U5301 (N_5301,N_3776,N_4103);
or U5302 (N_5302,N_3838,N_3197);
and U5303 (N_5303,N_4277,N_4565);
and U5304 (N_5304,N_4369,N_3893);
xor U5305 (N_5305,N_4022,N_3701);
and U5306 (N_5306,N_4407,N_4358);
and U5307 (N_5307,N_3286,N_2677);
xnor U5308 (N_5308,N_4430,N_3970);
and U5309 (N_5309,N_2648,N_4232);
xnor U5310 (N_5310,N_2691,N_4426);
nor U5311 (N_5311,N_4043,N_3864);
xnor U5312 (N_5312,N_3609,N_3266);
nor U5313 (N_5313,N_4231,N_4302);
nand U5314 (N_5314,N_3444,N_4680);
or U5315 (N_5315,N_4504,N_3750);
nand U5316 (N_5316,N_4649,N_3677);
and U5317 (N_5317,N_4287,N_3987);
and U5318 (N_5318,N_2910,N_3376);
xor U5319 (N_5319,N_2684,N_3961);
xor U5320 (N_5320,N_3895,N_4296);
and U5321 (N_5321,N_4607,N_3074);
xor U5322 (N_5322,N_3440,N_4114);
and U5323 (N_5323,N_3785,N_3078);
nor U5324 (N_5324,N_3519,N_2862);
xnor U5325 (N_5325,N_3974,N_3291);
nand U5326 (N_5326,N_4406,N_2913);
or U5327 (N_5327,N_2935,N_4073);
nor U5328 (N_5328,N_3804,N_3331);
xor U5329 (N_5329,N_3789,N_3878);
xor U5330 (N_5330,N_3738,N_3374);
and U5331 (N_5331,N_4351,N_3068);
or U5332 (N_5332,N_3019,N_4755);
and U5333 (N_5333,N_3518,N_4250);
xnor U5334 (N_5334,N_3976,N_2549);
nor U5335 (N_5335,N_4479,N_4337);
xor U5336 (N_5336,N_2938,N_3315);
or U5337 (N_5337,N_3057,N_4983);
xnor U5338 (N_5338,N_3207,N_4234);
nand U5339 (N_5339,N_3267,N_4486);
and U5340 (N_5340,N_2781,N_4601);
xnor U5341 (N_5341,N_4384,N_4963);
and U5342 (N_5342,N_2632,N_2539);
xnor U5343 (N_5343,N_3826,N_3105);
nand U5344 (N_5344,N_3821,N_3760);
and U5345 (N_5345,N_2904,N_4551);
or U5346 (N_5346,N_4113,N_2567);
or U5347 (N_5347,N_4808,N_3367);
nor U5348 (N_5348,N_4338,N_2841);
nand U5349 (N_5349,N_3992,N_2592);
and U5350 (N_5350,N_4522,N_4373);
nand U5351 (N_5351,N_2848,N_4940);
nor U5352 (N_5352,N_3777,N_4965);
xor U5353 (N_5353,N_4058,N_3718);
nor U5354 (N_5354,N_4527,N_3036);
nand U5355 (N_5355,N_2870,N_4300);
or U5356 (N_5356,N_4534,N_3332);
xor U5357 (N_5357,N_3020,N_3410);
xnor U5358 (N_5358,N_2656,N_4533);
nor U5359 (N_5359,N_3890,N_4572);
or U5360 (N_5360,N_3249,N_3651);
nand U5361 (N_5361,N_3049,N_3600);
xor U5362 (N_5362,N_3428,N_4222);
xnor U5363 (N_5363,N_3674,N_4979);
nor U5364 (N_5364,N_4767,N_2555);
and U5365 (N_5365,N_4318,N_3378);
and U5366 (N_5366,N_4245,N_4471);
nor U5367 (N_5367,N_3497,N_4064);
xnor U5368 (N_5368,N_3521,N_2630);
nand U5369 (N_5369,N_3195,N_4240);
xnor U5370 (N_5370,N_4770,N_3543);
or U5371 (N_5371,N_2665,N_2629);
nand U5372 (N_5372,N_3737,N_3744);
xnor U5373 (N_5373,N_2988,N_4897);
nand U5374 (N_5374,N_4626,N_4847);
nand U5375 (N_5375,N_2688,N_4651);
nor U5376 (N_5376,N_4570,N_3177);
nand U5377 (N_5377,N_4424,N_2740);
nand U5378 (N_5378,N_4674,N_2624);
or U5379 (N_5379,N_4271,N_3034);
nor U5380 (N_5380,N_4119,N_4068);
nand U5381 (N_5381,N_4684,N_3417);
nand U5382 (N_5382,N_4535,N_4889);
and U5383 (N_5383,N_3388,N_4306);
and U5384 (N_5384,N_4786,N_2915);
nand U5385 (N_5385,N_2681,N_3469);
nand U5386 (N_5386,N_2728,N_4322);
xnor U5387 (N_5387,N_3778,N_3903);
and U5388 (N_5388,N_3511,N_4138);
xor U5389 (N_5389,N_3964,N_2778);
and U5390 (N_5390,N_4297,N_4706);
nand U5391 (N_5391,N_4511,N_4953);
nor U5392 (N_5392,N_3076,N_3404);
and U5393 (N_5393,N_3392,N_2505);
nand U5394 (N_5394,N_4867,N_2966);
nand U5395 (N_5395,N_3095,N_2984);
or U5396 (N_5396,N_4813,N_3116);
nor U5397 (N_5397,N_4731,N_3604);
nand U5398 (N_5398,N_3090,N_3370);
nor U5399 (N_5399,N_3564,N_3953);
nand U5400 (N_5400,N_4576,N_4152);
or U5401 (N_5401,N_4021,N_3995);
nand U5402 (N_5402,N_2668,N_4636);
nor U5403 (N_5403,N_4800,N_4185);
nor U5404 (N_5404,N_2884,N_4461);
or U5405 (N_5405,N_2610,N_4195);
and U5406 (N_5406,N_3823,N_4072);
or U5407 (N_5407,N_4191,N_4090);
or U5408 (N_5408,N_4778,N_3608);
nor U5409 (N_5409,N_2912,N_2557);
nor U5410 (N_5410,N_4860,N_3928);
or U5411 (N_5411,N_2500,N_2738);
xor U5412 (N_5412,N_4941,N_4992);
and U5413 (N_5413,N_4620,N_2523);
and U5414 (N_5414,N_4681,N_2909);
nor U5415 (N_5415,N_2911,N_3208);
nand U5416 (N_5416,N_4356,N_3813);
or U5417 (N_5417,N_2849,N_3244);
nand U5418 (N_5418,N_3845,N_3787);
xor U5419 (N_5419,N_2808,N_4745);
xor U5420 (N_5420,N_3017,N_3719);
or U5421 (N_5421,N_3220,N_4314);
nand U5422 (N_5422,N_4252,N_3692);
and U5423 (N_5423,N_4002,N_3683);
and U5424 (N_5424,N_4835,N_3797);
nand U5425 (N_5425,N_3308,N_4417);
nand U5426 (N_5426,N_3144,N_4478);
and U5427 (N_5427,N_2536,N_3565);
xor U5428 (N_5428,N_3799,N_4515);
and U5429 (N_5429,N_3847,N_3221);
nor U5430 (N_5430,N_4432,N_3985);
and U5431 (N_5431,N_3421,N_4721);
or U5432 (N_5432,N_4371,N_2548);
nor U5433 (N_5433,N_2850,N_2767);
nor U5434 (N_5434,N_3199,N_3529);
nand U5435 (N_5435,N_3512,N_2878);
xor U5436 (N_5436,N_2887,N_3843);
xnor U5437 (N_5437,N_4613,N_3284);
nor U5438 (N_5438,N_4077,N_4402);
or U5439 (N_5439,N_4910,N_3264);
nor U5440 (N_5440,N_3923,N_2588);
nor U5441 (N_5441,N_2775,N_3492);
nand U5442 (N_5442,N_4415,N_3471);
xnor U5443 (N_5443,N_3769,N_4906);
or U5444 (N_5444,N_4921,N_3633);
xor U5445 (N_5445,N_2812,N_4469);
or U5446 (N_5446,N_3491,N_2867);
nor U5447 (N_5447,N_4362,N_4346);
nor U5448 (N_5448,N_4473,N_3579);
nor U5449 (N_5449,N_4270,N_4920);
nand U5450 (N_5450,N_2920,N_2537);
and U5451 (N_5451,N_2987,N_4420);
nor U5452 (N_5452,N_2819,N_3252);
nor U5453 (N_5453,N_2673,N_4327);
xor U5454 (N_5454,N_2710,N_3784);
and U5455 (N_5455,N_4929,N_3574);
xor U5456 (N_5456,N_2795,N_4949);
xnor U5457 (N_5457,N_4224,N_4648);
nand U5458 (N_5458,N_4331,N_4198);
nor U5459 (N_5459,N_3083,N_2991);
nor U5460 (N_5460,N_4054,N_4497);
xor U5461 (N_5461,N_4343,N_4342);
or U5462 (N_5462,N_3475,N_3549);
and U5463 (N_5463,N_3327,N_4563);
xnor U5464 (N_5464,N_2723,N_2919);
xnor U5465 (N_5465,N_2888,N_4263);
and U5466 (N_5466,N_3918,N_2527);
xor U5467 (N_5467,N_4879,N_2765);
nor U5468 (N_5468,N_3476,N_3802);
or U5469 (N_5469,N_2818,N_3586);
nor U5470 (N_5470,N_4111,N_3272);
or U5471 (N_5471,N_4392,N_4766);
nor U5472 (N_5472,N_2968,N_2664);
or U5473 (N_5473,N_3854,N_4503);
and U5474 (N_5474,N_4934,N_3661);
nand U5475 (N_5475,N_3980,N_3653);
and U5476 (N_5476,N_3914,N_3384);
xnor U5477 (N_5477,N_4107,N_4025);
nor U5478 (N_5478,N_2961,N_3731);
nand U5479 (N_5479,N_2957,N_4506);
or U5480 (N_5480,N_4733,N_4538);
nor U5481 (N_5481,N_2736,N_3660);
xnor U5482 (N_5482,N_2598,N_3235);
or U5483 (N_5483,N_3832,N_3024);
nand U5484 (N_5484,N_4575,N_2542);
and U5485 (N_5485,N_2758,N_4098);
xnor U5486 (N_5486,N_3919,N_4526);
or U5487 (N_5487,N_2670,N_2965);
and U5488 (N_5488,N_3030,N_3818);
and U5489 (N_5489,N_4853,N_4848);
or U5490 (N_5490,N_4552,N_3152);
xor U5491 (N_5491,N_3369,N_2792);
xor U5492 (N_5492,N_3840,N_3958);
nand U5493 (N_5493,N_2611,N_4482);
nor U5494 (N_5494,N_3707,N_3957);
nor U5495 (N_5495,N_3048,N_4326);
nor U5496 (N_5496,N_4622,N_3396);
and U5497 (N_5497,N_3502,N_4365);
nand U5498 (N_5498,N_4837,N_4991);
nor U5499 (N_5499,N_3183,N_4516);
and U5500 (N_5500,N_3016,N_4394);
nand U5501 (N_5501,N_3379,N_4488);
xnor U5502 (N_5502,N_3292,N_3907);
or U5503 (N_5503,N_4823,N_4737);
or U5504 (N_5504,N_3461,N_2924);
nand U5505 (N_5505,N_3570,N_3865);
nand U5506 (N_5506,N_4462,N_3730);
nand U5507 (N_5507,N_3081,N_3773);
nor U5508 (N_5508,N_4624,N_3464);
nor U5509 (N_5509,N_2694,N_3362);
xor U5510 (N_5510,N_3500,N_4230);
or U5511 (N_5511,N_3169,N_4170);
nor U5512 (N_5512,N_4692,N_3551);
nor U5513 (N_5513,N_3012,N_3422);
and U5514 (N_5514,N_4182,N_4980);
xor U5515 (N_5515,N_2873,N_2715);
nand U5516 (N_5516,N_2645,N_3694);
xor U5517 (N_5517,N_3310,N_2541);
nand U5518 (N_5518,N_3663,N_4872);
nand U5519 (N_5519,N_4132,N_3086);
and U5520 (N_5520,N_3058,N_3956);
nand U5521 (N_5521,N_3097,N_3753);
nor U5522 (N_5522,N_4937,N_4353);
or U5523 (N_5523,N_4183,N_4976);
xor U5524 (N_5524,N_4832,N_4226);
nand U5525 (N_5525,N_4390,N_3599);
nor U5526 (N_5526,N_2816,N_4454);
and U5527 (N_5527,N_4915,N_4429);
and U5528 (N_5528,N_2732,N_2761);
xor U5529 (N_5529,N_4055,N_2747);
and U5530 (N_5530,N_2712,N_3867);
or U5531 (N_5531,N_3704,N_4714);
nand U5532 (N_5532,N_3517,N_4760);
xor U5533 (N_5533,N_3913,N_3615);
nor U5534 (N_5534,N_2817,N_2620);
xor U5535 (N_5535,N_3216,N_3039);
nor U5536 (N_5536,N_4070,N_3578);
or U5537 (N_5537,N_4753,N_3356);
nor U5538 (N_5538,N_3652,N_3226);
or U5539 (N_5539,N_2793,N_3817);
nand U5540 (N_5540,N_4974,N_3839);
or U5541 (N_5541,N_4608,N_3842);
nor U5542 (N_5542,N_3171,N_4014);
and U5543 (N_5543,N_2789,N_4774);
nand U5544 (N_5544,N_4141,N_4746);
nor U5545 (N_5545,N_3897,N_2926);
nand U5546 (N_5546,N_2979,N_2847);
nor U5547 (N_5547,N_3300,N_4123);
nand U5548 (N_5548,N_3920,N_2619);
nor U5549 (N_5549,N_4761,N_3168);
and U5550 (N_5550,N_3085,N_4550);
and U5551 (N_5551,N_4628,N_3898);
nand U5552 (N_5552,N_2859,N_4606);
nand U5553 (N_5553,N_3515,N_3886);
xnor U5554 (N_5554,N_3088,N_2769);
or U5555 (N_5555,N_2949,N_4638);
or U5556 (N_5556,N_3952,N_2995);
or U5557 (N_5557,N_2826,N_3345);
nor U5558 (N_5558,N_2574,N_4716);
and U5559 (N_5559,N_3441,N_3334);
and U5560 (N_5560,N_2669,N_4878);
or U5561 (N_5561,N_4555,N_3077);
or U5562 (N_5562,N_3879,N_3128);
nand U5563 (N_5563,N_4556,N_3285);
nor U5564 (N_5564,N_2930,N_2783);
or U5565 (N_5565,N_3975,N_3951);
nor U5566 (N_5566,N_3686,N_4265);
nand U5567 (N_5567,N_2852,N_4229);
and U5568 (N_5568,N_4901,N_2768);
xnor U5569 (N_5569,N_4009,N_4094);
nand U5570 (N_5570,N_3612,N_4713);
nand U5571 (N_5571,N_4688,N_2559);
and U5572 (N_5572,N_3142,N_4932);
and U5573 (N_5573,N_3448,N_4584);
and U5574 (N_5574,N_2726,N_2655);
and U5575 (N_5575,N_3206,N_2890);
or U5576 (N_5576,N_4740,N_4248);
xnor U5577 (N_5577,N_3275,N_4850);
nor U5578 (N_5578,N_3723,N_2686);
xor U5579 (N_5579,N_3747,N_3260);
nand U5580 (N_5580,N_4401,N_3294);
or U5581 (N_5581,N_2868,N_4292);
xor U5582 (N_5582,N_4166,N_4614);
and U5583 (N_5583,N_3990,N_3714);
nor U5584 (N_5584,N_3513,N_3185);
and U5585 (N_5585,N_4789,N_3227);
nand U5586 (N_5586,N_4916,N_2820);
or U5587 (N_5587,N_3679,N_4599);
and U5588 (N_5588,N_3301,N_2622);
nand U5589 (N_5589,N_3230,N_2546);
nand U5590 (N_5590,N_2705,N_4637);
nor U5591 (N_5591,N_3669,N_3157);
xnor U5592 (N_5592,N_4391,N_2569);
and U5593 (N_5593,N_3270,N_3191);
nor U5594 (N_5594,N_3954,N_4776);
or U5595 (N_5595,N_3427,N_2886);
nand U5596 (N_5596,N_2744,N_2727);
or U5597 (N_5597,N_2840,N_3025);
nand U5598 (N_5598,N_2623,N_4091);
nor U5599 (N_5599,N_4811,N_4056);
and U5600 (N_5600,N_3638,N_2693);
or U5601 (N_5601,N_4944,N_4290);
nor U5602 (N_5602,N_4541,N_3094);
nor U5603 (N_5603,N_3602,N_4797);
nor U5604 (N_5604,N_4078,N_3029);
or U5605 (N_5605,N_4382,N_4079);
nand U5606 (N_5606,N_4155,N_4836);
nor U5607 (N_5607,N_2753,N_2832);
and U5608 (N_5608,N_4207,N_4312);
nand U5609 (N_5609,N_4457,N_4481);
or U5610 (N_5610,N_4596,N_3873);
nor U5611 (N_5611,N_4255,N_3628);
nor U5612 (N_5612,N_4543,N_3746);
and U5613 (N_5613,N_3209,N_3115);
xor U5614 (N_5614,N_3419,N_3592);
xor U5615 (N_5615,N_2916,N_4597);
xnor U5616 (N_5616,N_4377,N_4464);
and U5617 (N_5617,N_3871,N_4507);
or U5618 (N_5618,N_4927,N_4704);
nor U5619 (N_5619,N_4865,N_4589);
nand U5620 (N_5620,N_4677,N_4687);
nand U5621 (N_5621,N_3273,N_4440);
or U5622 (N_5622,N_4877,N_3542);
xnor U5623 (N_5623,N_3767,N_4443);
or U5624 (N_5624,N_3385,N_2627);
xor U5625 (N_5625,N_2524,N_4697);
nand U5626 (N_5626,N_2651,N_3625);
nand U5627 (N_5627,N_3150,N_3916);
or U5628 (N_5628,N_3153,N_4380);
xor U5629 (N_5629,N_2650,N_4554);
or U5630 (N_5630,N_4121,N_3408);
nand U5631 (N_5631,N_4973,N_3397);
nand U5632 (N_5632,N_3060,N_2899);
nand U5633 (N_5633,N_3891,N_4738);
nor U5634 (N_5634,N_4987,N_3742);
and U5635 (N_5635,N_4177,N_3959);
nor U5636 (N_5636,N_3977,N_4258);
and U5637 (N_5637,N_4793,N_4208);
nand U5638 (N_5638,N_2800,N_3506);
nor U5639 (N_5639,N_4388,N_4805);
xnor U5640 (N_5640,N_4173,N_4855);
and U5641 (N_5641,N_4763,N_4870);
or U5642 (N_5642,N_3936,N_4598);
nor U5643 (N_5643,N_2764,N_2553);
or U5644 (N_5644,N_3052,N_4799);
nor U5645 (N_5645,N_4124,N_4050);
or U5646 (N_5646,N_4190,N_3955);
nand U5647 (N_5647,N_4625,N_4046);
nor U5648 (N_5648,N_3646,N_3536);
nor U5649 (N_5649,N_4049,N_4108);
or U5650 (N_5650,N_3636,N_4668);
xor U5651 (N_5651,N_3280,N_4825);
xor U5652 (N_5652,N_3523,N_4463);
or U5653 (N_5653,N_3705,N_4741);
nor U5654 (N_5654,N_4447,N_2845);
and U5655 (N_5655,N_3346,N_3546);
or U5656 (N_5656,N_2992,N_4913);
nor U5657 (N_5657,N_4898,N_3111);
or U5658 (N_5658,N_2986,N_3166);
nand U5659 (N_5659,N_3482,N_3972);
or U5660 (N_5660,N_2571,N_4446);
nor U5661 (N_5661,N_3695,N_2803);
nor U5662 (N_5662,N_4852,N_4425);
xor U5663 (N_5663,N_2714,N_4011);
nand U5664 (N_5664,N_2901,N_4413);
nor U5665 (N_5665,N_2785,N_2628);
or U5666 (N_5666,N_4320,N_4374);
nand U5667 (N_5667,N_4724,N_4683);
nand U5668 (N_5668,N_3443,N_3027);
and U5669 (N_5669,N_4080,N_4370);
xor U5670 (N_5670,N_3232,N_3412);
xor U5671 (N_5671,N_3507,N_3141);
xnor U5672 (N_5672,N_4217,N_4631);
nor U5673 (N_5673,N_2519,N_4673);
xor U5674 (N_5674,N_2609,N_3413);
and U5675 (N_5675,N_2972,N_4313);
xnor U5676 (N_5676,N_2874,N_4015);
or U5677 (N_5677,N_4939,N_4238);
xor U5678 (N_5678,N_2725,N_2635);
and U5679 (N_5679,N_4873,N_3931);
and U5680 (N_5680,N_3269,N_3054);
xnor U5681 (N_5681,N_2654,N_4643);
nand U5682 (N_5682,N_2633,N_2956);
nand U5683 (N_5683,N_2696,N_3892);
and U5684 (N_5684,N_3391,N_2815);
xor U5685 (N_5685,N_3008,N_4333);
and U5686 (N_5686,N_3454,N_3837);
and U5687 (N_5687,N_2946,N_3998);
or U5688 (N_5688,N_3768,N_3394);
nand U5689 (N_5689,N_4148,N_3734);
xor U5690 (N_5690,N_4700,N_3993);
and U5691 (N_5691,N_2702,N_3358);
and U5692 (N_5692,N_2989,N_3556);
nor U5693 (N_5693,N_2550,N_2692);
nor U5694 (N_5694,N_2575,N_4118);
or U5695 (N_5695,N_3106,N_3472);
and U5696 (N_5696,N_3073,N_4989);
xnor U5697 (N_5697,N_3485,N_3589);
xnor U5698 (N_5698,N_3883,N_2877);
nand U5699 (N_5699,N_3164,N_2894);
or U5700 (N_5700,N_2683,N_4179);
nor U5701 (N_5701,N_2971,N_3991);
xor U5702 (N_5702,N_2804,N_3433);
xnor U5703 (N_5703,N_4485,N_2882);
and U5704 (N_5704,N_4176,N_4192);
nor U5705 (N_5705,N_4455,N_4409);
xnor U5706 (N_5706,N_4896,N_4585);
or U5707 (N_5707,N_4376,N_4798);
nor U5708 (N_5708,N_4588,N_4048);
nand U5709 (N_5709,N_3237,N_4935);
and U5710 (N_5710,N_4654,N_3423);
and U5711 (N_5711,N_4293,N_4517);
xor U5712 (N_5712,N_4129,N_4332);
nand U5713 (N_5713,N_4618,N_3357);
nand U5714 (N_5714,N_4757,N_3314);
or U5715 (N_5715,N_3909,N_3863);
nor U5716 (N_5716,N_3765,N_4282);
xnor U5717 (N_5717,N_2577,N_3555);
and U5718 (N_5718,N_4861,N_3757);
nor U5719 (N_5719,N_2649,N_3820);
or U5720 (N_5720,N_4883,N_3137);
and U5721 (N_5721,N_4082,N_3038);
or U5722 (N_5722,N_4187,N_2613);
or U5723 (N_5723,N_2960,N_2745);
and U5724 (N_5724,N_3870,N_3203);
nand U5725 (N_5725,N_2970,N_4734);
and U5726 (N_5726,N_2827,N_3156);
or U5727 (N_5727,N_4162,N_3299);
or U5728 (N_5728,N_3418,N_3801);
xnor U5729 (N_5729,N_3447,N_4412);
xnor U5730 (N_5730,N_4807,N_2953);
and U5731 (N_5731,N_4354,N_4722);
nor U5732 (N_5732,N_2638,N_4434);
nor U5733 (N_5733,N_3484,N_4421);
nand U5734 (N_5734,N_4205,N_3735);
nand U5735 (N_5735,N_3855,N_4595);
or U5736 (N_5736,N_2734,N_4719);
or U5737 (N_5737,N_4890,N_4914);
or U5738 (N_5738,N_3303,N_4665);
nand U5739 (N_5739,N_3274,N_2791);
nand U5740 (N_5740,N_4841,N_4892);
or U5741 (N_5741,N_3218,N_3779);
xor U5742 (N_5742,N_3333,N_3884);
xnor U5743 (N_5743,N_3988,N_3533);
or U5744 (N_5744,N_4026,N_3557);
or U5745 (N_5745,N_2662,N_2678);
nand U5746 (N_5746,N_2925,N_3561);
and U5747 (N_5747,N_4057,N_4945);
or U5748 (N_5748,N_3389,N_3535);
or U5749 (N_5749,N_3504,N_3581);
or U5750 (N_5750,N_3912,N_4936);
xor U5751 (N_5751,N_3772,N_4352);
nor U5752 (N_5752,N_3210,N_4329);
nand U5753 (N_5753,N_3415,N_2607);
nand U5754 (N_5754,N_2634,N_4069);
xor U5755 (N_5755,N_2568,N_4146);
or U5756 (N_5756,N_3005,N_3649);
nand U5757 (N_5757,N_3650,N_2790);
nand U5758 (N_5758,N_4694,N_3021);
nor U5759 (N_5759,N_3467,N_3498);
and U5760 (N_5760,N_2903,N_4967);
and U5761 (N_5761,N_4115,N_3107);
xnor U5762 (N_5762,N_2700,N_3337);
nand U5763 (N_5763,N_2530,N_3702);
or U5764 (N_5764,N_3184,N_4545);
or U5765 (N_5765,N_3493,N_2707);
or U5766 (N_5766,N_2839,N_4005);
xnor U5767 (N_5767,N_3253,N_4824);
nor U5768 (N_5768,N_3407,N_3148);
and U5769 (N_5769,N_2601,N_4514);
or U5770 (N_5770,N_4475,N_4105);
and U5771 (N_5771,N_2615,N_3261);
nand U5772 (N_5772,N_3576,N_3967);
nand U5773 (N_5773,N_3676,N_3302);
nand U5774 (N_5774,N_4946,N_4539);
and U5775 (N_5775,N_3224,N_4273);
or U5776 (N_5776,N_3182,N_4630);
nor U5777 (N_5777,N_2526,N_2501);
and U5778 (N_5778,N_4459,N_4403);
nand U5779 (N_5779,N_2853,N_4784);
and U5780 (N_5780,N_4203,N_3165);
and U5781 (N_5781,N_4995,N_4303);
xor U5782 (N_5782,N_4917,N_3587);
and U5783 (N_5783,N_4483,N_3899);
and U5784 (N_5784,N_3544,N_4316);
xnor U5785 (N_5785,N_3670,N_3834);
and U5786 (N_5786,N_3451,N_4661);
xnor U5787 (N_5787,N_3151,N_3037);
nand U5788 (N_5788,N_3630,N_4163);
or U5789 (N_5789,N_2980,N_3910);
nor U5790 (N_5790,N_4752,N_3572);
nand U5791 (N_5791,N_2658,N_4136);
or U5792 (N_5792,N_4308,N_3631);
nor U5793 (N_5793,N_3042,N_4075);
nand U5794 (N_5794,N_3340,N_3550);
and U5795 (N_5795,N_3902,N_4822);
nand U5796 (N_5796,N_3908,N_3641);
xnor U5797 (N_5797,N_3446,N_4204);
xor U5798 (N_5798,N_3129,N_3577);
nand U5799 (N_5799,N_4061,N_2708);
nor U5800 (N_5800,N_2514,N_2876);
and U5801 (N_5801,N_2842,N_4862);
xor U5802 (N_5802,N_3620,N_4087);
nand U5803 (N_5803,N_4691,N_4268);
or U5804 (N_5804,N_3033,N_4990);
nor U5805 (N_5805,N_4779,N_3118);
nor U5806 (N_5806,N_2998,N_3181);
and U5807 (N_5807,N_4718,N_4659);
nand U5808 (N_5808,N_3381,N_3335);
and U5809 (N_5809,N_4829,N_4510);
nor U5810 (N_5810,N_2813,N_3758);
nand U5811 (N_5811,N_4452,N_2720);
xor U5812 (N_5812,N_4281,N_4682);
nand U5813 (N_5813,N_3494,N_4159);
nand U5814 (N_5814,N_4172,N_2958);
or U5815 (N_5815,N_3473,N_4398);
and U5816 (N_5816,N_4518,N_3803);
or U5817 (N_5817,N_3828,N_4954);
xnor U5818 (N_5818,N_4605,N_2825);
nor U5819 (N_5819,N_3921,N_2735);
and U5820 (N_5820,N_4218,N_2978);
or U5821 (N_5821,N_3567,N_2891);
nor U5822 (N_5822,N_3426,N_4466);
nand U5823 (N_5823,N_2706,N_3277);
or U5824 (N_5824,N_3973,N_2625);
or U5825 (N_5825,N_3499,N_2558);
and U5826 (N_5826,N_4363,N_4144);
xor U5827 (N_5827,N_3904,N_2587);
xor U5828 (N_5828,N_4952,N_3163);
and U5829 (N_5829,N_3354,N_3905);
xor U5830 (N_5830,N_4328,N_4086);
xor U5831 (N_5831,N_2719,N_4427);
nand U5832 (N_5832,N_4416,N_4508);
nor U5833 (N_5833,N_3265,N_4233);
nand U5834 (N_5834,N_2964,N_2663);
or U5835 (N_5835,N_3596,N_4361);
xor U5836 (N_5836,N_3070,N_3349);
or U5837 (N_5837,N_2974,N_3896);
nor U5838 (N_5838,N_2612,N_2897);
and U5839 (N_5839,N_4938,N_3372);
or U5840 (N_5840,N_4020,N_4758);
and U5841 (N_5841,N_4264,N_4730);
nor U5842 (N_5842,N_3594,N_3968);
nor U5843 (N_5843,N_2529,N_3127);
or U5844 (N_5844,N_2535,N_4059);
nand U5845 (N_5845,N_3040,N_4484);
xnor U5846 (N_5846,N_2914,N_3343);
and U5847 (N_5847,N_4960,N_4071);
xnor U5848 (N_5848,N_3233,N_2947);
or U5849 (N_5849,N_3170,N_3283);
nor U5850 (N_5850,N_2830,N_4199);
nand U5851 (N_5851,N_2616,N_4635);
and U5852 (N_5852,N_4727,N_3811);
nand U5853 (N_5853,N_4658,N_3082);
nand U5854 (N_5854,N_3186,N_3262);
and U5855 (N_5855,N_3189,N_3637);
or U5856 (N_5856,N_3617,N_4235);
or U5857 (N_5857,N_4710,N_4476);
and U5858 (N_5858,N_3215,N_4215);
xor U5859 (N_5859,N_2544,N_4307);
and U5860 (N_5860,N_3647,N_4838);
nor U5861 (N_5861,N_3361,N_4819);
and U5862 (N_5862,N_4360,N_4627);
nand U5863 (N_5863,N_3969,N_3238);
or U5864 (N_5864,N_4431,N_2918);
nor U5865 (N_5865,N_4411,N_3348);
xor U5866 (N_5866,N_2510,N_4027);
or U5867 (N_5867,N_3825,N_3673);
or U5868 (N_5868,N_4869,N_3727);
and U5869 (N_5869,N_2518,N_2737);
and U5870 (N_5870,N_4640,N_3242);
or U5871 (N_5871,N_3809,N_3133);
nor U5872 (N_5872,N_3000,N_4574);
nand U5873 (N_5873,N_3271,N_3827);
xor U5874 (N_5874,N_4083,N_3124);
nand U5875 (N_5875,N_4134,N_2561);
or U5876 (N_5876,N_3202,N_3149);
nor U5877 (N_5877,N_4052,N_3243);
xnor U5878 (N_5878,N_4237,N_2823);
nor U5879 (N_5879,N_3495,N_3296);
or U5880 (N_5880,N_4866,N_3786);
and U5881 (N_5881,N_4396,N_3175);
nor U5882 (N_5882,N_2929,N_3295);
and U5883 (N_5883,N_2762,N_3962);
or U5884 (N_5884,N_4918,N_4695);
and U5885 (N_5885,N_3205,N_4404);
nor U5886 (N_5886,N_3004,N_3822);
nand U5887 (N_5887,N_3187,N_3055);
nand U5888 (N_5888,N_3212,N_4859);
xnor U5889 (N_5889,N_2718,N_4405);
or U5890 (N_5890,N_2509,N_2836);
nor U5891 (N_5891,N_4562,N_4969);
or U5892 (N_5892,N_3648,N_4289);
nor U5893 (N_5893,N_4547,N_3368);
or U5894 (N_5894,N_2948,N_4210);
or U5895 (N_5895,N_4812,N_3815);
nand U5896 (N_5896,N_3496,N_2835);
and U5897 (N_5897,N_3219,N_4803);
xor U5898 (N_5898,N_2973,N_3325);
xnor U5899 (N_5899,N_3880,N_4242);
or U5900 (N_5900,N_3806,N_4775);
xnor U5901 (N_5901,N_4593,N_2779);
nand U5902 (N_5902,N_3072,N_4010);
xnor U5903 (N_5903,N_3134,N_2560);
and U5904 (N_5904,N_3457,N_4559);
xor U5905 (N_5905,N_4045,N_4581);
nor U5906 (N_5906,N_4611,N_3795);
or U5907 (N_5907,N_3627,N_4340);
or U5908 (N_5908,N_2730,N_3963);
nand U5909 (N_5909,N_3366,N_3881);
nand U5910 (N_5910,N_4171,N_2690);
nor U5911 (N_5911,N_3289,N_4729);
xor U5912 (N_5912,N_2540,N_3940);
and U5913 (N_5913,N_2757,N_3680);
and U5914 (N_5914,N_4736,N_3508);
or U5915 (N_5915,N_3729,N_2583);
nor U5916 (N_5916,N_3585,N_3259);
xor U5917 (N_5917,N_4006,N_4467);
and U5918 (N_5918,N_3139,N_4787);
nor U5919 (N_5919,N_3708,N_3439);
nand U5920 (N_5920,N_2591,N_3736);
nor U5921 (N_5921,N_4520,N_3293);
nor U5922 (N_5922,N_3161,N_4804);
nand U5923 (N_5923,N_2967,N_3603);
xnor U5924 (N_5924,N_4041,N_4923);
nand U5925 (N_5925,N_4843,N_3480);
or U5926 (N_5926,N_4451,N_3196);
nor U5927 (N_5927,N_4619,N_3721);
nor U5928 (N_5928,N_4725,N_3486);
nor U5929 (N_5929,N_3401,N_4846);
nand U5930 (N_5930,N_4004,N_4422);
nand U5931 (N_5931,N_3687,N_2928);
xor U5932 (N_5932,N_4876,N_4686);
nand U5933 (N_5933,N_3009,N_3067);
nand U5934 (N_5934,N_4239,N_4127);
xnor U5935 (N_5935,N_3856,N_4349);
nor U5936 (N_5936,N_3614,N_2858);
and U5937 (N_5937,N_2572,N_2506);
xnor U5938 (N_5938,N_3122,N_2739);
nand U5939 (N_5939,N_3400,N_4335);
or U5940 (N_5940,N_4321,N_2584);
xor U5941 (N_5941,N_2905,N_4227);
and U5942 (N_5942,N_3245,N_4393);
xnor U5943 (N_5943,N_3509,N_4826);
and U5944 (N_5944,N_3015,N_4592);
nor U5945 (N_5945,N_4820,N_3399);
nor U5946 (N_5946,N_3051,N_2869);
nor U5947 (N_5947,N_3681,N_4178);
or U5948 (N_5948,N_2824,N_4583);
or U5949 (N_5949,N_4254,N_4344);
nand U5950 (N_5950,N_4495,N_4494);
nand U5951 (N_5951,N_3431,N_3353);
nand U5952 (N_5952,N_2922,N_2698);
xnor U5953 (N_5953,N_4213,N_3934);
nor U5954 (N_5954,N_2685,N_3198);
xor U5955 (N_5955,N_3131,N_3605);
xor U5956 (N_5956,N_3635,N_2756);
xor U5957 (N_5957,N_3875,N_4802);
nand U5958 (N_5958,N_3541,N_3553);
nand U5959 (N_5959,N_4251,N_3782);
nor U5960 (N_5960,N_4000,N_4436);
and U5961 (N_5961,N_2975,N_3812);
nor U5962 (N_5962,N_4366,N_4844);
nor U5963 (N_5963,N_3329,N_4632);
and U5964 (N_5964,N_3808,N_2573);
nor U5965 (N_5965,N_3064,N_4016);
or U5966 (N_5966,N_2955,N_3282);
nor U5967 (N_5967,N_2833,N_4037);
nand U5968 (N_5968,N_3986,N_4174);
xor U5969 (N_5969,N_3745,N_4833);
and U5970 (N_5970,N_2631,N_4548);
or U5971 (N_5971,N_3231,N_4571);
xor U5972 (N_5972,N_4894,N_3062);
and U5973 (N_5973,N_3678,N_4647);
and U5974 (N_5974,N_4646,N_2593);
nor U5975 (N_5975,N_3089,N_3125);
nor U5976 (N_5976,N_4815,N_4907);
nand U5977 (N_5977,N_2837,N_3682);
nor U5978 (N_5978,N_3398,N_3666);
or U5979 (N_5979,N_2906,N_4209);
and U5980 (N_5980,N_4221,N_4690);
nand U5981 (N_5981,N_4286,N_4168);
xor U5982 (N_5982,N_4262,N_3885);
nand U5983 (N_5983,N_3382,N_3790);
or U5984 (N_5984,N_3800,N_4319);
nand U5985 (N_5985,N_4882,N_3287);
nand U5986 (N_5986,N_3247,N_4272);
or U5987 (N_5987,N_2522,N_3317);
or U5988 (N_5988,N_2977,N_3297);
and U5989 (N_5989,N_3613,N_4544);
or U5990 (N_5990,N_3710,N_4193);
nor U5991 (N_5991,N_4959,N_4165);
nor U5992 (N_5992,N_4400,N_4754);
nand U5993 (N_5993,N_3014,N_3436);
nor U5994 (N_5994,N_2679,N_3759);
nor U5995 (N_5995,N_3755,N_3632);
or U5996 (N_5996,N_3724,N_3120);
or U5997 (N_5997,N_4602,N_4225);
nor U5998 (N_5998,N_4795,N_4645);
xor U5999 (N_5999,N_2532,N_3532);
nor U6000 (N_6000,N_3829,N_4678);
and U6001 (N_6001,N_3146,N_4600);
or U6002 (N_6002,N_4868,N_3126);
nand U6003 (N_6003,N_2602,N_4350);
nor U6004 (N_6004,N_2802,N_3223);
or U6005 (N_6005,N_4769,N_2697);
nand U6006 (N_6006,N_4849,N_4814);
xor U6007 (N_6007,N_3732,N_2855);
nand U6008 (N_6008,N_4097,N_3143);
xor U6009 (N_6009,N_2982,N_2944);
nor U6010 (N_6010,N_3393,N_4047);
nor U6011 (N_6011,N_3352,N_4044);
xnor U6012 (N_6012,N_4699,N_3853);
or U6013 (N_6013,N_4884,N_2932);
or U6014 (N_6014,N_4796,N_4275);
nand U6015 (N_6015,N_2512,N_3950);
xor U6016 (N_6016,N_3132,N_3538);
nor U6017 (N_6017,N_3465,N_4109);
nand U6018 (N_6018,N_3154,N_3848);
or U6019 (N_6019,N_4744,N_2643);
or U6020 (N_6020,N_3819,N_4372);
or U6021 (N_6021,N_2716,N_3091);
and U6022 (N_6022,N_3850,N_3006);
xnor U6023 (N_6023,N_4285,N_4007);
or U6024 (N_6024,N_4291,N_4294);
or U6025 (N_6025,N_2743,N_4283);
nand U6026 (N_6026,N_4996,N_2682);
nand U6027 (N_6027,N_4062,N_3360);
nor U6028 (N_6028,N_4367,N_3395);
or U6029 (N_6029,N_4040,N_4017);
xnor U6030 (N_6030,N_3026,N_4672);
nand U6031 (N_6031,N_3176,N_4978);
nand U6032 (N_6032,N_4003,N_3568);
nand U6033 (N_6033,N_4540,N_2809);
and U6034 (N_6034,N_2641,N_2900);
or U6035 (N_6035,N_3179,N_3121);
nand U6036 (N_6036,N_4066,N_3013);
nor U6037 (N_6037,N_4762,N_4886);
or U6038 (N_6038,N_3623,N_4759);
or U6039 (N_6039,N_4110,N_4964);
or U6040 (N_6040,N_4594,N_3943);
xnor U6041 (N_6041,N_4546,N_3619);
nand U6042 (N_6042,N_3947,N_4666);
nor U6043 (N_6043,N_4530,N_3639);
xnor U6044 (N_6044,N_3978,N_4984);
and U6045 (N_6045,N_4982,N_3869);
nand U6046 (N_6046,N_2604,N_3217);
nor U6047 (N_6047,N_3174,N_3640);
nand U6048 (N_6048,N_4169,N_4151);
or U6049 (N_6049,N_4261,N_4135);
or U6050 (N_6050,N_4629,N_3007);
or U6051 (N_6051,N_2534,N_3644);
nand U6052 (N_6052,N_4197,N_3047);
and U6053 (N_6053,N_3583,N_3824);
and U6054 (N_6054,N_3453,N_4355);
nand U6055 (N_6055,N_2843,N_3159);
nand U6056 (N_6056,N_4781,N_3691);
and U6057 (N_6057,N_2709,N_2857);
and U6058 (N_6058,N_2741,N_3981);
or U6059 (N_6059,N_3851,N_3540);
and U6060 (N_6060,N_2511,N_3690);
xor U6061 (N_6061,N_3318,N_3456);
or U6062 (N_6062,N_4139,N_3387);
nand U6063 (N_6063,N_2856,N_3061);
and U6064 (N_6064,N_3601,N_4669);
xor U6065 (N_6065,N_3685,N_3248);
nand U6066 (N_6066,N_4474,N_4751);
nor U6067 (N_6067,N_4791,N_2551);
nand U6068 (N_6068,N_4065,N_3836);
nor U6069 (N_6069,N_2713,N_3662);
xnor U6070 (N_6070,N_3307,N_4106);
nor U6071 (N_6071,N_2861,N_2748);
xor U6072 (N_6072,N_2579,N_3562);
or U6073 (N_6073,N_4922,N_3697);
nor U6074 (N_6074,N_2834,N_3911);
nand U6075 (N_6075,N_4441,N_3167);
and U6076 (N_6076,N_3258,N_2945);
nand U6077 (N_6077,N_2760,N_4439);
xor U6078 (N_6078,N_4558,N_4650);
or U6079 (N_6079,N_3933,N_3043);
xnor U6080 (N_6080,N_3050,N_3894);
nand U6081 (N_6081,N_3214,N_3762);
or U6082 (N_6082,N_2659,N_4810);
xor U6083 (N_6083,N_4500,N_4887);
or U6084 (N_6084,N_4298,N_4931);
or U6085 (N_6085,N_4509,N_3979);
or U6086 (N_6086,N_4067,N_3138);
or U6087 (N_6087,N_4553,N_4875);
nand U6088 (N_6088,N_4266,N_3771);
nand U6089 (N_6089,N_3582,N_4671);
xor U6090 (N_6090,N_4685,N_3193);
or U6091 (N_6091,N_4840,N_2703);
nor U6092 (N_6092,N_3751,N_2582);
nor U6093 (N_6093,N_3255,N_4948);
xnor U6094 (N_6094,N_3766,N_4038);
nor U6095 (N_6095,N_4301,N_3445);
and U6096 (N_6096,N_3528,N_4359);
xor U6097 (N_6097,N_4063,N_4018);
nand U6098 (N_6098,N_3188,N_3712);
nand U6099 (N_6099,N_3862,N_2786);
nand U6100 (N_6100,N_2731,N_4970);
xor U6101 (N_6101,N_3306,N_4241);
or U6102 (N_6102,N_2939,N_4131);
xor U6103 (N_6103,N_2570,N_4202);
or U6104 (N_6104,N_4657,N_4885);
nor U6105 (N_6105,N_3365,N_4039);
xnor U6106 (N_6106,N_4905,N_3537);
xnor U6107 (N_6107,N_2580,N_3590);
and U6108 (N_6108,N_3246,N_3110);
nor U6109 (N_6109,N_4792,N_3342);
or U6110 (N_6110,N_4304,N_4279);
or U6111 (N_6111,N_3298,N_4568);
nor U6112 (N_6112,N_3103,N_3487);
or U6113 (N_6113,N_3075,N_3018);
nor U6114 (N_6114,N_2828,N_3939);
xnor U6115 (N_6115,N_2644,N_2898);
or U6116 (N_6116,N_3035,N_3228);
or U6117 (N_6117,N_4723,N_3984);
nand U6118 (N_6118,N_4966,N_3098);
xor U6119 (N_6119,N_3654,N_4696);
xor U6120 (N_6120,N_4899,N_2533);
nor U6121 (N_6121,N_4149,N_3276);
xor U6122 (N_6122,N_4523,N_3522);
or U6123 (N_6123,N_4348,N_4243);
nor U6124 (N_6124,N_3411,N_3525);
or U6125 (N_6125,N_4580,N_2969);
xnor U6126 (N_6126,N_3868,N_4501);
and U6127 (N_6127,N_3575,N_3250);
nand U6128 (N_6128,N_3028,N_3876);
nand U6129 (N_6129,N_3882,N_4828);
xor U6130 (N_6130,N_4502,N_3598);
xor U6131 (N_6131,N_4315,N_2831);
nand U6132 (N_6132,N_2851,N_3621);
nor U6133 (N_6133,N_2936,N_4817);
nand U6134 (N_6134,N_3965,N_4717);
or U6135 (N_6135,N_3997,N_3622);
and U6136 (N_6136,N_2565,N_4612);
xor U6137 (N_6137,N_4772,N_4323);
and U6138 (N_6138,N_2798,N_3344);
nand U6139 (N_6139,N_3136,N_2811);
and U6140 (N_6140,N_2952,N_4157);
xnor U6141 (N_6141,N_4368,N_2860);
nor U6142 (N_6142,N_4278,N_3531);
xor U6143 (N_6143,N_3906,N_4334);
nand U6144 (N_6144,N_2667,N_3792);
xor U6145 (N_6145,N_4660,N_4201);
nand U6146 (N_6146,N_2821,N_4125);
nor U6147 (N_6147,N_3114,N_3459);
nand U6148 (N_6148,N_3626,N_4008);
nand U6149 (N_6149,N_2520,N_4957);
nand U6150 (N_6150,N_3377,N_3791);
nand U6151 (N_6151,N_2595,N_3655);
and U6152 (N_6152,N_3373,N_3278);
and U6153 (N_6153,N_4364,N_4444);
nor U6154 (N_6154,N_4881,N_2513);
or U6155 (N_6155,N_3949,N_2844);
nand U6156 (N_6156,N_2606,N_3709);
xnor U6157 (N_6157,N_2531,N_4470);
nor U6158 (N_6158,N_4675,N_3794);
nand U6159 (N_6159,N_2776,N_2954);
nor U6160 (N_6160,N_3481,N_3319);
nor U6161 (N_6161,N_4720,N_4582);
or U6162 (N_6162,N_4433,N_4419);
xor U6163 (N_6163,N_3833,N_3925);
nand U6164 (N_6164,N_4076,N_2994);
and U6165 (N_6165,N_3190,N_3489);
or U6166 (N_6166,N_2872,N_4088);
xor U6167 (N_6167,N_3927,N_2704);
xor U6168 (N_6168,N_3665,N_3066);
or U6169 (N_6169,N_4104,N_4655);
and U6170 (N_6170,N_3108,N_3741);
nor U6171 (N_6171,N_4389,N_3044);
nor U6172 (N_6172,N_3229,N_4150);
nor U6173 (N_6173,N_4013,N_2881);
and U6174 (N_6174,N_4708,N_3798);
nand U6175 (N_6175,N_2594,N_2596);
xnor U6176 (N_6176,N_4096,N_3645);
nand U6177 (N_6177,N_4117,N_4035);
nor U6178 (N_6178,N_4863,N_4460);
nand U6179 (N_6179,N_4743,N_3588);
nand U6180 (N_6180,N_3452,N_2889);
and U6181 (N_6181,N_2689,N_3046);
or U6182 (N_6182,N_2642,N_4375);
nand U6183 (N_6183,N_3323,N_2959);
or U6184 (N_6184,N_4942,N_3696);
or U6185 (N_6185,N_3178,N_4311);
nor U6186 (N_6186,N_4244,N_3534);
or U6187 (N_6187,N_4615,N_2636);
nor U6188 (N_6188,N_3162,N_2701);
nand U6189 (N_6189,N_2806,N_4498);
nand U6190 (N_6190,N_3434,N_2917);
and U6191 (N_6191,N_4305,N_4288);
nor U6192 (N_6192,N_3022,N_3715);
nand U6193 (N_6193,N_4496,N_3728);
or U6194 (N_6194,N_2652,N_2711);
nand U6195 (N_6195,N_4958,N_4116);
nand U6196 (N_6196,N_4536,N_2797);
nand U6197 (N_6197,N_4528,N_3350);
nor U6198 (N_6198,N_2614,N_3239);
nand U6199 (N_6199,N_3566,N_4560);
and U6200 (N_6200,N_4341,N_3616);
nand U6201 (N_6201,N_3901,N_4676);
nand U6202 (N_6202,N_4084,N_3326);
or U6203 (N_6203,N_4705,N_4981);
xor U6204 (N_6204,N_2981,N_4739);
nor U6205 (N_6205,N_3079,N_4267);
nor U6206 (N_6206,N_4472,N_3860);
nor U6207 (N_6207,N_3172,N_3263);
nor U6208 (N_6208,N_3383,N_2846);
xnor U6209 (N_6209,N_4891,N_2504);
or U6210 (N_6210,N_4962,N_3672);
xor U6211 (N_6211,N_2547,N_3312);
nor U6212 (N_6212,N_3322,N_3830);
xor U6213 (N_6213,N_4947,N_3201);
and U6214 (N_6214,N_3770,N_4986);
and U6215 (N_6215,N_3080,N_4634);
xor U6216 (N_6216,N_2895,N_4972);
nor U6217 (N_6217,N_4489,N_3416);
nand U6218 (N_6218,N_3425,N_3783);
xor U6219 (N_6219,N_3458,N_3944);
and U6220 (N_6220,N_2907,N_2983);
and U6221 (N_6221,N_2517,N_4908);
nand U6222 (N_6222,N_2780,N_3003);
nor U6223 (N_6223,N_4790,N_4513);
nor U6224 (N_6224,N_4997,N_2773);
nor U6225 (N_6225,N_4269,N_4030);
or U6226 (N_6226,N_2787,N_2742);
nand U6227 (N_6227,N_4140,N_4379);
nand U6228 (N_6228,N_2608,N_2521);
nor U6229 (N_6229,N_3703,N_4712);
or U6230 (N_6230,N_3338,N_4156);
or U6231 (N_6231,N_3816,N_4438);
and U6232 (N_6232,N_3844,N_2985);
or U6233 (N_6233,N_4325,N_3011);
nor U6234 (N_6234,N_2528,N_3807);
xor U6235 (N_6235,N_4909,N_3501);
nand U6236 (N_6236,N_3643,N_3403);
nand U6237 (N_6237,N_4487,N_3041);
and U6238 (N_6238,N_4525,N_2515);
and U6239 (N_6239,N_2879,N_3664);
or U6240 (N_6240,N_4211,N_3109);
nor U6241 (N_6241,N_3726,N_3241);
nor U6242 (N_6242,N_4656,N_3092);
nand U6243 (N_6243,N_2562,N_4701);
or U6244 (N_6244,N_2578,N_2902);
and U6245 (N_6245,N_4216,N_3234);
nor U6246 (N_6246,N_3371,N_4383);
nand U6247 (N_6247,N_3693,N_4652);
nor U6248 (N_6248,N_3560,N_2777);
nand U6249 (N_6249,N_4703,N_2754);
nand U6250 (N_6250,N_2792,N_3597);
nand U6251 (N_6251,N_4739,N_2905);
or U6252 (N_6252,N_4403,N_2682);
nor U6253 (N_6253,N_3197,N_4773);
nor U6254 (N_6254,N_3245,N_3423);
xor U6255 (N_6255,N_4543,N_3373);
xor U6256 (N_6256,N_2937,N_4030);
and U6257 (N_6257,N_3778,N_3943);
and U6258 (N_6258,N_4940,N_4884);
and U6259 (N_6259,N_4297,N_4134);
or U6260 (N_6260,N_2971,N_4189);
xor U6261 (N_6261,N_3054,N_3601);
nand U6262 (N_6262,N_4770,N_2752);
xnor U6263 (N_6263,N_3680,N_4468);
and U6264 (N_6264,N_4141,N_3069);
or U6265 (N_6265,N_4449,N_2632);
xor U6266 (N_6266,N_2931,N_2627);
xnor U6267 (N_6267,N_3709,N_4421);
and U6268 (N_6268,N_4682,N_4769);
nor U6269 (N_6269,N_3660,N_2868);
nor U6270 (N_6270,N_2775,N_2846);
nand U6271 (N_6271,N_3469,N_3597);
or U6272 (N_6272,N_2927,N_4679);
nor U6273 (N_6273,N_4542,N_4573);
and U6274 (N_6274,N_3948,N_3321);
nor U6275 (N_6275,N_3177,N_4574);
or U6276 (N_6276,N_4574,N_3968);
nand U6277 (N_6277,N_4656,N_3037);
nand U6278 (N_6278,N_4142,N_4784);
and U6279 (N_6279,N_3979,N_2537);
nor U6280 (N_6280,N_3379,N_2581);
or U6281 (N_6281,N_3744,N_3431);
nor U6282 (N_6282,N_3704,N_3991);
nand U6283 (N_6283,N_3115,N_4231);
and U6284 (N_6284,N_3732,N_3041);
nand U6285 (N_6285,N_3851,N_4281);
and U6286 (N_6286,N_4644,N_3079);
and U6287 (N_6287,N_2658,N_3775);
or U6288 (N_6288,N_3441,N_4023);
xor U6289 (N_6289,N_2591,N_4507);
nor U6290 (N_6290,N_3698,N_2872);
xor U6291 (N_6291,N_3933,N_4837);
and U6292 (N_6292,N_3777,N_4774);
xor U6293 (N_6293,N_3528,N_3919);
nand U6294 (N_6294,N_3913,N_3741);
and U6295 (N_6295,N_3706,N_4351);
xnor U6296 (N_6296,N_4520,N_3415);
nor U6297 (N_6297,N_3541,N_4493);
nand U6298 (N_6298,N_3670,N_3908);
or U6299 (N_6299,N_3810,N_4064);
or U6300 (N_6300,N_3666,N_4796);
nor U6301 (N_6301,N_2791,N_4444);
or U6302 (N_6302,N_3556,N_4481);
nand U6303 (N_6303,N_2743,N_3070);
or U6304 (N_6304,N_4480,N_4774);
nor U6305 (N_6305,N_4004,N_2949);
nor U6306 (N_6306,N_3318,N_4365);
and U6307 (N_6307,N_2722,N_4443);
and U6308 (N_6308,N_3980,N_3548);
xor U6309 (N_6309,N_4753,N_3039);
nor U6310 (N_6310,N_4799,N_3809);
or U6311 (N_6311,N_3034,N_4980);
or U6312 (N_6312,N_2636,N_3595);
nand U6313 (N_6313,N_3375,N_4040);
nand U6314 (N_6314,N_4199,N_2717);
or U6315 (N_6315,N_3987,N_3599);
nor U6316 (N_6316,N_4698,N_4330);
xnor U6317 (N_6317,N_4916,N_4113);
and U6318 (N_6318,N_4047,N_2768);
or U6319 (N_6319,N_4253,N_4230);
and U6320 (N_6320,N_2856,N_2816);
and U6321 (N_6321,N_2738,N_4604);
or U6322 (N_6322,N_4078,N_4086);
nor U6323 (N_6323,N_2961,N_2766);
or U6324 (N_6324,N_4185,N_4271);
nand U6325 (N_6325,N_2644,N_2955);
and U6326 (N_6326,N_2962,N_3666);
xor U6327 (N_6327,N_3965,N_2668);
nand U6328 (N_6328,N_4292,N_4648);
xnor U6329 (N_6329,N_3189,N_2742);
xnor U6330 (N_6330,N_4920,N_3424);
nand U6331 (N_6331,N_4504,N_3114);
nand U6332 (N_6332,N_3315,N_2752);
nor U6333 (N_6333,N_4017,N_3644);
and U6334 (N_6334,N_4710,N_3136);
or U6335 (N_6335,N_3158,N_4089);
or U6336 (N_6336,N_3748,N_3208);
and U6337 (N_6337,N_2558,N_4888);
xnor U6338 (N_6338,N_3944,N_2682);
and U6339 (N_6339,N_4516,N_2851);
nand U6340 (N_6340,N_2603,N_3463);
and U6341 (N_6341,N_4308,N_4300);
xnor U6342 (N_6342,N_4463,N_4983);
and U6343 (N_6343,N_3703,N_4810);
or U6344 (N_6344,N_3824,N_3755);
and U6345 (N_6345,N_3459,N_4119);
or U6346 (N_6346,N_3946,N_4808);
nor U6347 (N_6347,N_3280,N_3063);
nand U6348 (N_6348,N_2519,N_2617);
nor U6349 (N_6349,N_4777,N_4820);
nor U6350 (N_6350,N_3167,N_3638);
xnor U6351 (N_6351,N_2947,N_4768);
nor U6352 (N_6352,N_3752,N_3432);
xor U6353 (N_6353,N_4778,N_2645);
nand U6354 (N_6354,N_3895,N_3410);
xnor U6355 (N_6355,N_2693,N_3371);
nor U6356 (N_6356,N_4434,N_3694);
and U6357 (N_6357,N_3104,N_2512);
nor U6358 (N_6358,N_3390,N_4937);
nor U6359 (N_6359,N_2852,N_2666);
or U6360 (N_6360,N_3580,N_4395);
and U6361 (N_6361,N_3092,N_3830);
xor U6362 (N_6362,N_4564,N_3179);
or U6363 (N_6363,N_4427,N_2983);
nand U6364 (N_6364,N_4406,N_4784);
and U6365 (N_6365,N_4408,N_4711);
xor U6366 (N_6366,N_3541,N_4359);
or U6367 (N_6367,N_3152,N_3814);
and U6368 (N_6368,N_2605,N_4394);
nor U6369 (N_6369,N_4398,N_3375);
nor U6370 (N_6370,N_3057,N_3959);
and U6371 (N_6371,N_2678,N_2559);
nand U6372 (N_6372,N_3337,N_4964);
nor U6373 (N_6373,N_2792,N_4428);
nand U6374 (N_6374,N_4394,N_4921);
xor U6375 (N_6375,N_4248,N_3674);
xor U6376 (N_6376,N_4846,N_2740);
and U6377 (N_6377,N_3485,N_3526);
xor U6378 (N_6378,N_2520,N_2898);
and U6379 (N_6379,N_4368,N_4690);
xor U6380 (N_6380,N_4864,N_4520);
nand U6381 (N_6381,N_4463,N_4750);
nor U6382 (N_6382,N_4851,N_3218);
and U6383 (N_6383,N_4297,N_3445);
nor U6384 (N_6384,N_3836,N_2665);
xor U6385 (N_6385,N_4158,N_3722);
xnor U6386 (N_6386,N_4000,N_3654);
xor U6387 (N_6387,N_3031,N_2678);
xnor U6388 (N_6388,N_2978,N_2968);
nor U6389 (N_6389,N_2822,N_2724);
nor U6390 (N_6390,N_3675,N_3834);
or U6391 (N_6391,N_2997,N_4120);
xnor U6392 (N_6392,N_3578,N_3944);
nor U6393 (N_6393,N_4795,N_3738);
nand U6394 (N_6394,N_2667,N_4237);
nand U6395 (N_6395,N_4272,N_4239);
nor U6396 (N_6396,N_4834,N_3512);
xor U6397 (N_6397,N_3975,N_4178);
nor U6398 (N_6398,N_4249,N_3354);
or U6399 (N_6399,N_4840,N_4282);
nand U6400 (N_6400,N_3534,N_3902);
nand U6401 (N_6401,N_2530,N_3400);
nor U6402 (N_6402,N_3496,N_4438);
and U6403 (N_6403,N_2959,N_2746);
nand U6404 (N_6404,N_3799,N_4111);
nand U6405 (N_6405,N_3679,N_3777);
nor U6406 (N_6406,N_2539,N_3439);
and U6407 (N_6407,N_2869,N_2645);
and U6408 (N_6408,N_4147,N_3243);
nand U6409 (N_6409,N_2821,N_2946);
nor U6410 (N_6410,N_4319,N_3144);
and U6411 (N_6411,N_3111,N_2535);
xor U6412 (N_6412,N_4758,N_4840);
nand U6413 (N_6413,N_4164,N_4306);
nand U6414 (N_6414,N_4047,N_2844);
or U6415 (N_6415,N_2533,N_3466);
nand U6416 (N_6416,N_4232,N_4270);
nor U6417 (N_6417,N_2873,N_4576);
nor U6418 (N_6418,N_4172,N_3762);
nand U6419 (N_6419,N_3273,N_2652);
xnor U6420 (N_6420,N_2559,N_3363);
nand U6421 (N_6421,N_2602,N_4243);
or U6422 (N_6422,N_4582,N_3865);
xnor U6423 (N_6423,N_3166,N_4967);
or U6424 (N_6424,N_3628,N_3131);
nand U6425 (N_6425,N_3103,N_4018);
and U6426 (N_6426,N_2789,N_3799);
nor U6427 (N_6427,N_3729,N_4830);
nor U6428 (N_6428,N_3687,N_2540);
xnor U6429 (N_6429,N_4644,N_3397);
xor U6430 (N_6430,N_3674,N_3555);
or U6431 (N_6431,N_2923,N_3971);
xor U6432 (N_6432,N_3466,N_4015);
nor U6433 (N_6433,N_3848,N_2862);
xnor U6434 (N_6434,N_2741,N_3462);
nor U6435 (N_6435,N_4810,N_3784);
nor U6436 (N_6436,N_4103,N_2524);
and U6437 (N_6437,N_3494,N_3351);
xor U6438 (N_6438,N_4193,N_3393);
xnor U6439 (N_6439,N_4712,N_3721);
nand U6440 (N_6440,N_3578,N_2906);
xor U6441 (N_6441,N_4626,N_4132);
nor U6442 (N_6442,N_3897,N_3204);
xnor U6443 (N_6443,N_2582,N_3457);
xor U6444 (N_6444,N_2666,N_4741);
nand U6445 (N_6445,N_2713,N_3443);
nand U6446 (N_6446,N_3460,N_2801);
and U6447 (N_6447,N_3381,N_2718);
nor U6448 (N_6448,N_4287,N_3359);
and U6449 (N_6449,N_4042,N_3926);
or U6450 (N_6450,N_3269,N_4430);
nor U6451 (N_6451,N_2597,N_2980);
nand U6452 (N_6452,N_4154,N_2989);
nand U6453 (N_6453,N_2609,N_4314);
xnor U6454 (N_6454,N_4315,N_4300);
nand U6455 (N_6455,N_4253,N_3148);
xnor U6456 (N_6456,N_3893,N_4753);
nand U6457 (N_6457,N_3550,N_3007);
nor U6458 (N_6458,N_4923,N_3981);
xor U6459 (N_6459,N_3427,N_4279);
nor U6460 (N_6460,N_4095,N_4549);
xnor U6461 (N_6461,N_3422,N_4057);
xor U6462 (N_6462,N_2691,N_4452);
and U6463 (N_6463,N_4748,N_3071);
nand U6464 (N_6464,N_4648,N_3029);
or U6465 (N_6465,N_4517,N_3936);
nand U6466 (N_6466,N_4037,N_4040);
or U6467 (N_6467,N_4954,N_3919);
or U6468 (N_6468,N_4329,N_2852);
xor U6469 (N_6469,N_3209,N_2788);
nor U6470 (N_6470,N_3569,N_4814);
and U6471 (N_6471,N_3251,N_4606);
or U6472 (N_6472,N_3077,N_4892);
nand U6473 (N_6473,N_4382,N_2847);
nor U6474 (N_6474,N_2966,N_4606);
xor U6475 (N_6475,N_2937,N_4552);
and U6476 (N_6476,N_3841,N_3144);
or U6477 (N_6477,N_3431,N_2906);
or U6478 (N_6478,N_4155,N_4364);
nand U6479 (N_6479,N_4553,N_4021);
xnor U6480 (N_6480,N_3802,N_3696);
xor U6481 (N_6481,N_2500,N_4788);
or U6482 (N_6482,N_3412,N_3051);
nand U6483 (N_6483,N_4822,N_3845);
xor U6484 (N_6484,N_2836,N_2939);
nand U6485 (N_6485,N_4344,N_2937);
and U6486 (N_6486,N_4579,N_2555);
nor U6487 (N_6487,N_4634,N_4772);
nor U6488 (N_6488,N_2512,N_3297);
nor U6489 (N_6489,N_3294,N_2697);
xnor U6490 (N_6490,N_2914,N_3384);
and U6491 (N_6491,N_3027,N_2546);
nand U6492 (N_6492,N_3984,N_4929);
nand U6493 (N_6493,N_3853,N_3034);
nand U6494 (N_6494,N_3672,N_4237);
and U6495 (N_6495,N_3634,N_2576);
nor U6496 (N_6496,N_3330,N_2956);
and U6497 (N_6497,N_4070,N_2591);
xor U6498 (N_6498,N_4996,N_3305);
and U6499 (N_6499,N_2810,N_3891);
xor U6500 (N_6500,N_3422,N_2725);
nand U6501 (N_6501,N_2971,N_3868);
or U6502 (N_6502,N_2677,N_3574);
xor U6503 (N_6503,N_3538,N_3892);
xnor U6504 (N_6504,N_3669,N_3678);
xor U6505 (N_6505,N_4932,N_2871);
and U6506 (N_6506,N_3543,N_2845);
or U6507 (N_6507,N_3058,N_3457);
nor U6508 (N_6508,N_4646,N_2783);
nor U6509 (N_6509,N_3435,N_3677);
and U6510 (N_6510,N_3758,N_4132);
nor U6511 (N_6511,N_4020,N_4481);
nor U6512 (N_6512,N_4560,N_2569);
or U6513 (N_6513,N_3768,N_4618);
and U6514 (N_6514,N_4326,N_2641);
nand U6515 (N_6515,N_3201,N_2774);
nand U6516 (N_6516,N_4692,N_3894);
nand U6517 (N_6517,N_4047,N_3340);
or U6518 (N_6518,N_4118,N_4151);
nand U6519 (N_6519,N_3421,N_3956);
or U6520 (N_6520,N_4202,N_4438);
and U6521 (N_6521,N_3912,N_4064);
or U6522 (N_6522,N_3501,N_4822);
and U6523 (N_6523,N_3733,N_3765);
nor U6524 (N_6524,N_3204,N_4824);
or U6525 (N_6525,N_2927,N_2648);
or U6526 (N_6526,N_2561,N_2774);
xor U6527 (N_6527,N_4239,N_2734);
xor U6528 (N_6528,N_4452,N_3106);
nand U6529 (N_6529,N_4628,N_4293);
nand U6530 (N_6530,N_3166,N_3246);
nand U6531 (N_6531,N_4275,N_2894);
or U6532 (N_6532,N_3434,N_3605);
nor U6533 (N_6533,N_4351,N_4781);
nand U6534 (N_6534,N_3463,N_3893);
or U6535 (N_6535,N_3713,N_2936);
nand U6536 (N_6536,N_4403,N_3393);
xnor U6537 (N_6537,N_2989,N_4584);
or U6538 (N_6538,N_3413,N_4343);
and U6539 (N_6539,N_4999,N_3856);
and U6540 (N_6540,N_2630,N_3775);
nor U6541 (N_6541,N_4981,N_3023);
xnor U6542 (N_6542,N_4448,N_3571);
nor U6543 (N_6543,N_4718,N_3665);
xnor U6544 (N_6544,N_4448,N_3266);
or U6545 (N_6545,N_2926,N_2900);
xnor U6546 (N_6546,N_3739,N_3535);
or U6547 (N_6547,N_4124,N_2751);
nor U6548 (N_6548,N_2770,N_2551);
xor U6549 (N_6549,N_3228,N_4000);
or U6550 (N_6550,N_2738,N_3145);
nand U6551 (N_6551,N_3552,N_4973);
xnor U6552 (N_6552,N_2780,N_4411);
nand U6553 (N_6553,N_2506,N_2539);
nand U6554 (N_6554,N_3138,N_3568);
nor U6555 (N_6555,N_4703,N_2918);
or U6556 (N_6556,N_3541,N_3380);
or U6557 (N_6557,N_2634,N_3595);
xor U6558 (N_6558,N_3856,N_2629);
nand U6559 (N_6559,N_2631,N_4995);
nand U6560 (N_6560,N_4553,N_4283);
or U6561 (N_6561,N_4327,N_4259);
nor U6562 (N_6562,N_4370,N_2810);
xnor U6563 (N_6563,N_4419,N_3931);
xnor U6564 (N_6564,N_4830,N_4210);
and U6565 (N_6565,N_4067,N_4788);
nand U6566 (N_6566,N_4891,N_3111);
nor U6567 (N_6567,N_3529,N_3437);
nor U6568 (N_6568,N_3967,N_4091);
or U6569 (N_6569,N_3690,N_3253);
xnor U6570 (N_6570,N_2653,N_4504);
nand U6571 (N_6571,N_4775,N_3258);
and U6572 (N_6572,N_4474,N_4403);
xnor U6573 (N_6573,N_3623,N_2500);
xor U6574 (N_6574,N_3265,N_4065);
nor U6575 (N_6575,N_4095,N_3694);
nand U6576 (N_6576,N_2824,N_4132);
xor U6577 (N_6577,N_3796,N_3990);
and U6578 (N_6578,N_2547,N_2926);
nor U6579 (N_6579,N_2516,N_4027);
nand U6580 (N_6580,N_2822,N_4560);
nor U6581 (N_6581,N_2858,N_2574);
nor U6582 (N_6582,N_4443,N_4600);
nor U6583 (N_6583,N_4991,N_4655);
nor U6584 (N_6584,N_4669,N_3523);
and U6585 (N_6585,N_4451,N_3647);
nand U6586 (N_6586,N_2884,N_4122);
nand U6587 (N_6587,N_4825,N_3609);
xor U6588 (N_6588,N_4572,N_4611);
nand U6589 (N_6589,N_3437,N_4460);
nand U6590 (N_6590,N_4589,N_4253);
and U6591 (N_6591,N_4750,N_3441);
xnor U6592 (N_6592,N_2600,N_4332);
xor U6593 (N_6593,N_4756,N_3179);
nor U6594 (N_6594,N_4152,N_4452);
nand U6595 (N_6595,N_2606,N_2967);
nor U6596 (N_6596,N_2990,N_2828);
or U6597 (N_6597,N_2809,N_4822);
nand U6598 (N_6598,N_4474,N_2546);
xor U6599 (N_6599,N_4419,N_3422);
nand U6600 (N_6600,N_2509,N_3598);
nand U6601 (N_6601,N_3352,N_2799);
xor U6602 (N_6602,N_3329,N_2509);
xor U6603 (N_6603,N_3397,N_3055);
nand U6604 (N_6604,N_3964,N_3175);
nor U6605 (N_6605,N_2943,N_3071);
xnor U6606 (N_6606,N_2501,N_3592);
or U6607 (N_6607,N_3660,N_3035);
xor U6608 (N_6608,N_3947,N_4388);
xnor U6609 (N_6609,N_4003,N_4558);
and U6610 (N_6610,N_2822,N_2786);
or U6611 (N_6611,N_2520,N_3382);
nor U6612 (N_6612,N_3345,N_4298);
or U6613 (N_6613,N_4860,N_3665);
nand U6614 (N_6614,N_3693,N_4712);
and U6615 (N_6615,N_3577,N_3614);
and U6616 (N_6616,N_3570,N_3983);
nand U6617 (N_6617,N_4824,N_4160);
and U6618 (N_6618,N_3901,N_3508);
xnor U6619 (N_6619,N_3000,N_4345);
and U6620 (N_6620,N_4675,N_2965);
nor U6621 (N_6621,N_4539,N_4787);
xor U6622 (N_6622,N_2579,N_3914);
and U6623 (N_6623,N_4355,N_4860);
or U6624 (N_6624,N_4500,N_2728);
xnor U6625 (N_6625,N_2511,N_4003);
and U6626 (N_6626,N_4156,N_2702);
nor U6627 (N_6627,N_4947,N_2683);
nor U6628 (N_6628,N_3755,N_4418);
xnor U6629 (N_6629,N_2701,N_2588);
nand U6630 (N_6630,N_2666,N_3743);
nand U6631 (N_6631,N_3270,N_4189);
nor U6632 (N_6632,N_3949,N_3248);
and U6633 (N_6633,N_3036,N_4074);
or U6634 (N_6634,N_4532,N_4124);
and U6635 (N_6635,N_3999,N_2872);
and U6636 (N_6636,N_3961,N_4723);
and U6637 (N_6637,N_3912,N_2834);
and U6638 (N_6638,N_3366,N_4442);
and U6639 (N_6639,N_2895,N_4975);
or U6640 (N_6640,N_3644,N_3365);
nand U6641 (N_6641,N_3109,N_3425);
or U6642 (N_6642,N_3923,N_2777);
nand U6643 (N_6643,N_3549,N_4717);
or U6644 (N_6644,N_2621,N_3662);
xor U6645 (N_6645,N_3356,N_3160);
xor U6646 (N_6646,N_2684,N_2569);
xor U6647 (N_6647,N_4927,N_4664);
nor U6648 (N_6648,N_3332,N_4736);
xnor U6649 (N_6649,N_2618,N_2843);
nand U6650 (N_6650,N_2681,N_3750);
nand U6651 (N_6651,N_3354,N_3823);
nand U6652 (N_6652,N_4351,N_4992);
nand U6653 (N_6653,N_2631,N_3807);
xor U6654 (N_6654,N_4855,N_3224);
xor U6655 (N_6655,N_2641,N_4320);
or U6656 (N_6656,N_2510,N_4708);
and U6657 (N_6657,N_3272,N_3589);
xor U6658 (N_6658,N_4759,N_4496);
nand U6659 (N_6659,N_4999,N_4527);
or U6660 (N_6660,N_2967,N_3090);
xnor U6661 (N_6661,N_3023,N_3824);
nor U6662 (N_6662,N_4602,N_2648);
nor U6663 (N_6663,N_2893,N_3059);
nand U6664 (N_6664,N_4918,N_4205);
xor U6665 (N_6665,N_2765,N_3415);
nand U6666 (N_6666,N_2915,N_2826);
nor U6667 (N_6667,N_4722,N_4252);
nor U6668 (N_6668,N_2820,N_3160);
nand U6669 (N_6669,N_3187,N_4065);
or U6670 (N_6670,N_3629,N_2909);
nor U6671 (N_6671,N_2550,N_3103);
xnor U6672 (N_6672,N_3986,N_3761);
xor U6673 (N_6673,N_3930,N_2919);
and U6674 (N_6674,N_3559,N_4001);
xor U6675 (N_6675,N_4337,N_4211);
nor U6676 (N_6676,N_4775,N_3541);
or U6677 (N_6677,N_4407,N_4332);
and U6678 (N_6678,N_4697,N_4611);
xor U6679 (N_6679,N_3666,N_4585);
nand U6680 (N_6680,N_4093,N_2615);
or U6681 (N_6681,N_4626,N_4013);
nor U6682 (N_6682,N_3280,N_4964);
nand U6683 (N_6683,N_3156,N_4327);
and U6684 (N_6684,N_4948,N_3105);
nand U6685 (N_6685,N_3483,N_4582);
nand U6686 (N_6686,N_3485,N_4110);
xor U6687 (N_6687,N_2865,N_2707);
and U6688 (N_6688,N_2731,N_2592);
and U6689 (N_6689,N_4330,N_2926);
nor U6690 (N_6690,N_4527,N_3064);
and U6691 (N_6691,N_3379,N_4772);
or U6692 (N_6692,N_4899,N_4138);
or U6693 (N_6693,N_2912,N_3007);
nor U6694 (N_6694,N_4501,N_4834);
and U6695 (N_6695,N_3650,N_4564);
or U6696 (N_6696,N_4980,N_3012);
nand U6697 (N_6697,N_3850,N_4095);
or U6698 (N_6698,N_2834,N_3993);
nor U6699 (N_6699,N_4784,N_3169);
and U6700 (N_6700,N_3060,N_3601);
nand U6701 (N_6701,N_3202,N_4883);
and U6702 (N_6702,N_3609,N_3932);
or U6703 (N_6703,N_4264,N_3529);
nand U6704 (N_6704,N_2563,N_4451);
and U6705 (N_6705,N_2825,N_3714);
or U6706 (N_6706,N_4737,N_4175);
xor U6707 (N_6707,N_3419,N_4122);
nor U6708 (N_6708,N_2965,N_2746);
or U6709 (N_6709,N_2592,N_4004);
nor U6710 (N_6710,N_3973,N_3654);
nor U6711 (N_6711,N_4909,N_4240);
nand U6712 (N_6712,N_4034,N_4644);
and U6713 (N_6713,N_4927,N_3418);
or U6714 (N_6714,N_3970,N_4564);
nand U6715 (N_6715,N_2777,N_3636);
nand U6716 (N_6716,N_4934,N_3076);
and U6717 (N_6717,N_3780,N_4303);
xnor U6718 (N_6718,N_3128,N_3847);
and U6719 (N_6719,N_2613,N_4152);
xnor U6720 (N_6720,N_4051,N_2675);
or U6721 (N_6721,N_2732,N_2552);
xor U6722 (N_6722,N_2688,N_3504);
and U6723 (N_6723,N_2501,N_4819);
and U6724 (N_6724,N_4612,N_4367);
xnor U6725 (N_6725,N_4865,N_2837);
xor U6726 (N_6726,N_4829,N_4878);
nand U6727 (N_6727,N_3812,N_4142);
or U6728 (N_6728,N_4613,N_3872);
nand U6729 (N_6729,N_2798,N_4882);
or U6730 (N_6730,N_2976,N_4069);
or U6731 (N_6731,N_4100,N_2586);
nand U6732 (N_6732,N_4053,N_3215);
or U6733 (N_6733,N_2750,N_3344);
xnor U6734 (N_6734,N_4843,N_3962);
or U6735 (N_6735,N_3760,N_2887);
or U6736 (N_6736,N_4670,N_4866);
or U6737 (N_6737,N_2930,N_3960);
or U6738 (N_6738,N_4082,N_2907);
or U6739 (N_6739,N_4305,N_3782);
nor U6740 (N_6740,N_4172,N_4843);
nand U6741 (N_6741,N_4387,N_4042);
xor U6742 (N_6742,N_4819,N_3286);
nor U6743 (N_6743,N_4260,N_2916);
or U6744 (N_6744,N_4472,N_4568);
xnor U6745 (N_6745,N_4383,N_2749);
nor U6746 (N_6746,N_2596,N_3957);
nor U6747 (N_6747,N_4242,N_3510);
or U6748 (N_6748,N_2641,N_3138);
xnor U6749 (N_6749,N_4245,N_3376);
nand U6750 (N_6750,N_3483,N_4130);
xor U6751 (N_6751,N_3052,N_4853);
or U6752 (N_6752,N_4002,N_4288);
xor U6753 (N_6753,N_4638,N_3336);
xnor U6754 (N_6754,N_4941,N_4097);
and U6755 (N_6755,N_4268,N_3394);
nand U6756 (N_6756,N_4665,N_4701);
and U6757 (N_6757,N_4138,N_4624);
xor U6758 (N_6758,N_3898,N_3324);
nor U6759 (N_6759,N_2561,N_2593);
xor U6760 (N_6760,N_3300,N_3859);
or U6761 (N_6761,N_3123,N_2588);
and U6762 (N_6762,N_4828,N_3297);
xnor U6763 (N_6763,N_3248,N_3018);
nor U6764 (N_6764,N_3260,N_4628);
xor U6765 (N_6765,N_4308,N_3694);
or U6766 (N_6766,N_3114,N_4190);
xnor U6767 (N_6767,N_4009,N_3219);
xor U6768 (N_6768,N_4537,N_3477);
nor U6769 (N_6769,N_4969,N_2728);
nor U6770 (N_6770,N_2646,N_4302);
and U6771 (N_6771,N_2503,N_3372);
or U6772 (N_6772,N_2577,N_4903);
xor U6773 (N_6773,N_4304,N_3927);
or U6774 (N_6774,N_3550,N_4451);
and U6775 (N_6775,N_2666,N_3862);
or U6776 (N_6776,N_4087,N_2877);
xor U6777 (N_6777,N_2767,N_3743);
or U6778 (N_6778,N_3824,N_3694);
or U6779 (N_6779,N_4346,N_4904);
or U6780 (N_6780,N_4956,N_2944);
nor U6781 (N_6781,N_2719,N_4014);
nand U6782 (N_6782,N_4716,N_3799);
or U6783 (N_6783,N_2766,N_4009);
and U6784 (N_6784,N_4208,N_3610);
or U6785 (N_6785,N_3348,N_2785);
nor U6786 (N_6786,N_3294,N_2663);
nor U6787 (N_6787,N_3136,N_4255);
nand U6788 (N_6788,N_4348,N_4810);
and U6789 (N_6789,N_4039,N_4023);
nor U6790 (N_6790,N_2586,N_2647);
nor U6791 (N_6791,N_3538,N_4942);
and U6792 (N_6792,N_2626,N_2670);
or U6793 (N_6793,N_3386,N_2695);
nor U6794 (N_6794,N_4076,N_4584);
or U6795 (N_6795,N_4121,N_2527);
or U6796 (N_6796,N_4236,N_3819);
nand U6797 (N_6797,N_3655,N_3539);
or U6798 (N_6798,N_4040,N_3999);
or U6799 (N_6799,N_4922,N_4862);
xor U6800 (N_6800,N_3255,N_4122);
xnor U6801 (N_6801,N_4539,N_4567);
and U6802 (N_6802,N_4721,N_3631);
and U6803 (N_6803,N_2876,N_3078);
xnor U6804 (N_6804,N_4758,N_4216);
xor U6805 (N_6805,N_3607,N_3873);
nand U6806 (N_6806,N_3354,N_3530);
or U6807 (N_6807,N_4107,N_2914);
xor U6808 (N_6808,N_3926,N_4773);
and U6809 (N_6809,N_2500,N_3972);
and U6810 (N_6810,N_3267,N_3019);
xor U6811 (N_6811,N_4405,N_4655);
nor U6812 (N_6812,N_4731,N_3788);
xor U6813 (N_6813,N_3394,N_2683);
nand U6814 (N_6814,N_4603,N_4756);
nand U6815 (N_6815,N_2821,N_3184);
or U6816 (N_6816,N_3661,N_3045);
nor U6817 (N_6817,N_3150,N_3272);
nand U6818 (N_6818,N_4666,N_4708);
or U6819 (N_6819,N_2505,N_3853);
and U6820 (N_6820,N_2891,N_4809);
nand U6821 (N_6821,N_2571,N_3334);
and U6822 (N_6822,N_4771,N_4132);
nor U6823 (N_6823,N_3544,N_3863);
xor U6824 (N_6824,N_3073,N_3997);
xnor U6825 (N_6825,N_3097,N_2514);
xor U6826 (N_6826,N_3402,N_3740);
nor U6827 (N_6827,N_4713,N_3915);
xor U6828 (N_6828,N_3444,N_4664);
xnor U6829 (N_6829,N_2837,N_3092);
and U6830 (N_6830,N_4616,N_4253);
xor U6831 (N_6831,N_2985,N_3011);
nand U6832 (N_6832,N_3336,N_2837);
and U6833 (N_6833,N_3950,N_3319);
nand U6834 (N_6834,N_3007,N_4451);
xnor U6835 (N_6835,N_4151,N_4378);
and U6836 (N_6836,N_4106,N_3298);
nor U6837 (N_6837,N_2575,N_4889);
nor U6838 (N_6838,N_4218,N_2935);
or U6839 (N_6839,N_2794,N_4718);
and U6840 (N_6840,N_4663,N_4216);
xnor U6841 (N_6841,N_2838,N_3150);
and U6842 (N_6842,N_4619,N_4049);
and U6843 (N_6843,N_4257,N_3930);
or U6844 (N_6844,N_3107,N_4588);
xnor U6845 (N_6845,N_3716,N_3398);
nand U6846 (N_6846,N_3065,N_4880);
nor U6847 (N_6847,N_4798,N_3156);
xnor U6848 (N_6848,N_3984,N_4359);
nor U6849 (N_6849,N_3892,N_3962);
or U6850 (N_6850,N_3064,N_3492);
xor U6851 (N_6851,N_4967,N_3194);
nand U6852 (N_6852,N_4214,N_3298);
nand U6853 (N_6853,N_3603,N_2746);
or U6854 (N_6854,N_2730,N_3349);
nand U6855 (N_6855,N_4224,N_3039);
or U6856 (N_6856,N_4819,N_3403);
nor U6857 (N_6857,N_2526,N_3641);
nor U6858 (N_6858,N_4069,N_3492);
nand U6859 (N_6859,N_4179,N_4028);
nand U6860 (N_6860,N_2904,N_4983);
or U6861 (N_6861,N_2677,N_4205);
and U6862 (N_6862,N_3947,N_4485);
nand U6863 (N_6863,N_4492,N_3497);
or U6864 (N_6864,N_4075,N_4220);
or U6865 (N_6865,N_3464,N_4911);
or U6866 (N_6866,N_4270,N_4915);
xnor U6867 (N_6867,N_3786,N_3972);
nor U6868 (N_6868,N_3790,N_4472);
xnor U6869 (N_6869,N_3739,N_4937);
and U6870 (N_6870,N_4123,N_4161);
nand U6871 (N_6871,N_3681,N_3685);
nor U6872 (N_6872,N_2612,N_3629);
or U6873 (N_6873,N_3429,N_2567);
nor U6874 (N_6874,N_2634,N_4434);
nand U6875 (N_6875,N_4510,N_4304);
nand U6876 (N_6876,N_4151,N_4204);
nand U6877 (N_6877,N_2897,N_3825);
nor U6878 (N_6878,N_3082,N_4601);
nor U6879 (N_6879,N_4630,N_2683);
nor U6880 (N_6880,N_4675,N_4820);
and U6881 (N_6881,N_4144,N_2631);
xnor U6882 (N_6882,N_4291,N_4855);
or U6883 (N_6883,N_4040,N_4123);
xnor U6884 (N_6884,N_4322,N_3245);
nor U6885 (N_6885,N_2536,N_4231);
and U6886 (N_6886,N_3119,N_4899);
or U6887 (N_6887,N_4462,N_3758);
xor U6888 (N_6888,N_4630,N_4742);
nor U6889 (N_6889,N_4300,N_2672);
nand U6890 (N_6890,N_3489,N_3805);
and U6891 (N_6891,N_3124,N_3521);
xor U6892 (N_6892,N_4601,N_4792);
nor U6893 (N_6893,N_2912,N_3075);
or U6894 (N_6894,N_4884,N_4336);
or U6895 (N_6895,N_4627,N_4475);
nor U6896 (N_6896,N_2887,N_4628);
xor U6897 (N_6897,N_2594,N_4641);
nand U6898 (N_6898,N_2860,N_4273);
and U6899 (N_6899,N_2841,N_4613);
and U6900 (N_6900,N_2549,N_4113);
or U6901 (N_6901,N_4656,N_3193);
or U6902 (N_6902,N_4598,N_3813);
xor U6903 (N_6903,N_4641,N_3787);
nor U6904 (N_6904,N_4355,N_4731);
or U6905 (N_6905,N_4603,N_3551);
or U6906 (N_6906,N_4596,N_3217);
or U6907 (N_6907,N_2536,N_4598);
and U6908 (N_6908,N_3405,N_2809);
nand U6909 (N_6909,N_2938,N_2701);
nand U6910 (N_6910,N_2521,N_2591);
nor U6911 (N_6911,N_4687,N_3809);
nor U6912 (N_6912,N_2899,N_3069);
and U6913 (N_6913,N_4030,N_4864);
and U6914 (N_6914,N_2611,N_4179);
nor U6915 (N_6915,N_3590,N_3830);
nand U6916 (N_6916,N_3524,N_3357);
and U6917 (N_6917,N_3383,N_3705);
nand U6918 (N_6918,N_4131,N_3237);
or U6919 (N_6919,N_4831,N_3034);
nor U6920 (N_6920,N_3252,N_3907);
nand U6921 (N_6921,N_2927,N_4601);
nand U6922 (N_6922,N_3853,N_4778);
nand U6923 (N_6923,N_3359,N_3287);
nand U6924 (N_6924,N_2994,N_4304);
nor U6925 (N_6925,N_4727,N_3551);
nor U6926 (N_6926,N_3819,N_2626);
nor U6927 (N_6927,N_2650,N_3762);
nand U6928 (N_6928,N_3293,N_4543);
and U6929 (N_6929,N_3801,N_4418);
nor U6930 (N_6930,N_2760,N_3970);
nand U6931 (N_6931,N_4832,N_3326);
xnor U6932 (N_6932,N_3183,N_2678);
and U6933 (N_6933,N_2801,N_4549);
nand U6934 (N_6934,N_4025,N_3714);
nand U6935 (N_6935,N_3969,N_4426);
nor U6936 (N_6936,N_3384,N_4329);
nand U6937 (N_6937,N_3526,N_4812);
and U6938 (N_6938,N_2640,N_4301);
nor U6939 (N_6939,N_3887,N_3550);
nand U6940 (N_6940,N_3224,N_4943);
and U6941 (N_6941,N_4630,N_4159);
and U6942 (N_6942,N_3223,N_3651);
xnor U6943 (N_6943,N_4623,N_4982);
nand U6944 (N_6944,N_2820,N_3220);
and U6945 (N_6945,N_4739,N_3335);
nand U6946 (N_6946,N_3460,N_4726);
xor U6947 (N_6947,N_4520,N_3020);
xor U6948 (N_6948,N_2679,N_4867);
and U6949 (N_6949,N_3062,N_4188);
nor U6950 (N_6950,N_4656,N_2501);
nand U6951 (N_6951,N_4148,N_3461);
xor U6952 (N_6952,N_3395,N_4797);
nor U6953 (N_6953,N_2826,N_2624);
xnor U6954 (N_6954,N_3760,N_4958);
and U6955 (N_6955,N_3690,N_3325);
or U6956 (N_6956,N_3723,N_3957);
or U6957 (N_6957,N_4199,N_4175);
nor U6958 (N_6958,N_4619,N_2573);
or U6959 (N_6959,N_4094,N_3567);
nand U6960 (N_6960,N_4356,N_4919);
xnor U6961 (N_6961,N_2786,N_4226);
nor U6962 (N_6962,N_3610,N_4218);
nor U6963 (N_6963,N_4297,N_3330);
or U6964 (N_6964,N_3489,N_3337);
nand U6965 (N_6965,N_4460,N_3477);
xnor U6966 (N_6966,N_2619,N_3148);
and U6967 (N_6967,N_3748,N_3378);
or U6968 (N_6968,N_2750,N_4804);
nand U6969 (N_6969,N_2791,N_4185);
nor U6970 (N_6970,N_4330,N_4507);
xor U6971 (N_6971,N_2612,N_4046);
or U6972 (N_6972,N_4596,N_3082);
or U6973 (N_6973,N_3313,N_3696);
nand U6974 (N_6974,N_4715,N_3217);
xor U6975 (N_6975,N_3955,N_3768);
xnor U6976 (N_6976,N_3562,N_4590);
nand U6977 (N_6977,N_3556,N_4132);
xnor U6978 (N_6978,N_4924,N_3697);
nand U6979 (N_6979,N_2592,N_3266);
nand U6980 (N_6980,N_3419,N_4125);
nor U6981 (N_6981,N_4921,N_2620);
or U6982 (N_6982,N_3192,N_3449);
xor U6983 (N_6983,N_4545,N_4104);
or U6984 (N_6984,N_2663,N_4578);
xor U6985 (N_6985,N_2887,N_4202);
or U6986 (N_6986,N_4206,N_3892);
nor U6987 (N_6987,N_3775,N_3334);
or U6988 (N_6988,N_4528,N_4561);
and U6989 (N_6989,N_3752,N_4819);
or U6990 (N_6990,N_4319,N_2606);
nand U6991 (N_6991,N_2858,N_4135);
nor U6992 (N_6992,N_3228,N_3648);
xnor U6993 (N_6993,N_3638,N_3746);
or U6994 (N_6994,N_3631,N_4989);
or U6995 (N_6995,N_4454,N_3642);
nand U6996 (N_6996,N_4129,N_2767);
xnor U6997 (N_6997,N_4022,N_3996);
nand U6998 (N_6998,N_3861,N_4797);
or U6999 (N_6999,N_2935,N_4802);
and U7000 (N_7000,N_2709,N_4947);
or U7001 (N_7001,N_4815,N_2944);
xor U7002 (N_7002,N_2991,N_2779);
nand U7003 (N_7003,N_4416,N_3860);
nor U7004 (N_7004,N_3515,N_4582);
or U7005 (N_7005,N_2895,N_4110);
or U7006 (N_7006,N_4861,N_2945);
nand U7007 (N_7007,N_3236,N_4827);
nand U7008 (N_7008,N_4737,N_4527);
nand U7009 (N_7009,N_2709,N_4052);
or U7010 (N_7010,N_3852,N_3399);
xnor U7011 (N_7011,N_4734,N_4700);
nand U7012 (N_7012,N_2895,N_2756);
xor U7013 (N_7013,N_3985,N_2593);
or U7014 (N_7014,N_4565,N_3264);
nor U7015 (N_7015,N_4596,N_4288);
and U7016 (N_7016,N_2532,N_3020);
nor U7017 (N_7017,N_2936,N_4389);
xnor U7018 (N_7018,N_2885,N_4041);
nor U7019 (N_7019,N_4855,N_4280);
xnor U7020 (N_7020,N_4588,N_2980);
and U7021 (N_7021,N_3330,N_4397);
and U7022 (N_7022,N_3546,N_2954);
or U7023 (N_7023,N_4464,N_4332);
nand U7024 (N_7024,N_4993,N_2724);
nor U7025 (N_7025,N_4562,N_4346);
nor U7026 (N_7026,N_3612,N_4468);
nor U7027 (N_7027,N_3908,N_2801);
nor U7028 (N_7028,N_4405,N_4444);
or U7029 (N_7029,N_3868,N_4179);
or U7030 (N_7030,N_2810,N_4292);
and U7031 (N_7031,N_3359,N_3466);
nor U7032 (N_7032,N_4645,N_2744);
or U7033 (N_7033,N_4160,N_4746);
nand U7034 (N_7034,N_4919,N_4377);
and U7035 (N_7035,N_3845,N_4757);
and U7036 (N_7036,N_2615,N_3870);
xor U7037 (N_7037,N_2555,N_2800);
nand U7038 (N_7038,N_2657,N_4198);
nand U7039 (N_7039,N_4082,N_4712);
or U7040 (N_7040,N_3918,N_4883);
and U7041 (N_7041,N_2574,N_3643);
nor U7042 (N_7042,N_3607,N_4179);
or U7043 (N_7043,N_4053,N_2951);
nor U7044 (N_7044,N_4123,N_3564);
and U7045 (N_7045,N_4898,N_3395);
and U7046 (N_7046,N_4018,N_2773);
nor U7047 (N_7047,N_4797,N_2656);
nand U7048 (N_7048,N_2695,N_2899);
and U7049 (N_7049,N_4119,N_4618);
nand U7050 (N_7050,N_4642,N_3272);
xor U7051 (N_7051,N_4844,N_4261);
nor U7052 (N_7052,N_4636,N_4783);
nor U7053 (N_7053,N_3720,N_4792);
or U7054 (N_7054,N_3836,N_3640);
or U7055 (N_7055,N_4965,N_3190);
nand U7056 (N_7056,N_4989,N_3837);
nand U7057 (N_7057,N_2561,N_4032);
nor U7058 (N_7058,N_4096,N_4093);
or U7059 (N_7059,N_4829,N_3505);
xnor U7060 (N_7060,N_3901,N_4794);
and U7061 (N_7061,N_2791,N_3792);
nand U7062 (N_7062,N_4932,N_4674);
xor U7063 (N_7063,N_3474,N_4477);
or U7064 (N_7064,N_4121,N_4639);
and U7065 (N_7065,N_2525,N_3294);
nor U7066 (N_7066,N_4118,N_3429);
xor U7067 (N_7067,N_2993,N_4811);
or U7068 (N_7068,N_3814,N_4060);
nor U7069 (N_7069,N_4125,N_3329);
nand U7070 (N_7070,N_3372,N_3659);
xnor U7071 (N_7071,N_4636,N_3369);
or U7072 (N_7072,N_3880,N_4853);
and U7073 (N_7073,N_4122,N_4628);
nand U7074 (N_7074,N_3512,N_2615);
xor U7075 (N_7075,N_3264,N_4192);
nand U7076 (N_7076,N_4410,N_2631);
xor U7077 (N_7077,N_3386,N_4603);
nand U7078 (N_7078,N_3287,N_2629);
or U7079 (N_7079,N_3671,N_2945);
or U7080 (N_7080,N_3044,N_4100);
xnor U7081 (N_7081,N_4833,N_3394);
or U7082 (N_7082,N_4195,N_2762);
nand U7083 (N_7083,N_3246,N_3984);
xnor U7084 (N_7084,N_3507,N_2939);
and U7085 (N_7085,N_3527,N_4329);
or U7086 (N_7086,N_3318,N_3380);
xor U7087 (N_7087,N_2701,N_4266);
nor U7088 (N_7088,N_2536,N_4185);
and U7089 (N_7089,N_2742,N_3178);
nand U7090 (N_7090,N_3966,N_3797);
or U7091 (N_7091,N_3615,N_3352);
xor U7092 (N_7092,N_4258,N_3597);
nand U7093 (N_7093,N_2603,N_3132);
nand U7094 (N_7094,N_4690,N_3239);
and U7095 (N_7095,N_3945,N_3735);
nand U7096 (N_7096,N_3404,N_3699);
and U7097 (N_7097,N_4120,N_3067);
and U7098 (N_7098,N_4441,N_3675);
nor U7099 (N_7099,N_3818,N_3497);
nor U7100 (N_7100,N_4951,N_2779);
nor U7101 (N_7101,N_3931,N_2718);
nand U7102 (N_7102,N_4667,N_3012);
xnor U7103 (N_7103,N_3407,N_2998);
and U7104 (N_7104,N_2928,N_4657);
or U7105 (N_7105,N_4671,N_4757);
and U7106 (N_7106,N_4404,N_4533);
nor U7107 (N_7107,N_4432,N_3361);
xnor U7108 (N_7108,N_2573,N_2950);
or U7109 (N_7109,N_4445,N_4845);
nor U7110 (N_7110,N_3634,N_3947);
and U7111 (N_7111,N_4810,N_3868);
nor U7112 (N_7112,N_2593,N_3927);
xnor U7113 (N_7113,N_4428,N_2532);
and U7114 (N_7114,N_4749,N_4247);
nand U7115 (N_7115,N_3316,N_4224);
nor U7116 (N_7116,N_4932,N_2591);
nand U7117 (N_7117,N_4720,N_4159);
xor U7118 (N_7118,N_3576,N_4060);
nor U7119 (N_7119,N_4773,N_2649);
or U7120 (N_7120,N_4480,N_3170);
or U7121 (N_7121,N_3992,N_3136);
xor U7122 (N_7122,N_3075,N_3796);
or U7123 (N_7123,N_3481,N_4178);
and U7124 (N_7124,N_3336,N_4942);
and U7125 (N_7125,N_4669,N_3735);
nand U7126 (N_7126,N_3274,N_4855);
nor U7127 (N_7127,N_4725,N_3492);
and U7128 (N_7128,N_4204,N_3742);
nand U7129 (N_7129,N_2878,N_3396);
xnor U7130 (N_7130,N_4354,N_2714);
or U7131 (N_7131,N_4822,N_3846);
xnor U7132 (N_7132,N_3360,N_3267);
nor U7133 (N_7133,N_3618,N_3908);
nor U7134 (N_7134,N_3982,N_4296);
xor U7135 (N_7135,N_3038,N_2501);
nand U7136 (N_7136,N_4880,N_2756);
xnor U7137 (N_7137,N_4022,N_3534);
and U7138 (N_7138,N_4692,N_3332);
nor U7139 (N_7139,N_2682,N_3046);
xnor U7140 (N_7140,N_4706,N_4220);
nand U7141 (N_7141,N_3568,N_2605);
or U7142 (N_7142,N_4425,N_4838);
xor U7143 (N_7143,N_3903,N_4031);
xor U7144 (N_7144,N_3527,N_2822);
nor U7145 (N_7145,N_3430,N_3279);
and U7146 (N_7146,N_4724,N_3637);
nor U7147 (N_7147,N_3934,N_2845);
xnor U7148 (N_7148,N_3079,N_4121);
nor U7149 (N_7149,N_4324,N_4884);
xnor U7150 (N_7150,N_4338,N_2836);
and U7151 (N_7151,N_3563,N_3949);
nand U7152 (N_7152,N_4416,N_3936);
nor U7153 (N_7153,N_3689,N_2842);
nor U7154 (N_7154,N_2858,N_4044);
nor U7155 (N_7155,N_2503,N_2819);
and U7156 (N_7156,N_3010,N_4248);
nand U7157 (N_7157,N_2947,N_4203);
nor U7158 (N_7158,N_4857,N_4734);
nand U7159 (N_7159,N_4376,N_4167);
nand U7160 (N_7160,N_3171,N_4502);
and U7161 (N_7161,N_2774,N_3299);
nor U7162 (N_7162,N_2911,N_3575);
nor U7163 (N_7163,N_4026,N_4241);
or U7164 (N_7164,N_3487,N_4278);
and U7165 (N_7165,N_3170,N_4159);
and U7166 (N_7166,N_2599,N_3311);
and U7167 (N_7167,N_2959,N_3939);
and U7168 (N_7168,N_4564,N_3066);
and U7169 (N_7169,N_2714,N_2982);
nand U7170 (N_7170,N_4228,N_4199);
nor U7171 (N_7171,N_4817,N_4584);
or U7172 (N_7172,N_4283,N_2708);
or U7173 (N_7173,N_3298,N_4990);
xnor U7174 (N_7174,N_4086,N_4363);
and U7175 (N_7175,N_4650,N_2847);
nand U7176 (N_7176,N_3200,N_4593);
and U7177 (N_7177,N_4358,N_4338);
xor U7178 (N_7178,N_4614,N_4928);
xor U7179 (N_7179,N_3621,N_3673);
xor U7180 (N_7180,N_2589,N_3224);
or U7181 (N_7181,N_3281,N_2898);
and U7182 (N_7182,N_4822,N_4222);
nor U7183 (N_7183,N_2734,N_3937);
nor U7184 (N_7184,N_4947,N_4968);
nor U7185 (N_7185,N_3454,N_3108);
or U7186 (N_7186,N_3228,N_4465);
nor U7187 (N_7187,N_2734,N_3371);
and U7188 (N_7188,N_3979,N_2883);
and U7189 (N_7189,N_3162,N_3726);
nor U7190 (N_7190,N_4503,N_4298);
nand U7191 (N_7191,N_3250,N_3856);
or U7192 (N_7192,N_3928,N_4516);
nand U7193 (N_7193,N_3767,N_4681);
nand U7194 (N_7194,N_4404,N_2604);
nand U7195 (N_7195,N_4301,N_2630);
xor U7196 (N_7196,N_3494,N_2761);
nor U7197 (N_7197,N_3466,N_3754);
and U7198 (N_7198,N_3358,N_4213);
or U7199 (N_7199,N_4131,N_3008);
and U7200 (N_7200,N_4999,N_3410);
nand U7201 (N_7201,N_2654,N_3448);
nand U7202 (N_7202,N_2629,N_2825);
xor U7203 (N_7203,N_2541,N_4278);
xor U7204 (N_7204,N_4917,N_4034);
xnor U7205 (N_7205,N_3798,N_4941);
and U7206 (N_7206,N_4255,N_4741);
nor U7207 (N_7207,N_2803,N_3922);
and U7208 (N_7208,N_4287,N_2908);
nor U7209 (N_7209,N_4971,N_4392);
xnor U7210 (N_7210,N_3977,N_2522);
and U7211 (N_7211,N_3543,N_2913);
or U7212 (N_7212,N_4266,N_3175);
and U7213 (N_7213,N_3001,N_2520);
xor U7214 (N_7214,N_3952,N_3494);
and U7215 (N_7215,N_4346,N_3060);
xor U7216 (N_7216,N_4608,N_4554);
or U7217 (N_7217,N_3168,N_3586);
xnor U7218 (N_7218,N_4345,N_2586);
xor U7219 (N_7219,N_4250,N_2971);
nor U7220 (N_7220,N_2748,N_4653);
or U7221 (N_7221,N_2586,N_3811);
xnor U7222 (N_7222,N_4352,N_2848);
nor U7223 (N_7223,N_2718,N_3425);
and U7224 (N_7224,N_2807,N_3831);
and U7225 (N_7225,N_4389,N_2589);
or U7226 (N_7226,N_2619,N_4376);
xnor U7227 (N_7227,N_4766,N_4420);
xor U7228 (N_7228,N_3231,N_3452);
nand U7229 (N_7229,N_4083,N_3756);
nand U7230 (N_7230,N_3632,N_3515);
nor U7231 (N_7231,N_4597,N_3382);
nand U7232 (N_7232,N_3294,N_4467);
xnor U7233 (N_7233,N_3720,N_4753);
or U7234 (N_7234,N_3711,N_4375);
nor U7235 (N_7235,N_3631,N_3595);
xor U7236 (N_7236,N_4816,N_4730);
nand U7237 (N_7237,N_3653,N_3158);
and U7238 (N_7238,N_3759,N_2579);
and U7239 (N_7239,N_3043,N_3540);
xor U7240 (N_7240,N_2850,N_4617);
or U7241 (N_7241,N_4117,N_3089);
and U7242 (N_7242,N_4670,N_4874);
and U7243 (N_7243,N_3007,N_4608);
nand U7244 (N_7244,N_3541,N_3860);
nor U7245 (N_7245,N_3782,N_3052);
or U7246 (N_7246,N_3799,N_4033);
xor U7247 (N_7247,N_3462,N_3826);
nor U7248 (N_7248,N_3443,N_2622);
nand U7249 (N_7249,N_2798,N_2584);
or U7250 (N_7250,N_3997,N_2981);
nor U7251 (N_7251,N_4056,N_4911);
nand U7252 (N_7252,N_2689,N_3439);
or U7253 (N_7253,N_4592,N_3346);
nand U7254 (N_7254,N_2579,N_4703);
or U7255 (N_7255,N_3887,N_3137);
nor U7256 (N_7256,N_2903,N_4824);
and U7257 (N_7257,N_3222,N_3621);
and U7258 (N_7258,N_4748,N_4096);
and U7259 (N_7259,N_4762,N_3789);
nor U7260 (N_7260,N_3233,N_3360);
and U7261 (N_7261,N_4896,N_3655);
nand U7262 (N_7262,N_3369,N_2960);
nor U7263 (N_7263,N_4711,N_3820);
and U7264 (N_7264,N_2850,N_3610);
nor U7265 (N_7265,N_2808,N_2835);
nand U7266 (N_7266,N_4364,N_4841);
and U7267 (N_7267,N_4012,N_3105);
or U7268 (N_7268,N_4953,N_3246);
nand U7269 (N_7269,N_4752,N_3770);
or U7270 (N_7270,N_2879,N_4498);
or U7271 (N_7271,N_3845,N_2745);
nor U7272 (N_7272,N_4947,N_3071);
or U7273 (N_7273,N_3318,N_3619);
or U7274 (N_7274,N_3299,N_2801);
xor U7275 (N_7275,N_4729,N_4102);
nor U7276 (N_7276,N_3414,N_4172);
nor U7277 (N_7277,N_2595,N_2886);
or U7278 (N_7278,N_4338,N_4248);
xor U7279 (N_7279,N_4981,N_2709);
nand U7280 (N_7280,N_3986,N_3136);
nand U7281 (N_7281,N_3400,N_4869);
nand U7282 (N_7282,N_2542,N_3961);
and U7283 (N_7283,N_3791,N_2604);
and U7284 (N_7284,N_3188,N_3634);
and U7285 (N_7285,N_3311,N_4971);
nor U7286 (N_7286,N_3654,N_4097);
xor U7287 (N_7287,N_4782,N_2964);
xnor U7288 (N_7288,N_3016,N_4069);
or U7289 (N_7289,N_3936,N_3341);
xnor U7290 (N_7290,N_4437,N_2859);
and U7291 (N_7291,N_4842,N_2746);
nor U7292 (N_7292,N_3739,N_3727);
and U7293 (N_7293,N_4034,N_4728);
and U7294 (N_7294,N_3510,N_2569);
and U7295 (N_7295,N_4849,N_4738);
nor U7296 (N_7296,N_3063,N_2815);
and U7297 (N_7297,N_4770,N_4188);
and U7298 (N_7298,N_3803,N_4391);
or U7299 (N_7299,N_2569,N_3829);
and U7300 (N_7300,N_4411,N_2597);
and U7301 (N_7301,N_3503,N_4446);
and U7302 (N_7302,N_4119,N_4017);
and U7303 (N_7303,N_4493,N_4018);
nor U7304 (N_7304,N_4440,N_4268);
and U7305 (N_7305,N_3732,N_3754);
nor U7306 (N_7306,N_2622,N_4109);
nor U7307 (N_7307,N_4659,N_3206);
or U7308 (N_7308,N_4352,N_4802);
nor U7309 (N_7309,N_3379,N_2555);
and U7310 (N_7310,N_4947,N_3123);
nor U7311 (N_7311,N_4425,N_4352);
nor U7312 (N_7312,N_3019,N_3878);
or U7313 (N_7313,N_4066,N_2829);
nand U7314 (N_7314,N_4956,N_4852);
nor U7315 (N_7315,N_4395,N_3083);
and U7316 (N_7316,N_3244,N_4208);
and U7317 (N_7317,N_3780,N_3151);
and U7318 (N_7318,N_4199,N_3515);
xnor U7319 (N_7319,N_4475,N_2616);
or U7320 (N_7320,N_4525,N_3991);
or U7321 (N_7321,N_4703,N_4808);
xnor U7322 (N_7322,N_4691,N_3242);
xor U7323 (N_7323,N_2883,N_4780);
nor U7324 (N_7324,N_4859,N_3403);
xor U7325 (N_7325,N_4638,N_3621);
xor U7326 (N_7326,N_4048,N_3779);
xor U7327 (N_7327,N_4479,N_4646);
or U7328 (N_7328,N_4615,N_4142);
nor U7329 (N_7329,N_3573,N_4360);
xor U7330 (N_7330,N_3032,N_4876);
or U7331 (N_7331,N_4933,N_4173);
nand U7332 (N_7332,N_2531,N_2559);
xnor U7333 (N_7333,N_3585,N_3154);
or U7334 (N_7334,N_4154,N_4445);
xnor U7335 (N_7335,N_4402,N_4324);
xor U7336 (N_7336,N_4726,N_3067);
and U7337 (N_7337,N_2805,N_3391);
nor U7338 (N_7338,N_2582,N_4654);
xnor U7339 (N_7339,N_4121,N_2599);
and U7340 (N_7340,N_4432,N_2669);
nor U7341 (N_7341,N_2813,N_2630);
nand U7342 (N_7342,N_3635,N_3068);
or U7343 (N_7343,N_4525,N_3294);
nand U7344 (N_7344,N_3186,N_4649);
nand U7345 (N_7345,N_2700,N_3710);
xnor U7346 (N_7346,N_2726,N_3095);
and U7347 (N_7347,N_4620,N_3187);
nand U7348 (N_7348,N_4074,N_3413);
nor U7349 (N_7349,N_2618,N_3174);
or U7350 (N_7350,N_3792,N_4163);
and U7351 (N_7351,N_2997,N_2579);
and U7352 (N_7352,N_4156,N_3538);
nand U7353 (N_7353,N_3040,N_4872);
or U7354 (N_7354,N_3035,N_4332);
and U7355 (N_7355,N_2659,N_3126);
xor U7356 (N_7356,N_4185,N_3827);
nor U7357 (N_7357,N_3089,N_4062);
xnor U7358 (N_7358,N_4981,N_4813);
nor U7359 (N_7359,N_4166,N_4920);
or U7360 (N_7360,N_2903,N_3587);
nand U7361 (N_7361,N_4697,N_3913);
nand U7362 (N_7362,N_2638,N_3698);
or U7363 (N_7363,N_4891,N_3667);
or U7364 (N_7364,N_2617,N_3631);
or U7365 (N_7365,N_4127,N_4499);
or U7366 (N_7366,N_2911,N_3563);
and U7367 (N_7367,N_4857,N_3372);
xnor U7368 (N_7368,N_3151,N_2539);
and U7369 (N_7369,N_4964,N_3386);
nand U7370 (N_7370,N_3400,N_2811);
or U7371 (N_7371,N_3900,N_3426);
nor U7372 (N_7372,N_4474,N_2505);
nand U7373 (N_7373,N_3364,N_3944);
and U7374 (N_7374,N_2916,N_3267);
nand U7375 (N_7375,N_4859,N_2632);
nor U7376 (N_7376,N_2954,N_2600);
nand U7377 (N_7377,N_2770,N_4410);
or U7378 (N_7378,N_4588,N_3531);
xnor U7379 (N_7379,N_2900,N_3793);
nand U7380 (N_7380,N_3106,N_3352);
and U7381 (N_7381,N_4819,N_3833);
and U7382 (N_7382,N_4660,N_4593);
xnor U7383 (N_7383,N_3203,N_3586);
or U7384 (N_7384,N_3733,N_2792);
nand U7385 (N_7385,N_3026,N_2777);
xor U7386 (N_7386,N_2987,N_3797);
nor U7387 (N_7387,N_4057,N_4882);
or U7388 (N_7388,N_4120,N_2766);
nand U7389 (N_7389,N_2782,N_4342);
or U7390 (N_7390,N_4889,N_2800);
nor U7391 (N_7391,N_2648,N_4821);
and U7392 (N_7392,N_3785,N_3463);
nor U7393 (N_7393,N_3636,N_3655);
nor U7394 (N_7394,N_4098,N_4625);
and U7395 (N_7395,N_4401,N_4423);
nand U7396 (N_7396,N_3323,N_3324);
or U7397 (N_7397,N_2587,N_4574);
nand U7398 (N_7398,N_4658,N_4328);
and U7399 (N_7399,N_4566,N_4486);
or U7400 (N_7400,N_2885,N_2915);
and U7401 (N_7401,N_4323,N_3407);
nor U7402 (N_7402,N_2806,N_4030);
or U7403 (N_7403,N_4775,N_3101);
or U7404 (N_7404,N_4906,N_3201);
and U7405 (N_7405,N_3027,N_4537);
and U7406 (N_7406,N_4377,N_4642);
or U7407 (N_7407,N_3005,N_4422);
or U7408 (N_7408,N_4210,N_3929);
xnor U7409 (N_7409,N_3907,N_2792);
xor U7410 (N_7410,N_3538,N_3182);
xnor U7411 (N_7411,N_2952,N_3386);
and U7412 (N_7412,N_4093,N_4473);
xor U7413 (N_7413,N_4313,N_3089);
nand U7414 (N_7414,N_3628,N_2991);
and U7415 (N_7415,N_4087,N_2560);
and U7416 (N_7416,N_3208,N_4015);
nor U7417 (N_7417,N_4387,N_3453);
nor U7418 (N_7418,N_3602,N_4164);
nor U7419 (N_7419,N_4211,N_3586);
xnor U7420 (N_7420,N_4204,N_2582);
nand U7421 (N_7421,N_4690,N_2977);
xor U7422 (N_7422,N_2877,N_2801);
or U7423 (N_7423,N_3680,N_4358);
nand U7424 (N_7424,N_4534,N_3672);
nand U7425 (N_7425,N_4930,N_3957);
nor U7426 (N_7426,N_3436,N_2623);
nand U7427 (N_7427,N_4112,N_3642);
xnor U7428 (N_7428,N_3514,N_4440);
nand U7429 (N_7429,N_2844,N_4239);
nand U7430 (N_7430,N_4676,N_4228);
and U7431 (N_7431,N_3476,N_2525);
nand U7432 (N_7432,N_2692,N_2916);
nor U7433 (N_7433,N_2957,N_2709);
xor U7434 (N_7434,N_4938,N_4039);
and U7435 (N_7435,N_4993,N_4896);
and U7436 (N_7436,N_2884,N_3375);
nand U7437 (N_7437,N_2940,N_2907);
xor U7438 (N_7438,N_4615,N_4516);
or U7439 (N_7439,N_4970,N_4468);
and U7440 (N_7440,N_4576,N_4110);
nand U7441 (N_7441,N_4878,N_2815);
and U7442 (N_7442,N_3107,N_3262);
xor U7443 (N_7443,N_3731,N_2794);
nor U7444 (N_7444,N_2715,N_4852);
nor U7445 (N_7445,N_4150,N_2830);
or U7446 (N_7446,N_4228,N_4573);
xor U7447 (N_7447,N_2869,N_3999);
and U7448 (N_7448,N_3018,N_4920);
and U7449 (N_7449,N_3417,N_4592);
xnor U7450 (N_7450,N_3636,N_4933);
nor U7451 (N_7451,N_2844,N_3249);
or U7452 (N_7452,N_3066,N_3794);
or U7453 (N_7453,N_2735,N_3259);
xnor U7454 (N_7454,N_2586,N_2511);
or U7455 (N_7455,N_2702,N_3151);
and U7456 (N_7456,N_4928,N_3671);
nor U7457 (N_7457,N_3101,N_3116);
nor U7458 (N_7458,N_3878,N_4162);
and U7459 (N_7459,N_3368,N_4424);
nand U7460 (N_7460,N_3872,N_4557);
or U7461 (N_7461,N_3004,N_4168);
and U7462 (N_7462,N_3343,N_3258);
xnor U7463 (N_7463,N_2872,N_4996);
nand U7464 (N_7464,N_4515,N_4755);
nor U7465 (N_7465,N_4036,N_4519);
xor U7466 (N_7466,N_3628,N_4923);
nand U7467 (N_7467,N_4410,N_2752);
nand U7468 (N_7468,N_3392,N_3769);
or U7469 (N_7469,N_4309,N_2738);
nand U7470 (N_7470,N_4522,N_4206);
and U7471 (N_7471,N_4251,N_2653);
nand U7472 (N_7472,N_4626,N_2826);
and U7473 (N_7473,N_3442,N_2638);
nor U7474 (N_7474,N_4931,N_3281);
or U7475 (N_7475,N_4526,N_3231);
and U7476 (N_7476,N_3715,N_2558);
and U7477 (N_7477,N_4941,N_4810);
and U7478 (N_7478,N_3222,N_4724);
or U7479 (N_7479,N_4969,N_3841);
and U7480 (N_7480,N_3682,N_3757);
nand U7481 (N_7481,N_2936,N_4006);
xnor U7482 (N_7482,N_4222,N_2730);
xnor U7483 (N_7483,N_2756,N_4384);
or U7484 (N_7484,N_4214,N_3097);
nand U7485 (N_7485,N_3708,N_3997);
nand U7486 (N_7486,N_3835,N_3213);
or U7487 (N_7487,N_4904,N_4228);
and U7488 (N_7488,N_3089,N_3476);
nand U7489 (N_7489,N_4035,N_4285);
and U7490 (N_7490,N_3915,N_2826);
or U7491 (N_7491,N_4098,N_2621);
nor U7492 (N_7492,N_4363,N_3508);
or U7493 (N_7493,N_4478,N_2970);
or U7494 (N_7494,N_4559,N_3200);
xor U7495 (N_7495,N_4915,N_3142);
or U7496 (N_7496,N_4558,N_3879);
nand U7497 (N_7497,N_2598,N_3678);
or U7498 (N_7498,N_3622,N_2915);
nand U7499 (N_7499,N_2719,N_3704);
or U7500 (N_7500,N_6443,N_5139);
nor U7501 (N_7501,N_6015,N_5571);
xor U7502 (N_7502,N_5828,N_6772);
nor U7503 (N_7503,N_7094,N_7155);
xor U7504 (N_7504,N_6152,N_6936);
nand U7505 (N_7505,N_5770,N_6328);
or U7506 (N_7506,N_6161,N_6764);
and U7507 (N_7507,N_5366,N_5692);
or U7508 (N_7508,N_7389,N_6138);
xnor U7509 (N_7509,N_5167,N_5838);
nor U7510 (N_7510,N_6584,N_5782);
and U7511 (N_7511,N_7360,N_6830);
or U7512 (N_7512,N_5153,N_5271);
or U7513 (N_7513,N_6568,N_5641);
xor U7514 (N_7514,N_6230,N_5487);
xnor U7515 (N_7515,N_7107,N_5653);
xnor U7516 (N_7516,N_6991,N_7277);
xnor U7517 (N_7517,N_7001,N_6822);
or U7518 (N_7518,N_6877,N_5773);
and U7519 (N_7519,N_7264,N_7297);
nor U7520 (N_7520,N_7269,N_5588);
nor U7521 (N_7521,N_5951,N_7216);
xor U7522 (N_7522,N_6622,N_5372);
nor U7523 (N_7523,N_6789,N_5978);
or U7524 (N_7524,N_7368,N_7190);
or U7525 (N_7525,N_7146,N_6014);
xnor U7526 (N_7526,N_6605,N_6239);
or U7527 (N_7527,N_5999,N_5132);
or U7528 (N_7528,N_6232,N_5880);
or U7529 (N_7529,N_6905,N_6560);
nand U7530 (N_7530,N_5012,N_5154);
xor U7531 (N_7531,N_7351,N_5022);
or U7532 (N_7532,N_5244,N_5930);
and U7533 (N_7533,N_7486,N_6821);
xor U7534 (N_7534,N_7060,N_5331);
and U7535 (N_7535,N_6064,N_7141);
xnor U7536 (N_7536,N_5907,N_5579);
and U7537 (N_7537,N_6511,N_6653);
xor U7538 (N_7538,N_5870,N_5500);
xnor U7539 (N_7539,N_6059,N_6006);
xor U7540 (N_7540,N_6871,N_5281);
xor U7541 (N_7541,N_7230,N_6460);
or U7542 (N_7542,N_6953,N_6737);
xor U7543 (N_7543,N_7255,N_7312);
xnor U7544 (N_7544,N_7127,N_5850);
or U7545 (N_7545,N_6411,N_6414);
nand U7546 (N_7546,N_6795,N_6043);
xnor U7547 (N_7547,N_5456,N_5634);
xor U7548 (N_7548,N_6253,N_5373);
nand U7549 (N_7549,N_5530,N_6479);
nand U7550 (N_7550,N_7447,N_5582);
or U7551 (N_7551,N_7157,N_6222);
or U7552 (N_7552,N_5556,N_5338);
and U7553 (N_7553,N_6813,N_5702);
or U7554 (N_7554,N_6168,N_6675);
and U7555 (N_7555,N_5704,N_5156);
and U7556 (N_7556,N_6065,N_5750);
nand U7557 (N_7557,N_6782,N_6209);
nor U7558 (N_7558,N_5826,N_5229);
and U7559 (N_7559,N_6918,N_6869);
or U7560 (N_7560,N_7052,N_5399);
nor U7561 (N_7561,N_5248,N_6033);
or U7562 (N_7562,N_5426,N_7338);
nand U7563 (N_7563,N_5663,N_6097);
xor U7564 (N_7564,N_7038,N_5863);
nor U7565 (N_7565,N_7384,N_5474);
or U7566 (N_7566,N_5202,N_6706);
xnor U7567 (N_7567,N_5113,N_6722);
nand U7568 (N_7568,N_5486,N_5097);
nand U7569 (N_7569,N_7200,N_6888);
xor U7570 (N_7570,N_6304,N_5597);
and U7571 (N_7571,N_7032,N_5986);
nand U7572 (N_7572,N_5228,N_7182);
xor U7573 (N_7573,N_6023,N_6846);
and U7574 (N_7574,N_6543,N_5444);
and U7575 (N_7575,N_7379,N_6563);
and U7576 (N_7576,N_5578,N_6638);
nand U7577 (N_7577,N_6652,N_7362);
nand U7578 (N_7578,N_6602,N_6859);
xor U7579 (N_7579,N_5352,N_7130);
nand U7580 (N_7580,N_6494,N_7304);
and U7581 (N_7581,N_5844,N_6051);
xor U7582 (N_7582,N_5878,N_6704);
or U7583 (N_7583,N_6938,N_5059);
and U7584 (N_7584,N_7229,N_7162);
nor U7585 (N_7585,N_6200,N_6252);
nand U7586 (N_7586,N_6787,N_6480);
or U7587 (N_7587,N_5982,N_7075);
or U7588 (N_7588,N_7266,N_5861);
nor U7589 (N_7589,N_6967,N_5317);
or U7590 (N_7590,N_5548,N_5045);
or U7591 (N_7591,N_5542,N_6096);
and U7592 (N_7592,N_6405,N_6393);
nand U7593 (N_7593,N_5807,N_5533);
or U7594 (N_7594,N_5584,N_6113);
and U7595 (N_7595,N_7148,N_7281);
nor U7596 (N_7596,N_7406,N_5551);
xor U7597 (N_7597,N_6863,N_6753);
and U7598 (N_7598,N_6998,N_6768);
or U7599 (N_7599,N_6353,N_6710);
nor U7600 (N_7600,N_5383,N_6866);
nor U7601 (N_7601,N_7374,N_6736);
nor U7602 (N_7602,N_7298,N_6340);
xnor U7603 (N_7603,N_5976,N_6316);
nor U7604 (N_7604,N_5180,N_5420);
or U7605 (N_7605,N_5361,N_6713);
and U7606 (N_7606,N_5381,N_6774);
xnor U7607 (N_7607,N_5470,N_6453);
xnor U7608 (N_7608,N_6763,N_5693);
or U7609 (N_7609,N_5684,N_6211);
nand U7610 (N_7610,N_5145,N_6962);
nor U7611 (N_7611,N_6949,N_6449);
xnor U7612 (N_7612,N_6691,N_5447);
nand U7613 (N_7613,N_5897,N_5403);
nand U7614 (N_7614,N_6132,N_6357);
and U7615 (N_7615,N_5938,N_7345);
xor U7616 (N_7616,N_7414,N_7395);
xor U7617 (N_7617,N_6508,N_6192);
nand U7618 (N_7618,N_5708,N_6355);
and U7619 (N_7619,N_5882,N_5073);
nor U7620 (N_7620,N_5066,N_6326);
xor U7621 (N_7621,N_5287,N_6156);
nor U7622 (N_7622,N_5802,N_5360);
or U7623 (N_7623,N_5952,N_6876);
or U7624 (N_7624,N_5677,N_7472);
or U7625 (N_7625,N_5025,N_5659);
xor U7626 (N_7626,N_6714,N_5929);
and U7627 (N_7627,N_6378,N_5642);
nor U7628 (N_7628,N_5806,N_6044);
xnor U7629 (N_7629,N_6897,N_5491);
and U7630 (N_7630,N_6749,N_6053);
or U7631 (N_7631,N_6343,N_5939);
or U7632 (N_7632,N_5475,N_5747);
nand U7633 (N_7633,N_6016,N_7290);
and U7634 (N_7634,N_5004,N_7308);
or U7635 (N_7635,N_5068,N_6131);
and U7636 (N_7636,N_5232,N_5846);
or U7637 (N_7637,N_5165,N_7464);
xnor U7638 (N_7638,N_5780,N_5618);
and U7639 (N_7639,N_6269,N_6824);
nor U7640 (N_7640,N_5591,N_6784);
nand U7641 (N_7641,N_7084,N_7120);
nor U7642 (N_7642,N_5820,N_6093);
or U7643 (N_7643,N_5353,N_6498);
nor U7644 (N_7644,N_5107,N_5320);
or U7645 (N_7645,N_6671,N_7313);
nand U7646 (N_7646,N_6173,N_6860);
and U7647 (N_7647,N_5356,N_6060);
nor U7648 (N_7648,N_6471,N_6379);
or U7649 (N_7649,N_5606,N_7391);
nor U7650 (N_7650,N_7431,N_5080);
nor U7651 (N_7651,N_5029,N_7169);
and U7652 (N_7652,N_6927,N_6137);
or U7653 (N_7653,N_7006,N_5994);
xnor U7654 (N_7654,N_6042,N_5840);
nor U7655 (N_7655,N_5777,N_6332);
nand U7656 (N_7656,N_6094,N_5241);
and U7657 (N_7657,N_5410,N_5401);
xnor U7658 (N_7658,N_6155,N_6840);
or U7659 (N_7659,N_6867,N_6907);
xnor U7660 (N_7660,N_7133,N_6274);
nand U7661 (N_7661,N_7213,N_7128);
and U7662 (N_7662,N_6164,N_5147);
nand U7663 (N_7663,N_5753,N_6223);
and U7664 (N_7664,N_6424,N_5310);
and U7665 (N_7665,N_6726,N_7367);
or U7666 (N_7666,N_5215,N_5339);
nor U7667 (N_7667,N_7195,N_5944);
xor U7668 (N_7668,N_6818,N_6073);
or U7669 (N_7669,N_5564,N_7025);
and U7670 (N_7670,N_6327,N_5315);
nand U7671 (N_7671,N_6915,N_6878);
or U7672 (N_7672,N_7343,N_6587);
nand U7673 (N_7673,N_7115,N_5297);
and U7674 (N_7674,N_6122,N_7475);
or U7675 (N_7675,N_5687,N_6889);
nor U7676 (N_7676,N_6007,N_6448);
and U7677 (N_7677,N_6382,N_5843);
nand U7678 (N_7678,N_7069,N_6627);
xor U7679 (N_7679,N_7294,N_6573);
nand U7680 (N_7680,N_6788,N_5933);
and U7681 (N_7681,N_5057,N_6189);
xnor U7682 (N_7682,N_6997,N_6520);
xor U7683 (N_7683,N_7165,N_5868);
and U7684 (N_7684,N_7323,N_7329);
nand U7685 (N_7685,N_5342,N_6661);
nor U7686 (N_7686,N_7254,N_5871);
and U7687 (N_7687,N_6215,N_5607);
nand U7688 (N_7688,N_7090,N_5725);
or U7689 (N_7689,N_6906,N_6244);
or U7690 (N_7690,N_7106,N_5645);
or U7691 (N_7691,N_5830,N_6165);
xnor U7692 (N_7692,N_6839,N_5783);
and U7693 (N_7693,N_6350,N_5198);
nand U7694 (N_7694,N_6114,N_6974);
nand U7695 (N_7695,N_5809,N_6194);
nand U7696 (N_7696,N_6021,N_5576);
nor U7697 (N_7697,N_6851,N_6267);
nor U7698 (N_7698,N_7206,N_7174);
nor U7699 (N_7699,N_7272,N_7189);
nor U7700 (N_7700,N_6728,N_7054);
and U7701 (N_7701,N_6349,N_6817);
or U7702 (N_7702,N_5866,N_6538);
or U7703 (N_7703,N_6807,N_6625);
nor U7704 (N_7704,N_7253,N_5221);
nand U7705 (N_7705,N_6960,N_6098);
and U7706 (N_7706,N_5664,N_7402);
or U7707 (N_7707,N_5947,N_6542);
or U7708 (N_7708,N_5164,N_6124);
nor U7709 (N_7709,N_5098,N_5327);
and U7710 (N_7710,N_7187,N_5823);
xor U7711 (N_7711,N_6388,N_5408);
nor U7712 (N_7712,N_6410,N_7116);
and U7713 (N_7713,N_5449,N_7285);
nor U7714 (N_7714,N_7377,N_5799);
xnor U7715 (N_7715,N_5182,N_6146);
or U7716 (N_7716,N_7444,N_7415);
nand U7717 (N_7717,N_5977,N_7357);
or U7718 (N_7718,N_5330,N_6649);
xnor U7719 (N_7719,N_6808,N_7417);
xnor U7720 (N_7720,N_5920,N_6942);
nand U7721 (N_7721,N_6658,N_5661);
and U7722 (N_7722,N_7087,N_6743);
and U7723 (N_7723,N_7261,N_5540);
nor U7724 (N_7724,N_5008,N_5638);
xor U7725 (N_7725,N_5082,N_5083);
nand U7726 (N_7726,N_7467,N_5095);
and U7727 (N_7727,N_5586,N_6019);
nand U7728 (N_7728,N_5214,N_6760);
nand U7729 (N_7729,N_7493,N_7138);
or U7730 (N_7730,N_7341,N_7147);
xor U7731 (N_7731,N_7418,N_5608);
nor U7732 (N_7732,N_7441,N_6115);
nand U7733 (N_7733,N_7082,N_6207);
nor U7734 (N_7734,N_6005,N_5915);
nand U7735 (N_7735,N_5184,N_7434);
and U7736 (N_7736,N_5010,N_6497);
or U7737 (N_7737,N_6950,N_6903);
or U7738 (N_7738,N_5137,N_7086);
nand U7739 (N_7739,N_5031,N_5144);
nand U7740 (N_7740,N_6177,N_7018);
nand U7741 (N_7741,N_6249,N_7435);
xnor U7742 (N_7742,N_5231,N_6716);
or U7743 (N_7743,N_6112,N_5050);
nor U7744 (N_7744,N_5319,N_6488);
xor U7745 (N_7745,N_5676,N_7027);
or U7746 (N_7746,N_6070,N_6307);
nor U7747 (N_7747,N_5849,N_5890);
or U7748 (N_7748,N_5322,N_6086);
xnor U7749 (N_7749,N_6663,N_5262);
or U7750 (N_7750,N_5587,N_7160);
or U7751 (N_7751,N_5266,N_6794);
nand U7752 (N_7752,N_7301,N_5544);
nand U7753 (N_7753,N_6598,N_5289);
nor U7754 (N_7754,N_5974,N_5867);
nor U7755 (N_7755,N_6347,N_6407);
nand U7756 (N_7756,N_5836,N_5768);
nand U7757 (N_7757,N_7325,N_6937);
nand U7758 (N_7758,N_5932,N_7270);
or U7759 (N_7759,N_7008,N_5628);
nand U7760 (N_7760,N_5726,N_5743);
nor U7761 (N_7761,N_6681,N_6484);
nor U7762 (N_7762,N_6783,N_6721);
and U7763 (N_7763,N_7256,N_5392);
xnor U7764 (N_7764,N_6485,N_5419);
nor U7765 (N_7765,N_6752,N_5786);
and U7766 (N_7766,N_6101,N_5227);
or U7767 (N_7767,N_7173,N_6280);
or U7768 (N_7768,N_5854,N_6831);
and U7769 (N_7769,N_6812,N_5672);
and U7770 (N_7770,N_6169,N_6314);
and U7771 (N_7771,N_7470,N_7331);
nor U7772 (N_7772,N_5063,N_5957);
xor U7773 (N_7773,N_5762,N_5972);
and U7774 (N_7774,N_7224,N_5665);
xnor U7775 (N_7775,N_6133,N_5142);
or U7776 (N_7776,N_6444,N_5922);
nand U7777 (N_7777,N_5432,N_5696);
and U7778 (N_7778,N_7119,N_6946);
and U7779 (N_7779,N_6077,N_7283);
nand U7780 (N_7780,N_5111,N_6183);
and U7781 (N_7781,N_7359,N_7131);
and U7782 (N_7782,N_6342,N_5224);
nor U7783 (N_7783,N_6457,N_5463);
nand U7784 (N_7784,N_6723,N_7394);
nand U7785 (N_7785,N_5769,N_7429);
and U7786 (N_7786,N_7124,N_7179);
and U7787 (N_7787,N_5990,N_5539);
or U7788 (N_7788,N_6120,N_7023);
nor U7789 (N_7789,N_6154,N_7387);
and U7790 (N_7790,N_7263,N_6524);
nand U7791 (N_7791,N_5000,N_5494);
or U7792 (N_7792,N_6184,N_6853);
nor U7793 (N_7793,N_7020,N_6618);
and U7794 (N_7794,N_6972,N_6884);
nand U7795 (N_7795,N_7284,N_7476);
xnor U7796 (N_7796,N_5152,N_6694);
nor U7797 (N_7797,N_6487,N_6203);
and U7798 (N_7798,N_7478,N_5506);
nor U7799 (N_7799,N_6549,N_5728);
nor U7800 (N_7800,N_7352,N_6233);
or U7801 (N_7801,N_5928,N_5411);
xnor U7802 (N_7802,N_6761,N_7410);
xnor U7803 (N_7803,N_5461,N_6445);
or U7804 (N_7804,N_5223,N_5135);
nor U7805 (N_7805,N_7064,N_5968);
or U7806 (N_7806,N_6413,N_6447);
nor U7807 (N_7807,N_6049,N_6219);
and U7808 (N_7808,N_5033,N_5170);
and U7809 (N_7809,N_6909,N_5313);
or U7810 (N_7810,N_5916,N_6948);
nand U7811 (N_7811,N_5041,N_6231);
and U7812 (N_7812,N_6850,N_5163);
or U7813 (N_7813,N_5141,N_7028);
or U7814 (N_7814,N_5737,N_6957);
nor U7815 (N_7815,N_5812,N_7123);
nand U7816 (N_7816,N_6703,N_5208);
xor U7817 (N_7817,N_5964,N_6136);
nand U7818 (N_7818,N_5518,N_6188);
and U7819 (N_7819,N_5434,N_7227);
and U7820 (N_7820,N_5473,N_7457);
nand U7821 (N_7821,N_5765,N_6654);
nand U7822 (N_7822,N_6576,N_5171);
or U7823 (N_7823,N_7029,N_7488);
and U7824 (N_7824,N_7007,N_5872);
xor U7825 (N_7825,N_7428,N_6970);
nand U7826 (N_7826,N_5931,N_5176);
and U7827 (N_7827,N_5752,N_6791);
or U7828 (N_7828,N_5341,N_7365);
xor U7829 (N_7829,N_5568,N_5018);
xnor U7830 (N_7830,N_7065,N_5980);
nor U7831 (N_7831,N_6197,N_5336);
nor U7832 (N_7832,N_5776,N_6744);
xnor U7833 (N_7833,N_6930,N_6474);
xor U7834 (N_7834,N_5899,N_5102);
or U7835 (N_7835,N_6862,N_6462);
or U7836 (N_7836,N_6130,N_5669);
nand U7837 (N_7837,N_6275,N_7142);
nor U7838 (N_7838,N_5015,N_5819);
and U7839 (N_7839,N_5610,N_6557);
nand U7840 (N_7840,N_6592,N_7482);
nand U7841 (N_7841,N_5821,N_7150);
xnor U7842 (N_7842,N_6509,N_5927);
or U7843 (N_7843,N_5744,N_7209);
xor U7844 (N_7844,N_5671,N_5685);
nand U7845 (N_7845,N_5577,N_6922);
xnor U7846 (N_7846,N_5326,N_6535);
xnor U7847 (N_7847,N_6987,N_5894);
nor U7848 (N_7848,N_6740,N_6178);
nor U7849 (N_7849,N_6017,N_6291);
nor U7850 (N_7850,N_5742,N_5547);
and U7851 (N_7851,N_7337,N_6372);
nand U7852 (N_7852,N_7219,N_6153);
nand U7853 (N_7853,N_6456,N_7121);
xor U7854 (N_7854,N_7014,N_5344);
nor U7855 (N_7855,N_6100,N_6495);
or U7856 (N_7856,N_7423,N_5567);
xnor U7857 (N_7857,N_5283,N_7088);
or U7858 (N_7858,N_7140,N_7401);
and U7859 (N_7859,N_6331,N_5312);
nand U7860 (N_7860,N_6567,N_6078);
nand U7861 (N_7861,N_6301,N_6160);
nand U7862 (N_7862,N_7349,N_5496);
or U7863 (N_7863,N_6678,N_5575);
and U7864 (N_7864,N_6110,N_7045);
xnor U7865 (N_7865,N_7099,N_6548);
or U7866 (N_7866,N_5055,N_5125);
nand U7867 (N_7867,N_6384,N_7480);
nand U7868 (N_7868,N_6010,N_5794);
and U7869 (N_7869,N_6026,N_5296);
and U7870 (N_7870,N_5406,N_7332);
nand U7871 (N_7871,N_6258,N_7311);
or U7872 (N_7872,N_5954,N_7363);
or U7873 (N_7873,N_5950,N_7072);
nand U7874 (N_7874,N_7059,N_5829);
nand U7875 (N_7875,N_5531,N_6368);
xor U7876 (N_7876,N_7328,N_6606);
xor U7877 (N_7877,N_6395,N_5695);
xnor U7878 (N_7878,N_6297,N_5975);
nor U7879 (N_7879,N_5457,N_5417);
or U7880 (N_7880,N_5605,N_7288);
xnor U7881 (N_7881,N_6455,N_5604);
or U7882 (N_7882,N_5711,N_6874);
nand U7883 (N_7883,N_6002,N_6500);
nor U7884 (N_7884,N_6147,N_6356);
or U7885 (N_7885,N_5409,N_5757);
or U7886 (N_7886,N_6717,N_5797);
nand U7887 (N_7887,N_5323,N_6963);
nor U7888 (N_7888,N_7050,N_5959);
xor U7889 (N_7889,N_7404,N_6529);
and U7890 (N_7890,N_7421,N_5114);
and U7891 (N_7891,N_6739,N_6354);
nand U7892 (N_7892,N_6076,N_7348);
or U7893 (N_7893,N_5649,N_7129);
nor U7894 (N_7894,N_7320,N_7056);
and U7895 (N_7895,N_5825,N_5919);
and U7896 (N_7896,N_6913,N_6400);
or U7897 (N_7897,N_7246,N_5527);
nand U7898 (N_7898,N_6667,N_7275);
or U7899 (N_7899,N_6090,N_6000);
nand U7900 (N_7900,N_5077,N_6510);
and U7901 (N_7901,N_7234,N_5458);
or U7902 (N_7902,N_6063,N_5877);
nand U7903 (N_7903,N_6008,N_5620);
or U7904 (N_7904,N_5379,N_5442);
xnor U7905 (N_7905,N_6080,N_5632);
xor U7906 (N_7906,N_5790,N_6778);
nor U7907 (N_7907,N_6159,N_7035);
xor U7908 (N_7908,N_6095,N_6246);
or U7909 (N_7909,N_6170,N_5875);
or U7910 (N_7910,N_7026,N_5488);
nand U7911 (N_7911,N_6935,N_5013);
nand U7912 (N_7912,N_7296,N_6614);
and U7913 (N_7913,N_6259,N_5291);
or U7914 (N_7914,N_6346,N_5078);
xor U7915 (N_7915,N_6118,N_5534);
nor U7916 (N_7916,N_6483,N_6699);
or U7917 (N_7917,N_5913,N_5650);
nor U7918 (N_7918,N_5508,N_5199);
or U7919 (N_7919,N_5380,N_7137);
nand U7920 (N_7920,N_5949,N_6220);
nor U7921 (N_7921,N_7080,N_5699);
nand U7922 (N_7922,N_6797,N_6682);
xnor U7923 (N_7923,N_6245,N_5204);
xor U7924 (N_7924,N_6556,N_5358);
nor U7925 (N_7925,N_5321,N_7043);
nand U7926 (N_7926,N_7456,N_5679);
and U7927 (N_7927,N_6732,N_5636);
nand U7928 (N_7928,N_7228,N_6242);
nor U7929 (N_7929,N_7247,N_6106);
nand U7930 (N_7930,N_6037,N_7485);
nor U7931 (N_7931,N_6522,N_7199);
and U7932 (N_7932,N_7175,N_6011);
or U7933 (N_7933,N_6345,N_7490);
nand U7934 (N_7934,N_5722,N_6873);
nor U7935 (N_7935,N_7271,N_6525);
xor U7936 (N_7936,N_5479,N_5398);
nor U7937 (N_7937,N_6157,N_6381);
and U7938 (N_7938,N_5934,N_7412);
nand U7939 (N_7939,N_7222,N_5128);
nor U7940 (N_7940,N_7262,N_5914);
nand U7941 (N_7941,N_5953,N_5414);
nand U7942 (N_7942,N_7496,N_6558);
or U7943 (N_7943,N_7037,N_5332);
or U7944 (N_7944,N_6361,N_6046);
nor U7945 (N_7945,N_5595,N_6366);
nand U7946 (N_7946,N_5465,N_6908);
nor U7947 (N_7947,N_7408,N_6450);
xor U7948 (N_7948,N_7217,N_5079);
or U7949 (N_7949,N_5136,N_5759);
xor U7950 (N_7950,N_6452,N_6589);
xor U7951 (N_7951,N_5528,N_5335);
nand U7952 (N_7952,N_5749,N_6176);
and U7953 (N_7953,N_5637,N_5143);
and U7954 (N_7954,N_5503,N_6319);
xnor U7955 (N_7955,N_5306,N_7392);
and U7956 (N_7956,N_5691,N_5697);
xor U7957 (N_7957,N_6911,N_5084);
or U7958 (N_7958,N_5874,N_6641);
and U7959 (N_7959,N_5761,N_6647);
nor U7960 (N_7960,N_5804,N_6898);
or U7961 (N_7961,N_6885,N_6607);
and U7962 (N_7962,N_7382,N_5039);
xnor U7963 (N_7963,N_6143,N_6300);
and U7964 (N_7964,N_6254,N_5276);
and U7965 (N_7965,N_5881,N_6193);
xor U7966 (N_7966,N_6683,N_6854);
nor U7967 (N_7967,N_5583,N_5523);
nor U7968 (N_7968,N_6123,N_6527);
nand U7969 (N_7969,N_6061,N_5425);
xnor U7970 (N_7970,N_6550,N_6828);
nor U7971 (N_7971,N_5209,N_6872);
nand U7972 (N_7972,N_5350,N_6952);
xor U7973 (N_7973,N_6311,N_6707);
nand U7974 (N_7974,N_5158,N_6358);
or U7975 (N_7975,N_7451,N_7342);
nand U7976 (N_7976,N_6284,N_5443);
nor U7977 (N_7977,N_6276,N_7450);
and U7978 (N_7978,N_5061,N_5429);
and U7979 (N_7979,N_6746,N_5834);
xnor U7980 (N_7980,N_6074,N_6362);
nor U7981 (N_7981,N_6079,N_5853);
xor U7982 (N_7982,N_5477,N_7425);
xor U7983 (N_7983,N_6312,N_7442);
or U7984 (N_7984,N_6264,N_7321);
or U7985 (N_7985,N_5210,N_5510);
and U7986 (N_7986,N_5720,N_6621);
and U7987 (N_7987,N_6038,N_5075);
or U7988 (N_7988,N_6099,N_6265);
and U7989 (N_7989,N_5028,N_6816);
nor U7990 (N_7990,N_6486,N_6306);
nor U7991 (N_7991,N_5482,N_5424);
nor U7992 (N_7992,N_5521,N_5178);
nor U7993 (N_7993,N_6650,N_5601);
and U7994 (N_7994,N_7237,N_7170);
nor U7995 (N_7995,N_7193,N_6934);
or U7996 (N_7996,N_5355,N_5440);
nand U7997 (N_7997,N_5112,N_6171);
nor U7998 (N_7998,N_5557,N_7145);
nor U7999 (N_7999,N_5299,N_7369);
nor U8000 (N_8000,N_5104,N_5105);
and U8001 (N_8001,N_5755,N_5448);
and U8002 (N_8002,N_7031,N_6856);
nor U8003 (N_8003,N_6684,N_6213);
nand U8004 (N_8004,N_7117,N_5017);
nor U8005 (N_8005,N_5879,N_6091);
and U8006 (N_8006,N_6977,N_6442);
or U8007 (N_8007,N_6541,N_5668);
xor U8008 (N_8008,N_5689,N_5643);
xnor U8009 (N_8009,N_5249,N_6982);
xnor U8010 (N_8010,N_6947,N_7245);
nor U8011 (N_8011,N_5309,N_5284);
nand U8012 (N_8012,N_6464,N_6886);
and U8013 (N_8013,N_6570,N_6688);
nor U8014 (N_8014,N_5764,N_6506);
and U8015 (N_8015,N_6646,N_6376);
xor U8016 (N_8016,N_6092,N_7453);
nor U8017 (N_8017,N_5760,N_6552);
nor U8018 (N_8018,N_5437,N_6389);
nand U8019 (N_8019,N_7291,N_5280);
nor U8020 (N_8020,N_7232,N_5391);
and U8021 (N_8021,N_5775,N_5051);
xnor U8022 (N_8022,N_6283,N_6940);
or U8023 (N_8023,N_6435,N_6575);
or U8024 (N_8024,N_6196,N_6904);
and U8025 (N_8025,N_6923,N_5151);
or U8026 (N_8026,N_6664,N_6417);
and U8027 (N_8027,N_5225,N_7186);
nand U8028 (N_8028,N_6958,N_6458);
nor U8029 (N_8029,N_6374,N_5060);
or U8030 (N_8030,N_5325,N_7463);
or U8031 (N_8031,N_6582,N_5468);
xnor U8032 (N_8032,N_7248,N_5222);
nand U8033 (N_8033,N_6296,N_7449);
and U8034 (N_8034,N_7252,N_5115);
nor U8035 (N_8035,N_6882,N_5181);
nor U8036 (N_8036,N_6790,N_6968);
xnor U8037 (N_8037,N_7100,N_6126);
nand U8038 (N_8038,N_6633,N_5707);
nand U8039 (N_8039,N_5888,N_5285);
nand U8040 (N_8040,N_5454,N_5735);
nor U8041 (N_8041,N_6351,N_6864);
xnor U8042 (N_8042,N_7350,N_6980);
and U8043 (N_8043,N_5450,N_7210);
and U8044 (N_8044,N_5393,N_6674);
nand U8045 (N_8045,N_6827,N_7400);
xnor U8046 (N_8046,N_6518,N_5146);
nor U8047 (N_8047,N_7495,N_6755);
and U8048 (N_8048,N_5481,N_5859);
and U8049 (N_8049,N_7249,N_6425);
and U8050 (N_8050,N_6993,N_5624);
or U8051 (N_8051,N_7318,N_6191);
nand U8052 (N_8052,N_6377,N_6102);
or U8053 (N_8053,N_7113,N_5226);
and U8054 (N_8054,N_6881,N_5713);
xor U8055 (N_8055,N_6468,N_5382);
xnor U8056 (N_8056,N_6978,N_5027);
xor U8057 (N_8057,N_7197,N_7487);
and U8058 (N_8058,N_5791,N_7108);
and U8059 (N_8059,N_5295,N_5026);
nor U8060 (N_8060,N_6375,N_5729);
nor U8061 (N_8061,N_6656,N_5367);
or U8062 (N_8062,N_5376,N_6067);
xor U8063 (N_8063,N_7405,N_5700);
nor U8064 (N_8064,N_5889,N_7164);
xnor U8065 (N_8065,N_5842,N_5157);
or U8066 (N_8066,N_6365,N_6870);
or U8067 (N_8067,N_5988,N_5441);
nor U8068 (N_8068,N_6648,N_5763);
nand U8069 (N_8069,N_6914,N_7440);
nand U8070 (N_8070,N_6334,N_6562);
nand U8071 (N_8071,N_5270,N_7492);
nor U8072 (N_8072,N_6270,N_5946);
xor U8073 (N_8073,N_7494,N_7091);
nor U8074 (N_8074,N_5130,N_6397);
nand U8075 (N_8075,N_5340,N_5817);
nor U8076 (N_8076,N_6333,N_6204);
or U8077 (N_8077,N_6229,N_6048);
and U8078 (N_8078,N_6603,N_6762);
nor U8079 (N_8079,N_5796,N_5848);
nor U8080 (N_8080,N_6205,N_5851);
and U8081 (N_8081,N_7448,N_7104);
nand U8082 (N_8082,N_6227,N_5264);
or U8083 (N_8083,N_5492,N_6989);
xor U8084 (N_8084,N_6610,N_7201);
and U8085 (N_8085,N_7058,N_5810);
and U8086 (N_8086,N_5126,N_6917);
and U8087 (N_8087,N_6601,N_7071);
nand U8088 (N_8088,N_6243,N_5856);
nand U8089 (N_8089,N_6701,N_5909);
nand U8090 (N_8090,N_6055,N_5635);
and U8091 (N_8091,N_5580,N_6256);
xnor U8092 (N_8092,N_7221,N_6315);
nand U8093 (N_8093,N_5543,N_6235);
xnor U8094 (N_8094,N_6895,N_5252);
nand U8095 (N_8095,N_7017,N_5265);
nand U8096 (N_8096,N_6708,N_5189);
or U8097 (N_8097,N_6748,N_6632);
xnor U8098 (N_8098,N_7126,N_7167);
or U8099 (N_8099,N_5275,N_5839);
nor U8100 (N_8100,N_5886,N_5436);
nor U8101 (N_8101,N_6338,N_5710);
xnor U8102 (N_8102,N_7109,N_6050);
and U8103 (N_8103,N_6634,N_5172);
or U8104 (N_8104,N_6891,N_6117);
nand U8105 (N_8105,N_5688,N_7280);
xor U8106 (N_8106,N_6305,N_6580);
xor U8107 (N_8107,N_5852,N_6322);
nor U8108 (N_8108,N_6294,N_6491);
xnor U8109 (N_8109,N_6855,N_5598);
xor U8110 (N_8110,N_6473,N_5324);
or U8111 (N_8111,N_5658,N_6225);
nor U8112 (N_8112,N_5207,N_6181);
xnor U8113 (N_8113,N_5385,N_6800);
or U8114 (N_8114,N_6900,N_5374);
or U8115 (N_8115,N_7267,N_6437);
nand U8116 (N_8116,N_5002,N_5514);
and U8117 (N_8117,N_5100,N_5430);
and U8118 (N_8118,N_7443,N_5455);
and U8119 (N_8119,N_6672,N_6577);
xnor U8120 (N_8120,N_5278,N_6472);
nor U8121 (N_8121,N_6216,N_5905);
nand U8122 (N_8122,N_5499,N_6964);
or U8123 (N_8123,N_5970,N_5893);
nand U8124 (N_8124,N_6569,N_5065);
nor U8125 (N_8125,N_5626,N_5683);
nand U8126 (N_8126,N_6248,N_6369);
or U8127 (N_8127,N_5787,N_6547);
nand U8128 (N_8128,N_5599,N_5368);
or U8129 (N_8129,N_6594,N_7196);
xor U8130 (N_8130,N_7061,N_5246);
and U8131 (N_8131,N_6271,N_5462);
or U8132 (N_8132,N_5832,N_5816);
nand U8133 (N_8133,N_7289,N_7015);
nor U8134 (N_8134,N_7309,N_6320);
nand U8135 (N_8135,N_6711,N_6690);
xor U8136 (N_8136,N_6685,N_5501);
or U8137 (N_8137,N_7334,N_5040);
nor U8138 (N_8138,N_6657,N_5483);
nand U8139 (N_8139,N_7243,N_5633);
and U8140 (N_8140,N_5781,N_5719);
or U8141 (N_8141,N_7144,N_5921);
or U8142 (N_8142,N_7079,N_6660);
xnor U8143 (N_8143,N_5627,N_5989);
nand U8144 (N_8144,N_5122,N_5192);
nand U8145 (N_8145,N_5550,N_6363);
nor U8146 (N_8146,N_6292,N_6825);
nor U8147 (N_8147,N_5795,N_6910);
nand U8148 (N_8148,N_6961,N_6799);
and U8149 (N_8149,N_7156,N_6966);
and U8150 (N_8150,N_7143,N_6426);
nand U8151 (N_8151,N_5074,N_7286);
nor U8152 (N_8152,N_6172,N_5767);
or U8153 (N_8153,N_5570,N_5662);
nand U8154 (N_8154,N_5522,N_6835);
or U8155 (N_8155,N_5304,N_6403);
nor U8156 (N_8156,N_5991,N_7233);
nand U8157 (N_8157,N_6780,N_5149);
nor U8158 (N_8158,N_5504,N_5858);
nor U8159 (N_8159,N_5967,N_5788);
nor U8160 (N_8160,N_6396,N_6031);
nor U8161 (N_8161,N_7112,N_6720);
and U8162 (N_8162,N_6742,N_6677);
or U8163 (N_8163,N_7235,N_6698);
nand U8164 (N_8164,N_6103,N_5517);
xor U8165 (N_8165,N_6617,N_5005);
nand U8166 (N_8166,N_6446,N_5138);
or U8167 (N_8167,N_6089,N_6697);
xnor U8168 (N_8168,N_5049,N_5109);
nor U8169 (N_8169,N_5592,N_6507);
nor U8170 (N_8170,N_7326,N_5386);
nand U8171 (N_8171,N_6912,N_6609);
xnor U8172 (N_8172,N_5329,N_6841);
or U8173 (N_8173,N_6933,N_6775);
nand U8174 (N_8174,N_6528,N_6206);
nor U8175 (N_8175,N_6973,N_7236);
nor U8176 (N_8176,N_6013,N_5910);
and U8177 (N_8177,N_6260,N_5908);
and U8178 (N_8178,N_6637,N_7473);
xor U8179 (N_8179,N_7192,N_5801);
nor U8180 (N_8180,N_5316,N_5505);
or U8181 (N_8181,N_5640,N_5524);
nand U8182 (N_8182,N_7205,N_5709);
xnor U8183 (N_8183,N_7498,N_6024);
xor U8184 (N_8184,N_6140,N_5733);
nand U8185 (N_8185,N_5328,N_6734);
or U8186 (N_8186,N_5235,N_6999);
or U8187 (N_8187,N_5174,N_5096);
nor U8188 (N_8188,N_6921,N_6865);
nand U8189 (N_8189,N_6695,N_5212);
xnor U8190 (N_8190,N_5023,N_5286);
and U8191 (N_8191,N_5351,N_5175);
xor U8192 (N_8192,N_6599,N_6439);
xor U8193 (N_8193,N_5857,N_5585);
and U8194 (N_8194,N_6845,N_6250);
nor U8195 (N_8195,N_6939,N_6069);
or U8196 (N_8196,N_7432,N_5261);
nand U8197 (N_8197,N_6561,N_5402);
xnor U8198 (N_8198,N_7471,N_5290);
nor U8199 (N_8199,N_6371,N_6398);
nand U8200 (N_8200,N_5451,N_6988);
nand U8201 (N_8201,N_6290,N_6644);
nand U8202 (N_8202,N_5615,N_6955);
xnor U8203 (N_8203,N_5731,N_7077);
and U8204 (N_8204,N_5923,N_5942);
or U8205 (N_8205,N_6041,N_5394);
nand U8206 (N_8206,N_5407,N_5779);
xor U8207 (N_8207,N_6399,N_6985);
and U8208 (N_8208,N_7153,N_6492);
xor U8209 (N_8209,N_6127,N_5561);
xnor U8210 (N_8210,N_5519,N_7172);
nor U8211 (N_8211,N_5390,N_6792);
or U8212 (N_8212,N_6719,N_7000);
or U8213 (N_8213,N_6765,N_5433);
nor U8214 (N_8214,N_5581,N_5091);
and U8215 (N_8215,N_5800,N_7163);
nor U8216 (N_8216,N_5201,N_5525);
xnor U8217 (N_8217,N_7239,N_5250);
nor U8218 (N_8218,N_6893,N_7439);
nand U8219 (N_8219,N_5739,N_5814);
nand U8220 (N_8220,N_5529,N_5069);
or U8221 (N_8221,N_6591,N_5895);
nor U8222 (N_8222,N_5118,N_7039);
or U8223 (N_8223,N_6212,N_5766);
or U8224 (N_8224,N_6476,N_6255);
nor U8225 (N_8225,N_7204,N_7293);
and U8226 (N_8226,N_5831,N_5981);
nor U8227 (N_8227,N_5639,N_7066);
nand U8228 (N_8228,N_7242,N_5694);
nor U8229 (N_8229,N_5758,N_5948);
and U8230 (N_8230,N_6802,N_7386);
nand U8231 (N_8231,N_6545,N_6380);
nand U8232 (N_8232,N_5121,N_7183);
or U8233 (N_8233,N_5936,N_7111);
and U8234 (N_8234,N_5862,N_7016);
xor U8235 (N_8235,N_5898,N_5987);
nand U8236 (N_8236,N_5730,N_6626);
nand U8237 (N_8237,N_6519,N_5537);
nand U8238 (N_8238,N_6628,N_5070);
and U8239 (N_8239,N_5705,N_5446);
and U8240 (N_8240,N_6020,N_5555);
nand U8241 (N_8241,N_7282,N_6135);
nand U8242 (N_8242,N_6180,N_6776);
and U8243 (N_8243,N_6045,N_7335);
or U8244 (N_8244,N_6842,N_5048);
xor U8245 (N_8245,N_5973,N_6145);
and U8246 (N_8246,N_6572,N_5303);
nor U8247 (N_8247,N_5484,N_6536);
nand U8248 (N_8248,N_6385,N_6530);
nand U8249 (N_8249,N_5343,N_6036);
nand U8250 (N_8250,N_5546,N_5088);
and U8251 (N_8251,N_5007,N_7265);
xor U8252 (N_8252,N_5901,N_5203);
nand U8253 (N_8253,N_5785,N_7240);
or U8254 (N_8254,N_5423,N_6767);
and U8255 (N_8255,N_7207,N_6666);
or U8256 (N_8256,N_6210,N_6257);
nand U8257 (N_8257,N_6310,N_5535);
nand U8258 (N_8258,N_5101,N_5751);
nor U8259 (N_8259,N_5803,N_6034);
nor U8260 (N_8260,N_5734,N_6773);
or U8261 (N_8261,N_5120,N_6941);
nor U8262 (N_8262,N_6470,N_6218);
xnor U8263 (N_8263,N_5906,N_7468);
nand U8264 (N_8264,N_7499,N_5058);
or U8265 (N_8265,N_6083,N_7102);
or U8266 (N_8266,N_6513,N_6747);
and U8267 (N_8267,N_6995,N_6430);
nor U8268 (N_8268,N_5602,N_6919);
and U8269 (N_8269,N_7424,N_5254);
xor U8270 (N_8270,N_6287,N_5219);
nand U8271 (N_8271,N_6571,N_6805);
nor U8272 (N_8272,N_7316,N_6463);
nor U8273 (N_8273,N_6402,N_5062);
nand U8274 (N_8274,N_5099,N_5301);
nand U8275 (N_8275,N_5489,N_5675);
and U8276 (N_8276,N_5630,N_6693);
or U8277 (N_8277,N_6009,N_5962);
or U8278 (N_8278,N_5044,N_6623);
or U8279 (N_8279,N_6636,N_6066);
xnor U8280 (N_8280,N_7358,N_5003);
nor U8281 (N_8281,N_7419,N_5106);
and U8282 (N_8282,N_6052,N_5133);
and U8283 (N_8283,N_5016,N_5168);
nor U8284 (N_8284,N_5193,N_6620);
xor U8285 (N_8285,N_6809,N_7375);
xor U8286 (N_8286,N_6837,N_5439);
xor U8287 (N_8287,N_7469,N_5185);
nand U8288 (N_8288,N_6640,N_5076);
and U8289 (N_8289,N_7095,N_5251);
nor U8290 (N_8290,N_7040,N_7305);
or U8291 (N_8291,N_5160,N_5194);
nor U8292 (N_8292,N_7070,N_7276);
nor U8293 (N_8293,N_7479,N_6583);
nand U8294 (N_8294,N_5686,N_5869);
nand U8295 (N_8295,N_7399,N_6896);
xor U8296 (N_8296,N_7314,N_7445);
and U8297 (N_8297,N_5267,N_6829);
nor U8298 (N_8298,N_5622,N_5150);
or U8299 (N_8299,N_6676,N_7062);
nand U8300 (N_8300,N_7226,N_5384);
nand U8301 (N_8301,N_5526,N_6162);
nand U8302 (N_8302,N_7396,N_6104);
or U8303 (N_8303,N_5746,N_5239);
and U8304 (N_8304,N_6111,N_5148);
or U8305 (N_8305,N_6467,N_6344);
or U8306 (N_8306,N_5621,N_5553);
xnor U8307 (N_8307,N_6415,N_5904);
and U8308 (N_8308,N_6705,N_6976);
nor U8309 (N_8309,N_6887,N_6224);
nand U8310 (N_8310,N_7122,N_5258);
xnor U8311 (N_8311,N_7454,N_6221);
nand U8312 (N_8312,N_6826,N_7295);
nand U8313 (N_8313,N_7347,N_7353);
and U8314 (N_8314,N_6478,N_6521);
nor U8315 (N_8315,N_6925,N_7459);
nor U8316 (N_8316,N_6861,N_7383);
or U8317 (N_8317,N_7455,N_6731);
nor U8318 (N_8318,N_5498,N_5572);
or U8319 (N_8319,N_7344,N_5596);
nor U8320 (N_8320,N_5108,N_6422);
nand U8321 (N_8321,N_5260,N_5159);
or U8322 (N_8322,N_6986,N_6390);
nor U8323 (N_8323,N_7370,N_7046);
xor U8324 (N_8324,N_5305,N_6234);
xor U8325 (N_8325,N_5124,N_6056);
nor U8326 (N_8326,N_6022,N_6493);
nand U8327 (N_8327,N_6758,N_5205);
or U8328 (N_8328,N_7310,N_7110);
nand U8329 (N_8329,N_5110,N_6806);
and U8330 (N_8330,N_5230,N_7048);
nand U8331 (N_8331,N_5242,N_6751);
or U8332 (N_8332,N_6926,N_7327);
xor U8333 (N_8333,N_6238,N_6883);
and U8334 (N_8334,N_5560,N_6428);
nor U8335 (N_8335,N_6733,N_6469);
nand U8336 (N_8336,N_7166,N_5043);
nor U8337 (N_8337,N_5191,N_5778);
xnor U8338 (N_8338,N_7287,N_6564);
nor U8339 (N_8339,N_6735,N_5516);
nand U8340 (N_8340,N_5667,N_6228);
nor U8341 (N_8341,N_5616,N_6072);
and U8342 (N_8342,N_6531,N_6182);
or U8343 (N_8343,N_5740,N_5072);
nor U8344 (N_8344,N_5087,N_7214);
nand U8345 (N_8345,N_6951,N_6279);
and U8346 (N_8346,N_5086,N_5485);
xnor U8347 (N_8347,N_5090,N_5354);
or U8348 (N_8348,N_7260,N_6434);
and U8349 (N_8349,N_5035,N_5623);
or U8350 (N_8350,N_6278,N_7044);
xor U8351 (N_8351,N_5917,N_6943);
xnor U8352 (N_8352,N_5263,N_6128);
nor U8353 (N_8353,N_7279,N_7376);
and U8354 (N_8354,N_7067,N_7171);
or U8355 (N_8355,N_5318,N_7460);
nand U8356 (N_8356,N_5211,N_6559);
or U8357 (N_8357,N_5512,N_5197);
nor U8358 (N_8358,N_6324,N_5085);
and U8359 (N_8359,N_5955,N_6251);
nand U8360 (N_8360,N_5183,N_6715);
xnor U8361 (N_8361,N_7181,N_5670);
nor U8362 (N_8362,N_6803,N_5712);
nor U8363 (N_8363,N_6847,N_5721);
nor U8364 (N_8364,N_7051,N_5573);
nand U8365 (N_8365,N_7231,N_5123);
and U8366 (N_8366,N_5798,N_6759);
and U8367 (N_8367,N_5071,N_5298);
xnor U8368 (N_8368,N_5963,N_6811);
xnor U8369 (N_8369,N_6724,N_6929);
and U8370 (N_8370,N_6892,N_6323);
and U8371 (N_8371,N_6337,N_6429);
or U8372 (N_8372,N_6075,N_5617);
and U8373 (N_8373,N_6899,N_7159);
nor U8374 (N_8374,N_5240,N_5014);
or U8375 (N_8375,N_5841,N_7273);
nand U8376 (N_8376,N_5660,N_5466);
or U8377 (N_8377,N_5347,N_6639);
and U8378 (N_8378,N_7361,N_7114);
and U8379 (N_8379,N_6689,N_6588);
and U8380 (N_8380,N_6546,N_5220);
nor U8381 (N_8381,N_5369,N_5089);
or U8382 (N_8382,N_6983,N_6619);
nor U8383 (N_8383,N_5993,N_5961);
nand U8384 (N_8384,N_7436,N_7083);
xnor U8385 (N_8385,N_6858,N_6959);
xnor U8386 (N_8386,N_6418,N_6928);
nor U8387 (N_8387,N_6321,N_5651);
or U8388 (N_8388,N_5273,N_6475);
or U8389 (N_8389,N_6700,N_7268);
and U8390 (N_8390,N_7397,N_6148);
xor U8391 (N_8391,N_6370,N_7393);
nand U8392 (N_8392,N_7136,N_6604);
xnor U8393 (N_8393,N_6553,N_7089);
nor U8394 (N_8394,N_5237,N_7081);
nor U8395 (N_8395,N_5256,N_5179);
nand U8396 (N_8396,N_5093,N_6409);
or U8397 (N_8397,N_6836,N_5926);
nor U8398 (N_8398,N_6631,N_5827);
xnor U8399 (N_8399,N_6454,N_5348);
nor U8400 (N_8400,N_7315,N_5009);
nand U8401 (N_8401,N_6612,N_5397);
nand U8402 (N_8402,N_7356,N_6195);
or U8403 (N_8403,N_5892,N_6084);
nand U8404 (N_8404,N_7300,N_6595);
xnor U8405 (N_8405,N_5375,N_6709);
nand U8406 (N_8406,N_5925,N_6581);
or U8407 (N_8407,N_7009,N_5388);
and U8408 (N_8408,N_5460,N_6686);
xor U8409 (N_8409,N_7105,N_6574);
or U8410 (N_8410,N_7458,N_7178);
and U8411 (N_8411,N_6175,N_5495);
nand U8412 (N_8412,N_5603,N_6823);
nand U8413 (N_8413,N_7154,N_7381);
or U8414 (N_8414,N_7373,N_7340);
and U8415 (N_8415,N_7413,N_7085);
and U8416 (N_8416,N_5646,N_5903);
nand U8417 (N_8417,N_5493,N_5792);
nand U8418 (N_8418,N_5131,N_7257);
and U8419 (N_8419,N_6954,N_5238);
or U8420 (N_8420,N_5590,N_5155);
or U8421 (N_8421,N_7474,N_5716);
nor U8422 (N_8422,N_5119,N_5808);
and U8423 (N_8423,N_6273,N_6890);
nor U8424 (N_8424,N_7238,N_6615);
or U8425 (N_8425,N_6057,N_5277);
nor U8426 (N_8426,N_6082,N_7306);
or U8427 (N_8427,N_7211,N_6629);
nand U8428 (N_8428,N_5453,N_7191);
nor U8429 (N_8429,N_6071,N_5811);
xor U8430 (N_8430,N_6662,N_7218);
or U8431 (N_8431,N_5196,N_5476);
xor U8432 (N_8432,N_6624,N_6134);
and U8433 (N_8433,N_5698,N_6247);
and U8434 (N_8434,N_6262,N_7053);
nor U8435 (N_8435,N_6436,N_7022);
nor U8436 (N_8436,N_5431,N_7033);
and U8437 (N_8437,N_7317,N_6466);
nand U8438 (N_8438,N_6725,N_6670);
xnor U8439 (N_8439,N_5715,N_5370);
xor U8440 (N_8440,N_6745,N_5472);
nor U8441 (N_8441,N_6058,N_5818);
xnor U8442 (N_8442,N_7180,N_7466);
or U8443 (N_8443,N_5333,N_7407);
and U8444 (N_8444,N_5680,N_5037);
or U8445 (N_8445,N_6766,N_6975);
or U8446 (N_8446,N_5924,N_6298);
and U8447 (N_8447,N_5034,N_7185);
xnor U8448 (N_8448,N_6240,N_5593);
and U8449 (N_8449,N_6419,N_6924);
or U8450 (N_8450,N_5511,N_5562);
nand U8451 (N_8451,N_6796,N_6565);
or U8452 (N_8452,N_7063,N_5943);
xor U8453 (N_8453,N_5845,N_5815);
and U8454 (N_8454,N_5969,N_6187);
nor U8455 (N_8455,N_5911,N_6295);
and U8456 (N_8456,N_5985,N_5459);
xor U8457 (N_8457,N_5996,N_5140);
nor U8458 (N_8458,N_5945,N_6190);
or U8459 (N_8459,N_6108,N_6834);
xor U8460 (N_8460,N_6718,N_7427);
and U8461 (N_8461,N_6440,N_5103);
xor U8462 (N_8462,N_7168,N_6579);
nor U8463 (N_8463,N_6516,N_6754);
or U8464 (N_8464,N_6771,N_7491);
and U8465 (N_8465,N_5631,N_6432);
and U8466 (N_8466,N_5134,N_6302);
and U8467 (N_8467,N_5600,N_7462);
nor U8468 (N_8468,N_5116,N_5745);
or U8469 (N_8469,N_5019,N_5822);
nand U8470 (N_8470,N_7212,N_5835);
nor U8471 (N_8471,N_7101,N_6438);
xnor U8472 (N_8472,N_6944,N_5300);
nor U8473 (N_8473,N_7416,N_7096);
nor U8474 (N_8474,N_5415,N_6431);
nand U8475 (N_8475,N_5314,N_6325);
and U8476 (N_8476,N_6597,N_6144);
and U8477 (N_8477,N_6087,N_6848);
or U8478 (N_8478,N_5365,N_5216);
nand U8479 (N_8479,N_5438,N_5971);
or U8480 (N_8480,N_5984,N_7251);
nor U8481 (N_8481,N_5243,N_7333);
nand U8482 (N_8482,N_6383,N_7292);
nand U8483 (N_8483,N_5233,N_7055);
nor U8484 (N_8484,N_5377,N_5612);
nor U8485 (N_8485,N_7388,N_6819);
or U8486 (N_8486,N_6226,N_7223);
nor U8487 (N_8487,N_6198,N_5161);
or U8488 (N_8488,N_6266,N_5195);
nor U8489 (N_8489,N_5046,N_7034);
xnor U8490 (N_8490,N_5292,N_6317);
nand U8491 (N_8491,N_6427,N_5464);
or U8492 (N_8492,N_6105,N_5654);
or U8493 (N_8493,N_6129,N_6025);
and U8494 (N_8494,N_6916,N_6416);
and U8495 (N_8495,N_6001,N_5428);
xor U8496 (N_8496,N_5565,N_5884);
or U8497 (N_8497,N_5935,N_5302);
xor U8498 (N_8498,N_6730,N_7098);
nand U8499 (N_8499,N_6651,N_5789);
nand U8500 (N_8500,N_6241,N_6308);
and U8501 (N_8501,N_5703,N_5563);
nor U8502 (N_8502,N_5678,N_5594);
nor U8503 (N_8503,N_5253,N_7465);
nor U8504 (N_8504,N_6566,N_7346);
nor U8505 (N_8505,N_5771,N_5247);
xnor U8506 (N_8506,N_5569,N_6798);
or U8507 (N_8507,N_7259,N_5427);
or U8508 (N_8508,N_5021,N_7489);
and U8509 (N_8509,N_5349,N_7250);
or U8510 (N_8510,N_7208,N_7198);
or U8511 (N_8511,N_7036,N_5718);
nor U8512 (N_8512,N_5363,N_5053);
xnor U8513 (N_8513,N_5421,N_6018);
or U8514 (N_8514,N_7151,N_7481);
and U8515 (N_8515,N_6593,N_6272);
and U8516 (N_8516,N_7194,N_5983);
and U8517 (N_8517,N_5188,N_6875);
or U8518 (N_8518,N_6849,N_6504);
and U8519 (N_8519,N_5824,N_6679);
and U8520 (N_8520,N_5666,N_6441);
and U8521 (N_8521,N_5793,N_6318);
and U8522 (N_8522,N_7010,N_5359);
and U8523 (N_8523,N_5416,N_6613);
xor U8524 (N_8524,N_5418,N_5405);
nor U8525 (N_8525,N_5047,N_5001);
or U8526 (N_8526,N_5507,N_7324);
nand U8527 (N_8527,N_7042,N_6054);
nor U8528 (N_8528,N_6027,N_5200);
and U8529 (N_8529,N_6062,N_5308);
nor U8530 (N_8530,N_5177,N_5589);
xor U8531 (N_8531,N_6150,N_6852);
xnor U8532 (N_8532,N_5092,N_6503);
or U8533 (N_8533,N_5873,N_6359);
or U8534 (N_8534,N_6756,N_5245);
nor U8535 (N_8535,N_6673,N_5129);
and U8536 (N_8536,N_5648,N_5311);
xnor U8537 (N_8537,N_5236,N_6616);
and U8538 (N_8538,N_6879,N_6489);
xnor U8539 (N_8539,N_5912,N_6149);
or U8540 (N_8540,N_5545,N_6352);
or U8541 (N_8541,N_7420,N_6028);
or U8542 (N_8542,N_5865,N_5619);
and U8543 (N_8543,N_6392,N_6329);
nand U8544 (N_8544,N_5995,N_6665);
nor U8545 (N_8545,N_6303,N_5656);
xor U8546 (N_8546,N_6741,N_6004);
and U8547 (N_8547,N_7135,N_5652);
xor U8548 (N_8548,N_6293,N_6451);
xnor U8549 (N_8549,N_7354,N_7409);
nand U8550 (N_8550,N_6459,N_6214);
xor U8551 (N_8551,N_7461,N_7004);
nand U8552 (N_8552,N_5655,N_5288);
xor U8553 (N_8553,N_6729,N_6578);
nand U8554 (N_8554,N_6141,N_6777);
nand U8555 (N_8555,N_6109,N_5469);
or U8556 (N_8556,N_7398,N_7484);
xnor U8557 (N_8557,N_5011,N_5900);
and U8558 (N_8558,N_7330,N_6642);
xor U8559 (N_8559,N_6544,N_6843);
or U8560 (N_8560,N_6085,N_6030);
and U8561 (N_8561,N_5940,N_6596);
or U8562 (N_8562,N_5682,N_6282);
nand U8563 (N_8563,N_6902,N_6186);
nand U8564 (N_8564,N_5566,N_5805);
nand U8565 (N_8565,N_7068,N_7030);
or U8566 (N_8566,N_7097,N_5902);
nor U8567 (N_8567,N_6994,N_5064);
nor U8568 (N_8568,N_6502,N_7074);
nand U8569 (N_8569,N_7303,N_6496);
nand U8570 (N_8570,N_5860,N_7184);
nor U8571 (N_8571,N_6185,N_6341);
xor U8572 (N_8572,N_7002,N_5389);
or U8573 (N_8573,N_6360,N_6757);
or U8574 (N_8574,N_7452,N_7497);
xnor U8575 (N_8575,N_6526,N_5837);
nand U8576 (N_8576,N_5257,N_7073);
and U8577 (N_8577,N_6012,N_5883);
nand U8578 (N_8578,N_6477,N_6330);
and U8579 (N_8579,N_5268,N_7093);
or U8580 (N_8580,N_7422,N_5357);
and U8581 (N_8581,N_6501,N_5036);
nand U8582 (N_8582,N_5435,N_6920);
or U8583 (N_8583,N_6965,N_6481);
xnor U8584 (N_8584,N_6202,N_5732);
or U8585 (N_8585,N_6268,N_5056);
xnor U8586 (N_8586,N_6286,N_5772);
or U8587 (N_8587,N_6277,N_6590);
and U8588 (N_8588,N_6534,N_7225);
and U8589 (N_8589,N_7244,N_5395);
xnor U8590 (N_8590,N_6810,N_7364);
or U8591 (N_8591,N_6408,N_6263);
nor U8592 (N_8592,N_5480,N_5706);
nor U8593 (N_8593,N_5748,N_7011);
nor U8594 (N_8594,N_6433,N_5206);
nand U8595 (N_8595,N_6217,N_6738);
nand U8596 (N_8596,N_5162,N_6139);
xor U8597 (N_8597,N_7013,N_5614);
nand U8598 (N_8598,N_7024,N_6367);
and U8599 (N_8599,N_5186,N_5998);
nor U8600 (N_8600,N_6844,N_7403);
nor U8601 (N_8601,N_6540,N_7430);
xnor U8602 (N_8602,N_6281,N_7041);
xnor U8603 (N_8603,N_6119,N_5738);
nor U8604 (N_8604,N_5052,N_6364);
and U8605 (N_8605,N_6539,N_5117);
or U8606 (N_8606,N_5847,N_6373);
xnor U8607 (N_8607,N_5187,N_5515);
or U8608 (N_8608,N_5520,N_6979);
nand U8609 (N_8609,N_7161,N_5272);
or U8610 (N_8610,N_7125,N_5736);
nand U8611 (N_8611,N_6179,N_5345);
or U8612 (N_8612,N_5478,N_7078);
nor U8613 (N_8613,N_7322,N_6068);
xnor U8614 (N_8614,N_6981,N_5412);
nor U8615 (N_8615,N_6992,N_6659);
or U8616 (N_8616,N_7385,N_5674);
nand U8617 (N_8617,N_5701,N_6421);
and U8618 (N_8618,N_5997,N_5081);
xor U8619 (N_8619,N_6655,N_6142);
nor U8620 (N_8620,N_6555,N_6687);
nor U8621 (N_8621,N_5559,N_6158);
or U8622 (N_8622,N_7339,N_5497);
and U8623 (N_8623,N_7176,N_5030);
nor U8624 (N_8624,N_5625,N_6387);
nor U8625 (N_8625,N_6029,N_7258);
or U8626 (N_8626,N_6401,N_5038);
and U8627 (N_8627,N_5337,N_7477);
nand U8628 (N_8628,N_6533,N_6814);
and U8629 (N_8629,N_5094,N_6537);
or U8630 (N_8630,N_5334,N_5541);
nor U8631 (N_8631,N_7003,N_6585);
xor U8632 (N_8632,N_5422,N_5169);
nand U8633 (N_8633,N_5724,N_7299);
nand U8634 (N_8634,N_5396,N_6635);
and U8635 (N_8635,N_6166,N_5538);
nor U8636 (N_8636,N_6386,N_6820);
xnor U8637 (N_8637,N_5413,N_5190);
xnor U8638 (N_8638,N_7134,N_6969);
and U8639 (N_8639,N_5282,N_5371);
nand U8640 (N_8640,N_6335,N_6035);
or U8641 (N_8641,N_5234,N_6750);
xnor U8642 (N_8642,N_7372,N_6199);
or U8643 (N_8643,N_5387,N_6032);
xor U8644 (N_8644,N_5020,N_7438);
or U8645 (N_8645,N_5885,N_5958);
and U8646 (N_8646,N_6712,N_7005);
xor U8647 (N_8647,N_5213,N_6081);
xor U8648 (N_8648,N_7215,N_5813);
nand U8649 (N_8649,N_7371,N_6680);
xnor U8650 (N_8650,N_5269,N_6512);
nor U8651 (N_8651,N_6769,N_7446);
nor U8652 (N_8652,N_5613,N_5532);
nor U8653 (N_8653,N_5918,N_6702);
or U8654 (N_8654,N_5965,N_7019);
or U8655 (N_8655,N_5941,N_5979);
or U8656 (N_8656,N_6236,N_6174);
nand U8657 (N_8657,N_7220,N_5362);
nor U8658 (N_8658,N_6461,N_5032);
or U8659 (N_8659,N_5307,N_6554);
nand U8660 (N_8660,N_5166,N_5536);
and U8661 (N_8661,N_5502,N_7390);
or U8662 (N_8662,N_7047,N_5754);
nand U8663 (N_8663,N_5784,N_5509);
nand U8664 (N_8664,N_6880,N_6692);
nor U8665 (N_8665,N_6125,N_6523);
and U8666 (N_8666,N_5855,N_7139);
nor U8667 (N_8667,N_5549,N_5714);
nand U8668 (N_8668,N_7132,N_7433);
or U8669 (N_8669,N_5611,N_6313);
or U8670 (N_8670,N_7103,N_7307);
nor U8671 (N_8671,N_6412,N_6669);
and U8672 (N_8672,N_7302,N_6630);
nand U8673 (N_8673,N_5554,N_6404);
xor U8674 (N_8674,N_6971,N_5896);
xor U8675 (N_8675,N_5471,N_6391);
or U8676 (N_8676,N_6586,N_5681);
or U8677 (N_8677,N_6945,N_5717);
xnor U8678 (N_8678,N_6167,N_6151);
nor U8679 (N_8679,N_6668,N_6237);
nand U8680 (N_8680,N_7278,N_5255);
nor U8681 (N_8681,N_5054,N_5445);
or U8682 (N_8682,N_6107,N_5467);
nand U8683 (N_8683,N_6299,N_6786);
xor U8684 (N_8684,N_5217,N_5690);
nor U8685 (N_8685,N_7483,N_6868);
nor U8686 (N_8686,N_6990,N_6793);
nand U8687 (N_8687,N_5259,N_6645);
xnor U8688 (N_8688,N_6499,N_7049);
nand U8689 (N_8689,N_5173,N_6643);
and U8690 (N_8690,N_5956,N_5006);
xor U8691 (N_8691,N_5378,N_6394);
nand U8692 (N_8692,N_5364,N_7012);
nand U8693 (N_8693,N_5024,N_5552);
xnor U8694 (N_8694,N_6482,N_6336);
xnor U8695 (N_8695,N_6163,N_5887);
and U8696 (N_8696,N_6781,N_6116);
and U8697 (N_8697,N_6339,N_6040);
and U8698 (N_8698,N_7366,N_5513);
or U8699 (N_8699,N_5960,N_5876);
xor U8700 (N_8700,N_5647,N_5629);
xor U8701 (N_8701,N_6465,N_5723);
nor U8702 (N_8702,N_5067,N_6984);
nand U8703 (N_8703,N_5966,N_5833);
and U8704 (N_8704,N_5042,N_5741);
nor U8705 (N_8705,N_6838,N_7152);
xor U8706 (N_8706,N_7336,N_6815);
nor U8707 (N_8707,N_7092,N_7076);
nand U8708 (N_8708,N_5293,N_7426);
nand U8709 (N_8709,N_5346,N_5644);
or U8710 (N_8710,N_6406,N_6804);
or U8711 (N_8711,N_7411,N_7274);
and U8712 (N_8712,N_5400,N_7241);
nand U8713 (N_8713,N_6785,N_7149);
and U8714 (N_8714,N_6490,N_6505);
and U8715 (N_8715,N_6956,N_6514);
or U8716 (N_8716,N_7021,N_6423);
nor U8717 (N_8717,N_6832,N_6208);
or U8718 (N_8718,N_6727,N_7188);
and U8719 (N_8719,N_6833,N_5490);
or U8720 (N_8720,N_6517,N_6088);
or U8721 (N_8721,N_6047,N_6801);
and U8722 (N_8722,N_6309,N_7158);
and U8723 (N_8723,N_6289,N_6285);
nor U8724 (N_8724,N_5274,N_5452);
nand U8725 (N_8725,N_6201,N_5294);
or U8726 (N_8726,N_5774,N_6611);
nor U8727 (N_8727,N_7355,N_6288);
nand U8728 (N_8728,N_6857,N_7202);
xnor U8729 (N_8729,N_7057,N_5404);
nor U8730 (N_8730,N_6551,N_5558);
nor U8731 (N_8731,N_5864,N_6420);
nor U8732 (N_8732,N_5891,N_6608);
or U8733 (N_8733,N_6121,N_6600);
and U8734 (N_8734,N_5279,N_6894);
nor U8735 (N_8735,N_6931,N_5673);
nor U8736 (N_8736,N_5609,N_5937);
or U8737 (N_8737,N_7380,N_6532);
nor U8738 (N_8738,N_6261,N_6996);
and U8739 (N_8739,N_6039,N_6003);
xor U8740 (N_8740,N_5218,N_7319);
xor U8741 (N_8741,N_6515,N_6696);
xnor U8742 (N_8742,N_6779,N_7437);
and U8743 (N_8743,N_6348,N_6901);
nand U8744 (N_8744,N_5127,N_7203);
and U8745 (N_8745,N_5727,N_6932);
xnor U8746 (N_8746,N_7378,N_5756);
nand U8747 (N_8747,N_7118,N_5657);
nor U8748 (N_8748,N_5574,N_6770);
xor U8749 (N_8749,N_7177,N_5992);
nor U8750 (N_8750,N_5129,N_6735);
and U8751 (N_8751,N_7269,N_6099);
and U8752 (N_8752,N_5908,N_6464);
nand U8753 (N_8753,N_6870,N_6991);
xnor U8754 (N_8754,N_5097,N_7342);
xor U8755 (N_8755,N_5656,N_6026);
nor U8756 (N_8756,N_6145,N_6401);
nand U8757 (N_8757,N_5943,N_5545);
and U8758 (N_8758,N_6789,N_5787);
nor U8759 (N_8759,N_6087,N_7293);
or U8760 (N_8760,N_5719,N_6924);
and U8761 (N_8761,N_6427,N_6368);
nor U8762 (N_8762,N_6429,N_6215);
nand U8763 (N_8763,N_5575,N_6557);
nand U8764 (N_8764,N_7018,N_6335);
nand U8765 (N_8765,N_6226,N_5705);
nor U8766 (N_8766,N_6144,N_5324);
xor U8767 (N_8767,N_6408,N_6322);
or U8768 (N_8768,N_7409,N_6092);
nand U8769 (N_8769,N_5838,N_6971);
and U8770 (N_8770,N_7180,N_6235);
or U8771 (N_8771,N_7380,N_6540);
nand U8772 (N_8772,N_7060,N_6007);
xor U8773 (N_8773,N_7303,N_5953);
or U8774 (N_8774,N_6563,N_5961);
nor U8775 (N_8775,N_6913,N_5848);
or U8776 (N_8776,N_6164,N_5712);
nand U8777 (N_8777,N_5865,N_5442);
nor U8778 (N_8778,N_6881,N_5252);
nor U8779 (N_8779,N_6598,N_5054);
nor U8780 (N_8780,N_5256,N_6318);
nand U8781 (N_8781,N_6899,N_5738);
nor U8782 (N_8782,N_5916,N_5167);
nand U8783 (N_8783,N_5064,N_6320);
xor U8784 (N_8784,N_5119,N_6841);
or U8785 (N_8785,N_6410,N_5341);
or U8786 (N_8786,N_6784,N_5976);
xor U8787 (N_8787,N_5457,N_6144);
nor U8788 (N_8788,N_5662,N_6322);
xor U8789 (N_8789,N_6964,N_6307);
or U8790 (N_8790,N_5249,N_5637);
nor U8791 (N_8791,N_5506,N_5088);
or U8792 (N_8792,N_6256,N_7349);
or U8793 (N_8793,N_7148,N_5584);
nand U8794 (N_8794,N_6118,N_7237);
and U8795 (N_8795,N_5064,N_5814);
nand U8796 (N_8796,N_6890,N_6477);
and U8797 (N_8797,N_7445,N_5207);
nor U8798 (N_8798,N_5060,N_6170);
or U8799 (N_8799,N_6637,N_5225);
or U8800 (N_8800,N_6109,N_6695);
or U8801 (N_8801,N_5649,N_6982);
xor U8802 (N_8802,N_6218,N_6512);
xnor U8803 (N_8803,N_6831,N_6456);
nand U8804 (N_8804,N_5724,N_6790);
and U8805 (N_8805,N_5470,N_5883);
nor U8806 (N_8806,N_5860,N_5068);
nor U8807 (N_8807,N_5584,N_7421);
nor U8808 (N_8808,N_6052,N_6000);
nand U8809 (N_8809,N_5435,N_6233);
and U8810 (N_8810,N_5381,N_5269);
xnor U8811 (N_8811,N_6327,N_5334);
nor U8812 (N_8812,N_5023,N_5556);
or U8813 (N_8813,N_7151,N_7220);
nor U8814 (N_8814,N_6789,N_5096);
nand U8815 (N_8815,N_5751,N_5521);
and U8816 (N_8816,N_5091,N_6646);
nor U8817 (N_8817,N_5644,N_6559);
nand U8818 (N_8818,N_6550,N_5814);
or U8819 (N_8819,N_7215,N_6603);
or U8820 (N_8820,N_6586,N_6862);
xor U8821 (N_8821,N_5556,N_5092);
or U8822 (N_8822,N_6129,N_6348);
nor U8823 (N_8823,N_5168,N_6651);
nand U8824 (N_8824,N_6667,N_7400);
and U8825 (N_8825,N_5430,N_6955);
or U8826 (N_8826,N_7179,N_5696);
xor U8827 (N_8827,N_7430,N_5448);
nor U8828 (N_8828,N_6964,N_5997);
and U8829 (N_8829,N_6851,N_6314);
and U8830 (N_8830,N_5052,N_6939);
and U8831 (N_8831,N_6458,N_7202);
xor U8832 (N_8832,N_7183,N_5496);
nand U8833 (N_8833,N_5843,N_6322);
and U8834 (N_8834,N_7253,N_7134);
or U8835 (N_8835,N_6506,N_7492);
and U8836 (N_8836,N_5747,N_7039);
or U8837 (N_8837,N_5074,N_6898);
and U8838 (N_8838,N_6952,N_5261);
or U8839 (N_8839,N_6956,N_6243);
xor U8840 (N_8840,N_7317,N_6031);
nor U8841 (N_8841,N_7052,N_6947);
and U8842 (N_8842,N_5880,N_6604);
nand U8843 (N_8843,N_6895,N_5331);
nor U8844 (N_8844,N_5475,N_5534);
nor U8845 (N_8845,N_5607,N_5612);
or U8846 (N_8846,N_7082,N_5697);
and U8847 (N_8847,N_5409,N_5320);
xor U8848 (N_8848,N_5307,N_5812);
xor U8849 (N_8849,N_6452,N_5478);
and U8850 (N_8850,N_6627,N_7292);
nor U8851 (N_8851,N_7209,N_5317);
nand U8852 (N_8852,N_5262,N_5166);
or U8853 (N_8853,N_5197,N_7311);
xnor U8854 (N_8854,N_6478,N_7266);
or U8855 (N_8855,N_6159,N_6480);
xnor U8856 (N_8856,N_7017,N_6646);
or U8857 (N_8857,N_5508,N_5448);
and U8858 (N_8858,N_5140,N_6282);
and U8859 (N_8859,N_5594,N_6069);
nor U8860 (N_8860,N_6216,N_6215);
nand U8861 (N_8861,N_6290,N_6573);
nor U8862 (N_8862,N_7175,N_6008);
nor U8863 (N_8863,N_5260,N_5821);
nand U8864 (N_8864,N_5939,N_6316);
or U8865 (N_8865,N_6186,N_5445);
and U8866 (N_8866,N_5448,N_6265);
or U8867 (N_8867,N_7216,N_5088);
or U8868 (N_8868,N_5663,N_6949);
xor U8869 (N_8869,N_6100,N_6231);
or U8870 (N_8870,N_5156,N_7295);
xnor U8871 (N_8871,N_6503,N_6563);
or U8872 (N_8872,N_5817,N_6048);
nand U8873 (N_8873,N_7284,N_5720);
nor U8874 (N_8874,N_6284,N_5776);
or U8875 (N_8875,N_5102,N_6057);
and U8876 (N_8876,N_5487,N_7464);
xor U8877 (N_8877,N_5258,N_6548);
nor U8878 (N_8878,N_7491,N_6888);
nor U8879 (N_8879,N_5695,N_6363);
or U8880 (N_8880,N_7379,N_5273);
nand U8881 (N_8881,N_7149,N_6918);
xor U8882 (N_8882,N_5894,N_6086);
or U8883 (N_8883,N_5579,N_6805);
xor U8884 (N_8884,N_5069,N_5686);
and U8885 (N_8885,N_7393,N_6589);
xor U8886 (N_8886,N_7447,N_6039);
xnor U8887 (N_8887,N_6899,N_7458);
and U8888 (N_8888,N_6651,N_5769);
nor U8889 (N_8889,N_7083,N_6433);
nand U8890 (N_8890,N_5090,N_5590);
nand U8891 (N_8891,N_6859,N_7447);
and U8892 (N_8892,N_6947,N_5774);
or U8893 (N_8893,N_5280,N_6003);
and U8894 (N_8894,N_7119,N_7060);
or U8895 (N_8895,N_6586,N_5694);
and U8896 (N_8896,N_6436,N_5281);
and U8897 (N_8897,N_6683,N_6187);
or U8898 (N_8898,N_5951,N_5668);
nand U8899 (N_8899,N_5143,N_6128);
nor U8900 (N_8900,N_5838,N_5458);
and U8901 (N_8901,N_7479,N_7463);
or U8902 (N_8902,N_6965,N_5643);
xnor U8903 (N_8903,N_5521,N_5987);
nand U8904 (N_8904,N_5951,N_6457);
nand U8905 (N_8905,N_5325,N_7255);
and U8906 (N_8906,N_6296,N_5150);
nand U8907 (N_8907,N_6592,N_6273);
or U8908 (N_8908,N_5964,N_6064);
or U8909 (N_8909,N_6579,N_5584);
or U8910 (N_8910,N_6441,N_6004);
nor U8911 (N_8911,N_5622,N_7285);
xnor U8912 (N_8912,N_7200,N_6004);
nand U8913 (N_8913,N_5299,N_5968);
nor U8914 (N_8914,N_6047,N_5250);
or U8915 (N_8915,N_5007,N_5520);
and U8916 (N_8916,N_7261,N_5284);
nor U8917 (N_8917,N_5192,N_6573);
nor U8918 (N_8918,N_6145,N_6712);
nand U8919 (N_8919,N_5964,N_7034);
or U8920 (N_8920,N_7287,N_6616);
or U8921 (N_8921,N_7281,N_7420);
or U8922 (N_8922,N_7057,N_7416);
xnor U8923 (N_8923,N_6527,N_6811);
and U8924 (N_8924,N_6735,N_7190);
nor U8925 (N_8925,N_5209,N_6489);
nor U8926 (N_8926,N_6340,N_5966);
xnor U8927 (N_8927,N_6375,N_7358);
or U8928 (N_8928,N_6772,N_5286);
nor U8929 (N_8929,N_6718,N_7058);
nand U8930 (N_8930,N_5074,N_6312);
nor U8931 (N_8931,N_6797,N_7279);
nor U8932 (N_8932,N_7025,N_5749);
nor U8933 (N_8933,N_5366,N_6128);
xor U8934 (N_8934,N_5758,N_5751);
nor U8935 (N_8935,N_6872,N_5712);
and U8936 (N_8936,N_5923,N_6483);
or U8937 (N_8937,N_6526,N_7226);
nor U8938 (N_8938,N_6064,N_5726);
xnor U8939 (N_8939,N_5722,N_6794);
xnor U8940 (N_8940,N_6726,N_7215);
nand U8941 (N_8941,N_6800,N_5165);
or U8942 (N_8942,N_6158,N_6761);
xor U8943 (N_8943,N_7341,N_7081);
nand U8944 (N_8944,N_5817,N_7219);
nand U8945 (N_8945,N_6081,N_6629);
xnor U8946 (N_8946,N_6391,N_6990);
nand U8947 (N_8947,N_5926,N_6456);
nor U8948 (N_8948,N_5114,N_6229);
and U8949 (N_8949,N_6457,N_5838);
xnor U8950 (N_8950,N_6607,N_6381);
nor U8951 (N_8951,N_5730,N_5617);
and U8952 (N_8952,N_6251,N_5949);
nor U8953 (N_8953,N_5091,N_6835);
nor U8954 (N_8954,N_6689,N_5067);
and U8955 (N_8955,N_5458,N_6434);
xnor U8956 (N_8956,N_5861,N_7412);
nand U8957 (N_8957,N_6884,N_6286);
xnor U8958 (N_8958,N_7073,N_6957);
xnor U8959 (N_8959,N_5005,N_6667);
nor U8960 (N_8960,N_7104,N_6135);
or U8961 (N_8961,N_6016,N_6973);
xor U8962 (N_8962,N_6189,N_6839);
and U8963 (N_8963,N_6385,N_5106);
nor U8964 (N_8964,N_5370,N_7033);
nor U8965 (N_8965,N_7277,N_5506);
nand U8966 (N_8966,N_7213,N_5924);
nand U8967 (N_8967,N_5967,N_7367);
nand U8968 (N_8968,N_7422,N_5753);
nor U8969 (N_8969,N_6719,N_5177);
or U8970 (N_8970,N_5690,N_6331);
nor U8971 (N_8971,N_6632,N_6082);
and U8972 (N_8972,N_5064,N_6226);
xor U8973 (N_8973,N_5525,N_7203);
or U8974 (N_8974,N_6746,N_5070);
and U8975 (N_8975,N_7118,N_5171);
and U8976 (N_8976,N_6000,N_5426);
and U8977 (N_8977,N_6255,N_6340);
and U8978 (N_8978,N_5255,N_6160);
and U8979 (N_8979,N_5598,N_5898);
nor U8980 (N_8980,N_7059,N_6030);
and U8981 (N_8981,N_6410,N_5023);
nand U8982 (N_8982,N_5416,N_5489);
nand U8983 (N_8983,N_7281,N_6453);
nand U8984 (N_8984,N_6699,N_7451);
and U8985 (N_8985,N_7421,N_5503);
and U8986 (N_8986,N_7291,N_6235);
xor U8987 (N_8987,N_5582,N_5966);
nor U8988 (N_8988,N_6990,N_6835);
nand U8989 (N_8989,N_7276,N_5000);
xor U8990 (N_8990,N_6809,N_6260);
or U8991 (N_8991,N_6457,N_6549);
and U8992 (N_8992,N_7335,N_6863);
nor U8993 (N_8993,N_5708,N_6523);
nor U8994 (N_8994,N_6009,N_7351);
and U8995 (N_8995,N_6016,N_7488);
nand U8996 (N_8996,N_7391,N_7407);
nor U8997 (N_8997,N_6126,N_5736);
or U8998 (N_8998,N_6836,N_6209);
nand U8999 (N_8999,N_7167,N_6999);
nor U9000 (N_9000,N_6459,N_6346);
and U9001 (N_9001,N_5907,N_5398);
nand U9002 (N_9002,N_6956,N_5704);
nor U9003 (N_9003,N_5597,N_7404);
xor U9004 (N_9004,N_6045,N_6368);
or U9005 (N_9005,N_6595,N_6891);
nor U9006 (N_9006,N_5869,N_6113);
nor U9007 (N_9007,N_5448,N_7249);
and U9008 (N_9008,N_6300,N_7437);
and U9009 (N_9009,N_6754,N_7410);
or U9010 (N_9010,N_6226,N_7298);
xnor U9011 (N_9011,N_5327,N_5783);
nand U9012 (N_9012,N_6999,N_5592);
or U9013 (N_9013,N_6781,N_7193);
or U9014 (N_9014,N_7368,N_5208);
nor U9015 (N_9015,N_5495,N_5861);
or U9016 (N_9016,N_6832,N_5102);
nor U9017 (N_9017,N_5174,N_5567);
nor U9018 (N_9018,N_5846,N_5860);
or U9019 (N_9019,N_6034,N_6699);
xnor U9020 (N_9020,N_6006,N_5042);
and U9021 (N_9021,N_5092,N_6870);
nor U9022 (N_9022,N_5999,N_7464);
or U9023 (N_9023,N_6785,N_7090);
nand U9024 (N_9024,N_5959,N_6607);
nand U9025 (N_9025,N_5734,N_6973);
nand U9026 (N_9026,N_6278,N_5172);
nor U9027 (N_9027,N_5978,N_6763);
and U9028 (N_9028,N_5213,N_5468);
nand U9029 (N_9029,N_6696,N_6337);
nor U9030 (N_9030,N_5997,N_6552);
and U9031 (N_9031,N_6020,N_6522);
nand U9032 (N_9032,N_5193,N_7369);
or U9033 (N_9033,N_6503,N_7288);
or U9034 (N_9034,N_7025,N_7053);
nor U9035 (N_9035,N_6834,N_6738);
or U9036 (N_9036,N_6636,N_6758);
and U9037 (N_9037,N_5409,N_7096);
and U9038 (N_9038,N_7319,N_6205);
or U9039 (N_9039,N_6291,N_7385);
nor U9040 (N_9040,N_6692,N_6423);
xnor U9041 (N_9041,N_7025,N_5682);
nor U9042 (N_9042,N_7064,N_5335);
xor U9043 (N_9043,N_6990,N_5002);
nor U9044 (N_9044,N_5715,N_6177);
nor U9045 (N_9045,N_5130,N_6172);
nor U9046 (N_9046,N_6703,N_6575);
xnor U9047 (N_9047,N_5516,N_5847);
nor U9048 (N_9048,N_5790,N_5691);
and U9049 (N_9049,N_6861,N_5877);
and U9050 (N_9050,N_6143,N_5098);
nor U9051 (N_9051,N_6867,N_6151);
or U9052 (N_9052,N_7433,N_7350);
nor U9053 (N_9053,N_7429,N_7234);
and U9054 (N_9054,N_6982,N_6018);
nor U9055 (N_9055,N_5824,N_6179);
and U9056 (N_9056,N_6075,N_5997);
nand U9057 (N_9057,N_5092,N_5831);
nor U9058 (N_9058,N_6066,N_6053);
xor U9059 (N_9059,N_5847,N_5708);
and U9060 (N_9060,N_6800,N_5749);
nand U9061 (N_9061,N_5209,N_5088);
nand U9062 (N_9062,N_5549,N_5342);
nand U9063 (N_9063,N_5615,N_6904);
xnor U9064 (N_9064,N_7212,N_6774);
or U9065 (N_9065,N_6463,N_5550);
nor U9066 (N_9066,N_5630,N_5495);
and U9067 (N_9067,N_6460,N_6717);
or U9068 (N_9068,N_6475,N_5300);
xnor U9069 (N_9069,N_5245,N_6320);
xor U9070 (N_9070,N_7254,N_7229);
nand U9071 (N_9071,N_6967,N_6493);
nor U9072 (N_9072,N_6318,N_6701);
nor U9073 (N_9073,N_6788,N_6646);
or U9074 (N_9074,N_6463,N_7179);
and U9075 (N_9075,N_7471,N_6936);
nor U9076 (N_9076,N_7192,N_6650);
nand U9077 (N_9077,N_7215,N_6591);
or U9078 (N_9078,N_6196,N_5905);
or U9079 (N_9079,N_5167,N_5246);
or U9080 (N_9080,N_6811,N_5186);
nand U9081 (N_9081,N_5561,N_6415);
nor U9082 (N_9082,N_7496,N_7071);
nand U9083 (N_9083,N_6071,N_5943);
nor U9084 (N_9084,N_6474,N_6499);
or U9085 (N_9085,N_5615,N_5854);
nor U9086 (N_9086,N_5445,N_6263);
or U9087 (N_9087,N_5500,N_6711);
and U9088 (N_9088,N_6144,N_6228);
nand U9089 (N_9089,N_5828,N_6647);
xnor U9090 (N_9090,N_6696,N_7011);
and U9091 (N_9091,N_6883,N_5380);
xor U9092 (N_9092,N_6633,N_6218);
nor U9093 (N_9093,N_5536,N_6496);
and U9094 (N_9094,N_7109,N_5617);
or U9095 (N_9095,N_6711,N_6958);
xnor U9096 (N_9096,N_6936,N_5147);
nor U9097 (N_9097,N_5759,N_5822);
nor U9098 (N_9098,N_6633,N_5714);
nand U9099 (N_9099,N_7217,N_5374);
or U9100 (N_9100,N_6615,N_5112);
and U9101 (N_9101,N_6951,N_6881);
xnor U9102 (N_9102,N_5919,N_5065);
and U9103 (N_9103,N_5569,N_6886);
nand U9104 (N_9104,N_7327,N_7304);
or U9105 (N_9105,N_7045,N_7227);
xnor U9106 (N_9106,N_5459,N_6022);
or U9107 (N_9107,N_5150,N_7057);
nand U9108 (N_9108,N_5115,N_5929);
nand U9109 (N_9109,N_6159,N_5432);
and U9110 (N_9110,N_6984,N_6898);
nand U9111 (N_9111,N_7207,N_5856);
xor U9112 (N_9112,N_5759,N_5463);
nand U9113 (N_9113,N_5580,N_6690);
nand U9114 (N_9114,N_5246,N_7172);
or U9115 (N_9115,N_5903,N_5188);
or U9116 (N_9116,N_6574,N_5213);
and U9117 (N_9117,N_6568,N_5871);
xnor U9118 (N_9118,N_7325,N_5052);
and U9119 (N_9119,N_5840,N_5901);
nand U9120 (N_9120,N_6726,N_7183);
nand U9121 (N_9121,N_6601,N_6812);
nor U9122 (N_9122,N_5589,N_6016);
nor U9123 (N_9123,N_6792,N_7458);
and U9124 (N_9124,N_7194,N_5427);
xor U9125 (N_9125,N_7492,N_6544);
and U9126 (N_9126,N_5139,N_5902);
or U9127 (N_9127,N_6214,N_6813);
and U9128 (N_9128,N_7334,N_7489);
and U9129 (N_9129,N_5237,N_5842);
nor U9130 (N_9130,N_5091,N_6733);
nand U9131 (N_9131,N_6198,N_6700);
and U9132 (N_9132,N_5142,N_6153);
xor U9133 (N_9133,N_5885,N_7327);
or U9134 (N_9134,N_7434,N_5793);
xor U9135 (N_9135,N_5575,N_5397);
nand U9136 (N_9136,N_5343,N_5365);
xor U9137 (N_9137,N_5308,N_6259);
nand U9138 (N_9138,N_5144,N_6645);
and U9139 (N_9139,N_6867,N_6266);
or U9140 (N_9140,N_5577,N_5012);
nand U9141 (N_9141,N_5590,N_7188);
and U9142 (N_9142,N_5252,N_5564);
and U9143 (N_9143,N_5728,N_6552);
nand U9144 (N_9144,N_5314,N_5270);
xor U9145 (N_9145,N_6305,N_5767);
xnor U9146 (N_9146,N_5744,N_6410);
or U9147 (N_9147,N_6864,N_6615);
nand U9148 (N_9148,N_7305,N_5393);
and U9149 (N_9149,N_6599,N_6253);
nand U9150 (N_9150,N_5737,N_5309);
nor U9151 (N_9151,N_7340,N_5865);
xor U9152 (N_9152,N_5704,N_6040);
and U9153 (N_9153,N_6316,N_6794);
nor U9154 (N_9154,N_6243,N_6519);
xnor U9155 (N_9155,N_5614,N_5313);
nand U9156 (N_9156,N_6593,N_6322);
nand U9157 (N_9157,N_5795,N_5857);
xor U9158 (N_9158,N_5062,N_5480);
nor U9159 (N_9159,N_6921,N_6581);
and U9160 (N_9160,N_5697,N_6930);
nand U9161 (N_9161,N_6608,N_5864);
or U9162 (N_9162,N_5274,N_7359);
nor U9163 (N_9163,N_6253,N_7287);
xor U9164 (N_9164,N_5549,N_7182);
or U9165 (N_9165,N_5518,N_5260);
or U9166 (N_9166,N_7039,N_6972);
xor U9167 (N_9167,N_6249,N_6959);
nand U9168 (N_9168,N_5105,N_5518);
nand U9169 (N_9169,N_6535,N_5717);
nor U9170 (N_9170,N_5890,N_7104);
or U9171 (N_9171,N_6838,N_6299);
nand U9172 (N_9172,N_6979,N_6498);
xnor U9173 (N_9173,N_5648,N_6779);
nand U9174 (N_9174,N_7051,N_6023);
xor U9175 (N_9175,N_5652,N_6575);
nor U9176 (N_9176,N_7213,N_6889);
nand U9177 (N_9177,N_5673,N_5597);
nor U9178 (N_9178,N_7032,N_5661);
xor U9179 (N_9179,N_7214,N_7057);
xor U9180 (N_9180,N_6743,N_7017);
xor U9181 (N_9181,N_6206,N_5600);
nor U9182 (N_9182,N_7221,N_7430);
nand U9183 (N_9183,N_6961,N_5674);
nor U9184 (N_9184,N_5912,N_5109);
and U9185 (N_9185,N_7483,N_5191);
and U9186 (N_9186,N_5550,N_5941);
and U9187 (N_9187,N_6060,N_6285);
or U9188 (N_9188,N_5444,N_6409);
xor U9189 (N_9189,N_5131,N_5605);
or U9190 (N_9190,N_6317,N_7476);
or U9191 (N_9191,N_6257,N_6318);
and U9192 (N_9192,N_6223,N_5010);
and U9193 (N_9193,N_5350,N_6660);
and U9194 (N_9194,N_7454,N_6085);
xnor U9195 (N_9195,N_5167,N_6460);
and U9196 (N_9196,N_5779,N_5308);
or U9197 (N_9197,N_5615,N_5726);
nor U9198 (N_9198,N_6032,N_5755);
nand U9199 (N_9199,N_6144,N_6157);
and U9200 (N_9200,N_7051,N_5123);
and U9201 (N_9201,N_6759,N_7206);
and U9202 (N_9202,N_6488,N_6923);
or U9203 (N_9203,N_5598,N_5226);
nand U9204 (N_9204,N_6512,N_5339);
nand U9205 (N_9205,N_5791,N_7105);
nand U9206 (N_9206,N_5805,N_5560);
nand U9207 (N_9207,N_6051,N_5559);
or U9208 (N_9208,N_5790,N_5870);
nor U9209 (N_9209,N_6901,N_5722);
nand U9210 (N_9210,N_6552,N_7316);
or U9211 (N_9211,N_6967,N_7232);
and U9212 (N_9212,N_6401,N_6293);
xor U9213 (N_9213,N_7000,N_6441);
nor U9214 (N_9214,N_6926,N_6519);
or U9215 (N_9215,N_6300,N_5968);
and U9216 (N_9216,N_5594,N_5658);
xor U9217 (N_9217,N_5129,N_7189);
or U9218 (N_9218,N_7337,N_6884);
and U9219 (N_9219,N_5667,N_6132);
xor U9220 (N_9220,N_6612,N_6996);
or U9221 (N_9221,N_5348,N_7004);
xnor U9222 (N_9222,N_7445,N_6182);
or U9223 (N_9223,N_6203,N_7330);
or U9224 (N_9224,N_7165,N_5014);
and U9225 (N_9225,N_5556,N_6839);
xnor U9226 (N_9226,N_5773,N_6788);
or U9227 (N_9227,N_5382,N_7120);
xnor U9228 (N_9228,N_7152,N_6110);
and U9229 (N_9229,N_5940,N_5809);
nor U9230 (N_9230,N_7111,N_7141);
nand U9231 (N_9231,N_5416,N_6466);
nand U9232 (N_9232,N_5648,N_5353);
nor U9233 (N_9233,N_6222,N_5669);
nand U9234 (N_9234,N_5493,N_5545);
and U9235 (N_9235,N_5851,N_5219);
or U9236 (N_9236,N_7019,N_6562);
xor U9237 (N_9237,N_5636,N_5978);
xor U9238 (N_9238,N_7333,N_5630);
or U9239 (N_9239,N_5317,N_6045);
xor U9240 (N_9240,N_5824,N_6752);
and U9241 (N_9241,N_6914,N_5715);
nor U9242 (N_9242,N_6798,N_6178);
or U9243 (N_9243,N_5311,N_5712);
nand U9244 (N_9244,N_6575,N_5918);
nand U9245 (N_9245,N_5952,N_7326);
and U9246 (N_9246,N_6691,N_5819);
nor U9247 (N_9247,N_6810,N_5641);
and U9248 (N_9248,N_6778,N_6182);
xnor U9249 (N_9249,N_6079,N_5577);
nor U9250 (N_9250,N_6689,N_5629);
and U9251 (N_9251,N_5357,N_7091);
or U9252 (N_9252,N_7277,N_5886);
nand U9253 (N_9253,N_6606,N_6487);
and U9254 (N_9254,N_5238,N_5196);
nand U9255 (N_9255,N_6693,N_6637);
nand U9256 (N_9256,N_6101,N_6439);
xor U9257 (N_9257,N_7288,N_7285);
or U9258 (N_9258,N_5377,N_7141);
xnor U9259 (N_9259,N_5714,N_5218);
and U9260 (N_9260,N_5381,N_7096);
or U9261 (N_9261,N_5657,N_5563);
or U9262 (N_9262,N_5020,N_5746);
and U9263 (N_9263,N_5129,N_6428);
nor U9264 (N_9264,N_6704,N_7218);
or U9265 (N_9265,N_5277,N_7242);
nor U9266 (N_9266,N_5766,N_6864);
and U9267 (N_9267,N_6294,N_5583);
or U9268 (N_9268,N_6625,N_6411);
nor U9269 (N_9269,N_6711,N_6574);
or U9270 (N_9270,N_7454,N_6239);
nand U9271 (N_9271,N_6638,N_6772);
or U9272 (N_9272,N_6910,N_6816);
and U9273 (N_9273,N_7284,N_7078);
or U9274 (N_9274,N_5144,N_7127);
and U9275 (N_9275,N_5590,N_7283);
or U9276 (N_9276,N_5393,N_7013);
nor U9277 (N_9277,N_5687,N_6103);
and U9278 (N_9278,N_5441,N_5951);
or U9279 (N_9279,N_7334,N_5686);
xor U9280 (N_9280,N_5533,N_5216);
nor U9281 (N_9281,N_7464,N_6034);
or U9282 (N_9282,N_5816,N_6788);
nand U9283 (N_9283,N_6259,N_7102);
nor U9284 (N_9284,N_6285,N_5157);
or U9285 (N_9285,N_7112,N_7261);
or U9286 (N_9286,N_7030,N_5923);
xor U9287 (N_9287,N_5635,N_6730);
and U9288 (N_9288,N_6788,N_7026);
or U9289 (N_9289,N_5025,N_6162);
and U9290 (N_9290,N_6083,N_5145);
nand U9291 (N_9291,N_5223,N_6043);
xor U9292 (N_9292,N_5910,N_7261);
nand U9293 (N_9293,N_6625,N_5432);
xor U9294 (N_9294,N_6376,N_7184);
nand U9295 (N_9295,N_6181,N_5169);
and U9296 (N_9296,N_7378,N_5835);
or U9297 (N_9297,N_5926,N_5126);
and U9298 (N_9298,N_7369,N_5133);
xnor U9299 (N_9299,N_5846,N_7191);
nand U9300 (N_9300,N_7217,N_7142);
or U9301 (N_9301,N_7327,N_6945);
or U9302 (N_9302,N_6221,N_5567);
and U9303 (N_9303,N_6661,N_6588);
nand U9304 (N_9304,N_6615,N_5982);
nor U9305 (N_9305,N_7097,N_6569);
xor U9306 (N_9306,N_7464,N_6137);
or U9307 (N_9307,N_7404,N_6175);
xor U9308 (N_9308,N_5409,N_7072);
or U9309 (N_9309,N_6833,N_5599);
nand U9310 (N_9310,N_6531,N_6102);
nand U9311 (N_9311,N_6523,N_7185);
nor U9312 (N_9312,N_5217,N_5154);
nand U9313 (N_9313,N_5644,N_6996);
or U9314 (N_9314,N_5243,N_6431);
xor U9315 (N_9315,N_5205,N_5652);
nor U9316 (N_9316,N_5784,N_6800);
and U9317 (N_9317,N_5763,N_5395);
nand U9318 (N_9318,N_5282,N_5973);
or U9319 (N_9319,N_6081,N_5239);
or U9320 (N_9320,N_6401,N_7164);
nand U9321 (N_9321,N_5778,N_5477);
and U9322 (N_9322,N_7175,N_6056);
and U9323 (N_9323,N_5428,N_5824);
and U9324 (N_9324,N_6484,N_6279);
nand U9325 (N_9325,N_6455,N_6593);
nand U9326 (N_9326,N_7016,N_6805);
and U9327 (N_9327,N_6489,N_7260);
xnor U9328 (N_9328,N_6553,N_5183);
xor U9329 (N_9329,N_5948,N_6463);
nand U9330 (N_9330,N_5921,N_5521);
or U9331 (N_9331,N_5326,N_6656);
and U9332 (N_9332,N_6820,N_6153);
xor U9333 (N_9333,N_5216,N_5121);
xnor U9334 (N_9334,N_6735,N_5752);
or U9335 (N_9335,N_5769,N_7107);
nor U9336 (N_9336,N_5686,N_5631);
xnor U9337 (N_9337,N_7037,N_5682);
nor U9338 (N_9338,N_6174,N_5884);
or U9339 (N_9339,N_5583,N_5880);
xor U9340 (N_9340,N_5420,N_5765);
and U9341 (N_9341,N_6341,N_5670);
nor U9342 (N_9342,N_7136,N_6365);
nand U9343 (N_9343,N_6112,N_7074);
nand U9344 (N_9344,N_5565,N_5485);
nor U9345 (N_9345,N_7143,N_6231);
xnor U9346 (N_9346,N_6423,N_7335);
and U9347 (N_9347,N_5194,N_6364);
or U9348 (N_9348,N_6192,N_7248);
nand U9349 (N_9349,N_6203,N_6314);
nand U9350 (N_9350,N_5705,N_6243);
xnor U9351 (N_9351,N_6262,N_6409);
or U9352 (N_9352,N_6567,N_5909);
nand U9353 (N_9353,N_7366,N_7418);
nor U9354 (N_9354,N_6511,N_5674);
xnor U9355 (N_9355,N_5020,N_5598);
or U9356 (N_9356,N_7169,N_6816);
and U9357 (N_9357,N_5322,N_7088);
nand U9358 (N_9358,N_6615,N_6691);
xnor U9359 (N_9359,N_7128,N_7039);
xor U9360 (N_9360,N_5778,N_5426);
xor U9361 (N_9361,N_7006,N_6072);
nor U9362 (N_9362,N_6663,N_7332);
or U9363 (N_9363,N_5029,N_5134);
xnor U9364 (N_9364,N_6283,N_7248);
nand U9365 (N_9365,N_5965,N_6679);
nor U9366 (N_9366,N_7008,N_5483);
nand U9367 (N_9367,N_6431,N_6524);
xor U9368 (N_9368,N_6975,N_5839);
nor U9369 (N_9369,N_6612,N_6498);
and U9370 (N_9370,N_5766,N_5641);
xor U9371 (N_9371,N_5344,N_6495);
nor U9372 (N_9372,N_5022,N_6300);
xor U9373 (N_9373,N_5160,N_6687);
nand U9374 (N_9374,N_5747,N_7072);
and U9375 (N_9375,N_6583,N_6616);
and U9376 (N_9376,N_5452,N_6202);
nor U9377 (N_9377,N_7158,N_5349);
xnor U9378 (N_9378,N_5348,N_5707);
xor U9379 (N_9379,N_6478,N_5059);
nor U9380 (N_9380,N_6114,N_7198);
and U9381 (N_9381,N_5433,N_6630);
xor U9382 (N_9382,N_6943,N_6615);
nand U9383 (N_9383,N_5421,N_7045);
nand U9384 (N_9384,N_5599,N_5170);
or U9385 (N_9385,N_5164,N_5314);
xnor U9386 (N_9386,N_6963,N_7491);
xor U9387 (N_9387,N_7118,N_5754);
xnor U9388 (N_9388,N_6686,N_5333);
xor U9389 (N_9389,N_7087,N_5049);
xnor U9390 (N_9390,N_6436,N_5370);
nor U9391 (N_9391,N_6674,N_5527);
and U9392 (N_9392,N_6272,N_6893);
and U9393 (N_9393,N_6779,N_6397);
xor U9394 (N_9394,N_6869,N_6000);
nand U9395 (N_9395,N_7101,N_6178);
xnor U9396 (N_9396,N_6791,N_7486);
nand U9397 (N_9397,N_5503,N_5880);
xnor U9398 (N_9398,N_5122,N_6976);
or U9399 (N_9399,N_5498,N_6537);
xnor U9400 (N_9400,N_5243,N_6042);
xnor U9401 (N_9401,N_6686,N_6495);
or U9402 (N_9402,N_7010,N_6992);
or U9403 (N_9403,N_7330,N_7084);
or U9404 (N_9404,N_5249,N_6275);
or U9405 (N_9405,N_7187,N_6560);
xor U9406 (N_9406,N_5355,N_7291);
nand U9407 (N_9407,N_7337,N_5813);
xnor U9408 (N_9408,N_5790,N_6903);
xnor U9409 (N_9409,N_6637,N_6151);
and U9410 (N_9410,N_5978,N_7367);
xnor U9411 (N_9411,N_6043,N_7261);
nor U9412 (N_9412,N_6350,N_6814);
nor U9413 (N_9413,N_7383,N_7088);
nor U9414 (N_9414,N_7010,N_5114);
xor U9415 (N_9415,N_5042,N_5426);
nand U9416 (N_9416,N_5409,N_5967);
nand U9417 (N_9417,N_6530,N_5935);
nand U9418 (N_9418,N_6039,N_7142);
and U9419 (N_9419,N_7011,N_6432);
or U9420 (N_9420,N_7091,N_5076);
and U9421 (N_9421,N_7000,N_5762);
or U9422 (N_9422,N_6801,N_5464);
nand U9423 (N_9423,N_5121,N_7400);
nor U9424 (N_9424,N_5400,N_7321);
xnor U9425 (N_9425,N_7089,N_5709);
or U9426 (N_9426,N_5832,N_6132);
nor U9427 (N_9427,N_7380,N_5517);
xor U9428 (N_9428,N_6831,N_5737);
nand U9429 (N_9429,N_7157,N_6229);
or U9430 (N_9430,N_7347,N_5017);
or U9431 (N_9431,N_6617,N_5132);
xor U9432 (N_9432,N_6137,N_7110);
and U9433 (N_9433,N_5363,N_6536);
xnor U9434 (N_9434,N_6487,N_5667);
nor U9435 (N_9435,N_6029,N_5689);
and U9436 (N_9436,N_5274,N_5400);
nand U9437 (N_9437,N_5861,N_5221);
xor U9438 (N_9438,N_6783,N_6198);
nand U9439 (N_9439,N_5754,N_6858);
nand U9440 (N_9440,N_6605,N_5814);
or U9441 (N_9441,N_7429,N_5316);
nor U9442 (N_9442,N_5111,N_5884);
xnor U9443 (N_9443,N_5184,N_6274);
nor U9444 (N_9444,N_6835,N_6115);
or U9445 (N_9445,N_5164,N_5137);
xnor U9446 (N_9446,N_7201,N_7479);
nand U9447 (N_9447,N_5004,N_6237);
or U9448 (N_9448,N_5951,N_6494);
or U9449 (N_9449,N_7043,N_6830);
xor U9450 (N_9450,N_6752,N_7089);
or U9451 (N_9451,N_7282,N_7259);
or U9452 (N_9452,N_5565,N_5339);
nand U9453 (N_9453,N_5812,N_5201);
and U9454 (N_9454,N_6046,N_5055);
nand U9455 (N_9455,N_7093,N_5970);
nand U9456 (N_9456,N_5825,N_6234);
and U9457 (N_9457,N_5825,N_7402);
and U9458 (N_9458,N_6189,N_6016);
and U9459 (N_9459,N_6065,N_5341);
and U9460 (N_9460,N_5554,N_5566);
or U9461 (N_9461,N_7405,N_5745);
nor U9462 (N_9462,N_6472,N_6807);
nor U9463 (N_9463,N_6573,N_6992);
or U9464 (N_9464,N_7040,N_5817);
nor U9465 (N_9465,N_6180,N_6024);
or U9466 (N_9466,N_5599,N_5271);
and U9467 (N_9467,N_5965,N_6260);
or U9468 (N_9468,N_6974,N_6825);
nand U9469 (N_9469,N_7318,N_6339);
or U9470 (N_9470,N_5571,N_6408);
and U9471 (N_9471,N_6853,N_5808);
and U9472 (N_9472,N_5791,N_6221);
and U9473 (N_9473,N_6159,N_7000);
or U9474 (N_9474,N_5735,N_7324);
nand U9475 (N_9475,N_5440,N_7010);
nand U9476 (N_9476,N_5501,N_5408);
nand U9477 (N_9477,N_5302,N_5367);
and U9478 (N_9478,N_7263,N_5325);
xnor U9479 (N_9479,N_6249,N_5739);
xor U9480 (N_9480,N_5422,N_5448);
nor U9481 (N_9481,N_5749,N_7180);
or U9482 (N_9482,N_6045,N_6669);
and U9483 (N_9483,N_6869,N_5942);
or U9484 (N_9484,N_6258,N_6253);
or U9485 (N_9485,N_5878,N_6569);
xnor U9486 (N_9486,N_6201,N_6881);
or U9487 (N_9487,N_7326,N_5290);
nor U9488 (N_9488,N_6639,N_5475);
or U9489 (N_9489,N_6155,N_6004);
xor U9490 (N_9490,N_6418,N_6342);
xor U9491 (N_9491,N_7094,N_5998);
xor U9492 (N_9492,N_5866,N_7461);
and U9493 (N_9493,N_7195,N_5211);
nand U9494 (N_9494,N_6503,N_6162);
or U9495 (N_9495,N_5933,N_7324);
and U9496 (N_9496,N_6671,N_6458);
nor U9497 (N_9497,N_5316,N_6944);
nand U9498 (N_9498,N_5197,N_6492);
or U9499 (N_9499,N_5292,N_6489);
or U9500 (N_9500,N_6862,N_6839);
nand U9501 (N_9501,N_5374,N_5290);
and U9502 (N_9502,N_7109,N_7203);
and U9503 (N_9503,N_6848,N_6105);
nor U9504 (N_9504,N_7163,N_5121);
or U9505 (N_9505,N_7071,N_5526);
xnor U9506 (N_9506,N_5446,N_5515);
xor U9507 (N_9507,N_7215,N_5203);
xnor U9508 (N_9508,N_6744,N_5454);
and U9509 (N_9509,N_7444,N_5147);
nand U9510 (N_9510,N_5941,N_6985);
nor U9511 (N_9511,N_7167,N_6665);
and U9512 (N_9512,N_5221,N_6985);
nor U9513 (N_9513,N_6479,N_5235);
nor U9514 (N_9514,N_5491,N_5820);
and U9515 (N_9515,N_5003,N_7252);
xor U9516 (N_9516,N_5694,N_6908);
and U9517 (N_9517,N_5890,N_5220);
or U9518 (N_9518,N_5101,N_5200);
or U9519 (N_9519,N_6182,N_6417);
xor U9520 (N_9520,N_6786,N_6130);
xnor U9521 (N_9521,N_6403,N_6999);
or U9522 (N_9522,N_5790,N_6833);
nor U9523 (N_9523,N_6935,N_6611);
or U9524 (N_9524,N_5621,N_5432);
and U9525 (N_9525,N_6178,N_5477);
and U9526 (N_9526,N_6010,N_6418);
nor U9527 (N_9527,N_5647,N_6801);
or U9528 (N_9528,N_5261,N_5051);
xnor U9529 (N_9529,N_5779,N_7006);
nor U9530 (N_9530,N_7114,N_5672);
xnor U9531 (N_9531,N_6781,N_6871);
and U9532 (N_9532,N_7055,N_5485);
nand U9533 (N_9533,N_7156,N_6580);
or U9534 (N_9534,N_6194,N_6363);
nand U9535 (N_9535,N_7291,N_5615);
or U9536 (N_9536,N_5968,N_5741);
and U9537 (N_9537,N_5443,N_6360);
or U9538 (N_9538,N_6857,N_5282);
nor U9539 (N_9539,N_5219,N_5307);
or U9540 (N_9540,N_7259,N_6254);
and U9541 (N_9541,N_5041,N_5313);
or U9542 (N_9542,N_5697,N_5243);
or U9543 (N_9543,N_5211,N_7148);
or U9544 (N_9544,N_6076,N_5917);
and U9545 (N_9545,N_5236,N_6114);
and U9546 (N_9546,N_5731,N_5994);
or U9547 (N_9547,N_5942,N_5254);
xnor U9548 (N_9548,N_6792,N_7339);
xnor U9549 (N_9549,N_6817,N_7489);
or U9550 (N_9550,N_6869,N_5517);
or U9551 (N_9551,N_5575,N_6686);
xor U9552 (N_9552,N_6220,N_5383);
xnor U9553 (N_9553,N_6352,N_6910);
and U9554 (N_9554,N_6157,N_5123);
nand U9555 (N_9555,N_7066,N_5089);
nor U9556 (N_9556,N_6637,N_5879);
nand U9557 (N_9557,N_6129,N_7377);
nor U9558 (N_9558,N_5843,N_5069);
nor U9559 (N_9559,N_7356,N_7363);
or U9560 (N_9560,N_7434,N_5785);
nand U9561 (N_9561,N_7378,N_5414);
and U9562 (N_9562,N_6668,N_5087);
nand U9563 (N_9563,N_6432,N_6502);
and U9564 (N_9564,N_5504,N_6592);
nor U9565 (N_9565,N_5765,N_7080);
nand U9566 (N_9566,N_6562,N_6779);
nand U9567 (N_9567,N_6456,N_6591);
and U9568 (N_9568,N_7344,N_6310);
or U9569 (N_9569,N_5750,N_5553);
nand U9570 (N_9570,N_5432,N_6809);
or U9571 (N_9571,N_6355,N_5237);
nor U9572 (N_9572,N_5148,N_7287);
and U9573 (N_9573,N_6312,N_6405);
xor U9574 (N_9574,N_5675,N_7298);
nand U9575 (N_9575,N_5616,N_6602);
nand U9576 (N_9576,N_5860,N_7340);
xor U9577 (N_9577,N_6501,N_7330);
or U9578 (N_9578,N_5570,N_6082);
xor U9579 (N_9579,N_6490,N_7025);
or U9580 (N_9580,N_7231,N_5515);
and U9581 (N_9581,N_5973,N_5970);
or U9582 (N_9582,N_7300,N_5129);
nor U9583 (N_9583,N_6693,N_5779);
and U9584 (N_9584,N_5240,N_7461);
or U9585 (N_9585,N_6455,N_6909);
nor U9586 (N_9586,N_5776,N_6468);
and U9587 (N_9587,N_5530,N_6160);
or U9588 (N_9588,N_5812,N_7183);
nand U9589 (N_9589,N_5121,N_6850);
nor U9590 (N_9590,N_5633,N_7327);
nand U9591 (N_9591,N_6002,N_6568);
nor U9592 (N_9592,N_6072,N_6057);
xnor U9593 (N_9593,N_6484,N_6871);
or U9594 (N_9594,N_6524,N_5704);
xor U9595 (N_9595,N_5065,N_6006);
and U9596 (N_9596,N_6140,N_5391);
nor U9597 (N_9597,N_5140,N_5595);
or U9598 (N_9598,N_7312,N_6954);
or U9599 (N_9599,N_7365,N_5225);
nand U9600 (N_9600,N_5172,N_5454);
nand U9601 (N_9601,N_7345,N_7324);
nor U9602 (N_9602,N_6088,N_5063);
nor U9603 (N_9603,N_5673,N_5410);
xnor U9604 (N_9604,N_5344,N_5546);
xor U9605 (N_9605,N_6716,N_5937);
and U9606 (N_9606,N_5600,N_7434);
or U9607 (N_9607,N_6443,N_7040);
xnor U9608 (N_9608,N_5074,N_5768);
xnor U9609 (N_9609,N_6685,N_5827);
nand U9610 (N_9610,N_7307,N_5282);
nor U9611 (N_9611,N_6624,N_6284);
xnor U9612 (N_9612,N_7328,N_7469);
and U9613 (N_9613,N_6593,N_5140);
and U9614 (N_9614,N_6693,N_6267);
or U9615 (N_9615,N_6325,N_5422);
xnor U9616 (N_9616,N_5270,N_5587);
xor U9617 (N_9617,N_5023,N_5769);
and U9618 (N_9618,N_5875,N_6188);
nor U9619 (N_9619,N_7186,N_6321);
or U9620 (N_9620,N_6651,N_6760);
and U9621 (N_9621,N_5687,N_6076);
nor U9622 (N_9622,N_5618,N_7147);
xnor U9623 (N_9623,N_7448,N_5677);
nand U9624 (N_9624,N_6664,N_6204);
and U9625 (N_9625,N_5836,N_6359);
nand U9626 (N_9626,N_6831,N_6483);
xor U9627 (N_9627,N_6748,N_7412);
nand U9628 (N_9628,N_6156,N_7131);
and U9629 (N_9629,N_6886,N_5236);
and U9630 (N_9630,N_7486,N_6990);
and U9631 (N_9631,N_5920,N_6880);
nand U9632 (N_9632,N_6631,N_6535);
or U9633 (N_9633,N_5236,N_7085);
or U9634 (N_9634,N_7458,N_7375);
nor U9635 (N_9635,N_5300,N_6606);
and U9636 (N_9636,N_6445,N_6648);
nand U9637 (N_9637,N_6426,N_7185);
nand U9638 (N_9638,N_6378,N_7108);
nor U9639 (N_9639,N_6866,N_5858);
nand U9640 (N_9640,N_5971,N_5358);
and U9641 (N_9641,N_6640,N_6865);
nor U9642 (N_9642,N_7317,N_7478);
nand U9643 (N_9643,N_5175,N_6805);
and U9644 (N_9644,N_5896,N_5916);
and U9645 (N_9645,N_7418,N_6427);
nor U9646 (N_9646,N_5465,N_6917);
and U9647 (N_9647,N_6436,N_6017);
or U9648 (N_9648,N_7172,N_6936);
or U9649 (N_9649,N_5810,N_5619);
and U9650 (N_9650,N_6241,N_6424);
and U9651 (N_9651,N_6729,N_6672);
nand U9652 (N_9652,N_6469,N_7288);
or U9653 (N_9653,N_7159,N_7316);
nand U9654 (N_9654,N_5339,N_7322);
xnor U9655 (N_9655,N_7466,N_5104);
nor U9656 (N_9656,N_5278,N_5600);
and U9657 (N_9657,N_6411,N_5479);
and U9658 (N_9658,N_5775,N_5995);
or U9659 (N_9659,N_6073,N_7322);
nand U9660 (N_9660,N_6152,N_5397);
and U9661 (N_9661,N_5522,N_7032);
nor U9662 (N_9662,N_6022,N_7183);
or U9663 (N_9663,N_6628,N_5799);
or U9664 (N_9664,N_6473,N_7114);
and U9665 (N_9665,N_5620,N_6027);
or U9666 (N_9666,N_5249,N_5867);
nor U9667 (N_9667,N_6214,N_6931);
nor U9668 (N_9668,N_7425,N_6149);
or U9669 (N_9669,N_7082,N_6097);
or U9670 (N_9670,N_5391,N_6822);
nand U9671 (N_9671,N_5664,N_7271);
nand U9672 (N_9672,N_6876,N_6519);
or U9673 (N_9673,N_7019,N_6781);
xor U9674 (N_9674,N_5370,N_5027);
nor U9675 (N_9675,N_5533,N_6494);
or U9676 (N_9676,N_5987,N_5762);
nor U9677 (N_9677,N_6683,N_5892);
xor U9678 (N_9678,N_7129,N_7394);
nor U9679 (N_9679,N_5956,N_6082);
or U9680 (N_9680,N_7058,N_6646);
nand U9681 (N_9681,N_6743,N_7175);
xor U9682 (N_9682,N_7116,N_7286);
and U9683 (N_9683,N_5675,N_5687);
or U9684 (N_9684,N_5611,N_6787);
or U9685 (N_9685,N_7306,N_5545);
xnor U9686 (N_9686,N_6714,N_6391);
nand U9687 (N_9687,N_5076,N_6214);
nand U9688 (N_9688,N_6262,N_5723);
xor U9689 (N_9689,N_7480,N_5351);
nand U9690 (N_9690,N_6466,N_6654);
nor U9691 (N_9691,N_6088,N_7085);
nor U9692 (N_9692,N_6603,N_7159);
or U9693 (N_9693,N_6784,N_5572);
xnor U9694 (N_9694,N_5320,N_5690);
or U9695 (N_9695,N_6052,N_7394);
and U9696 (N_9696,N_7131,N_5804);
xnor U9697 (N_9697,N_5359,N_6959);
nor U9698 (N_9698,N_5566,N_6152);
and U9699 (N_9699,N_5598,N_5411);
or U9700 (N_9700,N_6906,N_5817);
nand U9701 (N_9701,N_6028,N_6482);
nand U9702 (N_9702,N_6955,N_5025);
or U9703 (N_9703,N_6481,N_5235);
nand U9704 (N_9704,N_6601,N_6024);
or U9705 (N_9705,N_6240,N_5375);
xor U9706 (N_9706,N_6890,N_7176);
xnor U9707 (N_9707,N_6528,N_6192);
xor U9708 (N_9708,N_6729,N_6818);
nor U9709 (N_9709,N_6355,N_6122);
nand U9710 (N_9710,N_6043,N_6847);
and U9711 (N_9711,N_6886,N_5493);
nor U9712 (N_9712,N_5330,N_5833);
and U9713 (N_9713,N_5308,N_7250);
and U9714 (N_9714,N_5955,N_6489);
nor U9715 (N_9715,N_7226,N_7145);
nor U9716 (N_9716,N_6235,N_6597);
or U9717 (N_9717,N_6711,N_7225);
nor U9718 (N_9718,N_7367,N_6311);
and U9719 (N_9719,N_6746,N_5625);
nor U9720 (N_9720,N_6190,N_5413);
nor U9721 (N_9721,N_5741,N_5885);
nand U9722 (N_9722,N_6116,N_5295);
xnor U9723 (N_9723,N_7250,N_6907);
nor U9724 (N_9724,N_6987,N_6686);
or U9725 (N_9725,N_5391,N_5183);
and U9726 (N_9726,N_6693,N_6427);
and U9727 (N_9727,N_5907,N_5380);
and U9728 (N_9728,N_6481,N_5090);
and U9729 (N_9729,N_5865,N_6619);
xnor U9730 (N_9730,N_5652,N_5162);
nor U9731 (N_9731,N_6805,N_5154);
nand U9732 (N_9732,N_5383,N_5357);
nor U9733 (N_9733,N_5179,N_6426);
xnor U9734 (N_9734,N_7378,N_6100);
nand U9735 (N_9735,N_7251,N_5748);
or U9736 (N_9736,N_6888,N_7264);
or U9737 (N_9737,N_5202,N_6366);
nand U9738 (N_9738,N_6863,N_5073);
nor U9739 (N_9739,N_6037,N_6606);
and U9740 (N_9740,N_6908,N_5082);
xor U9741 (N_9741,N_5778,N_5128);
xor U9742 (N_9742,N_5678,N_5018);
nand U9743 (N_9743,N_5924,N_5910);
xor U9744 (N_9744,N_7443,N_5136);
nor U9745 (N_9745,N_6721,N_5599);
nor U9746 (N_9746,N_6682,N_7296);
nor U9747 (N_9747,N_7160,N_5682);
nor U9748 (N_9748,N_5411,N_7480);
and U9749 (N_9749,N_6968,N_6467);
nor U9750 (N_9750,N_6546,N_6563);
and U9751 (N_9751,N_7032,N_5470);
xor U9752 (N_9752,N_6526,N_6490);
nand U9753 (N_9753,N_6439,N_6030);
nand U9754 (N_9754,N_6504,N_6883);
xor U9755 (N_9755,N_7039,N_6232);
nand U9756 (N_9756,N_6844,N_7263);
and U9757 (N_9757,N_7143,N_6125);
xnor U9758 (N_9758,N_6698,N_7046);
xor U9759 (N_9759,N_5837,N_5504);
nand U9760 (N_9760,N_6196,N_6676);
nor U9761 (N_9761,N_7312,N_7158);
xnor U9762 (N_9762,N_5140,N_6990);
xor U9763 (N_9763,N_6717,N_6196);
nor U9764 (N_9764,N_7192,N_6498);
or U9765 (N_9765,N_6839,N_7460);
and U9766 (N_9766,N_6680,N_5260);
xnor U9767 (N_9767,N_6773,N_7013);
or U9768 (N_9768,N_6777,N_7048);
nor U9769 (N_9769,N_6982,N_7301);
xnor U9770 (N_9770,N_5873,N_5584);
nand U9771 (N_9771,N_5343,N_6125);
xor U9772 (N_9772,N_7292,N_5015);
and U9773 (N_9773,N_5765,N_5623);
xnor U9774 (N_9774,N_5755,N_5459);
nor U9775 (N_9775,N_5450,N_5338);
nor U9776 (N_9776,N_7333,N_5958);
or U9777 (N_9777,N_5694,N_7403);
nand U9778 (N_9778,N_6996,N_5677);
nand U9779 (N_9779,N_6461,N_5001);
or U9780 (N_9780,N_7460,N_6853);
xor U9781 (N_9781,N_6630,N_6628);
and U9782 (N_9782,N_6428,N_6515);
and U9783 (N_9783,N_5503,N_5353);
and U9784 (N_9784,N_7244,N_5447);
nand U9785 (N_9785,N_5097,N_5585);
xor U9786 (N_9786,N_6978,N_6698);
nand U9787 (N_9787,N_7178,N_6954);
and U9788 (N_9788,N_5758,N_7131);
xnor U9789 (N_9789,N_6452,N_6168);
nand U9790 (N_9790,N_5059,N_7081);
nand U9791 (N_9791,N_7289,N_7119);
and U9792 (N_9792,N_5676,N_5099);
or U9793 (N_9793,N_5075,N_6476);
and U9794 (N_9794,N_6937,N_7019);
xor U9795 (N_9795,N_5532,N_5428);
nor U9796 (N_9796,N_7416,N_6384);
or U9797 (N_9797,N_5699,N_7122);
or U9798 (N_9798,N_5081,N_5744);
and U9799 (N_9799,N_5737,N_7149);
xnor U9800 (N_9800,N_6808,N_6681);
xnor U9801 (N_9801,N_5010,N_6541);
xnor U9802 (N_9802,N_5236,N_5976);
xnor U9803 (N_9803,N_7007,N_5084);
and U9804 (N_9804,N_6054,N_6408);
and U9805 (N_9805,N_6940,N_5678);
nand U9806 (N_9806,N_6099,N_6745);
and U9807 (N_9807,N_5578,N_5767);
or U9808 (N_9808,N_6818,N_6737);
xor U9809 (N_9809,N_7226,N_6292);
xor U9810 (N_9810,N_6958,N_6941);
nor U9811 (N_9811,N_6055,N_5624);
or U9812 (N_9812,N_7219,N_7209);
and U9813 (N_9813,N_6266,N_5504);
xnor U9814 (N_9814,N_6739,N_7151);
and U9815 (N_9815,N_5493,N_7159);
xor U9816 (N_9816,N_6135,N_5525);
or U9817 (N_9817,N_5925,N_6518);
or U9818 (N_9818,N_7435,N_5333);
nor U9819 (N_9819,N_6611,N_5455);
or U9820 (N_9820,N_7011,N_7197);
or U9821 (N_9821,N_7217,N_6787);
and U9822 (N_9822,N_7081,N_5267);
or U9823 (N_9823,N_6929,N_6483);
xnor U9824 (N_9824,N_6524,N_5193);
nor U9825 (N_9825,N_6257,N_6060);
nor U9826 (N_9826,N_6440,N_7284);
and U9827 (N_9827,N_6979,N_6070);
xor U9828 (N_9828,N_5805,N_7378);
or U9829 (N_9829,N_6369,N_5748);
nor U9830 (N_9830,N_6340,N_5210);
or U9831 (N_9831,N_5046,N_6691);
and U9832 (N_9832,N_5500,N_6075);
and U9833 (N_9833,N_6791,N_5212);
and U9834 (N_9834,N_5281,N_7374);
and U9835 (N_9835,N_6316,N_5398);
and U9836 (N_9836,N_5029,N_6389);
nand U9837 (N_9837,N_6855,N_5383);
nand U9838 (N_9838,N_5164,N_6236);
nand U9839 (N_9839,N_5846,N_6675);
xor U9840 (N_9840,N_5556,N_6185);
xor U9841 (N_9841,N_6364,N_5379);
and U9842 (N_9842,N_5740,N_6203);
nor U9843 (N_9843,N_5631,N_5256);
and U9844 (N_9844,N_6470,N_5322);
or U9845 (N_9845,N_6574,N_7185);
nand U9846 (N_9846,N_6083,N_6128);
xnor U9847 (N_9847,N_6109,N_5283);
nand U9848 (N_9848,N_6086,N_6131);
nand U9849 (N_9849,N_7480,N_6353);
and U9850 (N_9850,N_6652,N_5540);
and U9851 (N_9851,N_5795,N_5271);
xnor U9852 (N_9852,N_5277,N_6711);
nor U9853 (N_9853,N_7205,N_5004);
xnor U9854 (N_9854,N_5593,N_7303);
nor U9855 (N_9855,N_6665,N_7451);
nand U9856 (N_9856,N_7213,N_6589);
xnor U9857 (N_9857,N_7032,N_6401);
or U9858 (N_9858,N_6474,N_6107);
nand U9859 (N_9859,N_6731,N_6309);
and U9860 (N_9860,N_5586,N_6342);
or U9861 (N_9861,N_6875,N_5226);
or U9862 (N_9862,N_7143,N_5763);
nand U9863 (N_9863,N_6754,N_6641);
nor U9864 (N_9864,N_6039,N_5732);
xor U9865 (N_9865,N_6020,N_7024);
or U9866 (N_9866,N_5580,N_6238);
and U9867 (N_9867,N_6048,N_5003);
and U9868 (N_9868,N_5221,N_6559);
nor U9869 (N_9869,N_5944,N_5537);
nand U9870 (N_9870,N_7384,N_6538);
nor U9871 (N_9871,N_5740,N_6122);
xnor U9872 (N_9872,N_6362,N_6491);
xnor U9873 (N_9873,N_6176,N_6719);
nor U9874 (N_9874,N_6779,N_7355);
or U9875 (N_9875,N_5574,N_7007);
and U9876 (N_9876,N_6232,N_6130);
nor U9877 (N_9877,N_7259,N_6022);
xnor U9878 (N_9878,N_7201,N_6575);
nor U9879 (N_9879,N_5967,N_6120);
nand U9880 (N_9880,N_5079,N_6120);
xor U9881 (N_9881,N_5977,N_6769);
or U9882 (N_9882,N_6203,N_5714);
xnor U9883 (N_9883,N_5965,N_6533);
xnor U9884 (N_9884,N_5703,N_5426);
xnor U9885 (N_9885,N_7096,N_7388);
xnor U9886 (N_9886,N_5506,N_5949);
xnor U9887 (N_9887,N_6256,N_7253);
and U9888 (N_9888,N_5997,N_5288);
nor U9889 (N_9889,N_7365,N_5698);
xor U9890 (N_9890,N_6761,N_5096);
xor U9891 (N_9891,N_6341,N_6843);
nor U9892 (N_9892,N_7183,N_5910);
or U9893 (N_9893,N_5382,N_5221);
or U9894 (N_9894,N_7089,N_7457);
or U9895 (N_9895,N_6603,N_6367);
nor U9896 (N_9896,N_7388,N_7282);
nand U9897 (N_9897,N_6796,N_5798);
nor U9898 (N_9898,N_7414,N_6365);
xor U9899 (N_9899,N_5883,N_6089);
nor U9900 (N_9900,N_5804,N_7442);
nor U9901 (N_9901,N_5031,N_7486);
or U9902 (N_9902,N_6979,N_5238);
nor U9903 (N_9903,N_6358,N_5050);
nand U9904 (N_9904,N_6290,N_5846);
and U9905 (N_9905,N_6982,N_5286);
nor U9906 (N_9906,N_5301,N_6615);
xor U9907 (N_9907,N_6129,N_6819);
nand U9908 (N_9908,N_7140,N_5664);
xnor U9909 (N_9909,N_5047,N_5232);
nor U9910 (N_9910,N_7081,N_7365);
nand U9911 (N_9911,N_6592,N_5509);
xnor U9912 (N_9912,N_6266,N_5969);
nand U9913 (N_9913,N_6086,N_6512);
nand U9914 (N_9914,N_6465,N_7217);
nand U9915 (N_9915,N_5141,N_5055);
nand U9916 (N_9916,N_5776,N_5435);
nor U9917 (N_9917,N_6992,N_5670);
and U9918 (N_9918,N_6595,N_6175);
xor U9919 (N_9919,N_7206,N_7153);
xnor U9920 (N_9920,N_5075,N_5292);
or U9921 (N_9921,N_6830,N_7024);
nor U9922 (N_9922,N_6393,N_5655);
nor U9923 (N_9923,N_5283,N_6369);
or U9924 (N_9924,N_6844,N_5337);
and U9925 (N_9925,N_7072,N_5937);
nor U9926 (N_9926,N_5075,N_5745);
nand U9927 (N_9927,N_5691,N_5739);
and U9928 (N_9928,N_7383,N_6248);
or U9929 (N_9929,N_6821,N_6030);
nand U9930 (N_9930,N_5867,N_7360);
and U9931 (N_9931,N_7116,N_5836);
and U9932 (N_9932,N_5326,N_5099);
or U9933 (N_9933,N_7366,N_6161);
or U9934 (N_9934,N_5136,N_7336);
xnor U9935 (N_9935,N_6072,N_6885);
nor U9936 (N_9936,N_7096,N_7205);
nand U9937 (N_9937,N_6834,N_6643);
and U9938 (N_9938,N_6820,N_6119);
xor U9939 (N_9939,N_6827,N_5249);
nor U9940 (N_9940,N_6808,N_6789);
nor U9941 (N_9941,N_6246,N_5501);
nor U9942 (N_9942,N_7322,N_6368);
nand U9943 (N_9943,N_5823,N_5247);
nor U9944 (N_9944,N_5219,N_5510);
xor U9945 (N_9945,N_6895,N_6706);
and U9946 (N_9946,N_6426,N_5244);
xnor U9947 (N_9947,N_7127,N_5478);
or U9948 (N_9948,N_5176,N_6181);
xnor U9949 (N_9949,N_6912,N_6517);
nor U9950 (N_9950,N_6637,N_6524);
nor U9951 (N_9951,N_5129,N_6668);
nor U9952 (N_9952,N_6620,N_5762);
nor U9953 (N_9953,N_7448,N_5382);
or U9954 (N_9954,N_7069,N_5791);
nor U9955 (N_9955,N_6405,N_6250);
or U9956 (N_9956,N_5142,N_5221);
nand U9957 (N_9957,N_6222,N_7198);
and U9958 (N_9958,N_6515,N_6535);
nand U9959 (N_9959,N_5431,N_5161);
or U9960 (N_9960,N_5480,N_6056);
and U9961 (N_9961,N_6291,N_7245);
and U9962 (N_9962,N_6833,N_6444);
xnor U9963 (N_9963,N_7440,N_6129);
nand U9964 (N_9964,N_6666,N_6638);
xor U9965 (N_9965,N_5536,N_5604);
or U9966 (N_9966,N_7453,N_6419);
or U9967 (N_9967,N_6370,N_6533);
nand U9968 (N_9968,N_5546,N_6415);
or U9969 (N_9969,N_6799,N_6582);
xnor U9970 (N_9970,N_6300,N_5228);
or U9971 (N_9971,N_5129,N_5836);
and U9972 (N_9972,N_6719,N_7258);
and U9973 (N_9973,N_6116,N_6480);
or U9974 (N_9974,N_6463,N_6788);
or U9975 (N_9975,N_6723,N_6281);
xnor U9976 (N_9976,N_5009,N_5822);
nand U9977 (N_9977,N_6840,N_5117);
xor U9978 (N_9978,N_5795,N_6921);
and U9979 (N_9979,N_7004,N_7329);
or U9980 (N_9980,N_7071,N_5568);
nand U9981 (N_9981,N_6631,N_5786);
or U9982 (N_9982,N_7119,N_5994);
or U9983 (N_9983,N_7383,N_6436);
nand U9984 (N_9984,N_6270,N_5756);
xor U9985 (N_9985,N_5507,N_5922);
xor U9986 (N_9986,N_7262,N_5483);
nand U9987 (N_9987,N_6737,N_5440);
or U9988 (N_9988,N_5845,N_6055);
nor U9989 (N_9989,N_6352,N_5022);
or U9990 (N_9990,N_5420,N_6689);
and U9991 (N_9991,N_5375,N_5408);
and U9992 (N_9992,N_5077,N_7099);
or U9993 (N_9993,N_6682,N_5991);
nor U9994 (N_9994,N_5941,N_7008);
xnor U9995 (N_9995,N_7386,N_6642);
and U9996 (N_9996,N_6116,N_6823);
and U9997 (N_9997,N_6457,N_7295);
xnor U9998 (N_9998,N_7113,N_6612);
xor U9999 (N_9999,N_6563,N_6965);
nand UO_0 (O_0,N_8346,N_9328);
nor UO_1 (O_1,N_8364,N_9400);
and UO_2 (O_2,N_8746,N_7974);
nand UO_3 (O_3,N_8230,N_8443);
xor UO_4 (O_4,N_9936,N_9098);
nor UO_5 (O_5,N_7900,N_7919);
nand UO_6 (O_6,N_7680,N_8641);
and UO_7 (O_7,N_7952,N_8626);
and UO_8 (O_8,N_8127,N_9242);
nand UO_9 (O_9,N_8924,N_8069);
nand UO_10 (O_10,N_8500,N_9989);
or UO_11 (O_11,N_8254,N_9303);
nand UO_12 (O_12,N_8320,N_7679);
xnor UO_13 (O_13,N_7791,N_7997);
and UO_14 (O_14,N_9830,N_9299);
nand UO_15 (O_15,N_9636,N_8587);
nand UO_16 (O_16,N_8053,N_8605);
and UO_17 (O_17,N_9810,N_8431);
nand UO_18 (O_18,N_8942,N_7740);
nor UO_19 (O_19,N_8134,N_9865);
xor UO_20 (O_20,N_8283,N_7670);
xor UO_21 (O_21,N_9403,N_8154);
or UO_22 (O_22,N_7707,N_9512);
nor UO_23 (O_23,N_7854,N_7800);
nand UO_24 (O_24,N_7693,N_9150);
and UO_25 (O_25,N_7768,N_8063);
nor UO_26 (O_26,N_9545,N_9493);
nand UO_27 (O_27,N_7823,N_9111);
and UO_28 (O_28,N_7896,N_7603);
nand UO_29 (O_29,N_8397,N_9854);
xnor UO_30 (O_30,N_8041,N_9958);
and UO_31 (O_31,N_7810,N_8208);
and UO_32 (O_32,N_9286,N_9060);
or UO_33 (O_33,N_9185,N_9742);
or UO_34 (O_34,N_9506,N_8671);
or UO_35 (O_35,N_8452,N_7987);
and UO_36 (O_36,N_8610,N_8516);
or UO_37 (O_37,N_9215,N_9892);
nor UO_38 (O_38,N_8023,N_7792);
or UO_39 (O_39,N_8355,N_8559);
xor UO_40 (O_40,N_8373,N_8467);
or UO_41 (O_41,N_9095,N_9174);
and UO_42 (O_42,N_8710,N_9556);
nand UO_43 (O_43,N_8271,N_8335);
and UO_44 (O_44,N_9255,N_8534);
and UO_45 (O_45,N_7542,N_8143);
and UO_46 (O_46,N_9869,N_8140);
or UO_47 (O_47,N_8912,N_8814);
nor UO_48 (O_48,N_8943,N_9494);
and UO_49 (O_49,N_8082,N_8178);
and UO_50 (O_50,N_8648,N_8057);
or UO_51 (O_51,N_8078,N_9935);
xor UO_52 (O_52,N_9934,N_9139);
and UO_53 (O_53,N_8709,N_7733);
or UO_54 (O_54,N_8354,N_9689);
nor UO_55 (O_55,N_9718,N_8766);
and UO_56 (O_56,N_7774,N_8223);
and UO_57 (O_57,N_9559,N_9681);
or UO_58 (O_58,N_7538,N_7637);
nand UO_59 (O_59,N_9132,N_8358);
xnor UO_60 (O_60,N_9775,N_8582);
xor UO_61 (O_61,N_9282,N_8994);
nand UO_62 (O_62,N_8940,N_8332);
and UO_63 (O_63,N_9265,N_8586);
xnor UO_64 (O_64,N_7942,N_8611);
nand UO_65 (O_65,N_9089,N_9814);
and UO_66 (O_66,N_8929,N_9894);
or UO_67 (O_67,N_9912,N_8636);
xnor UO_68 (O_68,N_9991,N_9143);
nor UO_69 (O_69,N_8536,N_7561);
xnor UO_70 (O_70,N_8256,N_9340);
nor UO_71 (O_71,N_8333,N_7552);
and UO_72 (O_72,N_9858,N_8345);
nand UO_73 (O_73,N_9823,N_8732);
and UO_74 (O_74,N_9729,N_8010);
nand UO_75 (O_75,N_7698,N_8585);
or UO_76 (O_76,N_9219,N_8203);
xor UO_77 (O_77,N_9497,N_7647);
nand UO_78 (O_78,N_9479,N_8530);
and UO_79 (O_79,N_9076,N_9040);
xnor UO_80 (O_80,N_9369,N_9010);
and UO_81 (O_81,N_7711,N_8878);
nor UO_82 (O_82,N_8977,N_8105);
and UO_83 (O_83,N_7861,N_8511);
xnor UO_84 (O_84,N_9716,N_7777);
nor UO_85 (O_85,N_9474,N_9020);
nand UO_86 (O_86,N_9260,N_8347);
or UO_87 (O_87,N_9376,N_8250);
and UO_88 (O_88,N_8925,N_8522);
nand UO_89 (O_89,N_8549,N_8278);
xnor UO_90 (O_90,N_9356,N_7890);
or UO_91 (O_91,N_8150,N_7583);
nand UO_92 (O_92,N_7545,N_8176);
or UO_93 (O_93,N_7833,N_9832);
or UO_94 (O_94,N_9570,N_8820);
and UO_95 (O_95,N_8909,N_9438);
xor UO_96 (O_96,N_8160,N_9102);
nand UO_97 (O_97,N_8623,N_9240);
or UO_98 (O_98,N_7520,N_8319);
nor UO_99 (O_99,N_8003,N_8427);
and UO_100 (O_100,N_8677,N_9530);
nand UO_101 (O_101,N_7829,N_9104);
xnor UO_102 (O_102,N_7968,N_9468);
xor UO_103 (O_103,N_7834,N_9940);
nand UO_104 (O_104,N_8120,N_8778);
or UO_105 (O_105,N_9676,N_8324);
nand UO_106 (O_106,N_8029,N_8122);
or UO_107 (O_107,N_9730,N_9586);
nor UO_108 (O_108,N_8435,N_7534);
nand UO_109 (O_109,N_8341,N_8181);
xor UO_110 (O_110,N_8465,N_9033);
nor UO_111 (O_111,N_9529,N_9027);
or UO_112 (O_112,N_8987,N_7696);
xnor UO_113 (O_113,N_9843,N_7556);
and UO_114 (O_114,N_7627,N_9696);
and UO_115 (O_115,N_8436,N_8253);
xor UO_116 (O_116,N_7694,N_8863);
nor UO_117 (O_117,N_9756,N_7784);
nor UO_118 (O_118,N_7742,N_8696);
and UO_119 (O_119,N_9993,N_8566);
nor UO_120 (O_120,N_9527,N_8348);
and UO_121 (O_121,N_9152,N_9323);
or UO_122 (O_122,N_9607,N_9432);
nor UO_123 (O_123,N_8372,N_9650);
nor UO_124 (O_124,N_7775,N_9961);
and UO_125 (O_125,N_8818,N_8246);
or UO_126 (O_126,N_8414,N_9941);
nor UO_127 (O_127,N_9442,N_8706);
xor UO_128 (O_128,N_8875,N_8213);
nor UO_129 (O_129,N_9580,N_8043);
or UO_130 (O_130,N_8224,N_8855);
or UO_131 (O_131,N_8973,N_7855);
xor UO_132 (O_132,N_8758,N_7879);
nor UO_133 (O_133,N_9080,N_9051);
and UO_134 (O_134,N_8799,N_8212);
or UO_135 (O_135,N_9176,N_8039);
and UO_136 (O_136,N_8448,N_8386);
nand UO_137 (O_137,N_9598,N_7801);
xnor UO_138 (O_138,N_9500,N_9975);
or UO_139 (O_139,N_9999,N_9075);
and UO_140 (O_140,N_8817,N_7973);
or UO_141 (O_141,N_7803,N_7958);
nand UO_142 (O_142,N_9271,N_7736);
nand UO_143 (O_143,N_8411,N_8288);
or UO_144 (O_144,N_7675,N_9429);
xnor UO_145 (O_145,N_8784,N_9646);
nor UO_146 (O_146,N_7894,N_9608);
nor UO_147 (O_147,N_8051,N_8813);
xor UO_148 (O_148,N_9887,N_9879);
or UO_149 (O_149,N_9467,N_9722);
nand UO_150 (O_150,N_9754,N_9460);
nand UO_151 (O_151,N_7957,N_8665);
and UO_152 (O_152,N_8187,N_8954);
nor UO_153 (O_153,N_8395,N_8596);
or UO_154 (O_154,N_8849,N_9873);
nand UO_155 (O_155,N_9893,N_8316);
xnor UO_156 (O_156,N_7687,N_9984);
and UO_157 (O_157,N_9385,N_9433);
or UO_158 (O_158,N_8828,N_7532);
and UO_159 (O_159,N_9874,N_8872);
xnor UO_160 (O_160,N_9755,N_8770);
nand UO_161 (O_161,N_8811,N_9542);
xnor UO_162 (O_162,N_8357,N_7726);
or UO_163 (O_163,N_8231,N_7937);
nor UO_164 (O_164,N_9862,N_8115);
nand UO_165 (O_165,N_9985,N_9337);
or UO_166 (O_166,N_7773,N_7685);
or UO_167 (O_167,N_9844,N_8888);
xor UO_168 (O_168,N_8951,N_9245);
or UO_169 (O_169,N_9262,N_8824);
and UO_170 (O_170,N_9405,N_8966);
xor UO_171 (O_171,N_7660,N_9254);
nor UO_172 (O_172,N_7510,N_7554);
nor UO_173 (O_173,N_8403,N_9693);
and UO_174 (O_174,N_8591,N_8017);
nand UO_175 (O_175,N_8524,N_9485);
or UO_176 (O_176,N_9192,N_8106);
nor UO_177 (O_177,N_7850,N_8315);
nand UO_178 (O_178,N_9083,N_7537);
and UO_179 (O_179,N_7686,N_9634);
and UO_180 (O_180,N_7935,N_8180);
or UO_181 (O_181,N_9135,N_9523);
or UO_182 (O_182,N_7805,N_8701);
xnor UO_183 (O_183,N_7926,N_9914);
nand UO_184 (O_184,N_9436,N_8077);
or UO_185 (O_185,N_9908,N_7513);
and UO_186 (O_186,N_7518,N_7522);
nand UO_187 (O_187,N_9410,N_9937);
nand UO_188 (O_188,N_7710,N_8717);
nor UO_189 (O_189,N_9572,N_9759);
xor UO_190 (O_190,N_8862,N_9456);
or UO_191 (O_191,N_7663,N_7555);
or UO_192 (O_192,N_8833,N_9825);
or UO_193 (O_193,N_9939,N_8577);
or UO_194 (O_194,N_9236,N_9890);
or UO_195 (O_195,N_8287,N_7525);
nor UO_196 (O_196,N_9004,N_8290);
nand UO_197 (O_197,N_9656,N_7645);
or UO_198 (O_198,N_8282,N_8712);
xor UO_199 (O_199,N_9610,N_8590);
or UO_200 (O_200,N_7531,N_9671);
nor UO_201 (O_201,N_9443,N_9980);
and UO_202 (O_202,N_9791,N_8607);
and UO_203 (O_203,N_9588,N_8895);
xnor UO_204 (O_204,N_9166,N_7910);
nand UO_205 (O_205,N_7700,N_8441);
or UO_206 (O_206,N_8504,N_8344);
nor UO_207 (O_207,N_9628,N_8019);
or UO_208 (O_208,N_9522,N_9085);
xor UO_209 (O_209,N_9885,N_9228);
nand UO_210 (O_210,N_7843,N_8234);
nand UO_211 (O_211,N_9644,N_8228);
nand UO_212 (O_212,N_8484,N_9109);
nand UO_213 (O_213,N_7868,N_7960);
nor UO_214 (O_214,N_8184,N_7574);
or UO_215 (O_215,N_7604,N_8769);
xnor UO_216 (O_216,N_9952,N_8616);
or UO_217 (O_217,N_8734,N_8383);
xor UO_218 (O_218,N_7544,N_9402);
nor UO_219 (O_219,N_7811,N_9071);
or UO_220 (O_220,N_8462,N_9324);
nor UO_221 (O_221,N_9651,N_9048);
or UO_222 (O_222,N_9028,N_9330);
and UO_223 (O_223,N_9437,N_9649);
nand UO_224 (O_224,N_8891,N_9218);
and UO_225 (O_225,N_9054,N_9453);
xnor UO_226 (O_226,N_8464,N_8835);
xor UO_227 (O_227,N_8310,N_9744);
or UO_228 (O_228,N_8948,N_9964);
xnor UO_229 (O_229,N_9235,N_8752);
xnor UO_230 (O_230,N_8576,N_8666);
nand UO_231 (O_231,N_8406,N_9747);
and UO_232 (O_232,N_7760,N_7712);
or UO_233 (O_233,N_7503,N_9896);
nor UO_234 (O_234,N_9942,N_8356);
xor UO_235 (O_235,N_8437,N_8211);
nor UO_236 (O_236,N_9036,N_7920);
nor UO_237 (O_237,N_7962,N_9971);
nor UO_238 (O_238,N_7776,N_8667);
nor UO_239 (O_239,N_9346,N_8955);
or UO_240 (O_240,N_8601,N_9359);
nor UO_241 (O_241,N_8777,N_8661);
nand UO_242 (O_242,N_8497,N_7882);
xor UO_243 (O_243,N_8410,N_8119);
nand UO_244 (O_244,N_8844,N_7923);
and UO_245 (O_245,N_8620,N_7598);
nor UO_246 (O_246,N_8776,N_7543);
or UO_247 (O_247,N_8705,N_8961);
xnor UO_248 (O_248,N_8632,N_8939);
nor UO_249 (O_249,N_8259,N_9074);
xnor UO_250 (O_250,N_7977,N_8980);
xnor UO_251 (O_251,N_9837,N_8311);
nor UO_252 (O_252,N_8997,N_9505);
xor UO_253 (O_253,N_9031,N_8166);
xor UO_254 (O_254,N_8870,N_8771);
or UO_255 (O_255,N_8471,N_9956);
or UO_256 (O_256,N_9372,N_8300);
or UO_257 (O_257,N_8547,N_8475);
or UO_258 (O_258,N_8478,N_8727);
and UO_259 (O_259,N_9906,N_8136);
or UO_260 (O_260,N_8377,N_9576);
and UO_261 (O_261,N_7763,N_8907);
or UO_262 (O_262,N_9391,N_8753);
xor UO_263 (O_263,N_8135,N_9827);
xor UO_264 (O_264,N_9540,N_9470);
xnor UO_265 (O_265,N_9171,N_8487);
nand UO_266 (O_266,N_9574,N_8563);
nand UO_267 (O_267,N_8309,N_9960);
or UO_268 (O_268,N_8255,N_7783);
or UO_269 (O_269,N_8751,N_9435);
nor UO_270 (O_270,N_9558,N_8897);
and UO_271 (O_271,N_9127,N_8873);
nor UO_272 (O_272,N_9959,N_8655);
nor UO_273 (O_273,N_7963,N_7743);
and UO_274 (O_274,N_9969,N_9248);
nand UO_275 (O_275,N_9297,N_9230);
nand UO_276 (O_276,N_7989,N_8903);
xor UO_277 (O_277,N_8200,N_8656);
nand UO_278 (O_278,N_8550,N_9953);
and UO_279 (O_279,N_9302,N_8196);
and UO_280 (O_280,N_8056,N_8554);
or UO_281 (O_281,N_9712,N_7815);
xnor UO_282 (O_282,N_9763,N_8363);
nor UO_283 (O_283,N_8564,N_9995);
nand UO_284 (O_284,N_9792,N_8679);
xor UO_285 (O_285,N_9065,N_8353);
nor UO_286 (O_286,N_8092,N_9180);
xor UO_287 (O_287,N_8350,N_8318);
nor UO_288 (O_288,N_8738,N_8832);
and UO_289 (O_289,N_8236,N_7881);
xor UO_290 (O_290,N_8979,N_9804);
nand UO_291 (O_291,N_9162,N_8900);
and UO_292 (O_292,N_9536,N_9167);
xor UO_293 (O_293,N_8541,N_7580);
or UO_294 (O_294,N_9277,N_8768);
or UO_295 (O_295,N_8974,N_8993);
nor UO_296 (O_296,N_9888,N_9066);
xor UO_297 (O_297,N_9263,N_9341);
nand UO_298 (O_298,N_8146,N_7853);
xnor UO_299 (O_299,N_9809,N_7596);
nand UO_300 (O_300,N_9115,N_8412);
nor UO_301 (O_301,N_7579,N_7691);
and UO_302 (O_302,N_9283,N_8447);
nor UO_303 (O_303,N_8673,N_7812);
or UO_304 (O_304,N_7569,N_9211);
nand UO_305 (O_305,N_9731,N_8138);
and UO_306 (O_306,N_8201,N_9370);
nor UO_307 (O_307,N_8015,N_7669);
or UO_308 (O_308,N_9563,N_8739);
and UO_309 (O_309,N_9547,N_9491);
xnor UO_310 (O_310,N_9700,N_8243);
or UO_311 (O_311,N_8266,N_7618);
nand UO_312 (O_312,N_9769,N_8195);
nor UO_313 (O_313,N_8528,N_9399);
or UO_314 (O_314,N_8477,N_9029);
nor UO_315 (O_315,N_8006,N_8328);
nand UO_316 (O_316,N_9018,N_8568);
nand UO_317 (O_317,N_9968,N_8859);
nand UO_318 (O_318,N_7880,N_9762);
nand UO_319 (O_319,N_9582,N_9695);
nand UO_320 (O_320,N_9683,N_9383);
and UO_321 (O_321,N_9709,N_9510);
and UO_322 (O_322,N_9904,N_9087);
nor UO_323 (O_323,N_8574,N_9182);
xor UO_324 (O_324,N_9123,N_7820);
and UO_325 (O_325,N_7954,N_7657);
xor UO_326 (O_326,N_8635,N_8094);
xor UO_327 (O_327,N_7741,N_9519);
nand UO_328 (O_328,N_7844,N_7655);
nor UO_329 (O_329,N_8326,N_9239);
nor UO_330 (O_330,N_9928,N_8426);
xor UO_331 (O_331,N_7609,N_8953);
nand UO_332 (O_332,N_9156,N_7746);
or UO_333 (O_333,N_9070,N_8845);
xnor UO_334 (O_334,N_8906,N_8985);
nand UO_335 (O_335,N_9278,N_7750);
and UO_336 (O_336,N_7546,N_8887);
nor UO_337 (O_337,N_8747,N_9408);
nor UO_338 (O_338,N_8007,N_8647);
nor UO_339 (O_339,N_9032,N_8454);
or UO_340 (O_340,N_7914,N_8482);
nor UO_341 (O_341,N_8205,N_9378);
or UO_342 (O_342,N_9938,N_7563);
nand UO_343 (O_343,N_7903,N_9581);
xnor UO_344 (O_344,N_8731,N_7925);
and UO_345 (O_345,N_8698,N_9332);
nand UO_346 (O_346,N_9099,N_7908);
and UO_347 (O_347,N_9314,N_8640);
nand UO_348 (O_348,N_9309,N_7842);
nor UO_349 (O_349,N_8173,N_9499);
or UO_350 (O_350,N_8393,N_8931);
or UO_351 (O_351,N_9014,N_8399);
or UO_352 (O_352,N_8472,N_8113);
nand UO_353 (O_353,N_7749,N_8837);
xnor UO_354 (O_354,N_8233,N_9243);
xnor UO_355 (O_355,N_9623,N_8096);
xor UO_356 (O_356,N_9049,N_8904);
nor UO_357 (O_357,N_9390,N_7643);
nand UO_358 (O_358,N_9905,N_7929);
xor UO_359 (O_359,N_9599,N_9318);
and UO_360 (O_360,N_8327,N_9772);
xnor UO_361 (O_361,N_7828,N_8513);
and UO_362 (O_362,N_8546,N_9112);
nand UO_363 (O_363,N_9119,N_9268);
xor UO_364 (O_364,N_8539,N_7507);
xnor UO_365 (O_365,N_8579,N_8240);
or UO_366 (O_366,N_9382,N_8059);
xor UO_367 (O_367,N_9699,N_9566);
and UO_368 (O_368,N_8194,N_9196);
and UO_369 (O_369,N_7547,N_9678);
and UO_370 (O_370,N_9535,N_9720);
nand UO_371 (O_371,N_9125,N_7993);
and UO_372 (O_372,N_9415,N_7995);
nor UO_373 (O_373,N_7658,N_8526);
xor UO_374 (O_374,N_9949,N_8680);
xnor UO_375 (O_375,N_7994,N_8235);
xor UO_376 (O_376,N_8144,N_8790);
or UO_377 (O_377,N_9767,N_8918);
nor UO_378 (O_378,N_7761,N_9884);
nand UO_379 (O_379,N_7584,N_9172);
nor UO_380 (O_380,N_8580,N_9261);
nand UO_381 (O_381,N_7864,N_7949);
nand UO_382 (O_382,N_7869,N_8681);
nand UO_383 (O_383,N_7876,N_8996);
nor UO_384 (O_384,N_9840,N_7511);
nor UO_385 (O_385,N_9761,N_7759);
nand UO_386 (O_386,N_9600,N_9101);
nor UO_387 (O_387,N_7909,N_9721);
xnor UO_388 (O_388,N_9963,N_7593);
nand UO_389 (O_389,N_8274,N_9684);
or UO_390 (O_390,N_8428,N_9137);
or UO_391 (O_391,N_9223,N_9508);
nor UO_392 (O_392,N_8198,N_8062);
nor UO_393 (O_393,N_9351,N_9913);
xor UO_394 (O_394,N_8400,N_8329);
or UO_395 (O_395,N_9670,N_9872);
and UO_396 (O_396,N_7639,N_9451);
nand UO_397 (O_397,N_7568,N_8091);
and UO_398 (O_398,N_9238,N_9648);
nor UO_399 (O_399,N_8207,N_7838);
nand UO_400 (O_400,N_9414,N_8773);
and UO_401 (O_401,N_9787,N_9147);
or UO_402 (O_402,N_9903,N_8026);
and UO_403 (O_403,N_9190,N_9525);
and UO_404 (O_404,N_9045,N_8131);
and UO_405 (O_405,N_9226,N_8483);
nand UO_406 (O_406,N_7804,N_7671);
xnor UO_407 (O_407,N_7500,N_9622);
or UO_408 (O_408,N_8459,N_8141);
nor UO_409 (O_409,N_8562,N_9669);
xnor UO_410 (O_410,N_8080,N_8998);
and UO_411 (O_411,N_9360,N_8794);
nand UO_412 (O_412,N_8286,N_7617);
or UO_413 (O_413,N_9821,N_8296);
nor UO_414 (O_414,N_8651,N_9533);
nand UO_415 (O_415,N_9770,N_8978);
or UO_416 (O_416,N_8759,N_9674);
and UO_417 (O_417,N_7560,N_9298);
xnor UO_418 (O_418,N_9401,N_8085);
nor UO_419 (O_419,N_7817,N_7874);
or UO_420 (O_420,N_9998,N_9394);
and UO_421 (O_421,N_9024,N_8889);
or UO_422 (O_422,N_8070,N_7631);
nand UO_423 (O_423,N_9428,N_7689);
and UO_424 (O_424,N_9838,N_9796);
and UO_425 (O_425,N_8672,N_9710);
or UO_426 (O_426,N_9170,N_7644);
or UO_427 (O_427,N_9153,N_8075);
xnor UO_428 (O_428,N_8061,N_9590);
or UO_429 (O_429,N_8202,N_8446);
xor UO_430 (O_430,N_9551,N_8217);
nor UO_431 (O_431,N_8033,N_8947);
nand UO_432 (O_432,N_8485,N_8034);
or UO_433 (O_433,N_8957,N_8273);
xor UO_434 (O_434,N_8658,N_7826);
nor UO_435 (O_435,N_7541,N_8368);
xor UO_436 (O_436,N_8689,N_8046);
or UO_437 (O_437,N_9619,N_9016);
nand UO_438 (O_438,N_8389,N_7931);
nor UO_439 (O_439,N_8417,N_8894);
and UO_440 (O_440,N_9735,N_9274);
or UO_441 (O_441,N_8843,N_9350);
and UO_442 (O_442,N_9727,N_8460);
and UO_443 (O_443,N_8491,N_9348);
nor UO_444 (O_444,N_9055,N_9396);
xor UO_445 (O_445,N_9777,N_8660);
xnor UO_446 (O_446,N_9117,N_9808);
and UO_447 (O_447,N_7690,N_7846);
or UO_448 (O_448,N_9141,N_9633);
xnor UO_449 (O_449,N_9625,N_7688);
nand UO_450 (O_450,N_7790,N_7744);
nor UO_451 (O_451,N_9822,N_8518);
or UO_452 (O_452,N_9951,N_8058);
and UO_453 (O_453,N_8220,N_9943);
or UO_454 (O_454,N_7992,N_9849);
or UO_455 (O_455,N_9441,N_7916);
or UO_456 (O_456,N_8294,N_9084);
or UO_457 (O_457,N_8645,N_8219);
or UO_458 (O_458,N_8707,N_9295);
and UO_459 (O_459,N_9275,N_9142);
nand UO_460 (O_460,N_8713,N_8992);
or UO_461 (O_461,N_8038,N_9698);
nand UO_462 (O_462,N_9131,N_8186);
or UO_463 (O_463,N_7754,N_9257);
nand UO_464 (O_464,N_8162,N_9758);
and UO_465 (O_465,N_8425,N_8830);
nand UO_466 (O_466,N_9826,N_8825);
nand UO_467 (O_467,N_9354,N_9812);
xor UO_468 (O_468,N_8434,N_8970);
and UO_469 (O_469,N_9774,N_9480);
and UO_470 (O_470,N_8101,N_8451);
and UO_471 (O_471,N_8826,N_8239);
nor UO_472 (O_472,N_8741,N_7682);
and UO_473 (O_473,N_8089,N_8958);
nor UO_474 (O_474,N_9713,N_7905);
nor UO_475 (O_475,N_9657,N_9554);
or UO_476 (O_476,N_7703,N_9059);
xor UO_477 (O_477,N_9082,N_7831);
xor UO_478 (O_478,N_9465,N_9011);
or UO_479 (O_479,N_8480,N_8692);
nand UO_480 (O_480,N_8542,N_7738);
nor UO_481 (O_481,N_9452,N_9645);
or UO_482 (O_482,N_8962,N_8916);
nand UO_483 (O_483,N_8737,N_9457);
nand UO_484 (O_484,N_8432,N_9555);
nand UO_485 (O_485,N_9439,N_8720);
nand UO_486 (O_486,N_8225,N_7619);
xnor UO_487 (O_487,N_9629,N_9269);
and UO_488 (O_488,N_7573,N_8561);
and UO_489 (O_489,N_9972,N_7620);
or UO_490 (O_490,N_9259,N_9454);
xnor UO_491 (O_491,N_7924,N_9151);
xnor UO_492 (O_492,N_9092,N_9595);
nand UO_493 (O_493,N_9327,N_7592);
nor UO_494 (O_494,N_8722,N_7965);
nor UO_495 (O_495,N_8869,N_8760);
or UO_496 (O_496,N_8009,N_9108);
and UO_497 (O_497,N_8387,N_8370);
nand UO_498 (O_498,N_9785,N_9397);
xnor UO_499 (O_499,N_7767,N_7684);
and UO_500 (O_500,N_8474,N_9638);
and UO_501 (O_501,N_8210,N_7936);
nor UO_502 (O_502,N_9373,N_9864);
nor UO_503 (O_503,N_9685,N_7845);
xnor UO_504 (O_504,N_9022,N_7616);
nor UO_505 (O_505,N_8686,N_8339);
nand UO_506 (O_506,N_8054,N_8527);
nor UO_507 (O_507,N_8949,N_8989);
or UO_508 (O_508,N_9285,N_8637);
nand UO_509 (O_509,N_8735,N_8102);
nor UO_510 (O_510,N_9715,N_8492);
xnor UO_511 (O_511,N_8165,N_8976);
nor UO_512 (O_512,N_9578,N_9977);
xor UO_513 (O_513,N_7588,N_8573);
xor UO_514 (O_514,N_8408,N_9692);
or UO_515 (O_515,N_7966,N_9426);
xor UO_516 (O_516,N_9154,N_9375);
nand UO_517 (O_517,N_9947,N_9208);
nor UO_518 (O_518,N_9541,N_8109);
nand UO_519 (O_519,N_9305,N_8226);
nor UO_520 (O_520,N_8685,N_9902);
nor UO_521 (O_521,N_8430,N_9495);
nor UO_522 (O_522,N_9764,N_8456);
nor UO_523 (O_523,N_7857,N_8514);
or UO_524 (O_524,N_8821,N_8517);
and UO_525 (O_525,N_8649,N_9381);
and UO_526 (O_526,N_7967,N_9739);
xor UO_527 (O_527,N_9752,N_8643);
nand UO_528 (O_528,N_8185,N_7873);
nand UO_529 (O_529,N_9103,N_9835);
and UO_530 (O_530,N_9640,N_8908);
xor UO_531 (O_531,N_9138,N_9845);
nor UO_532 (O_532,N_9349,N_9380);
xor UO_533 (O_533,N_9877,N_8232);
nor UO_534 (O_534,N_7877,N_9232);
nor UO_535 (O_535,N_7692,N_9312);
nor UO_536 (O_536,N_8774,N_7508);
xnor UO_537 (O_537,N_9210,N_9534);
or UO_538 (O_538,N_9895,N_7901);
and UO_539 (O_539,N_9163,N_9665);
nand UO_540 (O_540,N_9005,N_7591);
xnor UO_541 (O_541,N_7567,N_9281);
nand UO_542 (O_542,N_9169,N_7887);
nor UO_543 (O_543,N_8714,N_7731);
and UO_544 (O_544,N_7708,N_8986);
or UO_545 (O_545,N_9184,N_9773);
nand UO_546 (O_546,N_8361,N_9929);
or UO_547 (O_547,N_7668,N_9725);
nand UO_548 (O_548,N_9464,N_9419);
and UO_549 (O_549,N_7794,N_8726);
nand UO_550 (O_550,N_7517,N_9335);
nand UO_551 (O_551,N_8001,N_7878);
nor UO_552 (O_552,N_9565,N_9795);
nand UO_553 (O_553,N_7893,N_8762);
or UO_554 (O_554,N_9253,N_7664);
or UO_555 (O_555,N_8678,N_7529);
xor UO_556 (O_556,N_7888,N_7808);
or UO_557 (O_557,N_8885,N_9987);
xnor UO_558 (O_558,N_9000,N_8983);
nor UO_559 (O_559,N_8927,N_8012);
xor UO_560 (O_560,N_8708,N_9532);
nor UO_561 (O_561,N_7615,N_7720);
nor UO_562 (O_562,N_7628,N_7747);
or UO_563 (O_563,N_8756,N_8642);
or UO_564 (O_564,N_7938,N_9883);
nor UO_565 (O_565,N_9252,N_8126);
and UO_566 (O_566,N_9475,N_9757);
or UO_567 (O_567,N_8052,N_7653);
nand UO_568 (O_568,N_8874,N_9292);
nor UO_569 (O_569,N_8449,N_8390);
and UO_570 (O_570,N_9168,N_9591);
and UO_571 (O_571,N_8779,N_8245);
nor UO_572 (O_572,N_9078,N_8555);
xnor UO_573 (O_573,N_8381,N_8036);
xor UO_574 (O_574,N_9697,N_8964);
xnor UO_575 (O_575,N_9604,N_8693);
nor UO_576 (O_576,N_7526,N_9144);
nand UO_577 (O_577,N_8764,N_8107);
or UO_578 (O_578,N_9866,N_9760);
and UO_579 (O_579,N_8157,N_9973);
or UO_580 (O_580,N_9355,N_8950);
nor UO_581 (O_581,N_8968,N_9160);
or UO_582 (O_582,N_9043,N_8783);
xor UO_583 (O_583,N_8215,N_7928);
and UO_584 (O_584,N_9291,N_9481);
nor UO_585 (O_585,N_8510,N_9217);
nand UO_586 (O_586,N_9155,N_9026);
xor UO_587 (O_587,N_9813,N_7944);
nor UO_588 (O_588,N_9331,N_8704);
and UO_589 (O_589,N_8937,N_7551);
nor UO_590 (O_590,N_9881,N_8171);
xnor UO_591 (O_591,N_9136,N_9272);
or UO_592 (O_592,N_8880,N_8772);
and UO_593 (O_593,N_7521,N_7895);
or UO_594 (O_594,N_8422,N_7504);
or UO_595 (O_595,N_7600,N_9105);
and UO_596 (O_596,N_9128,N_9411);
nor UO_597 (O_597,N_8503,N_8788);
or UO_598 (O_598,N_9925,N_7638);
and UO_599 (O_599,N_9501,N_8864);
and UO_600 (O_600,N_9107,N_9420);
nor UO_601 (O_601,N_8172,N_9158);
nor UO_602 (O_602,N_8780,N_8807);
and UO_603 (O_603,N_8694,N_9539);
or UO_604 (O_604,N_8104,N_8330);
xor UO_605 (O_605,N_9081,N_9407);
and UO_606 (O_606,N_7998,N_8935);
or UO_607 (O_607,N_9063,N_9164);
nand UO_608 (O_608,N_8670,N_9749);
or UO_609 (O_609,N_9140,N_8652);
xor UO_610 (O_610,N_9842,N_9690);
nor UO_611 (O_611,N_9594,N_8164);
nor UO_612 (O_612,N_7779,N_8360);
or UO_613 (O_613,N_8209,N_9876);
and UO_614 (O_614,N_9047,N_8675);
xnor UO_615 (O_615,N_8110,N_9584);
nor UO_616 (O_616,N_9948,N_7640);
and UO_617 (O_617,N_8384,N_9422);
nor UO_618 (O_618,N_8301,N_8299);
xor UO_619 (O_619,N_8834,N_8926);
nand UO_620 (O_620,N_9280,N_9361);
xnor UO_621 (O_621,N_9743,N_8183);
or UO_622 (O_622,N_9507,N_8501);
xor UO_623 (O_623,N_8529,N_9266);
and UO_624 (O_624,N_9463,N_9201);
and UO_625 (O_625,N_7884,N_8005);
or UO_626 (O_626,N_8860,N_8856);
and UO_627 (O_627,N_9122,N_8815);
nor UO_628 (O_628,N_7902,N_8068);
xnor UO_629 (O_629,N_7523,N_9041);
xor UO_630 (O_630,N_8438,N_8458);
or UO_631 (O_631,N_9284,N_8850);
or UO_632 (O_632,N_9726,N_8382);
or UO_633 (O_633,N_9733,N_8822);
and UO_634 (O_634,N_8702,N_9477);
or UO_635 (O_635,N_8519,N_9717);
nor UO_636 (O_636,N_9237,N_9601);
nor UO_637 (O_637,N_7676,N_7892);
xnor UO_638 (O_638,N_8132,N_7756);
nor UO_639 (O_639,N_9231,N_8402);
nor UO_640 (O_640,N_9320,N_9015);
xnor UO_641 (O_641,N_7535,N_7732);
and UO_642 (O_642,N_9994,N_8011);
nor UO_643 (O_643,N_9630,N_8802);
nand UO_644 (O_644,N_9675,N_8548);
and UO_645 (O_645,N_9990,N_7991);
and UO_646 (O_646,N_8946,N_8999);
xor UO_647 (O_647,N_8169,N_8631);
and UO_648 (O_648,N_8045,N_9514);
or UO_649 (O_649,N_8981,N_9526);
and UO_650 (O_650,N_8249,N_8775);
xor UO_651 (O_651,N_9276,N_9802);
or UO_652 (O_652,N_9067,N_8048);
and UO_653 (O_653,N_8570,N_8086);
nor UO_654 (O_654,N_8791,N_8657);
or UO_655 (O_655,N_7978,N_8420);
or UO_656 (O_656,N_8306,N_8921);
and UO_657 (O_657,N_9557,N_8468);
nor UO_658 (O_658,N_9899,N_8823);
or UO_659 (O_659,N_9639,N_8540);
or UO_660 (O_660,N_9365,N_9856);
xor UO_661 (O_661,N_8782,N_8721);
and UO_662 (O_662,N_8571,N_7590);
nor UO_663 (O_663,N_8604,N_9006);
and UO_664 (O_664,N_7656,N_9363);
nor UO_665 (O_665,N_8936,N_8008);
nor UO_666 (O_666,N_8795,N_8598);
xor UO_667 (O_667,N_8004,N_8902);
or UO_668 (O_668,N_9886,N_7933);
and UO_669 (O_669,N_9264,N_7558);
and UO_670 (O_670,N_7999,N_8088);
nand UO_671 (O_671,N_7961,N_9801);
xnor UO_672 (O_672,N_8365,N_8098);
and UO_673 (O_673,N_7699,N_7852);
xnor UO_674 (O_674,N_7858,N_9549);
and UO_675 (O_675,N_9221,N_7539);
nand UO_676 (O_676,N_8450,N_9966);
and UO_677 (O_677,N_7948,N_7837);
and UO_678 (O_678,N_9724,N_9848);
or UO_679 (O_679,N_7940,N_9434);
or UO_680 (O_680,N_9148,N_9146);
nor UO_681 (O_681,N_8663,N_9069);
nor UO_682 (O_682,N_8396,N_9461);
and UO_683 (O_683,N_8409,N_7613);
nor UO_684 (O_684,N_8398,N_8595);
nor UO_685 (O_685,N_7721,N_9666);
nor UO_686 (O_686,N_8060,N_8816);
nor UO_687 (O_687,N_9035,N_9300);
or UO_688 (O_688,N_9258,N_8277);
nor UO_689 (O_689,N_8928,N_8803);
xnor UO_690 (O_690,N_9012,N_8499);
or UO_691 (O_691,N_7950,N_7886);
xor UO_692 (O_692,N_9819,N_8493);
or UO_693 (O_693,N_9921,N_9197);
xor UO_694 (O_694,N_9621,N_8687);
and UO_695 (O_695,N_8603,N_9333);
nor UO_696 (O_696,N_9911,N_8617);
and UO_697 (O_697,N_8543,N_9244);
and UO_698 (O_698,N_8016,N_9427);
or UO_699 (O_699,N_9857,N_7506);
and UO_700 (O_700,N_9204,N_7972);
nand UO_701 (O_701,N_9296,N_9548);
or UO_702 (O_702,N_7899,N_9393);
nor UO_703 (O_703,N_9459,N_8349);
nor UO_704 (O_704,N_7809,N_9106);
or UO_705 (O_705,N_7728,N_8757);
nand UO_706 (O_706,N_9632,N_7714);
and UO_707 (O_707,N_8796,N_9919);
and UO_708 (O_708,N_8808,N_9384);
nand UO_709 (O_709,N_8413,N_7512);
nor UO_710 (O_710,N_8153,N_9882);
nand UO_711 (O_711,N_9771,N_9714);
nor UO_712 (O_712,N_9828,N_7630);
xnor UO_713 (O_713,N_8963,N_9867);
and UO_714 (O_714,N_7943,N_7898);
or UO_715 (O_715,N_8244,N_8911);
or UO_716 (O_716,N_7959,N_8050);
and UO_717 (O_717,N_9915,N_8700);
nor UO_718 (O_718,N_8071,N_9423);
or UO_719 (O_719,N_8125,N_8806);
and UO_720 (O_720,N_8884,N_8690);
nor UO_721 (O_721,N_9229,N_9062);
and UO_722 (O_722,N_9614,N_9515);
nor UO_723 (O_723,N_9776,N_9793);
or UO_724 (O_724,N_8750,N_9079);
nand UO_725 (O_725,N_8614,N_8111);
xor UO_726 (O_726,N_8959,N_9342);
and UO_727 (O_727,N_9308,N_9173);
nand UO_728 (O_728,N_9357,N_7818);
or UO_729 (O_729,N_8876,N_7667);
xnor UO_730 (O_730,N_9672,N_9037);
nor UO_731 (O_731,N_9543,N_7872);
xnor UO_732 (O_732,N_9694,N_8108);
and UO_733 (O_733,N_9897,N_7832);
xnor UO_734 (O_734,N_8292,N_8083);
nand UO_735 (O_735,N_7576,N_8087);
nor UO_736 (O_736,N_8404,N_9064);
xnor UO_737 (O_737,N_9021,N_7654);
xor UO_738 (O_738,N_9833,N_8279);
xor UO_739 (O_739,N_8237,N_8740);
or UO_740 (O_740,N_9306,N_8618);
and UO_741 (O_741,N_7625,N_7870);
xnor UO_742 (O_742,N_8801,N_8619);
nand UO_743 (O_743,N_7587,N_8179);
and UO_744 (O_744,N_8691,N_9870);
xor UO_745 (O_745,N_9738,N_7941);
nand UO_746 (O_746,N_9329,N_9191);
xor UO_747 (O_747,N_7565,N_9165);
or UO_748 (O_748,N_8133,N_8688);
xor UO_749 (O_749,N_8281,N_9377);
xnor UO_750 (O_750,N_8730,N_9846);
nand UO_751 (O_751,N_8967,N_8247);
or UO_752 (O_752,N_7982,N_8295);
nand UO_753 (O_753,N_8161,N_8167);
nand UO_754 (O_754,N_7641,N_9517);
xnor UO_755 (O_755,N_9528,N_8890);
xnor UO_756 (O_756,N_9686,N_9931);
xor UO_757 (O_757,N_9946,N_9326);
nand UO_758 (O_758,N_7988,N_9424);
nor UO_759 (O_759,N_9178,N_9784);
nand UO_760 (O_760,N_8293,N_9737);
or UO_761 (O_761,N_7757,N_8421);
nor UO_762 (O_762,N_8322,N_7610);
xnor UO_763 (O_763,N_7990,N_8336);
or UO_764 (O_764,N_7635,N_8995);
nor UO_765 (O_765,N_8812,N_9290);
nor UO_766 (O_766,N_8567,N_9110);
or UO_767 (O_767,N_7629,N_9707);
or UO_768 (O_768,N_9056,N_9982);
nand UO_769 (O_769,N_9198,N_8216);
nand UO_770 (O_770,N_7718,N_9183);
nor UO_771 (O_771,N_7798,N_8206);
nor UO_772 (O_772,N_7704,N_9446);
or UO_773 (O_773,N_8930,N_7540);
nor UO_774 (O_774,N_9044,N_8578);
nand UO_775 (O_775,N_9486,N_8507);
nand UO_776 (O_776,N_9663,N_9492);
nor UO_777 (O_777,N_7766,N_9798);
and UO_778 (O_778,N_8074,N_9635);
or UO_779 (O_779,N_8175,N_9789);
nor UO_780 (O_780,N_8137,N_9781);
nand UO_781 (O_781,N_8723,N_9564);
nand UO_782 (O_782,N_8289,N_7621);
or UO_783 (O_783,N_8905,N_9611);
and UO_784 (O_784,N_8629,N_7825);
or UO_785 (O_785,N_7753,N_9072);
or UO_786 (O_786,N_8415,N_9212);
nor UO_787 (O_787,N_9924,N_9907);
nor UO_788 (O_788,N_8883,N_8917);
or UO_789 (O_789,N_7678,N_9880);
nand UO_790 (O_790,N_9444,N_7705);
xnor UO_791 (O_791,N_8040,N_8521);
and UO_792 (O_792,N_8112,N_9023);
or UO_793 (O_793,N_7934,N_9509);
nand UO_794 (O_794,N_8748,N_9202);
xnor UO_795 (O_795,N_9224,N_9579);
and UO_796 (O_796,N_9778,N_9871);
nor UO_797 (O_797,N_8638,N_9398);
nor UO_798 (O_798,N_9592,N_9898);
xor UO_799 (O_799,N_8952,N_9945);
nor UO_800 (O_800,N_9818,N_9585);
nand UO_801 (O_801,N_8659,N_9920);
nand UO_802 (O_802,N_7911,N_9199);
or UO_803 (O_803,N_8093,N_8442);
xnor UO_804 (O_804,N_7939,N_8258);
xnor UO_805 (O_805,N_7782,N_9293);
nor UO_806 (O_806,N_8305,N_7581);
or UO_807 (O_807,N_8476,N_8551);
xor UO_808 (O_808,N_8800,N_9404);
xor UO_809 (O_809,N_9352,N_9347);
or UO_810 (O_810,N_9159,N_9050);
xor UO_811 (O_811,N_9025,N_7841);
and UO_812 (O_812,N_8188,N_8313);
nor UO_813 (O_813,N_9310,N_8754);
or UO_814 (O_814,N_9358,N_8733);
and UO_815 (O_815,N_9786,N_7827);
and UO_816 (O_816,N_8486,N_8848);
nand UO_817 (O_817,N_9647,N_7595);
or UO_818 (O_818,N_9668,N_7605);
nor UO_819 (O_819,N_7575,N_9130);
xnor UO_820 (O_820,N_9641,N_7976);
xor UO_821 (O_821,N_7723,N_9294);
nand UO_822 (O_822,N_8031,N_8520);
nand UO_823 (O_823,N_8781,N_9120);
or UO_824 (O_824,N_8291,N_8265);
xor UO_825 (O_825,N_8565,N_8067);
xor UO_826 (O_826,N_9345,N_8027);
or UO_827 (O_827,N_9817,N_8128);
nand UO_828 (O_828,N_8505,N_7673);
xnor UO_829 (O_829,N_8024,N_9524);
nor UO_830 (O_830,N_9976,N_8847);
nand UO_831 (O_831,N_8025,N_7661);
and UO_832 (O_832,N_8502,N_8915);
nor UO_833 (O_833,N_9719,N_9473);
nor UO_834 (O_834,N_9086,N_8602);
xor UO_835 (O_835,N_9455,N_8984);
and UO_836 (O_836,N_8072,N_8190);
or UO_837 (O_837,N_7807,N_7701);
nor UO_838 (O_838,N_9705,N_8214);
nand UO_839 (O_839,N_8965,N_8079);
nor UO_840 (O_840,N_9097,N_8334);
nor UO_841 (O_841,N_9094,N_8934);
and UO_842 (O_842,N_8960,N_7652);
or UO_843 (O_843,N_9740,N_8037);
xnor UO_844 (O_844,N_8479,N_9322);
nand UO_845 (O_845,N_7927,N_9301);
or UO_846 (O_846,N_8552,N_9496);
or UO_847 (O_847,N_9901,N_7819);
nand UO_848 (O_848,N_8049,N_7788);
nor UO_849 (O_849,N_8938,N_9406);
nand UO_850 (O_850,N_7636,N_8715);
nor UO_851 (O_851,N_8597,N_8589);
or UO_852 (O_852,N_9193,N_7955);
or UO_853 (O_853,N_8285,N_7848);
nor UO_854 (O_854,N_8378,N_9469);
nor UO_855 (O_855,N_9440,N_7979);
nor UO_856 (O_856,N_9596,N_9417);
nor UO_857 (O_857,N_8622,N_9392);
nor UO_858 (O_858,N_8913,N_8674);
nand UO_859 (O_859,N_8392,N_9926);
or UO_860 (O_860,N_7646,N_8910);
xor UO_861 (O_861,N_8394,N_8901);
or UO_862 (O_862,N_9177,N_9805);
and UO_863 (O_863,N_9746,N_9482);
nor UO_864 (O_864,N_8340,N_8703);
and UO_865 (O_865,N_9847,N_9561);
xnor UO_866 (O_866,N_9616,N_9658);
nor UO_867 (O_867,N_8022,N_8745);
and UO_868 (O_868,N_8625,N_9483);
xor UO_869 (O_869,N_9797,N_8654);
nor UO_870 (O_870,N_8081,N_9251);
nand UO_871 (O_871,N_7932,N_7797);
xor UO_872 (O_872,N_9811,N_9019);
xnor UO_873 (O_873,N_7772,N_8268);
or UO_874 (O_874,N_9851,N_8343);
nor UO_875 (O_875,N_7786,N_7796);
or UO_876 (O_876,N_8839,N_8260);
or UO_877 (O_877,N_9965,N_7729);
nor UO_878 (O_878,N_8798,N_9974);
or UO_879 (O_879,N_8831,N_9311);
and UO_880 (O_880,N_9338,N_7715);
and UO_881 (O_881,N_9216,N_8276);
or UO_882 (O_882,N_8145,N_8919);
xor UO_883 (O_883,N_9544,N_7956);
nor UO_884 (O_884,N_9325,N_8325);
and UO_885 (O_885,N_8263,N_9704);
or UO_886 (O_886,N_9979,N_7904);
or UO_887 (O_887,N_8466,N_7549);
nor UO_888 (O_888,N_9803,N_7751);
or UO_889 (O_889,N_9552,N_9967);
xor UO_890 (O_890,N_8170,N_7824);
and UO_891 (O_891,N_8374,N_8262);
and UO_892 (O_892,N_9289,N_9395);
and UO_893 (O_893,N_7516,N_9661);
xor UO_894 (O_894,N_9997,N_9950);
and UO_895 (O_895,N_9815,N_8793);
xor UO_896 (O_896,N_8512,N_9571);
nor UO_897 (O_897,N_7971,N_8893);
nor UO_898 (O_898,N_8199,N_8035);
xor UO_899 (O_899,N_9577,N_7983);
nand UO_900 (O_900,N_8114,N_7502);
nor UO_901 (O_901,N_9124,N_9910);
or UO_902 (O_902,N_7524,N_9503);
xnor UO_903 (O_903,N_9256,N_9189);
or UO_904 (O_904,N_8391,N_7806);
nor UO_905 (O_905,N_8767,N_8827);
xnor UO_906 (O_906,N_9655,N_8506);
nand UO_907 (O_907,N_9476,N_8021);
nor UO_908 (O_908,N_9096,N_9918);
nor UO_909 (O_909,N_7632,N_8489);
nor UO_910 (O_910,N_8065,N_9605);
and UO_911 (O_911,N_9319,N_8174);
nor UO_912 (O_912,N_7816,N_7622);
xnor UO_913 (O_913,N_7871,N_9829);
or UO_914 (O_914,N_8191,N_8572);
nand UO_915 (O_915,N_9748,N_8149);
nor UO_916 (O_916,N_9077,N_9186);
nor UO_917 (O_917,N_9531,N_9703);
xnor UO_918 (O_918,N_9820,N_7651);
nor UO_919 (O_919,N_9250,N_9241);
and UO_920 (O_920,N_8453,N_8388);
nor UO_921 (O_921,N_9642,N_8941);
or UO_922 (O_922,N_8644,N_9583);
xor UO_923 (O_923,N_8853,N_7606);
and UO_924 (O_924,N_9708,N_9917);
xnor UO_925 (O_925,N_7659,N_9606);
nor UO_926 (O_926,N_8866,N_9836);
xor UO_927 (O_927,N_8755,N_7589);
xor UO_928 (O_928,N_9513,N_7608);
or UO_929 (O_929,N_8627,N_9129);
nand UO_930 (O_930,N_8116,N_9736);
nor UO_931 (O_931,N_8419,N_9550);
and UO_932 (O_932,N_8861,N_9954);
xnor UO_933 (O_933,N_8317,N_8945);
nor UO_934 (O_934,N_8401,N_8842);
or UO_935 (O_935,N_9009,N_8218);
nand UO_936 (O_936,N_9181,N_8241);
and UO_937 (O_937,N_9839,N_8307);
nand UO_938 (O_938,N_9790,N_8569);
nor UO_939 (O_939,N_8841,N_8152);
nand UO_940 (O_940,N_8594,N_9878);
or UO_941 (O_941,N_9121,N_9618);
xnor UO_942 (O_942,N_9652,N_7566);
and UO_943 (O_943,N_8797,N_9213);
and UO_944 (O_944,N_9788,N_9039);
xnor UO_945 (O_945,N_7859,N_9662);
nand UO_946 (O_946,N_8494,N_8337);
nand UO_947 (O_947,N_9834,N_9593);
xor UO_948 (O_948,N_8030,N_8238);
xor UO_949 (O_949,N_9568,N_9841);
or UO_950 (O_950,N_9315,N_7866);
xnor UO_951 (O_951,N_8189,N_8423);
and UO_952 (O_952,N_7722,N_9728);
or UO_953 (O_953,N_8609,N_8531);
nand UO_954 (O_954,N_8371,N_8197);
nor UO_955 (O_955,N_8182,N_9783);
xor UO_956 (O_956,N_9498,N_7799);
or UO_957 (O_957,N_7996,N_7719);
or UO_958 (O_958,N_9782,N_8407);
and UO_959 (O_959,N_8405,N_9624);
or UO_960 (O_960,N_8676,N_8786);
nand UO_961 (O_961,N_9449,N_7964);
nand UO_962 (O_962,N_9850,N_8117);
and UO_963 (O_963,N_9179,N_8130);
or UO_964 (O_964,N_8303,N_8156);
nor UO_965 (O_965,N_9304,N_7785);
and UO_966 (O_966,N_7706,N_8819);
and UO_967 (O_967,N_7907,N_9205);
and UO_968 (O_968,N_7802,N_7725);
or UO_969 (O_969,N_8084,N_7856);
nand UO_970 (O_970,N_9225,N_9418);
nor UO_971 (O_971,N_9214,N_8898);
nand UO_972 (O_972,N_7913,N_8718);
and UO_973 (O_973,N_8284,N_9597);
xnor UO_974 (O_974,N_9516,N_9916);
or UO_975 (O_975,N_8538,N_8321);
nand UO_976 (O_976,N_7623,N_9490);
nor UO_977 (O_977,N_8865,N_7930);
or UO_978 (O_978,N_8743,N_8809);
or UO_979 (O_979,N_9667,N_9001);
or UO_980 (O_980,N_8155,N_7509);
xnor UO_981 (O_981,N_9472,N_8533);
nor UO_982 (O_982,N_7891,N_9537);
nor UO_983 (O_983,N_8684,N_8765);
xnor UO_984 (O_984,N_9471,N_8455);
or UO_985 (O_985,N_7553,N_9889);
xnor UO_986 (O_986,N_8055,N_7780);
and UO_987 (O_987,N_8653,N_7793);
or UO_988 (O_988,N_9891,N_9100);
nor UO_989 (O_989,N_9379,N_8558);
and UO_990 (O_990,N_9187,N_8914);
nor UO_991 (O_991,N_9068,N_8639);
or UO_992 (O_992,N_8525,N_8090);
nor UO_993 (O_993,N_9637,N_9569);
xnor UO_994 (O_994,N_9750,N_7836);
and UO_995 (O_995,N_9389,N_8593);
nor UO_996 (O_996,N_7533,N_9981);
nand UO_997 (O_997,N_9613,N_9992);
nand UO_998 (O_998,N_9053,N_9688);
nand UO_999 (O_999,N_7918,N_9807);
nor UO_1000 (O_1000,N_7969,N_7986);
nor UO_1001 (O_1001,N_7985,N_8682);
xor UO_1002 (O_1002,N_9955,N_9367);
or UO_1003 (O_1003,N_8867,N_9673);
and UO_1004 (O_1004,N_7642,N_9511);
xnor UO_1005 (O_1005,N_8557,N_8857);
nor UO_1006 (O_1006,N_7889,N_7528);
or UO_1007 (O_1007,N_7599,N_8810);
or UO_1008 (O_1008,N_7771,N_7970);
xnor UO_1009 (O_1009,N_9861,N_8634);
nand UO_1010 (O_1010,N_7851,N_9222);
or UO_1011 (O_1011,N_9362,N_7624);
nand UO_1012 (O_1012,N_9923,N_7953);
and UO_1013 (O_1013,N_7839,N_9057);
or UO_1014 (O_1014,N_8787,N_9134);
nor UO_1015 (O_1015,N_7849,N_9587);
nand UO_1016 (O_1016,N_7683,N_9371);
xor UO_1017 (O_1017,N_7716,N_7607);
xnor UO_1018 (O_1018,N_9466,N_8416);
or UO_1019 (O_1019,N_8376,N_8066);
and UO_1020 (O_1020,N_9233,N_9052);
or UO_1021 (O_1021,N_8366,N_7662);
or UO_1022 (O_1022,N_8975,N_7677);
nand UO_1023 (O_1023,N_8251,N_9659);
or UO_1024 (O_1024,N_7752,N_8662);
or UO_1025 (O_1025,N_8148,N_8495);
or UO_1026 (O_1026,N_7717,N_7594);
and UO_1027 (O_1027,N_7912,N_9336);
or UO_1028 (O_1028,N_8375,N_8892);
nand UO_1029 (O_1029,N_8719,N_9560);
or UO_1030 (O_1030,N_9933,N_7650);
nor UO_1031 (O_1031,N_9734,N_8990);
nor UO_1032 (O_1032,N_8600,N_8103);
xor UO_1033 (O_1033,N_8323,N_8379);
and UO_1034 (O_1034,N_9504,N_8724);
xnor UO_1035 (O_1035,N_7582,N_7770);
nand UO_1036 (O_1036,N_9711,N_9868);
nand UO_1037 (O_1037,N_9766,N_9003);
or UO_1038 (O_1038,N_9317,N_8697);
nor UO_1039 (O_1039,N_7527,N_8646);
and UO_1040 (O_1040,N_8544,N_9234);
nor UO_1041 (O_1041,N_8922,N_9909);
xnor UO_1042 (O_1042,N_8972,N_9209);
nand UO_1043 (O_1043,N_9421,N_8064);
nor UO_1044 (O_1044,N_8248,N_8463);
and UO_1045 (O_1045,N_8257,N_9448);
nor UO_1046 (O_1046,N_9058,N_7840);
nand UO_1047 (O_1047,N_7602,N_9157);
nand UO_1048 (O_1048,N_8858,N_9988);
nor UO_1049 (O_1049,N_9046,N_8280);
xor UO_1050 (O_1050,N_8868,N_9643);
nand UO_1051 (O_1051,N_8881,N_7570);
or UO_1052 (O_1052,N_8628,N_7814);
xor UO_1053 (O_1053,N_9800,N_8789);
nor UO_1054 (O_1054,N_8923,N_9983);
and UO_1055 (O_1055,N_9090,N_8469);
or UO_1056 (O_1056,N_8275,N_7614);
nor UO_1057 (O_1057,N_8840,N_9620);
nor UO_1058 (O_1058,N_8899,N_8805);
nor UO_1059 (O_1059,N_8630,N_8575);
and UO_1060 (O_1060,N_8624,N_7813);
nand UO_1061 (O_1061,N_9575,N_8020);
and UO_1062 (O_1062,N_7739,N_7597);
and UO_1063 (O_1063,N_9706,N_9900);
nor UO_1064 (O_1064,N_9765,N_9612);
and UO_1065 (O_1065,N_8129,N_9374);
nand UO_1066 (O_1066,N_9664,N_8532);
nand UO_1067 (O_1067,N_7980,N_9745);
nand UO_1068 (O_1068,N_8042,N_8242);
and UO_1069 (O_1069,N_9518,N_9484);
nor UO_1070 (O_1070,N_8583,N_8711);
nand UO_1071 (O_1071,N_7536,N_9723);
nand UO_1072 (O_1072,N_8229,N_9321);
or UO_1073 (O_1073,N_8359,N_7572);
nand UO_1074 (O_1074,N_8424,N_8097);
xor UO_1075 (O_1075,N_9149,N_9602);
or UO_1076 (O_1076,N_8429,N_7921);
or UO_1077 (O_1077,N_8592,N_8457);
or UO_1078 (O_1078,N_7666,N_9175);
nand UO_1079 (O_1079,N_7585,N_8100);
nor UO_1080 (O_1080,N_9631,N_8272);
nor UO_1081 (O_1081,N_9553,N_9013);
nand UO_1082 (O_1082,N_9957,N_8664);
or UO_1083 (O_1083,N_7550,N_8351);
nand UO_1084 (O_1084,N_9386,N_7922);
and UO_1085 (O_1085,N_9831,N_9038);
and UO_1086 (O_1086,N_8545,N_7865);
or UO_1087 (O_1087,N_7519,N_8308);
nand UO_1088 (O_1088,N_9030,N_9930);
nor UO_1089 (O_1089,N_7789,N_9751);
xor UO_1090 (O_1090,N_8846,N_8877);
and UO_1091 (O_1091,N_8267,N_9116);
xnor UO_1092 (O_1092,N_8920,N_7769);
nand UO_1093 (O_1093,N_9932,N_9615);
nor UO_1094 (O_1094,N_9779,N_9220);
and UO_1095 (O_1095,N_7781,N_8362);
nor UO_1096 (O_1096,N_8380,N_9687);
xor UO_1097 (O_1097,N_9677,N_7681);
or UO_1098 (O_1098,N_8854,N_8047);
xnor UO_1099 (O_1099,N_8227,N_7586);
xnor UO_1100 (O_1100,N_7821,N_9996);
and UO_1101 (O_1101,N_9617,N_7758);
and UO_1102 (O_1102,N_8615,N_8699);
xnor UO_1103 (O_1103,N_8297,N_8338);
nor UO_1104 (O_1104,N_9353,N_9203);
or UO_1105 (O_1105,N_8886,N_7787);
xnor UO_1106 (O_1106,N_9660,N_8270);
xnor UO_1107 (O_1107,N_8804,N_9806);
nand UO_1108 (O_1108,N_9855,N_8633);
nand UO_1109 (O_1109,N_7875,N_9113);
nand UO_1110 (O_1110,N_7674,N_7951);
xnor UO_1111 (O_1111,N_8481,N_9207);
xnor UO_1112 (O_1112,N_7734,N_8725);
and UO_1113 (O_1113,N_9126,N_9450);
nor UO_1114 (O_1114,N_8785,N_9195);
and UO_1115 (O_1115,N_8331,N_9194);
nand UO_1116 (O_1116,N_8124,N_9368);
xnor UO_1117 (O_1117,N_9447,N_9387);
and UO_1118 (O_1118,N_8168,N_9538);
or UO_1119 (O_1119,N_9339,N_9279);
nand UO_1120 (O_1120,N_9603,N_7947);
and UO_1121 (O_1121,N_9753,N_8044);
nand UO_1122 (O_1122,N_8669,N_8829);
or UO_1123 (O_1123,N_8608,N_8193);
and UO_1124 (O_1124,N_8073,N_7577);
xor UO_1125 (O_1125,N_7515,N_9478);
and UO_1126 (O_1126,N_9416,N_9732);
nand UO_1127 (O_1127,N_7727,N_8584);
and UO_1128 (O_1128,N_8944,N_8508);
xnor UO_1129 (O_1129,N_9431,N_9249);
nor UO_1130 (O_1130,N_9691,N_7915);
or UO_1131 (O_1131,N_8896,N_7505);
or UO_1132 (O_1132,N_7514,N_7724);
nor UO_1133 (O_1133,N_8369,N_8956);
nand UO_1134 (O_1134,N_7822,N_9430);
xor UO_1135 (O_1135,N_7897,N_8650);
xnor UO_1136 (O_1136,N_8385,N_9313);
or UO_1137 (O_1137,N_7847,N_9863);
nand UO_1138 (O_1138,N_9145,N_7559);
xor UO_1139 (O_1139,N_8204,N_9502);
xnor UO_1140 (O_1140,N_9042,N_8496);
xor UO_1141 (O_1141,N_9962,N_8879);
xnor UO_1142 (O_1142,N_7795,N_9860);
xnor UO_1143 (O_1143,N_9413,N_8470);
nand UO_1144 (O_1144,N_9462,N_9609);
and UO_1145 (O_1145,N_9679,N_8159);
or UO_1146 (O_1146,N_7835,N_9206);
nor UO_1147 (O_1147,N_8490,N_8014);
or UO_1148 (O_1148,N_8298,N_9944);
xor UO_1149 (O_1149,N_8192,N_9200);
or UO_1150 (O_1150,N_9008,N_8151);
and UO_1151 (O_1151,N_8991,N_9344);
or UO_1152 (O_1152,N_7562,N_8736);
and UO_1153 (O_1153,N_9875,N_9114);
or UO_1154 (O_1154,N_8728,N_7665);
nor UO_1155 (O_1155,N_7917,N_9034);
xor UO_1156 (O_1156,N_8418,N_9227);
nor UO_1157 (O_1157,N_9267,N_9188);
xor UO_1158 (O_1158,N_7778,N_9270);
nand UO_1159 (O_1159,N_9002,N_9567);
or UO_1160 (O_1160,N_7737,N_8763);
nor UO_1161 (O_1161,N_8851,N_8537);
and UO_1162 (O_1162,N_9488,N_8099);
nand UO_1163 (O_1163,N_7885,N_8683);
nor UO_1164 (O_1164,N_8095,N_8488);
nand UO_1165 (O_1165,N_7830,N_7713);
nor UO_1166 (O_1166,N_7634,N_8982);
nand UO_1167 (O_1167,N_7860,N_9425);
and UO_1168 (O_1168,N_9626,N_8018);
or UO_1169 (O_1169,N_9366,N_9489);
nand UO_1170 (O_1170,N_7702,N_8716);
or UO_1171 (O_1171,N_7709,N_8588);
nor UO_1172 (O_1172,N_9017,N_9161);
xor UO_1173 (O_1173,N_7764,N_8252);
and UO_1174 (O_1174,N_7867,N_7649);
or UO_1175 (O_1175,N_8792,N_9986);
xnor UO_1176 (O_1176,N_8000,N_8581);
or UO_1177 (O_1177,N_9061,N_9246);
and UO_1178 (O_1178,N_9680,N_8744);
or UO_1179 (O_1179,N_7557,N_7863);
nor UO_1180 (O_1180,N_8933,N_9702);
and UO_1181 (O_1181,N_9093,N_8668);
or UO_1182 (O_1182,N_9654,N_8749);
or UO_1183 (O_1183,N_9409,N_8302);
or UO_1184 (O_1184,N_9816,N_9627);
and UO_1185 (O_1185,N_9273,N_8118);
xor UO_1186 (O_1186,N_7697,N_9521);
nor UO_1187 (O_1187,N_7975,N_9118);
or UO_1188 (O_1188,N_8264,N_9133);
nand UO_1189 (O_1189,N_8367,N_8142);
and UO_1190 (O_1190,N_9343,N_8002);
nor UO_1191 (O_1191,N_9573,N_8342);
xnor UO_1192 (O_1192,N_7745,N_8222);
or UO_1193 (O_1193,N_8969,N_8445);
and UO_1194 (O_1194,N_7530,N_8013);
and UO_1195 (O_1195,N_8433,N_9852);
xor UO_1196 (O_1196,N_8352,N_8553);
or UO_1197 (O_1197,N_9412,N_7548);
nand UO_1198 (O_1198,N_8444,N_7762);
and UO_1199 (O_1199,N_8612,N_8742);
nand UO_1200 (O_1200,N_9589,N_9562);
and UO_1201 (O_1201,N_7648,N_8439);
xor UO_1202 (O_1202,N_9768,N_9741);
nand UO_1203 (O_1203,N_7906,N_9445);
nor UO_1204 (O_1204,N_8621,N_8076);
nor UO_1205 (O_1205,N_7730,N_9701);
nand UO_1206 (O_1206,N_8314,N_7695);
nor UO_1207 (O_1207,N_8461,N_7611);
or UO_1208 (O_1208,N_7564,N_8440);
or UO_1209 (O_1209,N_8269,N_8163);
and UO_1210 (O_1210,N_9824,N_8606);
or UO_1211 (O_1211,N_9091,N_7981);
nor UO_1212 (O_1212,N_8729,N_8304);
and UO_1213 (O_1213,N_9546,N_7501);
nor UO_1214 (O_1214,N_7862,N_7946);
nor UO_1215 (O_1215,N_8523,N_9364);
nand UO_1216 (O_1216,N_7571,N_9780);
and UO_1217 (O_1217,N_9307,N_9653);
or UO_1218 (O_1218,N_9388,N_9073);
and UO_1219 (O_1219,N_9794,N_8515);
xor UO_1220 (O_1220,N_8158,N_8147);
xnor UO_1221 (O_1221,N_7626,N_8871);
nor UO_1222 (O_1222,N_8535,N_8838);
nor UO_1223 (O_1223,N_9978,N_9458);
or UO_1224 (O_1224,N_8988,N_8932);
nand UO_1225 (O_1225,N_8139,N_7984);
nor UO_1226 (O_1226,N_9853,N_9316);
nor UO_1227 (O_1227,N_7735,N_8560);
nand UO_1228 (O_1228,N_8498,N_7883);
nand UO_1229 (O_1229,N_9288,N_9334);
and UO_1230 (O_1230,N_7633,N_7748);
nor UO_1231 (O_1231,N_8177,N_8613);
nand UO_1232 (O_1232,N_7578,N_9927);
or UO_1233 (O_1233,N_8312,N_8971);
and UO_1234 (O_1234,N_8473,N_8123);
nand UO_1235 (O_1235,N_7755,N_9287);
and UO_1236 (O_1236,N_7672,N_8852);
nand UO_1237 (O_1237,N_7612,N_9922);
nand UO_1238 (O_1238,N_7945,N_8599);
or UO_1239 (O_1239,N_8221,N_8032);
nor UO_1240 (O_1240,N_8836,N_8028);
nor UO_1241 (O_1241,N_8761,N_9088);
nor UO_1242 (O_1242,N_9970,N_8695);
xor UO_1243 (O_1243,N_8121,N_8261);
nand UO_1244 (O_1244,N_9799,N_7765);
or UO_1245 (O_1245,N_9007,N_7601);
nand UO_1246 (O_1246,N_9247,N_8882);
xnor UO_1247 (O_1247,N_9859,N_8509);
nand UO_1248 (O_1248,N_8556,N_9520);
and UO_1249 (O_1249,N_9487,N_9682);
and UO_1250 (O_1250,N_9147,N_7898);
nor UO_1251 (O_1251,N_7516,N_8444);
or UO_1252 (O_1252,N_8387,N_9507);
or UO_1253 (O_1253,N_8922,N_9224);
or UO_1254 (O_1254,N_7754,N_9547);
xnor UO_1255 (O_1255,N_8881,N_9188);
or UO_1256 (O_1256,N_8092,N_7864);
nor UO_1257 (O_1257,N_8121,N_8566);
xor UO_1258 (O_1258,N_7552,N_8444);
and UO_1259 (O_1259,N_9187,N_8191);
nor UO_1260 (O_1260,N_9926,N_9466);
or UO_1261 (O_1261,N_9745,N_7611);
or UO_1262 (O_1262,N_8852,N_8429);
or UO_1263 (O_1263,N_9590,N_9584);
and UO_1264 (O_1264,N_7931,N_8919);
xor UO_1265 (O_1265,N_8416,N_9550);
and UO_1266 (O_1266,N_9256,N_9999);
or UO_1267 (O_1267,N_9647,N_9678);
nor UO_1268 (O_1268,N_9178,N_8800);
and UO_1269 (O_1269,N_9317,N_9018);
nand UO_1270 (O_1270,N_8873,N_9659);
or UO_1271 (O_1271,N_8596,N_8681);
nand UO_1272 (O_1272,N_8007,N_9642);
nand UO_1273 (O_1273,N_8333,N_8525);
or UO_1274 (O_1274,N_8285,N_9764);
and UO_1275 (O_1275,N_9721,N_8905);
nor UO_1276 (O_1276,N_9822,N_8358);
or UO_1277 (O_1277,N_9805,N_8127);
and UO_1278 (O_1278,N_8520,N_7893);
or UO_1279 (O_1279,N_9969,N_8121);
xor UO_1280 (O_1280,N_9813,N_9351);
nand UO_1281 (O_1281,N_8210,N_9791);
and UO_1282 (O_1282,N_8333,N_8352);
and UO_1283 (O_1283,N_8387,N_9716);
and UO_1284 (O_1284,N_8239,N_7770);
or UO_1285 (O_1285,N_8476,N_8069);
and UO_1286 (O_1286,N_9280,N_7529);
xnor UO_1287 (O_1287,N_8951,N_8994);
nand UO_1288 (O_1288,N_8471,N_8264);
nand UO_1289 (O_1289,N_7988,N_9749);
and UO_1290 (O_1290,N_9316,N_7691);
and UO_1291 (O_1291,N_9063,N_8254);
xor UO_1292 (O_1292,N_9707,N_7829);
nor UO_1293 (O_1293,N_9621,N_8064);
xor UO_1294 (O_1294,N_7986,N_7603);
nor UO_1295 (O_1295,N_8884,N_8015);
or UO_1296 (O_1296,N_7778,N_7931);
xor UO_1297 (O_1297,N_9943,N_8346);
nand UO_1298 (O_1298,N_8297,N_7545);
nor UO_1299 (O_1299,N_7855,N_7831);
or UO_1300 (O_1300,N_7733,N_8400);
and UO_1301 (O_1301,N_9336,N_7641);
and UO_1302 (O_1302,N_9745,N_8286);
and UO_1303 (O_1303,N_7523,N_9106);
nand UO_1304 (O_1304,N_8629,N_7878);
xnor UO_1305 (O_1305,N_9056,N_9132);
xnor UO_1306 (O_1306,N_8270,N_8699);
nor UO_1307 (O_1307,N_9079,N_9556);
and UO_1308 (O_1308,N_9190,N_8644);
xor UO_1309 (O_1309,N_8946,N_9138);
nand UO_1310 (O_1310,N_8057,N_8443);
nand UO_1311 (O_1311,N_8796,N_9833);
xor UO_1312 (O_1312,N_9512,N_8443);
and UO_1313 (O_1313,N_7771,N_8098);
nand UO_1314 (O_1314,N_7534,N_9973);
or UO_1315 (O_1315,N_9606,N_9682);
or UO_1316 (O_1316,N_9827,N_8455);
or UO_1317 (O_1317,N_9349,N_7740);
xor UO_1318 (O_1318,N_8983,N_9033);
nand UO_1319 (O_1319,N_8227,N_9300);
and UO_1320 (O_1320,N_8143,N_7590);
xor UO_1321 (O_1321,N_9205,N_8115);
nand UO_1322 (O_1322,N_8355,N_8746);
nor UO_1323 (O_1323,N_8058,N_9316);
nor UO_1324 (O_1324,N_9764,N_7500);
xor UO_1325 (O_1325,N_9189,N_8940);
xor UO_1326 (O_1326,N_8646,N_8375);
and UO_1327 (O_1327,N_8185,N_9709);
nor UO_1328 (O_1328,N_7762,N_8855);
xor UO_1329 (O_1329,N_9962,N_7937);
and UO_1330 (O_1330,N_8935,N_7637);
nand UO_1331 (O_1331,N_7642,N_8328);
nor UO_1332 (O_1332,N_9673,N_8605);
nor UO_1333 (O_1333,N_9403,N_9670);
xor UO_1334 (O_1334,N_8952,N_7949);
and UO_1335 (O_1335,N_8685,N_8256);
nor UO_1336 (O_1336,N_8372,N_9827);
nand UO_1337 (O_1337,N_7703,N_8497);
nor UO_1338 (O_1338,N_7981,N_7615);
xor UO_1339 (O_1339,N_7817,N_8025);
nand UO_1340 (O_1340,N_7539,N_8642);
and UO_1341 (O_1341,N_7575,N_9701);
xnor UO_1342 (O_1342,N_9724,N_9774);
nand UO_1343 (O_1343,N_8711,N_8543);
xnor UO_1344 (O_1344,N_8168,N_7528);
nand UO_1345 (O_1345,N_9358,N_8137);
nor UO_1346 (O_1346,N_7924,N_9425);
xor UO_1347 (O_1347,N_7741,N_8094);
nor UO_1348 (O_1348,N_9784,N_7711);
nor UO_1349 (O_1349,N_7675,N_7557);
and UO_1350 (O_1350,N_9609,N_8770);
nor UO_1351 (O_1351,N_8199,N_9583);
nor UO_1352 (O_1352,N_9471,N_9636);
nor UO_1353 (O_1353,N_7503,N_8028);
nor UO_1354 (O_1354,N_9525,N_7739);
and UO_1355 (O_1355,N_9810,N_9125);
nand UO_1356 (O_1356,N_8617,N_9639);
and UO_1357 (O_1357,N_8571,N_7967);
xnor UO_1358 (O_1358,N_7611,N_8803);
nand UO_1359 (O_1359,N_8049,N_8731);
nand UO_1360 (O_1360,N_7972,N_9353);
and UO_1361 (O_1361,N_7598,N_9544);
or UO_1362 (O_1362,N_9276,N_7536);
and UO_1363 (O_1363,N_9078,N_8379);
nor UO_1364 (O_1364,N_8043,N_9963);
nand UO_1365 (O_1365,N_9357,N_9050);
nand UO_1366 (O_1366,N_9971,N_7909);
and UO_1367 (O_1367,N_9969,N_8380);
nor UO_1368 (O_1368,N_9113,N_9569);
and UO_1369 (O_1369,N_8486,N_9592);
nand UO_1370 (O_1370,N_8656,N_9879);
nor UO_1371 (O_1371,N_8962,N_9707);
xor UO_1372 (O_1372,N_7766,N_8888);
xnor UO_1373 (O_1373,N_9907,N_8441);
nor UO_1374 (O_1374,N_8157,N_8102);
or UO_1375 (O_1375,N_8242,N_7518);
nand UO_1376 (O_1376,N_9019,N_8805);
and UO_1377 (O_1377,N_9632,N_9142);
nand UO_1378 (O_1378,N_8205,N_8623);
and UO_1379 (O_1379,N_8569,N_7755);
nand UO_1380 (O_1380,N_9636,N_7684);
nor UO_1381 (O_1381,N_9243,N_9887);
xnor UO_1382 (O_1382,N_8864,N_9306);
nand UO_1383 (O_1383,N_9121,N_9182);
nor UO_1384 (O_1384,N_7696,N_9214);
and UO_1385 (O_1385,N_9778,N_8043);
nand UO_1386 (O_1386,N_9268,N_9539);
or UO_1387 (O_1387,N_8272,N_9323);
or UO_1388 (O_1388,N_9775,N_8356);
nand UO_1389 (O_1389,N_9253,N_9428);
or UO_1390 (O_1390,N_8756,N_9620);
nor UO_1391 (O_1391,N_8043,N_8516);
and UO_1392 (O_1392,N_9395,N_8473);
xor UO_1393 (O_1393,N_8623,N_8654);
and UO_1394 (O_1394,N_9373,N_7620);
nor UO_1395 (O_1395,N_8332,N_9575);
and UO_1396 (O_1396,N_9264,N_7764);
xnor UO_1397 (O_1397,N_9855,N_9394);
and UO_1398 (O_1398,N_7504,N_9620);
and UO_1399 (O_1399,N_9273,N_8011);
xnor UO_1400 (O_1400,N_9454,N_7826);
nand UO_1401 (O_1401,N_8137,N_9623);
and UO_1402 (O_1402,N_8230,N_9930);
xor UO_1403 (O_1403,N_8873,N_7839);
nor UO_1404 (O_1404,N_7997,N_9082);
nor UO_1405 (O_1405,N_8195,N_8263);
or UO_1406 (O_1406,N_7905,N_8333);
nor UO_1407 (O_1407,N_9433,N_9465);
or UO_1408 (O_1408,N_9758,N_9417);
or UO_1409 (O_1409,N_8323,N_9773);
or UO_1410 (O_1410,N_7901,N_8328);
nor UO_1411 (O_1411,N_9685,N_9521);
and UO_1412 (O_1412,N_8766,N_9816);
and UO_1413 (O_1413,N_7584,N_9938);
or UO_1414 (O_1414,N_8082,N_8133);
or UO_1415 (O_1415,N_8089,N_8721);
and UO_1416 (O_1416,N_8050,N_7887);
nor UO_1417 (O_1417,N_8897,N_8669);
nor UO_1418 (O_1418,N_7840,N_9491);
xnor UO_1419 (O_1419,N_8671,N_8001);
or UO_1420 (O_1420,N_9956,N_7643);
and UO_1421 (O_1421,N_8168,N_8081);
nand UO_1422 (O_1422,N_9673,N_8816);
nand UO_1423 (O_1423,N_9129,N_7703);
or UO_1424 (O_1424,N_7741,N_8571);
nor UO_1425 (O_1425,N_9485,N_8253);
or UO_1426 (O_1426,N_9559,N_8895);
xnor UO_1427 (O_1427,N_7988,N_8397);
nand UO_1428 (O_1428,N_9982,N_9435);
or UO_1429 (O_1429,N_7901,N_8806);
nor UO_1430 (O_1430,N_7651,N_8115);
or UO_1431 (O_1431,N_9403,N_7600);
and UO_1432 (O_1432,N_8503,N_8475);
xnor UO_1433 (O_1433,N_8974,N_9436);
xor UO_1434 (O_1434,N_8112,N_8784);
nand UO_1435 (O_1435,N_8229,N_7821);
and UO_1436 (O_1436,N_8544,N_7774);
xnor UO_1437 (O_1437,N_8256,N_7656);
nor UO_1438 (O_1438,N_8516,N_9820);
nand UO_1439 (O_1439,N_8824,N_9002);
nand UO_1440 (O_1440,N_8903,N_8867);
and UO_1441 (O_1441,N_8033,N_8975);
and UO_1442 (O_1442,N_9596,N_9302);
xor UO_1443 (O_1443,N_9459,N_8952);
nor UO_1444 (O_1444,N_8990,N_8648);
nor UO_1445 (O_1445,N_9188,N_7747);
or UO_1446 (O_1446,N_8937,N_9565);
nor UO_1447 (O_1447,N_8027,N_7589);
nor UO_1448 (O_1448,N_9968,N_8333);
xnor UO_1449 (O_1449,N_9199,N_8539);
xor UO_1450 (O_1450,N_8603,N_8713);
or UO_1451 (O_1451,N_9876,N_9454);
xnor UO_1452 (O_1452,N_8019,N_9578);
and UO_1453 (O_1453,N_8721,N_8591);
and UO_1454 (O_1454,N_8766,N_9801);
xor UO_1455 (O_1455,N_8185,N_8327);
or UO_1456 (O_1456,N_8016,N_9793);
xor UO_1457 (O_1457,N_9108,N_8303);
nand UO_1458 (O_1458,N_7579,N_7869);
and UO_1459 (O_1459,N_8513,N_9241);
nor UO_1460 (O_1460,N_8761,N_8397);
and UO_1461 (O_1461,N_7927,N_7676);
xor UO_1462 (O_1462,N_9274,N_7736);
xnor UO_1463 (O_1463,N_9223,N_8773);
or UO_1464 (O_1464,N_8282,N_8718);
or UO_1465 (O_1465,N_7687,N_7551);
or UO_1466 (O_1466,N_8400,N_8075);
nand UO_1467 (O_1467,N_9382,N_7624);
xor UO_1468 (O_1468,N_9159,N_8619);
xor UO_1469 (O_1469,N_9470,N_7805);
or UO_1470 (O_1470,N_8221,N_8271);
nand UO_1471 (O_1471,N_9899,N_8066);
nand UO_1472 (O_1472,N_9305,N_8406);
nor UO_1473 (O_1473,N_9583,N_7759);
xnor UO_1474 (O_1474,N_7769,N_8263);
nand UO_1475 (O_1475,N_9288,N_7589);
nor UO_1476 (O_1476,N_7957,N_7824);
or UO_1477 (O_1477,N_8751,N_7570);
and UO_1478 (O_1478,N_9328,N_7931);
or UO_1479 (O_1479,N_7972,N_8540);
nor UO_1480 (O_1480,N_7562,N_9161);
or UO_1481 (O_1481,N_8733,N_9675);
or UO_1482 (O_1482,N_8332,N_9962);
or UO_1483 (O_1483,N_8905,N_7770);
xor UO_1484 (O_1484,N_8573,N_7934);
nor UO_1485 (O_1485,N_9289,N_8055);
or UO_1486 (O_1486,N_8524,N_8538);
nand UO_1487 (O_1487,N_9753,N_7783);
xor UO_1488 (O_1488,N_7820,N_9900);
and UO_1489 (O_1489,N_8273,N_9268);
nor UO_1490 (O_1490,N_8286,N_8514);
nand UO_1491 (O_1491,N_9246,N_7929);
nor UO_1492 (O_1492,N_7794,N_8191);
or UO_1493 (O_1493,N_7653,N_8176);
and UO_1494 (O_1494,N_9780,N_9109);
nor UO_1495 (O_1495,N_8839,N_9978);
xnor UO_1496 (O_1496,N_8354,N_9113);
nand UO_1497 (O_1497,N_9234,N_7830);
nand UO_1498 (O_1498,N_7965,N_7968);
nor UO_1499 (O_1499,N_9214,N_9858);
endmodule