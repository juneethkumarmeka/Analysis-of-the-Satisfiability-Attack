module basic_500_3000_500_4_levels_1xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_91,In_281);
nand U1 (N_1,In_46,In_127);
nand U2 (N_2,In_13,In_263);
nor U3 (N_3,In_339,In_429);
nor U4 (N_4,In_311,In_114);
and U5 (N_5,In_85,In_470);
nor U6 (N_6,In_428,In_289);
or U7 (N_7,In_58,In_391);
xor U8 (N_8,In_39,In_76);
nand U9 (N_9,In_186,In_217);
and U10 (N_10,In_237,In_47);
nor U11 (N_11,In_243,In_312);
nor U12 (N_12,In_204,In_31);
and U13 (N_13,In_455,In_279);
nand U14 (N_14,In_146,In_474);
or U15 (N_15,In_215,In_187);
or U16 (N_16,In_54,In_7);
nor U17 (N_17,In_388,In_172);
nand U18 (N_18,In_229,In_275);
and U19 (N_19,In_11,In_40);
nand U20 (N_20,In_409,In_41);
nand U21 (N_21,In_469,In_177);
nand U22 (N_22,In_163,In_90);
nor U23 (N_23,In_287,In_235);
and U24 (N_24,In_483,In_396);
or U25 (N_25,In_443,In_228);
nand U26 (N_26,In_352,In_107);
and U27 (N_27,In_299,In_53);
nor U28 (N_28,In_486,In_225);
nor U29 (N_29,In_449,In_110);
or U30 (N_30,In_322,In_448);
and U31 (N_31,In_340,In_245);
xor U32 (N_32,In_176,In_387);
or U33 (N_33,In_249,In_250);
and U34 (N_34,In_231,In_456);
and U35 (N_35,In_179,In_205);
or U36 (N_36,In_355,In_270);
and U37 (N_37,In_414,In_104);
nor U38 (N_38,In_178,In_478);
nor U39 (N_39,In_402,In_431);
and U40 (N_40,In_211,In_12);
and U41 (N_41,In_441,In_410);
nand U42 (N_42,In_248,In_463);
nor U43 (N_43,In_439,In_454);
nand U44 (N_44,In_109,In_238);
and U45 (N_45,In_379,In_111);
and U46 (N_46,In_383,In_203);
and U47 (N_47,In_244,In_297);
nand U48 (N_48,In_406,In_128);
nand U49 (N_49,In_384,In_267);
nor U50 (N_50,In_349,In_133);
nor U51 (N_51,In_315,In_298);
nor U52 (N_52,In_376,In_347);
and U53 (N_53,In_28,In_135);
nor U54 (N_54,In_476,In_481);
nor U55 (N_55,In_78,In_398);
nor U56 (N_56,In_434,In_462);
nand U57 (N_57,In_75,In_356);
and U58 (N_58,In_116,In_62);
and U59 (N_59,In_381,In_389);
nand U60 (N_60,In_268,In_223);
nand U61 (N_61,In_233,In_145);
or U62 (N_62,In_288,In_149);
nor U63 (N_63,In_98,In_188);
and U64 (N_64,In_363,In_351);
nand U65 (N_65,In_296,In_258);
nor U66 (N_66,In_30,In_499);
nand U67 (N_67,In_423,In_309);
nand U68 (N_68,In_79,In_252);
nand U69 (N_69,In_304,In_152);
and U70 (N_70,In_446,In_106);
or U71 (N_71,In_416,In_120);
or U72 (N_72,In_200,In_329);
nand U73 (N_73,In_208,In_0);
nand U74 (N_74,In_21,In_447);
or U75 (N_75,In_220,In_422);
nand U76 (N_76,In_404,In_300);
nor U77 (N_77,In_256,In_490);
nand U78 (N_78,In_372,In_22);
nor U79 (N_79,In_344,In_253);
nor U80 (N_80,In_335,In_320);
nor U81 (N_81,In_35,In_317);
nor U82 (N_82,In_264,In_292);
xor U83 (N_83,In_360,In_239);
nor U84 (N_84,In_494,In_165);
or U85 (N_85,In_394,In_15);
or U86 (N_86,In_489,In_313);
nor U87 (N_87,In_419,In_147);
nor U88 (N_88,In_430,In_332);
or U89 (N_89,In_385,In_52);
nand U90 (N_90,In_411,In_8);
or U91 (N_91,In_471,In_255);
and U92 (N_92,In_453,In_173);
nand U93 (N_93,In_260,In_36);
nand U94 (N_94,In_399,In_14);
or U95 (N_95,In_166,In_161);
nor U96 (N_96,In_94,In_466);
nor U97 (N_97,In_190,In_373);
and U98 (N_98,In_89,In_459);
nand U99 (N_99,In_464,In_103);
nand U100 (N_100,In_9,In_207);
or U101 (N_101,In_336,In_440);
or U102 (N_102,In_37,In_63);
or U103 (N_103,In_353,In_43);
nand U104 (N_104,In_272,In_427);
and U105 (N_105,In_195,In_236);
nor U106 (N_106,In_6,In_38);
and U107 (N_107,In_445,In_5);
nor U108 (N_108,In_60,In_265);
or U109 (N_109,In_362,In_84);
nor U110 (N_110,In_242,In_475);
nand U111 (N_111,In_50,In_150);
or U112 (N_112,In_283,In_171);
or U113 (N_113,In_44,In_465);
nand U114 (N_114,In_66,In_302);
or U115 (N_115,In_433,In_153);
nand U116 (N_116,In_167,In_99);
nor U117 (N_117,In_139,In_1);
nand U118 (N_118,In_3,In_259);
and U119 (N_119,In_97,In_48);
and U120 (N_120,In_125,In_286);
and U121 (N_121,In_59,In_222);
nor U122 (N_122,In_407,In_393);
nor U123 (N_123,In_293,In_359);
nand U124 (N_124,In_276,In_61);
or U125 (N_125,In_226,In_174);
nand U126 (N_126,In_444,In_20);
nor U127 (N_127,In_71,In_274);
or U128 (N_128,In_131,In_34);
nor U129 (N_129,In_333,In_129);
and U130 (N_130,In_366,In_180);
and U131 (N_131,In_306,In_350);
and U132 (N_132,In_56,In_113);
nor U133 (N_133,In_155,In_325);
xor U134 (N_134,In_301,In_370);
nor U135 (N_135,In_137,In_277);
or U136 (N_136,In_123,In_375);
or U137 (N_137,In_294,In_158);
nor U138 (N_138,In_168,In_432);
nand U139 (N_139,In_421,In_266);
nor U140 (N_140,In_81,In_122);
or U141 (N_141,In_377,In_191);
nand U142 (N_142,In_197,In_487);
and U143 (N_143,In_418,In_392);
or U144 (N_144,In_307,In_33);
nand U145 (N_145,In_65,In_284);
nand U146 (N_146,In_210,In_282);
or U147 (N_147,In_119,In_68);
nand U148 (N_148,In_209,In_214);
nor U149 (N_149,In_397,In_118);
nand U150 (N_150,In_403,In_257);
nand U151 (N_151,In_357,In_87);
nand U152 (N_152,In_450,In_202);
and U153 (N_153,In_380,In_460);
nand U154 (N_154,In_479,In_124);
nand U155 (N_155,In_201,In_467);
nor U156 (N_156,In_323,In_221);
or U157 (N_157,In_148,In_251);
nor U158 (N_158,In_151,In_80);
nor U159 (N_159,In_115,In_371);
nand U160 (N_160,In_185,In_121);
nor U161 (N_161,In_194,In_159);
and U162 (N_162,In_192,In_224);
or U163 (N_163,In_425,In_227);
nand U164 (N_164,In_219,In_10);
nand U165 (N_165,In_438,In_183);
nor U166 (N_166,In_426,In_241);
or U167 (N_167,In_358,In_18);
or U168 (N_168,In_442,In_361);
nor U169 (N_169,In_319,In_25);
or U170 (N_170,In_206,In_324);
or U171 (N_171,In_346,In_310);
or U172 (N_172,In_458,In_278);
nand U173 (N_173,In_51,In_23);
nor U174 (N_174,In_101,In_285);
nand U175 (N_175,In_473,In_72);
and U176 (N_176,In_420,In_436);
nand U177 (N_177,In_364,In_74);
nor U178 (N_178,In_378,In_316);
nand U179 (N_179,In_457,In_156);
nand U180 (N_180,In_218,In_196);
nor U181 (N_181,In_343,In_412);
and U182 (N_182,In_73,In_117);
or U183 (N_183,In_184,In_138);
nand U184 (N_184,In_82,In_247);
and U185 (N_185,In_484,In_273);
nand U186 (N_186,In_141,In_77);
nand U187 (N_187,In_102,In_16);
nand U188 (N_188,In_374,In_482);
nand U189 (N_189,In_493,In_400);
nand U190 (N_190,In_395,In_485);
nor U191 (N_191,In_345,In_417);
or U192 (N_192,In_198,In_17);
or U193 (N_193,In_154,In_271);
nand U194 (N_194,In_334,In_435);
or U195 (N_195,In_86,In_480);
nand U196 (N_196,In_369,In_327);
nand U197 (N_197,In_144,In_240);
nand U198 (N_198,In_164,In_24);
nor U199 (N_199,In_130,In_95);
or U200 (N_200,In_108,In_280);
nand U201 (N_201,In_488,In_230);
and U202 (N_202,In_367,In_262);
xnor U203 (N_203,In_492,In_193);
xnor U204 (N_204,In_100,In_496);
nor U205 (N_205,In_472,In_326);
nand U206 (N_206,In_143,In_468);
nand U207 (N_207,In_27,In_338);
or U208 (N_208,In_452,In_2);
or U209 (N_209,In_386,In_497);
nand U210 (N_210,In_42,In_112);
nor U211 (N_211,In_162,In_365);
nand U212 (N_212,In_136,In_498);
nor U213 (N_213,In_330,In_390);
nor U214 (N_214,In_408,In_269);
or U215 (N_215,In_182,In_437);
nor U216 (N_216,In_199,In_477);
nor U217 (N_217,In_69,In_415);
or U218 (N_218,In_290,In_140);
nand U219 (N_219,In_134,In_83);
nand U220 (N_220,In_105,In_451);
nor U221 (N_221,In_189,In_295);
or U222 (N_222,In_382,In_405);
nand U223 (N_223,In_216,In_93);
nand U224 (N_224,In_169,In_45);
and U225 (N_225,In_337,In_261);
nor U226 (N_226,In_368,In_126);
or U227 (N_227,In_70,In_55);
and U228 (N_228,In_64,In_160);
and U229 (N_229,In_234,In_96);
or U230 (N_230,In_342,In_341);
nor U231 (N_231,In_328,In_157);
or U232 (N_232,In_303,In_321);
nor U233 (N_233,In_461,In_331);
and U234 (N_234,In_19,In_291);
xnor U235 (N_235,In_213,In_308);
nor U236 (N_236,In_175,In_413);
and U237 (N_237,In_142,In_181);
nand U238 (N_238,In_305,In_67);
nand U239 (N_239,In_88,In_92);
and U240 (N_240,In_232,In_348);
and U241 (N_241,In_57,In_354);
or U242 (N_242,In_26,In_49);
nor U243 (N_243,In_424,In_212);
nor U244 (N_244,In_132,In_32);
and U245 (N_245,In_318,In_170);
and U246 (N_246,In_4,In_401);
and U247 (N_247,In_246,In_491);
or U248 (N_248,In_495,In_314);
and U249 (N_249,In_254,In_29);
or U250 (N_250,In_303,In_371);
and U251 (N_251,In_267,In_295);
and U252 (N_252,In_432,In_214);
nand U253 (N_253,In_366,In_72);
nand U254 (N_254,In_173,In_444);
or U255 (N_255,In_329,In_452);
or U256 (N_256,In_363,In_63);
and U257 (N_257,In_363,In_26);
and U258 (N_258,In_408,In_22);
nand U259 (N_259,In_175,In_147);
nand U260 (N_260,In_447,In_253);
nor U261 (N_261,In_234,In_362);
nand U262 (N_262,In_264,In_43);
nand U263 (N_263,In_104,In_377);
nor U264 (N_264,In_289,In_287);
nor U265 (N_265,In_407,In_299);
nor U266 (N_266,In_351,In_418);
and U267 (N_267,In_172,In_88);
or U268 (N_268,In_142,In_35);
and U269 (N_269,In_34,In_243);
or U270 (N_270,In_302,In_91);
or U271 (N_271,In_459,In_359);
nand U272 (N_272,In_447,In_241);
nor U273 (N_273,In_238,In_56);
nor U274 (N_274,In_490,In_104);
and U275 (N_275,In_460,In_80);
and U276 (N_276,In_129,In_326);
nand U277 (N_277,In_465,In_77);
or U278 (N_278,In_180,In_438);
nor U279 (N_279,In_471,In_190);
nand U280 (N_280,In_485,In_150);
and U281 (N_281,In_326,In_51);
and U282 (N_282,In_364,In_414);
and U283 (N_283,In_292,In_59);
nor U284 (N_284,In_473,In_411);
nand U285 (N_285,In_499,In_24);
nand U286 (N_286,In_100,In_76);
or U287 (N_287,In_325,In_83);
and U288 (N_288,In_408,In_262);
or U289 (N_289,In_254,In_43);
nor U290 (N_290,In_172,In_430);
nand U291 (N_291,In_294,In_297);
nor U292 (N_292,In_313,In_343);
and U293 (N_293,In_458,In_238);
nor U294 (N_294,In_17,In_496);
and U295 (N_295,In_102,In_173);
nand U296 (N_296,In_421,In_380);
and U297 (N_297,In_248,In_150);
xnor U298 (N_298,In_23,In_234);
or U299 (N_299,In_458,In_409);
nand U300 (N_300,In_116,In_474);
and U301 (N_301,In_460,In_1);
and U302 (N_302,In_445,In_432);
nand U303 (N_303,In_490,In_159);
nor U304 (N_304,In_192,In_290);
nand U305 (N_305,In_425,In_81);
or U306 (N_306,In_15,In_381);
and U307 (N_307,In_196,In_60);
or U308 (N_308,In_340,In_141);
nor U309 (N_309,In_74,In_363);
and U310 (N_310,In_56,In_160);
nor U311 (N_311,In_174,In_437);
nand U312 (N_312,In_66,In_408);
or U313 (N_313,In_478,In_138);
nor U314 (N_314,In_404,In_52);
and U315 (N_315,In_431,In_2);
nand U316 (N_316,In_314,In_470);
and U317 (N_317,In_175,In_233);
or U318 (N_318,In_189,In_80);
nand U319 (N_319,In_60,In_371);
or U320 (N_320,In_312,In_84);
nor U321 (N_321,In_22,In_65);
and U322 (N_322,In_64,In_273);
nand U323 (N_323,In_142,In_269);
nor U324 (N_324,In_26,In_499);
and U325 (N_325,In_266,In_495);
or U326 (N_326,In_133,In_223);
nand U327 (N_327,In_32,In_485);
and U328 (N_328,In_112,In_415);
and U329 (N_329,In_318,In_88);
nand U330 (N_330,In_458,In_490);
nand U331 (N_331,In_337,In_42);
or U332 (N_332,In_459,In_45);
and U333 (N_333,In_173,In_349);
xor U334 (N_334,In_355,In_159);
nor U335 (N_335,In_1,In_282);
or U336 (N_336,In_359,In_114);
or U337 (N_337,In_319,In_175);
nor U338 (N_338,In_55,In_53);
nor U339 (N_339,In_16,In_315);
nand U340 (N_340,In_143,In_247);
or U341 (N_341,In_77,In_266);
or U342 (N_342,In_101,In_429);
xor U343 (N_343,In_209,In_137);
or U344 (N_344,In_342,In_81);
nand U345 (N_345,In_437,In_31);
and U346 (N_346,In_355,In_321);
nand U347 (N_347,In_385,In_136);
and U348 (N_348,In_156,In_404);
and U349 (N_349,In_6,In_94);
and U350 (N_350,In_475,In_66);
nand U351 (N_351,In_385,In_316);
nand U352 (N_352,In_204,In_3);
or U353 (N_353,In_315,In_367);
nand U354 (N_354,In_52,In_152);
or U355 (N_355,In_318,In_34);
or U356 (N_356,In_354,In_121);
and U357 (N_357,In_492,In_188);
or U358 (N_358,In_275,In_472);
or U359 (N_359,In_409,In_363);
nor U360 (N_360,In_179,In_133);
nor U361 (N_361,In_289,In_470);
nor U362 (N_362,In_457,In_227);
or U363 (N_363,In_389,In_370);
nor U364 (N_364,In_234,In_383);
or U365 (N_365,In_231,In_167);
nand U366 (N_366,In_366,In_356);
nor U367 (N_367,In_185,In_370);
or U368 (N_368,In_210,In_32);
and U369 (N_369,In_149,In_426);
nand U370 (N_370,In_499,In_485);
or U371 (N_371,In_146,In_370);
and U372 (N_372,In_337,In_242);
nand U373 (N_373,In_12,In_413);
nor U374 (N_374,In_391,In_207);
or U375 (N_375,In_22,In_407);
and U376 (N_376,In_8,In_320);
or U377 (N_377,In_451,In_60);
nor U378 (N_378,In_160,In_262);
and U379 (N_379,In_166,In_320);
or U380 (N_380,In_237,In_119);
or U381 (N_381,In_129,In_299);
nor U382 (N_382,In_349,In_378);
nor U383 (N_383,In_488,In_157);
and U384 (N_384,In_385,In_209);
nand U385 (N_385,In_130,In_215);
and U386 (N_386,In_141,In_5);
nor U387 (N_387,In_90,In_422);
nand U388 (N_388,In_328,In_449);
and U389 (N_389,In_23,In_174);
nor U390 (N_390,In_179,In_456);
or U391 (N_391,In_37,In_186);
nor U392 (N_392,In_243,In_342);
or U393 (N_393,In_49,In_243);
nor U394 (N_394,In_261,In_431);
nor U395 (N_395,In_355,In_54);
or U396 (N_396,In_281,In_419);
nor U397 (N_397,In_54,In_339);
nor U398 (N_398,In_111,In_144);
and U399 (N_399,In_428,In_283);
nand U400 (N_400,In_84,In_272);
nand U401 (N_401,In_422,In_88);
and U402 (N_402,In_470,In_78);
and U403 (N_403,In_152,In_437);
and U404 (N_404,In_168,In_192);
nand U405 (N_405,In_117,In_443);
and U406 (N_406,In_380,In_241);
or U407 (N_407,In_226,In_211);
nor U408 (N_408,In_220,In_150);
or U409 (N_409,In_491,In_225);
nor U410 (N_410,In_455,In_165);
nor U411 (N_411,In_368,In_45);
and U412 (N_412,In_387,In_395);
or U413 (N_413,In_197,In_1);
and U414 (N_414,In_276,In_313);
nand U415 (N_415,In_24,In_410);
nor U416 (N_416,In_489,In_233);
nand U417 (N_417,In_386,In_82);
and U418 (N_418,In_399,In_493);
nand U419 (N_419,In_137,In_376);
and U420 (N_420,In_165,In_438);
or U421 (N_421,In_279,In_290);
nand U422 (N_422,In_104,In_307);
nand U423 (N_423,In_455,In_86);
or U424 (N_424,In_317,In_477);
nand U425 (N_425,In_464,In_117);
and U426 (N_426,In_440,In_94);
and U427 (N_427,In_249,In_85);
and U428 (N_428,In_7,In_398);
nor U429 (N_429,In_412,In_455);
nor U430 (N_430,In_68,In_126);
or U431 (N_431,In_244,In_490);
or U432 (N_432,In_428,In_315);
and U433 (N_433,In_148,In_132);
nand U434 (N_434,In_94,In_178);
and U435 (N_435,In_12,In_177);
nand U436 (N_436,In_489,In_91);
and U437 (N_437,In_276,In_2);
and U438 (N_438,In_44,In_420);
and U439 (N_439,In_431,In_72);
nor U440 (N_440,In_117,In_415);
nand U441 (N_441,In_285,In_67);
nor U442 (N_442,In_344,In_374);
nor U443 (N_443,In_224,In_119);
or U444 (N_444,In_356,In_448);
nand U445 (N_445,In_354,In_122);
nand U446 (N_446,In_467,In_10);
and U447 (N_447,In_241,In_99);
or U448 (N_448,In_30,In_398);
or U449 (N_449,In_138,In_360);
and U450 (N_450,In_75,In_188);
xnor U451 (N_451,In_104,In_203);
or U452 (N_452,In_365,In_469);
nor U453 (N_453,In_399,In_297);
nand U454 (N_454,In_327,In_171);
nand U455 (N_455,In_437,In_433);
and U456 (N_456,In_304,In_96);
and U457 (N_457,In_187,In_66);
nand U458 (N_458,In_299,In_92);
or U459 (N_459,In_280,In_250);
and U460 (N_460,In_333,In_219);
nor U461 (N_461,In_418,In_362);
and U462 (N_462,In_402,In_258);
nand U463 (N_463,In_380,In_191);
nand U464 (N_464,In_288,In_272);
or U465 (N_465,In_371,In_297);
nand U466 (N_466,In_238,In_132);
or U467 (N_467,In_277,In_498);
nor U468 (N_468,In_422,In_473);
nand U469 (N_469,In_165,In_113);
or U470 (N_470,In_139,In_414);
nor U471 (N_471,In_49,In_240);
or U472 (N_472,In_220,In_107);
and U473 (N_473,In_495,In_36);
or U474 (N_474,In_214,In_328);
or U475 (N_475,In_494,In_155);
nand U476 (N_476,In_118,In_292);
nand U477 (N_477,In_156,In_464);
or U478 (N_478,In_56,In_415);
nand U479 (N_479,In_471,In_227);
nor U480 (N_480,In_445,In_344);
or U481 (N_481,In_323,In_380);
nor U482 (N_482,In_410,In_28);
and U483 (N_483,In_52,In_107);
or U484 (N_484,In_199,In_396);
nor U485 (N_485,In_473,In_23);
nor U486 (N_486,In_53,In_353);
nor U487 (N_487,In_407,In_330);
or U488 (N_488,In_410,In_361);
nor U489 (N_489,In_461,In_160);
or U490 (N_490,In_346,In_147);
or U491 (N_491,In_418,In_97);
nor U492 (N_492,In_203,In_498);
and U493 (N_493,In_463,In_82);
and U494 (N_494,In_290,In_153);
or U495 (N_495,In_22,In_260);
nor U496 (N_496,In_225,In_344);
and U497 (N_497,In_175,In_367);
nand U498 (N_498,In_86,In_402);
or U499 (N_499,In_187,In_475);
nand U500 (N_500,In_45,In_188);
nor U501 (N_501,In_181,In_407);
nand U502 (N_502,In_42,In_87);
or U503 (N_503,In_108,In_378);
and U504 (N_504,In_424,In_2);
and U505 (N_505,In_386,In_456);
nor U506 (N_506,In_391,In_285);
xor U507 (N_507,In_206,In_294);
or U508 (N_508,In_360,In_325);
and U509 (N_509,In_85,In_418);
nor U510 (N_510,In_188,In_220);
nand U511 (N_511,In_84,In_183);
or U512 (N_512,In_52,In_440);
xor U513 (N_513,In_445,In_349);
and U514 (N_514,In_381,In_43);
nand U515 (N_515,In_42,In_309);
or U516 (N_516,In_432,In_294);
nor U517 (N_517,In_212,In_309);
nor U518 (N_518,In_19,In_465);
nor U519 (N_519,In_280,In_290);
or U520 (N_520,In_51,In_210);
nand U521 (N_521,In_337,In_349);
nand U522 (N_522,In_92,In_14);
and U523 (N_523,In_295,In_137);
or U524 (N_524,In_457,In_278);
nor U525 (N_525,In_189,In_101);
or U526 (N_526,In_303,In_151);
nand U527 (N_527,In_188,In_204);
or U528 (N_528,In_257,In_489);
and U529 (N_529,In_315,In_453);
or U530 (N_530,In_204,In_207);
nor U531 (N_531,In_131,In_270);
nand U532 (N_532,In_204,In_88);
nor U533 (N_533,In_441,In_4);
and U534 (N_534,In_438,In_115);
nand U535 (N_535,In_274,In_212);
or U536 (N_536,In_470,In_184);
or U537 (N_537,In_133,In_74);
nand U538 (N_538,In_410,In_178);
or U539 (N_539,In_453,In_3);
nor U540 (N_540,In_339,In_64);
nor U541 (N_541,In_150,In_166);
nor U542 (N_542,In_335,In_240);
nor U543 (N_543,In_393,In_229);
nand U544 (N_544,In_369,In_392);
nand U545 (N_545,In_325,In_418);
or U546 (N_546,In_240,In_8);
or U547 (N_547,In_354,In_213);
or U548 (N_548,In_7,In_208);
and U549 (N_549,In_145,In_376);
and U550 (N_550,In_494,In_255);
nand U551 (N_551,In_308,In_311);
and U552 (N_552,In_53,In_187);
nor U553 (N_553,In_478,In_224);
or U554 (N_554,In_448,In_272);
or U555 (N_555,In_466,In_74);
xor U556 (N_556,In_222,In_269);
and U557 (N_557,In_419,In_12);
and U558 (N_558,In_475,In_80);
nand U559 (N_559,In_190,In_321);
nor U560 (N_560,In_429,In_178);
nor U561 (N_561,In_32,In_398);
and U562 (N_562,In_431,In_194);
or U563 (N_563,In_245,In_391);
and U564 (N_564,In_141,In_293);
and U565 (N_565,In_258,In_153);
and U566 (N_566,In_38,In_114);
and U567 (N_567,In_156,In_302);
and U568 (N_568,In_462,In_436);
nor U569 (N_569,In_111,In_249);
or U570 (N_570,In_26,In_32);
or U571 (N_571,In_358,In_465);
nand U572 (N_572,In_395,In_92);
and U573 (N_573,In_324,In_298);
and U574 (N_574,In_412,In_269);
or U575 (N_575,In_352,In_195);
and U576 (N_576,In_434,In_179);
nand U577 (N_577,In_263,In_98);
and U578 (N_578,In_227,In_472);
or U579 (N_579,In_118,In_359);
nand U580 (N_580,In_304,In_63);
nor U581 (N_581,In_158,In_234);
or U582 (N_582,In_429,In_193);
or U583 (N_583,In_36,In_295);
and U584 (N_584,In_464,In_345);
nor U585 (N_585,In_231,In_182);
or U586 (N_586,In_204,In_170);
and U587 (N_587,In_77,In_388);
and U588 (N_588,In_271,In_31);
or U589 (N_589,In_370,In_226);
and U590 (N_590,In_241,In_353);
or U591 (N_591,In_334,In_409);
and U592 (N_592,In_392,In_269);
nor U593 (N_593,In_132,In_197);
and U594 (N_594,In_139,In_439);
nand U595 (N_595,In_45,In_351);
nor U596 (N_596,In_17,In_211);
or U597 (N_597,In_15,In_150);
nand U598 (N_598,In_193,In_89);
or U599 (N_599,In_225,In_106);
nor U600 (N_600,In_386,In_293);
nand U601 (N_601,In_461,In_434);
and U602 (N_602,In_425,In_61);
nand U603 (N_603,In_385,In_293);
or U604 (N_604,In_183,In_107);
nand U605 (N_605,In_192,In_169);
or U606 (N_606,In_304,In_256);
or U607 (N_607,In_299,In_150);
or U608 (N_608,In_318,In_338);
nand U609 (N_609,In_110,In_407);
nor U610 (N_610,In_223,In_356);
nor U611 (N_611,In_337,In_227);
nor U612 (N_612,In_465,In_40);
nand U613 (N_613,In_20,In_8);
nand U614 (N_614,In_111,In_108);
nor U615 (N_615,In_17,In_70);
or U616 (N_616,In_110,In_2);
or U617 (N_617,In_386,In_349);
nand U618 (N_618,In_208,In_73);
nand U619 (N_619,In_193,In_329);
nor U620 (N_620,In_276,In_240);
and U621 (N_621,In_192,In_359);
or U622 (N_622,In_9,In_62);
and U623 (N_623,In_481,In_174);
nand U624 (N_624,In_68,In_44);
or U625 (N_625,In_384,In_160);
or U626 (N_626,In_96,In_484);
nor U627 (N_627,In_77,In_329);
nand U628 (N_628,In_18,In_69);
or U629 (N_629,In_262,In_157);
or U630 (N_630,In_300,In_46);
nand U631 (N_631,In_351,In_328);
nand U632 (N_632,In_296,In_208);
or U633 (N_633,In_375,In_134);
xnor U634 (N_634,In_134,In_187);
nor U635 (N_635,In_333,In_392);
nand U636 (N_636,In_474,In_405);
and U637 (N_637,In_132,In_144);
and U638 (N_638,In_266,In_208);
and U639 (N_639,In_59,In_296);
or U640 (N_640,In_26,In_192);
nand U641 (N_641,In_456,In_108);
nor U642 (N_642,In_297,In_300);
or U643 (N_643,In_363,In_249);
and U644 (N_644,In_391,In_46);
nor U645 (N_645,In_388,In_474);
and U646 (N_646,In_414,In_85);
and U647 (N_647,In_72,In_493);
or U648 (N_648,In_404,In_13);
and U649 (N_649,In_2,In_86);
nor U650 (N_650,In_1,In_278);
nand U651 (N_651,In_281,In_134);
or U652 (N_652,In_289,In_45);
and U653 (N_653,In_447,In_246);
nor U654 (N_654,In_343,In_432);
nand U655 (N_655,In_163,In_311);
nor U656 (N_656,In_43,In_482);
and U657 (N_657,In_226,In_175);
and U658 (N_658,In_364,In_434);
and U659 (N_659,In_362,In_247);
and U660 (N_660,In_57,In_421);
nor U661 (N_661,In_101,In_0);
or U662 (N_662,In_357,In_39);
and U663 (N_663,In_364,In_371);
nand U664 (N_664,In_282,In_488);
nand U665 (N_665,In_382,In_297);
or U666 (N_666,In_375,In_393);
and U667 (N_667,In_378,In_84);
nor U668 (N_668,In_178,In_236);
nor U669 (N_669,In_156,In_284);
nor U670 (N_670,In_304,In_42);
and U671 (N_671,In_338,In_147);
and U672 (N_672,In_329,In_109);
nand U673 (N_673,In_0,In_435);
nand U674 (N_674,In_476,In_478);
or U675 (N_675,In_299,In_459);
nor U676 (N_676,In_483,In_41);
nor U677 (N_677,In_247,In_24);
or U678 (N_678,In_227,In_197);
and U679 (N_679,In_446,In_179);
and U680 (N_680,In_356,In_162);
and U681 (N_681,In_226,In_42);
nor U682 (N_682,In_29,In_179);
nor U683 (N_683,In_0,In_481);
nor U684 (N_684,In_248,In_239);
nand U685 (N_685,In_257,In_416);
and U686 (N_686,In_96,In_308);
and U687 (N_687,In_442,In_383);
and U688 (N_688,In_304,In_40);
nor U689 (N_689,In_69,In_355);
nand U690 (N_690,In_471,In_361);
or U691 (N_691,In_496,In_300);
or U692 (N_692,In_102,In_354);
or U693 (N_693,In_353,In_36);
nand U694 (N_694,In_86,In_416);
or U695 (N_695,In_130,In_78);
nor U696 (N_696,In_24,In_194);
or U697 (N_697,In_481,In_444);
nand U698 (N_698,In_264,In_309);
or U699 (N_699,In_380,In_496);
nand U700 (N_700,In_112,In_74);
nor U701 (N_701,In_52,In_10);
nor U702 (N_702,In_19,In_96);
and U703 (N_703,In_121,In_462);
or U704 (N_704,In_76,In_219);
or U705 (N_705,In_80,In_8);
or U706 (N_706,In_97,In_184);
nor U707 (N_707,In_122,In_469);
or U708 (N_708,In_474,In_79);
nor U709 (N_709,In_363,In_224);
or U710 (N_710,In_381,In_213);
nor U711 (N_711,In_456,In_147);
nor U712 (N_712,In_359,In_9);
xnor U713 (N_713,In_0,In_64);
xnor U714 (N_714,In_40,In_485);
and U715 (N_715,In_432,In_472);
xor U716 (N_716,In_118,In_456);
nor U717 (N_717,In_309,In_47);
nand U718 (N_718,In_208,In_38);
or U719 (N_719,In_62,In_56);
or U720 (N_720,In_338,In_371);
nor U721 (N_721,In_56,In_365);
nand U722 (N_722,In_165,In_140);
xnor U723 (N_723,In_293,In_250);
nor U724 (N_724,In_250,In_146);
or U725 (N_725,In_217,In_3);
nor U726 (N_726,In_185,In_14);
nand U727 (N_727,In_319,In_244);
and U728 (N_728,In_287,In_168);
nor U729 (N_729,In_497,In_120);
or U730 (N_730,In_400,In_175);
and U731 (N_731,In_483,In_472);
or U732 (N_732,In_0,In_199);
and U733 (N_733,In_185,In_451);
nand U734 (N_734,In_434,In_320);
nand U735 (N_735,In_487,In_134);
nor U736 (N_736,In_269,In_51);
nor U737 (N_737,In_174,In_258);
nor U738 (N_738,In_429,In_161);
and U739 (N_739,In_33,In_294);
and U740 (N_740,In_31,In_7);
nor U741 (N_741,In_37,In_383);
and U742 (N_742,In_47,In_423);
or U743 (N_743,In_259,In_201);
or U744 (N_744,In_327,In_212);
and U745 (N_745,In_118,In_296);
and U746 (N_746,In_392,In_275);
or U747 (N_747,In_489,In_428);
nand U748 (N_748,In_281,In_300);
nand U749 (N_749,In_30,In_350);
or U750 (N_750,N_322,N_593);
nor U751 (N_751,N_583,N_329);
or U752 (N_752,N_594,N_668);
nand U753 (N_753,N_584,N_542);
nor U754 (N_754,N_655,N_224);
nor U755 (N_755,N_433,N_264);
nor U756 (N_756,N_174,N_181);
nand U757 (N_757,N_740,N_696);
or U758 (N_758,N_465,N_480);
or U759 (N_759,N_199,N_641);
nor U760 (N_760,N_253,N_614);
or U761 (N_761,N_451,N_527);
nand U762 (N_762,N_581,N_724);
xnor U763 (N_763,N_151,N_164);
nand U764 (N_764,N_82,N_96);
nand U765 (N_765,N_715,N_679);
nor U766 (N_766,N_11,N_667);
and U767 (N_767,N_179,N_472);
and U768 (N_768,N_684,N_633);
nor U769 (N_769,N_540,N_454);
and U770 (N_770,N_222,N_304);
nor U771 (N_771,N_44,N_694);
nor U772 (N_772,N_336,N_533);
nor U773 (N_773,N_499,N_689);
and U774 (N_774,N_207,N_28);
or U775 (N_775,N_463,N_648);
or U776 (N_776,N_241,N_640);
nor U777 (N_777,N_685,N_229);
nand U778 (N_778,N_61,N_574);
or U779 (N_779,N_323,N_80);
nand U780 (N_780,N_344,N_482);
or U781 (N_781,N_575,N_682);
or U782 (N_782,N_391,N_255);
or U783 (N_783,N_320,N_49);
nand U784 (N_784,N_675,N_595);
nand U785 (N_785,N_328,N_136);
nand U786 (N_786,N_494,N_307);
nor U787 (N_787,N_627,N_268);
and U788 (N_788,N_739,N_182);
or U789 (N_789,N_205,N_147);
or U790 (N_790,N_672,N_467);
nor U791 (N_791,N_298,N_321);
or U792 (N_792,N_156,N_259);
nand U793 (N_793,N_230,N_635);
nor U794 (N_794,N_416,N_319);
nor U795 (N_795,N_507,N_741);
nor U796 (N_796,N_159,N_619);
nor U797 (N_797,N_726,N_204);
nor U798 (N_798,N_611,N_92);
nand U799 (N_799,N_330,N_16);
nand U800 (N_800,N_504,N_585);
and U801 (N_801,N_210,N_364);
or U802 (N_802,N_237,N_101);
and U803 (N_803,N_70,N_380);
or U804 (N_804,N_162,N_200);
nand U805 (N_805,N_34,N_352);
nand U806 (N_806,N_612,N_500);
nor U807 (N_807,N_282,N_40);
nand U808 (N_808,N_447,N_299);
nand U809 (N_809,N_456,N_664);
nand U810 (N_810,N_77,N_291);
nand U811 (N_811,N_64,N_128);
or U812 (N_812,N_48,N_26);
or U813 (N_813,N_252,N_520);
or U814 (N_814,N_471,N_38);
and U815 (N_815,N_130,N_506);
nand U816 (N_816,N_24,N_603);
nand U817 (N_817,N_529,N_290);
nand U818 (N_818,N_530,N_260);
nand U819 (N_819,N_123,N_634);
and U820 (N_820,N_599,N_459);
nor U821 (N_821,N_676,N_42);
or U822 (N_822,N_343,N_281);
or U823 (N_823,N_98,N_478);
nand U824 (N_824,N_414,N_541);
nor U825 (N_825,N_663,N_335);
nand U826 (N_826,N_466,N_671);
or U827 (N_827,N_324,N_188);
nand U828 (N_828,N_526,N_395);
nand U829 (N_829,N_242,N_607);
and U830 (N_830,N_382,N_310);
and U831 (N_831,N_216,N_749);
and U832 (N_832,N_318,N_432);
nand U833 (N_833,N_625,N_7);
and U834 (N_834,N_286,N_536);
nor U835 (N_835,N_458,N_251);
nand U836 (N_836,N_347,N_680);
or U837 (N_837,N_449,N_355);
and U838 (N_838,N_0,N_103);
nand U839 (N_839,N_415,N_538);
or U840 (N_840,N_484,N_651);
nor U841 (N_841,N_231,N_398);
or U842 (N_842,N_201,N_440);
or U843 (N_843,N_544,N_687);
nor U844 (N_844,N_58,N_600);
nor U845 (N_845,N_591,N_125);
and U846 (N_846,N_621,N_656);
nand U847 (N_847,N_191,N_562);
and U848 (N_848,N_501,N_121);
or U849 (N_849,N_345,N_617);
nor U850 (N_850,N_327,N_309);
nand U851 (N_851,N_144,N_618);
or U852 (N_852,N_218,N_273);
or U853 (N_853,N_637,N_378);
nor U854 (N_854,N_220,N_427);
nand U855 (N_855,N_550,N_226);
nor U856 (N_856,N_570,N_735);
and U857 (N_857,N_187,N_175);
or U858 (N_858,N_576,N_69);
nor U859 (N_859,N_517,N_403);
and U860 (N_860,N_742,N_236);
or U861 (N_861,N_620,N_557);
or U862 (N_862,N_301,N_5);
and U863 (N_863,N_111,N_35);
nand U864 (N_864,N_359,N_71);
nor U865 (N_865,N_485,N_346);
and U866 (N_866,N_443,N_525);
xor U867 (N_867,N_196,N_184);
or U868 (N_868,N_261,N_721);
and U869 (N_869,N_45,N_654);
or U870 (N_870,N_582,N_592);
or U871 (N_871,N_561,N_502);
or U872 (N_872,N_413,N_624);
nand U873 (N_873,N_228,N_59);
nor U874 (N_874,N_25,N_510);
nor U875 (N_875,N_183,N_217);
nor U876 (N_876,N_375,N_243);
and U877 (N_877,N_356,N_89);
or U878 (N_878,N_528,N_531);
and U879 (N_879,N_445,N_461);
or U880 (N_880,N_138,N_41);
nand U881 (N_881,N_386,N_155);
or U882 (N_882,N_744,N_95);
nand U883 (N_883,N_513,N_73);
nand U884 (N_884,N_3,N_703);
nand U885 (N_885,N_509,N_590);
and U886 (N_886,N_537,N_404);
nor U887 (N_887,N_94,N_438);
and U888 (N_888,N_350,N_234);
or U889 (N_889,N_137,N_43);
nand U890 (N_890,N_332,N_565);
nor U891 (N_891,N_6,N_662);
or U892 (N_892,N_300,N_367);
or U893 (N_893,N_645,N_748);
and U894 (N_894,N_709,N_453);
nand U895 (N_895,N_686,N_288);
and U896 (N_896,N_280,N_305);
nor U897 (N_897,N_396,N_102);
nor U898 (N_898,N_149,N_161);
nand U899 (N_899,N_247,N_314);
or U900 (N_900,N_189,N_642);
nor U901 (N_901,N_609,N_361);
or U902 (N_902,N_365,N_420);
or U903 (N_903,N_15,N_468);
and U904 (N_904,N_503,N_475);
and U905 (N_905,N_418,N_295);
nand U906 (N_906,N_691,N_362);
nor U907 (N_907,N_14,N_407);
nand U908 (N_908,N_248,N_57);
or U909 (N_909,N_400,N_37);
or U910 (N_910,N_177,N_695);
and U911 (N_911,N_489,N_81);
or U912 (N_912,N_732,N_46);
and U913 (N_913,N_688,N_197);
nand U914 (N_914,N_498,N_644);
or U915 (N_915,N_434,N_613);
nand U916 (N_916,N_341,N_276);
xnor U917 (N_917,N_4,N_518);
nand U918 (N_918,N_457,N_342);
nor U919 (N_919,N_545,N_674);
or U920 (N_920,N_158,N_532);
nor U921 (N_921,N_622,N_496);
and U922 (N_922,N_254,N_65);
nand U923 (N_923,N_154,N_631);
and U924 (N_924,N_589,N_139);
nor U925 (N_925,N_269,N_579);
or U926 (N_926,N_711,N_134);
nand U927 (N_927,N_474,N_441);
nand U928 (N_928,N_317,N_293);
or U929 (N_929,N_12,N_444);
nor U930 (N_930,N_133,N_745);
nand U931 (N_931,N_374,N_165);
or U932 (N_932,N_135,N_90);
nand U933 (N_933,N_402,N_713);
and U934 (N_934,N_554,N_258);
or U935 (N_935,N_580,N_512);
or U936 (N_936,N_727,N_649);
and U937 (N_937,N_166,N_308);
xor U938 (N_938,N_129,N_50);
nand U939 (N_939,N_194,N_481);
or U940 (N_940,N_521,N_412);
and U941 (N_941,N_112,N_53);
or U942 (N_942,N_702,N_22);
or U943 (N_943,N_326,N_516);
or U944 (N_944,N_647,N_140);
or U945 (N_945,N_373,N_431);
or U946 (N_946,N_477,N_747);
and U947 (N_947,N_708,N_54);
or U948 (N_948,N_523,N_608);
nor U949 (N_949,N_132,N_249);
nor U950 (N_950,N_665,N_553);
and U951 (N_951,N_473,N_256);
nor U952 (N_952,N_208,N_240);
or U953 (N_953,N_569,N_389);
or U954 (N_954,N_172,N_435);
or U955 (N_955,N_30,N_723);
and U956 (N_956,N_535,N_211);
or U957 (N_957,N_601,N_598);
nor U958 (N_958,N_491,N_572);
nand U959 (N_959,N_85,N_377);
and U960 (N_960,N_490,N_60);
and U961 (N_961,N_623,N_267);
and U962 (N_962,N_296,N_738);
or U963 (N_963,N_388,N_351);
and U964 (N_964,N_119,N_354);
nand U965 (N_965,N_366,N_549);
nand U966 (N_966,N_636,N_392);
and U967 (N_967,N_17,N_659);
nand U968 (N_968,N_99,N_720);
nor U969 (N_969,N_455,N_728);
or U970 (N_970,N_712,N_100);
nand U971 (N_971,N_105,N_209);
nand U972 (N_972,N_730,N_657);
and U973 (N_973,N_331,N_272);
nor U974 (N_974,N_180,N_107);
nor U975 (N_975,N_47,N_719);
or U976 (N_976,N_171,N_312);
nand U977 (N_977,N_571,N_379);
nand U978 (N_978,N_376,N_79);
nor U979 (N_979,N_556,N_394);
nand U980 (N_980,N_120,N_63);
nor U981 (N_981,N_587,N_145);
nand U982 (N_982,N_437,N_313);
or U983 (N_983,N_9,N_408);
nor U984 (N_984,N_195,N_646);
nor U985 (N_985,N_371,N_124);
nor U986 (N_986,N_479,N_372);
and U987 (N_987,N_238,N_212);
or U988 (N_988,N_84,N_652);
nand U989 (N_989,N_153,N_469);
nand U990 (N_990,N_419,N_339);
nor U991 (N_991,N_606,N_737);
nand U992 (N_992,N_68,N_401);
and U993 (N_993,N_148,N_353);
and U994 (N_994,N_409,N_495);
or U995 (N_995,N_639,N_425);
or U996 (N_996,N_493,N_424);
nand U997 (N_997,N_460,N_152);
and U998 (N_998,N_660,N_340);
or U999 (N_999,N_397,N_223);
nor U1000 (N_1000,N_524,N_337);
nand U1001 (N_1001,N_275,N_422);
nor U1002 (N_1002,N_446,N_734);
or U1003 (N_1003,N_170,N_487);
nor U1004 (N_1004,N_733,N_439);
and U1005 (N_1005,N_505,N_245);
or U1006 (N_1006,N_710,N_650);
nand U1007 (N_1007,N_97,N_262);
nor U1008 (N_1008,N_227,N_178);
or U1009 (N_1009,N_514,N_126);
nand U1010 (N_1010,N_198,N_629);
nand U1011 (N_1011,N_705,N_190);
and U1012 (N_1012,N_368,N_157);
nor U1013 (N_1013,N_108,N_29);
nor U1014 (N_1014,N_219,N_552);
nand U1015 (N_1015,N_39,N_743);
or U1016 (N_1016,N_610,N_605);
or U1017 (N_1017,N_274,N_143);
nand U1018 (N_1018,N_76,N_193);
or U1019 (N_1019,N_638,N_677);
and U1020 (N_1020,N_548,N_736);
or U1021 (N_1021,N_192,N_692);
or U1022 (N_1022,N_32,N_597);
or U1023 (N_1023,N_430,N_289);
or U1024 (N_1024,N_673,N_716);
nor U1025 (N_1025,N_360,N_405);
nand U1026 (N_1026,N_348,N_244);
nor U1027 (N_1027,N_52,N_106);
nand U1028 (N_1028,N_141,N_543);
nor U1029 (N_1029,N_383,N_511);
nor U1030 (N_1030,N_349,N_225);
nor U1031 (N_1031,N_169,N_232);
nor U1032 (N_1032,N_86,N_567);
nand U1033 (N_1033,N_150,N_257);
or U1034 (N_1034,N_653,N_566);
or U1035 (N_1035,N_508,N_577);
nor U1036 (N_1036,N_555,N_303);
or U1037 (N_1037,N_701,N_338);
nand U1038 (N_1038,N_486,N_729);
or U1039 (N_1039,N_693,N_110);
xor U1040 (N_1040,N_573,N_423);
or U1041 (N_1041,N_55,N_370);
nor U1042 (N_1042,N_588,N_604);
nand U1043 (N_1043,N_700,N_292);
nand U1044 (N_1044,N_669,N_203);
or U1045 (N_1045,N_746,N_142);
and U1046 (N_1046,N_357,N_221);
or U1047 (N_1047,N_714,N_421);
or U1048 (N_1048,N_88,N_315);
nand U1049 (N_1049,N_411,N_160);
or U1050 (N_1050,N_287,N_596);
nand U1051 (N_1051,N_83,N_534);
nand U1052 (N_1052,N_306,N_19);
or U1053 (N_1053,N_515,N_442);
nor U1054 (N_1054,N_202,N_699);
and U1055 (N_1055,N_114,N_628);
nor U1056 (N_1056,N_185,N_213);
nor U1057 (N_1057,N_20,N_75);
or U1058 (N_1058,N_186,N_704);
nand U1059 (N_1059,N_426,N_78);
nand U1060 (N_1060,N_390,N_13);
nor U1061 (N_1061,N_559,N_118);
or U1062 (N_1062,N_146,N_586);
nor U1063 (N_1063,N_233,N_564);
nor U1064 (N_1064,N_492,N_235);
or U1065 (N_1065,N_632,N_681);
and U1066 (N_1066,N_263,N_464);
or U1067 (N_1067,N_18,N_115);
nor U1068 (N_1068,N_363,N_277);
nand U1069 (N_1069,N_74,N_578);
nand U1070 (N_1070,N_283,N_91);
nand U1071 (N_1071,N_393,N_476);
nor U1072 (N_1072,N_302,N_630);
or U1073 (N_1073,N_163,N_36);
nor U1074 (N_1074,N_33,N_72);
and U1075 (N_1075,N_278,N_131);
or U1076 (N_1076,N_399,N_568);
nor U1077 (N_1077,N_462,N_488);
nand U1078 (N_1078,N_558,N_683);
and U1079 (N_1079,N_250,N_547);
nor U1080 (N_1080,N_717,N_27);
or U1081 (N_1081,N_725,N_10);
and U1082 (N_1082,N_690,N_246);
nand U1083 (N_1083,N_678,N_104);
nand U1084 (N_1084,N_560,N_661);
nand U1085 (N_1085,N_718,N_522);
nor U1086 (N_1086,N_2,N_436);
or U1087 (N_1087,N_551,N_271);
nor U1088 (N_1088,N_429,N_270);
nand U1089 (N_1089,N_722,N_381);
nor U1090 (N_1090,N_8,N_23);
or U1091 (N_1091,N_116,N_670);
nor U1092 (N_1092,N_616,N_239);
and U1093 (N_1093,N_539,N_67);
nand U1094 (N_1094,N_21,N_168);
nand U1095 (N_1095,N_31,N_707);
xor U1096 (N_1096,N_284,N_215);
nor U1097 (N_1097,N_167,N_731);
nand U1098 (N_1098,N_87,N_93);
or U1099 (N_1099,N_697,N_56);
nor U1100 (N_1100,N_265,N_66);
or U1101 (N_1101,N_297,N_698);
nor U1102 (N_1102,N_410,N_706);
or U1103 (N_1103,N_626,N_519);
and U1104 (N_1104,N_214,N_483);
or U1105 (N_1105,N_369,N_109);
nand U1106 (N_1106,N_384,N_385);
nand U1107 (N_1107,N_448,N_122);
and U1108 (N_1108,N_285,N_266);
or U1109 (N_1109,N_417,N_602);
or U1110 (N_1110,N_563,N_316);
nor U1111 (N_1111,N_127,N_406);
or U1112 (N_1112,N_117,N_666);
and U1113 (N_1113,N_546,N_311);
nand U1114 (N_1114,N_643,N_173);
nor U1115 (N_1115,N_325,N_387);
or U1116 (N_1116,N_113,N_62);
nor U1117 (N_1117,N_1,N_615);
nand U1118 (N_1118,N_452,N_279);
nand U1119 (N_1119,N_206,N_428);
nor U1120 (N_1120,N_294,N_358);
nand U1121 (N_1121,N_450,N_176);
nor U1122 (N_1122,N_658,N_333);
nand U1123 (N_1123,N_51,N_497);
or U1124 (N_1124,N_334,N_470);
or U1125 (N_1125,N_49,N_638);
or U1126 (N_1126,N_597,N_575);
nand U1127 (N_1127,N_239,N_487);
nand U1128 (N_1128,N_538,N_97);
and U1129 (N_1129,N_592,N_662);
and U1130 (N_1130,N_224,N_313);
nor U1131 (N_1131,N_41,N_107);
and U1132 (N_1132,N_419,N_268);
nand U1133 (N_1133,N_93,N_123);
nor U1134 (N_1134,N_222,N_151);
or U1135 (N_1135,N_247,N_489);
or U1136 (N_1136,N_28,N_450);
nand U1137 (N_1137,N_119,N_288);
and U1138 (N_1138,N_349,N_395);
and U1139 (N_1139,N_413,N_308);
nor U1140 (N_1140,N_59,N_293);
or U1141 (N_1141,N_714,N_508);
nor U1142 (N_1142,N_569,N_638);
nor U1143 (N_1143,N_63,N_54);
nand U1144 (N_1144,N_590,N_194);
and U1145 (N_1145,N_329,N_540);
or U1146 (N_1146,N_237,N_624);
or U1147 (N_1147,N_558,N_679);
nand U1148 (N_1148,N_488,N_681);
nor U1149 (N_1149,N_132,N_361);
nand U1150 (N_1150,N_116,N_599);
nand U1151 (N_1151,N_79,N_27);
or U1152 (N_1152,N_165,N_703);
nand U1153 (N_1153,N_400,N_167);
xnor U1154 (N_1154,N_82,N_108);
nand U1155 (N_1155,N_92,N_105);
nand U1156 (N_1156,N_310,N_349);
or U1157 (N_1157,N_565,N_278);
nor U1158 (N_1158,N_18,N_748);
nand U1159 (N_1159,N_631,N_81);
and U1160 (N_1160,N_6,N_109);
or U1161 (N_1161,N_24,N_346);
or U1162 (N_1162,N_296,N_55);
nand U1163 (N_1163,N_409,N_374);
nor U1164 (N_1164,N_23,N_662);
or U1165 (N_1165,N_59,N_559);
nand U1166 (N_1166,N_41,N_425);
and U1167 (N_1167,N_559,N_503);
nor U1168 (N_1168,N_98,N_647);
and U1169 (N_1169,N_716,N_611);
or U1170 (N_1170,N_493,N_255);
and U1171 (N_1171,N_316,N_354);
and U1172 (N_1172,N_230,N_358);
and U1173 (N_1173,N_675,N_24);
nor U1174 (N_1174,N_595,N_288);
nand U1175 (N_1175,N_88,N_284);
and U1176 (N_1176,N_505,N_206);
or U1177 (N_1177,N_212,N_339);
and U1178 (N_1178,N_36,N_515);
nor U1179 (N_1179,N_638,N_303);
nor U1180 (N_1180,N_422,N_727);
and U1181 (N_1181,N_528,N_64);
or U1182 (N_1182,N_594,N_248);
nor U1183 (N_1183,N_415,N_2);
nand U1184 (N_1184,N_260,N_362);
nor U1185 (N_1185,N_469,N_322);
nor U1186 (N_1186,N_346,N_144);
nand U1187 (N_1187,N_744,N_357);
nand U1188 (N_1188,N_204,N_75);
and U1189 (N_1189,N_594,N_717);
and U1190 (N_1190,N_620,N_482);
nor U1191 (N_1191,N_602,N_3);
nand U1192 (N_1192,N_415,N_333);
or U1193 (N_1193,N_107,N_491);
or U1194 (N_1194,N_280,N_3);
or U1195 (N_1195,N_5,N_528);
and U1196 (N_1196,N_547,N_371);
nand U1197 (N_1197,N_677,N_608);
and U1198 (N_1198,N_400,N_383);
or U1199 (N_1199,N_639,N_322);
or U1200 (N_1200,N_10,N_366);
and U1201 (N_1201,N_110,N_6);
nor U1202 (N_1202,N_704,N_693);
nand U1203 (N_1203,N_124,N_271);
nand U1204 (N_1204,N_94,N_133);
nor U1205 (N_1205,N_332,N_42);
and U1206 (N_1206,N_104,N_186);
nand U1207 (N_1207,N_686,N_627);
nand U1208 (N_1208,N_68,N_666);
or U1209 (N_1209,N_142,N_387);
nand U1210 (N_1210,N_266,N_565);
or U1211 (N_1211,N_200,N_164);
nand U1212 (N_1212,N_541,N_393);
and U1213 (N_1213,N_117,N_408);
nor U1214 (N_1214,N_60,N_240);
nand U1215 (N_1215,N_680,N_666);
nor U1216 (N_1216,N_322,N_258);
and U1217 (N_1217,N_709,N_16);
xor U1218 (N_1218,N_506,N_557);
or U1219 (N_1219,N_494,N_643);
nor U1220 (N_1220,N_122,N_328);
xnor U1221 (N_1221,N_638,N_589);
or U1222 (N_1222,N_404,N_678);
or U1223 (N_1223,N_299,N_81);
nand U1224 (N_1224,N_279,N_707);
nand U1225 (N_1225,N_198,N_438);
or U1226 (N_1226,N_221,N_230);
nand U1227 (N_1227,N_111,N_469);
and U1228 (N_1228,N_432,N_29);
nand U1229 (N_1229,N_459,N_75);
and U1230 (N_1230,N_702,N_72);
and U1231 (N_1231,N_438,N_473);
or U1232 (N_1232,N_732,N_392);
and U1233 (N_1233,N_623,N_496);
nand U1234 (N_1234,N_233,N_239);
or U1235 (N_1235,N_633,N_467);
nand U1236 (N_1236,N_561,N_391);
nand U1237 (N_1237,N_419,N_749);
and U1238 (N_1238,N_409,N_153);
nor U1239 (N_1239,N_361,N_241);
or U1240 (N_1240,N_532,N_453);
or U1241 (N_1241,N_601,N_239);
and U1242 (N_1242,N_327,N_79);
nor U1243 (N_1243,N_495,N_196);
xor U1244 (N_1244,N_95,N_29);
nor U1245 (N_1245,N_53,N_733);
or U1246 (N_1246,N_532,N_322);
nor U1247 (N_1247,N_606,N_118);
nand U1248 (N_1248,N_238,N_465);
and U1249 (N_1249,N_555,N_118);
or U1250 (N_1250,N_96,N_508);
nor U1251 (N_1251,N_736,N_69);
nand U1252 (N_1252,N_217,N_381);
or U1253 (N_1253,N_384,N_103);
nor U1254 (N_1254,N_616,N_0);
nand U1255 (N_1255,N_624,N_611);
and U1256 (N_1256,N_315,N_292);
nand U1257 (N_1257,N_286,N_392);
or U1258 (N_1258,N_257,N_180);
nand U1259 (N_1259,N_382,N_313);
and U1260 (N_1260,N_281,N_161);
nand U1261 (N_1261,N_407,N_409);
or U1262 (N_1262,N_55,N_14);
nor U1263 (N_1263,N_20,N_346);
nor U1264 (N_1264,N_238,N_355);
or U1265 (N_1265,N_689,N_321);
xor U1266 (N_1266,N_730,N_34);
nand U1267 (N_1267,N_716,N_313);
or U1268 (N_1268,N_357,N_649);
nor U1269 (N_1269,N_218,N_502);
or U1270 (N_1270,N_6,N_230);
or U1271 (N_1271,N_42,N_73);
or U1272 (N_1272,N_338,N_644);
xnor U1273 (N_1273,N_339,N_714);
nand U1274 (N_1274,N_567,N_30);
and U1275 (N_1275,N_268,N_466);
nand U1276 (N_1276,N_426,N_663);
nor U1277 (N_1277,N_502,N_692);
or U1278 (N_1278,N_386,N_23);
nand U1279 (N_1279,N_330,N_742);
or U1280 (N_1280,N_313,N_670);
and U1281 (N_1281,N_519,N_710);
or U1282 (N_1282,N_138,N_139);
nand U1283 (N_1283,N_474,N_461);
and U1284 (N_1284,N_652,N_498);
nor U1285 (N_1285,N_432,N_512);
nor U1286 (N_1286,N_736,N_431);
nor U1287 (N_1287,N_735,N_409);
and U1288 (N_1288,N_656,N_43);
and U1289 (N_1289,N_521,N_578);
nand U1290 (N_1290,N_716,N_733);
nor U1291 (N_1291,N_510,N_28);
or U1292 (N_1292,N_316,N_300);
nand U1293 (N_1293,N_735,N_509);
or U1294 (N_1294,N_400,N_249);
nor U1295 (N_1295,N_4,N_218);
nor U1296 (N_1296,N_429,N_480);
nor U1297 (N_1297,N_152,N_484);
and U1298 (N_1298,N_319,N_184);
nand U1299 (N_1299,N_545,N_660);
nor U1300 (N_1300,N_13,N_139);
and U1301 (N_1301,N_117,N_448);
nor U1302 (N_1302,N_603,N_542);
xor U1303 (N_1303,N_557,N_319);
nand U1304 (N_1304,N_239,N_544);
nand U1305 (N_1305,N_560,N_196);
nor U1306 (N_1306,N_272,N_620);
nor U1307 (N_1307,N_423,N_728);
and U1308 (N_1308,N_564,N_601);
nand U1309 (N_1309,N_44,N_701);
and U1310 (N_1310,N_749,N_687);
nor U1311 (N_1311,N_10,N_2);
nor U1312 (N_1312,N_67,N_185);
nor U1313 (N_1313,N_220,N_590);
or U1314 (N_1314,N_459,N_355);
and U1315 (N_1315,N_49,N_360);
nand U1316 (N_1316,N_328,N_275);
or U1317 (N_1317,N_284,N_343);
and U1318 (N_1318,N_616,N_138);
or U1319 (N_1319,N_288,N_484);
or U1320 (N_1320,N_94,N_440);
nor U1321 (N_1321,N_243,N_505);
nand U1322 (N_1322,N_417,N_551);
nand U1323 (N_1323,N_386,N_528);
nor U1324 (N_1324,N_25,N_294);
or U1325 (N_1325,N_83,N_332);
or U1326 (N_1326,N_359,N_382);
nand U1327 (N_1327,N_122,N_738);
and U1328 (N_1328,N_37,N_238);
nor U1329 (N_1329,N_641,N_616);
and U1330 (N_1330,N_470,N_664);
nor U1331 (N_1331,N_474,N_116);
xor U1332 (N_1332,N_463,N_206);
and U1333 (N_1333,N_211,N_290);
nor U1334 (N_1334,N_530,N_746);
or U1335 (N_1335,N_379,N_446);
nor U1336 (N_1336,N_282,N_362);
nor U1337 (N_1337,N_467,N_153);
nand U1338 (N_1338,N_190,N_59);
and U1339 (N_1339,N_101,N_77);
nand U1340 (N_1340,N_129,N_193);
or U1341 (N_1341,N_489,N_730);
and U1342 (N_1342,N_402,N_708);
or U1343 (N_1343,N_332,N_113);
and U1344 (N_1344,N_549,N_695);
nand U1345 (N_1345,N_51,N_512);
nor U1346 (N_1346,N_141,N_350);
nand U1347 (N_1347,N_312,N_534);
nand U1348 (N_1348,N_463,N_689);
nand U1349 (N_1349,N_372,N_673);
or U1350 (N_1350,N_13,N_15);
and U1351 (N_1351,N_612,N_523);
nor U1352 (N_1352,N_371,N_27);
nor U1353 (N_1353,N_210,N_63);
nor U1354 (N_1354,N_287,N_664);
and U1355 (N_1355,N_316,N_632);
or U1356 (N_1356,N_362,N_281);
nor U1357 (N_1357,N_236,N_428);
or U1358 (N_1358,N_6,N_365);
or U1359 (N_1359,N_35,N_184);
nand U1360 (N_1360,N_207,N_219);
nor U1361 (N_1361,N_357,N_187);
and U1362 (N_1362,N_273,N_508);
nand U1363 (N_1363,N_488,N_519);
and U1364 (N_1364,N_325,N_436);
nor U1365 (N_1365,N_725,N_73);
nor U1366 (N_1366,N_619,N_34);
and U1367 (N_1367,N_225,N_356);
and U1368 (N_1368,N_19,N_239);
or U1369 (N_1369,N_92,N_424);
xor U1370 (N_1370,N_623,N_34);
nor U1371 (N_1371,N_132,N_672);
nor U1372 (N_1372,N_563,N_82);
nor U1373 (N_1373,N_513,N_272);
nor U1374 (N_1374,N_394,N_408);
or U1375 (N_1375,N_3,N_246);
and U1376 (N_1376,N_315,N_647);
nor U1377 (N_1377,N_363,N_89);
nor U1378 (N_1378,N_468,N_515);
nand U1379 (N_1379,N_716,N_420);
nand U1380 (N_1380,N_225,N_365);
or U1381 (N_1381,N_728,N_433);
and U1382 (N_1382,N_546,N_400);
nand U1383 (N_1383,N_656,N_702);
and U1384 (N_1384,N_735,N_596);
nand U1385 (N_1385,N_563,N_500);
nand U1386 (N_1386,N_742,N_645);
nand U1387 (N_1387,N_96,N_137);
and U1388 (N_1388,N_514,N_367);
nor U1389 (N_1389,N_193,N_3);
and U1390 (N_1390,N_298,N_645);
nand U1391 (N_1391,N_721,N_144);
or U1392 (N_1392,N_541,N_329);
or U1393 (N_1393,N_508,N_282);
or U1394 (N_1394,N_680,N_292);
and U1395 (N_1395,N_342,N_366);
or U1396 (N_1396,N_384,N_674);
nor U1397 (N_1397,N_32,N_489);
nand U1398 (N_1398,N_293,N_743);
and U1399 (N_1399,N_704,N_43);
and U1400 (N_1400,N_93,N_329);
or U1401 (N_1401,N_109,N_640);
nor U1402 (N_1402,N_144,N_729);
and U1403 (N_1403,N_227,N_171);
and U1404 (N_1404,N_552,N_392);
or U1405 (N_1405,N_22,N_111);
and U1406 (N_1406,N_686,N_305);
or U1407 (N_1407,N_527,N_645);
and U1408 (N_1408,N_481,N_220);
nand U1409 (N_1409,N_100,N_369);
nor U1410 (N_1410,N_189,N_527);
or U1411 (N_1411,N_645,N_22);
nand U1412 (N_1412,N_116,N_201);
and U1413 (N_1413,N_134,N_105);
or U1414 (N_1414,N_500,N_534);
or U1415 (N_1415,N_465,N_342);
and U1416 (N_1416,N_36,N_558);
or U1417 (N_1417,N_562,N_22);
nand U1418 (N_1418,N_243,N_585);
nand U1419 (N_1419,N_381,N_230);
nand U1420 (N_1420,N_272,N_292);
and U1421 (N_1421,N_152,N_123);
and U1422 (N_1422,N_677,N_42);
nand U1423 (N_1423,N_434,N_716);
and U1424 (N_1424,N_143,N_1);
nand U1425 (N_1425,N_205,N_457);
nor U1426 (N_1426,N_299,N_58);
nor U1427 (N_1427,N_285,N_395);
or U1428 (N_1428,N_447,N_200);
nor U1429 (N_1429,N_192,N_402);
and U1430 (N_1430,N_173,N_237);
and U1431 (N_1431,N_412,N_625);
nand U1432 (N_1432,N_409,N_265);
nand U1433 (N_1433,N_720,N_231);
nor U1434 (N_1434,N_220,N_460);
or U1435 (N_1435,N_597,N_49);
or U1436 (N_1436,N_411,N_691);
nand U1437 (N_1437,N_39,N_345);
or U1438 (N_1438,N_114,N_561);
nor U1439 (N_1439,N_139,N_40);
nand U1440 (N_1440,N_159,N_298);
nor U1441 (N_1441,N_130,N_525);
or U1442 (N_1442,N_240,N_748);
nor U1443 (N_1443,N_625,N_173);
nor U1444 (N_1444,N_397,N_719);
or U1445 (N_1445,N_744,N_189);
nor U1446 (N_1446,N_453,N_52);
and U1447 (N_1447,N_695,N_210);
nand U1448 (N_1448,N_330,N_551);
or U1449 (N_1449,N_427,N_226);
and U1450 (N_1450,N_426,N_512);
or U1451 (N_1451,N_376,N_112);
and U1452 (N_1452,N_440,N_421);
and U1453 (N_1453,N_716,N_643);
nand U1454 (N_1454,N_441,N_271);
xnor U1455 (N_1455,N_606,N_72);
nor U1456 (N_1456,N_544,N_594);
nand U1457 (N_1457,N_686,N_143);
nor U1458 (N_1458,N_718,N_170);
or U1459 (N_1459,N_489,N_737);
nand U1460 (N_1460,N_296,N_0);
or U1461 (N_1461,N_340,N_629);
nand U1462 (N_1462,N_135,N_528);
or U1463 (N_1463,N_627,N_748);
nor U1464 (N_1464,N_19,N_389);
nand U1465 (N_1465,N_742,N_169);
nor U1466 (N_1466,N_379,N_365);
xnor U1467 (N_1467,N_545,N_583);
and U1468 (N_1468,N_319,N_212);
nor U1469 (N_1469,N_395,N_26);
and U1470 (N_1470,N_257,N_122);
nand U1471 (N_1471,N_220,N_192);
nand U1472 (N_1472,N_136,N_498);
nand U1473 (N_1473,N_632,N_594);
and U1474 (N_1474,N_369,N_307);
nand U1475 (N_1475,N_509,N_716);
nand U1476 (N_1476,N_405,N_722);
nand U1477 (N_1477,N_403,N_675);
and U1478 (N_1478,N_713,N_173);
nor U1479 (N_1479,N_353,N_303);
or U1480 (N_1480,N_338,N_636);
or U1481 (N_1481,N_393,N_671);
or U1482 (N_1482,N_263,N_598);
xor U1483 (N_1483,N_82,N_153);
or U1484 (N_1484,N_82,N_686);
or U1485 (N_1485,N_339,N_650);
or U1486 (N_1486,N_488,N_57);
and U1487 (N_1487,N_548,N_681);
xnor U1488 (N_1488,N_715,N_519);
or U1489 (N_1489,N_405,N_380);
nor U1490 (N_1490,N_19,N_736);
and U1491 (N_1491,N_43,N_125);
or U1492 (N_1492,N_31,N_365);
and U1493 (N_1493,N_466,N_281);
or U1494 (N_1494,N_745,N_445);
nand U1495 (N_1495,N_366,N_586);
and U1496 (N_1496,N_331,N_337);
and U1497 (N_1497,N_620,N_722);
nor U1498 (N_1498,N_483,N_622);
nor U1499 (N_1499,N_532,N_480);
and U1500 (N_1500,N_1439,N_1383);
and U1501 (N_1501,N_1021,N_1233);
and U1502 (N_1502,N_1365,N_1429);
or U1503 (N_1503,N_1153,N_1098);
nand U1504 (N_1504,N_1472,N_984);
nor U1505 (N_1505,N_1020,N_1097);
and U1506 (N_1506,N_1101,N_973);
and U1507 (N_1507,N_1404,N_980);
and U1508 (N_1508,N_1119,N_1156);
or U1509 (N_1509,N_905,N_1494);
nand U1510 (N_1510,N_1238,N_840);
nand U1511 (N_1511,N_810,N_1287);
and U1512 (N_1512,N_953,N_1093);
and U1513 (N_1513,N_1416,N_963);
nand U1514 (N_1514,N_1169,N_762);
and U1515 (N_1515,N_1307,N_1133);
and U1516 (N_1516,N_1055,N_871);
or U1517 (N_1517,N_1442,N_1464);
nor U1518 (N_1518,N_879,N_1474);
or U1519 (N_1519,N_1209,N_955);
nand U1520 (N_1520,N_1360,N_1006);
nor U1521 (N_1521,N_1345,N_944);
nand U1522 (N_1522,N_870,N_885);
and U1523 (N_1523,N_881,N_1427);
nand U1524 (N_1524,N_825,N_792);
and U1525 (N_1525,N_814,N_1099);
nor U1526 (N_1526,N_1108,N_1452);
nor U1527 (N_1527,N_1149,N_750);
nand U1528 (N_1528,N_993,N_1341);
and U1529 (N_1529,N_793,N_927);
nand U1530 (N_1530,N_800,N_805);
nor U1531 (N_1531,N_1285,N_1009);
or U1532 (N_1532,N_1181,N_835);
or U1533 (N_1533,N_802,N_847);
or U1534 (N_1534,N_1121,N_1184);
and U1535 (N_1535,N_1432,N_1188);
nand U1536 (N_1536,N_796,N_1202);
nand U1537 (N_1537,N_985,N_1322);
and U1538 (N_1538,N_1206,N_1003);
nand U1539 (N_1539,N_1444,N_1157);
and U1540 (N_1540,N_755,N_1131);
nor U1541 (N_1541,N_1094,N_1061);
and U1542 (N_1542,N_1314,N_1254);
or U1543 (N_1543,N_1288,N_1273);
or U1544 (N_1544,N_1445,N_1414);
xor U1545 (N_1545,N_1419,N_1195);
nor U1546 (N_1546,N_1053,N_1304);
nor U1547 (N_1547,N_1028,N_1168);
or U1548 (N_1548,N_859,N_854);
and U1549 (N_1549,N_931,N_1357);
and U1550 (N_1550,N_756,N_1215);
or U1551 (N_1551,N_757,N_1362);
nand U1552 (N_1552,N_938,N_892);
nor U1553 (N_1553,N_777,N_783);
nor U1554 (N_1554,N_883,N_1323);
nand U1555 (N_1555,N_982,N_1282);
and U1556 (N_1556,N_1438,N_804);
and U1557 (N_1557,N_1155,N_1249);
nor U1558 (N_1558,N_781,N_1090);
nor U1559 (N_1559,N_1096,N_752);
and U1560 (N_1560,N_1493,N_1110);
nand U1561 (N_1561,N_1344,N_776);
and U1562 (N_1562,N_1312,N_1183);
nor U1563 (N_1563,N_1479,N_754);
or U1564 (N_1564,N_965,N_1011);
nand U1565 (N_1565,N_1402,N_1234);
and U1566 (N_1566,N_1431,N_1269);
or U1567 (N_1567,N_780,N_911);
and U1568 (N_1568,N_1358,N_1240);
nand U1569 (N_1569,N_1275,N_1276);
or U1570 (N_1570,N_1399,N_1220);
nor U1571 (N_1571,N_1029,N_1083);
nor U1572 (N_1572,N_994,N_832);
nor U1573 (N_1573,N_1247,N_1042);
nor U1574 (N_1574,N_1385,N_1498);
and U1575 (N_1575,N_1130,N_1303);
xor U1576 (N_1576,N_1278,N_1052);
nand U1577 (N_1577,N_1469,N_1377);
or U1578 (N_1578,N_917,N_978);
nor U1579 (N_1579,N_1113,N_1010);
nor U1580 (N_1580,N_1400,N_1151);
or U1581 (N_1581,N_1465,N_808);
and U1582 (N_1582,N_864,N_988);
and U1583 (N_1583,N_1016,N_1422);
and U1584 (N_1584,N_857,N_1332);
nand U1585 (N_1585,N_989,N_774);
nor U1586 (N_1586,N_1253,N_763);
nand U1587 (N_1587,N_1216,N_926);
and U1588 (N_1588,N_923,N_765);
nand U1589 (N_1589,N_1441,N_1271);
or U1590 (N_1590,N_1380,N_1397);
nand U1591 (N_1591,N_1144,N_1082);
and U1592 (N_1592,N_948,N_1415);
and U1593 (N_1593,N_821,N_895);
nand U1594 (N_1594,N_1484,N_1018);
and U1595 (N_1595,N_972,N_1428);
nor U1596 (N_1596,N_1281,N_971);
or U1597 (N_1597,N_1409,N_1036);
nor U1598 (N_1598,N_1148,N_891);
and U1599 (N_1599,N_1395,N_875);
nand U1600 (N_1600,N_819,N_1482);
nand U1601 (N_1601,N_1125,N_1239);
nor U1602 (N_1602,N_1297,N_934);
and U1603 (N_1603,N_760,N_913);
or U1604 (N_1604,N_924,N_1179);
or U1605 (N_1605,N_856,N_1346);
and U1606 (N_1606,N_1353,N_919);
nand U1607 (N_1607,N_1392,N_974);
nor U1608 (N_1608,N_1235,N_1229);
nor U1609 (N_1609,N_874,N_809);
or U1610 (N_1610,N_823,N_1451);
and U1611 (N_1611,N_1176,N_1057);
and U1612 (N_1612,N_1252,N_1471);
nand U1613 (N_1613,N_956,N_970);
and U1614 (N_1614,N_1076,N_1190);
nand U1615 (N_1615,N_1313,N_1124);
nor U1616 (N_1616,N_1194,N_966);
nor U1617 (N_1617,N_794,N_799);
nor U1618 (N_1618,N_1266,N_1059);
or U1619 (N_1619,N_1213,N_1349);
nand U1620 (N_1620,N_1129,N_789);
xnor U1621 (N_1621,N_795,N_1408);
nor U1622 (N_1622,N_1136,N_1167);
and U1623 (N_1623,N_1350,N_1069);
and U1624 (N_1624,N_1001,N_1348);
and U1625 (N_1625,N_1047,N_957);
and U1626 (N_1626,N_1066,N_1111);
nor U1627 (N_1627,N_1426,N_1091);
or U1628 (N_1628,N_867,N_1352);
or U1629 (N_1629,N_1489,N_910);
xor U1630 (N_1630,N_824,N_1241);
nor U1631 (N_1631,N_1243,N_837);
nor U1632 (N_1632,N_1460,N_1401);
or U1633 (N_1633,N_845,N_888);
nor U1634 (N_1634,N_1347,N_1192);
or U1635 (N_1635,N_798,N_1497);
nand U1636 (N_1636,N_1141,N_1396);
or U1637 (N_1637,N_1309,N_967);
nor U1638 (N_1638,N_1072,N_868);
or U1639 (N_1639,N_898,N_986);
nand U1640 (N_1640,N_815,N_1205);
or U1641 (N_1641,N_1175,N_813);
nor U1642 (N_1642,N_1259,N_915);
and U1643 (N_1643,N_886,N_1318);
nand U1644 (N_1644,N_1255,N_1244);
nor U1645 (N_1645,N_921,N_977);
nor U1646 (N_1646,N_1490,N_1035);
nor U1647 (N_1647,N_1476,N_1054);
or U1648 (N_1648,N_1280,N_1267);
or U1649 (N_1649,N_1319,N_1411);
nand U1650 (N_1650,N_940,N_1262);
and U1651 (N_1651,N_872,N_1370);
or U1652 (N_1652,N_1120,N_1436);
nand U1653 (N_1653,N_818,N_1227);
and U1654 (N_1654,N_1290,N_785);
and U1655 (N_1655,N_1039,N_1012);
and U1656 (N_1656,N_1116,N_1228);
nor U1657 (N_1657,N_1211,N_1456);
nor U1658 (N_1658,N_863,N_1475);
xor U1659 (N_1659,N_1005,N_849);
or U1660 (N_1660,N_1308,N_1242);
nand U1661 (N_1661,N_1163,N_894);
nand U1662 (N_1662,N_852,N_1374);
nor U1663 (N_1663,N_1434,N_1306);
or U1664 (N_1664,N_1388,N_1070);
nor U1665 (N_1665,N_1296,N_1334);
nand U1666 (N_1666,N_877,N_790);
and U1667 (N_1667,N_983,N_1300);
and U1668 (N_1668,N_1390,N_1173);
nand U1669 (N_1669,N_772,N_889);
or U1670 (N_1670,N_1421,N_1461);
or U1671 (N_1671,N_1232,N_1495);
nor U1672 (N_1672,N_1088,N_1369);
and U1673 (N_1673,N_1087,N_838);
nor U1674 (N_1674,N_860,N_811);
or U1675 (N_1675,N_1193,N_1062);
or U1676 (N_1676,N_861,N_1270);
or U1677 (N_1677,N_1305,N_1126);
nor U1678 (N_1678,N_1433,N_968);
and U1679 (N_1679,N_1201,N_1044);
nor U1680 (N_1680,N_841,N_1218);
and U1681 (N_1681,N_1085,N_1177);
nor U1682 (N_1682,N_1185,N_1407);
nand U1683 (N_1683,N_991,N_1147);
nor U1684 (N_1684,N_1260,N_908);
and U1685 (N_1685,N_1364,N_1468);
nand U1686 (N_1686,N_1135,N_1283);
nor U1687 (N_1687,N_1182,N_1132);
nand U1688 (N_1688,N_946,N_828);
nand U1689 (N_1689,N_1310,N_806);
and U1690 (N_1690,N_975,N_995);
or U1691 (N_1691,N_928,N_1292);
and U1692 (N_1692,N_1045,N_833);
and U1693 (N_1693,N_1014,N_1197);
or U1694 (N_1694,N_865,N_869);
nand U1695 (N_1695,N_941,N_1221);
or U1696 (N_1696,N_1118,N_1467);
nand U1697 (N_1697,N_1217,N_866);
or U1698 (N_1698,N_1450,N_1378);
or U1699 (N_1699,N_1140,N_1316);
nor U1700 (N_1700,N_1462,N_1100);
or U1701 (N_1701,N_1178,N_987);
or U1702 (N_1702,N_1106,N_1160);
nand U1703 (N_1703,N_1320,N_902);
or U1704 (N_1704,N_1406,N_951);
and U1705 (N_1705,N_1105,N_1298);
nor U1706 (N_1706,N_759,N_1258);
nand U1707 (N_1707,N_878,N_1373);
or U1708 (N_1708,N_1204,N_850);
or U1709 (N_1709,N_930,N_767);
nand U1710 (N_1710,N_1446,N_1079);
or U1711 (N_1711,N_1230,N_1154);
and U1712 (N_1712,N_1343,N_1123);
or U1713 (N_1713,N_803,N_1102);
nand U1714 (N_1714,N_880,N_893);
or U1715 (N_1715,N_1355,N_1004);
and U1716 (N_1716,N_788,N_769);
and U1717 (N_1717,N_1488,N_1448);
and U1718 (N_1718,N_925,N_904);
or U1719 (N_1719,N_1114,N_1339);
or U1720 (N_1720,N_1128,N_1379);
nor U1721 (N_1721,N_1172,N_1024);
nor U1722 (N_1722,N_1257,N_1331);
nand U1723 (N_1723,N_1051,N_899);
nor U1724 (N_1724,N_1231,N_969);
or U1725 (N_1725,N_1071,N_1338);
nor U1726 (N_1726,N_1226,N_1381);
nand U1727 (N_1727,N_1189,N_1470);
and U1728 (N_1728,N_914,N_1478);
nor U1729 (N_1729,N_1040,N_1394);
and U1730 (N_1730,N_1214,N_822);
or U1731 (N_1731,N_1063,N_1321);
nor U1732 (N_1732,N_1073,N_900);
nor U1733 (N_1733,N_1065,N_1127);
nand U1734 (N_1734,N_1351,N_1095);
nand U1735 (N_1735,N_1284,N_812);
nand U1736 (N_1736,N_839,N_1048);
nand U1737 (N_1737,N_1389,N_764);
nand U1738 (N_1738,N_1174,N_1222);
nor U1739 (N_1739,N_1480,N_1107);
nand U1740 (N_1740,N_920,N_801);
nand U1741 (N_1741,N_1186,N_1295);
nor U1742 (N_1742,N_1324,N_1137);
and U1743 (N_1743,N_1092,N_906);
and U1744 (N_1744,N_1210,N_1033);
or U1745 (N_1745,N_1486,N_1293);
or U1746 (N_1746,N_1064,N_981);
or U1747 (N_1747,N_1263,N_1150);
or U1748 (N_1748,N_1081,N_1405);
nand U1749 (N_1749,N_1041,N_1152);
or U1750 (N_1750,N_1356,N_922);
or U1751 (N_1751,N_836,N_844);
and U1752 (N_1752,N_964,N_1393);
or U1753 (N_1753,N_1371,N_1437);
nor U1754 (N_1754,N_761,N_1117);
or U1755 (N_1755,N_787,N_1080);
nor U1756 (N_1756,N_846,N_1315);
and U1757 (N_1757,N_829,N_990);
and U1758 (N_1758,N_943,N_1329);
nor U1759 (N_1759,N_820,N_1376);
nor U1760 (N_1760,N_1264,N_826);
and U1761 (N_1761,N_1142,N_1325);
nand U1762 (N_1762,N_1212,N_1311);
or U1763 (N_1763,N_768,N_960);
nand U1764 (N_1764,N_1291,N_1139);
nand U1765 (N_1765,N_1068,N_1333);
nor U1766 (N_1766,N_751,N_979);
or U1767 (N_1767,N_1219,N_1375);
nand U1768 (N_1768,N_1279,N_896);
or U1769 (N_1769,N_937,N_843);
or U1770 (N_1770,N_1002,N_1122);
nor U1771 (N_1771,N_1328,N_1487);
nor U1772 (N_1772,N_1340,N_918);
and U1773 (N_1773,N_1491,N_853);
or U1774 (N_1774,N_1146,N_1038);
or U1775 (N_1775,N_855,N_936);
xor U1776 (N_1776,N_1046,N_1466);
nor U1777 (N_1777,N_831,N_1089);
or U1778 (N_1778,N_1198,N_830);
nor U1779 (N_1779,N_1074,N_773);
or U1780 (N_1780,N_1224,N_1265);
nand U1781 (N_1781,N_1037,N_753);
or U1782 (N_1782,N_1457,N_1420);
nand U1783 (N_1783,N_1447,N_1022);
or U1784 (N_1784,N_1171,N_929);
or U1785 (N_1785,N_848,N_1007);
nor U1786 (N_1786,N_1200,N_1166);
and U1787 (N_1787,N_1477,N_1086);
and U1788 (N_1788,N_876,N_827);
and U1789 (N_1789,N_1372,N_935);
or U1790 (N_1790,N_947,N_976);
or U1791 (N_1791,N_1058,N_1245);
or U1792 (N_1792,N_961,N_1115);
nand U1793 (N_1793,N_1337,N_887);
nand U1794 (N_1794,N_932,N_778);
nor U1795 (N_1795,N_1251,N_1162);
nor U1796 (N_1796,N_1109,N_882);
or U1797 (N_1797,N_1361,N_1084);
or U1798 (N_1798,N_1459,N_1104);
nand U1799 (N_1799,N_766,N_1424);
nand U1800 (N_1800,N_817,N_1384);
or U1801 (N_1801,N_1391,N_916);
nand U1802 (N_1802,N_1026,N_797);
and U1803 (N_1803,N_1112,N_1196);
nand U1804 (N_1804,N_1425,N_771);
or U1805 (N_1805,N_992,N_1499);
and U1806 (N_1806,N_1056,N_912);
nor U1807 (N_1807,N_1237,N_1277);
or U1808 (N_1808,N_1386,N_1000);
or U1809 (N_1809,N_901,N_1049);
and U1810 (N_1810,N_1032,N_1492);
nor U1811 (N_1811,N_1013,N_1294);
nand U1812 (N_1812,N_1134,N_1025);
or U1813 (N_1813,N_1286,N_1027);
or U1814 (N_1814,N_1443,N_1354);
or U1815 (N_1815,N_1417,N_1382);
or U1816 (N_1816,N_1077,N_952);
nand U1817 (N_1817,N_1398,N_1256);
or U1818 (N_1818,N_770,N_1272);
and U1819 (N_1819,N_851,N_1299);
nand U1820 (N_1820,N_884,N_939);
xor U1821 (N_1821,N_816,N_1031);
nand U1822 (N_1822,N_1225,N_897);
nand U1823 (N_1823,N_784,N_1236);
nor U1824 (N_1824,N_1268,N_1145);
and U1825 (N_1825,N_1078,N_909);
or U1826 (N_1826,N_1335,N_1015);
nor U1827 (N_1827,N_1138,N_1327);
nor U1828 (N_1828,N_1423,N_958);
nand U1829 (N_1829,N_942,N_1103);
and U1830 (N_1830,N_959,N_903);
nand U1831 (N_1831,N_1199,N_1359);
or U1832 (N_1832,N_842,N_1017);
nand U1833 (N_1833,N_1060,N_1449);
nand U1834 (N_1834,N_1336,N_1250);
or U1835 (N_1835,N_1418,N_1159);
and U1836 (N_1836,N_775,N_873);
and U1837 (N_1837,N_999,N_1208);
nor U1838 (N_1838,N_1342,N_1203);
or U1839 (N_1839,N_1403,N_1248);
nand U1840 (N_1840,N_1410,N_1030);
nor U1841 (N_1841,N_834,N_907);
nand U1842 (N_1842,N_1170,N_1207);
nand U1843 (N_1843,N_1454,N_1440);
nor U1844 (N_1844,N_782,N_1330);
or U1845 (N_1845,N_1165,N_1023);
or U1846 (N_1846,N_1143,N_758);
and U1847 (N_1847,N_1075,N_1034);
nor U1848 (N_1848,N_1246,N_1161);
and U1849 (N_1849,N_1326,N_1453);
and U1850 (N_1850,N_1413,N_1067);
nand U1851 (N_1851,N_1180,N_1019);
and U1852 (N_1852,N_890,N_1455);
or U1853 (N_1853,N_1158,N_1463);
nand U1854 (N_1854,N_1301,N_1368);
nand U1855 (N_1855,N_1458,N_996);
or U1856 (N_1856,N_1164,N_1412);
or U1857 (N_1857,N_786,N_1302);
or U1858 (N_1858,N_1387,N_1481);
and U1859 (N_1859,N_950,N_1317);
nand U1860 (N_1860,N_779,N_1483);
and U1861 (N_1861,N_862,N_1261);
nand U1862 (N_1862,N_1289,N_962);
and U1863 (N_1863,N_997,N_1430);
nand U1864 (N_1864,N_1366,N_1274);
nand U1865 (N_1865,N_954,N_945);
nor U1866 (N_1866,N_1496,N_1191);
nor U1867 (N_1867,N_1435,N_1043);
nand U1868 (N_1868,N_1363,N_858);
nor U1869 (N_1869,N_933,N_1008);
nand U1870 (N_1870,N_791,N_998);
nand U1871 (N_1871,N_1485,N_1187);
and U1872 (N_1872,N_1473,N_1050);
and U1873 (N_1873,N_807,N_1367);
nand U1874 (N_1874,N_949,N_1223);
nor U1875 (N_1875,N_1477,N_1309);
nand U1876 (N_1876,N_1226,N_1258);
nand U1877 (N_1877,N_976,N_1468);
nor U1878 (N_1878,N_1207,N_1024);
nor U1879 (N_1879,N_796,N_1429);
or U1880 (N_1880,N_1382,N_1366);
nor U1881 (N_1881,N_1097,N_1349);
nor U1882 (N_1882,N_1382,N_1252);
and U1883 (N_1883,N_872,N_1156);
nand U1884 (N_1884,N_1003,N_891);
nand U1885 (N_1885,N_1236,N_1136);
nor U1886 (N_1886,N_959,N_1010);
and U1887 (N_1887,N_865,N_826);
or U1888 (N_1888,N_1002,N_1076);
or U1889 (N_1889,N_1466,N_1091);
nor U1890 (N_1890,N_978,N_1374);
nor U1891 (N_1891,N_1023,N_1100);
nand U1892 (N_1892,N_750,N_1413);
nor U1893 (N_1893,N_1029,N_1480);
nor U1894 (N_1894,N_1025,N_961);
and U1895 (N_1895,N_841,N_1272);
and U1896 (N_1896,N_1437,N_1029);
and U1897 (N_1897,N_1472,N_1462);
nand U1898 (N_1898,N_1246,N_1075);
nor U1899 (N_1899,N_1236,N_1384);
nor U1900 (N_1900,N_897,N_1097);
and U1901 (N_1901,N_753,N_1246);
and U1902 (N_1902,N_1318,N_828);
or U1903 (N_1903,N_1304,N_1355);
and U1904 (N_1904,N_827,N_1103);
nor U1905 (N_1905,N_1012,N_1051);
nand U1906 (N_1906,N_1008,N_1058);
nand U1907 (N_1907,N_974,N_1343);
and U1908 (N_1908,N_873,N_1183);
or U1909 (N_1909,N_906,N_1146);
or U1910 (N_1910,N_1273,N_1136);
and U1911 (N_1911,N_761,N_1495);
nor U1912 (N_1912,N_838,N_805);
nand U1913 (N_1913,N_1411,N_991);
nor U1914 (N_1914,N_1147,N_1375);
nor U1915 (N_1915,N_1279,N_1141);
xnor U1916 (N_1916,N_1209,N_1151);
nor U1917 (N_1917,N_1411,N_1204);
and U1918 (N_1918,N_1170,N_1112);
nand U1919 (N_1919,N_795,N_881);
nand U1920 (N_1920,N_1447,N_1269);
nor U1921 (N_1921,N_1465,N_1428);
nor U1922 (N_1922,N_1449,N_760);
nor U1923 (N_1923,N_752,N_1385);
nor U1924 (N_1924,N_913,N_1215);
and U1925 (N_1925,N_1484,N_1349);
nand U1926 (N_1926,N_896,N_761);
nand U1927 (N_1927,N_1135,N_842);
nand U1928 (N_1928,N_1284,N_1249);
nor U1929 (N_1929,N_1277,N_1325);
nor U1930 (N_1930,N_1115,N_1387);
and U1931 (N_1931,N_867,N_1197);
nand U1932 (N_1932,N_1386,N_956);
nand U1933 (N_1933,N_1262,N_1438);
nand U1934 (N_1934,N_1449,N_1483);
or U1935 (N_1935,N_1253,N_1085);
xnor U1936 (N_1936,N_1402,N_1448);
or U1937 (N_1937,N_1189,N_1145);
nor U1938 (N_1938,N_1214,N_1295);
nor U1939 (N_1939,N_1161,N_1255);
and U1940 (N_1940,N_1132,N_1463);
nor U1941 (N_1941,N_1187,N_1324);
nand U1942 (N_1942,N_791,N_1168);
nor U1943 (N_1943,N_842,N_1202);
nor U1944 (N_1944,N_1102,N_1154);
nand U1945 (N_1945,N_1143,N_1382);
and U1946 (N_1946,N_1409,N_1276);
or U1947 (N_1947,N_1343,N_937);
and U1948 (N_1948,N_1306,N_1128);
nand U1949 (N_1949,N_1068,N_1069);
and U1950 (N_1950,N_1021,N_873);
nand U1951 (N_1951,N_1040,N_1116);
nor U1952 (N_1952,N_1298,N_993);
nor U1953 (N_1953,N_769,N_1303);
nand U1954 (N_1954,N_1305,N_1096);
xor U1955 (N_1955,N_1426,N_913);
nor U1956 (N_1956,N_1214,N_1280);
or U1957 (N_1957,N_1300,N_1113);
nand U1958 (N_1958,N_1355,N_1123);
and U1959 (N_1959,N_993,N_1321);
or U1960 (N_1960,N_958,N_1343);
xor U1961 (N_1961,N_803,N_900);
nor U1962 (N_1962,N_1472,N_1194);
nand U1963 (N_1963,N_940,N_1442);
and U1964 (N_1964,N_1117,N_1013);
or U1965 (N_1965,N_1446,N_1017);
nor U1966 (N_1966,N_1141,N_897);
nand U1967 (N_1967,N_970,N_886);
and U1968 (N_1968,N_855,N_797);
and U1969 (N_1969,N_811,N_1019);
or U1970 (N_1970,N_805,N_1369);
nor U1971 (N_1971,N_1466,N_761);
or U1972 (N_1972,N_1478,N_883);
and U1973 (N_1973,N_898,N_1110);
nand U1974 (N_1974,N_1026,N_1177);
or U1975 (N_1975,N_1296,N_760);
or U1976 (N_1976,N_1283,N_811);
or U1977 (N_1977,N_1381,N_1121);
nand U1978 (N_1978,N_1051,N_1313);
nor U1979 (N_1979,N_811,N_996);
nor U1980 (N_1980,N_1496,N_776);
nand U1981 (N_1981,N_958,N_1009);
or U1982 (N_1982,N_1443,N_1379);
and U1983 (N_1983,N_1168,N_938);
or U1984 (N_1984,N_1357,N_1394);
nor U1985 (N_1985,N_977,N_1412);
nor U1986 (N_1986,N_1285,N_1252);
nor U1987 (N_1987,N_1054,N_940);
nand U1988 (N_1988,N_1317,N_1244);
nand U1989 (N_1989,N_1317,N_1102);
and U1990 (N_1990,N_1488,N_1009);
or U1991 (N_1991,N_1220,N_1002);
nand U1992 (N_1992,N_1071,N_1207);
or U1993 (N_1993,N_950,N_819);
or U1994 (N_1994,N_1420,N_1337);
nor U1995 (N_1995,N_1161,N_1006);
nand U1996 (N_1996,N_898,N_824);
nor U1997 (N_1997,N_874,N_1122);
nand U1998 (N_1998,N_751,N_1310);
nand U1999 (N_1999,N_1001,N_1095);
nand U2000 (N_2000,N_1049,N_850);
or U2001 (N_2001,N_1015,N_1370);
or U2002 (N_2002,N_1052,N_1041);
or U2003 (N_2003,N_890,N_1458);
nand U2004 (N_2004,N_1128,N_898);
nand U2005 (N_2005,N_1436,N_1110);
or U2006 (N_2006,N_1470,N_1377);
and U2007 (N_2007,N_1279,N_1182);
and U2008 (N_2008,N_1018,N_1180);
nor U2009 (N_2009,N_798,N_954);
and U2010 (N_2010,N_1206,N_1160);
and U2011 (N_2011,N_1467,N_1204);
and U2012 (N_2012,N_1167,N_1012);
nor U2013 (N_2013,N_1322,N_1393);
nand U2014 (N_2014,N_1033,N_1080);
or U2015 (N_2015,N_778,N_1321);
and U2016 (N_2016,N_1237,N_1273);
nand U2017 (N_2017,N_959,N_1155);
nand U2018 (N_2018,N_918,N_861);
and U2019 (N_2019,N_1249,N_1313);
or U2020 (N_2020,N_1394,N_951);
nor U2021 (N_2021,N_1121,N_792);
nand U2022 (N_2022,N_928,N_1340);
nand U2023 (N_2023,N_1240,N_1315);
and U2024 (N_2024,N_1115,N_814);
nor U2025 (N_2025,N_1369,N_857);
or U2026 (N_2026,N_852,N_1393);
nor U2027 (N_2027,N_1399,N_999);
or U2028 (N_2028,N_885,N_993);
and U2029 (N_2029,N_954,N_1001);
nor U2030 (N_2030,N_1008,N_1409);
or U2031 (N_2031,N_832,N_933);
and U2032 (N_2032,N_940,N_1093);
nor U2033 (N_2033,N_919,N_1088);
nor U2034 (N_2034,N_1466,N_915);
nor U2035 (N_2035,N_797,N_954);
or U2036 (N_2036,N_914,N_986);
nand U2037 (N_2037,N_1064,N_1229);
and U2038 (N_2038,N_813,N_1421);
or U2039 (N_2039,N_1380,N_892);
nand U2040 (N_2040,N_1344,N_1261);
and U2041 (N_2041,N_916,N_1313);
xor U2042 (N_2042,N_1306,N_803);
xnor U2043 (N_2043,N_997,N_1391);
nand U2044 (N_2044,N_1111,N_1095);
nand U2045 (N_2045,N_843,N_1420);
nand U2046 (N_2046,N_1302,N_1247);
and U2047 (N_2047,N_1428,N_1490);
or U2048 (N_2048,N_1225,N_1326);
nand U2049 (N_2049,N_1439,N_867);
nand U2050 (N_2050,N_865,N_1052);
nor U2051 (N_2051,N_1314,N_870);
nand U2052 (N_2052,N_1347,N_853);
and U2053 (N_2053,N_1348,N_1168);
nor U2054 (N_2054,N_1053,N_1323);
nor U2055 (N_2055,N_1037,N_1022);
nand U2056 (N_2056,N_1221,N_1043);
nand U2057 (N_2057,N_1497,N_1352);
nor U2058 (N_2058,N_1049,N_1403);
nor U2059 (N_2059,N_1086,N_1471);
nand U2060 (N_2060,N_1216,N_945);
nand U2061 (N_2061,N_1235,N_837);
nor U2062 (N_2062,N_862,N_1472);
nand U2063 (N_2063,N_836,N_953);
or U2064 (N_2064,N_1108,N_930);
nor U2065 (N_2065,N_892,N_1405);
nand U2066 (N_2066,N_938,N_1475);
nand U2067 (N_2067,N_1312,N_902);
or U2068 (N_2068,N_918,N_1144);
and U2069 (N_2069,N_1218,N_1108);
nand U2070 (N_2070,N_809,N_1257);
nor U2071 (N_2071,N_1444,N_781);
or U2072 (N_2072,N_753,N_1089);
and U2073 (N_2073,N_975,N_1455);
nor U2074 (N_2074,N_864,N_1452);
and U2075 (N_2075,N_1152,N_1134);
or U2076 (N_2076,N_1046,N_1125);
nand U2077 (N_2077,N_804,N_1013);
nand U2078 (N_2078,N_1434,N_1484);
and U2079 (N_2079,N_1227,N_1441);
and U2080 (N_2080,N_1493,N_932);
and U2081 (N_2081,N_917,N_1133);
or U2082 (N_2082,N_1075,N_1256);
or U2083 (N_2083,N_1352,N_1222);
nor U2084 (N_2084,N_1459,N_1274);
or U2085 (N_2085,N_1054,N_765);
nand U2086 (N_2086,N_825,N_1404);
nand U2087 (N_2087,N_927,N_1102);
and U2088 (N_2088,N_1076,N_839);
nor U2089 (N_2089,N_1224,N_1413);
nor U2090 (N_2090,N_1395,N_1445);
xor U2091 (N_2091,N_795,N_1397);
nor U2092 (N_2092,N_835,N_1199);
or U2093 (N_2093,N_841,N_832);
nor U2094 (N_2094,N_1362,N_1378);
and U2095 (N_2095,N_920,N_1324);
nand U2096 (N_2096,N_792,N_1242);
nor U2097 (N_2097,N_1390,N_1284);
nor U2098 (N_2098,N_1140,N_1024);
nor U2099 (N_2099,N_899,N_1009);
nand U2100 (N_2100,N_1101,N_1410);
nand U2101 (N_2101,N_1247,N_856);
nor U2102 (N_2102,N_855,N_949);
or U2103 (N_2103,N_1389,N_1121);
or U2104 (N_2104,N_1186,N_1242);
nor U2105 (N_2105,N_1476,N_970);
nor U2106 (N_2106,N_1052,N_789);
or U2107 (N_2107,N_1371,N_1021);
and U2108 (N_2108,N_1089,N_1096);
or U2109 (N_2109,N_1199,N_1384);
nand U2110 (N_2110,N_1196,N_1187);
or U2111 (N_2111,N_998,N_1044);
or U2112 (N_2112,N_1224,N_1373);
and U2113 (N_2113,N_1184,N_1220);
nand U2114 (N_2114,N_752,N_1049);
nor U2115 (N_2115,N_1364,N_1464);
nand U2116 (N_2116,N_936,N_1170);
and U2117 (N_2117,N_1038,N_759);
and U2118 (N_2118,N_1496,N_1209);
nand U2119 (N_2119,N_1071,N_1136);
or U2120 (N_2120,N_963,N_1261);
or U2121 (N_2121,N_1274,N_1410);
xor U2122 (N_2122,N_1006,N_844);
or U2123 (N_2123,N_1190,N_1265);
nor U2124 (N_2124,N_828,N_1295);
or U2125 (N_2125,N_1284,N_763);
or U2126 (N_2126,N_1360,N_1365);
or U2127 (N_2127,N_853,N_1098);
nor U2128 (N_2128,N_1346,N_962);
or U2129 (N_2129,N_1307,N_963);
or U2130 (N_2130,N_1213,N_1148);
nand U2131 (N_2131,N_1320,N_957);
or U2132 (N_2132,N_1167,N_1201);
or U2133 (N_2133,N_884,N_1303);
and U2134 (N_2134,N_1126,N_1341);
nor U2135 (N_2135,N_1398,N_1358);
nand U2136 (N_2136,N_1481,N_1261);
nor U2137 (N_2137,N_837,N_1430);
nor U2138 (N_2138,N_795,N_1450);
nor U2139 (N_2139,N_1279,N_1080);
or U2140 (N_2140,N_929,N_1045);
and U2141 (N_2141,N_1157,N_1347);
nor U2142 (N_2142,N_910,N_872);
and U2143 (N_2143,N_888,N_1158);
nand U2144 (N_2144,N_825,N_794);
nand U2145 (N_2145,N_1312,N_1063);
nor U2146 (N_2146,N_1471,N_762);
and U2147 (N_2147,N_1215,N_858);
or U2148 (N_2148,N_1462,N_1207);
nand U2149 (N_2149,N_844,N_1041);
and U2150 (N_2150,N_849,N_902);
or U2151 (N_2151,N_1380,N_1440);
or U2152 (N_2152,N_783,N_821);
nand U2153 (N_2153,N_846,N_1231);
nand U2154 (N_2154,N_819,N_1466);
nor U2155 (N_2155,N_1149,N_1341);
or U2156 (N_2156,N_827,N_1360);
nor U2157 (N_2157,N_820,N_1359);
or U2158 (N_2158,N_1243,N_1199);
nor U2159 (N_2159,N_1352,N_1093);
nor U2160 (N_2160,N_1322,N_1222);
and U2161 (N_2161,N_1420,N_770);
or U2162 (N_2162,N_1132,N_1017);
and U2163 (N_2163,N_1343,N_966);
and U2164 (N_2164,N_890,N_1135);
and U2165 (N_2165,N_1050,N_832);
nand U2166 (N_2166,N_941,N_1406);
and U2167 (N_2167,N_1317,N_1143);
and U2168 (N_2168,N_1234,N_852);
nor U2169 (N_2169,N_1090,N_978);
and U2170 (N_2170,N_1288,N_913);
nand U2171 (N_2171,N_1420,N_1026);
nor U2172 (N_2172,N_1325,N_951);
nand U2173 (N_2173,N_1258,N_774);
and U2174 (N_2174,N_870,N_760);
xnor U2175 (N_2175,N_1427,N_1402);
nand U2176 (N_2176,N_1073,N_1011);
nand U2177 (N_2177,N_828,N_1291);
nand U2178 (N_2178,N_843,N_1443);
nor U2179 (N_2179,N_1018,N_1037);
or U2180 (N_2180,N_1240,N_1127);
or U2181 (N_2181,N_1336,N_834);
nand U2182 (N_2182,N_764,N_1239);
xor U2183 (N_2183,N_1218,N_1245);
and U2184 (N_2184,N_863,N_1484);
or U2185 (N_2185,N_1066,N_1466);
or U2186 (N_2186,N_785,N_1219);
nand U2187 (N_2187,N_946,N_1267);
or U2188 (N_2188,N_1022,N_910);
nand U2189 (N_2189,N_1022,N_1067);
nand U2190 (N_2190,N_1189,N_1324);
nand U2191 (N_2191,N_1394,N_1237);
nor U2192 (N_2192,N_1099,N_755);
nor U2193 (N_2193,N_1287,N_1196);
xnor U2194 (N_2194,N_1463,N_810);
nor U2195 (N_2195,N_781,N_1066);
nor U2196 (N_2196,N_1088,N_936);
nand U2197 (N_2197,N_1158,N_1442);
nand U2198 (N_2198,N_1273,N_819);
xor U2199 (N_2199,N_1353,N_1290);
nor U2200 (N_2200,N_1002,N_1234);
nor U2201 (N_2201,N_1166,N_994);
and U2202 (N_2202,N_1105,N_1232);
and U2203 (N_2203,N_894,N_1367);
nand U2204 (N_2204,N_1330,N_946);
and U2205 (N_2205,N_1482,N_1031);
and U2206 (N_2206,N_769,N_1162);
nor U2207 (N_2207,N_910,N_1324);
nor U2208 (N_2208,N_1242,N_1157);
and U2209 (N_2209,N_1371,N_1436);
nand U2210 (N_2210,N_791,N_1451);
and U2211 (N_2211,N_1426,N_1345);
nor U2212 (N_2212,N_1470,N_1105);
and U2213 (N_2213,N_1205,N_1189);
nor U2214 (N_2214,N_772,N_1343);
or U2215 (N_2215,N_1053,N_995);
and U2216 (N_2216,N_757,N_1043);
or U2217 (N_2217,N_1125,N_1481);
and U2218 (N_2218,N_1110,N_1117);
nand U2219 (N_2219,N_990,N_1020);
nand U2220 (N_2220,N_892,N_1397);
or U2221 (N_2221,N_1454,N_972);
and U2222 (N_2222,N_1154,N_1477);
nor U2223 (N_2223,N_1041,N_865);
nand U2224 (N_2224,N_801,N_1376);
nand U2225 (N_2225,N_1231,N_1104);
nand U2226 (N_2226,N_1059,N_869);
and U2227 (N_2227,N_1460,N_945);
or U2228 (N_2228,N_1440,N_1231);
nand U2229 (N_2229,N_1013,N_1353);
or U2230 (N_2230,N_1263,N_907);
nand U2231 (N_2231,N_1339,N_1383);
or U2232 (N_2232,N_887,N_1426);
nor U2233 (N_2233,N_1129,N_1319);
and U2234 (N_2234,N_1300,N_1194);
and U2235 (N_2235,N_1243,N_815);
nand U2236 (N_2236,N_888,N_1311);
nand U2237 (N_2237,N_1109,N_1060);
xnor U2238 (N_2238,N_1083,N_1000);
or U2239 (N_2239,N_1070,N_1146);
nand U2240 (N_2240,N_1131,N_803);
or U2241 (N_2241,N_819,N_966);
and U2242 (N_2242,N_993,N_1096);
nand U2243 (N_2243,N_1189,N_1144);
or U2244 (N_2244,N_1131,N_1114);
or U2245 (N_2245,N_1200,N_939);
or U2246 (N_2246,N_1151,N_1360);
nand U2247 (N_2247,N_929,N_1164);
nand U2248 (N_2248,N_859,N_1270);
nor U2249 (N_2249,N_1165,N_1321);
nand U2250 (N_2250,N_1950,N_1947);
nor U2251 (N_2251,N_1753,N_2181);
or U2252 (N_2252,N_1906,N_1583);
and U2253 (N_2253,N_2086,N_1995);
nand U2254 (N_2254,N_1930,N_1652);
or U2255 (N_2255,N_1576,N_1986);
nand U2256 (N_2256,N_2162,N_1566);
and U2257 (N_2257,N_1650,N_1554);
nor U2258 (N_2258,N_1864,N_1748);
nor U2259 (N_2259,N_2075,N_1861);
xnor U2260 (N_2260,N_1700,N_1636);
or U2261 (N_2261,N_1705,N_1832);
and U2262 (N_2262,N_1506,N_2087);
or U2263 (N_2263,N_1970,N_1779);
nor U2264 (N_2264,N_1967,N_2018);
and U2265 (N_2265,N_1815,N_1546);
nor U2266 (N_2266,N_2141,N_1642);
and U2267 (N_2267,N_2208,N_1920);
and U2268 (N_2268,N_1818,N_1616);
and U2269 (N_2269,N_1573,N_1527);
nor U2270 (N_2270,N_2022,N_1728);
nor U2271 (N_2271,N_2182,N_2165);
or U2272 (N_2272,N_1846,N_1773);
nor U2273 (N_2273,N_2079,N_1828);
nor U2274 (N_2274,N_2111,N_1688);
and U2275 (N_2275,N_1678,N_2107);
and U2276 (N_2276,N_2068,N_1833);
and U2277 (N_2277,N_2012,N_2130);
nor U2278 (N_2278,N_2136,N_1741);
or U2279 (N_2279,N_2209,N_1765);
or U2280 (N_2280,N_1579,N_1683);
nor U2281 (N_2281,N_1876,N_2194);
nor U2282 (N_2282,N_1697,N_1751);
nor U2283 (N_2283,N_1989,N_2016);
nor U2284 (N_2284,N_1682,N_1591);
nand U2285 (N_2285,N_1851,N_1507);
and U2286 (N_2286,N_1707,N_1919);
and U2287 (N_2287,N_1536,N_2216);
or U2288 (N_2288,N_2221,N_1586);
nand U2289 (N_2289,N_1676,N_1848);
and U2290 (N_2290,N_1831,N_1973);
nor U2291 (N_2291,N_2051,N_1549);
nand U2292 (N_2292,N_1626,N_1900);
or U2293 (N_2293,N_1834,N_1996);
or U2294 (N_2294,N_2071,N_1574);
nand U2295 (N_2295,N_1843,N_1913);
and U2296 (N_2296,N_1879,N_2242);
nand U2297 (N_2297,N_2233,N_1835);
and U2298 (N_2298,N_1607,N_2142);
nand U2299 (N_2299,N_1839,N_1551);
or U2300 (N_2300,N_1729,N_2043);
nor U2301 (N_2301,N_1824,N_2057);
nand U2302 (N_2302,N_1608,N_2210);
nor U2303 (N_2303,N_1672,N_1597);
xor U2304 (N_2304,N_1810,N_1780);
nor U2305 (N_2305,N_1965,N_2054);
nand U2306 (N_2306,N_1770,N_2153);
nor U2307 (N_2307,N_1885,N_2037);
or U2308 (N_2308,N_1886,N_2249);
nand U2309 (N_2309,N_1977,N_2244);
nor U2310 (N_2310,N_1580,N_2188);
nor U2311 (N_2311,N_2005,N_1987);
and U2312 (N_2312,N_1685,N_1908);
and U2313 (N_2313,N_1840,N_1791);
nor U2314 (N_2314,N_1658,N_1881);
or U2315 (N_2315,N_1797,N_1830);
nand U2316 (N_2316,N_1804,N_2118);
nand U2317 (N_2317,N_1960,N_1798);
and U2318 (N_2318,N_1620,N_2083);
nor U2319 (N_2319,N_1905,N_2028);
nor U2320 (N_2320,N_1531,N_2225);
nand U2321 (N_2321,N_2157,N_1736);
nor U2322 (N_2322,N_2082,N_1638);
nor U2323 (N_2323,N_1602,N_1558);
nor U2324 (N_2324,N_2186,N_1954);
nor U2325 (N_2325,N_2085,N_2236);
and U2326 (N_2326,N_2205,N_2102);
or U2327 (N_2327,N_1647,N_1553);
nor U2328 (N_2328,N_1624,N_1855);
xor U2329 (N_2329,N_1568,N_1702);
and U2330 (N_2330,N_2040,N_2036);
and U2331 (N_2331,N_1789,N_1595);
nor U2332 (N_2332,N_1587,N_1541);
or U2333 (N_2333,N_2089,N_2062);
and U2334 (N_2334,N_1726,N_2219);
nand U2335 (N_2335,N_1867,N_2148);
or U2336 (N_2336,N_2121,N_2227);
and U2337 (N_2337,N_1860,N_1699);
nand U2338 (N_2338,N_2211,N_1788);
or U2339 (N_2339,N_1966,N_2047);
nor U2340 (N_2340,N_1775,N_1984);
nand U2341 (N_2341,N_1863,N_2055);
nor U2342 (N_2342,N_2127,N_1749);
and U2343 (N_2343,N_1983,N_1763);
nor U2344 (N_2344,N_1552,N_2091);
nor U2345 (N_2345,N_2061,N_1991);
and U2346 (N_2346,N_1884,N_1785);
nor U2347 (N_2347,N_2008,N_1817);
nand U2348 (N_2348,N_1777,N_1956);
or U2349 (N_2349,N_2046,N_1899);
xor U2350 (N_2350,N_2222,N_2017);
and U2351 (N_2351,N_1515,N_1730);
nor U2352 (N_2352,N_2213,N_1878);
and U2353 (N_2353,N_2030,N_1517);
or U2354 (N_2354,N_1963,N_1644);
nand U2355 (N_2355,N_2131,N_1868);
nor U2356 (N_2356,N_2101,N_2137);
and U2357 (N_2357,N_1955,N_1819);
nand U2358 (N_2358,N_1961,N_1656);
nor U2359 (N_2359,N_1992,N_1520);
nand U2360 (N_2360,N_2093,N_2139);
or U2361 (N_2361,N_2167,N_1938);
and U2362 (N_2362,N_1888,N_1945);
nor U2363 (N_2363,N_2041,N_1891);
nand U2364 (N_2364,N_2081,N_1925);
nand U2365 (N_2365,N_1928,N_1927);
or U2366 (N_2366,N_1567,N_1661);
or U2367 (N_2367,N_1714,N_1572);
and U2368 (N_2368,N_1924,N_2064);
or U2369 (N_2369,N_1903,N_1766);
and U2370 (N_2370,N_2066,N_1752);
and U2371 (N_2371,N_1943,N_2033);
or U2372 (N_2372,N_1663,N_2224);
nor U2373 (N_2373,N_1942,N_1525);
or U2374 (N_2374,N_1666,N_1933);
nand U2375 (N_2375,N_2007,N_2193);
or U2376 (N_2376,N_2214,N_1904);
nor U2377 (N_2377,N_1994,N_1631);
and U2378 (N_2378,N_1964,N_1865);
nand U2379 (N_2379,N_2078,N_2246);
nand U2380 (N_2380,N_1962,N_1600);
and U2381 (N_2381,N_1706,N_1821);
nor U2382 (N_2382,N_2060,N_1915);
nand U2383 (N_2383,N_2084,N_1719);
and U2384 (N_2384,N_1853,N_1912);
nor U2385 (N_2385,N_1701,N_1800);
nand U2386 (N_2386,N_1784,N_1612);
nor U2387 (N_2387,N_2226,N_2126);
nand U2388 (N_2388,N_1738,N_1548);
nor U2389 (N_2389,N_1570,N_1849);
and U2390 (N_2390,N_1988,N_1764);
and U2391 (N_2391,N_2109,N_1922);
nor U2392 (N_2392,N_2110,N_1571);
nand U2393 (N_2393,N_1926,N_1618);
or U2394 (N_2394,N_1794,N_1911);
and U2395 (N_2395,N_1841,N_1510);
nand U2396 (N_2396,N_2166,N_1617);
and U2397 (N_2397,N_1565,N_1603);
nor U2398 (N_2398,N_1890,N_1621);
or U2399 (N_2399,N_2147,N_2014);
and U2400 (N_2400,N_1660,N_1653);
or U2401 (N_2401,N_1781,N_2088);
nor U2402 (N_2402,N_1792,N_2095);
nand U2403 (N_2403,N_2099,N_1873);
or U2404 (N_2404,N_1856,N_1916);
nor U2405 (N_2405,N_2065,N_1585);
nor U2406 (N_2406,N_2230,N_1783);
or U2407 (N_2407,N_2070,N_1556);
nor U2408 (N_2408,N_1669,N_1655);
nor U2409 (N_2409,N_1921,N_1615);
nor U2410 (N_2410,N_1543,N_1858);
nor U2411 (N_2411,N_1874,N_1667);
and U2412 (N_2412,N_1664,N_2117);
nor U2413 (N_2413,N_1599,N_2234);
nor U2414 (N_2414,N_2027,N_2056);
nor U2415 (N_2415,N_1695,N_1809);
nor U2416 (N_2416,N_2123,N_1820);
nor U2417 (N_2417,N_1540,N_1516);
or U2418 (N_2418,N_1501,N_1716);
nor U2419 (N_2419,N_1949,N_2052);
xnor U2420 (N_2420,N_1518,N_1997);
nand U2421 (N_2421,N_1657,N_2164);
or U2422 (N_2422,N_1936,N_2067);
or U2423 (N_2423,N_1643,N_2145);
nand U2424 (N_2424,N_1625,N_2231);
nand U2425 (N_2425,N_1931,N_1768);
nor U2426 (N_2426,N_1774,N_1606);
or U2427 (N_2427,N_2152,N_1569);
nand U2428 (N_2428,N_1948,N_2198);
nand U2429 (N_2429,N_1604,N_1564);
and U2430 (N_2430,N_1668,N_2232);
nor U2431 (N_2431,N_1634,N_2175);
or U2432 (N_2432,N_1557,N_1715);
nor U2433 (N_2433,N_1723,N_1806);
nor U2434 (N_2434,N_1718,N_1635);
and U2435 (N_2435,N_1929,N_2160);
nor U2436 (N_2436,N_1639,N_1584);
nand U2437 (N_2437,N_2245,N_2158);
nand U2438 (N_2438,N_2090,N_2119);
nand U2439 (N_2439,N_1629,N_1980);
or U2440 (N_2440,N_1681,N_1786);
nand U2441 (N_2441,N_1686,N_1665);
and U2442 (N_2442,N_2223,N_1513);
nor U2443 (N_2443,N_1852,N_1526);
or U2444 (N_2444,N_1838,N_2228);
or U2445 (N_2445,N_1578,N_1892);
nand U2446 (N_2446,N_1522,N_1757);
or U2447 (N_2447,N_2034,N_1512);
nand U2448 (N_2448,N_1827,N_2023);
nor U2449 (N_2449,N_2106,N_1914);
and U2450 (N_2450,N_1503,N_1857);
nor U2451 (N_2451,N_1813,N_1509);
and U2452 (N_2452,N_2200,N_1596);
and U2453 (N_2453,N_2020,N_1673);
and U2454 (N_2454,N_1850,N_2132);
nor U2455 (N_2455,N_2206,N_2176);
and U2456 (N_2456,N_1589,N_2026);
nand U2457 (N_2457,N_2174,N_1897);
and U2458 (N_2458,N_2044,N_2006);
nor U2459 (N_2459,N_1677,N_1659);
or U2460 (N_2460,N_1999,N_2019);
or U2461 (N_2461,N_1799,N_1769);
nor U2462 (N_2462,N_2190,N_1590);
nand U2463 (N_2463,N_1880,N_1941);
nand U2464 (N_2464,N_1862,N_2191);
nand U2465 (N_2465,N_1684,N_1918);
nor U2466 (N_2466,N_1692,N_1993);
xor U2467 (N_2467,N_1640,N_1633);
or U2468 (N_2468,N_2024,N_1611);
or U2469 (N_2469,N_2077,N_1743);
or U2470 (N_2470,N_1796,N_1981);
nand U2471 (N_2471,N_1776,N_2204);
and U2472 (N_2472,N_1645,N_2217);
nand U2473 (N_2473,N_1690,N_1829);
and U2474 (N_2474,N_1519,N_1812);
and U2475 (N_2475,N_1917,N_2021);
and U2476 (N_2476,N_1720,N_2015);
nand U2477 (N_2477,N_2159,N_1985);
and U2478 (N_2478,N_1560,N_1674);
nand U2479 (N_2479,N_1952,N_1725);
or U2480 (N_2480,N_2241,N_1538);
or U2481 (N_2481,N_2058,N_1555);
nand U2482 (N_2482,N_2180,N_2049);
nand U2483 (N_2483,N_1883,N_1935);
nand U2484 (N_2484,N_1907,N_2187);
nand U2485 (N_2485,N_2002,N_1593);
and U2486 (N_2486,N_2154,N_1524);
and U2487 (N_2487,N_2185,N_2025);
nand U2488 (N_2488,N_1958,N_1610);
or U2489 (N_2489,N_1708,N_2150);
and U2490 (N_2490,N_1940,N_1641);
and U2491 (N_2491,N_2218,N_1619);
and U2492 (N_2492,N_2120,N_1544);
and U2493 (N_2493,N_2240,N_2010);
nor U2494 (N_2494,N_2011,N_2161);
and U2495 (N_2495,N_1649,N_1713);
xor U2496 (N_2496,N_1782,N_2146);
nor U2497 (N_2497,N_1790,N_1795);
and U2498 (N_2498,N_1547,N_2009);
and U2499 (N_2499,N_1894,N_2196);
and U2500 (N_2500,N_2094,N_2122);
nand U2501 (N_2501,N_1534,N_1530);
and U2502 (N_2502,N_2202,N_1953);
nand U2503 (N_2503,N_2097,N_2201);
and U2504 (N_2504,N_2113,N_1500);
or U2505 (N_2505,N_2247,N_1968);
nor U2506 (N_2506,N_2104,N_1528);
nor U2507 (N_2507,N_1979,N_1703);
nor U2508 (N_2508,N_2173,N_1837);
or U2509 (N_2509,N_2013,N_2172);
or U2510 (N_2510,N_2069,N_2238);
nor U2511 (N_2511,N_1577,N_1654);
and U2512 (N_2512,N_1651,N_2135);
nor U2513 (N_2513,N_2073,N_2045);
nand U2514 (N_2514,N_1533,N_1711);
nand U2515 (N_2515,N_2098,N_1733);
nand U2516 (N_2516,N_2092,N_2129);
nor U2517 (N_2517,N_1724,N_1825);
nor U2518 (N_2518,N_1679,N_2053);
and U2519 (N_2519,N_1539,N_1693);
or U2520 (N_2520,N_1755,N_1628);
nor U2521 (N_2521,N_1737,N_2063);
and U2522 (N_2522,N_1759,N_1974);
nor U2523 (N_2523,N_1854,N_1923);
nor U2524 (N_2524,N_1767,N_2115);
nand U2525 (N_2525,N_1739,N_1605);
and U2526 (N_2526,N_1866,N_1982);
nor U2527 (N_2527,N_1882,N_1717);
and U2528 (N_2528,N_1823,N_1559);
nand U2529 (N_2529,N_1502,N_1563);
and U2530 (N_2530,N_2163,N_2103);
nor U2531 (N_2531,N_1756,N_1762);
and U2532 (N_2532,N_1601,N_2229);
or U2533 (N_2533,N_1511,N_1870);
or U2534 (N_2534,N_2171,N_1869);
and U2535 (N_2535,N_2004,N_1550);
nand U2536 (N_2536,N_1895,N_2000);
and U2537 (N_2537,N_1978,N_2042);
nand U2538 (N_2538,N_2177,N_1807);
nor U2539 (N_2539,N_2212,N_2105);
or U2540 (N_2540,N_1801,N_1630);
or U2541 (N_2541,N_2003,N_2203);
and U2542 (N_2542,N_1562,N_2235);
and U2543 (N_2543,N_1902,N_2001);
or U2544 (N_2544,N_2100,N_1646);
and U2545 (N_2545,N_2133,N_1529);
and U2546 (N_2546,N_1910,N_1976);
or U2547 (N_2547,N_1814,N_2168);
and U2548 (N_2548,N_1742,N_1722);
and U2549 (N_2549,N_1731,N_1893);
nand U2550 (N_2550,N_1842,N_1712);
and U2551 (N_2551,N_1581,N_1521);
and U2552 (N_2552,N_2108,N_1632);
and U2553 (N_2553,N_1710,N_2125);
nor U2554 (N_2554,N_1747,N_1746);
or U2555 (N_2555,N_2134,N_1836);
and U2556 (N_2556,N_1575,N_1592);
and U2557 (N_2557,N_1946,N_1847);
nand U2558 (N_2558,N_1696,N_1594);
nand U2559 (N_2559,N_1990,N_1998);
nor U2560 (N_2560,N_1505,N_1971);
nor U2561 (N_2561,N_2038,N_1959);
nand U2562 (N_2562,N_2207,N_1871);
nand U2563 (N_2563,N_1735,N_1901);
or U2564 (N_2564,N_2059,N_1535);
and U2565 (N_2565,N_2076,N_2050);
nor U2566 (N_2566,N_1537,N_2029);
or U2567 (N_2567,N_1808,N_2156);
or U2568 (N_2568,N_2215,N_2128);
nand U2569 (N_2569,N_2143,N_1859);
nand U2570 (N_2570,N_1627,N_2197);
nand U2571 (N_2571,N_1691,N_1675);
nand U2572 (N_2572,N_2032,N_1803);
nand U2573 (N_2573,N_1637,N_1889);
and U2574 (N_2574,N_1523,N_1898);
nand U2575 (N_2575,N_1771,N_1740);
or U2576 (N_2576,N_1614,N_2114);
or U2577 (N_2577,N_1975,N_1877);
nor U2578 (N_2578,N_1793,N_1772);
or U2579 (N_2579,N_1758,N_2124);
and U2580 (N_2580,N_1802,N_1745);
and U2581 (N_2581,N_1778,N_2096);
or U2582 (N_2582,N_2195,N_1545);
nand U2583 (N_2583,N_2192,N_1582);
and U2584 (N_2584,N_1875,N_1721);
nand U2585 (N_2585,N_2243,N_2035);
nand U2586 (N_2586,N_1613,N_1887);
and U2587 (N_2587,N_2199,N_1687);
and U2588 (N_2588,N_1727,N_2183);
nand U2589 (N_2589,N_2072,N_2151);
nand U2590 (N_2590,N_1542,N_1909);
or U2591 (N_2591,N_1532,N_1972);
and U2592 (N_2592,N_2144,N_2138);
nand U2593 (N_2593,N_1732,N_1514);
and U2594 (N_2594,N_1761,N_1957);
nand U2595 (N_2595,N_1934,N_1760);
nand U2596 (N_2596,N_1932,N_1623);
nand U2597 (N_2597,N_1822,N_1845);
xor U2598 (N_2598,N_1671,N_2155);
nand U2599 (N_2599,N_1704,N_1844);
nor U2600 (N_2600,N_1670,N_1504);
nor U2601 (N_2601,N_2149,N_2039);
nand U2602 (N_2602,N_2048,N_1694);
and U2603 (N_2603,N_1937,N_1939);
xnor U2604 (N_2604,N_2074,N_1750);
and U2605 (N_2605,N_1689,N_1969);
nand U2606 (N_2606,N_2178,N_2179);
nand U2607 (N_2607,N_1944,N_2220);
or U2608 (N_2608,N_2031,N_1734);
and U2609 (N_2609,N_2237,N_1662);
nor U2610 (N_2610,N_1805,N_2248);
nor U2611 (N_2611,N_1787,N_1826);
nor U2612 (N_2612,N_2112,N_1648);
nor U2613 (N_2613,N_2239,N_1588);
and U2614 (N_2614,N_1811,N_2189);
nor U2615 (N_2615,N_1698,N_2116);
and U2616 (N_2616,N_1754,N_1561);
nand U2617 (N_2617,N_2080,N_1816);
nand U2618 (N_2618,N_2140,N_1951);
nand U2619 (N_2619,N_1744,N_2170);
nor U2620 (N_2620,N_1622,N_1609);
nor U2621 (N_2621,N_1508,N_1872);
nor U2622 (N_2622,N_1709,N_1598);
nand U2623 (N_2623,N_1680,N_1896);
or U2624 (N_2624,N_2169,N_2184);
nand U2625 (N_2625,N_1849,N_1868);
or U2626 (N_2626,N_1571,N_1880);
or U2627 (N_2627,N_2036,N_1548);
and U2628 (N_2628,N_2135,N_1588);
or U2629 (N_2629,N_1902,N_1855);
nor U2630 (N_2630,N_2076,N_1740);
and U2631 (N_2631,N_1803,N_1514);
and U2632 (N_2632,N_1542,N_2249);
or U2633 (N_2633,N_1950,N_2110);
nor U2634 (N_2634,N_2074,N_1951);
and U2635 (N_2635,N_1969,N_1585);
or U2636 (N_2636,N_1869,N_2161);
nor U2637 (N_2637,N_1570,N_1868);
and U2638 (N_2638,N_1852,N_2102);
and U2639 (N_2639,N_1535,N_2240);
nand U2640 (N_2640,N_2041,N_1563);
nor U2641 (N_2641,N_1905,N_2121);
or U2642 (N_2642,N_1802,N_1644);
nor U2643 (N_2643,N_1666,N_1511);
or U2644 (N_2644,N_2160,N_2090);
and U2645 (N_2645,N_1962,N_1722);
nor U2646 (N_2646,N_1562,N_1843);
or U2647 (N_2647,N_1562,N_1509);
nand U2648 (N_2648,N_1701,N_1771);
or U2649 (N_2649,N_2044,N_1741);
nor U2650 (N_2650,N_1769,N_1601);
or U2651 (N_2651,N_2030,N_2137);
and U2652 (N_2652,N_1951,N_1852);
or U2653 (N_2653,N_2002,N_1697);
nor U2654 (N_2654,N_2245,N_1763);
nor U2655 (N_2655,N_1634,N_1546);
and U2656 (N_2656,N_1950,N_1869);
and U2657 (N_2657,N_2020,N_1975);
and U2658 (N_2658,N_2102,N_2240);
nor U2659 (N_2659,N_1535,N_2086);
nor U2660 (N_2660,N_1678,N_1697);
nor U2661 (N_2661,N_1684,N_1815);
nor U2662 (N_2662,N_1892,N_2131);
or U2663 (N_2663,N_1763,N_2237);
nor U2664 (N_2664,N_1659,N_1883);
and U2665 (N_2665,N_2057,N_2088);
nor U2666 (N_2666,N_1614,N_2011);
and U2667 (N_2667,N_1791,N_1704);
nand U2668 (N_2668,N_2119,N_2015);
nand U2669 (N_2669,N_1978,N_1574);
nor U2670 (N_2670,N_1983,N_1639);
nor U2671 (N_2671,N_1939,N_2069);
nor U2672 (N_2672,N_1558,N_2054);
or U2673 (N_2673,N_1681,N_2203);
and U2674 (N_2674,N_2207,N_1697);
nand U2675 (N_2675,N_1597,N_1894);
nand U2676 (N_2676,N_1682,N_1859);
nor U2677 (N_2677,N_1790,N_1512);
nand U2678 (N_2678,N_1636,N_1983);
and U2679 (N_2679,N_2036,N_1946);
nor U2680 (N_2680,N_1618,N_1880);
nand U2681 (N_2681,N_1954,N_1751);
or U2682 (N_2682,N_2240,N_1642);
nand U2683 (N_2683,N_1768,N_2017);
and U2684 (N_2684,N_1985,N_1830);
nand U2685 (N_2685,N_1827,N_1524);
nand U2686 (N_2686,N_1500,N_1754);
nand U2687 (N_2687,N_1916,N_1858);
nor U2688 (N_2688,N_1863,N_1755);
nand U2689 (N_2689,N_2225,N_1756);
nand U2690 (N_2690,N_1748,N_1606);
and U2691 (N_2691,N_1864,N_1839);
and U2692 (N_2692,N_1714,N_2063);
nor U2693 (N_2693,N_1619,N_1834);
or U2694 (N_2694,N_1571,N_1831);
nand U2695 (N_2695,N_2104,N_1709);
and U2696 (N_2696,N_1999,N_2196);
or U2697 (N_2697,N_2107,N_1970);
nand U2698 (N_2698,N_1717,N_1867);
nor U2699 (N_2699,N_1525,N_1687);
nand U2700 (N_2700,N_2202,N_1815);
nor U2701 (N_2701,N_1509,N_2229);
nor U2702 (N_2702,N_1606,N_1753);
or U2703 (N_2703,N_1535,N_1839);
nand U2704 (N_2704,N_1589,N_2012);
nor U2705 (N_2705,N_1561,N_2017);
nand U2706 (N_2706,N_1992,N_2228);
and U2707 (N_2707,N_1718,N_1961);
nand U2708 (N_2708,N_1717,N_2102);
and U2709 (N_2709,N_1838,N_1969);
nor U2710 (N_2710,N_1575,N_2146);
or U2711 (N_2711,N_2197,N_1735);
or U2712 (N_2712,N_2237,N_1882);
or U2713 (N_2713,N_1696,N_2117);
or U2714 (N_2714,N_1901,N_1944);
or U2715 (N_2715,N_2072,N_2066);
nand U2716 (N_2716,N_1651,N_1945);
and U2717 (N_2717,N_1720,N_1515);
or U2718 (N_2718,N_2010,N_2101);
or U2719 (N_2719,N_2008,N_1937);
and U2720 (N_2720,N_1665,N_2246);
nor U2721 (N_2721,N_2143,N_2059);
and U2722 (N_2722,N_1586,N_1575);
nor U2723 (N_2723,N_1778,N_1598);
nor U2724 (N_2724,N_1909,N_1664);
and U2725 (N_2725,N_1675,N_2062);
nand U2726 (N_2726,N_2082,N_2135);
or U2727 (N_2727,N_1906,N_2104);
or U2728 (N_2728,N_1837,N_1588);
or U2729 (N_2729,N_2088,N_1897);
or U2730 (N_2730,N_1571,N_1617);
or U2731 (N_2731,N_1780,N_2221);
nor U2732 (N_2732,N_2199,N_1532);
and U2733 (N_2733,N_2030,N_2064);
nand U2734 (N_2734,N_2051,N_1742);
nor U2735 (N_2735,N_1920,N_1863);
or U2736 (N_2736,N_1625,N_1538);
nand U2737 (N_2737,N_1919,N_2239);
nor U2738 (N_2738,N_1561,N_1961);
nor U2739 (N_2739,N_1762,N_1989);
nand U2740 (N_2740,N_1748,N_2108);
nor U2741 (N_2741,N_2030,N_1747);
nand U2742 (N_2742,N_1996,N_1853);
or U2743 (N_2743,N_1945,N_1691);
nand U2744 (N_2744,N_1508,N_1636);
nor U2745 (N_2745,N_1724,N_1878);
or U2746 (N_2746,N_2241,N_1725);
or U2747 (N_2747,N_1633,N_1842);
and U2748 (N_2748,N_1624,N_1566);
and U2749 (N_2749,N_2099,N_2246);
and U2750 (N_2750,N_1976,N_2093);
nor U2751 (N_2751,N_1721,N_2242);
nor U2752 (N_2752,N_2132,N_1759);
and U2753 (N_2753,N_1867,N_1820);
nor U2754 (N_2754,N_1581,N_1740);
nand U2755 (N_2755,N_1783,N_2074);
nor U2756 (N_2756,N_1507,N_1862);
nor U2757 (N_2757,N_1579,N_2162);
nor U2758 (N_2758,N_1810,N_1797);
nor U2759 (N_2759,N_1763,N_1833);
and U2760 (N_2760,N_2047,N_1519);
or U2761 (N_2761,N_1913,N_1840);
or U2762 (N_2762,N_1900,N_2147);
nor U2763 (N_2763,N_1648,N_1588);
nor U2764 (N_2764,N_2097,N_1669);
nand U2765 (N_2765,N_1958,N_1832);
or U2766 (N_2766,N_2176,N_1759);
nor U2767 (N_2767,N_1691,N_1609);
nand U2768 (N_2768,N_1759,N_1790);
nor U2769 (N_2769,N_2248,N_1745);
or U2770 (N_2770,N_1849,N_1735);
nor U2771 (N_2771,N_1829,N_2243);
and U2772 (N_2772,N_2086,N_1542);
and U2773 (N_2773,N_2042,N_1602);
nand U2774 (N_2774,N_1953,N_2085);
nand U2775 (N_2775,N_2149,N_1728);
nor U2776 (N_2776,N_1630,N_2249);
and U2777 (N_2777,N_2079,N_1904);
and U2778 (N_2778,N_1969,N_1512);
and U2779 (N_2779,N_1890,N_1770);
nor U2780 (N_2780,N_1931,N_1724);
and U2781 (N_2781,N_2087,N_1641);
nand U2782 (N_2782,N_1876,N_2002);
or U2783 (N_2783,N_1572,N_1682);
and U2784 (N_2784,N_1679,N_1663);
nand U2785 (N_2785,N_1549,N_1778);
nand U2786 (N_2786,N_1578,N_1973);
nor U2787 (N_2787,N_2208,N_1567);
nand U2788 (N_2788,N_2017,N_1973);
or U2789 (N_2789,N_2012,N_2062);
and U2790 (N_2790,N_1722,N_1804);
nor U2791 (N_2791,N_2079,N_1513);
nand U2792 (N_2792,N_2089,N_1966);
nor U2793 (N_2793,N_1765,N_2120);
and U2794 (N_2794,N_1566,N_1710);
nor U2795 (N_2795,N_1904,N_1812);
or U2796 (N_2796,N_1607,N_1530);
and U2797 (N_2797,N_1585,N_1895);
nand U2798 (N_2798,N_1625,N_1976);
nand U2799 (N_2799,N_1737,N_1883);
or U2800 (N_2800,N_1876,N_2167);
and U2801 (N_2801,N_1776,N_2035);
nor U2802 (N_2802,N_2021,N_1874);
and U2803 (N_2803,N_1876,N_1596);
nand U2804 (N_2804,N_1686,N_1965);
nand U2805 (N_2805,N_1727,N_1742);
nand U2806 (N_2806,N_1967,N_1972);
nand U2807 (N_2807,N_1895,N_1902);
or U2808 (N_2808,N_1933,N_1793);
xor U2809 (N_2809,N_2059,N_1761);
or U2810 (N_2810,N_2160,N_1996);
or U2811 (N_2811,N_2066,N_1826);
nor U2812 (N_2812,N_2091,N_1951);
nor U2813 (N_2813,N_1739,N_1592);
nand U2814 (N_2814,N_1849,N_2157);
or U2815 (N_2815,N_1672,N_1795);
nand U2816 (N_2816,N_2028,N_1794);
and U2817 (N_2817,N_2223,N_1579);
or U2818 (N_2818,N_1957,N_1710);
nor U2819 (N_2819,N_1892,N_1957);
nor U2820 (N_2820,N_1619,N_1773);
and U2821 (N_2821,N_2160,N_2004);
nand U2822 (N_2822,N_2087,N_1587);
nand U2823 (N_2823,N_2073,N_1921);
nand U2824 (N_2824,N_1714,N_2154);
nor U2825 (N_2825,N_1596,N_1611);
nor U2826 (N_2826,N_2068,N_2038);
nor U2827 (N_2827,N_2078,N_1878);
or U2828 (N_2828,N_1725,N_1507);
nand U2829 (N_2829,N_2005,N_2173);
nor U2830 (N_2830,N_1988,N_1830);
nor U2831 (N_2831,N_1805,N_1721);
nor U2832 (N_2832,N_1910,N_1539);
nand U2833 (N_2833,N_1767,N_1747);
or U2834 (N_2834,N_1851,N_1903);
nor U2835 (N_2835,N_1714,N_1814);
and U2836 (N_2836,N_1534,N_1622);
nor U2837 (N_2837,N_1840,N_1636);
or U2838 (N_2838,N_2168,N_1871);
nor U2839 (N_2839,N_2036,N_2133);
or U2840 (N_2840,N_1769,N_2198);
and U2841 (N_2841,N_1922,N_1865);
nor U2842 (N_2842,N_2222,N_1864);
nor U2843 (N_2843,N_1862,N_1593);
nor U2844 (N_2844,N_1903,N_2173);
or U2845 (N_2845,N_1530,N_1813);
nand U2846 (N_2846,N_1679,N_1764);
and U2847 (N_2847,N_2099,N_1985);
nand U2848 (N_2848,N_2133,N_1627);
or U2849 (N_2849,N_1652,N_1845);
nand U2850 (N_2850,N_1567,N_1586);
and U2851 (N_2851,N_1545,N_2007);
nor U2852 (N_2852,N_1504,N_1626);
and U2853 (N_2853,N_1772,N_1717);
or U2854 (N_2854,N_2080,N_2014);
or U2855 (N_2855,N_2151,N_1996);
nor U2856 (N_2856,N_1940,N_1637);
nand U2857 (N_2857,N_2188,N_1678);
or U2858 (N_2858,N_1808,N_2199);
nand U2859 (N_2859,N_1632,N_2139);
xor U2860 (N_2860,N_1531,N_1984);
and U2861 (N_2861,N_2124,N_1756);
nand U2862 (N_2862,N_1769,N_1503);
nand U2863 (N_2863,N_1610,N_2032);
nor U2864 (N_2864,N_1851,N_1515);
nor U2865 (N_2865,N_2224,N_1779);
and U2866 (N_2866,N_2200,N_2070);
nor U2867 (N_2867,N_1835,N_1846);
nand U2868 (N_2868,N_2146,N_2064);
or U2869 (N_2869,N_1657,N_1857);
nand U2870 (N_2870,N_1928,N_2093);
nor U2871 (N_2871,N_2146,N_2231);
nand U2872 (N_2872,N_1756,N_1869);
nor U2873 (N_2873,N_2006,N_1736);
nor U2874 (N_2874,N_1973,N_1732);
nand U2875 (N_2875,N_1508,N_1510);
nand U2876 (N_2876,N_1864,N_1957);
nand U2877 (N_2877,N_1789,N_1567);
and U2878 (N_2878,N_1970,N_2102);
nand U2879 (N_2879,N_2081,N_1679);
nor U2880 (N_2880,N_2056,N_1540);
and U2881 (N_2881,N_1957,N_1735);
and U2882 (N_2882,N_2003,N_1616);
and U2883 (N_2883,N_2140,N_2099);
and U2884 (N_2884,N_1664,N_1735);
and U2885 (N_2885,N_1923,N_2060);
nand U2886 (N_2886,N_1522,N_1842);
nand U2887 (N_2887,N_2144,N_2054);
or U2888 (N_2888,N_1789,N_1809);
nand U2889 (N_2889,N_2146,N_1711);
or U2890 (N_2890,N_1867,N_1767);
or U2891 (N_2891,N_1970,N_2244);
and U2892 (N_2892,N_1734,N_1895);
nand U2893 (N_2893,N_1846,N_1518);
and U2894 (N_2894,N_1967,N_2203);
or U2895 (N_2895,N_1595,N_1719);
nand U2896 (N_2896,N_2092,N_2135);
or U2897 (N_2897,N_1622,N_1808);
or U2898 (N_2898,N_1719,N_1650);
nor U2899 (N_2899,N_1626,N_1660);
or U2900 (N_2900,N_1681,N_1860);
and U2901 (N_2901,N_2178,N_1741);
xnor U2902 (N_2902,N_1829,N_1653);
and U2903 (N_2903,N_1794,N_1973);
and U2904 (N_2904,N_1902,N_1949);
and U2905 (N_2905,N_1650,N_1528);
nand U2906 (N_2906,N_1540,N_1961);
and U2907 (N_2907,N_1677,N_1635);
nand U2908 (N_2908,N_2080,N_1659);
nor U2909 (N_2909,N_1656,N_1808);
nand U2910 (N_2910,N_1865,N_1955);
and U2911 (N_2911,N_1689,N_2092);
or U2912 (N_2912,N_1660,N_1667);
nand U2913 (N_2913,N_2147,N_1573);
nand U2914 (N_2914,N_2085,N_1826);
or U2915 (N_2915,N_1960,N_1535);
nand U2916 (N_2916,N_1707,N_2018);
nor U2917 (N_2917,N_1864,N_1824);
nand U2918 (N_2918,N_1858,N_1734);
and U2919 (N_2919,N_1975,N_2034);
nor U2920 (N_2920,N_1965,N_1626);
or U2921 (N_2921,N_1782,N_1874);
nor U2922 (N_2922,N_1837,N_1684);
and U2923 (N_2923,N_1901,N_2148);
and U2924 (N_2924,N_1976,N_1689);
nor U2925 (N_2925,N_2037,N_1755);
nor U2926 (N_2926,N_1823,N_1698);
nand U2927 (N_2927,N_1515,N_2231);
or U2928 (N_2928,N_2191,N_1516);
and U2929 (N_2929,N_1842,N_1514);
nand U2930 (N_2930,N_2027,N_1578);
or U2931 (N_2931,N_2164,N_1864);
or U2932 (N_2932,N_2079,N_1619);
and U2933 (N_2933,N_1742,N_1664);
or U2934 (N_2934,N_1600,N_2085);
and U2935 (N_2935,N_1587,N_1985);
nor U2936 (N_2936,N_2237,N_1779);
nor U2937 (N_2937,N_2122,N_1866);
nor U2938 (N_2938,N_1593,N_1806);
nor U2939 (N_2939,N_1800,N_1745);
nand U2940 (N_2940,N_1807,N_2247);
nand U2941 (N_2941,N_1588,N_1832);
nor U2942 (N_2942,N_1996,N_1630);
nor U2943 (N_2943,N_1885,N_1545);
nor U2944 (N_2944,N_2205,N_1516);
xnor U2945 (N_2945,N_1829,N_1662);
or U2946 (N_2946,N_2131,N_2194);
nor U2947 (N_2947,N_1993,N_2175);
or U2948 (N_2948,N_2228,N_2050);
nor U2949 (N_2949,N_1709,N_2186);
nor U2950 (N_2950,N_1609,N_2118);
and U2951 (N_2951,N_2051,N_1979);
nand U2952 (N_2952,N_2091,N_1694);
and U2953 (N_2953,N_2123,N_1664);
or U2954 (N_2954,N_1834,N_2206);
or U2955 (N_2955,N_1613,N_1636);
or U2956 (N_2956,N_2028,N_1808);
xnor U2957 (N_2957,N_1689,N_2166);
or U2958 (N_2958,N_1870,N_2163);
nand U2959 (N_2959,N_2156,N_2169);
and U2960 (N_2960,N_1601,N_1971);
nor U2961 (N_2961,N_2037,N_1670);
nand U2962 (N_2962,N_1573,N_1554);
nand U2963 (N_2963,N_2062,N_2134);
or U2964 (N_2964,N_1504,N_1981);
and U2965 (N_2965,N_1811,N_2244);
nor U2966 (N_2966,N_1876,N_1809);
nor U2967 (N_2967,N_1587,N_1811);
and U2968 (N_2968,N_1910,N_2216);
nor U2969 (N_2969,N_1970,N_1871);
and U2970 (N_2970,N_1536,N_2052);
nand U2971 (N_2971,N_1727,N_1540);
and U2972 (N_2972,N_1967,N_1514);
nor U2973 (N_2973,N_1674,N_1626);
and U2974 (N_2974,N_1588,N_1722);
and U2975 (N_2975,N_1953,N_1756);
and U2976 (N_2976,N_1631,N_2083);
nand U2977 (N_2977,N_2022,N_1720);
and U2978 (N_2978,N_2087,N_1747);
and U2979 (N_2979,N_1685,N_1985);
nand U2980 (N_2980,N_1879,N_2066);
or U2981 (N_2981,N_2132,N_2056);
nand U2982 (N_2982,N_1629,N_2033);
nand U2983 (N_2983,N_1628,N_2035);
and U2984 (N_2984,N_2077,N_1956);
and U2985 (N_2985,N_1641,N_1824);
nand U2986 (N_2986,N_1904,N_1653);
or U2987 (N_2987,N_1766,N_1617);
and U2988 (N_2988,N_2216,N_1999);
or U2989 (N_2989,N_1893,N_1670);
and U2990 (N_2990,N_2150,N_1582);
or U2991 (N_2991,N_1862,N_1826);
or U2992 (N_2992,N_1746,N_1625);
nand U2993 (N_2993,N_1730,N_1644);
nand U2994 (N_2994,N_1743,N_1528);
or U2995 (N_2995,N_1867,N_2039);
nor U2996 (N_2996,N_2007,N_2164);
nand U2997 (N_2997,N_1834,N_1714);
nand U2998 (N_2998,N_1909,N_1924);
and U2999 (N_2999,N_2121,N_2186);
and UO_0 (O_0,N_2494,N_2635);
and UO_1 (O_1,N_2641,N_2532);
and UO_2 (O_2,N_2385,N_2302);
and UO_3 (O_3,N_2814,N_2539);
nor UO_4 (O_4,N_2914,N_2825);
nand UO_5 (O_5,N_2732,N_2350);
and UO_6 (O_6,N_2605,N_2794);
or UO_7 (O_7,N_2256,N_2366);
nand UO_8 (O_8,N_2606,N_2254);
or UO_9 (O_9,N_2857,N_2855);
nand UO_10 (O_10,N_2511,N_2685);
nand UO_11 (O_11,N_2592,N_2772);
and UO_12 (O_12,N_2562,N_2341);
nand UO_13 (O_13,N_2580,N_2472);
nor UO_14 (O_14,N_2691,N_2623);
and UO_15 (O_15,N_2858,N_2423);
or UO_16 (O_16,N_2682,N_2823);
xnor UO_17 (O_17,N_2558,N_2339);
nand UO_18 (O_18,N_2513,N_2671);
or UO_19 (O_19,N_2953,N_2566);
nor UO_20 (O_20,N_2454,N_2841);
or UO_21 (O_21,N_2673,N_2431);
and UO_22 (O_22,N_2518,N_2743);
nor UO_23 (O_23,N_2546,N_2901);
or UO_24 (O_24,N_2946,N_2838);
or UO_25 (O_25,N_2676,N_2443);
nand UO_26 (O_26,N_2972,N_2775);
nand UO_27 (O_27,N_2528,N_2644);
and UO_28 (O_28,N_2432,N_2464);
nor UO_29 (O_29,N_2418,N_2403);
and UO_30 (O_30,N_2709,N_2821);
and UO_31 (O_31,N_2404,N_2527);
nand UO_32 (O_32,N_2614,N_2813);
nor UO_33 (O_33,N_2983,N_2738);
and UO_34 (O_34,N_2899,N_2979);
or UO_35 (O_35,N_2425,N_2756);
nor UO_36 (O_36,N_2663,N_2291);
or UO_37 (O_37,N_2474,N_2834);
nand UO_38 (O_38,N_2283,N_2752);
nor UO_39 (O_39,N_2519,N_2434);
nor UO_40 (O_40,N_2694,N_2278);
nor UO_41 (O_41,N_2660,N_2701);
or UO_42 (O_42,N_2757,N_2289);
nand UO_43 (O_43,N_2295,N_2723);
or UO_44 (O_44,N_2711,N_2894);
and UO_45 (O_45,N_2255,N_2553);
nand UO_46 (O_46,N_2864,N_2311);
and UO_47 (O_47,N_2355,N_2479);
nor UO_48 (O_48,N_2905,N_2521);
nor UO_49 (O_49,N_2465,N_2356);
or UO_50 (O_50,N_2453,N_2508);
nand UO_51 (O_51,N_2651,N_2514);
nor UO_52 (O_52,N_2570,N_2380);
and UO_53 (O_53,N_2804,N_2360);
nand UO_54 (O_54,N_2702,N_2354);
and UO_55 (O_55,N_2344,N_2374);
and UO_56 (O_56,N_2578,N_2446);
nand UO_57 (O_57,N_2524,N_2799);
nand UO_58 (O_58,N_2634,N_2590);
nor UO_59 (O_59,N_2357,N_2611);
nor UO_60 (O_60,N_2338,N_2603);
nor UO_61 (O_61,N_2674,N_2268);
and UO_62 (O_62,N_2891,N_2954);
nor UO_63 (O_63,N_2293,N_2964);
and UO_64 (O_64,N_2797,N_2997);
nor UO_65 (O_65,N_2492,N_2907);
nand UO_66 (O_66,N_2428,N_2800);
or UO_67 (O_67,N_2913,N_2776);
nand UO_68 (O_68,N_2625,N_2333);
or UO_69 (O_69,N_2657,N_2897);
nand UO_70 (O_70,N_2792,N_2369);
and UO_71 (O_71,N_2787,N_2725);
or UO_72 (O_72,N_2822,N_2739);
nor UO_73 (O_73,N_2544,N_2309);
nor UO_74 (O_74,N_2928,N_2378);
nand UO_75 (O_75,N_2462,N_2895);
or UO_76 (O_76,N_2960,N_2535);
nor UO_77 (O_77,N_2741,N_2285);
nor UO_78 (O_78,N_2370,N_2517);
nor UO_79 (O_79,N_2693,N_2912);
nand UO_80 (O_80,N_2733,N_2627);
and UO_81 (O_81,N_2990,N_2999);
or UO_82 (O_82,N_2873,N_2643);
and UO_83 (O_83,N_2729,N_2368);
and UO_84 (O_84,N_2600,N_2461);
or UO_85 (O_85,N_2300,N_2444);
nor UO_86 (O_86,N_2515,N_2886);
or UO_87 (O_87,N_2542,N_2654);
and UO_88 (O_88,N_2639,N_2933);
and UO_89 (O_89,N_2351,N_2932);
and UO_90 (O_90,N_2778,N_2640);
and UO_91 (O_91,N_2966,N_2384);
nor UO_92 (O_92,N_2938,N_2690);
nand UO_93 (O_93,N_2407,N_2261);
or UO_94 (O_94,N_2576,N_2608);
nand UO_95 (O_95,N_2317,N_2981);
or UO_96 (O_96,N_2998,N_2318);
nor UO_97 (O_97,N_2885,N_2442);
nor UO_98 (O_98,N_2844,N_2664);
and UO_99 (O_99,N_2531,N_2398);
and UO_100 (O_100,N_2985,N_2489);
nand UO_101 (O_101,N_2386,N_2719);
and UO_102 (O_102,N_2807,N_2468);
or UO_103 (O_103,N_2439,N_2417);
nand UO_104 (O_104,N_2884,N_2696);
nor UO_105 (O_105,N_2632,N_2727);
or UO_106 (O_106,N_2502,N_2324);
nand UO_107 (O_107,N_2896,N_2745);
nand UO_108 (O_108,N_2935,N_2506);
or UO_109 (O_109,N_2780,N_2371);
or UO_110 (O_110,N_2348,N_2383);
nor UO_111 (O_111,N_2267,N_2722);
nor UO_112 (O_112,N_2862,N_2301);
nand UO_113 (O_113,N_2326,N_2548);
nor UO_114 (O_114,N_2924,N_2342);
nor UO_115 (O_115,N_2646,N_2626);
and UO_116 (O_116,N_2617,N_2781);
and UO_117 (O_117,N_2773,N_2850);
nand UO_118 (O_118,N_2304,N_2771);
nand UO_119 (O_119,N_2397,N_2853);
or UO_120 (O_120,N_2943,N_2993);
or UO_121 (O_121,N_2496,N_2543);
and UO_122 (O_122,N_2422,N_2868);
and UO_123 (O_123,N_2828,N_2467);
nand UO_124 (O_124,N_2699,N_2487);
or UO_125 (O_125,N_2426,N_2598);
nand UO_126 (O_126,N_2959,N_2835);
and UO_127 (O_127,N_2609,N_2929);
nand UO_128 (O_128,N_2367,N_2485);
nor UO_129 (O_129,N_2604,N_2796);
or UO_130 (O_130,N_2402,N_2433);
nor UO_131 (O_131,N_2840,N_2497);
or UO_132 (O_132,N_2883,N_2991);
nand UO_133 (O_133,N_2619,N_2642);
and UO_134 (O_134,N_2949,N_2483);
and UO_135 (O_135,N_2675,N_2286);
or UO_136 (O_136,N_2656,N_2353);
or UO_137 (O_137,N_2320,N_2806);
or UO_138 (O_138,N_2591,N_2334);
and UO_139 (O_139,N_2303,N_2538);
nand UO_140 (O_140,N_2473,N_2662);
and UO_141 (O_141,N_2345,N_2970);
nor UO_142 (O_142,N_2500,N_2533);
or UO_143 (O_143,N_2659,N_2887);
or UO_144 (O_144,N_2352,N_2541);
and UO_145 (O_145,N_2365,N_2961);
nor UO_146 (O_146,N_2389,N_2612);
and UO_147 (O_147,N_2764,N_2495);
and UO_148 (O_148,N_2451,N_2584);
and UO_149 (O_149,N_2452,N_2670);
and UO_150 (O_150,N_2849,N_2572);
nand UO_151 (O_151,N_2388,N_2296);
nand UO_152 (O_152,N_2534,N_2455);
nor UO_153 (O_153,N_2692,N_2892);
or UO_154 (O_154,N_2652,N_2755);
nor UO_155 (O_155,N_2810,N_2842);
or UO_156 (O_156,N_2504,N_2890);
nand UO_157 (O_157,N_2488,N_2965);
or UO_158 (O_158,N_2758,N_2681);
and UO_159 (O_159,N_2536,N_2280);
or UO_160 (O_160,N_2613,N_2951);
and UO_161 (O_161,N_2471,N_2337);
and UO_162 (O_162,N_2686,N_2866);
or UO_163 (O_163,N_2688,N_2715);
and UO_164 (O_164,N_2375,N_2327);
and UO_165 (O_165,N_2503,N_2974);
or UO_166 (O_166,N_2395,N_2730);
nand UO_167 (O_167,N_2331,N_2622);
or UO_168 (O_168,N_2759,N_2499);
nand UO_169 (O_169,N_2941,N_2530);
and UO_170 (O_170,N_2836,N_2358);
and UO_171 (O_171,N_2429,N_2271);
or UO_172 (O_172,N_2879,N_2266);
and UO_173 (O_173,N_2803,N_2273);
and UO_174 (O_174,N_2955,N_2768);
nor UO_175 (O_175,N_2469,N_2491);
or UO_176 (O_176,N_2290,N_2336);
nand UO_177 (O_177,N_2708,N_2560);
nand UO_178 (O_178,N_2852,N_2948);
nor UO_179 (O_179,N_2512,N_2881);
nand UO_180 (O_180,N_2843,N_2315);
nor UO_181 (O_181,N_2921,N_2270);
or UO_182 (O_182,N_2870,N_2906);
and UO_183 (O_183,N_2585,N_2409);
nor UO_184 (O_184,N_2364,N_2889);
and UO_185 (O_185,N_2459,N_2615);
or UO_186 (O_186,N_2437,N_2861);
or UO_187 (O_187,N_2550,N_2616);
nor UO_188 (O_188,N_2340,N_2299);
and UO_189 (O_189,N_2769,N_2482);
nor UO_190 (O_190,N_2274,N_2737);
or UO_191 (O_191,N_2904,N_2281);
and UO_192 (O_192,N_2902,N_2963);
nand UO_193 (O_193,N_2330,N_2820);
nand UO_194 (O_194,N_2687,N_2925);
and UO_195 (O_195,N_2684,N_2636);
or UO_196 (O_196,N_2783,N_2677);
nor UO_197 (O_197,N_2851,N_2556);
nor UO_198 (O_198,N_2449,N_2396);
nor UO_199 (O_199,N_2854,N_2440);
or UO_200 (O_200,N_2728,N_2798);
nor UO_201 (O_201,N_2791,N_2582);
nand UO_202 (O_202,N_2313,N_2975);
nor UO_203 (O_203,N_2329,N_2490);
nand UO_204 (O_204,N_2774,N_2312);
nor UO_205 (O_205,N_2265,N_2287);
nor UO_206 (O_206,N_2765,N_2874);
nor UO_207 (O_207,N_2391,N_2420);
nor UO_208 (O_208,N_2856,N_2706);
or UO_209 (O_209,N_2577,N_2898);
or UO_210 (O_210,N_2478,N_2569);
nor UO_211 (O_211,N_2481,N_2470);
nand UO_212 (O_212,N_2638,N_2314);
nor UO_213 (O_213,N_2272,N_2379);
or UO_214 (O_214,N_2475,N_2363);
or UO_215 (O_215,N_2373,N_2698);
nand UO_216 (O_216,N_2305,N_2766);
nor UO_217 (O_217,N_2669,N_2666);
nand UO_218 (O_218,N_2310,N_2911);
nand UO_219 (O_219,N_2631,N_2450);
or UO_220 (O_220,N_2917,N_2588);
or UO_221 (O_221,N_2689,N_2316);
nand UO_222 (O_222,N_2498,N_2815);
and UO_223 (O_223,N_2658,N_2647);
nor UO_224 (O_224,N_2322,N_2257);
and UO_225 (O_225,N_2968,N_2996);
and UO_226 (O_226,N_2387,N_2760);
nor UO_227 (O_227,N_2637,N_2980);
nor UO_228 (O_228,N_2973,N_2476);
nand UO_229 (O_229,N_2667,N_2571);
or UO_230 (O_230,N_2650,N_2845);
or UO_231 (O_231,N_2258,N_2847);
nand UO_232 (O_232,N_2731,N_2816);
nor UO_233 (O_233,N_2335,N_2493);
nor UO_234 (O_234,N_2712,N_2665);
and UO_235 (O_235,N_2726,N_2922);
and UO_236 (O_236,N_2819,N_2882);
nor UO_237 (O_237,N_2522,N_2962);
nor UO_238 (O_238,N_2995,N_2441);
or UO_239 (O_239,N_2749,N_2695);
or UO_240 (O_240,N_2307,N_2332);
nor UO_241 (O_241,N_2872,N_2567);
nand UO_242 (O_242,N_2435,N_2831);
nor UO_243 (O_243,N_2923,N_2957);
or UO_244 (O_244,N_2782,N_2501);
or UO_245 (O_245,N_2477,N_2865);
or UO_246 (O_246,N_2940,N_2926);
nor UO_247 (O_247,N_2523,N_2648);
nand UO_248 (O_248,N_2833,N_2460);
nor UO_249 (O_249,N_2977,N_2735);
and UO_250 (O_250,N_2408,N_2786);
and UO_251 (O_251,N_2325,N_2292);
and UO_252 (O_252,N_2628,N_2958);
nor UO_253 (O_253,N_2565,N_2372);
or UO_254 (O_254,N_2262,N_2457);
or UO_255 (O_255,N_2545,N_2581);
or UO_256 (O_256,N_2406,N_2555);
nor UO_257 (O_257,N_2875,N_2392);
nand UO_258 (O_258,N_2599,N_2405);
nor UO_259 (O_259,N_2306,N_2829);
nand UO_260 (O_260,N_2805,N_2621);
or UO_261 (O_261,N_2716,N_2401);
and UO_262 (O_262,N_2509,N_2377);
nor UO_263 (O_263,N_2410,N_2826);
nor UO_264 (O_264,N_2987,N_2763);
nor UO_265 (O_265,N_2448,N_2414);
and UO_266 (O_266,N_2575,N_2264);
nand UO_267 (O_267,N_2263,N_2863);
nor UO_268 (O_268,N_2624,N_2947);
or UO_269 (O_269,N_2607,N_2994);
and UO_270 (O_270,N_2678,N_2988);
nand UO_271 (O_271,N_2789,N_2679);
nand UO_272 (O_272,N_2750,N_2547);
and UO_273 (O_273,N_2610,N_2579);
or UO_274 (O_274,N_2554,N_2910);
nand UO_275 (O_275,N_2564,N_2986);
nor UO_276 (O_276,N_2936,N_2359);
nand UO_277 (O_277,N_2746,N_2930);
and UO_278 (O_278,N_2620,N_2721);
nor UO_279 (O_279,N_2552,N_2419);
or UO_280 (O_280,N_2458,N_2507);
or UO_281 (O_281,N_2880,N_2276);
and UO_282 (O_282,N_2400,N_2394);
and UO_283 (O_283,N_2253,N_2574);
nor UO_284 (O_284,N_2871,N_2812);
or UO_285 (O_285,N_2415,N_2744);
nand UO_286 (O_286,N_2297,N_2393);
nor UO_287 (O_287,N_2633,N_2793);
nor UO_288 (O_288,N_2361,N_2416);
nand UO_289 (O_289,N_2978,N_2480);
and UO_290 (O_290,N_2802,N_2298);
nor UO_291 (O_291,N_2992,N_2937);
and UO_292 (O_292,N_2790,N_2779);
xor UO_293 (O_293,N_2645,N_2630);
xnor UO_294 (O_294,N_2308,N_2767);
nor UO_295 (O_295,N_2927,N_2751);
nor UO_296 (O_296,N_2944,N_2346);
or UO_297 (O_297,N_2700,N_2284);
nand UO_298 (O_298,N_2718,N_2279);
nand UO_299 (O_299,N_2893,N_2436);
nand UO_300 (O_300,N_2427,N_2390);
nor UO_301 (O_301,N_2655,N_2668);
or UO_302 (O_302,N_2918,N_2411);
nand UO_303 (O_303,N_2413,N_2876);
nand UO_304 (O_304,N_2595,N_2589);
or UO_305 (O_305,N_2587,N_2740);
nand UO_306 (O_306,N_2559,N_2707);
nor UO_307 (O_307,N_2549,N_2399);
nand UO_308 (O_308,N_2754,N_2969);
nand UO_309 (O_309,N_2717,N_2683);
and UO_310 (O_310,N_2529,N_2830);
and UO_311 (O_311,N_2971,N_2586);
nor UO_312 (O_312,N_2456,N_2260);
nor UO_313 (O_313,N_2724,N_2252);
or UO_314 (O_314,N_2869,N_2915);
and UO_315 (O_315,N_2382,N_2596);
nand UO_316 (O_316,N_2801,N_2878);
and UO_317 (O_317,N_2505,N_2563);
and UO_318 (O_318,N_2704,N_2321);
or UO_319 (O_319,N_2967,N_2900);
nor UO_320 (O_320,N_2705,N_2447);
and UO_321 (O_321,N_2710,N_2984);
nand UO_322 (O_322,N_2463,N_2583);
and UO_323 (O_323,N_2445,N_2788);
nand UO_324 (O_324,N_2747,N_2777);
xnor UO_325 (O_325,N_2323,N_2294);
or UO_326 (O_326,N_2976,N_2680);
nor UO_327 (O_327,N_2661,N_2343);
or UO_328 (O_328,N_2839,N_2697);
nor UO_329 (O_329,N_2525,N_2275);
or UO_330 (O_330,N_2618,N_2277);
nand UO_331 (O_331,N_2561,N_2832);
nand UO_332 (O_332,N_2486,N_2795);
or UO_333 (O_333,N_2817,N_2753);
or UO_334 (O_334,N_2860,N_2282);
nor UO_335 (O_335,N_2466,N_2848);
and UO_336 (O_336,N_2908,N_2748);
nand UO_337 (O_337,N_2557,N_2376);
and UO_338 (O_338,N_2424,N_2288);
nand UO_339 (O_339,N_2438,N_2672);
nor UO_340 (O_340,N_2594,N_2713);
nor UO_341 (O_341,N_2808,N_2945);
nand UO_342 (O_342,N_2846,N_2362);
and UO_343 (O_343,N_2597,N_2430);
and UO_344 (O_344,N_2877,N_2785);
nor UO_345 (O_345,N_2837,N_2734);
nand UO_346 (O_346,N_2888,N_2516);
or UO_347 (O_347,N_2982,N_2601);
and UO_348 (O_348,N_2931,N_2950);
nand UO_349 (O_349,N_2939,N_2349);
and UO_350 (O_350,N_2942,N_2784);
nand UO_351 (O_351,N_2381,N_2551);
nand UO_352 (O_352,N_2250,N_2934);
and UO_353 (O_353,N_2269,N_2867);
or UO_354 (O_354,N_2703,N_2919);
and UO_355 (O_355,N_2720,N_2649);
and UO_356 (O_356,N_2770,N_2818);
nor UO_357 (O_357,N_2811,N_2568);
or UO_358 (O_358,N_2920,N_2573);
or UO_359 (O_359,N_2809,N_2526);
nand UO_360 (O_360,N_2510,N_2602);
nor UO_361 (O_361,N_2714,N_2761);
and UO_362 (O_362,N_2903,N_2956);
nand UO_363 (O_363,N_2421,N_2251);
nor UO_364 (O_364,N_2520,N_2827);
or UO_365 (O_365,N_2629,N_2909);
or UO_366 (O_366,N_2593,N_2319);
nor UO_367 (O_367,N_2537,N_2762);
and UO_368 (O_368,N_2328,N_2484);
nand UO_369 (O_369,N_2259,N_2347);
nand UO_370 (O_370,N_2653,N_2916);
nor UO_371 (O_371,N_2412,N_2989);
and UO_372 (O_372,N_2824,N_2736);
nor UO_373 (O_373,N_2859,N_2952);
nand UO_374 (O_374,N_2540,N_2742);
or UO_375 (O_375,N_2251,N_2366);
and UO_376 (O_376,N_2587,N_2463);
nor UO_377 (O_377,N_2632,N_2856);
or UO_378 (O_378,N_2559,N_2742);
and UO_379 (O_379,N_2559,N_2364);
and UO_380 (O_380,N_2588,N_2923);
and UO_381 (O_381,N_2881,N_2653);
and UO_382 (O_382,N_2532,N_2573);
nor UO_383 (O_383,N_2902,N_2753);
nor UO_384 (O_384,N_2550,N_2482);
nor UO_385 (O_385,N_2717,N_2690);
nand UO_386 (O_386,N_2536,N_2748);
nor UO_387 (O_387,N_2548,N_2912);
or UO_388 (O_388,N_2981,N_2938);
nor UO_389 (O_389,N_2975,N_2691);
nand UO_390 (O_390,N_2260,N_2429);
nand UO_391 (O_391,N_2464,N_2951);
nor UO_392 (O_392,N_2885,N_2651);
and UO_393 (O_393,N_2339,N_2938);
nand UO_394 (O_394,N_2838,N_2817);
nor UO_395 (O_395,N_2455,N_2526);
or UO_396 (O_396,N_2784,N_2440);
nand UO_397 (O_397,N_2658,N_2354);
and UO_398 (O_398,N_2530,N_2355);
nor UO_399 (O_399,N_2612,N_2555);
or UO_400 (O_400,N_2908,N_2358);
or UO_401 (O_401,N_2503,N_2988);
nand UO_402 (O_402,N_2999,N_2412);
or UO_403 (O_403,N_2622,N_2956);
and UO_404 (O_404,N_2556,N_2961);
and UO_405 (O_405,N_2928,N_2755);
or UO_406 (O_406,N_2658,N_2447);
nand UO_407 (O_407,N_2791,N_2905);
nand UO_408 (O_408,N_2758,N_2511);
or UO_409 (O_409,N_2773,N_2716);
nor UO_410 (O_410,N_2813,N_2525);
and UO_411 (O_411,N_2404,N_2942);
nand UO_412 (O_412,N_2951,N_2967);
or UO_413 (O_413,N_2739,N_2471);
and UO_414 (O_414,N_2333,N_2763);
and UO_415 (O_415,N_2844,N_2715);
and UO_416 (O_416,N_2834,N_2534);
nor UO_417 (O_417,N_2611,N_2680);
nor UO_418 (O_418,N_2816,N_2842);
nor UO_419 (O_419,N_2667,N_2678);
nand UO_420 (O_420,N_2314,N_2336);
nand UO_421 (O_421,N_2437,N_2825);
nand UO_422 (O_422,N_2518,N_2398);
nor UO_423 (O_423,N_2643,N_2650);
nand UO_424 (O_424,N_2920,N_2251);
or UO_425 (O_425,N_2268,N_2692);
nor UO_426 (O_426,N_2957,N_2782);
and UO_427 (O_427,N_2573,N_2629);
nor UO_428 (O_428,N_2633,N_2592);
or UO_429 (O_429,N_2348,N_2632);
nand UO_430 (O_430,N_2316,N_2573);
or UO_431 (O_431,N_2958,N_2287);
nor UO_432 (O_432,N_2715,N_2890);
and UO_433 (O_433,N_2814,N_2998);
nor UO_434 (O_434,N_2680,N_2506);
nor UO_435 (O_435,N_2365,N_2302);
or UO_436 (O_436,N_2537,N_2506);
and UO_437 (O_437,N_2688,N_2851);
nand UO_438 (O_438,N_2984,N_2616);
and UO_439 (O_439,N_2614,N_2536);
nor UO_440 (O_440,N_2715,N_2960);
or UO_441 (O_441,N_2907,N_2937);
nor UO_442 (O_442,N_2858,N_2416);
nor UO_443 (O_443,N_2573,N_2624);
nor UO_444 (O_444,N_2840,N_2514);
or UO_445 (O_445,N_2920,N_2502);
and UO_446 (O_446,N_2651,N_2761);
nand UO_447 (O_447,N_2641,N_2908);
and UO_448 (O_448,N_2764,N_2462);
or UO_449 (O_449,N_2855,N_2260);
or UO_450 (O_450,N_2338,N_2898);
and UO_451 (O_451,N_2432,N_2655);
and UO_452 (O_452,N_2784,N_2992);
and UO_453 (O_453,N_2486,N_2472);
xnor UO_454 (O_454,N_2703,N_2907);
nand UO_455 (O_455,N_2799,N_2378);
and UO_456 (O_456,N_2558,N_2801);
or UO_457 (O_457,N_2698,N_2992);
nor UO_458 (O_458,N_2549,N_2307);
nand UO_459 (O_459,N_2313,N_2445);
or UO_460 (O_460,N_2376,N_2942);
nor UO_461 (O_461,N_2360,N_2673);
or UO_462 (O_462,N_2642,N_2279);
or UO_463 (O_463,N_2802,N_2516);
and UO_464 (O_464,N_2402,N_2703);
nor UO_465 (O_465,N_2460,N_2848);
nor UO_466 (O_466,N_2268,N_2509);
nand UO_467 (O_467,N_2321,N_2850);
or UO_468 (O_468,N_2622,N_2964);
nor UO_469 (O_469,N_2834,N_2772);
and UO_470 (O_470,N_2985,N_2574);
nand UO_471 (O_471,N_2731,N_2909);
or UO_472 (O_472,N_2464,N_2543);
or UO_473 (O_473,N_2858,N_2498);
nand UO_474 (O_474,N_2680,N_2668);
nand UO_475 (O_475,N_2585,N_2484);
or UO_476 (O_476,N_2470,N_2999);
and UO_477 (O_477,N_2492,N_2727);
or UO_478 (O_478,N_2537,N_2656);
nor UO_479 (O_479,N_2882,N_2770);
and UO_480 (O_480,N_2414,N_2936);
nor UO_481 (O_481,N_2301,N_2807);
nor UO_482 (O_482,N_2681,N_2349);
nand UO_483 (O_483,N_2677,N_2992);
nand UO_484 (O_484,N_2311,N_2315);
and UO_485 (O_485,N_2874,N_2539);
or UO_486 (O_486,N_2629,N_2520);
nor UO_487 (O_487,N_2532,N_2607);
or UO_488 (O_488,N_2322,N_2758);
nand UO_489 (O_489,N_2574,N_2765);
and UO_490 (O_490,N_2545,N_2913);
nand UO_491 (O_491,N_2515,N_2931);
or UO_492 (O_492,N_2907,N_2770);
or UO_493 (O_493,N_2815,N_2626);
nand UO_494 (O_494,N_2330,N_2912);
and UO_495 (O_495,N_2399,N_2788);
and UO_496 (O_496,N_2675,N_2250);
nor UO_497 (O_497,N_2858,N_2310);
or UO_498 (O_498,N_2507,N_2947);
nand UO_499 (O_499,N_2649,N_2794);
endmodule