module basic_2000_20000_2500_10_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
xor U0 (N_0,In_1487,In_165);
and U1 (N_1,In_436,In_1895);
and U2 (N_2,In_1491,In_134);
or U3 (N_3,In_1857,In_290);
nor U4 (N_4,In_698,In_60);
xnor U5 (N_5,In_1434,In_250);
and U6 (N_6,In_1409,In_992);
and U7 (N_7,In_202,In_805);
nor U8 (N_8,In_1072,In_937);
nand U9 (N_9,In_509,In_1464);
nor U10 (N_10,In_1831,In_1360);
or U11 (N_11,In_350,In_489);
xnor U12 (N_12,In_1701,In_961);
xor U13 (N_13,In_652,In_1397);
nand U14 (N_14,In_367,In_1079);
xor U15 (N_15,In_731,In_1158);
or U16 (N_16,In_1558,In_575);
and U17 (N_17,In_1728,In_1340);
xnor U18 (N_18,In_856,In_671);
nand U19 (N_19,In_889,In_829);
and U20 (N_20,In_708,In_982);
nor U21 (N_21,In_1297,In_98);
and U22 (N_22,In_1383,In_71);
or U23 (N_23,In_905,In_1544);
xnor U24 (N_24,In_726,In_1919);
and U25 (N_25,In_611,In_1962);
xnor U26 (N_26,In_1458,In_1386);
or U27 (N_27,In_1234,In_1592);
xor U28 (N_28,In_1042,In_1039);
nand U29 (N_29,In_1175,In_1308);
and U30 (N_30,In_1553,In_542);
or U31 (N_31,In_954,In_1767);
xor U32 (N_32,In_125,In_818);
xor U33 (N_33,In_1226,In_345);
or U34 (N_34,In_395,In_128);
or U35 (N_35,In_841,In_942);
xor U36 (N_36,In_577,In_162);
nand U37 (N_37,In_1820,In_298);
xor U38 (N_38,In_300,In_623);
nand U39 (N_39,In_1684,In_490);
or U40 (N_40,In_810,In_933);
xor U41 (N_41,In_464,In_46);
nand U42 (N_42,In_1631,In_392);
or U43 (N_43,In_636,In_1860);
nand U44 (N_44,In_221,In_585);
nand U45 (N_45,In_494,In_1939);
and U46 (N_46,In_1247,In_146);
xnor U47 (N_47,In_1817,In_424);
nor U48 (N_48,In_772,In_349);
xor U49 (N_49,In_1431,In_723);
nand U50 (N_50,In_1593,In_292);
and U51 (N_51,In_1290,In_1634);
and U52 (N_52,In_958,In_439);
xor U53 (N_53,In_1059,In_1452);
nor U54 (N_54,In_1578,In_285);
or U55 (N_55,In_1594,In_348);
xor U56 (N_56,In_709,In_1913);
and U57 (N_57,In_1187,In_1012);
or U58 (N_58,In_1246,In_18);
nand U59 (N_59,In_56,In_273);
nor U60 (N_60,In_133,In_1688);
and U61 (N_61,In_1752,In_1912);
nand U62 (N_62,In_38,In_1848);
or U63 (N_63,In_84,In_352);
or U64 (N_64,In_1643,In_507);
xor U65 (N_65,In_520,In_983);
or U66 (N_66,In_676,In_1148);
nor U67 (N_67,In_1310,In_1950);
nor U68 (N_68,In_1502,In_76);
xor U69 (N_69,In_1797,In_1610);
or U70 (N_70,In_1024,In_602);
or U71 (N_71,In_789,In_1471);
or U72 (N_72,In_160,In_242);
xnor U73 (N_73,In_1103,In_540);
and U74 (N_74,In_1959,In_1743);
nand U75 (N_75,In_287,In_1614);
and U76 (N_76,In_1045,In_1987);
nand U77 (N_77,In_1798,In_1381);
nor U78 (N_78,In_1724,In_956);
and U79 (N_79,In_1160,In_1238);
or U80 (N_80,In_884,In_231);
and U81 (N_81,In_1077,In_337);
or U82 (N_82,In_1055,In_206);
nor U83 (N_83,In_262,In_1010);
nand U84 (N_84,In_478,In_776);
or U85 (N_85,In_307,In_305);
xnor U86 (N_86,In_814,In_747);
nand U87 (N_87,In_1164,In_1653);
or U88 (N_88,In_842,In_1616);
nor U89 (N_89,In_695,In_1730);
nand U90 (N_90,In_1140,In_1672);
nand U91 (N_91,In_283,In_1147);
nor U92 (N_92,In_846,In_249);
nor U93 (N_93,In_1493,In_0);
nor U94 (N_94,In_1359,In_386);
nor U95 (N_95,In_852,In_50);
nand U96 (N_96,In_208,In_1159);
nand U97 (N_97,In_1395,In_265);
nand U98 (N_98,In_1889,In_1056);
and U99 (N_99,In_529,In_1398);
and U100 (N_100,In_931,In_1648);
or U101 (N_101,In_1851,In_631);
nand U102 (N_102,In_421,In_241);
xnor U103 (N_103,In_936,In_573);
xor U104 (N_104,In_83,In_826);
nor U105 (N_105,In_1520,In_645);
nand U106 (N_106,In_39,In_278);
or U107 (N_107,In_1030,In_123);
xnor U108 (N_108,In_666,In_1532);
and U109 (N_109,In_1036,In_1348);
nor U110 (N_110,In_1833,In_1920);
xor U111 (N_111,In_209,In_1715);
nor U112 (N_112,In_1953,In_1215);
or U113 (N_113,In_1985,In_739);
and U114 (N_114,In_322,In_1534);
nand U115 (N_115,In_391,In_899);
and U116 (N_116,In_1506,In_354);
nor U117 (N_117,In_190,In_1572);
or U118 (N_118,In_1830,In_1071);
and U119 (N_119,In_948,In_416);
nor U120 (N_120,In_1457,In_1037);
xor U121 (N_121,In_1515,In_1638);
and U122 (N_122,In_1760,In_748);
nor U123 (N_123,In_728,In_1635);
nor U124 (N_124,In_1043,In_1890);
nor U125 (N_125,In_1976,In_622);
and U126 (N_126,In_959,In_1120);
xnor U127 (N_127,In_677,In_336);
nor U128 (N_128,In_1839,In_1863);
nand U129 (N_129,In_245,In_1067);
xor U130 (N_130,In_1352,In_106);
nor U131 (N_131,In_735,In_1891);
or U132 (N_132,In_407,In_1300);
nor U133 (N_133,In_661,In_444);
and U134 (N_134,In_216,In_1086);
xnor U135 (N_135,In_1664,In_77);
nor U136 (N_136,In_1883,In_574);
xor U137 (N_137,In_660,In_1733);
nor U138 (N_138,In_1134,In_702);
xor U139 (N_139,In_1231,In_1549);
and U140 (N_140,In_343,In_627);
xor U141 (N_141,In_1218,In_1963);
nand U142 (N_142,In_1429,In_1837);
nand U143 (N_143,In_1214,In_868);
nand U144 (N_144,In_1362,In_442);
and U145 (N_145,In_1015,In_1796);
nand U146 (N_146,In_503,In_1321);
nor U147 (N_147,In_299,In_1034);
and U148 (N_148,In_451,In_1825);
and U149 (N_149,In_239,In_733);
nand U150 (N_150,In_1898,In_806);
nand U151 (N_151,In_1979,In_586);
and U152 (N_152,In_819,In_272);
or U153 (N_153,In_893,In_16);
or U154 (N_154,In_374,In_515);
and U155 (N_155,In_502,In_263);
xnor U156 (N_156,In_475,In_716);
xnor U157 (N_157,In_560,In_775);
nor U158 (N_158,In_1689,In_521);
xor U159 (N_159,In_1580,In_1991);
or U160 (N_160,In_519,In_820);
nand U161 (N_161,In_617,In_719);
nor U162 (N_162,In_154,In_1318);
xnor U163 (N_163,In_1675,In_1106);
nor U164 (N_164,In_1367,In_1233);
nand U165 (N_165,In_2,In_1376);
or U166 (N_166,In_1373,In_1249);
and U167 (N_167,In_1566,In_67);
nand U168 (N_168,In_222,In_1834);
and U169 (N_169,In_1986,In_1776);
nand U170 (N_170,In_1972,In_981);
or U171 (N_171,In_1301,In_441);
xor U172 (N_172,In_1074,In_510);
nand U173 (N_173,In_1240,In_1438);
and U174 (N_174,In_1169,In_749);
and U175 (N_175,In_1408,In_1660);
nor U176 (N_176,In_1914,In_1922);
or U177 (N_177,In_356,In_1859);
and U178 (N_178,In_555,In_911);
xor U179 (N_179,In_616,In_750);
xnor U180 (N_180,In_754,In_92);
and U181 (N_181,In_1542,In_147);
nand U182 (N_182,In_646,In_1375);
nand U183 (N_183,In_1726,In_865);
or U184 (N_184,In_411,In_674);
nor U185 (N_185,In_1101,In_1165);
xnor U186 (N_186,In_1563,In_452);
nor U187 (N_187,In_675,In_831);
nor U188 (N_188,In_1112,In_331);
and U189 (N_189,In_773,In_1430);
or U190 (N_190,In_1190,In_1209);
nand U191 (N_191,In_512,In_1974);
nor U192 (N_192,In_59,In_833);
nand U193 (N_193,In_493,In_977);
xor U194 (N_194,In_261,In_1117);
nand U195 (N_195,In_720,In_181);
nor U196 (N_196,In_528,In_908);
or U197 (N_197,In_1138,In_1007);
nand U198 (N_198,In_1858,In_1317);
xnor U199 (N_199,In_1577,In_1327);
and U200 (N_200,In_801,In_780);
nand U201 (N_201,In_1069,In_1738);
and U202 (N_202,In_766,In_1569);
nor U203 (N_203,In_1132,In_979);
xnor U204 (N_204,In_972,In_1719);
and U205 (N_205,In_40,In_843);
or U206 (N_206,In_1687,In_481);
and U207 (N_207,In_1691,In_741);
and U208 (N_208,In_1501,In_1556);
xor U209 (N_209,In_1358,In_866);
nand U210 (N_210,In_1057,In_426);
xor U211 (N_211,In_547,In_1661);
and U212 (N_212,In_70,In_1720);
xor U213 (N_213,In_718,In_1279);
and U214 (N_214,In_1873,In_1800);
or U215 (N_215,In_1149,In_873);
nor U216 (N_216,In_694,In_1781);
and U217 (N_217,In_27,In_1746);
xnor U218 (N_218,In_929,In_1507);
xor U219 (N_219,In_1678,In_1893);
or U220 (N_220,In_1186,In_1029);
nor U221 (N_221,In_1811,In_1311);
xor U222 (N_222,In_987,In_1482);
xnor U223 (N_223,In_119,In_303);
or U224 (N_224,In_580,In_1870);
and U225 (N_225,In_1052,In_969);
xnor U226 (N_226,In_1718,In_1999);
nand U227 (N_227,In_1338,In_1528);
and U228 (N_228,In_1004,In_150);
or U229 (N_229,In_308,In_362);
or U230 (N_230,In_579,In_472);
xor U231 (N_231,In_377,In_217);
nand U232 (N_232,In_934,In_994);
or U233 (N_233,In_497,In_971);
nand U234 (N_234,In_581,In_1651);
nor U235 (N_235,In_1454,In_86);
xnor U236 (N_236,In_1992,In_1641);
nor U237 (N_237,In_795,In_790);
nor U238 (N_238,In_1885,In_900);
nand U239 (N_239,In_986,In_340);
or U240 (N_240,In_357,In_1068);
xor U241 (N_241,In_508,In_1299);
nor U242 (N_242,In_706,In_429);
and U243 (N_243,In_1787,In_313);
or U244 (N_244,In_1144,In_1038);
nor U245 (N_245,In_1545,In_764);
and U246 (N_246,In_1667,In_136);
and U247 (N_247,In_1474,In_615);
nor U248 (N_248,In_328,In_1490);
or U249 (N_249,In_1258,In_15);
nand U250 (N_250,In_270,In_1183);
xor U251 (N_251,In_904,In_1705);
and U252 (N_252,In_1928,In_1418);
and U253 (N_253,In_743,In_1958);
and U254 (N_254,In_1948,In_189);
xor U255 (N_255,In_450,In_387);
nand U256 (N_256,In_1590,In_192);
nand U257 (N_257,In_1685,In_148);
or U258 (N_258,In_872,In_605);
nor U259 (N_259,In_112,In_1343);
nor U260 (N_260,In_632,In_753);
or U261 (N_261,In_651,In_1780);
xnor U262 (N_262,In_5,In_4);
nor U263 (N_263,In_1264,In_435);
xnor U264 (N_264,In_985,In_1192);
and U265 (N_265,In_1777,In_998);
nand U266 (N_266,In_1512,In_1040);
or U267 (N_267,In_906,In_1014);
nor U268 (N_268,In_1326,In_1330);
and U269 (N_269,In_1740,In_1424);
xnor U270 (N_270,In_315,In_1335);
and U271 (N_271,In_1287,In_34);
or U272 (N_272,In_408,In_103);
nand U273 (N_273,In_830,In_779);
or U274 (N_274,In_109,In_736);
nand U275 (N_275,In_1998,In_434);
or U276 (N_276,In_476,In_368);
or U277 (N_277,In_210,In_1339);
or U278 (N_278,In_1931,In_1508);
or U279 (N_279,In_1449,In_1598);
xnor U280 (N_280,In_1178,In_1682);
nor U281 (N_281,In_1773,In_761);
nor U282 (N_282,In_898,In_118);
nor U283 (N_283,In_401,In_1447);
nand U284 (N_284,In_1576,In_832);
and U285 (N_285,In_1530,In_896);
nor U286 (N_286,In_358,In_275);
xnor U287 (N_287,In_1462,In_57);
or U288 (N_288,In_114,In_1531);
nand U289 (N_289,In_1561,In_201);
or U290 (N_290,In_1096,In_124);
and U291 (N_291,In_1771,In_1076);
xnor U292 (N_292,In_69,In_1082);
or U293 (N_293,In_1141,In_840);
and U294 (N_294,In_544,In_1422);
nor U295 (N_295,In_566,In_653);
or U296 (N_296,In_1053,In_1690);
and U297 (N_297,In_304,In_1814);
and U298 (N_298,In_1081,In_859);
and U299 (N_299,In_1254,In_714);
xor U300 (N_300,In_1374,In_1803);
xnor U301 (N_301,In_1763,In_62);
or U302 (N_302,In_168,In_480);
xnor U303 (N_303,In_1717,In_1145);
and U304 (N_304,In_707,In_1697);
xor U305 (N_305,In_504,In_782);
and U306 (N_306,In_685,In_774);
nor U307 (N_307,In_1866,In_659);
or U308 (N_308,In_1960,In_297);
xor U309 (N_309,In_1621,In_734);
or U310 (N_310,In_1115,In_690);
nor U311 (N_311,In_1843,In_477);
nand U312 (N_312,In_1821,In_967);
nand U313 (N_313,In_268,In_468);
nand U314 (N_314,In_1748,In_45);
nor U315 (N_315,In_500,In_1645);
and U316 (N_316,In_794,In_557);
and U317 (N_317,In_61,In_1560);
or U318 (N_318,In_562,In_175);
xnor U319 (N_319,In_1571,In_1319);
and U320 (N_320,In_1329,In_1868);
or U321 (N_321,In_712,In_1706);
and U322 (N_322,In_1085,In_380);
or U323 (N_323,In_663,In_1731);
and U324 (N_324,In_1517,In_1927);
or U325 (N_325,In_141,In_1827);
or U326 (N_326,In_1849,In_1722);
and U327 (N_327,In_301,In_17);
nand U328 (N_328,In_54,In_1923);
and U329 (N_329,In_131,In_1900);
or U330 (N_330,In_1166,In_932);
or U331 (N_331,In_311,In_235);
or U332 (N_332,In_51,In_266);
nand U333 (N_333,In_1880,In_1309);
nand U334 (N_334,In_1448,In_179);
nor U335 (N_335,In_486,In_182);
xor U336 (N_336,In_1713,In_1286);
nand U337 (N_337,In_332,In_306);
xnor U338 (N_338,In_1088,In_447);
and U339 (N_339,In_1554,In_1184);
and U340 (N_340,In_1200,In_379);
and U341 (N_341,In_1704,In_888);
xor U342 (N_342,In_129,In_1990);
nand U343 (N_343,In_1437,In_229);
or U344 (N_344,In_467,In_144);
or U345 (N_345,In_1167,In_891);
or U346 (N_346,In_1975,In_1845);
and U347 (N_347,In_445,In_1608);
and U348 (N_348,In_1472,In_1765);
nand U349 (N_349,In_180,In_219);
xnor U350 (N_350,In_1801,In_1989);
nand U351 (N_351,In_1073,In_634);
or U352 (N_352,In_822,In_492);
or U353 (N_353,In_662,In_912);
nor U354 (N_354,In_804,In_215);
and U355 (N_355,In_1562,In_1202);
or U356 (N_356,In_1619,In_1951);
nand U357 (N_357,In_1881,In_1646);
and U358 (N_358,In_641,In_1712);
or U359 (N_359,In_836,In_746);
nor U360 (N_360,In_1273,In_531);
nand U361 (N_361,In_1944,In_1842);
nand U362 (N_362,In_1427,In_1952);
or U363 (N_363,In_1742,In_1041);
or U364 (N_364,In_1394,In_309);
nor U365 (N_365,In_240,In_1625);
nand U366 (N_366,In_276,In_163);
nand U367 (N_367,In_1371,In_1354);
xnor U368 (N_368,In_1032,In_1624);
and U369 (N_369,In_966,In_258);
or U370 (N_370,In_1812,In_454);
xor U371 (N_371,In_1936,In_366);
nand U372 (N_372,In_1419,In_960);
or U373 (N_373,In_1650,In_253);
nor U374 (N_374,In_564,In_1198);
nor U375 (N_375,In_1173,In_1152);
and U376 (N_376,In_570,In_1058);
or U377 (N_377,In_406,In_802);
xor U378 (N_378,In_920,In_1275);
nor U379 (N_379,In_1680,In_1599);
and U380 (N_380,In_922,In_130);
and U381 (N_381,In_974,In_758);
xor U382 (N_382,In_1337,In_1177);
nand U383 (N_383,In_543,In_1806);
or U384 (N_384,In_226,In_296);
xor U385 (N_385,In_1442,In_957);
or U386 (N_386,In_1961,In_534);
nor U387 (N_387,In_1872,In_807);
xor U388 (N_388,In_597,In_1629);
xor U389 (N_389,In_390,In_1465);
and U390 (N_390,In_1504,In_563);
nand U391 (N_391,In_1445,In_590);
nand U392 (N_392,In_1874,In_913);
and U393 (N_393,In_576,In_110);
and U394 (N_394,In_1212,In_1230);
nand U395 (N_395,In_870,In_1201);
nand U396 (N_396,In_1783,In_43);
nand U397 (N_397,In_1089,In_280);
and U398 (N_398,In_1251,In_1105);
and U399 (N_399,In_950,In_1581);
nor U400 (N_400,In_824,In_1652);
or U401 (N_401,In_1320,In_556);
xnor U402 (N_402,In_1984,In_1196);
and U403 (N_403,In_996,In_598);
nor U404 (N_404,In_1481,In_1372);
nor U405 (N_405,In_102,In_638);
or U406 (N_406,In_1925,In_256);
xnor U407 (N_407,In_1412,In_1476);
nand U408 (N_408,In_1864,In_1421);
or U409 (N_409,In_1679,In_730);
nor U410 (N_410,In_1968,In_1107);
nand U411 (N_411,In_784,In_871);
or U412 (N_412,In_251,In_364);
xnor U413 (N_413,In_1400,In_770);
xnor U414 (N_414,In_882,In_284);
and U415 (N_415,In_153,In_1229);
or U416 (N_416,In_277,In_654);
or U417 (N_417,In_1496,In_1709);
nor U418 (N_418,In_1256,In_1500);
nand U419 (N_419,In_1867,In_501);
or U420 (N_420,In_1216,In_1150);
nand U421 (N_421,In_1411,In_828);
xor U422 (N_422,In_1516,In_1905);
xnor U423 (N_423,In_907,In_755);
or U424 (N_424,In_1921,In_1632);
nor U425 (N_425,In_588,In_1574);
or U426 (N_426,In_1875,In_1478);
and U427 (N_427,In_113,In_1802);
or U428 (N_428,In_1463,In_725);
nor U429 (N_429,In_680,In_196);
or U430 (N_430,In_630,In_962);
nor U431 (N_431,In_1739,In_341);
nand U432 (N_432,In_1791,In_1217);
or U433 (N_433,In_729,In_1020);
and U434 (N_434,In_1477,In_1716);
and U435 (N_435,In_993,In_234);
nand U436 (N_436,In_1916,In_1877);
or U437 (N_437,In_1353,In_1813);
nand U438 (N_438,In_1930,In_811);
xnor U439 (N_439,In_1901,In_1884);
or U440 (N_440,In_781,In_796);
xnor U441 (N_441,In_1940,In_1659);
or U442 (N_442,In_1698,In_673);
nand U443 (N_443,In_1239,In_1283);
xnor U444 (N_444,In_1673,In_470);
and U445 (N_445,In_458,In_1988);
nand U446 (N_446,In_78,In_317);
or U447 (N_447,In_541,In_1271);
xnor U448 (N_448,In_667,In_637);
xnor U449 (N_449,In_1527,In_446);
xor U450 (N_450,In_978,In_885);
and U451 (N_451,In_672,In_1483);
or U452 (N_452,In_973,In_1696);
or U453 (N_453,In_530,In_704);
nand U454 (N_454,In_1023,In_37);
nor U455 (N_455,In_1793,In_727);
xor U456 (N_456,In_571,In_1784);
or U457 (N_457,In_517,In_693);
or U458 (N_458,In_744,In_132);
nor U459 (N_459,In_1788,In_35);
or U460 (N_460,In_752,In_1102);
nand U461 (N_461,In_22,In_1126);
or U462 (N_462,In_32,In_1695);
nand U463 (N_463,In_918,In_759);
xnor U464 (N_464,In_1826,In_1656);
xor U465 (N_465,In_705,In_1633);
or U466 (N_466,In_1161,In_402);
or U467 (N_467,In_6,In_1266);
or U468 (N_468,In_183,In_1824);
and U469 (N_469,In_247,In_1840);
nor U470 (N_470,In_798,In_1080);
nor U471 (N_471,In_227,In_522);
and U472 (N_472,In_1918,In_66);
xor U473 (N_473,In_448,In_413);
and U474 (N_474,In_1586,In_1046);
nand U475 (N_475,In_643,In_1091);
nor U476 (N_476,In_1794,In_1174);
or U477 (N_477,In_1658,In_1929);
nand U478 (N_478,In_771,In_1910);
nor U479 (N_479,In_629,In_1302);
nand U480 (N_480,In_552,In_624);
nand U481 (N_481,In_1996,In_1692);
and U482 (N_482,In_765,In_1006);
or U483 (N_483,In_1288,In_1087);
and U484 (N_484,In_1022,In_1924);
nor U485 (N_485,In_785,In_878);
xor U486 (N_486,In_419,In_1220);
or U487 (N_487,In_1917,In_686);
and U488 (N_488,In_1810,In_417);
nor U489 (N_489,In_1162,In_1026);
nand U490 (N_490,In_1155,In_384);
xnor U491 (N_491,In_457,In_1276);
nor U492 (N_492,In_117,In_1946);
and U493 (N_493,In_1331,In_42);
or U494 (N_494,In_516,In_471);
nand U495 (N_495,In_1681,In_10);
and U496 (N_496,In_1540,In_269);
xor U497 (N_497,In_264,In_1642);
or U498 (N_498,In_549,In_1861);
xor U499 (N_499,In_1446,In_901);
or U500 (N_500,In_1779,In_52);
nor U501 (N_501,In_428,In_533);
and U502 (N_502,In_1346,In_1334);
and U503 (N_503,In_152,In_649);
nor U504 (N_504,In_1983,In_53);
xor U505 (N_505,In_1171,In_1129);
and U506 (N_506,In_1061,In_334);
nor U507 (N_507,In_1050,In_485);
and U508 (N_508,In_594,In_1436);
or U509 (N_509,In_1176,In_1090);
or U510 (N_510,In_167,In_1649);
nand U511 (N_511,In_928,In_1755);
nand U512 (N_512,In_1350,In_1503);
and U513 (N_513,In_1965,In_1257);
xor U514 (N_514,In_1272,In_1314);
xnor U515 (N_515,In_1093,In_1766);
or U516 (N_516,In_31,In_1469);
or U517 (N_517,In_925,In_1060);
xnor U518 (N_518,In_1832,In_1522);
and U519 (N_519,In_463,In_1139);
xor U520 (N_520,In_681,In_383);
or U521 (N_521,In_561,In_1909);
nor U522 (N_522,In_438,In_756);
xor U523 (N_523,In_228,In_174);
and U524 (N_524,In_388,In_1142);
nor U525 (N_525,In_837,In_955);
and U526 (N_526,In_1296,In_1391);
nand U527 (N_527,In_244,In_1293);
nor U528 (N_528,In_938,In_1564);
or U529 (N_529,In_312,In_496);
nor U530 (N_530,In_139,In_1304);
and U531 (N_531,In_1714,In_342);
or U532 (N_532,In_1168,In_121);
and U533 (N_533,In_1466,In_791);
nor U534 (N_534,In_115,In_1414);
and U535 (N_535,In_513,In_821);
nand U536 (N_536,In_1741,In_606);
xor U537 (N_537,In_1432,In_834);
or U538 (N_538,In_116,In_149);
and U539 (N_539,In_1894,In_1510);
and U540 (N_540,In_614,In_869);
nor U541 (N_541,In_1282,In_887);
xor U542 (N_542,In_404,In_1307);
xor U543 (N_543,In_1479,In_1970);
or U544 (N_544,In_1003,In_620);
nand U545 (N_545,In_257,In_1541);
nor U546 (N_546,In_1365,In_860);
nor U547 (N_547,In_696,In_799);
or U548 (N_548,In_1906,In_1955);
or U549 (N_549,In_1829,In_572);
xnor U550 (N_550,In_1768,In_1135);
and U551 (N_551,In_1332,In_101);
nand U552 (N_552,In_1406,In_1322);
nor U553 (N_553,In_1441,In_96);
or U554 (N_554,In_1349,In_647);
nand U555 (N_555,In_1185,In_1389);
nand U556 (N_556,In_1815,In_487);
nor U557 (N_557,In_1298,In_1189);
nor U558 (N_558,In_224,In_664);
or U559 (N_559,In_923,In_1982);
nor U560 (N_560,In_1981,In_1151);
and U561 (N_561,In_1355,In_628);
and U562 (N_562,In_1031,In_1723);
nand U563 (N_563,In_1127,In_145);
nor U564 (N_564,In_381,In_786);
xnor U565 (N_565,In_425,In_584);
xnor U566 (N_566,In_1265,In_769);
nor U567 (N_567,In_1312,In_1044);
nand U568 (N_568,In_223,In_532);
or U569 (N_569,In_9,In_1677);
nand U570 (N_570,In_1662,In_1604);
and U571 (N_571,In_1747,In_7);
nor U572 (N_572,In_460,In_88);
or U573 (N_573,In_1492,In_1325);
and U574 (N_574,In_185,In_839);
or U575 (N_575,In_135,In_1131);
nor U576 (N_576,In_1363,In_951);
nand U577 (N_577,In_414,In_225);
nand U578 (N_578,In_1762,In_1423);
and U579 (N_579,In_1823,In_850);
and U580 (N_580,In_1347,In_212);
nand U581 (N_581,In_495,In_1847);
nand U582 (N_582,In_177,In_1933);
and U583 (N_583,In_293,In_1612);
xor U584 (N_584,In_1255,In_1786);
xnor U585 (N_585,In_1390,In_1180);
nand U586 (N_586,In_164,In_127);
xor U587 (N_587,In_194,In_1850);
nand U588 (N_588,In_155,In_558);
nor U589 (N_589,In_1876,In_1489);
nand U590 (N_590,In_1597,In_267);
nor U591 (N_591,In_1345,In_399);
and U592 (N_592,In_204,In_140);
nor U593 (N_593,In_619,In_1904);
xor U594 (N_594,In_108,In_762);
nand U595 (N_595,In_610,In_1486);
xnor U596 (N_596,In_363,In_976);
xor U597 (N_597,In_927,In_330);
nor U598 (N_598,In_855,In_604);
and U599 (N_599,In_63,In_760);
or U600 (N_600,In_55,In_176);
or U601 (N_601,In_793,In_1613);
and U602 (N_602,In_120,In_1035);
or U603 (N_603,In_1336,In_385);
nand U604 (N_604,In_601,In_85);
and U605 (N_605,In_514,In_997);
nand U606 (N_606,In_473,In_1809);
or U607 (N_607,In_724,In_64);
and U608 (N_608,In_1770,In_1025);
nor U609 (N_609,In_1380,In_286);
nor U610 (N_610,In_1208,In_949);
xor U611 (N_611,In_484,In_608);
and U612 (N_612,In_1790,In_943);
or U613 (N_613,In_1644,In_143);
nor U614 (N_614,In_845,In_583);
xnor U615 (N_615,In_1602,In_1062);
nor U616 (N_616,In_890,In_1453);
xnor U617 (N_617,In_1242,In_1595);
nor U618 (N_618,In_1879,In_36);
and U619 (N_619,In_1892,In_1323);
nand U620 (N_620,In_876,In_1782);
nor U621 (N_621,In_626,In_188);
and U622 (N_622,In_1559,In_142);
or U623 (N_623,In_159,In_1609);
nand U624 (N_624,In_1498,In_1244);
or U625 (N_625,In_1495,In_1405);
nor U626 (N_626,In_1888,In_89);
or U627 (N_627,In_838,In_1221);
nand U628 (N_628,In_1443,In_919);
nand U629 (N_629,In_440,In_65);
nor U630 (N_630,In_1828,In_1509);
nor U631 (N_631,In_1745,In_1710);
or U632 (N_632,In_930,In_1676);
nand U633 (N_633,In_1754,In_988);
nor U634 (N_634,In_200,In_657);
xor U635 (N_635,In_1260,In_372);
nand U636 (N_636,In_207,In_1146);
xor U637 (N_637,In_1361,In_410);
nor U638 (N_638,In_1392,In_991);
nand U639 (N_639,In_926,In_1245);
and U640 (N_640,In_431,In_1587);
nor U641 (N_641,In_483,In_1799);
or U642 (N_642,In_274,In_1816);
or U643 (N_643,In_1637,In_1665);
nor U644 (N_644,In_233,In_1225);
xor U645 (N_645,In_1205,In_862);
and U646 (N_646,In_1097,In_1707);
or U647 (N_647,In_1468,In_184);
nor U648 (N_648,In_238,In_1639);
xor U649 (N_649,In_8,In_1211);
or U650 (N_650,In_655,In_1818);
xnor U651 (N_651,In_44,In_405);
nand U652 (N_652,In_1401,In_669);
and U653 (N_653,In_1997,In_326);
nor U654 (N_654,In_1137,In_1557);
and U655 (N_655,In_1001,In_1499);
or U656 (N_656,In_80,In_700);
nand U657 (N_657,In_857,In_41);
nor U658 (N_658,In_68,In_1513);
or U659 (N_659,In_847,In_591);
nor U660 (N_660,In_232,In_1596);
nor U661 (N_661,In_721,In_1623);
nand U662 (N_662,In_939,In_715);
nor U663 (N_663,In_1744,In_1751);
and U664 (N_664,In_1536,In_1618);
nand U665 (N_665,In_1756,In_751);
and U666 (N_666,In_107,In_1013);
nand U667 (N_667,In_397,In_246);
or U668 (N_668,In_1341,In_1461);
xnor U669 (N_669,In_1402,In_917);
nand U670 (N_670,In_186,In_879);
and U671 (N_671,In_1529,In_193);
xor U672 (N_672,In_1605,In_964);
and U673 (N_673,In_635,In_678);
nand U674 (N_674,In_1385,In_1551);
nand U675 (N_675,In_808,In_73);
or U676 (N_676,In_953,In_491);
nor U677 (N_677,In_1525,In_545);
or U678 (N_678,In_1807,In_1666);
or U679 (N_679,In_1943,In_1838);
nor U680 (N_680,In_1377,In_314);
nor U681 (N_681,In_625,In_389);
and U682 (N_682,In_346,In_1699);
xor U683 (N_683,In_1019,In_1455);
nor U684 (N_684,In_980,In_1370);
nor U685 (N_685,In_1083,In_58);
nand U686 (N_686,In_1732,In_849);
xor U687 (N_687,In_524,In_1203);
nor U688 (N_688,In_1002,In_1973);
and U689 (N_689,In_1757,In_259);
nor U690 (N_690,In_1911,In_455);
and U691 (N_691,In_371,In_1324);
nand U692 (N_692,In_1603,In_236);
xor U693 (N_693,In_1399,In_1333);
and U694 (N_694,In_418,In_1285);
and U695 (N_695,In_1094,In_1686);
nor U696 (N_696,In_1396,In_1795);
nor U697 (N_697,In_1969,In_1364);
nand U698 (N_698,In_1075,In_713);
and U699 (N_699,In_535,In_1368);
or U700 (N_700,In_1125,In_1382);
and U701 (N_701,In_737,In_1450);
and U702 (N_702,In_1248,In_420);
nor U703 (N_703,In_378,In_1128);
or U704 (N_704,In_187,In_1425);
nor U705 (N_705,In_1475,In_665);
xor U706 (N_706,In_995,In_1711);
xor U707 (N_707,In_321,In_1444);
xnor U708 (N_708,In_199,In_1435);
nor U709 (N_709,In_1018,In_546);
and U710 (N_710,In_230,In_1000);
nand U711 (N_711,In_13,In_897);
xnor U712 (N_712,In_1417,In_797);
nand U713 (N_713,In_1538,In_1);
or U714 (N_714,In_861,In_1670);
or U715 (N_715,In_1759,In_203);
nand U716 (N_716,In_1518,In_1207);
or U717 (N_717,In_506,In_1197);
or U718 (N_718,In_1626,In_1407);
nand U719 (N_719,In_640,In_1388);
and U720 (N_720,In_1114,In_327);
nor U721 (N_721,In_742,In_817);
and U722 (N_722,In_138,In_668);
nor U723 (N_723,In_423,In_1313);
or U724 (N_724,In_569,In_1846);
nor U725 (N_725,In_763,In_1778);
xnor U726 (N_726,In_437,In_1170);
and U727 (N_727,In_568,In_375);
and U728 (N_728,In_1957,In_1734);
xnor U729 (N_729,In_1582,In_218);
nor U730 (N_730,In_1535,In_1926);
nor U731 (N_731,In_803,In_1100);
nand U732 (N_732,In_963,In_1514);
or U733 (N_733,In_49,In_432);
xnor U734 (N_734,In_1737,In_1005);
and U735 (N_735,In_1278,In_1259);
xnor U736 (N_736,In_525,In_1379);
nand U737 (N_737,In_26,In_82);
xor U738 (N_738,In_1181,In_722);
and U739 (N_739,In_1223,In_1433);
nand U740 (N_740,In_1280,In_1654);
and U741 (N_741,In_394,In_1484);
and U742 (N_742,In_1063,In_329);
or U743 (N_743,In_1292,In_1066);
or U744 (N_744,In_1907,In_1123);
nor U745 (N_745,In_1727,In_24);
and U746 (N_746,In_351,In_1552);
xor U747 (N_747,In_319,In_1344);
nor U748 (N_748,In_474,In_553);
and U749 (N_749,In_248,In_965);
or U750 (N_750,In_1947,In_639);
or U751 (N_751,In_1938,In_1281);
xnor U752 (N_752,In_1977,In_1694);
or U753 (N_753,In_1964,In_1854);
xnor U754 (N_754,In_1267,In_339);
nand U755 (N_755,In_1274,In_1195);
nor U756 (N_756,In_166,In_302);
or U757 (N_757,In_427,In_1488);
nor U758 (N_758,In_1702,In_1725);
and U759 (N_759,In_323,In_745);
nand U760 (N_760,In_335,In_1792);
or U761 (N_761,In_1819,In_592);
or U762 (N_762,In_1182,In_172);
nor U763 (N_763,In_1456,In_924);
or U764 (N_764,In_596,In_944);
xnor U765 (N_765,In_679,In_844);
nand U766 (N_766,In_1294,In_1822);
and U767 (N_767,In_1937,In_688);
xor U768 (N_768,In_271,In_1841);
nand U769 (N_769,In_1607,In_1769);
nand U770 (N_770,In_333,In_1878);
xnor U771 (N_771,In_935,In_650);
nor U772 (N_772,In_1882,In_1051);
and U773 (N_773,In_777,In_1539);
or U774 (N_774,In_767,In_848);
or U775 (N_775,In_642,In_1869);
or U776 (N_776,In_433,In_1932);
xor U777 (N_777,In_456,In_1550);
xnor U778 (N_778,In_324,In_282);
xor U779 (N_779,In_1683,In_1615);
xnor U780 (N_780,In_916,In_361);
nand U781 (N_781,In_1172,In_867);
nand U782 (N_782,In_600,In_1862);
or U783 (N_783,In_940,In_809);
or U784 (N_784,In_1836,In_1585);
and U785 (N_785,In_703,In_81);
nor U786 (N_786,In_295,In_902);
or U787 (N_787,In_701,In_344);
and U788 (N_788,In_740,In_946);
nand U789 (N_789,In_894,In_1967);
nor U790 (N_790,In_880,In_1284);
xor U791 (N_791,In_1413,In_941);
nor U792 (N_792,In_551,In_1956);
or U793 (N_793,In_104,In_195);
xnor U794 (N_794,In_1896,In_1121);
and U795 (N_795,In_1356,In_1110);
nor U796 (N_796,In_578,In_466);
or U797 (N_797,In_254,In_518);
xnor U798 (N_798,In_815,In_892);
and U799 (N_799,In_1547,In_1403);
nor U800 (N_800,In_910,In_1573);
nor U801 (N_801,In_851,In_1485);
nor U802 (N_802,In_252,In_1415);
and U803 (N_803,In_970,In_1393);
nand U804 (N_804,In_1567,In_294);
and U805 (N_805,In_376,In_670);
or U806 (N_806,In_1611,In_1119);
or U807 (N_807,In_644,In_593);
xor U808 (N_808,In_1749,In_1048);
nand U809 (N_809,In_1440,In_75);
nand U810 (N_810,In_835,In_1565);
xnor U811 (N_811,In_1526,In_157);
xor U812 (N_812,In_29,In_787);
and U813 (N_813,In_1303,In_1533);
and U814 (N_814,In_1934,In_30);
xor U815 (N_815,In_1617,In_255);
nand U816 (N_816,In_11,In_21);
nand U817 (N_817,In_1219,In_211);
nand U818 (N_818,In_1143,In_1378);
xor U819 (N_819,In_1736,In_1124);
xor U820 (N_820,In_170,In_373);
nor U821 (N_821,In_1118,In_1154);
nor U822 (N_822,In_288,In_1157);
or U823 (N_823,In_393,In_565);
nor U824 (N_824,In_1647,In_858);
xor U825 (N_825,In_20,In_582);
nand U826 (N_826,In_1268,In_122);
nand U827 (N_827,In_1021,In_369);
or U828 (N_828,In_1627,In_1113);
nand U829 (N_829,In_1663,In_827);
nand U830 (N_830,In_197,In_1213);
nand U831 (N_831,In_415,In_1428);
xnor U832 (N_832,In_1622,In_1669);
and U833 (N_833,In_289,In_1136);
xnor U834 (N_834,In_1224,In_511);
and U835 (N_835,In_800,In_1584);
and U836 (N_836,In_237,In_156);
nor U837 (N_837,In_90,In_1591);
xnor U838 (N_838,In_465,In_1579);
nand U839 (N_839,In_1116,In_812);
xor U840 (N_840,In_105,In_325);
nand U841 (N_841,In_1505,In_94);
nor U842 (N_842,In_1568,In_449);
xnor U843 (N_843,In_1589,In_1104);
and U844 (N_844,In_710,In_875);
or U845 (N_845,In_914,In_1369);
xor U846 (N_846,In_79,In_550);
nor U847 (N_847,In_99,In_1270);
nand U848 (N_848,In_1078,In_1099);
nand U849 (N_849,In_260,In_1289);
xnor U850 (N_850,In_1404,In_768);
or U851 (N_851,In_595,In_1805);
xor U852 (N_852,In_567,In_1342);
or U853 (N_853,In_279,In_1277);
nor U854 (N_854,In_1753,In_1011);
or U855 (N_855,In_874,In_952);
or U856 (N_856,In_1903,In_1758);
nor U857 (N_857,In_1199,In_1459);
nand U858 (N_858,In_536,In_1084);
and U859 (N_859,In_1640,In_1416);
and U860 (N_860,In_1575,In_430);
xor U861 (N_861,In_403,In_1206);
nor U862 (N_862,In_1628,In_347);
xnor U863 (N_863,In_1935,In_191);
xor U864 (N_864,In_1583,In_864);
or U865 (N_865,In_360,In_365);
nand U866 (N_866,In_1735,In_968);
or U867 (N_867,In_74,In_1785);
xor U868 (N_868,In_443,In_1460);
xor U869 (N_869,In_539,In_1945);
xor U870 (N_870,In_1570,In_999);
nor U871 (N_871,In_1008,In_1188);
xor U872 (N_872,In_886,In_1387);
xor U873 (N_873,In_1049,In_1236);
or U874 (N_874,In_854,In_1232);
and U875 (N_875,In_1519,In_396);
nand U876 (N_876,In_823,In_788);
nor U877 (N_877,In_587,In_97);
and U878 (N_878,In_1721,In_697);
and U879 (N_879,In_213,In_1630);
nor U880 (N_880,In_1671,In_1111);
and U881 (N_881,In_618,In_462);
and U882 (N_882,In_91,In_1410);
and U883 (N_883,In_684,In_482);
or U884 (N_884,In_461,In_310);
and U885 (N_885,In_1855,In_95);
nand U886 (N_886,In_479,In_682);
and U887 (N_887,In_1384,In_1473);
nor U888 (N_888,In_989,In_1098);
xnor U889 (N_889,In_1252,In_214);
xnor U890 (N_890,In_1601,In_1261);
xor U891 (N_891,In_178,In_1761);
xnor U892 (N_892,In_1054,In_1703);
or U893 (N_893,In_738,In_1902);
or U894 (N_894,In_1253,In_1070);
or U895 (N_895,In_1636,In_1366);
nand U896 (N_896,In_1620,In_633);
nor U897 (N_897,In_1269,In_1708);
nand U898 (N_898,In_825,In_1470);
nand U899 (N_899,In_1480,In_559);
nand U900 (N_900,In_158,In_1439);
xnor U901 (N_901,In_687,In_47);
and U902 (N_902,In_1016,In_1210);
or U903 (N_903,In_1017,In_909);
nor U904 (N_904,In_488,In_683);
nor U905 (N_905,In_1657,In_691);
and U906 (N_906,In_1524,In_370);
xor U907 (N_907,In_1954,In_711);
nor U908 (N_908,In_1774,In_1750);
nand U909 (N_909,In_863,In_903);
nand U910 (N_910,In_422,In_1426);
and U911 (N_911,In_1130,In_1808);
and U912 (N_912,In_1451,In_48);
or U913 (N_913,In_1156,In_498);
nor U914 (N_914,In_453,In_607);
nor U915 (N_915,In_1194,In_538);
nand U916 (N_916,In_984,In_881);
or U917 (N_917,In_1065,In_1122);
and U918 (N_918,In_1306,In_169);
xnor U919 (N_919,In_1193,In_93);
nand U920 (N_920,In_1179,In_853);
nor U921 (N_921,In_316,In_732);
and U922 (N_922,In_589,In_1009);
nor U923 (N_923,In_398,In_658);
xor U924 (N_924,In_1980,In_1693);
and U925 (N_925,In_459,In_523);
xnor U926 (N_926,In_1235,In_137);
or U927 (N_927,In_1305,In_1064);
nand U928 (N_928,In_1511,In_1844);
xor U929 (N_929,In_161,In_1543);
xnor U930 (N_930,In_783,In_1095);
xor U931 (N_931,In_1897,In_1243);
xor U932 (N_932,In_1241,In_72);
and U933 (N_933,In_609,In_599);
and U934 (N_934,In_990,In_126);
nand U935 (N_935,In_947,In_1163);
or U936 (N_936,In_699,In_281);
nor U937 (N_937,In_1228,In_359);
nand U938 (N_938,In_1942,In_1941);
nand U939 (N_939,In_1655,In_505);
nor U940 (N_940,In_1871,In_171);
and U941 (N_941,In_1028,In_1772);
xor U942 (N_942,In_1700,In_945);
nor U943 (N_943,In_243,In_621);
nand U944 (N_944,In_1357,In_291);
nand U945 (N_945,In_1915,In_612);
nand U946 (N_946,In_1887,In_603);
or U947 (N_947,In_353,In_400);
nand U948 (N_948,In_1856,In_1852);
and U949 (N_949,In_883,In_1316);
nand U950 (N_950,In_412,In_757);
or U951 (N_951,In_198,In_1995);
nand U952 (N_952,In_111,In_19);
nor U953 (N_953,In_1133,In_320);
nor U954 (N_954,In_554,In_87);
or U955 (N_955,In_656,In_1537);
or U956 (N_956,In_1521,In_1588);
nand U957 (N_957,In_921,In_1971);
nor U958 (N_958,In_1993,In_1295);
and U959 (N_959,In_1351,In_1949);
nor U960 (N_960,In_1804,In_23);
nand U961 (N_961,In_1789,In_12);
nand U962 (N_962,In_1033,In_1420);
nand U963 (N_963,In_1109,In_537);
nand U964 (N_964,In_613,In_1153);
nor U965 (N_965,In_1191,In_1027);
xnor U966 (N_966,In_499,In_382);
nand U967 (N_967,In_915,In_792);
or U968 (N_968,In_1606,In_220);
or U969 (N_969,In_1674,In_1865);
nand U970 (N_970,In_1994,In_1886);
or U971 (N_971,In_14,In_151);
and U972 (N_972,In_25,In_1899);
and U973 (N_973,In_1494,In_205);
xnor U974 (N_974,In_469,In_1555);
or U975 (N_975,In_1092,In_548);
nor U976 (N_976,In_877,In_355);
and U977 (N_977,In_3,In_526);
xor U978 (N_978,In_1835,In_173);
nand U979 (N_979,In_527,In_100);
xor U980 (N_980,In_1262,In_975);
nor U981 (N_981,In_28,In_1497);
nor U982 (N_982,In_1853,In_692);
nor U983 (N_983,In_813,In_1546);
and U984 (N_984,In_1204,In_1222);
and U985 (N_985,In_1263,In_1908);
xor U986 (N_986,In_1227,In_1523);
nand U987 (N_987,In_1775,In_409);
xor U988 (N_988,In_1250,In_338);
and U989 (N_989,In_1764,In_1328);
or U990 (N_990,In_689,In_1978);
xnor U991 (N_991,In_1600,In_1237);
nand U992 (N_992,In_1467,In_318);
and U993 (N_993,In_1047,In_816);
or U994 (N_994,In_717,In_1108);
nor U995 (N_995,In_1966,In_1291);
nand U996 (N_996,In_1315,In_1548);
nand U997 (N_997,In_1668,In_895);
nand U998 (N_998,In_33,In_648);
and U999 (N_999,In_1729,In_778);
and U1000 (N_1000,In_1789,In_1191);
xor U1001 (N_1001,In_1698,In_836);
nand U1002 (N_1002,In_1285,In_1906);
nor U1003 (N_1003,In_304,In_1162);
nor U1004 (N_1004,In_1858,In_459);
or U1005 (N_1005,In_1928,In_1071);
nor U1006 (N_1006,In_1933,In_1756);
nor U1007 (N_1007,In_1131,In_28);
xor U1008 (N_1008,In_1826,In_1290);
xnor U1009 (N_1009,In_763,In_1999);
nor U1010 (N_1010,In_381,In_1390);
nand U1011 (N_1011,In_1552,In_1590);
nand U1012 (N_1012,In_1171,In_670);
xor U1013 (N_1013,In_1615,In_184);
and U1014 (N_1014,In_1422,In_986);
nor U1015 (N_1015,In_969,In_1729);
or U1016 (N_1016,In_1936,In_1760);
nand U1017 (N_1017,In_174,In_1999);
nor U1018 (N_1018,In_582,In_1475);
or U1019 (N_1019,In_1372,In_1860);
and U1020 (N_1020,In_340,In_405);
nand U1021 (N_1021,In_585,In_1689);
or U1022 (N_1022,In_1164,In_786);
or U1023 (N_1023,In_1678,In_1550);
nand U1024 (N_1024,In_541,In_1177);
xnor U1025 (N_1025,In_137,In_1158);
or U1026 (N_1026,In_1215,In_1545);
or U1027 (N_1027,In_11,In_222);
nand U1028 (N_1028,In_786,In_1554);
nand U1029 (N_1029,In_1415,In_1247);
xnor U1030 (N_1030,In_26,In_1706);
and U1031 (N_1031,In_389,In_1210);
and U1032 (N_1032,In_347,In_839);
and U1033 (N_1033,In_603,In_1609);
xnor U1034 (N_1034,In_1087,In_24);
or U1035 (N_1035,In_497,In_1769);
nand U1036 (N_1036,In_1767,In_380);
nand U1037 (N_1037,In_49,In_651);
xor U1038 (N_1038,In_263,In_1433);
nor U1039 (N_1039,In_1669,In_1877);
or U1040 (N_1040,In_785,In_1298);
or U1041 (N_1041,In_570,In_212);
nand U1042 (N_1042,In_1870,In_1796);
and U1043 (N_1043,In_996,In_1347);
nand U1044 (N_1044,In_1879,In_750);
nor U1045 (N_1045,In_327,In_642);
nor U1046 (N_1046,In_728,In_1447);
xnor U1047 (N_1047,In_718,In_831);
xnor U1048 (N_1048,In_226,In_1582);
or U1049 (N_1049,In_344,In_264);
and U1050 (N_1050,In_381,In_1148);
nand U1051 (N_1051,In_194,In_738);
and U1052 (N_1052,In_637,In_86);
and U1053 (N_1053,In_580,In_1998);
or U1054 (N_1054,In_1300,In_1464);
nor U1055 (N_1055,In_1109,In_1711);
xnor U1056 (N_1056,In_1441,In_912);
and U1057 (N_1057,In_1913,In_1908);
nand U1058 (N_1058,In_1810,In_1959);
nor U1059 (N_1059,In_1914,In_444);
nor U1060 (N_1060,In_832,In_803);
nor U1061 (N_1061,In_1772,In_573);
nor U1062 (N_1062,In_372,In_1849);
or U1063 (N_1063,In_1932,In_1008);
nor U1064 (N_1064,In_1788,In_1795);
nand U1065 (N_1065,In_830,In_1914);
nor U1066 (N_1066,In_1421,In_1173);
nand U1067 (N_1067,In_1295,In_1101);
and U1068 (N_1068,In_305,In_726);
or U1069 (N_1069,In_502,In_1956);
and U1070 (N_1070,In_366,In_560);
or U1071 (N_1071,In_213,In_1552);
and U1072 (N_1072,In_1471,In_807);
xnor U1073 (N_1073,In_246,In_16);
and U1074 (N_1074,In_470,In_1233);
xnor U1075 (N_1075,In_1302,In_692);
nor U1076 (N_1076,In_1664,In_1398);
xor U1077 (N_1077,In_153,In_1354);
xnor U1078 (N_1078,In_1055,In_1034);
nand U1079 (N_1079,In_606,In_1194);
nand U1080 (N_1080,In_875,In_340);
or U1081 (N_1081,In_523,In_1046);
or U1082 (N_1082,In_983,In_346);
nand U1083 (N_1083,In_1336,In_1825);
and U1084 (N_1084,In_1741,In_1536);
xnor U1085 (N_1085,In_504,In_1641);
nand U1086 (N_1086,In_477,In_680);
or U1087 (N_1087,In_1223,In_509);
nand U1088 (N_1088,In_1724,In_152);
nor U1089 (N_1089,In_977,In_1818);
nor U1090 (N_1090,In_1624,In_103);
or U1091 (N_1091,In_1497,In_574);
and U1092 (N_1092,In_29,In_953);
nand U1093 (N_1093,In_433,In_424);
nor U1094 (N_1094,In_156,In_1442);
or U1095 (N_1095,In_1121,In_1203);
xnor U1096 (N_1096,In_1573,In_1991);
and U1097 (N_1097,In_1924,In_1926);
and U1098 (N_1098,In_1795,In_1823);
nor U1099 (N_1099,In_1397,In_970);
nor U1100 (N_1100,In_385,In_1588);
and U1101 (N_1101,In_354,In_346);
nand U1102 (N_1102,In_286,In_870);
xnor U1103 (N_1103,In_27,In_1743);
nand U1104 (N_1104,In_1763,In_583);
nand U1105 (N_1105,In_151,In_1209);
nand U1106 (N_1106,In_634,In_1283);
or U1107 (N_1107,In_1331,In_1324);
nor U1108 (N_1108,In_310,In_969);
nor U1109 (N_1109,In_1006,In_1274);
and U1110 (N_1110,In_1819,In_502);
nand U1111 (N_1111,In_177,In_1334);
and U1112 (N_1112,In_102,In_1473);
xor U1113 (N_1113,In_1778,In_916);
xor U1114 (N_1114,In_1117,In_1171);
or U1115 (N_1115,In_675,In_1165);
nand U1116 (N_1116,In_674,In_1257);
or U1117 (N_1117,In_87,In_1298);
nor U1118 (N_1118,In_1994,In_563);
nand U1119 (N_1119,In_1040,In_710);
or U1120 (N_1120,In_1099,In_1589);
and U1121 (N_1121,In_596,In_1062);
and U1122 (N_1122,In_1009,In_122);
xor U1123 (N_1123,In_494,In_269);
xnor U1124 (N_1124,In_1134,In_881);
nor U1125 (N_1125,In_396,In_592);
nor U1126 (N_1126,In_118,In_1992);
nand U1127 (N_1127,In_1077,In_779);
nand U1128 (N_1128,In_210,In_938);
or U1129 (N_1129,In_496,In_1053);
nor U1130 (N_1130,In_421,In_1762);
nand U1131 (N_1131,In_1494,In_1412);
nand U1132 (N_1132,In_818,In_1938);
nand U1133 (N_1133,In_981,In_179);
or U1134 (N_1134,In_568,In_1440);
nand U1135 (N_1135,In_1420,In_864);
nand U1136 (N_1136,In_1653,In_1183);
or U1137 (N_1137,In_3,In_65);
nor U1138 (N_1138,In_948,In_1607);
xor U1139 (N_1139,In_352,In_1238);
xor U1140 (N_1140,In_323,In_428);
nor U1141 (N_1141,In_1963,In_145);
and U1142 (N_1142,In_1522,In_224);
nand U1143 (N_1143,In_600,In_742);
nor U1144 (N_1144,In_407,In_523);
and U1145 (N_1145,In_1481,In_201);
or U1146 (N_1146,In_1043,In_457);
nor U1147 (N_1147,In_680,In_1885);
nor U1148 (N_1148,In_463,In_769);
and U1149 (N_1149,In_415,In_1727);
xnor U1150 (N_1150,In_1488,In_38);
nand U1151 (N_1151,In_1699,In_498);
or U1152 (N_1152,In_767,In_1257);
or U1153 (N_1153,In_1464,In_1954);
nor U1154 (N_1154,In_1863,In_1703);
xnor U1155 (N_1155,In_1180,In_1817);
and U1156 (N_1156,In_83,In_81);
nor U1157 (N_1157,In_972,In_385);
nor U1158 (N_1158,In_575,In_1978);
nand U1159 (N_1159,In_1466,In_1226);
or U1160 (N_1160,In_862,In_456);
xor U1161 (N_1161,In_1769,In_1419);
nor U1162 (N_1162,In_1386,In_1314);
nor U1163 (N_1163,In_366,In_227);
nand U1164 (N_1164,In_188,In_1615);
xor U1165 (N_1165,In_797,In_1446);
xor U1166 (N_1166,In_1086,In_1582);
and U1167 (N_1167,In_1893,In_1180);
and U1168 (N_1168,In_55,In_1187);
and U1169 (N_1169,In_1710,In_591);
xor U1170 (N_1170,In_884,In_1140);
xor U1171 (N_1171,In_153,In_1934);
xor U1172 (N_1172,In_294,In_688);
and U1173 (N_1173,In_1259,In_1640);
or U1174 (N_1174,In_1984,In_73);
xor U1175 (N_1175,In_775,In_1400);
nand U1176 (N_1176,In_1744,In_280);
or U1177 (N_1177,In_1118,In_1189);
and U1178 (N_1178,In_1906,In_1190);
nor U1179 (N_1179,In_83,In_1560);
or U1180 (N_1180,In_205,In_563);
and U1181 (N_1181,In_1421,In_70);
nand U1182 (N_1182,In_453,In_1693);
nand U1183 (N_1183,In_660,In_1204);
nand U1184 (N_1184,In_1941,In_1128);
and U1185 (N_1185,In_796,In_63);
or U1186 (N_1186,In_206,In_552);
or U1187 (N_1187,In_592,In_845);
or U1188 (N_1188,In_1005,In_1135);
and U1189 (N_1189,In_932,In_1760);
nand U1190 (N_1190,In_1457,In_1917);
or U1191 (N_1191,In_864,In_1943);
or U1192 (N_1192,In_1414,In_1481);
or U1193 (N_1193,In_398,In_725);
and U1194 (N_1194,In_1359,In_860);
nor U1195 (N_1195,In_1995,In_980);
or U1196 (N_1196,In_19,In_1737);
or U1197 (N_1197,In_1921,In_617);
and U1198 (N_1198,In_1519,In_1795);
nand U1199 (N_1199,In_655,In_313);
nor U1200 (N_1200,In_692,In_312);
nand U1201 (N_1201,In_1597,In_1868);
and U1202 (N_1202,In_401,In_308);
nor U1203 (N_1203,In_572,In_1579);
or U1204 (N_1204,In_283,In_142);
or U1205 (N_1205,In_1711,In_1474);
or U1206 (N_1206,In_1315,In_742);
nor U1207 (N_1207,In_1257,In_826);
nor U1208 (N_1208,In_212,In_1674);
and U1209 (N_1209,In_1194,In_1491);
and U1210 (N_1210,In_268,In_1198);
or U1211 (N_1211,In_1864,In_1022);
nand U1212 (N_1212,In_1750,In_1386);
xnor U1213 (N_1213,In_1771,In_1509);
xor U1214 (N_1214,In_1127,In_1275);
xnor U1215 (N_1215,In_1962,In_1871);
nor U1216 (N_1216,In_28,In_926);
nor U1217 (N_1217,In_216,In_22);
nand U1218 (N_1218,In_242,In_1954);
nor U1219 (N_1219,In_1313,In_89);
nor U1220 (N_1220,In_1935,In_13);
xnor U1221 (N_1221,In_1040,In_1256);
and U1222 (N_1222,In_996,In_148);
xnor U1223 (N_1223,In_283,In_1240);
nand U1224 (N_1224,In_437,In_342);
or U1225 (N_1225,In_948,In_1547);
or U1226 (N_1226,In_1055,In_380);
and U1227 (N_1227,In_778,In_917);
xnor U1228 (N_1228,In_99,In_523);
nor U1229 (N_1229,In_658,In_1682);
xnor U1230 (N_1230,In_1463,In_667);
xnor U1231 (N_1231,In_748,In_1567);
and U1232 (N_1232,In_886,In_818);
or U1233 (N_1233,In_780,In_1039);
and U1234 (N_1234,In_520,In_537);
nand U1235 (N_1235,In_371,In_849);
xor U1236 (N_1236,In_1036,In_1121);
and U1237 (N_1237,In_1022,In_1397);
nor U1238 (N_1238,In_1751,In_1164);
xnor U1239 (N_1239,In_831,In_1508);
and U1240 (N_1240,In_457,In_1979);
nand U1241 (N_1241,In_1541,In_20);
xor U1242 (N_1242,In_773,In_1903);
and U1243 (N_1243,In_1588,In_248);
nor U1244 (N_1244,In_37,In_842);
and U1245 (N_1245,In_623,In_761);
xor U1246 (N_1246,In_127,In_929);
nand U1247 (N_1247,In_242,In_8);
nand U1248 (N_1248,In_1091,In_735);
xor U1249 (N_1249,In_819,In_828);
xnor U1250 (N_1250,In_1036,In_1344);
or U1251 (N_1251,In_846,In_781);
nor U1252 (N_1252,In_176,In_1273);
nand U1253 (N_1253,In_182,In_390);
nor U1254 (N_1254,In_546,In_1954);
and U1255 (N_1255,In_49,In_1511);
nand U1256 (N_1256,In_1774,In_1567);
nor U1257 (N_1257,In_101,In_708);
nand U1258 (N_1258,In_1537,In_418);
xnor U1259 (N_1259,In_619,In_748);
or U1260 (N_1260,In_1343,In_1759);
or U1261 (N_1261,In_164,In_85);
or U1262 (N_1262,In_1276,In_1146);
and U1263 (N_1263,In_1606,In_1292);
and U1264 (N_1264,In_1402,In_529);
and U1265 (N_1265,In_613,In_132);
nor U1266 (N_1266,In_42,In_299);
xnor U1267 (N_1267,In_759,In_70);
xor U1268 (N_1268,In_1448,In_168);
nand U1269 (N_1269,In_1430,In_582);
nor U1270 (N_1270,In_1889,In_666);
or U1271 (N_1271,In_746,In_368);
nand U1272 (N_1272,In_1117,In_1267);
and U1273 (N_1273,In_15,In_694);
nand U1274 (N_1274,In_1426,In_1908);
and U1275 (N_1275,In_645,In_236);
and U1276 (N_1276,In_756,In_1550);
nand U1277 (N_1277,In_94,In_669);
or U1278 (N_1278,In_110,In_1977);
and U1279 (N_1279,In_1266,In_355);
or U1280 (N_1280,In_508,In_631);
xnor U1281 (N_1281,In_1566,In_861);
nand U1282 (N_1282,In_1969,In_226);
and U1283 (N_1283,In_1253,In_1023);
xnor U1284 (N_1284,In_1886,In_1188);
and U1285 (N_1285,In_1153,In_68);
or U1286 (N_1286,In_375,In_1089);
nand U1287 (N_1287,In_963,In_1544);
nor U1288 (N_1288,In_1264,In_922);
and U1289 (N_1289,In_1455,In_554);
or U1290 (N_1290,In_281,In_1668);
nor U1291 (N_1291,In_849,In_1097);
and U1292 (N_1292,In_1487,In_188);
or U1293 (N_1293,In_1396,In_1015);
and U1294 (N_1294,In_376,In_1044);
and U1295 (N_1295,In_1262,In_1800);
nand U1296 (N_1296,In_865,In_1621);
nor U1297 (N_1297,In_1751,In_875);
or U1298 (N_1298,In_213,In_971);
or U1299 (N_1299,In_695,In_1372);
nand U1300 (N_1300,In_1224,In_1111);
or U1301 (N_1301,In_1639,In_1450);
nor U1302 (N_1302,In_847,In_912);
nand U1303 (N_1303,In_537,In_1528);
and U1304 (N_1304,In_1534,In_396);
nor U1305 (N_1305,In_1102,In_1841);
nor U1306 (N_1306,In_1608,In_964);
xnor U1307 (N_1307,In_1875,In_904);
or U1308 (N_1308,In_1607,In_1208);
nand U1309 (N_1309,In_1139,In_286);
and U1310 (N_1310,In_1038,In_922);
nor U1311 (N_1311,In_6,In_371);
and U1312 (N_1312,In_1356,In_1944);
and U1313 (N_1313,In_71,In_1390);
nor U1314 (N_1314,In_1401,In_285);
nor U1315 (N_1315,In_1513,In_467);
and U1316 (N_1316,In_1798,In_882);
xnor U1317 (N_1317,In_1028,In_347);
nor U1318 (N_1318,In_1894,In_1602);
and U1319 (N_1319,In_751,In_1020);
xor U1320 (N_1320,In_1960,In_1020);
or U1321 (N_1321,In_70,In_912);
xor U1322 (N_1322,In_1435,In_1649);
and U1323 (N_1323,In_440,In_1802);
nor U1324 (N_1324,In_255,In_333);
xnor U1325 (N_1325,In_1806,In_437);
and U1326 (N_1326,In_1923,In_255);
xnor U1327 (N_1327,In_796,In_784);
nor U1328 (N_1328,In_713,In_1649);
or U1329 (N_1329,In_1882,In_1563);
xnor U1330 (N_1330,In_1963,In_836);
or U1331 (N_1331,In_1425,In_1014);
and U1332 (N_1332,In_314,In_181);
nor U1333 (N_1333,In_1731,In_252);
nand U1334 (N_1334,In_1346,In_1876);
nand U1335 (N_1335,In_392,In_333);
nor U1336 (N_1336,In_708,In_1647);
or U1337 (N_1337,In_1040,In_352);
and U1338 (N_1338,In_1579,In_827);
xor U1339 (N_1339,In_792,In_1948);
and U1340 (N_1340,In_454,In_548);
nor U1341 (N_1341,In_205,In_415);
nor U1342 (N_1342,In_526,In_856);
xnor U1343 (N_1343,In_1956,In_1144);
or U1344 (N_1344,In_1949,In_1283);
nor U1345 (N_1345,In_560,In_517);
nand U1346 (N_1346,In_658,In_1166);
xnor U1347 (N_1347,In_675,In_804);
nand U1348 (N_1348,In_656,In_579);
nand U1349 (N_1349,In_515,In_1547);
xor U1350 (N_1350,In_1651,In_888);
xor U1351 (N_1351,In_408,In_1030);
nand U1352 (N_1352,In_282,In_460);
nand U1353 (N_1353,In_1716,In_1959);
nand U1354 (N_1354,In_1803,In_396);
or U1355 (N_1355,In_1960,In_1684);
nor U1356 (N_1356,In_769,In_1571);
nor U1357 (N_1357,In_637,In_1044);
or U1358 (N_1358,In_352,In_1566);
or U1359 (N_1359,In_1157,In_1534);
nand U1360 (N_1360,In_1568,In_1697);
and U1361 (N_1361,In_1382,In_216);
nor U1362 (N_1362,In_1725,In_917);
xor U1363 (N_1363,In_1571,In_1960);
and U1364 (N_1364,In_74,In_897);
or U1365 (N_1365,In_1647,In_208);
xor U1366 (N_1366,In_1775,In_1249);
nand U1367 (N_1367,In_1467,In_1017);
and U1368 (N_1368,In_75,In_1681);
or U1369 (N_1369,In_417,In_1844);
or U1370 (N_1370,In_446,In_1574);
or U1371 (N_1371,In_1396,In_78);
and U1372 (N_1372,In_1160,In_1542);
and U1373 (N_1373,In_1338,In_1399);
nand U1374 (N_1374,In_1865,In_485);
nor U1375 (N_1375,In_760,In_143);
nand U1376 (N_1376,In_1414,In_1571);
nor U1377 (N_1377,In_216,In_625);
xnor U1378 (N_1378,In_1571,In_1955);
nor U1379 (N_1379,In_849,In_1457);
nand U1380 (N_1380,In_1453,In_1126);
or U1381 (N_1381,In_1992,In_695);
nor U1382 (N_1382,In_1258,In_1448);
or U1383 (N_1383,In_730,In_412);
xor U1384 (N_1384,In_419,In_479);
xnor U1385 (N_1385,In_471,In_1347);
or U1386 (N_1386,In_178,In_1344);
or U1387 (N_1387,In_1017,In_367);
and U1388 (N_1388,In_1929,In_482);
and U1389 (N_1389,In_1170,In_1487);
or U1390 (N_1390,In_1683,In_34);
nand U1391 (N_1391,In_62,In_1210);
xor U1392 (N_1392,In_1344,In_1308);
nand U1393 (N_1393,In_1647,In_1234);
and U1394 (N_1394,In_1016,In_196);
nor U1395 (N_1395,In_1039,In_1508);
and U1396 (N_1396,In_700,In_1296);
or U1397 (N_1397,In_1939,In_923);
or U1398 (N_1398,In_742,In_854);
xor U1399 (N_1399,In_1053,In_771);
or U1400 (N_1400,In_971,In_1569);
nor U1401 (N_1401,In_1663,In_387);
xor U1402 (N_1402,In_1924,In_32);
xor U1403 (N_1403,In_341,In_1449);
nor U1404 (N_1404,In_1367,In_384);
or U1405 (N_1405,In_379,In_1106);
or U1406 (N_1406,In_465,In_1713);
and U1407 (N_1407,In_1027,In_194);
xnor U1408 (N_1408,In_1846,In_1077);
xor U1409 (N_1409,In_1127,In_862);
and U1410 (N_1410,In_203,In_1282);
nor U1411 (N_1411,In_22,In_124);
and U1412 (N_1412,In_1057,In_345);
or U1413 (N_1413,In_1216,In_172);
nor U1414 (N_1414,In_460,In_1044);
nand U1415 (N_1415,In_675,In_673);
nor U1416 (N_1416,In_1848,In_1213);
and U1417 (N_1417,In_1446,In_999);
or U1418 (N_1418,In_1381,In_1986);
nor U1419 (N_1419,In_467,In_285);
nand U1420 (N_1420,In_554,In_1058);
nand U1421 (N_1421,In_823,In_442);
nand U1422 (N_1422,In_1032,In_427);
nand U1423 (N_1423,In_882,In_1873);
nand U1424 (N_1424,In_1054,In_545);
xor U1425 (N_1425,In_483,In_890);
xor U1426 (N_1426,In_1451,In_538);
nor U1427 (N_1427,In_782,In_215);
nor U1428 (N_1428,In_578,In_1212);
nor U1429 (N_1429,In_1657,In_1920);
and U1430 (N_1430,In_907,In_1977);
xor U1431 (N_1431,In_782,In_1861);
nand U1432 (N_1432,In_1572,In_1134);
xor U1433 (N_1433,In_1920,In_1761);
or U1434 (N_1434,In_1234,In_115);
nor U1435 (N_1435,In_1028,In_25);
nand U1436 (N_1436,In_1279,In_708);
nand U1437 (N_1437,In_647,In_1820);
nand U1438 (N_1438,In_766,In_351);
nand U1439 (N_1439,In_1591,In_125);
and U1440 (N_1440,In_13,In_150);
nor U1441 (N_1441,In_361,In_522);
xnor U1442 (N_1442,In_931,In_1794);
nand U1443 (N_1443,In_79,In_1455);
nand U1444 (N_1444,In_696,In_1192);
or U1445 (N_1445,In_1107,In_1194);
or U1446 (N_1446,In_1624,In_991);
or U1447 (N_1447,In_1808,In_967);
or U1448 (N_1448,In_1871,In_1185);
and U1449 (N_1449,In_348,In_1706);
nor U1450 (N_1450,In_909,In_274);
nand U1451 (N_1451,In_518,In_537);
nor U1452 (N_1452,In_527,In_1257);
nor U1453 (N_1453,In_1766,In_1381);
and U1454 (N_1454,In_254,In_1371);
xnor U1455 (N_1455,In_1434,In_1772);
and U1456 (N_1456,In_1155,In_436);
nand U1457 (N_1457,In_387,In_1961);
xor U1458 (N_1458,In_1352,In_307);
xor U1459 (N_1459,In_641,In_1720);
and U1460 (N_1460,In_306,In_881);
and U1461 (N_1461,In_1277,In_722);
nand U1462 (N_1462,In_734,In_10);
or U1463 (N_1463,In_167,In_1276);
nor U1464 (N_1464,In_1232,In_1834);
nor U1465 (N_1465,In_783,In_851);
and U1466 (N_1466,In_1034,In_1841);
or U1467 (N_1467,In_973,In_1593);
and U1468 (N_1468,In_1957,In_1688);
or U1469 (N_1469,In_611,In_1221);
xnor U1470 (N_1470,In_827,In_1166);
nor U1471 (N_1471,In_390,In_425);
and U1472 (N_1472,In_1247,In_1020);
or U1473 (N_1473,In_465,In_635);
nand U1474 (N_1474,In_86,In_1582);
nand U1475 (N_1475,In_358,In_1769);
xor U1476 (N_1476,In_1566,In_1254);
nand U1477 (N_1477,In_343,In_1053);
or U1478 (N_1478,In_62,In_1967);
nand U1479 (N_1479,In_1246,In_327);
nor U1480 (N_1480,In_1489,In_42);
nor U1481 (N_1481,In_832,In_1496);
and U1482 (N_1482,In_265,In_295);
nand U1483 (N_1483,In_1964,In_325);
and U1484 (N_1484,In_1608,In_1974);
and U1485 (N_1485,In_291,In_1265);
nor U1486 (N_1486,In_1474,In_1118);
and U1487 (N_1487,In_1029,In_748);
nor U1488 (N_1488,In_1630,In_694);
nor U1489 (N_1489,In_346,In_745);
xor U1490 (N_1490,In_1367,In_1729);
and U1491 (N_1491,In_627,In_1105);
and U1492 (N_1492,In_848,In_116);
nor U1493 (N_1493,In_1969,In_72);
nand U1494 (N_1494,In_307,In_1912);
nor U1495 (N_1495,In_1287,In_718);
nor U1496 (N_1496,In_324,In_1816);
or U1497 (N_1497,In_1548,In_1784);
and U1498 (N_1498,In_689,In_315);
nand U1499 (N_1499,In_1646,In_1721);
and U1500 (N_1500,In_1934,In_210);
xor U1501 (N_1501,In_331,In_1181);
xor U1502 (N_1502,In_887,In_1023);
xor U1503 (N_1503,In_1092,In_758);
nor U1504 (N_1504,In_1887,In_663);
or U1505 (N_1505,In_1053,In_85);
nor U1506 (N_1506,In_1230,In_15);
and U1507 (N_1507,In_669,In_1042);
or U1508 (N_1508,In_238,In_721);
nand U1509 (N_1509,In_138,In_876);
or U1510 (N_1510,In_424,In_1130);
xor U1511 (N_1511,In_368,In_193);
nor U1512 (N_1512,In_1244,In_134);
xor U1513 (N_1513,In_1673,In_25);
and U1514 (N_1514,In_1297,In_1659);
xnor U1515 (N_1515,In_101,In_1285);
or U1516 (N_1516,In_601,In_1915);
xnor U1517 (N_1517,In_1185,In_239);
xor U1518 (N_1518,In_824,In_1523);
or U1519 (N_1519,In_1893,In_1804);
and U1520 (N_1520,In_409,In_743);
or U1521 (N_1521,In_1735,In_320);
nand U1522 (N_1522,In_168,In_1718);
and U1523 (N_1523,In_637,In_1310);
nand U1524 (N_1524,In_1761,In_1860);
nor U1525 (N_1525,In_1560,In_413);
nor U1526 (N_1526,In_529,In_1243);
nor U1527 (N_1527,In_1005,In_337);
nor U1528 (N_1528,In_1896,In_1960);
and U1529 (N_1529,In_1760,In_539);
xor U1530 (N_1530,In_714,In_833);
and U1531 (N_1531,In_2,In_1673);
xnor U1532 (N_1532,In_884,In_1188);
or U1533 (N_1533,In_1952,In_1193);
nand U1534 (N_1534,In_1005,In_1705);
xor U1535 (N_1535,In_1076,In_204);
and U1536 (N_1536,In_1830,In_964);
xnor U1537 (N_1537,In_359,In_1243);
and U1538 (N_1538,In_166,In_1042);
xnor U1539 (N_1539,In_934,In_602);
or U1540 (N_1540,In_7,In_1442);
nor U1541 (N_1541,In_1117,In_513);
nand U1542 (N_1542,In_1284,In_1979);
nand U1543 (N_1543,In_182,In_279);
and U1544 (N_1544,In_1647,In_1453);
or U1545 (N_1545,In_1796,In_1021);
nor U1546 (N_1546,In_1310,In_1182);
or U1547 (N_1547,In_1647,In_902);
and U1548 (N_1548,In_106,In_949);
nor U1549 (N_1549,In_1544,In_38);
nand U1550 (N_1550,In_1011,In_1850);
nor U1551 (N_1551,In_930,In_1797);
or U1552 (N_1552,In_1558,In_1194);
nor U1553 (N_1553,In_1101,In_489);
nor U1554 (N_1554,In_1551,In_982);
nor U1555 (N_1555,In_1716,In_368);
xnor U1556 (N_1556,In_1125,In_1489);
nor U1557 (N_1557,In_297,In_955);
or U1558 (N_1558,In_648,In_1986);
nand U1559 (N_1559,In_1218,In_549);
nor U1560 (N_1560,In_1099,In_1071);
or U1561 (N_1561,In_1759,In_738);
nor U1562 (N_1562,In_174,In_1558);
xor U1563 (N_1563,In_1296,In_229);
nor U1564 (N_1564,In_214,In_1695);
and U1565 (N_1565,In_1700,In_1679);
nor U1566 (N_1566,In_170,In_563);
xnor U1567 (N_1567,In_1733,In_681);
and U1568 (N_1568,In_1843,In_202);
and U1569 (N_1569,In_1034,In_701);
or U1570 (N_1570,In_1761,In_690);
xor U1571 (N_1571,In_1766,In_562);
and U1572 (N_1572,In_331,In_1634);
and U1573 (N_1573,In_1565,In_54);
or U1574 (N_1574,In_812,In_1351);
or U1575 (N_1575,In_1948,In_1674);
and U1576 (N_1576,In_279,In_248);
nor U1577 (N_1577,In_924,In_1128);
xor U1578 (N_1578,In_1327,In_1986);
nand U1579 (N_1579,In_782,In_781);
or U1580 (N_1580,In_454,In_1491);
or U1581 (N_1581,In_671,In_1947);
or U1582 (N_1582,In_472,In_1096);
and U1583 (N_1583,In_1855,In_62);
nor U1584 (N_1584,In_72,In_1871);
nand U1585 (N_1585,In_1597,In_754);
xnor U1586 (N_1586,In_1992,In_1809);
xor U1587 (N_1587,In_243,In_1072);
nand U1588 (N_1588,In_1739,In_355);
and U1589 (N_1589,In_1801,In_1197);
or U1590 (N_1590,In_914,In_1524);
nand U1591 (N_1591,In_1127,In_923);
and U1592 (N_1592,In_1096,In_573);
or U1593 (N_1593,In_378,In_1276);
xnor U1594 (N_1594,In_1754,In_844);
xor U1595 (N_1595,In_1784,In_177);
nor U1596 (N_1596,In_743,In_142);
and U1597 (N_1597,In_522,In_1676);
nand U1598 (N_1598,In_557,In_1032);
nand U1599 (N_1599,In_315,In_1305);
nand U1600 (N_1600,In_672,In_1696);
and U1601 (N_1601,In_1449,In_531);
xor U1602 (N_1602,In_1373,In_463);
xor U1603 (N_1603,In_736,In_195);
nand U1604 (N_1604,In_1390,In_743);
nor U1605 (N_1605,In_506,In_1476);
xnor U1606 (N_1606,In_1740,In_593);
or U1607 (N_1607,In_1646,In_413);
or U1608 (N_1608,In_1187,In_733);
nor U1609 (N_1609,In_461,In_163);
and U1610 (N_1610,In_1329,In_6);
xor U1611 (N_1611,In_1919,In_820);
nand U1612 (N_1612,In_790,In_1661);
or U1613 (N_1613,In_449,In_237);
and U1614 (N_1614,In_1990,In_19);
or U1615 (N_1615,In_1885,In_1038);
nor U1616 (N_1616,In_551,In_849);
and U1617 (N_1617,In_438,In_1098);
or U1618 (N_1618,In_29,In_494);
nand U1619 (N_1619,In_1474,In_846);
or U1620 (N_1620,In_137,In_1240);
nor U1621 (N_1621,In_1098,In_1256);
nand U1622 (N_1622,In_861,In_860);
and U1623 (N_1623,In_1877,In_1795);
nand U1624 (N_1624,In_650,In_1663);
nand U1625 (N_1625,In_227,In_1445);
and U1626 (N_1626,In_1123,In_587);
xnor U1627 (N_1627,In_988,In_890);
nand U1628 (N_1628,In_1784,In_787);
nand U1629 (N_1629,In_117,In_1959);
nor U1630 (N_1630,In_1794,In_679);
nor U1631 (N_1631,In_1390,In_201);
nand U1632 (N_1632,In_532,In_882);
or U1633 (N_1633,In_1851,In_91);
nand U1634 (N_1634,In_1999,In_1888);
or U1635 (N_1635,In_1953,In_582);
and U1636 (N_1636,In_821,In_1848);
xnor U1637 (N_1637,In_1785,In_678);
nand U1638 (N_1638,In_1095,In_1291);
and U1639 (N_1639,In_1517,In_365);
xnor U1640 (N_1640,In_973,In_1841);
nor U1641 (N_1641,In_1584,In_185);
xnor U1642 (N_1642,In_967,In_1734);
xor U1643 (N_1643,In_1525,In_688);
nand U1644 (N_1644,In_1777,In_98);
nor U1645 (N_1645,In_964,In_1542);
nand U1646 (N_1646,In_1532,In_1407);
and U1647 (N_1647,In_592,In_1694);
nor U1648 (N_1648,In_1213,In_1833);
or U1649 (N_1649,In_1809,In_1130);
nand U1650 (N_1650,In_579,In_761);
or U1651 (N_1651,In_1227,In_1351);
nor U1652 (N_1652,In_1718,In_1823);
nand U1653 (N_1653,In_1594,In_1660);
nand U1654 (N_1654,In_1427,In_1089);
nand U1655 (N_1655,In_304,In_1336);
and U1656 (N_1656,In_879,In_1532);
xnor U1657 (N_1657,In_1507,In_872);
or U1658 (N_1658,In_1942,In_883);
and U1659 (N_1659,In_1675,In_370);
xor U1660 (N_1660,In_1552,In_755);
xnor U1661 (N_1661,In_38,In_1715);
nor U1662 (N_1662,In_1724,In_1232);
xor U1663 (N_1663,In_1455,In_410);
and U1664 (N_1664,In_1587,In_481);
and U1665 (N_1665,In_911,In_1465);
and U1666 (N_1666,In_420,In_566);
nand U1667 (N_1667,In_1270,In_263);
and U1668 (N_1668,In_1362,In_394);
or U1669 (N_1669,In_192,In_411);
and U1670 (N_1670,In_1717,In_1542);
nor U1671 (N_1671,In_618,In_239);
or U1672 (N_1672,In_313,In_125);
nor U1673 (N_1673,In_635,In_434);
or U1674 (N_1674,In_1050,In_1140);
nor U1675 (N_1675,In_383,In_1329);
or U1676 (N_1676,In_759,In_1641);
xor U1677 (N_1677,In_225,In_1420);
nor U1678 (N_1678,In_1977,In_1288);
nor U1679 (N_1679,In_855,In_277);
nor U1680 (N_1680,In_1657,In_73);
nand U1681 (N_1681,In_152,In_824);
or U1682 (N_1682,In_1416,In_1654);
or U1683 (N_1683,In_1001,In_1165);
or U1684 (N_1684,In_1255,In_1278);
and U1685 (N_1685,In_1973,In_409);
xnor U1686 (N_1686,In_1331,In_1471);
nor U1687 (N_1687,In_710,In_552);
or U1688 (N_1688,In_909,In_1476);
or U1689 (N_1689,In_408,In_442);
xor U1690 (N_1690,In_1037,In_1502);
nand U1691 (N_1691,In_282,In_326);
and U1692 (N_1692,In_1588,In_429);
xnor U1693 (N_1693,In_886,In_1591);
nand U1694 (N_1694,In_1905,In_405);
and U1695 (N_1695,In_524,In_924);
nand U1696 (N_1696,In_1368,In_1966);
xor U1697 (N_1697,In_1013,In_1646);
and U1698 (N_1698,In_1144,In_1856);
xnor U1699 (N_1699,In_247,In_753);
nand U1700 (N_1700,In_236,In_634);
nand U1701 (N_1701,In_499,In_709);
nand U1702 (N_1702,In_823,In_1219);
or U1703 (N_1703,In_833,In_1707);
nor U1704 (N_1704,In_438,In_1161);
xor U1705 (N_1705,In_1948,In_1807);
xnor U1706 (N_1706,In_1006,In_988);
xor U1707 (N_1707,In_1033,In_1683);
or U1708 (N_1708,In_1825,In_550);
xor U1709 (N_1709,In_891,In_984);
or U1710 (N_1710,In_1607,In_1219);
nand U1711 (N_1711,In_1319,In_198);
nor U1712 (N_1712,In_838,In_1864);
nand U1713 (N_1713,In_662,In_169);
nor U1714 (N_1714,In_247,In_342);
xnor U1715 (N_1715,In_1976,In_1723);
nor U1716 (N_1716,In_1726,In_291);
nand U1717 (N_1717,In_1245,In_1812);
xor U1718 (N_1718,In_376,In_1490);
and U1719 (N_1719,In_222,In_1687);
nand U1720 (N_1720,In_227,In_1656);
and U1721 (N_1721,In_668,In_294);
xor U1722 (N_1722,In_882,In_1126);
nand U1723 (N_1723,In_904,In_417);
or U1724 (N_1724,In_1753,In_550);
nand U1725 (N_1725,In_680,In_1264);
nand U1726 (N_1726,In_1909,In_1569);
or U1727 (N_1727,In_185,In_1341);
or U1728 (N_1728,In_571,In_921);
and U1729 (N_1729,In_701,In_1492);
and U1730 (N_1730,In_1476,In_1754);
nand U1731 (N_1731,In_495,In_1386);
nand U1732 (N_1732,In_1475,In_1717);
nor U1733 (N_1733,In_1102,In_510);
nand U1734 (N_1734,In_1686,In_513);
nand U1735 (N_1735,In_1612,In_800);
nor U1736 (N_1736,In_353,In_13);
and U1737 (N_1737,In_155,In_928);
or U1738 (N_1738,In_373,In_1622);
xnor U1739 (N_1739,In_84,In_925);
and U1740 (N_1740,In_1634,In_1946);
or U1741 (N_1741,In_488,In_1870);
xnor U1742 (N_1742,In_1292,In_916);
nand U1743 (N_1743,In_1423,In_1943);
xor U1744 (N_1744,In_639,In_1390);
nor U1745 (N_1745,In_1676,In_1184);
nand U1746 (N_1746,In_602,In_1295);
and U1747 (N_1747,In_540,In_1983);
and U1748 (N_1748,In_770,In_1704);
nand U1749 (N_1749,In_1924,In_259);
nand U1750 (N_1750,In_755,In_1008);
or U1751 (N_1751,In_300,In_1559);
and U1752 (N_1752,In_1995,In_513);
nor U1753 (N_1753,In_106,In_849);
and U1754 (N_1754,In_902,In_61);
nor U1755 (N_1755,In_438,In_13);
nand U1756 (N_1756,In_385,In_1783);
xnor U1757 (N_1757,In_1347,In_1353);
or U1758 (N_1758,In_1388,In_1257);
or U1759 (N_1759,In_580,In_68);
nand U1760 (N_1760,In_82,In_675);
or U1761 (N_1761,In_1797,In_615);
and U1762 (N_1762,In_157,In_534);
xor U1763 (N_1763,In_1849,In_683);
and U1764 (N_1764,In_1573,In_913);
xor U1765 (N_1765,In_856,In_16);
nor U1766 (N_1766,In_1191,In_1814);
and U1767 (N_1767,In_1273,In_112);
xnor U1768 (N_1768,In_1335,In_1819);
nor U1769 (N_1769,In_3,In_1007);
and U1770 (N_1770,In_1510,In_1795);
nand U1771 (N_1771,In_784,In_537);
xnor U1772 (N_1772,In_1846,In_1211);
or U1773 (N_1773,In_847,In_550);
nand U1774 (N_1774,In_1130,In_1524);
or U1775 (N_1775,In_44,In_1186);
xor U1776 (N_1776,In_1274,In_480);
nand U1777 (N_1777,In_1487,In_1562);
nor U1778 (N_1778,In_313,In_950);
xor U1779 (N_1779,In_1315,In_248);
or U1780 (N_1780,In_1616,In_169);
xnor U1781 (N_1781,In_1616,In_287);
or U1782 (N_1782,In_426,In_1703);
or U1783 (N_1783,In_1149,In_1284);
nor U1784 (N_1784,In_1636,In_1398);
and U1785 (N_1785,In_1898,In_1611);
nand U1786 (N_1786,In_1364,In_1140);
nor U1787 (N_1787,In_168,In_675);
and U1788 (N_1788,In_1260,In_1304);
and U1789 (N_1789,In_834,In_246);
nor U1790 (N_1790,In_1920,In_1604);
or U1791 (N_1791,In_1588,In_1251);
xnor U1792 (N_1792,In_649,In_1054);
nor U1793 (N_1793,In_1584,In_351);
xnor U1794 (N_1794,In_833,In_842);
nor U1795 (N_1795,In_1131,In_989);
xor U1796 (N_1796,In_1628,In_1000);
and U1797 (N_1797,In_1649,In_412);
xnor U1798 (N_1798,In_1726,In_200);
nand U1799 (N_1799,In_1576,In_1403);
or U1800 (N_1800,In_445,In_1897);
nand U1801 (N_1801,In_388,In_470);
or U1802 (N_1802,In_1218,In_980);
and U1803 (N_1803,In_1781,In_515);
nand U1804 (N_1804,In_1835,In_1757);
nand U1805 (N_1805,In_1439,In_1270);
nand U1806 (N_1806,In_676,In_1484);
or U1807 (N_1807,In_1454,In_953);
and U1808 (N_1808,In_714,In_451);
or U1809 (N_1809,In_1940,In_254);
xnor U1810 (N_1810,In_1471,In_412);
or U1811 (N_1811,In_660,In_117);
nor U1812 (N_1812,In_1396,In_1242);
or U1813 (N_1813,In_838,In_852);
and U1814 (N_1814,In_1058,In_35);
and U1815 (N_1815,In_138,In_996);
and U1816 (N_1816,In_1371,In_1107);
nor U1817 (N_1817,In_220,In_1912);
nand U1818 (N_1818,In_137,In_1463);
or U1819 (N_1819,In_203,In_265);
nor U1820 (N_1820,In_1640,In_1412);
nand U1821 (N_1821,In_1420,In_844);
xnor U1822 (N_1822,In_1594,In_1430);
or U1823 (N_1823,In_1843,In_1282);
nor U1824 (N_1824,In_1971,In_1577);
or U1825 (N_1825,In_1578,In_1782);
xor U1826 (N_1826,In_296,In_1372);
and U1827 (N_1827,In_1074,In_1581);
or U1828 (N_1828,In_1053,In_858);
xnor U1829 (N_1829,In_1472,In_953);
and U1830 (N_1830,In_6,In_1499);
nand U1831 (N_1831,In_1242,In_585);
nor U1832 (N_1832,In_1621,In_1293);
or U1833 (N_1833,In_1860,In_198);
or U1834 (N_1834,In_377,In_1807);
and U1835 (N_1835,In_190,In_588);
nand U1836 (N_1836,In_25,In_963);
or U1837 (N_1837,In_1310,In_592);
nand U1838 (N_1838,In_161,In_1062);
nand U1839 (N_1839,In_741,In_1295);
xnor U1840 (N_1840,In_1501,In_1980);
nand U1841 (N_1841,In_660,In_922);
or U1842 (N_1842,In_615,In_1364);
xnor U1843 (N_1843,In_1382,In_1388);
nand U1844 (N_1844,In_205,In_1816);
xor U1845 (N_1845,In_840,In_410);
nand U1846 (N_1846,In_956,In_1420);
and U1847 (N_1847,In_1409,In_1987);
and U1848 (N_1848,In_1060,In_1019);
xnor U1849 (N_1849,In_1877,In_618);
and U1850 (N_1850,In_1462,In_1602);
xnor U1851 (N_1851,In_797,In_712);
nand U1852 (N_1852,In_1590,In_1830);
nand U1853 (N_1853,In_1242,In_1766);
and U1854 (N_1854,In_676,In_293);
nor U1855 (N_1855,In_935,In_767);
nand U1856 (N_1856,In_1679,In_1118);
nand U1857 (N_1857,In_1749,In_321);
nor U1858 (N_1858,In_493,In_572);
xnor U1859 (N_1859,In_92,In_1278);
and U1860 (N_1860,In_1868,In_1788);
nand U1861 (N_1861,In_968,In_90);
and U1862 (N_1862,In_883,In_419);
and U1863 (N_1863,In_1270,In_1654);
nor U1864 (N_1864,In_1438,In_1936);
and U1865 (N_1865,In_61,In_1583);
nor U1866 (N_1866,In_1327,In_460);
nor U1867 (N_1867,In_1659,In_276);
nor U1868 (N_1868,In_295,In_1630);
nor U1869 (N_1869,In_1755,In_1647);
and U1870 (N_1870,In_1749,In_1679);
nand U1871 (N_1871,In_611,In_1637);
nor U1872 (N_1872,In_1992,In_1030);
nor U1873 (N_1873,In_604,In_1739);
or U1874 (N_1874,In_451,In_1070);
and U1875 (N_1875,In_571,In_1703);
or U1876 (N_1876,In_1900,In_1167);
and U1877 (N_1877,In_1111,In_1914);
xor U1878 (N_1878,In_567,In_513);
nor U1879 (N_1879,In_347,In_490);
xnor U1880 (N_1880,In_1674,In_1210);
nor U1881 (N_1881,In_447,In_1887);
or U1882 (N_1882,In_629,In_346);
nor U1883 (N_1883,In_1366,In_830);
or U1884 (N_1884,In_429,In_1161);
xor U1885 (N_1885,In_1527,In_187);
nand U1886 (N_1886,In_1762,In_174);
xor U1887 (N_1887,In_174,In_478);
nand U1888 (N_1888,In_461,In_719);
nor U1889 (N_1889,In_962,In_1825);
or U1890 (N_1890,In_1851,In_1695);
and U1891 (N_1891,In_1755,In_230);
nor U1892 (N_1892,In_1522,In_1566);
or U1893 (N_1893,In_1238,In_1893);
nor U1894 (N_1894,In_1736,In_1437);
nand U1895 (N_1895,In_1120,In_111);
and U1896 (N_1896,In_1635,In_995);
nor U1897 (N_1897,In_322,In_1998);
nand U1898 (N_1898,In_1211,In_960);
nand U1899 (N_1899,In_776,In_1362);
nand U1900 (N_1900,In_1677,In_230);
nand U1901 (N_1901,In_1691,In_716);
xor U1902 (N_1902,In_863,In_1789);
and U1903 (N_1903,In_788,In_567);
xor U1904 (N_1904,In_1902,In_1941);
nand U1905 (N_1905,In_1229,In_762);
and U1906 (N_1906,In_545,In_1436);
and U1907 (N_1907,In_405,In_1193);
xnor U1908 (N_1908,In_188,In_671);
nand U1909 (N_1909,In_629,In_198);
nand U1910 (N_1910,In_739,In_238);
and U1911 (N_1911,In_1618,In_797);
and U1912 (N_1912,In_1523,In_419);
nor U1913 (N_1913,In_1298,In_1075);
and U1914 (N_1914,In_1284,In_1970);
nand U1915 (N_1915,In_1728,In_780);
or U1916 (N_1916,In_909,In_1494);
nor U1917 (N_1917,In_466,In_1702);
or U1918 (N_1918,In_584,In_1515);
xnor U1919 (N_1919,In_640,In_1237);
xnor U1920 (N_1920,In_151,In_1575);
nor U1921 (N_1921,In_14,In_1085);
nand U1922 (N_1922,In_1350,In_1601);
or U1923 (N_1923,In_1994,In_203);
nand U1924 (N_1924,In_71,In_204);
xnor U1925 (N_1925,In_1320,In_167);
and U1926 (N_1926,In_1558,In_1368);
or U1927 (N_1927,In_38,In_586);
and U1928 (N_1928,In_241,In_146);
and U1929 (N_1929,In_482,In_379);
nor U1930 (N_1930,In_1534,In_1778);
xnor U1931 (N_1931,In_365,In_1032);
nand U1932 (N_1932,In_574,In_301);
nor U1933 (N_1933,In_613,In_438);
or U1934 (N_1934,In_1915,In_1314);
or U1935 (N_1935,In_1102,In_823);
xor U1936 (N_1936,In_1469,In_1979);
nor U1937 (N_1937,In_1652,In_25);
xor U1938 (N_1938,In_231,In_1687);
nor U1939 (N_1939,In_67,In_761);
xor U1940 (N_1940,In_730,In_628);
nand U1941 (N_1941,In_1919,In_802);
and U1942 (N_1942,In_1714,In_82);
and U1943 (N_1943,In_55,In_1552);
nand U1944 (N_1944,In_322,In_1515);
or U1945 (N_1945,In_1527,In_1799);
and U1946 (N_1946,In_578,In_880);
and U1947 (N_1947,In_618,In_1622);
xor U1948 (N_1948,In_1568,In_1351);
or U1949 (N_1949,In_1724,In_55);
xor U1950 (N_1950,In_1697,In_1993);
xor U1951 (N_1951,In_1520,In_321);
or U1952 (N_1952,In_1780,In_1075);
xor U1953 (N_1953,In_1982,In_1580);
or U1954 (N_1954,In_1090,In_1601);
nor U1955 (N_1955,In_1023,In_1668);
and U1956 (N_1956,In_1637,In_1949);
xnor U1957 (N_1957,In_363,In_980);
nand U1958 (N_1958,In_163,In_1930);
nand U1959 (N_1959,In_1202,In_1722);
and U1960 (N_1960,In_1679,In_259);
or U1961 (N_1961,In_1064,In_435);
nand U1962 (N_1962,In_1376,In_144);
and U1963 (N_1963,In_160,In_113);
or U1964 (N_1964,In_1325,In_1639);
nor U1965 (N_1965,In_1231,In_1408);
nor U1966 (N_1966,In_688,In_839);
and U1967 (N_1967,In_1881,In_14);
nor U1968 (N_1968,In_1512,In_1189);
and U1969 (N_1969,In_573,In_1138);
xor U1970 (N_1970,In_1778,In_447);
xor U1971 (N_1971,In_1995,In_979);
or U1972 (N_1972,In_946,In_185);
xor U1973 (N_1973,In_1394,In_542);
and U1974 (N_1974,In_1281,In_1952);
or U1975 (N_1975,In_653,In_558);
or U1976 (N_1976,In_406,In_102);
or U1977 (N_1977,In_1932,In_893);
nor U1978 (N_1978,In_1438,In_1586);
nand U1979 (N_1979,In_283,In_1058);
or U1980 (N_1980,In_104,In_337);
xor U1981 (N_1981,In_1699,In_1702);
nand U1982 (N_1982,In_1676,In_1874);
or U1983 (N_1983,In_69,In_749);
nor U1984 (N_1984,In_1740,In_658);
and U1985 (N_1985,In_1385,In_922);
nor U1986 (N_1986,In_1128,In_1494);
or U1987 (N_1987,In_1303,In_1537);
nand U1988 (N_1988,In_1810,In_1666);
or U1989 (N_1989,In_294,In_204);
or U1990 (N_1990,In_379,In_1823);
and U1991 (N_1991,In_1536,In_469);
nor U1992 (N_1992,In_1856,In_1791);
xnor U1993 (N_1993,In_1062,In_1157);
xor U1994 (N_1994,In_982,In_962);
or U1995 (N_1995,In_467,In_811);
or U1996 (N_1996,In_289,In_783);
nand U1997 (N_1997,In_1215,In_1941);
xnor U1998 (N_1998,In_1565,In_1215);
and U1999 (N_1999,In_278,In_368);
and U2000 (N_2000,N_1982,N_615);
nand U2001 (N_2001,N_282,N_151);
and U2002 (N_2002,N_1902,N_727);
or U2003 (N_2003,N_477,N_1043);
or U2004 (N_2004,N_382,N_1145);
and U2005 (N_2005,N_1657,N_709);
xnor U2006 (N_2006,N_1614,N_1236);
and U2007 (N_2007,N_1883,N_105);
nor U2008 (N_2008,N_165,N_1223);
xor U2009 (N_2009,N_1068,N_867);
and U2010 (N_2010,N_770,N_1267);
and U2011 (N_2011,N_560,N_685);
nor U2012 (N_2012,N_1014,N_1460);
xor U2013 (N_2013,N_712,N_1035);
nand U2014 (N_2014,N_932,N_1978);
xnor U2015 (N_2015,N_1436,N_447);
or U2016 (N_2016,N_1893,N_296);
nor U2017 (N_2017,N_1767,N_844);
xnor U2018 (N_2018,N_622,N_1384);
nor U2019 (N_2019,N_1988,N_1316);
xnor U2020 (N_2020,N_1344,N_40);
nor U2021 (N_2021,N_1432,N_543);
nand U2022 (N_2022,N_723,N_1322);
nor U2023 (N_2023,N_1063,N_1134);
nor U2024 (N_2024,N_832,N_629);
and U2025 (N_2025,N_1163,N_1435);
or U2026 (N_2026,N_612,N_1601);
or U2027 (N_2027,N_1324,N_998);
nor U2028 (N_2028,N_547,N_1291);
nand U2029 (N_2029,N_1864,N_1470);
nor U2030 (N_2030,N_1418,N_1443);
nor U2031 (N_2031,N_1456,N_1559);
and U2032 (N_2032,N_1633,N_1830);
or U2033 (N_2033,N_850,N_780);
nor U2034 (N_2034,N_1345,N_371);
xnor U2035 (N_2035,N_12,N_1957);
nand U2036 (N_2036,N_191,N_1707);
nor U2037 (N_2037,N_1701,N_854);
and U2038 (N_2038,N_1116,N_529);
nand U2039 (N_2039,N_652,N_1403);
nor U2040 (N_2040,N_1503,N_640);
nand U2041 (N_2041,N_799,N_820);
and U2042 (N_2042,N_1030,N_1508);
and U2043 (N_2043,N_213,N_1581);
and U2044 (N_2044,N_696,N_455);
and U2045 (N_2045,N_1362,N_1187);
and U2046 (N_2046,N_931,N_933);
nor U2047 (N_2047,N_1142,N_1033);
nand U2048 (N_2048,N_1516,N_147);
xnor U2049 (N_2049,N_1064,N_753);
xnor U2050 (N_2050,N_194,N_9);
nor U2051 (N_2051,N_1549,N_504);
nand U2052 (N_2052,N_1492,N_199);
xnor U2053 (N_2053,N_107,N_620);
xor U2054 (N_2054,N_1476,N_1059);
nand U2055 (N_2055,N_1552,N_901);
and U2056 (N_2056,N_419,N_1620);
nor U2057 (N_2057,N_965,N_1929);
or U2058 (N_2058,N_1479,N_1792);
nor U2059 (N_2059,N_270,N_818);
or U2060 (N_2060,N_1130,N_1350);
nand U2061 (N_2061,N_76,N_83);
nor U2062 (N_2062,N_292,N_370);
nor U2063 (N_2063,N_1689,N_390);
and U2064 (N_2064,N_523,N_1832);
or U2065 (N_2065,N_877,N_956);
xnor U2066 (N_2066,N_995,N_689);
nor U2067 (N_2067,N_1222,N_861);
nor U2068 (N_2068,N_801,N_1773);
nor U2069 (N_2069,N_130,N_1131);
nand U2070 (N_2070,N_377,N_1625);
nand U2071 (N_2071,N_373,N_168);
and U2072 (N_2072,N_857,N_1061);
nor U2073 (N_2073,N_1193,N_954);
nor U2074 (N_2074,N_407,N_1320);
or U2075 (N_2075,N_1598,N_28);
xnor U2076 (N_2076,N_1986,N_1786);
xnor U2077 (N_2077,N_276,N_410);
and U2078 (N_2078,N_44,N_911);
nand U2079 (N_2079,N_1356,N_684);
or U2080 (N_2080,N_581,N_1167);
or U2081 (N_2081,N_866,N_1968);
nor U2082 (N_2082,N_1155,N_1090);
or U2083 (N_2083,N_298,N_680);
nand U2084 (N_2084,N_843,N_1154);
and U2085 (N_2085,N_1829,N_1042);
nand U2086 (N_2086,N_449,N_1333);
or U2087 (N_2087,N_1168,N_1989);
xnor U2088 (N_2088,N_120,N_608);
xor U2089 (N_2089,N_1106,N_895);
xnor U2090 (N_2090,N_495,N_1956);
or U2091 (N_2091,N_490,N_1218);
and U2092 (N_2092,N_1458,N_1279);
xor U2093 (N_2093,N_1727,N_1245);
and U2094 (N_2094,N_1232,N_720);
nor U2095 (N_2095,N_344,N_1780);
xor U2096 (N_2096,N_481,N_1983);
nand U2097 (N_2097,N_1138,N_1505);
nor U2098 (N_2098,N_334,N_133);
or U2099 (N_2099,N_1611,N_1381);
nand U2100 (N_2100,N_636,N_74);
nor U2101 (N_2101,N_1979,N_862);
and U2102 (N_2102,N_1740,N_891);
xor U2103 (N_2103,N_1778,N_84);
or U2104 (N_2104,N_1367,N_1238);
or U2105 (N_2105,N_457,N_1874);
nand U2106 (N_2106,N_1490,N_1056);
nor U2107 (N_2107,N_602,N_453);
nor U2108 (N_2108,N_324,N_1420);
or U2109 (N_2109,N_1817,N_626);
or U2110 (N_2110,N_531,N_450);
and U2111 (N_2111,N_916,N_331);
nor U2112 (N_2112,N_1317,N_678);
nor U2113 (N_2113,N_628,N_573);
xnor U2114 (N_2114,N_971,N_1634);
and U2115 (N_2115,N_150,N_880);
or U2116 (N_2116,N_1535,N_217);
and U2117 (N_2117,N_722,N_1920);
nor U2118 (N_2118,N_214,N_1724);
nor U2119 (N_2119,N_119,N_472);
or U2120 (N_2120,N_1734,N_915);
xnor U2121 (N_2121,N_1579,N_1121);
and U2122 (N_2122,N_1797,N_108);
and U2123 (N_2123,N_1020,N_1784);
nand U2124 (N_2124,N_1843,N_1307);
nor U2125 (N_2125,N_632,N_1569);
or U2126 (N_2126,N_1256,N_1966);
and U2127 (N_2127,N_238,N_1704);
nand U2128 (N_2128,N_1336,N_333);
nand U2129 (N_2129,N_17,N_1233);
nor U2130 (N_2130,N_614,N_922);
or U2131 (N_2131,N_1450,N_555);
nor U2132 (N_2132,N_1449,N_658);
xor U2133 (N_2133,N_1177,N_1866);
xor U2134 (N_2134,N_374,N_483);
nand U2135 (N_2135,N_461,N_1998);
xor U2136 (N_2136,N_22,N_823);
and U2137 (N_2137,N_1757,N_1198);
nor U2138 (N_2138,N_1143,N_834);
nand U2139 (N_2139,N_772,N_1802);
nand U2140 (N_2140,N_1854,N_175);
and U2141 (N_2141,N_397,N_185);
or U2142 (N_2142,N_819,N_91);
nand U2143 (N_2143,N_750,N_353);
xnor U2144 (N_2144,N_323,N_1082);
xor U2145 (N_2145,N_1749,N_767);
or U2146 (N_2146,N_766,N_1609);
and U2147 (N_2147,N_928,N_1621);
nor U2148 (N_2148,N_1343,N_577);
xnor U2149 (N_2149,N_777,N_209);
and U2150 (N_2150,N_283,N_365);
nor U2151 (N_2151,N_1885,N_1045);
or U2152 (N_2152,N_475,N_1523);
nand U2153 (N_2153,N_1341,N_790);
and U2154 (N_2154,N_1103,N_1700);
or U2155 (N_2155,N_921,N_502);
and U2156 (N_2156,N_786,N_1354);
xnor U2157 (N_2157,N_1007,N_1884);
nor U2158 (N_2158,N_75,N_118);
nor U2159 (N_2159,N_1246,N_386);
and U2160 (N_2160,N_1386,N_812);
and U2161 (N_2161,N_436,N_1921);
and U2162 (N_2162,N_853,N_1050);
xor U2163 (N_2163,N_35,N_1464);
and U2164 (N_2164,N_1448,N_984);
xnor U2165 (N_2165,N_1809,N_400);
or U2166 (N_2166,N_1735,N_317);
nor U2167 (N_2167,N_788,N_1912);
nor U2168 (N_2168,N_380,N_1995);
or U2169 (N_2169,N_73,N_856);
xor U2170 (N_2170,N_1889,N_215);
and U2171 (N_2171,N_1109,N_286);
nand U2172 (N_2172,N_1877,N_439);
nand U2173 (N_2173,N_1655,N_1563);
xor U2174 (N_2174,N_198,N_879);
nand U2175 (N_2175,N_1416,N_960);
xnor U2176 (N_2176,N_1152,N_166);
nand U2177 (N_2177,N_1880,N_917);
nand U2178 (N_2178,N_1406,N_1365);
nand U2179 (N_2179,N_1895,N_19);
or U2180 (N_2180,N_695,N_1065);
nand U2181 (N_2181,N_1954,N_739);
nand U2182 (N_2182,N_875,N_228);
and U2183 (N_2183,N_1610,N_944);
nor U2184 (N_2184,N_1274,N_1718);
nand U2185 (N_2185,N_1815,N_1251);
or U2186 (N_2186,N_332,N_18);
and U2187 (N_2187,N_563,N_508);
or U2188 (N_2188,N_1841,N_1157);
nor U2189 (N_2189,N_1188,N_113);
and U2190 (N_2190,N_1544,N_237);
nor U2191 (N_2191,N_1328,N_546);
xnor U2192 (N_2192,N_1916,N_797);
or U2193 (N_2193,N_466,N_1574);
xor U2194 (N_2194,N_654,N_905);
nand U2195 (N_2195,N_1099,N_184);
and U2196 (N_2196,N_699,N_51);
or U2197 (N_2197,N_1126,N_236);
and U2198 (N_2198,N_1713,N_972);
or U2199 (N_2199,N_576,N_1339);
nand U2200 (N_2200,N_366,N_1482);
nand U2201 (N_2201,N_1237,N_242);
nor U2202 (N_2202,N_1278,N_735);
or U2203 (N_2203,N_463,N_1510);
xor U2204 (N_2204,N_1419,N_1340);
nand U2205 (N_2205,N_381,N_210);
or U2206 (N_2206,N_1473,N_517);
nand U2207 (N_2207,N_258,N_160);
and U2208 (N_2208,N_605,N_886);
xnor U2209 (N_2209,N_499,N_756);
and U2210 (N_2210,N_1779,N_1720);
xor U2211 (N_2211,N_312,N_1536);
or U2212 (N_2212,N_146,N_262);
xor U2213 (N_2213,N_48,N_1211);
nand U2214 (N_2214,N_661,N_945);
nor U2215 (N_2215,N_1684,N_1863);
xnor U2216 (N_2216,N_1851,N_122);
nand U2217 (N_2217,N_460,N_465);
and U2218 (N_2218,N_761,N_1692);
and U2219 (N_2219,N_1423,N_1617);
nor U2220 (N_2220,N_1129,N_1695);
nor U2221 (N_2221,N_1015,N_1359);
nor U2222 (N_2222,N_1772,N_47);
and U2223 (N_2223,N_1886,N_322);
nor U2224 (N_2224,N_746,N_1133);
xnor U2225 (N_2225,N_538,N_1243);
nand U2226 (N_2226,N_230,N_1537);
or U2227 (N_2227,N_686,N_1387);
xor U2228 (N_2228,N_1839,N_1694);
xnor U2229 (N_2229,N_1319,N_1346);
or U2230 (N_2230,N_550,N_526);
and U2231 (N_2231,N_1461,N_1970);
nand U2232 (N_2232,N_205,N_1010);
or U2233 (N_2233,N_976,N_1687);
xor U2234 (N_2234,N_142,N_1628);
or U2235 (N_2235,N_1946,N_1967);
and U2236 (N_2236,N_4,N_343);
xnor U2237 (N_2237,N_707,N_1931);
nand U2238 (N_2238,N_1214,N_1870);
nand U2239 (N_2239,N_422,N_702);
nand U2240 (N_2240,N_1375,N_1029);
nand U2241 (N_2241,N_434,N_432);
nor U2242 (N_2242,N_1545,N_1011);
nor U2243 (N_2243,N_1977,N_1051);
nor U2244 (N_2244,N_1244,N_1891);
xnor U2245 (N_2245,N_471,N_816);
nand U2246 (N_2246,N_1226,N_1395);
or U2247 (N_2247,N_849,N_631);
or U2248 (N_2248,N_1626,N_32);
and U2249 (N_2249,N_768,N_571);
xor U2250 (N_2250,N_1485,N_327);
or U2251 (N_2251,N_528,N_473);
and U2252 (N_2252,N_1148,N_25);
or U2253 (N_2253,N_1558,N_584);
nand U2254 (N_2254,N_745,N_817);
nand U2255 (N_2255,N_1021,N_551);
nor U2256 (N_2256,N_1093,N_683);
nand U2257 (N_2257,N_1282,N_1737);
and U2258 (N_2258,N_1721,N_868);
or U2259 (N_2259,N_1229,N_212);
and U2260 (N_2260,N_649,N_749);
nor U2261 (N_2261,N_46,N_294);
nand U2262 (N_2262,N_394,N_938);
nand U2263 (N_2263,N_1589,N_603);
nand U2264 (N_2264,N_1927,N_355);
xnor U2265 (N_2265,N_694,N_1108);
xnor U2266 (N_2266,N_1202,N_1997);
nand U2267 (N_2267,N_741,N_549);
nand U2268 (N_2268,N_1821,N_800);
xnor U2269 (N_2269,N_1981,N_1225);
or U2270 (N_2270,N_804,N_598);
and U2271 (N_2271,N_1411,N_1994);
xnor U2272 (N_2272,N_1452,N_1373);
and U2273 (N_2273,N_653,N_1196);
or U2274 (N_2274,N_1046,N_306);
xor U2275 (N_2275,N_1642,N_315);
and U2276 (N_2276,N_1437,N_0);
xnor U2277 (N_2277,N_1331,N_1622);
nor U2278 (N_2278,N_186,N_1658);
xor U2279 (N_2279,N_257,N_117);
or U2280 (N_2280,N_493,N_1216);
nor U2281 (N_2281,N_1496,N_145);
nand U2282 (N_2282,N_1872,N_1442);
or U2283 (N_2283,N_1421,N_906);
nand U2284 (N_2284,N_1629,N_1999);
nand U2285 (N_2285,N_1417,N_997);
nand U2286 (N_2286,N_89,N_1774);
xor U2287 (N_2287,N_218,N_641);
nor U2288 (N_2288,N_1383,N_656);
nand U2289 (N_2289,N_1299,N_41);
and U2290 (N_2290,N_1867,N_1984);
nor U2291 (N_2291,N_1819,N_95);
xnor U2292 (N_2292,N_273,N_1190);
nand U2293 (N_2293,N_1572,N_1494);
and U2294 (N_2294,N_926,N_744);
nand U2295 (N_2295,N_1665,N_607);
nand U2296 (N_2296,N_1399,N_1078);
nor U2297 (N_2297,N_1682,N_530);
and U2298 (N_2298,N_1451,N_1207);
xnor U2299 (N_2299,N_1221,N_1660);
xor U2300 (N_2300,N_527,N_1673);
xor U2301 (N_2301,N_356,N_635);
nor U2302 (N_2302,N_1650,N_1052);
and U2303 (N_2303,N_1358,N_1105);
nand U2304 (N_2304,N_359,N_525);
and U2305 (N_2305,N_1186,N_710);
and U2306 (N_2306,N_587,N_1112);
or U2307 (N_2307,N_1087,N_1044);
or U2308 (N_2308,N_263,N_1702);
nor U2309 (N_2309,N_1446,N_1659);
xnor U2310 (N_2310,N_1349,N_1976);
and U2311 (N_2311,N_1288,N_624);
xor U2312 (N_2312,N_458,N_1250);
xnor U2313 (N_2313,N_1260,N_618);
nand U2314 (N_2314,N_1493,N_1264);
and U2315 (N_2315,N_1812,N_250);
or U2316 (N_2316,N_1026,N_301);
or U2317 (N_2317,N_303,N_604);
xor U2318 (N_2318,N_1136,N_1258);
and U2319 (N_2319,N_398,N_1235);
nand U2320 (N_2320,N_893,N_1661);
or U2321 (N_2321,N_31,N_1756);
or U2322 (N_2322,N_1636,N_609);
xnor U2323 (N_2323,N_1228,N_63);
and U2324 (N_2324,N_348,N_672);
or U2325 (N_2325,N_1876,N_364);
nand U2326 (N_2326,N_1807,N_1615);
and U2327 (N_2327,N_106,N_1306);
and U2328 (N_2328,N_53,N_1725);
nor U2329 (N_2329,N_1638,N_743);
xnor U2330 (N_2330,N_590,N_1783);
nor U2331 (N_2331,N_1987,N_1040);
and U2332 (N_2332,N_1666,N_1888);
or U2333 (N_2333,N_1135,N_402);
nand U2334 (N_2334,N_994,N_1798);
and U2335 (N_2335,N_88,N_887);
nor U2336 (N_2336,N_1781,N_408);
nand U2337 (N_2337,N_77,N_562);
nand U2338 (N_2338,N_56,N_201);
xnor U2339 (N_2339,N_831,N_548);
xnor U2340 (N_2340,N_1879,N_1653);
or U2341 (N_2341,N_1468,N_281);
nor U2342 (N_2342,N_58,N_1507);
xnor U2343 (N_2343,N_1215,N_698);
nand U2344 (N_2344,N_1810,N_1670);
nand U2345 (N_2345,N_503,N_321);
and U2346 (N_2346,N_1486,N_96);
nor U2347 (N_2347,N_1431,N_894);
or U2348 (N_2348,N_583,N_1089);
xnor U2349 (N_2349,N_93,N_1624);
or U2350 (N_2350,N_1820,N_623);
nor U2351 (N_2351,N_1060,N_1481);
xor U2352 (N_2352,N_657,N_1826);
and U2353 (N_2353,N_486,N_290);
xor U2354 (N_2354,N_715,N_1709);
or U2355 (N_2355,N_101,N_542);
xnor U2356 (N_2356,N_1407,N_884);
nor U2357 (N_2357,N_521,N_757);
nand U2358 (N_2358,N_260,N_1677);
xnor U2359 (N_2359,N_769,N_1938);
or U2360 (N_2360,N_470,N_898);
xor U2361 (N_2361,N_1122,N_1227);
and U2362 (N_2362,N_1396,N_835);
nand U2363 (N_2363,N_919,N_1019);
and U2364 (N_2364,N_372,N_1933);
xnor U2365 (N_2365,N_480,N_1500);
nor U2366 (N_2366,N_1438,N_229);
xor U2367 (N_2367,N_115,N_1645);
nor U2368 (N_2368,N_1806,N_29);
and U2369 (N_2369,N_78,N_1348);
xnor U2370 (N_2370,N_1801,N_600);
and U2371 (N_2371,N_703,N_1255);
and U2372 (N_2372,N_1374,N_1849);
nor U2373 (N_2373,N_10,N_224);
nor U2374 (N_2374,N_1393,N_1489);
nor U2375 (N_2375,N_1220,N_968);
xnor U2376 (N_2376,N_38,N_1000);
or U2377 (N_2377,N_586,N_822);
or U2378 (N_2378,N_1147,N_1965);
nand U2379 (N_2379,N_392,N_1858);
nor U2380 (N_2380,N_1269,N_1003);
and U2381 (N_2381,N_54,N_388);
nand U2382 (N_2382,N_37,N_1647);
nand U2383 (N_2383,N_1942,N_1234);
or U2384 (N_2384,N_1771,N_1961);
and U2385 (N_2385,N_411,N_474);
nand U2386 (N_2386,N_742,N_520);
nor U2387 (N_2387,N_1459,N_1539);
nand U2388 (N_2388,N_318,N_1799);
nand U2389 (N_2389,N_1445,N_1730);
and U2390 (N_2390,N_1791,N_1731);
nand U2391 (N_2391,N_729,N_1049);
xnor U2392 (N_2392,N_248,N_1074);
nand U2393 (N_2393,N_863,N_1372);
xnor U2394 (N_2394,N_1913,N_1275);
nand U2395 (N_2395,N_1491,N_650);
xnor U2396 (N_2396,N_287,N_183);
or U2397 (N_2397,N_1675,N_1554);
nor U2398 (N_2398,N_103,N_445);
xnor U2399 (N_2399,N_1032,N_1753);
xor U2400 (N_2400,N_255,N_732);
nor U2401 (N_2401,N_143,N_665);
or U2402 (N_2402,N_924,N_125);
xnor U2403 (N_2403,N_1910,N_98);
and U2404 (N_2404,N_1656,N_1189);
xor U2405 (N_2405,N_1855,N_1137);
xnor U2406 (N_2406,N_50,N_1915);
and U2407 (N_2407,N_279,N_1975);
xor U2408 (N_2408,N_99,N_1295);
nor U2409 (N_2409,N_265,N_264);
nand U2410 (N_2410,N_363,N_606);
or U2411 (N_2411,N_713,N_1006);
xor U2412 (N_2412,N_81,N_983);
xnor U2413 (N_2413,N_939,N_1334);
and U2414 (N_2414,N_1919,N_429);
nand U2415 (N_2415,N_1859,N_779);
or U2416 (N_2416,N_1887,N_1414);
or U2417 (N_2417,N_1405,N_240);
xnor U2418 (N_2418,N_759,N_1277);
nor U2419 (N_2419,N_1591,N_269);
and U2420 (N_2420,N_482,N_1146);
nor U2421 (N_2421,N_467,N_1752);
nand U2422 (N_2422,N_1909,N_1648);
and U2423 (N_2423,N_1101,N_711);
nand U2424 (N_2424,N_1321,N_1848);
xor U2425 (N_2425,N_846,N_929);
or U2426 (N_2426,N_1497,N_266);
or U2427 (N_2427,N_1602,N_302);
or U2428 (N_2428,N_1805,N_487);
nor U2429 (N_2429,N_452,N_1002);
nor U2430 (N_2430,N_1833,N_319);
or U2431 (N_2431,N_1197,N_1896);
xor U2432 (N_2432,N_1018,N_1422);
and U2433 (N_2433,N_676,N_778);
xnor U2434 (N_2434,N_825,N_736);
or U2435 (N_2435,N_1878,N_1242);
and U2436 (N_2436,N_1769,N_599);
nor U2437 (N_2437,N_986,N_501);
nand U2438 (N_2438,N_1203,N_152);
and U2439 (N_2439,N_1041,N_578);
or U2440 (N_2440,N_1310,N_308);
nand U2441 (N_2441,N_881,N_1415);
and U2442 (N_2442,N_1294,N_1787);
xor U2443 (N_2443,N_1327,N_902);
or U2444 (N_2444,N_1009,N_1838);
nor U2445 (N_2445,N_1795,N_347);
nor U2446 (N_2446,N_64,N_1499);
nor U2447 (N_2447,N_936,N_1290);
xor U2448 (N_2448,N_104,N_1715);
nand U2449 (N_2449,N_488,N_1576);
nand U2450 (N_2450,N_1114,N_651);
or U2451 (N_2451,N_1249,N_1127);
and U2452 (N_2452,N_1181,N_1153);
or U2453 (N_2453,N_1522,N_1538);
or U2454 (N_2454,N_498,N_1678);
and U2455 (N_2455,N_907,N_459);
or U2456 (N_2456,N_163,N_341);
and U2457 (N_2457,N_62,N_1487);
nor U2458 (N_2458,N_771,N_655);
nor U2459 (N_2459,N_1401,N_1651);
nand U2460 (N_2460,N_339,N_1325);
or U2461 (N_2461,N_580,N_1710);
or U2462 (N_2462,N_1219,N_1330);
nand U2463 (N_2463,N_1712,N_889);
or U2464 (N_2464,N_1828,N_1604);
nand U2465 (N_2465,N_1788,N_1113);
or U2466 (N_2466,N_1212,N_764);
nor U2467 (N_2467,N_848,N_1366);
or U2468 (N_2468,N_513,N_1398);
nor U2469 (N_2469,N_337,N_216);
and U2470 (N_2470,N_162,N_1547);
nand U2471 (N_2471,N_838,N_914);
nor U2472 (N_2472,N_588,N_518);
and U2473 (N_2473,N_1402,N_506);
nor U2474 (N_2474,N_11,N_534);
and U2475 (N_2475,N_1462,N_1501);
xor U2476 (N_2476,N_593,N_730);
and U2477 (N_2477,N_1681,N_313);
xor U2478 (N_2478,N_663,N_26);
xnor U2479 (N_2479,N_845,N_1760);
xor U2480 (N_2480,N_338,N_1900);
nand U2481 (N_2481,N_1038,N_20);
nor U2482 (N_2482,N_991,N_1498);
xor U2483 (N_2483,N_23,N_1557);
and U2484 (N_2484,N_393,N_52);
or U2485 (N_2485,N_1400,N_885);
nand U2486 (N_2486,N_329,N_721);
nor U2487 (N_2487,N_579,N_1945);
and U2488 (N_2488,N_1081,N_802);
xor U2489 (N_2489,N_1281,N_1166);
or U2490 (N_2490,N_784,N_1764);
nand U2491 (N_2491,N_1635,N_1066);
nand U2492 (N_2492,N_1048,N_1315);
xnor U2493 (N_2493,N_1397,N_1102);
or U2494 (N_2494,N_1488,N_454);
and U2495 (N_2495,N_564,N_934);
nor U2496 (N_2496,N_172,N_85);
and U2497 (N_2497,N_575,N_1191);
xnor U2498 (N_2498,N_1567,N_33);
or U2499 (N_2499,N_140,N_1616);
nand U2500 (N_2500,N_1388,N_1164);
nand U2501 (N_2501,N_1901,N_137);
nand U2502 (N_2502,N_1241,N_1054);
nor U2503 (N_2503,N_648,N_154);
and U2504 (N_2504,N_1844,N_187);
xnor U2505 (N_2505,N_1894,N_1096);
or U2506 (N_2506,N_1690,N_384);
and U2507 (N_2507,N_1263,N_1286);
nor U2508 (N_2508,N_1741,N_1782);
and U2509 (N_2509,N_14,N_1951);
nand U2510 (N_2510,N_874,N_1016);
and U2511 (N_2511,N_1284,N_1326);
or U2512 (N_2512,N_307,N_1719);
nor U2513 (N_2513,N_1176,N_342);
nand U2514 (N_2514,N_491,N_1025);
and U2515 (N_2515,N_1930,N_49);
xor U2516 (N_2516,N_837,N_1526);
and U2517 (N_2517,N_990,N_1162);
nand U2518 (N_2518,N_708,N_1253);
or U2519 (N_2519,N_793,N_174);
xor U2520 (N_2520,N_1012,N_196);
or U2521 (N_2521,N_1079,N_1144);
nor U2522 (N_2522,N_737,N_139);
or U2523 (N_2523,N_978,N_1845);
nand U2524 (N_2524,N_775,N_541);
nand U2525 (N_2525,N_985,N_1935);
nand U2526 (N_2526,N_1342,N_1963);
or U2527 (N_2527,N_1751,N_1644);
and U2528 (N_2528,N_1693,N_507);
xor U2529 (N_2529,N_336,N_829);
nand U2530 (N_2530,N_1502,N_1847);
or U2531 (N_2531,N_1672,N_442);
nand U2532 (N_2532,N_256,N_167);
nand U2533 (N_2533,N_1355,N_1761);
nand U2534 (N_2534,N_690,N_1297);
and U2535 (N_2535,N_1301,N_1204);
nor U2536 (N_2536,N_1905,N_1776);
or U2537 (N_2537,N_225,N_1180);
nand U2538 (N_2538,N_958,N_677);
nor U2539 (N_2539,N_1639,N_72);
nor U2540 (N_2540,N_222,N_539);
and U2541 (N_2541,N_957,N_1053);
nor U2542 (N_2542,N_616,N_153);
or U2543 (N_2543,N_70,N_1904);
xor U2544 (N_2544,N_1723,N_1871);
or U2545 (N_2545,N_668,N_430);
nor U2546 (N_2546,N_1231,N_582);
nand U2547 (N_2547,N_1314,N_1717);
nor U2548 (N_2548,N_328,N_1903);
nor U2549 (N_2549,N_1513,N_1364);
nor U2550 (N_2550,N_1150,N_36);
xor U2551 (N_2551,N_252,N_1941);
and U2552 (N_2552,N_1674,N_763);
xnor U2553 (N_2553,N_155,N_638);
xnor U2554 (N_2554,N_1834,N_869);
and U2555 (N_2555,N_65,N_1803);
and U2556 (N_2556,N_937,N_385);
and U2557 (N_2557,N_842,N_1151);
nor U2558 (N_2558,N_1506,N_289);
and U2559 (N_2559,N_1543,N_1627);
nor U2560 (N_2560,N_1914,N_1943);
nor U2561 (N_2561,N_1816,N_1156);
and U2562 (N_2562,N_21,N_1923);
or U2563 (N_2563,N_435,N_533);
or U2564 (N_2564,N_613,N_462);
xnor U2565 (N_2565,N_717,N_963);
xor U2566 (N_2566,N_1969,N_1382);
nand U2567 (N_2567,N_1329,N_1512);
and U2568 (N_2568,N_500,N_141);
nand U2569 (N_2569,N_320,N_989);
and U2570 (N_2570,N_219,N_1571);
or U2571 (N_2571,N_941,N_5);
nand U2572 (N_2572,N_949,N_409);
xor U2573 (N_2573,N_1313,N_1534);
and U2574 (N_2574,N_27,N_272);
nor U2575 (N_2575,N_833,N_512);
nor U2576 (N_2576,N_316,N_693);
and U2577 (N_2577,N_387,N_660);
nand U2578 (N_2578,N_1770,N_293);
and U2579 (N_2579,N_1555,N_1261);
xnor U2580 (N_2580,N_157,N_1560);
xor U2581 (N_2581,N_1729,N_1743);
xor U2582 (N_2582,N_952,N_311);
or U2583 (N_2583,N_200,N_828);
or U2584 (N_2584,N_1599,N_1484);
nand U2585 (N_2585,N_627,N_478);
nand U2586 (N_2586,N_805,N_1711);
and U2587 (N_2587,N_1224,N_1069);
xor U2588 (N_2588,N_1822,N_1098);
nor U2589 (N_2589,N_1521,N_433);
xor U2590 (N_2590,N_1254,N_1973);
or U2591 (N_2591,N_494,N_559);
or U2592 (N_2592,N_1055,N_79);
nor U2593 (N_2593,N_871,N_1793);
nor U2594 (N_2594,N_299,N_1862);
and U2595 (N_2595,N_1922,N_948);
xnor U2596 (N_2596,N_1952,N_813);
or U2597 (N_2597,N_1305,N_803);
xnor U2598 (N_2598,N_159,N_275);
and U2599 (N_2599,N_417,N_92);
nand U2600 (N_2600,N_1149,N_232);
nor U2601 (N_2601,N_1027,N_1210);
and U2602 (N_2602,N_1944,N_1519);
or U2603 (N_2603,N_1262,N_807);
nor U2604 (N_2604,N_673,N_1296);
and U2605 (N_2605,N_345,N_135);
or U2606 (N_2606,N_992,N_30);
or U2607 (N_2607,N_247,N_1239);
and U2608 (N_2608,N_918,N_1777);
or U2609 (N_2609,N_1183,N_1654);
or U2610 (N_2610,N_1906,N_1947);
nor U2611 (N_2611,N_1104,N_389);
xor U2612 (N_2612,N_1426,N_1062);
nor U2613 (N_2613,N_540,N_1705);
nand U2614 (N_2614,N_516,N_1008);
and U2615 (N_2615,N_116,N_1107);
nand U2616 (N_2616,N_795,N_271);
nor U2617 (N_2617,N_1824,N_1159);
nand U2618 (N_2618,N_127,N_1580);
or U2619 (N_2619,N_1568,N_1039);
or U2620 (N_2620,N_1111,N_1643);
nor U2621 (N_2621,N_1527,N_897);
xnor U2622 (N_2622,N_1562,N_231);
and U2623 (N_2623,N_1257,N_1308);
nand U2624 (N_2624,N_558,N_734);
xnor U2625 (N_2625,N_725,N_1533);
nand U2626 (N_2626,N_1934,N_57);
or U2627 (N_2627,N_1869,N_621);
nand U2628 (N_2628,N_1283,N_278);
or U2629 (N_2629,N_190,N_565);
nor U2630 (N_2630,N_794,N_892);
or U2631 (N_2631,N_357,N_1899);
nor U2632 (N_2632,N_68,N_1165);
nand U2633 (N_2633,N_1515,N_953);
or U2634 (N_2634,N_1641,N_1285);
or U2635 (N_2635,N_112,N_1679);
or U2636 (N_2636,N_1022,N_351);
or U2637 (N_2637,N_126,N_1206);
and U2638 (N_2638,N_444,N_688);
and U2639 (N_2639,N_404,N_376);
nand U2640 (N_2640,N_1077,N_1683);
xor U2641 (N_2641,N_304,N_1950);
nor U2642 (N_2642,N_1668,N_1584);
nor U2643 (N_2643,N_1747,N_241);
xnor U2644 (N_2644,N_1953,N_1875);
and U2645 (N_2645,N_251,N_1857);
and U2646 (N_2646,N_1971,N_675);
nor U2647 (N_2647,N_1408,N_1608);
xnor U2648 (N_2648,N_979,N_999);
xor U2649 (N_2649,N_1546,N_509);
and U2650 (N_2650,N_239,N_1471);
nor U2651 (N_2651,N_1357,N_925);
nand U2652 (N_2652,N_1728,N_596);
xnor U2653 (N_2653,N_920,N_1831);
or U2654 (N_2654,N_1005,N_1664);
and U2655 (N_2655,N_589,N_1467);
nand U2656 (N_2656,N_1955,N_1881);
or U2657 (N_2657,N_1890,N_585);
nand U2658 (N_2658,N_1575,N_601);
or U2659 (N_2659,N_246,N_1477);
nand U2660 (N_2660,N_1413,N_1287);
xnor U2661 (N_2661,N_1265,N_361);
nor U2662 (N_2662,N_1818,N_959);
or U2663 (N_2663,N_1175,N_208);
nor U2664 (N_2664,N_687,N_1091);
and U2665 (N_2665,N_760,N_416);
nor U2666 (N_2666,N_1630,N_630);
nor U2667 (N_2667,N_1266,N_738);
nor U2668 (N_2668,N_1835,N_1972);
xnor U2669 (N_2669,N_642,N_497);
nor U2670 (N_2670,N_1303,N_1140);
or U2671 (N_2671,N_354,N_977);
nor U2672 (N_2672,N_443,N_1304);
nand U2673 (N_2673,N_277,N_1474);
nand U2674 (N_2674,N_535,N_1394);
or U2675 (N_2675,N_1173,N_1746);
nand U2676 (N_2676,N_1483,N_1391);
xnor U2677 (N_2677,N_1248,N_102);
or U2678 (N_2678,N_982,N_1846);
or U2679 (N_2679,N_149,N_295);
and U2680 (N_2680,N_1201,N_66);
and U2681 (N_2681,N_401,N_249);
and U2682 (N_2682,N_1318,N_375);
and U2683 (N_2683,N_67,N_136);
or U2684 (N_2684,N_1323,N_1379);
nor U2685 (N_2685,N_597,N_1924);
nand U2686 (N_2686,N_1856,N_1028);
xor U2687 (N_2687,N_39,N_679);
or U2688 (N_2688,N_940,N_1637);
nor U2689 (N_2689,N_858,N_86);
and U2690 (N_2690,N_1428,N_1199);
xor U2691 (N_2691,N_572,N_288);
nand U2692 (N_2692,N_492,N_1444);
nor U2693 (N_2693,N_1853,N_15);
xor U2694 (N_2694,N_261,N_1551);
or U2695 (N_2695,N_1,N_1588);
or U2696 (N_2696,N_1813,N_352);
nand U2697 (N_2697,N_1528,N_872);
xnor U2698 (N_2698,N_747,N_1478);
nand U2699 (N_2699,N_69,N_860);
and U2700 (N_2700,N_758,N_156);
nand U2701 (N_2701,N_1057,N_464);
or U2702 (N_2702,N_1991,N_1745);
and U2703 (N_2703,N_193,N_61);
nand U2704 (N_2704,N_424,N_227);
xnor U2705 (N_2705,N_1128,N_847);
nand U2706 (N_2706,N_1688,N_515);
or U2707 (N_2707,N_1842,N_909);
nor U2708 (N_2708,N_1990,N_740);
xor U2709 (N_2709,N_291,N_697);
and U2710 (N_2710,N_552,N_1441);
nand U2711 (N_2711,N_639,N_876);
or U2712 (N_2712,N_970,N_1184);
nor U2713 (N_2713,N_1369,N_1606);
nand U2714 (N_2714,N_1058,N_1280);
and U2715 (N_2715,N_418,N_1542);
and U2716 (N_2716,N_728,N_109);
nand U2717 (N_2717,N_1940,N_1075);
nand U2718 (N_2718,N_413,N_438);
nor U2719 (N_2719,N_1532,N_82);
xor U2720 (N_2720,N_314,N_1596);
and U2721 (N_2721,N_1936,N_568);
and U2722 (N_2722,N_1619,N_1472);
nand U2723 (N_2723,N_1247,N_643);
and U2724 (N_2724,N_988,N_1708);
xnor U2725 (N_2725,N_1583,N_280);
or U2726 (N_2726,N_1429,N_1495);
or U2727 (N_2727,N_1332,N_1733);
or U2728 (N_2728,N_1192,N_1640);
nand U2729 (N_2729,N_821,N_967);
xnor U2730 (N_2730,N_1161,N_1556);
xor U2731 (N_2731,N_814,N_1697);
nand U2732 (N_2732,N_692,N_368);
and U2733 (N_2733,N_765,N_888);
nor U2734 (N_2734,N_1948,N_1685);
nor U2735 (N_2735,N_1031,N_751);
and U2736 (N_2736,N_870,N_611);
or U2737 (N_2737,N_1739,N_810);
nor U2738 (N_2738,N_634,N_1425);
nand U2739 (N_2739,N_950,N_1351);
xor U2740 (N_2740,N_1804,N_1073);
nor U2741 (N_2741,N_1993,N_59);
nand U2742 (N_2742,N_1171,N_904);
nand U2743 (N_2743,N_1932,N_431);
nor U2744 (N_2744,N_1001,N_180);
nand U2745 (N_2745,N_1352,N_748);
and U2746 (N_2746,N_391,N_669);
or U2747 (N_2747,N_1182,N_1085);
or U2748 (N_2748,N_90,N_340);
nand U2749 (N_2749,N_1376,N_94);
nand U2750 (N_2750,N_798,N_6);
nor U2751 (N_2751,N_176,N_1646);
and U2752 (N_2752,N_1663,N_864);
xnor U2753 (N_2753,N_1706,N_1985);
nor U2754 (N_2754,N_1347,N_1463);
xor U2755 (N_2755,N_1742,N_1125);
and U2756 (N_2756,N_633,N_1240);
and U2757 (N_2757,N_378,N_610);
or U2758 (N_2758,N_561,N_1312);
nor U2759 (N_2759,N_851,N_1808);
and U2760 (N_2760,N_1004,N_1992);
nor U2761 (N_2761,N_1440,N_544);
xor U2762 (N_2762,N_1427,N_204);
nand U2763 (N_2763,N_1465,N_8);
nand U2764 (N_2764,N_1453,N_1268);
and U2765 (N_2765,N_852,N_197);
or U2766 (N_2766,N_253,N_192);
and U2767 (N_2767,N_865,N_1169);
xnor U2768 (N_2768,N_1892,N_646);
or U2769 (N_2769,N_1390,N_128);
nand U2770 (N_2770,N_226,N_489);
and U2771 (N_2771,N_1252,N_681);
and U2772 (N_2772,N_132,N_244);
or U2773 (N_2773,N_1141,N_181);
and U2774 (N_2774,N_1083,N_310);
and U2775 (N_2775,N_406,N_859);
or U2776 (N_2776,N_1338,N_595);
or U2777 (N_2777,N_1024,N_1768);
or U2778 (N_2778,N_1873,N_1517);
nor U2779 (N_2779,N_808,N_195);
and U2780 (N_2780,N_7,N_836);
nor U2781 (N_2781,N_1118,N_1353);
nor U2782 (N_2782,N_809,N_1613);
or U2783 (N_2783,N_569,N_899);
xor U2784 (N_2784,N_285,N_1300);
and U2785 (N_2785,N_996,N_1865);
xor U2786 (N_2786,N_1738,N_1385);
xnor U2787 (N_2787,N_1213,N_1524);
or U2788 (N_2788,N_1964,N_705);
and U2789 (N_2789,N_423,N_131);
nand U2790 (N_2790,N_537,N_1530);
and U2791 (N_2791,N_1926,N_556);
xor U2792 (N_2792,N_903,N_1755);
or U2793 (N_2793,N_1292,N_594);
xor U2794 (N_2794,N_1917,N_1088);
xnor U2795 (N_2795,N_16,N_1311);
or U2796 (N_2796,N_220,N_1800);
nor U2797 (N_2797,N_1789,N_134);
or U2798 (N_2798,N_1360,N_267);
nand U2799 (N_2799,N_456,N_1744);
xnor U2800 (N_2800,N_1092,N_440);
or U2801 (N_2801,N_754,N_1949);
nand U2802 (N_2802,N_1600,N_1270);
nor U2803 (N_2803,N_1597,N_1529);
nand U2804 (N_2804,N_514,N_1785);
or U2805 (N_2805,N_1958,N_3);
xnor U2806 (N_2806,N_203,N_1918);
xnor U2807 (N_2807,N_1531,N_981);
nor U2808 (N_2808,N_80,N_114);
nor U2809 (N_2809,N_1424,N_617);
and U2810 (N_2810,N_980,N_259);
xnor U2811 (N_2811,N_97,N_1825);
xor U2812 (N_2812,N_900,N_987);
xor U2813 (N_2813,N_1194,N_309);
or U2814 (N_2814,N_1698,N_719);
and U2815 (N_2815,N_645,N_1080);
nand U2816 (N_2816,N_164,N_110);
xnor U2817 (N_2817,N_785,N_947);
or U2818 (N_2818,N_554,N_330);
and U2819 (N_2819,N_1017,N_300);
or U2820 (N_2820,N_1185,N_706);
xnor U2821 (N_2821,N_664,N_1907);
xnor U2822 (N_2822,N_233,N_855);
and U2823 (N_2823,N_158,N_1208);
or U2824 (N_2824,N_1750,N_1409);
nor U2825 (N_2825,N_1861,N_1363);
nand U2826 (N_2826,N_1174,N_1691);
or U2827 (N_2827,N_666,N_1023);
nand U2828 (N_2828,N_441,N_1937);
and U2829 (N_2829,N_567,N_420);
or U2830 (N_2830,N_144,N_414);
or U2831 (N_2831,N_1762,N_1577);
and U2832 (N_2832,N_100,N_935);
xor U2833 (N_2833,N_1067,N_1766);
xor U2834 (N_2834,N_667,N_1410);
and U2835 (N_2835,N_412,N_1172);
and U2836 (N_2836,N_726,N_245);
nand U2837 (N_2837,N_923,N_1582);
xor U2838 (N_2838,N_124,N_71);
nand U2839 (N_2839,N_1775,N_975);
nor U2840 (N_2840,N_1790,N_1205);
nand U2841 (N_2841,N_783,N_1928);
and U2842 (N_2842,N_1160,N_1573);
xor U2843 (N_2843,N_796,N_731);
or U2844 (N_2844,N_659,N_841);
nand U2845 (N_2845,N_1392,N_1652);
nand U2846 (N_2846,N_1882,N_234);
nand U2847 (N_2847,N_349,N_1076);
or U2848 (N_2848,N_60,N_1475);
or U2849 (N_2849,N_1680,N_1939);
xor U2850 (N_2850,N_1748,N_1561);
and U2851 (N_2851,N_566,N_1550);
nand U2852 (N_2852,N_350,N_1195);
xor U2853 (N_2853,N_243,N_1699);
or U2854 (N_2854,N_1980,N_1592);
xor U2855 (N_2855,N_592,N_806);
nor U2856 (N_2856,N_55,N_1548);
xor U2857 (N_2857,N_1736,N_1361);
nor U2858 (N_2858,N_570,N_479);
and U2859 (N_2859,N_718,N_781);
nor U2860 (N_2860,N_1714,N_1170);
nor U2861 (N_2861,N_752,N_1850);
nand U2862 (N_2862,N_1852,N_121);
nor U2863 (N_2863,N_24,N_427);
xnor U2864 (N_2864,N_811,N_792);
or U2865 (N_2865,N_1837,N_1593);
nor U2866 (N_2866,N_545,N_1447);
nand U2867 (N_2867,N_1758,N_426);
nand U2868 (N_2868,N_34,N_883);
nor U2869 (N_2869,N_670,N_358);
nor U2870 (N_2870,N_476,N_207);
nand U2871 (N_2871,N_1586,N_170);
nor U2872 (N_2872,N_1511,N_890);
and U2873 (N_2873,N_1605,N_1996);
and U2874 (N_2874,N_701,N_591);
nor U2875 (N_2875,N_505,N_774);
xor U2876 (N_2876,N_437,N_574);
or U2877 (N_2877,N_428,N_787);
or U2878 (N_2878,N_1298,N_827);
and U2879 (N_2879,N_1631,N_1585);
and U2880 (N_2880,N_446,N_396);
and U2881 (N_2881,N_1230,N_1732);
or U2882 (N_2882,N_421,N_383);
and U2883 (N_2883,N_830,N_1566);
xor U2884 (N_2884,N_733,N_1094);
xor U2885 (N_2885,N_1962,N_469);
and U2886 (N_2886,N_305,N_221);
or U2887 (N_2887,N_882,N_1117);
or U2888 (N_2888,N_346,N_1259);
or U2889 (N_2889,N_1454,N_1084);
or U2890 (N_2890,N_1036,N_962);
nand U2891 (N_2891,N_13,N_1811);
or U2892 (N_2892,N_1669,N_1565);
nand U2893 (N_2893,N_369,N_966);
nor U2894 (N_2894,N_1289,N_815);
or U2895 (N_2895,N_789,N_671);
nor U2896 (N_2896,N_553,N_1412);
or U2897 (N_2897,N_188,N_1370);
or U2898 (N_2898,N_1827,N_1273);
and U2899 (N_2899,N_682,N_961);
and U2900 (N_2900,N_714,N_1518);
xnor U2901 (N_2901,N_1271,N_189);
or U2902 (N_2902,N_360,N_1814);
or U2903 (N_2903,N_1509,N_297);
nor U2904 (N_2904,N_1540,N_1564);
xnor U2905 (N_2905,N_1335,N_1726);
or U2906 (N_2906,N_1722,N_123);
or U2907 (N_2907,N_910,N_1868);
or U2908 (N_2908,N_1671,N_1119);
nand U2909 (N_2909,N_173,N_993);
nor U2910 (N_2910,N_1897,N_1377);
xnor U2911 (N_2911,N_1457,N_1480);
nor U2912 (N_2912,N_148,N_1139);
and U2913 (N_2913,N_1603,N_1309);
nor U2914 (N_2914,N_878,N_1123);
xnor U2915 (N_2915,N_1925,N_1466);
and U2916 (N_2916,N_522,N_1754);
nand U2917 (N_2917,N_1070,N_1037);
nor U2918 (N_2918,N_776,N_1371);
and U2919 (N_2919,N_724,N_930);
nor U2920 (N_2920,N_1217,N_524);
xor U2921 (N_2921,N_927,N_1612);
or U2922 (N_2922,N_1618,N_1623);
and U2923 (N_2923,N_1293,N_519);
xor U2924 (N_2924,N_326,N_1115);
and U2925 (N_2925,N_178,N_1796);
nand U2926 (N_2926,N_974,N_951);
and U2927 (N_2927,N_1430,N_1632);
or U2928 (N_2928,N_325,N_274);
xnor U2929 (N_2929,N_1200,N_206);
and U2930 (N_2930,N_1696,N_1607);
and U2931 (N_2931,N_1514,N_284);
nor U2932 (N_2932,N_415,N_1404);
and U2933 (N_2933,N_362,N_1570);
or U2934 (N_2934,N_973,N_1434);
and U2935 (N_2935,N_335,N_111);
nand U2936 (N_2936,N_1525,N_536);
xor U2937 (N_2937,N_912,N_969);
or U2938 (N_2938,N_1439,N_896);
nor U2939 (N_2939,N_1703,N_367);
and U2940 (N_2940,N_791,N_700);
nand U2941 (N_2941,N_762,N_691);
or U2942 (N_2942,N_1716,N_1840);
or U2943 (N_2943,N_1765,N_43);
nor U2944 (N_2944,N_1100,N_161);
and U2945 (N_2945,N_1110,N_1072);
or U2946 (N_2946,N_211,N_1595);
nand U2947 (N_2947,N_177,N_908);
nor U2948 (N_2948,N_1959,N_129);
or U2949 (N_2949,N_1686,N_138);
and U2950 (N_2950,N_1095,N_202);
nand U2951 (N_2951,N_1047,N_955);
and U2952 (N_2952,N_773,N_647);
and U2953 (N_2953,N_511,N_1908);
nand U2954 (N_2954,N_1013,N_403);
nor U2955 (N_2955,N_395,N_45);
nor U2956 (N_2956,N_182,N_451);
nor U2957 (N_2957,N_873,N_942);
xnor U2958 (N_2958,N_716,N_510);
nand U2959 (N_2959,N_946,N_782);
nand U2960 (N_2960,N_268,N_405);
xnor U2961 (N_2961,N_1455,N_425);
xor U2962 (N_2962,N_1469,N_1794);
and U2963 (N_2963,N_171,N_1759);
nand U2964 (N_2964,N_399,N_1504);
or U2965 (N_2965,N_1520,N_1594);
or U2966 (N_2966,N_1553,N_179);
or U2967 (N_2967,N_964,N_42);
xor U2968 (N_2968,N_1034,N_557);
or U2969 (N_2969,N_379,N_468);
nor U2970 (N_2970,N_755,N_1179);
nor U2971 (N_2971,N_1587,N_223);
and U2972 (N_2972,N_839,N_1898);
nor U2973 (N_2973,N_169,N_2);
and U2974 (N_2974,N_1389,N_235);
or U2975 (N_2975,N_674,N_1097);
or U2976 (N_2976,N_913,N_1302);
and U2977 (N_2977,N_1578,N_254);
nand U2978 (N_2978,N_1132,N_1124);
nor U2979 (N_2979,N_1662,N_943);
xor U2980 (N_2980,N_1911,N_87);
nand U2981 (N_2981,N_625,N_1209);
nor U2982 (N_2982,N_532,N_1071);
and U2983 (N_2983,N_1960,N_496);
or U2984 (N_2984,N_1836,N_637);
and U2985 (N_2985,N_662,N_1378);
and U2986 (N_2986,N_1158,N_1667);
or U2987 (N_2987,N_824,N_826);
or U2988 (N_2988,N_1086,N_644);
nand U2989 (N_2989,N_619,N_1590);
nand U2990 (N_2990,N_1368,N_1120);
nor U2991 (N_2991,N_448,N_1380);
or U2992 (N_2992,N_1860,N_1823);
and U2993 (N_2993,N_484,N_840);
or U2994 (N_2994,N_1676,N_1974);
nand U2995 (N_2995,N_704,N_1178);
xor U2996 (N_2996,N_1649,N_1276);
nor U2997 (N_2997,N_1272,N_1541);
nor U2998 (N_2998,N_1763,N_485);
and U2999 (N_2999,N_1433,N_1337);
or U3000 (N_3000,N_779,N_105);
nor U3001 (N_3001,N_1914,N_803);
nor U3002 (N_3002,N_1543,N_1583);
xnor U3003 (N_3003,N_1009,N_266);
or U3004 (N_3004,N_1258,N_715);
xor U3005 (N_3005,N_1002,N_1850);
nand U3006 (N_3006,N_111,N_1324);
or U3007 (N_3007,N_1189,N_37);
or U3008 (N_3008,N_462,N_1597);
and U3009 (N_3009,N_590,N_1866);
xor U3010 (N_3010,N_1930,N_1938);
or U3011 (N_3011,N_1412,N_147);
and U3012 (N_3012,N_137,N_1213);
nand U3013 (N_3013,N_429,N_1538);
or U3014 (N_3014,N_363,N_690);
and U3015 (N_3015,N_1157,N_1067);
xor U3016 (N_3016,N_1604,N_339);
nand U3017 (N_3017,N_980,N_602);
nand U3018 (N_3018,N_835,N_201);
nand U3019 (N_3019,N_148,N_743);
nor U3020 (N_3020,N_1536,N_158);
nor U3021 (N_3021,N_313,N_1688);
xor U3022 (N_3022,N_127,N_1502);
xnor U3023 (N_3023,N_1873,N_482);
or U3024 (N_3024,N_1081,N_1655);
or U3025 (N_3025,N_1590,N_1253);
xor U3026 (N_3026,N_1816,N_1629);
or U3027 (N_3027,N_180,N_351);
or U3028 (N_3028,N_1405,N_1120);
or U3029 (N_3029,N_1699,N_327);
nand U3030 (N_3030,N_1186,N_1937);
xor U3031 (N_3031,N_1113,N_1399);
or U3032 (N_3032,N_923,N_1673);
nor U3033 (N_3033,N_66,N_1549);
nand U3034 (N_3034,N_701,N_699);
xor U3035 (N_3035,N_1477,N_1981);
nor U3036 (N_3036,N_1741,N_1968);
or U3037 (N_3037,N_1075,N_1600);
and U3038 (N_3038,N_470,N_226);
and U3039 (N_3039,N_229,N_1348);
and U3040 (N_3040,N_412,N_1178);
nand U3041 (N_3041,N_1981,N_465);
xor U3042 (N_3042,N_262,N_863);
nand U3043 (N_3043,N_810,N_19);
nor U3044 (N_3044,N_768,N_457);
and U3045 (N_3045,N_1757,N_1932);
and U3046 (N_3046,N_968,N_1785);
nand U3047 (N_3047,N_202,N_1064);
xor U3048 (N_3048,N_1277,N_436);
nand U3049 (N_3049,N_804,N_577);
nor U3050 (N_3050,N_1587,N_486);
xnor U3051 (N_3051,N_323,N_1917);
xnor U3052 (N_3052,N_1497,N_1600);
nand U3053 (N_3053,N_975,N_1502);
nand U3054 (N_3054,N_252,N_1620);
nand U3055 (N_3055,N_1923,N_796);
or U3056 (N_3056,N_1021,N_786);
nor U3057 (N_3057,N_1723,N_332);
or U3058 (N_3058,N_1480,N_553);
nand U3059 (N_3059,N_1959,N_1726);
or U3060 (N_3060,N_1377,N_1039);
and U3061 (N_3061,N_428,N_1861);
xor U3062 (N_3062,N_306,N_965);
nand U3063 (N_3063,N_425,N_28);
nor U3064 (N_3064,N_732,N_934);
or U3065 (N_3065,N_159,N_1251);
xor U3066 (N_3066,N_778,N_1426);
xor U3067 (N_3067,N_993,N_371);
and U3068 (N_3068,N_1384,N_1170);
xnor U3069 (N_3069,N_486,N_553);
xor U3070 (N_3070,N_1020,N_168);
xnor U3071 (N_3071,N_373,N_1432);
or U3072 (N_3072,N_1959,N_805);
nand U3073 (N_3073,N_22,N_1342);
nand U3074 (N_3074,N_1137,N_726);
or U3075 (N_3075,N_903,N_818);
xor U3076 (N_3076,N_90,N_1117);
nand U3077 (N_3077,N_1186,N_171);
nor U3078 (N_3078,N_1725,N_48);
nor U3079 (N_3079,N_1052,N_1630);
nor U3080 (N_3080,N_44,N_639);
nand U3081 (N_3081,N_207,N_1253);
nor U3082 (N_3082,N_1726,N_946);
nor U3083 (N_3083,N_1454,N_1862);
nand U3084 (N_3084,N_295,N_1111);
nand U3085 (N_3085,N_1096,N_311);
nand U3086 (N_3086,N_647,N_1347);
nor U3087 (N_3087,N_1734,N_384);
and U3088 (N_3088,N_371,N_1725);
nor U3089 (N_3089,N_1558,N_1707);
nor U3090 (N_3090,N_148,N_1720);
xor U3091 (N_3091,N_924,N_1211);
and U3092 (N_3092,N_507,N_1652);
and U3093 (N_3093,N_404,N_1324);
xor U3094 (N_3094,N_723,N_664);
and U3095 (N_3095,N_1017,N_387);
nor U3096 (N_3096,N_367,N_1875);
and U3097 (N_3097,N_321,N_1562);
and U3098 (N_3098,N_1689,N_109);
xnor U3099 (N_3099,N_608,N_337);
or U3100 (N_3100,N_1067,N_1202);
nor U3101 (N_3101,N_419,N_1102);
nor U3102 (N_3102,N_1947,N_1105);
and U3103 (N_3103,N_397,N_1830);
or U3104 (N_3104,N_1049,N_468);
xnor U3105 (N_3105,N_1487,N_579);
nor U3106 (N_3106,N_1269,N_1465);
or U3107 (N_3107,N_846,N_1820);
xnor U3108 (N_3108,N_955,N_1069);
and U3109 (N_3109,N_1042,N_857);
nand U3110 (N_3110,N_383,N_1940);
xor U3111 (N_3111,N_129,N_1883);
and U3112 (N_3112,N_500,N_375);
nand U3113 (N_3113,N_1211,N_870);
and U3114 (N_3114,N_1479,N_678);
xnor U3115 (N_3115,N_1798,N_1779);
or U3116 (N_3116,N_1471,N_181);
or U3117 (N_3117,N_87,N_156);
nor U3118 (N_3118,N_1720,N_1834);
or U3119 (N_3119,N_1203,N_167);
nor U3120 (N_3120,N_1425,N_4);
and U3121 (N_3121,N_764,N_1043);
and U3122 (N_3122,N_761,N_1491);
or U3123 (N_3123,N_1386,N_731);
nand U3124 (N_3124,N_1598,N_1818);
nand U3125 (N_3125,N_527,N_193);
and U3126 (N_3126,N_1500,N_1016);
nand U3127 (N_3127,N_1505,N_1679);
nor U3128 (N_3128,N_1327,N_1372);
nor U3129 (N_3129,N_666,N_1918);
xor U3130 (N_3130,N_320,N_1156);
and U3131 (N_3131,N_1300,N_263);
xnor U3132 (N_3132,N_269,N_194);
and U3133 (N_3133,N_1473,N_1476);
and U3134 (N_3134,N_965,N_1161);
nand U3135 (N_3135,N_857,N_1861);
nand U3136 (N_3136,N_1097,N_6);
and U3137 (N_3137,N_1254,N_482);
nand U3138 (N_3138,N_151,N_303);
nor U3139 (N_3139,N_255,N_428);
xor U3140 (N_3140,N_1654,N_676);
nand U3141 (N_3141,N_687,N_1255);
xnor U3142 (N_3142,N_1296,N_323);
and U3143 (N_3143,N_1401,N_922);
nand U3144 (N_3144,N_57,N_823);
xor U3145 (N_3145,N_1804,N_1498);
nor U3146 (N_3146,N_588,N_8);
and U3147 (N_3147,N_717,N_188);
or U3148 (N_3148,N_444,N_1717);
nand U3149 (N_3149,N_503,N_1263);
or U3150 (N_3150,N_852,N_752);
xor U3151 (N_3151,N_1435,N_496);
and U3152 (N_3152,N_1017,N_1498);
nor U3153 (N_3153,N_1524,N_747);
nor U3154 (N_3154,N_808,N_1344);
nand U3155 (N_3155,N_1919,N_875);
or U3156 (N_3156,N_68,N_298);
and U3157 (N_3157,N_1337,N_467);
nand U3158 (N_3158,N_1045,N_1925);
nor U3159 (N_3159,N_291,N_1820);
xnor U3160 (N_3160,N_1771,N_989);
or U3161 (N_3161,N_1964,N_97);
nand U3162 (N_3162,N_944,N_1697);
nor U3163 (N_3163,N_162,N_1761);
nand U3164 (N_3164,N_542,N_755);
or U3165 (N_3165,N_1557,N_1932);
and U3166 (N_3166,N_1171,N_499);
and U3167 (N_3167,N_300,N_312);
and U3168 (N_3168,N_59,N_768);
nor U3169 (N_3169,N_732,N_1527);
nor U3170 (N_3170,N_1600,N_652);
nor U3171 (N_3171,N_1056,N_1249);
xor U3172 (N_3172,N_1297,N_1477);
xnor U3173 (N_3173,N_924,N_81);
or U3174 (N_3174,N_1875,N_1681);
and U3175 (N_3175,N_896,N_1918);
and U3176 (N_3176,N_1535,N_1493);
xor U3177 (N_3177,N_1205,N_1063);
and U3178 (N_3178,N_104,N_1117);
nand U3179 (N_3179,N_1841,N_767);
or U3180 (N_3180,N_510,N_1879);
and U3181 (N_3181,N_377,N_1368);
or U3182 (N_3182,N_1514,N_1378);
or U3183 (N_3183,N_1814,N_272);
nand U3184 (N_3184,N_1615,N_1037);
or U3185 (N_3185,N_1093,N_262);
and U3186 (N_3186,N_1992,N_598);
xor U3187 (N_3187,N_1654,N_1607);
xnor U3188 (N_3188,N_42,N_147);
xor U3189 (N_3189,N_1736,N_1772);
xor U3190 (N_3190,N_474,N_133);
nor U3191 (N_3191,N_1131,N_335);
or U3192 (N_3192,N_323,N_574);
and U3193 (N_3193,N_494,N_196);
xor U3194 (N_3194,N_930,N_134);
nor U3195 (N_3195,N_1879,N_267);
xnor U3196 (N_3196,N_1527,N_809);
or U3197 (N_3197,N_1609,N_1837);
xor U3198 (N_3198,N_1752,N_1436);
or U3199 (N_3199,N_1679,N_169);
or U3200 (N_3200,N_1910,N_1447);
xnor U3201 (N_3201,N_378,N_1488);
nand U3202 (N_3202,N_1749,N_317);
nand U3203 (N_3203,N_506,N_1219);
nand U3204 (N_3204,N_1450,N_311);
xor U3205 (N_3205,N_468,N_1846);
nor U3206 (N_3206,N_37,N_1048);
nor U3207 (N_3207,N_541,N_134);
nor U3208 (N_3208,N_409,N_1795);
xor U3209 (N_3209,N_1,N_788);
xnor U3210 (N_3210,N_543,N_255);
and U3211 (N_3211,N_10,N_125);
nor U3212 (N_3212,N_1208,N_1270);
and U3213 (N_3213,N_398,N_807);
nand U3214 (N_3214,N_169,N_1868);
nor U3215 (N_3215,N_840,N_1090);
nand U3216 (N_3216,N_792,N_1516);
xnor U3217 (N_3217,N_21,N_1418);
nand U3218 (N_3218,N_1347,N_1528);
or U3219 (N_3219,N_1827,N_1132);
nor U3220 (N_3220,N_1919,N_959);
nand U3221 (N_3221,N_1700,N_1698);
xor U3222 (N_3222,N_874,N_716);
nor U3223 (N_3223,N_1788,N_466);
nor U3224 (N_3224,N_316,N_1917);
nand U3225 (N_3225,N_1071,N_694);
nand U3226 (N_3226,N_1171,N_1227);
or U3227 (N_3227,N_961,N_718);
or U3228 (N_3228,N_901,N_515);
or U3229 (N_3229,N_1598,N_370);
and U3230 (N_3230,N_1601,N_569);
nand U3231 (N_3231,N_1449,N_123);
or U3232 (N_3232,N_680,N_720);
nand U3233 (N_3233,N_84,N_1825);
or U3234 (N_3234,N_1547,N_974);
nand U3235 (N_3235,N_251,N_1160);
or U3236 (N_3236,N_645,N_216);
and U3237 (N_3237,N_1933,N_985);
or U3238 (N_3238,N_632,N_349);
xor U3239 (N_3239,N_1415,N_691);
nor U3240 (N_3240,N_1530,N_879);
nand U3241 (N_3241,N_453,N_478);
nand U3242 (N_3242,N_1509,N_971);
or U3243 (N_3243,N_932,N_1837);
or U3244 (N_3244,N_885,N_737);
or U3245 (N_3245,N_1236,N_1598);
and U3246 (N_3246,N_1507,N_1045);
nor U3247 (N_3247,N_869,N_528);
nor U3248 (N_3248,N_737,N_1089);
nand U3249 (N_3249,N_1838,N_1539);
and U3250 (N_3250,N_1954,N_412);
or U3251 (N_3251,N_987,N_1788);
or U3252 (N_3252,N_623,N_348);
and U3253 (N_3253,N_1662,N_1028);
xnor U3254 (N_3254,N_1558,N_1696);
or U3255 (N_3255,N_1322,N_1228);
xnor U3256 (N_3256,N_1937,N_1520);
nor U3257 (N_3257,N_1672,N_16);
or U3258 (N_3258,N_1350,N_358);
and U3259 (N_3259,N_830,N_86);
or U3260 (N_3260,N_1645,N_1799);
nand U3261 (N_3261,N_1742,N_1013);
or U3262 (N_3262,N_212,N_1125);
or U3263 (N_3263,N_255,N_1934);
or U3264 (N_3264,N_1000,N_979);
nor U3265 (N_3265,N_1467,N_602);
and U3266 (N_3266,N_557,N_848);
or U3267 (N_3267,N_797,N_1454);
xnor U3268 (N_3268,N_107,N_232);
nand U3269 (N_3269,N_1129,N_519);
xnor U3270 (N_3270,N_901,N_997);
and U3271 (N_3271,N_216,N_1062);
xnor U3272 (N_3272,N_1297,N_1851);
xnor U3273 (N_3273,N_1190,N_526);
nor U3274 (N_3274,N_566,N_877);
nor U3275 (N_3275,N_941,N_108);
nor U3276 (N_3276,N_1058,N_1927);
and U3277 (N_3277,N_1775,N_1490);
nand U3278 (N_3278,N_1407,N_751);
and U3279 (N_3279,N_1974,N_1863);
and U3280 (N_3280,N_1282,N_1314);
nor U3281 (N_3281,N_1816,N_1761);
nand U3282 (N_3282,N_413,N_1200);
and U3283 (N_3283,N_1439,N_1724);
and U3284 (N_3284,N_227,N_545);
nor U3285 (N_3285,N_230,N_657);
xor U3286 (N_3286,N_943,N_1973);
nand U3287 (N_3287,N_190,N_43);
and U3288 (N_3288,N_1449,N_360);
xnor U3289 (N_3289,N_1445,N_1574);
and U3290 (N_3290,N_624,N_1090);
and U3291 (N_3291,N_901,N_1802);
nor U3292 (N_3292,N_188,N_318);
or U3293 (N_3293,N_1506,N_67);
and U3294 (N_3294,N_988,N_381);
and U3295 (N_3295,N_1174,N_521);
or U3296 (N_3296,N_106,N_1185);
and U3297 (N_3297,N_1966,N_586);
nand U3298 (N_3298,N_1772,N_1174);
and U3299 (N_3299,N_318,N_1400);
nand U3300 (N_3300,N_14,N_441);
or U3301 (N_3301,N_66,N_1379);
nand U3302 (N_3302,N_1640,N_169);
or U3303 (N_3303,N_426,N_1088);
and U3304 (N_3304,N_1314,N_1180);
nand U3305 (N_3305,N_645,N_134);
xnor U3306 (N_3306,N_1489,N_647);
or U3307 (N_3307,N_774,N_29);
and U3308 (N_3308,N_1773,N_1298);
xnor U3309 (N_3309,N_1556,N_1011);
xor U3310 (N_3310,N_656,N_618);
xor U3311 (N_3311,N_1606,N_1292);
nand U3312 (N_3312,N_1211,N_1154);
and U3313 (N_3313,N_576,N_727);
nor U3314 (N_3314,N_1411,N_328);
and U3315 (N_3315,N_1033,N_1608);
or U3316 (N_3316,N_1618,N_543);
nand U3317 (N_3317,N_1399,N_1189);
nand U3318 (N_3318,N_1672,N_1468);
or U3319 (N_3319,N_639,N_1555);
and U3320 (N_3320,N_1695,N_1678);
nand U3321 (N_3321,N_1207,N_173);
nand U3322 (N_3322,N_151,N_1596);
nand U3323 (N_3323,N_1622,N_1330);
or U3324 (N_3324,N_896,N_263);
nand U3325 (N_3325,N_505,N_425);
or U3326 (N_3326,N_1701,N_1249);
or U3327 (N_3327,N_1493,N_1532);
nor U3328 (N_3328,N_297,N_852);
nor U3329 (N_3329,N_463,N_868);
xor U3330 (N_3330,N_530,N_2);
xor U3331 (N_3331,N_548,N_1715);
or U3332 (N_3332,N_904,N_99);
and U3333 (N_3333,N_1868,N_1837);
nor U3334 (N_3334,N_1208,N_121);
xor U3335 (N_3335,N_1405,N_1201);
or U3336 (N_3336,N_917,N_149);
xor U3337 (N_3337,N_1236,N_624);
xor U3338 (N_3338,N_1281,N_1980);
and U3339 (N_3339,N_135,N_1897);
and U3340 (N_3340,N_501,N_1081);
xnor U3341 (N_3341,N_1044,N_901);
nand U3342 (N_3342,N_1310,N_845);
and U3343 (N_3343,N_827,N_1142);
or U3344 (N_3344,N_1278,N_1303);
or U3345 (N_3345,N_119,N_25);
nand U3346 (N_3346,N_415,N_1526);
xor U3347 (N_3347,N_1361,N_928);
nand U3348 (N_3348,N_1774,N_1422);
and U3349 (N_3349,N_1499,N_1178);
or U3350 (N_3350,N_1106,N_446);
or U3351 (N_3351,N_893,N_1915);
or U3352 (N_3352,N_1775,N_1192);
xor U3353 (N_3353,N_129,N_1414);
xnor U3354 (N_3354,N_1839,N_531);
nand U3355 (N_3355,N_649,N_1364);
nand U3356 (N_3356,N_1246,N_486);
or U3357 (N_3357,N_160,N_1955);
and U3358 (N_3358,N_1113,N_1909);
and U3359 (N_3359,N_1209,N_390);
and U3360 (N_3360,N_1603,N_216);
nor U3361 (N_3361,N_1550,N_435);
xnor U3362 (N_3362,N_1362,N_1330);
and U3363 (N_3363,N_1113,N_1713);
xor U3364 (N_3364,N_437,N_578);
and U3365 (N_3365,N_179,N_774);
nand U3366 (N_3366,N_1939,N_600);
nand U3367 (N_3367,N_125,N_717);
xnor U3368 (N_3368,N_85,N_170);
nand U3369 (N_3369,N_1861,N_1059);
or U3370 (N_3370,N_483,N_1787);
and U3371 (N_3371,N_112,N_145);
nand U3372 (N_3372,N_1347,N_490);
or U3373 (N_3373,N_1490,N_18);
and U3374 (N_3374,N_1878,N_480);
nor U3375 (N_3375,N_1885,N_591);
nand U3376 (N_3376,N_1555,N_169);
and U3377 (N_3377,N_673,N_179);
nand U3378 (N_3378,N_1594,N_1199);
xnor U3379 (N_3379,N_1819,N_696);
nand U3380 (N_3380,N_1112,N_1704);
nand U3381 (N_3381,N_1705,N_1280);
or U3382 (N_3382,N_50,N_476);
xor U3383 (N_3383,N_1386,N_33);
nor U3384 (N_3384,N_717,N_1504);
xnor U3385 (N_3385,N_151,N_1220);
and U3386 (N_3386,N_1145,N_1990);
nand U3387 (N_3387,N_761,N_815);
and U3388 (N_3388,N_1988,N_666);
nor U3389 (N_3389,N_1931,N_1279);
and U3390 (N_3390,N_111,N_1510);
xor U3391 (N_3391,N_833,N_257);
nand U3392 (N_3392,N_1842,N_1329);
and U3393 (N_3393,N_1483,N_1963);
nor U3394 (N_3394,N_1673,N_1494);
nor U3395 (N_3395,N_372,N_1581);
xnor U3396 (N_3396,N_219,N_290);
nor U3397 (N_3397,N_1247,N_1414);
xor U3398 (N_3398,N_1330,N_1466);
xor U3399 (N_3399,N_299,N_867);
nand U3400 (N_3400,N_1822,N_60);
and U3401 (N_3401,N_1149,N_1316);
and U3402 (N_3402,N_1282,N_1729);
xor U3403 (N_3403,N_1730,N_1519);
and U3404 (N_3404,N_1790,N_20);
or U3405 (N_3405,N_1676,N_747);
xnor U3406 (N_3406,N_1303,N_281);
xor U3407 (N_3407,N_910,N_874);
and U3408 (N_3408,N_789,N_511);
xnor U3409 (N_3409,N_65,N_1366);
nand U3410 (N_3410,N_233,N_1022);
or U3411 (N_3411,N_78,N_334);
nand U3412 (N_3412,N_496,N_1486);
or U3413 (N_3413,N_853,N_435);
xor U3414 (N_3414,N_1832,N_1058);
nor U3415 (N_3415,N_770,N_111);
nor U3416 (N_3416,N_1882,N_1275);
nand U3417 (N_3417,N_275,N_1484);
xor U3418 (N_3418,N_489,N_1258);
and U3419 (N_3419,N_1826,N_272);
or U3420 (N_3420,N_1760,N_1133);
or U3421 (N_3421,N_1505,N_488);
and U3422 (N_3422,N_940,N_722);
and U3423 (N_3423,N_1452,N_1555);
xnor U3424 (N_3424,N_1493,N_1587);
nand U3425 (N_3425,N_1592,N_128);
and U3426 (N_3426,N_426,N_1133);
and U3427 (N_3427,N_773,N_1426);
xor U3428 (N_3428,N_1190,N_1267);
nor U3429 (N_3429,N_504,N_1035);
nand U3430 (N_3430,N_223,N_1525);
nand U3431 (N_3431,N_871,N_735);
nor U3432 (N_3432,N_1134,N_1744);
xnor U3433 (N_3433,N_770,N_1808);
xor U3434 (N_3434,N_1675,N_171);
and U3435 (N_3435,N_1104,N_770);
xor U3436 (N_3436,N_47,N_1840);
and U3437 (N_3437,N_189,N_1659);
and U3438 (N_3438,N_849,N_1957);
or U3439 (N_3439,N_442,N_576);
or U3440 (N_3440,N_1960,N_211);
xnor U3441 (N_3441,N_1138,N_521);
nand U3442 (N_3442,N_1023,N_94);
or U3443 (N_3443,N_664,N_1013);
nor U3444 (N_3444,N_1645,N_962);
or U3445 (N_3445,N_804,N_1259);
and U3446 (N_3446,N_705,N_437);
nand U3447 (N_3447,N_600,N_193);
xor U3448 (N_3448,N_1810,N_1130);
and U3449 (N_3449,N_450,N_889);
and U3450 (N_3450,N_1671,N_1990);
nand U3451 (N_3451,N_1601,N_54);
nor U3452 (N_3452,N_440,N_207);
nand U3453 (N_3453,N_1230,N_1176);
and U3454 (N_3454,N_1797,N_358);
nor U3455 (N_3455,N_485,N_1446);
nor U3456 (N_3456,N_266,N_1692);
xnor U3457 (N_3457,N_741,N_626);
xnor U3458 (N_3458,N_1317,N_1779);
or U3459 (N_3459,N_773,N_1197);
xnor U3460 (N_3460,N_256,N_269);
nor U3461 (N_3461,N_610,N_1732);
xnor U3462 (N_3462,N_97,N_1978);
nor U3463 (N_3463,N_822,N_886);
xor U3464 (N_3464,N_1478,N_505);
or U3465 (N_3465,N_306,N_1822);
xnor U3466 (N_3466,N_632,N_1605);
xnor U3467 (N_3467,N_202,N_1561);
and U3468 (N_3468,N_1714,N_1926);
and U3469 (N_3469,N_356,N_474);
nor U3470 (N_3470,N_1875,N_1065);
or U3471 (N_3471,N_802,N_41);
nand U3472 (N_3472,N_1396,N_1811);
nor U3473 (N_3473,N_247,N_723);
nand U3474 (N_3474,N_1706,N_1198);
or U3475 (N_3475,N_985,N_1675);
and U3476 (N_3476,N_800,N_1635);
xnor U3477 (N_3477,N_1125,N_1229);
or U3478 (N_3478,N_475,N_301);
or U3479 (N_3479,N_1413,N_935);
nand U3480 (N_3480,N_792,N_802);
xor U3481 (N_3481,N_445,N_1837);
or U3482 (N_3482,N_252,N_1365);
xnor U3483 (N_3483,N_278,N_533);
nand U3484 (N_3484,N_1385,N_1102);
xnor U3485 (N_3485,N_604,N_1738);
xnor U3486 (N_3486,N_899,N_1845);
or U3487 (N_3487,N_924,N_150);
nor U3488 (N_3488,N_953,N_1282);
nand U3489 (N_3489,N_184,N_1175);
xnor U3490 (N_3490,N_1596,N_1898);
or U3491 (N_3491,N_1606,N_1498);
or U3492 (N_3492,N_1845,N_1353);
and U3493 (N_3493,N_349,N_440);
xnor U3494 (N_3494,N_1107,N_911);
or U3495 (N_3495,N_1472,N_392);
xor U3496 (N_3496,N_1928,N_1845);
nor U3497 (N_3497,N_833,N_1977);
and U3498 (N_3498,N_1529,N_673);
nand U3499 (N_3499,N_812,N_1309);
nor U3500 (N_3500,N_387,N_261);
xnor U3501 (N_3501,N_1269,N_159);
and U3502 (N_3502,N_244,N_1754);
nor U3503 (N_3503,N_921,N_1644);
or U3504 (N_3504,N_539,N_771);
nand U3505 (N_3505,N_791,N_918);
xnor U3506 (N_3506,N_815,N_204);
xor U3507 (N_3507,N_537,N_266);
nand U3508 (N_3508,N_909,N_1925);
and U3509 (N_3509,N_316,N_1417);
or U3510 (N_3510,N_1660,N_615);
and U3511 (N_3511,N_1023,N_1617);
or U3512 (N_3512,N_1053,N_27);
and U3513 (N_3513,N_670,N_532);
or U3514 (N_3514,N_313,N_1202);
nand U3515 (N_3515,N_994,N_848);
nor U3516 (N_3516,N_197,N_401);
or U3517 (N_3517,N_1449,N_1161);
or U3518 (N_3518,N_1529,N_1370);
nand U3519 (N_3519,N_1418,N_778);
nand U3520 (N_3520,N_139,N_1103);
nor U3521 (N_3521,N_434,N_1652);
or U3522 (N_3522,N_983,N_432);
and U3523 (N_3523,N_956,N_785);
nor U3524 (N_3524,N_825,N_1167);
nor U3525 (N_3525,N_885,N_1509);
or U3526 (N_3526,N_1152,N_1713);
nand U3527 (N_3527,N_1013,N_529);
or U3528 (N_3528,N_1137,N_483);
xor U3529 (N_3529,N_564,N_142);
xor U3530 (N_3530,N_970,N_290);
xor U3531 (N_3531,N_489,N_1822);
nand U3532 (N_3532,N_926,N_825);
xnor U3533 (N_3533,N_17,N_985);
nand U3534 (N_3534,N_180,N_1094);
and U3535 (N_3535,N_40,N_460);
xnor U3536 (N_3536,N_1529,N_1519);
nor U3537 (N_3537,N_1112,N_1612);
nand U3538 (N_3538,N_1169,N_1252);
or U3539 (N_3539,N_1667,N_1125);
or U3540 (N_3540,N_1698,N_412);
xnor U3541 (N_3541,N_1413,N_788);
nand U3542 (N_3542,N_373,N_1619);
nand U3543 (N_3543,N_1609,N_1938);
nand U3544 (N_3544,N_1221,N_426);
xor U3545 (N_3545,N_359,N_32);
nor U3546 (N_3546,N_1272,N_973);
nand U3547 (N_3547,N_1787,N_1968);
and U3548 (N_3548,N_1429,N_137);
and U3549 (N_3549,N_435,N_353);
nand U3550 (N_3550,N_490,N_1370);
nor U3551 (N_3551,N_840,N_1237);
nand U3552 (N_3552,N_621,N_1697);
and U3553 (N_3553,N_1085,N_1809);
or U3554 (N_3554,N_715,N_1118);
nand U3555 (N_3555,N_1255,N_447);
xnor U3556 (N_3556,N_1108,N_699);
xnor U3557 (N_3557,N_779,N_120);
nand U3558 (N_3558,N_1558,N_1384);
or U3559 (N_3559,N_526,N_603);
nor U3560 (N_3560,N_1674,N_520);
and U3561 (N_3561,N_565,N_818);
or U3562 (N_3562,N_1280,N_1625);
xnor U3563 (N_3563,N_490,N_833);
or U3564 (N_3564,N_842,N_511);
or U3565 (N_3565,N_1674,N_71);
nand U3566 (N_3566,N_441,N_290);
or U3567 (N_3567,N_1330,N_1030);
nand U3568 (N_3568,N_857,N_57);
or U3569 (N_3569,N_1084,N_54);
xnor U3570 (N_3570,N_1529,N_775);
or U3571 (N_3571,N_1454,N_217);
nor U3572 (N_3572,N_225,N_1299);
and U3573 (N_3573,N_1993,N_579);
or U3574 (N_3574,N_972,N_1329);
xnor U3575 (N_3575,N_215,N_1919);
nor U3576 (N_3576,N_563,N_429);
and U3577 (N_3577,N_163,N_1915);
or U3578 (N_3578,N_710,N_1814);
nor U3579 (N_3579,N_1898,N_1);
or U3580 (N_3580,N_1307,N_498);
and U3581 (N_3581,N_1845,N_263);
xnor U3582 (N_3582,N_663,N_1912);
and U3583 (N_3583,N_778,N_1409);
nor U3584 (N_3584,N_1941,N_170);
nor U3585 (N_3585,N_1698,N_1916);
and U3586 (N_3586,N_1974,N_644);
or U3587 (N_3587,N_985,N_1171);
nand U3588 (N_3588,N_841,N_1907);
xor U3589 (N_3589,N_1028,N_1723);
nor U3590 (N_3590,N_1945,N_1827);
xnor U3591 (N_3591,N_1027,N_1368);
nand U3592 (N_3592,N_1473,N_1861);
xnor U3593 (N_3593,N_1831,N_1312);
and U3594 (N_3594,N_1564,N_1546);
nor U3595 (N_3595,N_1120,N_36);
or U3596 (N_3596,N_901,N_204);
nor U3597 (N_3597,N_167,N_716);
or U3598 (N_3598,N_67,N_433);
and U3599 (N_3599,N_724,N_811);
xnor U3600 (N_3600,N_1758,N_967);
nor U3601 (N_3601,N_431,N_1741);
nor U3602 (N_3602,N_476,N_211);
nand U3603 (N_3603,N_716,N_957);
or U3604 (N_3604,N_1741,N_1375);
xor U3605 (N_3605,N_728,N_672);
xor U3606 (N_3606,N_1197,N_24);
or U3607 (N_3607,N_1377,N_717);
xor U3608 (N_3608,N_1576,N_52);
xor U3609 (N_3609,N_1161,N_311);
nor U3610 (N_3610,N_1957,N_42);
nand U3611 (N_3611,N_1876,N_1024);
and U3612 (N_3612,N_1285,N_1697);
or U3613 (N_3613,N_1266,N_522);
xnor U3614 (N_3614,N_1243,N_441);
or U3615 (N_3615,N_1587,N_1256);
nand U3616 (N_3616,N_459,N_1575);
nand U3617 (N_3617,N_762,N_809);
and U3618 (N_3618,N_1673,N_17);
or U3619 (N_3619,N_1711,N_1702);
nand U3620 (N_3620,N_1516,N_477);
or U3621 (N_3621,N_1551,N_1434);
or U3622 (N_3622,N_912,N_1732);
or U3623 (N_3623,N_556,N_394);
nand U3624 (N_3624,N_1343,N_5);
nor U3625 (N_3625,N_568,N_1114);
or U3626 (N_3626,N_1283,N_1844);
nor U3627 (N_3627,N_685,N_988);
nand U3628 (N_3628,N_1886,N_1742);
xor U3629 (N_3629,N_491,N_1272);
nor U3630 (N_3630,N_1182,N_426);
and U3631 (N_3631,N_1251,N_535);
nand U3632 (N_3632,N_58,N_295);
nand U3633 (N_3633,N_970,N_1238);
nand U3634 (N_3634,N_1756,N_510);
and U3635 (N_3635,N_1895,N_1267);
xor U3636 (N_3636,N_1138,N_1631);
nand U3637 (N_3637,N_1419,N_1373);
xnor U3638 (N_3638,N_1392,N_1157);
nand U3639 (N_3639,N_676,N_396);
or U3640 (N_3640,N_286,N_1420);
and U3641 (N_3641,N_156,N_1079);
nor U3642 (N_3642,N_1790,N_217);
nor U3643 (N_3643,N_897,N_847);
nor U3644 (N_3644,N_275,N_641);
xor U3645 (N_3645,N_55,N_696);
nor U3646 (N_3646,N_1578,N_1656);
nor U3647 (N_3647,N_421,N_273);
nor U3648 (N_3648,N_1856,N_1594);
xnor U3649 (N_3649,N_1188,N_851);
xor U3650 (N_3650,N_1060,N_535);
nand U3651 (N_3651,N_1873,N_1786);
or U3652 (N_3652,N_761,N_667);
or U3653 (N_3653,N_274,N_944);
or U3654 (N_3654,N_940,N_1599);
and U3655 (N_3655,N_948,N_401);
or U3656 (N_3656,N_1519,N_874);
and U3657 (N_3657,N_1220,N_267);
nor U3658 (N_3658,N_1110,N_787);
nand U3659 (N_3659,N_194,N_1825);
xnor U3660 (N_3660,N_1337,N_813);
nand U3661 (N_3661,N_909,N_1223);
or U3662 (N_3662,N_1073,N_1310);
xor U3663 (N_3663,N_609,N_499);
and U3664 (N_3664,N_1459,N_1439);
nand U3665 (N_3665,N_1496,N_933);
nor U3666 (N_3666,N_77,N_1125);
or U3667 (N_3667,N_1571,N_890);
nor U3668 (N_3668,N_526,N_95);
or U3669 (N_3669,N_1584,N_112);
and U3670 (N_3670,N_1394,N_1118);
xnor U3671 (N_3671,N_193,N_1563);
and U3672 (N_3672,N_920,N_1380);
or U3673 (N_3673,N_384,N_1370);
and U3674 (N_3674,N_716,N_692);
nand U3675 (N_3675,N_714,N_957);
and U3676 (N_3676,N_1558,N_77);
or U3677 (N_3677,N_193,N_1261);
or U3678 (N_3678,N_1518,N_1572);
nand U3679 (N_3679,N_155,N_965);
nand U3680 (N_3680,N_1135,N_229);
xnor U3681 (N_3681,N_1855,N_1499);
nand U3682 (N_3682,N_317,N_120);
nand U3683 (N_3683,N_924,N_1856);
nand U3684 (N_3684,N_1429,N_1247);
nand U3685 (N_3685,N_1012,N_1381);
nand U3686 (N_3686,N_781,N_242);
nand U3687 (N_3687,N_418,N_1000);
nand U3688 (N_3688,N_867,N_1049);
nor U3689 (N_3689,N_1866,N_1890);
nor U3690 (N_3690,N_194,N_1166);
or U3691 (N_3691,N_1648,N_301);
xnor U3692 (N_3692,N_1177,N_1302);
or U3693 (N_3693,N_816,N_1490);
and U3694 (N_3694,N_1231,N_691);
or U3695 (N_3695,N_1103,N_25);
xor U3696 (N_3696,N_1585,N_1841);
nand U3697 (N_3697,N_1417,N_1442);
or U3698 (N_3698,N_1044,N_601);
and U3699 (N_3699,N_744,N_201);
and U3700 (N_3700,N_1501,N_1629);
or U3701 (N_3701,N_1317,N_1984);
xnor U3702 (N_3702,N_739,N_916);
and U3703 (N_3703,N_1949,N_387);
xnor U3704 (N_3704,N_1756,N_1478);
nand U3705 (N_3705,N_801,N_1204);
nor U3706 (N_3706,N_1621,N_1785);
and U3707 (N_3707,N_26,N_1794);
xnor U3708 (N_3708,N_1565,N_1997);
nand U3709 (N_3709,N_1715,N_1676);
and U3710 (N_3710,N_1415,N_876);
and U3711 (N_3711,N_372,N_935);
xnor U3712 (N_3712,N_1699,N_318);
or U3713 (N_3713,N_913,N_615);
and U3714 (N_3714,N_17,N_1268);
xor U3715 (N_3715,N_766,N_126);
or U3716 (N_3716,N_999,N_615);
nor U3717 (N_3717,N_1442,N_723);
and U3718 (N_3718,N_696,N_955);
or U3719 (N_3719,N_1159,N_1268);
nand U3720 (N_3720,N_88,N_1354);
and U3721 (N_3721,N_129,N_133);
nor U3722 (N_3722,N_483,N_431);
or U3723 (N_3723,N_436,N_635);
or U3724 (N_3724,N_169,N_174);
or U3725 (N_3725,N_269,N_416);
nand U3726 (N_3726,N_1874,N_580);
nor U3727 (N_3727,N_1643,N_49);
and U3728 (N_3728,N_1773,N_347);
and U3729 (N_3729,N_1753,N_1502);
nor U3730 (N_3730,N_1670,N_838);
and U3731 (N_3731,N_67,N_228);
nand U3732 (N_3732,N_1226,N_581);
or U3733 (N_3733,N_967,N_358);
or U3734 (N_3734,N_511,N_471);
nor U3735 (N_3735,N_818,N_1824);
and U3736 (N_3736,N_596,N_516);
or U3737 (N_3737,N_702,N_1059);
nand U3738 (N_3738,N_1530,N_561);
nand U3739 (N_3739,N_393,N_250);
or U3740 (N_3740,N_1374,N_818);
nand U3741 (N_3741,N_90,N_407);
or U3742 (N_3742,N_277,N_1038);
or U3743 (N_3743,N_1238,N_1929);
and U3744 (N_3744,N_455,N_1547);
and U3745 (N_3745,N_1936,N_1440);
nor U3746 (N_3746,N_1322,N_626);
nor U3747 (N_3747,N_534,N_1784);
xnor U3748 (N_3748,N_784,N_520);
and U3749 (N_3749,N_485,N_1503);
nor U3750 (N_3750,N_1455,N_661);
nand U3751 (N_3751,N_1538,N_913);
or U3752 (N_3752,N_1521,N_1441);
nand U3753 (N_3753,N_388,N_669);
or U3754 (N_3754,N_1037,N_1340);
or U3755 (N_3755,N_188,N_1121);
or U3756 (N_3756,N_450,N_1405);
nand U3757 (N_3757,N_1282,N_1881);
and U3758 (N_3758,N_271,N_810);
xor U3759 (N_3759,N_291,N_208);
and U3760 (N_3760,N_1546,N_159);
or U3761 (N_3761,N_773,N_1733);
nor U3762 (N_3762,N_803,N_314);
or U3763 (N_3763,N_1293,N_596);
nor U3764 (N_3764,N_538,N_26);
nand U3765 (N_3765,N_1155,N_1741);
and U3766 (N_3766,N_1634,N_1852);
or U3767 (N_3767,N_1122,N_1733);
or U3768 (N_3768,N_252,N_1448);
or U3769 (N_3769,N_1701,N_1862);
nand U3770 (N_3770,N_448,N_251);
nor U3771 (N_3771,N_588,N_1571);
xor U3772 (N_3772,N_244,N_1007);
nor U3773 (N_3773,N_1622,N_435);
or U3774 (N_3774,N_1300,N_726);
nor U3775 (N_3775,N_1566,N_893);
or U3776 (N_3776,N_548,N_663);
or U3777 (N_3777,N_1376,N_20);
nand U3778 (N_3778,N_1700,N_454);
nor U3779 (N_3779,N_353,N_9);
nor U3780 (N_3780,N_1567,N_144);
nand U3781 (N_3781,N_1064,N_803);
xor U3782 (N_3782,N_319,N_1263);
nand U3783 (N_3783,N_1189,N_1761);
or U3784 (N_3784,N_587,N_567);
or U3785 (N_3785,N_1493,N_781);
xor U3786 (N_3786,N_1743,N_1947);
or U3787 (N_3787,N_738,N_351);
nand U3788 (N_3788,N_1256,N_1430);
and U3789 (N_3789,N_1438,N_1961);
or U3790 (N_3790,N_658,N_981);
xnor U3791 (N_3791,N_921,N_1590);
and U3792 (N_3792,N_1974,N_1357);
nand U3793 (N_3793,N_190,N_994);
and U3794 (N_3794,N_1690,N_166);
xnor U3795 (N_3795,N_1253,N_851);
nand U3796 (N_3796,N_1122,N_1289);
nand U3797 (N_3797,N_1283,N_1106);
nand U3798 (N_3798,N_1041,N_1992);
xnor U3799 (N_3799,N_503,N_832);
xor U3800 (N_3800,N_1224,N_659);
nor U3801 (N_3801,N_1680,N_370);
nor U3802 (N_3802,N_725,N_155);
xor U3803 (N_3803,N_1012,N_1944);
or U3804 (N_3804,N_17,N_1607);
or U3805 (N_3805,N_236,N_1075);
xor U3806 (N_3806,N_1722,N_1076);
nand U3807 (N_3807,N_1676,N_103);
or U3808 (N_3808,N_1681,N_191);
nor U3809 (N_3809,N_1292,N_1637);
nand U3810 (N_3810,N_96,N_872);
or U3811 (N_3811,N_1985,N_1401);
nor U3812 (N_3812,N_1823,N_751);
and U3813 (N_3813,N_803,N_924);
and U3814 (N_3814,N_760,N_135);
xnor U3815 (N_3815,N_1383,N_1197);
xor U3816 (N_3816,N_1255,N_124);
nor U3817 (N_3817,N_1974,N_1661);
nand U3818 (N_3818,N_171,N_588);
nand U3819 (N_3819,N_28,N_681);
xnor U3820 (N_3820,N_1094,N_485);
nor U3821 (N_3821,N_635,N_1528);
xnor U3822 (N_3822,N_132,N_60);
nor U3823 (N_3823,N_1623,N_1073);
nor U3824 (N_3824,N_1572,N_633);
nor U3825 (N_3825,N_1338,N_1773);
xnor U3826 (N_3826,N_47,N_1949);
or U3827 (N_3827,N_1975,N_1120);
and U3828 (N_3828,N_1159,N_1697);
nor U3829 (N_3829,N_68,N_1985);
or U3830 (N_3830,N_1829,N_1714);
or U3831 (N_3831,N_1893,N_893);
xnor U3832 (N_3832,N_1929,N_470);
nand U3833 (N_3833,N_1649,N_630);
nor U3834 (N_3834,N_273,N_737);
nor U3835 (N_3835,N_1236,N_81);
nand U3836 (N_3836,N_780,N_215);
or U3837 (N_3837,N_1558,N_231);
nand U3838 (N_3838,N_418,N_1515);
nor U3839 (N_3839,N_1253,N_1163);
xor U3840 (N_3840,N_797,N_530);
nand U3841 (N_3841,N_655,N_1780);
or U3842 (N_3842,N_144,N_550);
or U3843 (N_3843,N_920,N_1012);
nor U3844 (N_3844,N_1061,N_157);
xnor U3845 (N_3845,N_1734,N_138);
and U3846 (N_3846,N_1448,N_1308);
xor U3847 (N_3847,N_165,N_1503);
xnor U3848 (N_3848,N_1744,N_348);
xor U3849 (N_3849,N_30,N_1087);
and U3850 (N_3850,N_1958,N_556);
nor U3851 (N_3851,N_675,N_1449);
nand U3852 (N_3852,N_1682,N_771);
nor U3853 (N_3853,N_1890,N_1744);
or U3854 (N_3854,N_6,N_1191);
nor U3855 (N_3855,N_1324,N_991);
and U3856 (N_3856,N_488,N_325);
and U3857 (N_3857,N_1791,N_529);
nand U3858 (N_3858,N_1642,N_906);
and U3859 (N_3859,N_1959,N_1617);
xnor U3860 (N_3860,N_307,N_1792);
nor U3861 (N_3861,N_725,N_645);
xnor U3862 (N_3862,N_1507,N_1137);
and U3863 (N_3863,N_793,N_1199);
or U3864 (N_3864,N_1031,N_1435);
xnor U3865 (N_3865,N_788,N_1236);
and U3866 (N_3866,N_393,N_484);
nor U3867 (N_3867,N_1773,N_582);
xor U3868 (N_3868,N_973,N_785);
or U3869 (N_3869,N_546,N_500);
nor U3870 (N_3870,N_1742,N_1078);
or U3871 (N_3871,N_1498,N_1059);
nand U3872 (N_3872,N_298,N_136);
and U3873 (N_3873,N_1404,N_1001);
nor U3874 (N_3874,N_1541,N_1604);
nor U3875 (N_3875,N_878,N_1596);
xnor U3876 (N_3876,N_1438,N_923);
or U3877 (N_3877,N_571,N_363);
nor U3878 (N_3878,N_1058,N_330);
xor U3879 (N_3879,N_419,N_1710);
and U3880 (N_3880,N_1427,N_1148);
nand U3881 (N_3881,N_1828,N_808);
nor U3882 (N_3882,N_1204,N_1657);
xnor U3883 (N_3883,N_1419,N_88);
nor U3884 (N_3884,N_937,N_99);
nand U3885 (N_3885,N_1684,N_1025);
nor U3886 (N_3886,N_556,N_1074);
nor U3887 (N_3887,N_1631,N_1236);
nand U3888 (N_3888,N_1669,N_663);
nor U3889 (N_3889,N_817,N_1067);
xor U3890 (N_3890,N_1415,N_1124);
nand U3891 (N_3891,N_929,N_1153);
xor U3892 (N_3892,N_578,N_235);
or U3893 (N_3893,N_582,N_785);
nand U3894 (N_3894,N_1043,N_1466);
nand U3895 (N_3895,N_1718,N_1846);
or U3896 (N_3896,N_540,N_405);
nor U3897 (N_3897,N_1268,N_1442);
xnor U3898 (N_3898,N_360,N_279);
and U3899 (N_3899,N_736,N_1357);
or U3900 (N_3900,N_178,N_4);
or U3901 (N_3901,N_1937,N_1462);
nand U3902 (N_3902,N_1573,N_436);
and U3903 (N_3903,N_1572,N_1463);
and U3904 (N_3904,N_788,N_491);
or U3905 (N_3905,N_513,N_1160);
and U3906 (N_3906,N_570,N_1075);
nor U3907 (N_3907,N_1573,N_1586);
nand U3908 (N_3908,N_267,N_174);
nor U3909 (N_3909,N_1058,N_587);
nor U3910 (N_3910,N_309,N_1573);
and U3911 (N_3911,N_1863,N_1583);
and U3912 (N_3912,N_1593,N_9);
nand U3913 (N_3913,N_1726,N_1775);
or U3914 (N_3914,N_1985,N_291);
nand U3915 (N_3915,N_993,N_1662);
or U3916 (N_3916,N_949,N_699);
and U3917 (N_3917,N_650,N_924);
xor U3918 (N_3918,N_1505,N_1293);
xnor U3919 (N_3919,N_104,N_9);
and U3920 (N_3920,N_1246,N_1807);
and U3921 (N_3921,N_1778,N_79);
nand U3922 (N_3922,N_1969,N_800);
or U3923 (N_3923,N_622,N_34);
xnor U3924 (N_3924,N_733,N_1481);
or U3925 (N_3925,N_292,N_984);
and U3926 (N_3926,N_181,N_1514);
xor U3927 (N_3927,N_1413,N_1071);
xnor U3928 (N_3928,N_767,N_1457);
nand U3929 (N_3929,N_1857,N_68);
or U3930 (N_3930,N_1307,N_800);
xor U3931 (N_3931,N_769,N_289);
or U3932 (N_3932,N_1689,N_1316);
nor U3933 (N_3933,N_85,N_1944);
xnor U3934 (N_3934,N_1395,N_1831);
xnor U3935 (N_3935,N_227,N_292);
and U3936 (N_3936,N_580,N_1945);
xor U3937 (N_3937,N_1495,N_1747);
xor U3938 (N_3938,N_1410,N_659);
nor U3939 (N_3939,N_229,N_1088);
and U3940 (N_3940,N_279,N_1966);
and U3941 (N_3941,N_410,N_1352);
xnor U3942 (N_3942,N_811,N_30);
xor U3943 (N_3943,N_1303,N_534);
or U3944 (N_3944,N_1909,N_317);
or U3945 (N_3945,N_1221,N_1420);
nor U3946 (N_3946,N_382,N_1834);
and U3947 (N_3947,N_1049,N_1694);
nor U3948 (N_3948,N_970,N_1986);
nor U3949 (N_3949,N_196,N_507);
nand U3950 (N_3950,N_1007,N_390);
nor U3951 (N_3951,N_1385,N_237);
xor U3952 (N_3952,N_1897,N_272);
or U3953 (N_3953,N_512,N_1387);
or U3954 (N_3954,N_1135,N_494);
or U3955 (N_3955,N_728,N_466);
and U3956 (N_3956,N_604,N_136);
nor U3957 (N_3957,N_899,N_145);
nand U3958 (N_3958,N_222,N_115);
nor U3959 (N_3959,N_1851,N_1584);
xnor U3960 (N_3960,N_1081,N_1692);
or U3961 (N_3961,N_1909,N_1452);
or U3962 (N_3962,N_9,N_832);
nor U3963 (N_3963,N_1635,N_637);
or U3964 (N_3964,N_337,N_391);
nand U3965 (N_3965,N_1957,N_1244);
nor U3966 (N_3966,N_932,N_1490);
nor U3967 (N_3967,N_763,N_651);
nand U3968 (N_3968,N_793,N_861);
nor U3969 (N_3969,N_1864,N_452);
xor U3970 (N_3970,N_1407,N_1864);
and U3971 (N_3971,N_765,N_388);
nand U3972 (N_3972,N_1057,N_371);
nand U3973 (N_3973,N_593,N_354);
or U3974 (N_3974,N_1028,N_1641);
nand U3975 (N_3975,N_1235,N_1292);
or U3976 (N_3976,N_1132,N_1098);
xor U3977 (N_3977,N_1438,N_1371);
xnor U3978 (N_3978,N_1010,N_820);
or U3979 (N_3979,N_1788,N_1234);
nor U3980 (N_3980,N_722,N_85);
nor U3981 (N_3981,N_1793,N_671);
nand U3982 (N_3982,N_689,N_934);
nand U3983 (N_3983,N_1700,N_1843);
nand U3984 (N_3984,N_1766,N_202);
and U3985 (N_3985,N_1946,N_1971);
nor U3986 (N_3986,N_1559,N_55);
nor U3987 (N_3987,N_636,N_451);
or U3988 (N_3988,N_328,N_1252);
and U3989 (N_3989,N_667,N_914);
or U3990 (N_3990,N_176,N_730);
and U3991 (N_3991,N_1426,N_126);
xnor U3992 (N_3992,N_1048,N_105);
xor U3993 (N_3993,N_782,N_101);
and U3994 (N_3994,N_468,N_303);
and U3995 (N_3995,N_1524,N_559);
and U3996 (N_3996,N_1862,N_207);
xnor U3997 (N_3997,N_1394,N_473);
nand U3998 (N_3998,N_1557,N_1510);
nor U3999 (N_3999,N_204,N_369);
and U4000 (N_4000,N_2085,N_2853);
nor U4001 (N_4001,N_2268,N_3294);
nor U4002 (N_4002,N_2764,N_2871);
or U4003 (N_4003,N_2667,N_3930);
and U4004 (N_4004,N_3380,N_3298);
nand U4005 (N_4005,N_3467,N_2478);
nand U4006 (N_4006,N_3046,N_2099);
or U4007 (N_4007,N_3417,N_3780);
or U4008 (N_4008,N_3256,N_2513);
nand U4009 (N_4009,N_3817,N_3051);
nor U4010 (N_4010,N_2790,N_2011);
nand U4011 (N_4011,N_3798,N_3788);
nand U4012 (N_4012,N_2287,N_2492);
and U4013 (N_4013,N_3497,N_2774);
nor U4014 (N_4014,N_2383,N_3522);
and U4015 (N_4015,N_3992,N_3269);
nor U4016 (N_4016,N_3106,N_3213);
nand U4017 (N_4017,N_2999,N_3799);
or U4018 (N_4018,N_3535,N_3323);
xor U4019 (N_4019,N_2658,N_3519);
nor U4020 (N_4020,N_2425,N_3361);
nor U4021 (N_4021,N_2820,N_2054);
nor U4022 (N_4022,N_2012,N_2958);
or U4023 (N_4023,N_3072,N_2750);
xnor U4024 (N_4024,N_2039,N_2541);
xor U4025 (N_4025,N_3069,N_2595);
xnor U4026 (N_4026,N_2980,N_3291);
and U4027 (N_4027,N_2118,N_3881);
nand U4028 (N_4028,N_3452,N_3117);
or U4029 (N_4029,N_2366,N_2622);
and U4030 (N_4030,N_2198,N_3946);
nor U4031 (N_4031,N_2013,N_3325);
xnor U4032 (N_4032,N_2866,N_2852);
xor U4033 (N_4033,N_3561,N_3065);
nand U4034 (N_4034,N_3079,N_3095);
nor U4035 (N_4035,N_2452,N_3469);
or U4036 (N_4036,N_3709,N_3237);
nor U4037 (N_4037,N_2566,N_2361);
or U4038 (N_4038,N_3114,N_3701);
xnor U4039 (N_4039,N_3165,N_3658);
nand U4040 (N_4040,N_2607,N_3133);
and U4041 (N_4041,N_3542,N_3883);
and U4042 (N_4042,N_3007,N_2426);
nor U4043 (N_4043,N_2728,N_3252);
or U4044 (N_4044,N_2526,N_3707);
or U4045 (N_4045,N_3887,N_3867);
nand U4046 (N_4046,N_2092,N_2620);
nor U4047 (N_4047,N_2134,N_3851);
nor U4048 (N_4048,N_3430,N_3878);
nand U4049 (N_4049,N_3692,N_2613);
and U4050 (N_4050,N_3124,N_2501);
and U4051 (N_4051,N_3951,N_2281);
xnor U4052 (N_4052,N_2831,N_3217);
xor U4053 (N_4053,N_3405,N_2090);
nor U4054 (N_4054,N_3498,N_3178);
xor U4055 (N_4055,N_3993,N_2982);
nand U4056 (N_4056,N_2377,N_3943);
nor U4057 (N_4057,N_2972,N_3604);
nor U4058 (N_4058,N_2941,N_3964);
and U4059 (N_4059,N_3110,N_3848);
xnor U4060 (N_4060,N_2898,N_3534);
xor U4061 (N_4061,N_3460,N_2989);
or U4062 (N_4062,N_2666,N_2060);
nor U4063 (N_4063,N_3232,N_2945);
nor U4064 (N_4064,N_2462,N_2807);
or U4065 (N_4065,N_3333,N_3419);
nor U4066 (N_4066,N_2741,N_2389);
nand U4067 (N_4067,N_3438,N_2202);
nand U4068 (N_4068,N_2496,N_2736);
nor U4069 (N_4069,N_2662,N_2149);
nor U4070 (N_4070,N_2307,N_3487);
xor U4071 (N_4071,N_3674,N_2178);
and U4072 (N_4072,N_2127,N_3465);
nor U4073 (N_4073,N_3281,N_3215);
or U4074 (N_4074,N_2507,N_3547);
nor U4075 (N_4075,N_2519,N_2598);
nand U4076 (N_4076,N_2890,N_3462);
xor U4077 (N_4077,N_2348,N_3698);
or U4078 (N_4078,N_3950,N_2991);
or U4079 (N_4079,N_2376,N_3092);
nor U4080 (N_4080,N_2318,N_3713);
xnor U4081 (N_4081,N_3546,N_2707);
nor U4082 (N_4082,N_3440,N_2182);
nand U4083 (N_4083,N_3821,N_2749);
xor U4084 (N_4084,N_3398,N_3639);
nand U4085 (N_4085,N_2035,N_3394);
or U4086 (N_4086,N_2811,N_3379);
nand U4087 (N_4087,N_3491,N_3610);
nand U4088 (N_4088,N_3620,N_3180);
nand U4089 (N_4089,N_2649,N_2244);
or U4090 (N_4090,N_3279,N_2443);
or U4091 (N_4091,N_2734,N_2372);
or U4092 (N_4092,N_2485,N_2765);
nor U4093 (N_4093,N_2309,N_3345);
xor U4094 (N_4094,N_2763,N_2726);
nand U4095 (N_4095,N_2788,N_2909);
nor U4096 (N_4096,N_3302,N_2575);
or U4097 (N_4097,N_3933,N_2358);
and U4098 (N_4098,N_2881,N_3995);
xor U4099 (N_4099,N_2018,N_3927);
xor U4100 (N_4100,N_3742,N_3564);
nand U4101 (N_4101,N_3907,N_3598);
and U4102 (N_4102,N_3945,N_3810);
and U4103 (N_4103,N_3804,N_2861);
or U4104 (N_4104,N_3093,N_3349);
xor U4105 (N_4105,N_2642,N_3682);
nor U4106 (N_4106,N_2423,N_2283);
or U4107 (N_4107,N_2604,N_2023);
or U4108 (N_4108,N_2838,N_3724);
nand U4109 (N_4109,N_2296,N_2706);
xnor U4110 (N_4110,N_3515,N_3014);
or U4111 (N_4111,N_3317,N_3952);
nor U4112 (N_4112,N_2179,N_2711);
and U4113 (N_4113,N_3705,N_2094);
nor U4114 (N_4114,N_2534,N_2992);
nand U4115 (N_4115,N_2165,N_2556);
nor U4116 (N_4116,N_2248,N_3937);
xnor U4117 (N_4117,N_3406,N_3026);
or U4118 (N_4118,N_2834,N_2160);
and U4119 (N_4119,N_3550,N_3024);
nand U4120 (N_4120,N_2727,N_2238);
and U4121 (N_4121,N_2056,N_3665);
nand U4122 (N_4122,N_3220,N_3625);
nand U4123 (N_4123,N_2785,N_3488);
xor U4124 (N_4124,N_2457,N_3480);
nor U4125 (N_4125,N_3548,N_2282);
and U4126 (N_4126,N_3301,N_2122);
nor U4127 (N_4127,N_2091,N_3085);
nand U4128 (N_4128,N_2928,N_3594);
and U4129 (N_4129,N_3576,N_3310);
nand U4130 (N_4130,N_2276,N_2944);
and U4131 (N_4131,N_3496,N_3395);
nand U4132 (N_4132,N_2614,N_3805);
or U4133 (N_4133,N_2044,N_2180);
or U4134 (N_4134,N_2842,N_3882);
nand U4135 (N_4135,N_2812,N_3212);
nand U4136 (N_4136,N_3154,N_3533);
nor U4137 (N_4137,N_2596,N_3711);
and U4138 (N_4138,N_2747,N_3872);
or U4139 (N_4139,N_3344,N_2483);
and U4140 (N_4140,N_3649,N_3559);
or U4141 (N_4141,N_2223,N_3292);
or U4142 (N_4142,N_2632,N_2967);
and U4143 (N_4143,N_2494,N_3677);
nor U4144 (N_4144,N_3408,N_2095);
xor U4145 (N_4145,N_3094,N_3241);
and U4146 (N_4146,N_3222,N_2561);
nor U4147 (N_4147,N_3637,N_2137);
or U4148 (N_4148,N_2002,N_2200);
xor U4149 (N_4149,N_3869,N_2518);
and U4150 (N_4150,N_3048,N_2186);
nand U4151 (N_4151,N_2552,N_3544);
nand U4152 (N_4152,N_2136,N_3695);
xor U4153 (N_4153,N_3211,N_3941);
nor U4154 (N_4154,N_2337,N_3795);
and U4155 (N_4155,N_2690,N_2597);
or U4156 (N_4156,N_2684,N_2681);
nor U4157 (N_4157,N_2862,N_3012);
nand U4158 (N_4158,N_3486,N_3224);
and U4159 (N_4159,N_2675,N_3456);
or U4160 (N_4160,N_2610,N_3179);
xnor U4161 (N_4161,N_3131,N_2833);
nor U4162 (N_4162,N_2627,N_2919);
and U4163 (N_4163,N_3636,N_2147);
and U4164 (N_4164,N_2902,N_2123);
or U4165 (N_4165,N_2379,N_2752);
xor U4166 (N_4166,N_3870,N_3989);
xnor U4167 (N_4167,N_2599,N_3979);
nand U4168 (N_4168,N_3615,N_3797);
xnor U4169 (N_4169,N_2509,N_2738);
and U4170 (N_4170,N_2456,N_3953);
or U4171 (N_4171,N_2381,N_3647);
and U4172 (N_4172,N_3243,N_3088);
xor U4173 (N_4173,N_3410,N_3084);
nor U4174 (N_4174,N_2697,N_3808);
or U4175 (N_4175,N_2406,N_2638);
nand U4176 (N_4176,N_2336,N_3402);
nor U4177 (N_4177,N_3105,N_3028);
xor U4178 (N_4178,N_2399,N_3833);
nor U4179 (N_4179,N_2175,N_3322);
nor U4180 (N_4180,N_2105,N_2724);
nand U4181 (N_4181,N_3321,N_3512);
or U4182 (N_4182,N_2387,N_3538);
nor U4183 (N_4183,N_3573,N_3358);
nor U4184 (N_4184,N_3409,N_2077);
nor U4185 (N_4185,N_2959,N_3956);
or U4186 (N_4186,N_3645,N_2537);
nor U4187 (N_4187,N_3021,N_2592);
nand U4188 (N_4188,N_3142,N_3416);
and U4189 (N_4189,N_2289,N_2760);
nand U4190 (N_4190,N_3689,N_2663);
and U4191 (N_4191,N_3303,N_2395);
nand U4192 (N_4192,N_3109,N_2646);
xnor U4193 (N_4193,N_3511,N_3628);
or U4194 (N_4194,N_2292,N_3958);
xnor U4195 (N_4195,N_2647,N_3167);
nand U4196 (N_4196,N_2947,N_2643);
xor U4197 (N_4197,N_3924,N_3577);
and U4198 (N_4198,N_3818,N_3214);
and U4199 (N_4199,N_2181,N_2516);
or U4200 (N_4200,N_3599,N_2064);
and U4201 (N_4201,N_3976,N_2532);
nor U4202 (N_4202,N_3686,N_3068);
xnor U4203 (N_4203,N_2885,N_2975);
nor U4204 (N_4204,N_3146,N_2352);
nand U4205 (N_4205,N_3553,N_3827);
and U4206 (N_4206,N_3987,N_2653);
or U4207 (N_4207,N_2086,N_2657);
and U4208 (N_4208,N_2015,N_3514);
nand U4209 (N_4209,N_2199,N_3911);
nor U4210 (N_4210,N_2828,N_2355);
nand U4211 (N_4211,N_3499,N_2293);
or U4212 (N_4212,N_2045,N_3368);
nand U4213 (N_4213,N_2799,N_2994);
xor U4214 (N_4214,N_3735,N_2081);
and U4215 (N_4215,N_2824,N_2163);
xnor U4216 (N_4216,N_3441,N_3337);
and U4217 (N_4217,N_3016,N_2350);
nand U4218 (N_4218,N_2401,N_2326);
xor U4219 (N_4219,N_3740,N_3595);
nor U4220 (N_4220,N_2382,N_2708);
nor U4221 (N_4221,N_2264,N_2036);
and U4222 (N_4222,N_3009,N_3596);
nand U4223 (N_4223,N_2906,N_2347);
nand U4224 (N_4224,N_2792,N_2325);
nand U4225 (N_4225,N_3169,N_2404);
or U4226 (N_4226,N_2682,N_3889);
xor U4227 (N_4227,N_2611,N_3572);
or U4228 (N_4228,N_2024,N_3531);
xnor U4229 (N_4229,N_2428,N_2568);
xnor U4230 (N_4230,N_3994,N_3723);
nor U4231 (N_4231,N_2574,N_3503);
xor U4232 (N_4232,N_3928,N_2623);
nand U4233 (N_4233,N_2484,N_3374);
or U4234 (N_4234,N_3489,N_3721);
nor U4235 (N_4235,N_3308,N_3838);
and U4236 (N_4236,N_3540,N_3664);
or U4237 (N_4237,N_3904,N_3287);
nor U4238 (N_4238,N_3749,N_2508);
nor U4239 (N_4239,N_3173,N_2804);
and U4240 (N_4240,N_3988,N_2718);
and U4241 (N_4241,N_2965,N_3769);
nor U4242 (N_4242,N_2783,N_2710);
and U4243 (N_4243,N_3481,N_2315);
nand U4244 (N_4244,N_2413,N_3569);
xnor U4245 (N_4245,N_2071,N_3900);
and U4246 (N_4246,N_3171,N_2939);
or U4247 (N_4247,N_2761,N_2052);
xnor U4248 (N_4248,N_2261,N_3874);
nand U4249 (N_4249,N_3074,N_3143);
nand U4250 (N_4250,N_2059,N_3717);
nand U4251 (N_4251,N_2089,N_3790);
and U4252 (N_4252,N_3737,N_2083);
nand U4253 (N_4253,N_3209,N_3318);
nand U4254 (N_4254,N_2343,N_2290);
xor U4255 (N_4255,N_3013,N_2116);
or U4256 (N_4256,N_2349,N_2733);
and U4257 (N_4257,N_2897,N_3836);
or U4258 (N_4258,N_3841,N_3612);
nor U4259 (N_4259,N_3244,N_3255);
xnor U4260 (N_4260,N_2161,N_2988);
xnor U4261 (N_4261,N_2243,N_2873);
and U4262 (N_4262,N_2633,N_2530);
and U4263 (N_4263,N_2709,N_3120);
xor U4264 (N_4264,N_3376,N_2856);
nand U4265 (N_4265,N_2584,N_2234);
nand U4266 (N_4266,N_3475,N_2998);
nand U4267 (N_4267,N_3396,N_2419);
and U4268 (N_4268,N_3485,N_3034);
and U4269 (N_4269,N_2275,N_2335);
and U4270 (N_4270,N_2021,N_3254);
or U4271 (N_4271,N_3585,N_2970);
nand U4272 (N_4272,N_2170,N_2801);
or U4273 (N_4273,N_3083,N_3917);
nor U4274 (N_4274,N_3231,N_2380);
nor U4275 (N_4275,N_2976,N_3570);
nand U4276 (N_4276,N_2864,N_2194);
or U4277 (N_4277,N_2969,N_2590);
nand U4278 (N_4278,N_2886,N_3446);
nand U4279 (N_4279,N_2114,N_2961);
and U4280 (N_4280,N_3293,N_2061);
nor U4281 (N_4281,N_2816,N_2257);
and U4282 (N_4282,N_3830,N_3815);
nand U4283 (N_4283,N_2051,N_3360);
nand U4284 (N_4284,N_2437,N_2087);
nor U4285 (N_4285,N_3066,N_3587);
and U4286 (N_4286,N_2628,N_2713);
and U4287 (N_4287,N_3736,N_3336);
nor U4288 (N_4288,N_2593,N_3918);
xor U4289 (N_4289,N_2907,N_3184);
and U4290 (N_4290,N_2735,N_3972);
and U4291 (N_4291,N_2030,N_2321);
nor U4292 (N_4292,N_2288,N_3159);
or U4293 (N_4293,N_3239,N_3329);
or U4294 (N_4294,N_2217,N_3306);
nand U4295 (N_4295,N_3706,N_3166);
xor U4296 (N_4296,N_3896,N_3346);
nor U4297 (N_4297,N_3839,N_2385);
xnor U4298 (N_4298,N_2922,N_2847);
and U4299 (N_4299,N_3565,N_3442);
xor U4300 (N_4300,N_2908,N_3716);
xnor U4301 (N_4301,N_3877,N_3632);
or U4302 (N_4302,N_3479,N_3875);
nor U4303 (N_4303,N_2803,N_3352);
or U4304 (N_4304,N_2910,N_2111);
or U4305 (N_4305,N_2522,N_2327);
and U4306 (N_4306,N_2344,N_2316);
or U4307 (N_4307,N_2931,N_2057);
nand U4308 (N_4308,N_2101,N_2434);
xor U4309 (N_4309,N_3247,N_2031);
and U4310 (N_4310,N_2600,N_2468);
or U4311 (N_4311,N_2211,N_3545);
nor U4312 (N_4312,N_2840,N_2313);
and U4313 (N_4313,N_3794,N_3055);
xor U4314 (N_4314,N_2514,N_3864);
and U4315 (N_4315,N_2798,N_3315);
or U4316 (N_4316,N_3053,N_2477);
xnor U4317 (N_4317,N_2544,N_2505);
nor U4318 (N_4318,N_3458,N_3132);
nor U4319 (N_4319,N_2974,N_3763);
nand U4320 (N_4320,N_2026,N_2453);
or U4321 (N_4321,N_3414,N_2677);
or U4322 (N_4322,N_2454,N_3865);
and U4323 (N_4323,N_3299,N_2010);
nand U4324 (N_4324,N_2725,N_3111);
nand U4325 (N_4325,N_2569,N_2768);
xor U4326 (N_4326,N_3773,N_2844);
xor U4327 (N_4327,N_2153,N_2210);
nand U4328 (N_4328,N_3603,N_3641);
and U4329 (N_4329,N_3746,N_3986);
or U4330 (N_4330,N_3957,N_2073);
nor U4331 (N_4331,N_2778,N_2096);
xor U4332 (N_4332,N_2656,N_3786);
xor U4333 (N_4333,N_2332,N_2331);
xor U4334 (N_4334,N_2701,N_2055);
or U4335 (N_4335,N_3835,N_2850);
or U4336 (N_4336,N_3283,N_2564);
and U4337 (N_4337,N_2417,N_3768);
xor U4338 (N_4338,N_2551,N_2324);
nor U4339 (N_4339,N_3385,N_3364);
or U4340 (N_4340,N_3863,N_2237);
nand U4341 (N_4341,N_3278,N_2040);
and U4342 (N_4342,N_2319,N_3353);
and U4343 (N_4343,N_3052,N_2767);
xor U4344 (N_4344,N_3858,N_3675);
and U4345 (N_4345,N_2305,N_3144);
nor U4346 (N_4346,N_2203,N_3050);
nand U4347 (N_4347,N_2692,N_3022);
and U4348 (N_4348,N_2363,N_3296);
and U4349 (N_4349,N_2762,N_2142);
nand U4350 (N_4350,N_2235,N_3605);
or U4351 (N_4351,N_3468,N_2354);
nor U4352 (N_4352,N_3999,N_2705);
or U4353 (N_4353,N_2263,N_2482);
xnor U4354 (N_4354,N_2185,N_2612);
nand U4355 (N_4355,N_3728,N_2860);
or U4356 (N_4356,N_2069,N_2571);
nor U4357 (N_4357,N_3152,N_2641);
or U4358 (N_4358,N_3560,N_2345);
or U4359 (N_4359,N_2849,N_3125);
xnor U4360 (N_4360,N_2639,N_3567);
or U4361 (N_4361,N_3582,N_2731);
nand U4362 (N_4362,N_2635,N_3849);
xor U4363 (N_4363,N_3776,N_2904);
and U4364 (N_4364,N_3648,N_2184);
xor U4365 (N_4365,N_2894,N_2751);
nand U4366 (N_4366,N_3549,N_3388);
or U4367 (N_4367,N_2365,N_2899);
and U4368 (N_4368,N_2841,N_3857);
nand U4369 (N_4369,N_3642,N_3473);
or U4370 (N_4370,N_2716,N_2351);
nor U4371 (N_4371,N_3562,N_3261);
xnor U4372 (N_4372,N_3873,N_3422);
or U4373 (N_4373,N_2837,N_2393);
xor U4374 (N_4374,N_3436,N_3777);
nand U4375 (N_4375,N_2102,N_2775);
and U4376 (N_4376,N_2278,N_2458);
and U4377 (N_4377,N_2151,N_2900);
xor U4378 (N_4378,N_2495,N_3043);
or U4379 (N_4379,N_3258,N_2594);
nor U4380 (N_4380,N_3655,N_2813);
xor U4381 (N_4381,N_3868,N_3973);
nor U4382 (N_4382,N_2895,N_2913);
nor U4383 (N_4383,N_2542,N_2493);
xnor U4384 (N_4384,N_3614,N_3340);
and U4385 (N_4385,N_2722,N_3206);
xnor U4386 (N_4386,N_2587,N_3734);
or U4387 (N_4387,N_2782,N_2949);
nand U4388 (N_4388,N_2250,N_2442);
nor U4389 (N_4389,N_3161,N_2191);
nor U4390 (N_4390,N_3025,N_2927);
xor U4391 (N_4391,N_3381,N_2397);
and U4392 (N_4392,N_2753,N_3676);
or U4393 (N_4393,N_3634,N_2815);
and U4394 (N_4394,N_3588,N_3495);
or U4395 (N_4395,N_3922,N_2481);
nand U4396 (N_4396,N_3850,N_3197);
or U4397 (N_4397,N_3741,N_3657);
nand U4398 (N_4398,N_2000,N_3899);
xor U4399 (N_4399,N_2872,N_2488);
and U4400 (N_4400,N_3983,N_3650);
and U4401 (N_4401,N_3704,N_3913);
or U4402 (N_4402,N_2424,N_2236);
or U4403 (N_4403,N_3947,N_2152);
nor U4404 (N_4404,N_2444,N_3163);
or U4405 (N_4405,N_2270,N_2131);
and U4406 (N_4406,N_3793,N_2414);
xnor U4407 (N_4407,N_2500,N_2121);
or U4408 (N_4408,N_3528,N_3201);
or U4409 (N_4409,N_3643,N_3807);
and U4410 (N_4410,N_2219,N_3493);
and U4411 (N_4411,N_2440,N_2227);
xnor U4412 (N_4412,N_2648,N_3929);
and U4413 (N_4413,N_3806,N_3203);
or U4414 (N_4414,N_3834,N_3482);
nand U4415 (N_4415,N_3425,N_3890);
or U4416 (N_4416,N_2075,N_2173);
nand U4417 (N_4417,N_3621,N_3242);
or U4418 (N_4418,N_2580,N_3627);
and U4419 (N_4419,N_3400,N_2323);
or U4420 (N_4420,N_3667,N_3792);
nand U4421 (N_4421,N_2698,N_3583);
or U4422 (N_4422,N_3775,N_2557);
nand U4423 (N_4423,N_2341,N_2626);
xor U4424 (N_4424,N_3392,N_2375);
or U4425 (N_4425,N_3448,N_3006);
nand U4426 (N_4426,N_3866,N_2957);
and U4427 (N_4427,N_2421,N_3432);
nand U4428 (N_4428,N_3193,N_3760);
and U4429 (N_4429,N_3502,N_3355);
nand U4430 (N_4430,N_2691,N_2043);
and U4431 (N_4431,N_2130,N_3801);
and U4432 (N_4432,N_3263,N_2441);
nor U4433 (N_4433,N_2362,N_3932);
nor U4434 (N_4434,N_2135,N_2249);
or U4435 (N_4435,N_3136,N_2814);
nand U4436 (N_4436,N_3977,N_3003);
or U4437 (N_4437,N_2269,N_2543);
nand U4438 (N_4438,N_2132,N_3811);
or U4439 (N_4439,N_3182,N_2167);
nand U4440 (N_4440,N_3731,N_2601);
nor U4441 (N_4441,N_3314,N_3871);
and U4442 (N_4442,N_2805,N_2112);
nor U4443 (N_4443,N_2929,N_3424);
or U4444 (N_4444,N_2531,N_3662);
and U4445 (N_4445,N_2286,N_3415);
and U4446 (N_4446,N_2322,N_2033);
and U4447 (N_4447,N_2515,N_2755);
xnor U4448 (N_4448,N_2960,N_3158);
nor U4449 (N_4449,N_2408,N_2356);
xor U4450 (N_4450,N_3524,N_2330);
xnor U4451 (N_4451,N_2963,N_2048);
or U4452 (N_4452,N_2744,N_3509);
and U4453 (N_4453,N_3238,N_3149);
xnor U4454 (N_4454,N_3919,N_3284);
and U4455 (N_4455,N_2088,N_3816);
or U4456 (N_4456,N_3134,N_2739);
and U4457 (N_4457,N_3663,N_2721);
or U4458 (N_4458,N_3608,N_3076);
xor U4459 (N_4459,N_3700,N_3463);
nand U4460 (N_4460,N_3991,N_3225);
xnor U4461 (N_4461,N_3812,N_2241);
nand U4462 (N_4462,N_2139,N_3885);
nor U4463 (N_4463,N_2978,N_3748);
and U4464 (N_4464,N_3348,N_3027);
nand U4465 (N_4465,N_3309,N_2480);
xor U4466 (N_4466,N_2209,N_3316);
nor U4467 (N_4467,N_2216,N_2328);
or U4468 (N_4468,N_3753,N_3304);
nor U4469 (N_4469,N_2757,N_3453);
or U4470 (N_4470,N_2588,N_2825);
nor U4471 (N_4471,N_2369,N_2025);
xnor U4472 (N_4472,N_2038,N_3529);
or U4473 (N_4473,N_2231,N_2986);
xor U4474 (N_4474,N_3579,N_3997);
nor U4475 (N_4475,N_2312,N_3350);
nand U4476 (N_4476,N_3008,N_3130);
xnor U4477 (N_4477,N_2213,N_3145);
xor U4478 (N_4478,N_3936,N_3845);
xor U4479 (N_4479,N_3483,N_2606);
xnor U4480 (N_4480,N_2683,N_2918);
and U4481 (N_4481,N_3556,N_3586);
and U4482 (N_4482,N_2390,N_2695);
or U4483 (N_4483,N_2171,N_2679);
and U4484 (N_4484,N_2702,N_2472);
nand U4485 (N_4485,N_3412,N_3445);
and U4486 (N_4486,N_2984,N_2113);
nand U4487 (N_4487,N_3045,N_2221);
xor U4488 (N_4488,N_2743,N_2933);
xnor U4489 (N_4489,N_3752,N_3060);
nand U4490 (N_4490,N_2545,N_2476);
and U4491 (N_4491,N_2370,N_3669);
nor U4492 (N_4492,N_2155,N_3508);
nand U4493 (N_4493,N_2388,N_3371);
xnor U4494 (N_4494,N_3277,N_2581);
and U4495 (N_4495,N_2993,N_3756);
nor U4496 (N_4496,N_2229,N_3824);
and U4497 (N_4497,N_3063,N_3273);
or U4498 (N_4498,N_3590,N_3326);
or U4499 (N_4499,N_2005,N_2891);
nor U4500 (N_4500,N_3673,N_3010);
nand U4501 (N_4501,N_3974,N_3591);
and U4502 (N_4502,N_3411,N_3127);
and U4503 (N_4503,N_2616,N_3981);
or U4504 (N_4504,N_3840,N_2981);
nand U4505 (N_4505,N_2636,N_2776);
nor U4506 (N_4506,N_3819,N_3341);
xor U4507 (N_4507,N_3901,N_2935);
nand U4508 (N_4508,N_2084,N_3948);
and U4509 (N_4509,N_2378,N_2072);
and U4510 (N_4510,N_2740,N_2859);
or U4511 (N_4511,N_3234,N_3847);
and U4512 (N_4512,N_3119,N_2197);
nand U4513 (N_4513,N_3905,N_3121);
and U4514 (N_4514,N_2915,N_3477);
or U4515 (N_4515,N_2037,N_2995);
xnor U4516 (N_4516,N_2644,N_3982);
or U4517 (N_4517,N_2800,N_3443);
nor U4518 (N_4518,N_3123,N_3955);
xnor U4519 (N_4519,N_2273,N_3574);
or U4520 (N_4520,N_3391,N_3190);
or U4521 (N_4521,N_3537,N_3581);
nor U4522 (N_4522,N_3478,N_3000);
nor U4523 (N_4523,N_3253,N_2830);
nand U4524 (N_4524,N_3172,N_3005);
or U4525 (N_4525,N_3399,N_2912);
xor U4526 (N_4526,N_3040,N_2391);
nand U4527 (N_4527,N_2570,N_2166);
nor U4528 (N_4528,N_2143,N_2810);
nand U4529 (N_4529,N_3802,N_3616);
or U4530 (N_4530,N_3101,N_2586);
or U4531 (N_4531,N_3061,N_3372);
nor U4532 (N_4532,N_2409,N_3039);
or U4533 (N_4533,N_3199,N_2070);
nand U4534 (N_4534,N_3726,N_3638);
or U4535 (N_4535,N_2074,N_2271);
and U4536 (N_4536,N_3272,N_3619);
xor U4537 (N_4537,N_2893,N_2789);
and U4538 (N_4538,N_3725,N_3837);
xor U4539 (N_4539,N_3099,N_2498);
and U4540 (N_4540,N_3520,N_2795);
xor U4541 (N_4541,N_3047,N_2857);
nand U4542 (N_4542,N_3710,N_2676);
or U4543 (N_4543,N_3020,N_2009);
or U4544 (N_4544,N_2979,N_2602);
or U4545 (N_4545,N_3970,N_2430);
xor U4546 (N_4546,N_3803,N_3687);
nor U4547 (N_4547,N_2068,N_2855);
nand U4548 (N_4548,N_2954,N_2572);
nor U4549 (N_4549,N_2342,N_3971);
xor U4550 (N_4550,N_2109,N_2934);
or U4551 (N_4551,N_2125,N_2003);
and U4552 (N_4552,N_2688,N_3832);
nand U4553 (N_4553,N_2615,N_3041);
nand U4554 (N_4554,N_3606,N_2098);
or U4555 (N_4555,N_2460,N_3139);
nand U4556 (N_4556,N_3831,N_3843);
nand U4557 (N_4557,N_3210,N_2863);
xnor U4558 (N_4558,N_3450,N_3334);
nand U4559 (N_4559,N_3397,N_3688);
and U4560 (N_4560,N_2374,N_3359);
xnor U4561 (N_4561,N_3939,N_3646);
nand U4562 (N_4562,N_2285,N_3037);
nor U4563 (N_4563,N_2432,N_2078);
nand U4564 (N_4564,N_2925,N_2272);
and U4565 (N_4565,N_2364,N_2650);
xor U4566 (N_4566,N_3787,N_3772);
and U4567 (N_4567,N_3789,N_2256);
and U4568 (N_4568,N_2433,N_3931);
xor U4569 (N_4569,N_2333,N_2867);
and U4570 (N_4570,N_3357,N_3200);
or U4571 (N_4571,N_3501,N_3954);
xor U4572 (N_4572,N_2188,N_2334);
or U4573 (N_4573,N_3476,N_2346);
and U4574 (N_4574,N_2156,N_3090);
xor U4575 (N_4575,N_2438,N_3030);
or U4576 (N_4576,N_2246,N_2884);
nand U4577 (N_4577,N_2461,N_3903);
and U4578 (N_4578,N_3282,N_2671);
nand U4579 (N_4579,N_3276,N_3343);
and U4580 (N_4580,N_2239,N_3738);
nand U4581 (N_4581,N_3204,N_3897);
nor U4582 (N_4582,N_3771,N_3207);
nor U4583 (N_4583,N_3386,N_2896);
nand U4584 (N_4584,N_2654,N_2138);
nand U4585 (N_4585,N_2554,N_3966);
or U4586 (N_4586,N_2512,N_3527);
xor U4587 (N_4587,N_3194,N_3920);
or U4588 (N_4588,N_2553,N_2962);
nor U4589 (N_4589,N_3510,N_3484);
xor U4590 (N_4590,N_3170,N_3653);
or U4591 (N_4591,N_3175,N_2809);
nor U4592 (N_4592,N_3285,N_3168);
and U4593 (N_4593,N_2067,N_2467);
nor U4594 (N_4594,N_3064,N_3312);
nand U4595 (N_4595,N_3855,N_3233);
or U4596 (N_4596,N_2529,N_2550);
nand U4597 (N_4597,N_2892,N_2260);
nor U4598 (N_4598,N_2669,N_3219);
and U4599 (N_4599,N_2533,N_3814);
nand U4600 (N_4600,N_3265,N_2119);
xnor U4601 (N_4601,N_3969,N_3494);
xnor U4602 (N_4602,N_3555,N_2524);
and U4603 (N_4603,N_2206,N_3525);
xnor U4604 (N_4604,N_2392,N_2538);
xor U4605 (N_4605,N_2106,N_3221);
or U4606 (N_4606,N_3563,N_3373);
xor U4607 (N_4607,N_3218,N_3668);
and U4608 (N_4608,N_3141,N_2159);
nand U4609 (N_4609,N_2422,N_2196);
nor U4610 (N_4610,N_2802,N_3058);
or U4611 (N_4611,N_3447,N_3800);
and U4612 (N_4612,N_2573,N_3062);
and U4613 (N_4613,N_2784,N_3192);
and U4614 (N_4614,N_3426,N_2201);
nand U4615 (N_4615,N_2817,N_3102);
nor U4616 (N_4616,N_2110,N_3418);
nand U4617 (N_4617,N_3551,N_3347);
nand U4618 (N_4618,N_3319,N_3137);
nand U4619 (N_4619,N_3332,N_2253);
nor U4620 (N_4620,N_3338,N_2266);
xor U4621 (N_4621,N_3474,N_2845);
or U4622 (N_4622,N_2558,N_2145);
xor U4623 (N_4623,N_2407,N_3774);
xnor U4624 (N_4624,N_3745,N_3428);
nand U4625 (N_4625,N_2546,N_2547);
xnor U4626 (N_4626,N_3331,N_2169);
nor U4627 (N_4627,N_3683,N_3019);
xor U4628 (N_4628,N_2228,N_3004);
and U4629 (N_4629,N_3829,N_3968);
xnor U4630 (N_4630,N_3086,N_3115);
or U4631 (N_4631,N_3859,N_2053);
nor U4632 (N_4632,N_3521,N_3626);
nand U4633 (N_4633,N_2310,N_3264);
xnor U4634 (N_4634,N_2506,N_3216);
nor U4635 (N_4635,N_3696,N_3906);
xor U4636 (N_4636,N_2129,N_2412);
or U4637 (N_4637,N_3195,N_3965);
nor U4638 (N_4638,N_2063,N_3978);
nand U4639 (N_4639,N_2001,N_3886);
nor U4640 (N_4640,N_2208,N_2793);
and U4641 (N_4641,N_3518,N_3071);
nor U4642 (N_4642,N_2420,N_3571);
and U4643 (N_4643,N_3313,N_2486);
and U4644 (N_4644,N_3162,N_3038);
and U4645 (N_4645,N_2511,N_3032);
or U4646 (N_4646,N_2042,N_2565);
nor U4647 (N_4647,N_2629,N_3393);
nand U4648 (N_4648,N_3543,N_2368);
or U4649 (N_4649,N_2771,N_2489);
nor U4650 (N_4650,N_2955,N_3733);
and U4651 (N_4651,N_3249,N_2589);
nand U4652 (N_4652,N_2359,N_2174);
nor U4653 (N_4653,N_2189,N_3081);
xor U4654 (N_4654,N_2766,N_2050);
nor U4655 (N_4655,N_2625,N_3635);
xor U4656 (N_4656,N_3506,N_3670);
or U4657 (N_4657,N_3297,N_2563);
nand U4658 (N_4658,N_2769,N_3435);
or U4659 (N_4659,N_3059,N_2193);
or U4660 (N_4660,N_2903,N_2146);
xor U4661 (N_4661,N_2339,N_2535);
or U4662 (N_4662,N_2353,N_2668);
xor U4663 (N_4663,N_2665,N_2259);
and U4664 (N_4664,N_3680,N_2664);
and U4665 (N_4665,N_2689,N_2966);
or U4666 (N_4666,N_2714,N_2338);
xor U4667 (N_4667,N_2464,N_2624);
or U4668 (N_4668,N_2888,N_2280);
nor U4669 (N_4669,N_2770,N_3327);
xnor U4670 (N_4670,N_2304,N_2497);
xnor U4671 (N_4671,N_2618,N_2704);
or U4672 (N_4672,N_2267,N_3504);
or U4673 (N_4673,N_3492,N_2007);
xnor U4674 (N_4674,N_3176,N_3286);
nor U4675 (N_4675,N_2373,N_2258);
nor U4676 (N_4676,N_3031,N_2445);
nand U4677 (N_4677,N_3324,N_2661);
nand U4678 (N_4678,N_3967,N_2694);
and U4679 (N_4679,N_2990,N_2415);
xnor U4680 (N_4680,N_2128,N_2527);
or U4681 (N_4681,N_2487,N_3690);
xor U4682 (N_4682,N_2712,N_3767);
and U4683 (N_4683,N_3597,N_3235);
and U4684 (N_4684,N_3305,N_3715);
and U4685 (N_4685,N_3075,N_3925);
xnor U4686 (N_4686,N_2400,N_2510);
nor U4687 (N_4687,N_3135,N_3378);
nor U4688 (N_4688,N_3098,N_2997);
nand U4689 (N_4689,N_3880,N_3893);
or U4690 (N_4690,N_2103,N_2473);
nor U4691 (N_4691,N_3684,N_2148);
nand U4692 (N_4692,N_3909,N_2192);
nand U4693 (N_4693,N_3714,N_3813);
nor U4694 (N_4694,N_2754,N_3472);
nand U4695 (N_4695,N_2796,N_3708);
xor U4696 (N_4696,N_2780,N_3910);
or U4697 (N_4697,N_2948,N_3914);
and U4698 (N_4698,N_2971,N_3148);
nand U4699 (N_4699,N_3250,N_3678);
nand U4700 (N_4700,N_2459,N_2218);
or U4701 (N_4701,N_3823,N_3963);
or U4702 (N_4702,N_2608,N_2555);
and U4703 (N_4703,N_2004,N_3017);
nor U4704 (N_4704,N_3681,N_3236);
and U4705 (N_4705,N_3782,N_2491);
and U4706 (N_4706,N_3082,N_3363);
nor U4707 (N_4707,N_2226,N_2823);
nand U4708 (N_4708,N_3765,N_3892);
or U4709 (N_4709,N_2357,N_2678);
xor U4710 (N_4710,N_2539,N_3722);
nor U4711 (N_4711,N_3434,N_3852);
and U4712 (N_4712,N_2047,N_2693);
nor U4713 (N_4713,N_3617,N_3470);
or U4714 (N_4714,N_3633,N_2080);
and U4715 (N_4715,N_2474,N_3661);
or U4716 (N_4716,N_2224,N_2742);
and U4717 (N_4717,N_2117,N_3274);
or U4718 (N_4718,N_3067,N_3001);
nand U4719 (N_4719,N_2028,N_3985);
nor U4720 (N_4720,N_2937,N_2670);
or U4721 (N_4721,N_2956,N_3825);
and U4722 (N_4722,N_3097,N_2603);
nor U4723 (N_4723,N_2940,N_2252);
and U4724 (N_4724,N_3023,N_2195);
and U4725 (N_4725,N_3600,N_3539);
nor U4726 (N_4726,N_2848,N_2066);
or U4727 (N_4727,N_2220,N_3362);
or U4728 (N_4728,N_3592,N_2806);
nor U4729 (N_4729,N_2205,N_3248);
and U4730 (N_4730,N_3116,N_2717);
xor U4731 (N_4731,N_3270,N_2839);
and U4732 (N_4732,N_2140,N_2887);
xnor U4733 (N_4733,N_3268,N_2582);
xnor U4734 (N_4734,N_2439,N_3744);
xnor U4735 (N_4735,N_3049,N_3153);
nor U4736 (N_4736,N_3070,N_2911);
nor U4737 (N_4737,N_2640,N_2384);
nand U4738 (N_4738,N_3764,N_3390);
nand U4739 (N_4739,N_2503,N_2133);
and U4740 (N_4740,N_2469,N_3589);
nand U4741 (N_4741,N_2475,N_3356);
nor U4742 (N_4742,N_2781,N_2818);
nand U4743 (N_4743,N_3500,N_2851);
and U4744 (N_4744,N_3654,N_2254);
xor U4745 (N_4745,N_2017,N_3601);
xor U4746 (N_4746,N_3575,N_2854);
nand U4747 (N_4747,N_2020,N_2204);
nand U4748 (N_4748,N_3940,N_3666);
nand U4749 (N_4749,N_2274,N_3240);
nor U4750 (N_4750,N_3516,N_3461);
nand U4751 (N_4751,N_3685,N_3862);
or U4752 (N_4752,N_3879,N_3389);
nand U4753 (N_4753,N_2973,N_2465);
xor U4754 (N_4754,N_2041,N_2162);
nor U4755 (N_4755,N_3113,N_3757);
and U4756 (N_4756,N_2540,N_2560);
or U4757 (N_4757,N_3747,N_3490);
xnor U4758 (N_4758,N_2521,N_3054);
and U4759 (N_4759,N_2920,N_2164);
nor U4760 (N_4760,N_3809,N_3433);
nand U4761 (N_4761,N_2977,N_2062);
and U4762 (N_4762,N_2396,N_2773);
nand U4763 (N_4763,N_2737,N_2504);
nor U4764 (N_4764,N_2405,N_2079);
nand U4765 (N_4765,N_2924,N_3584);
nand U4766 (N_4766,N_2049,N_3464);
and U4767 (N_4767,N_3157,N_2772);
nand U4768 (N_4768,N_2548,N_2846);
nand U4769 (N_4769,N_2297,N_3421);
and U4770 (N_4770,N_3342,N_2797);
nand U4771 (N_4771,N_3754,N_3087);
or U4772 (N_4772,N_3112,N_2964);
nand U4773 (N_4773,N_3245,N_2791);
xor U4774 (N_4774,N_3387,N_3762);
xor U4775 (N_4775,N_2411,N_2889);
and U4776 (N_4776,N_2499,N_3938);
or U4777 (N_4777,N_3962,N_2298);
nor U4778 (N_4778,N_2938,N_3750);
or U4779 (N_4779,N_2672,N_2150);
xnor U4780 (N_4780,N_2410,N_2076);
nand U4781 (N_4781,N_2230,N_3660);
xor U4782 (N_4782,N_2936,N_2299);
xor U4783 (N_4783,N_3697,N_2882);
nand U4784 (N_4784,N_2652,N_3078);
or U4785 (N_4785,N_3507,N_3727);
xnor U4786 (N_4786,N_3280,N_3884);
nor U4787 (N_4787,N_3290,N_3536);
or U4788 (N_4788,N_3513,N_3164);
nor U4789 (N_4789,N_3679,N_2758);
or U4790 (N_4790,N_2429,N_3781);
and U4791 (N_4791,N_2832,N_3459);
and U4792 (N_4792,N_3108,N_2014);
nor U4793 (N_4793,N_2046,N_3251);
nand U4794 (N_4794,N_2279,N_2247);
xnor U4795 (N_4795,N_2794,N_3652);
nor U4796 (N_4796,N_3311,N_3694);
and U4797 (N_4797,N_3126,N_2723);
or U4798 (N_4798,N_2284,N_3703);
and U4799 (N_4799,N_2868,N_2120);
xor U4800 (N_4800,N_3150,N_3128);
nand U4801 (N_4801,N_3934,N_3288);
nor U4802 (N_4802,N_2295,N_3826);
nand U4803 (N_4803,N_2065,N_3783);
nor U4804 (N_4804,N_2630,N_2987);
nor U4805 (N_4805,N_2865,N_2168);
nand U4806 (N_4806,N_3057,N_3187);
nor U4807 (N_4807,N_3205,N_2302);
and U4808 (N_4808,N_2877,N_3926);
xnor U4809 (N_4809,N_3365,N_2926);
nor U4810 (N_4810,N_3077,N_3672);
xnor U4811 (N_4811,N_3246,N_3260);
xor U4812 (N_4812,N_3923,N_2591);
xnor U4813 (N_4813,N_2619,N_3651);
nor U4814 (N_4814,N_2124,N_2436);
or U4815 (N_4815,N_2930,N_3844);
or U4816 (N_4816,N_3791,N_3100);
and U4817 (N_4817,N_3568,N_2471);
or U4818 (N_4818,N_2329,N_2100);
nor U4819 (N_4819,N_2386,N_3185);
and U4820 (N_4820,N_2836,N_2583);
xor U4821 (N_4821,N_3558,N_2416);
or U4822 (N_4822,N_2637,N_2659);
or U4823 (N_4823,N_3266,N_2746);
nor U4824 (N_4824,N_3607,N_3033);
nand U4825 (N_4825,N_3103,N_3915);
nand U4826 (N_4826,N_3407,N_2277);
and U4827 (N_4827,N_3761,N_2523);
or U4828 (N_4828,N_2869,N_2779);
nor U4829 (N_4829,N_2455,N_2144);
nand U4830 (N_4830,N_3729,N_2631);
nand U4831 (N_4831,N_2262,N_2108);
nor U4832 (N_4832,N_3147,N_3056);
and U4833 (N_4833,N_2008,N_2905);
xor U4834 (N_4834,N_3138,N_2034);
and U4835 (N_4835,N_3427,N_3384);
nor U4836 (N_4836,N_3449,N_2951);
nand U4837 (N_4837,N_3018,N_3856);
xnor U4838 (N_4838,N_2686,N_3593);
or U4839 (N_4839,N_3339,N_3895);
and U4840 (N_4840,N_3289,N_3259);
xor U4841 (N_4841,N_2645,N_3894);
xnor U4842 (N_4842,N_2634,N_3404);
xor U4843 (N_4843,N_2306,N_3640);
xnor U4844 (N_4844,N_2923,N_3779);
and U4845 (N_4845,N_2435,N_3613);
nand U4846 (N_4846,N_3718,N_2294);
and U4847 (N_4847,N_3751,N_3042);
nand U4848 (N_4848,N_2567,N_2605);
xnor U4849 (N_4849,N_3796,N_3949);
or U4850 (N_4850,N_3702,N_3228);
and U4851 (N_4851,N_3198,N_2255);
and U4852 (N_4852,N_2729,N_2158);
or U4853 (N_4853,N_2943,N_3189);
nand U4854 (N_4854,N_3623,N_2858);
and U4855 (N_4855,N_3860,N_2207);
and U4856 (N_4856,N_3403,N_3262);
and U4857 (N_4857,N_2371,N_3413);
xnor U4858 (N_4858,N_3377,N_2154);
nor U4859 (N_4859,N_3307,N_3523);
nand U4860 (N_4860,N_2748,N_3451);
and U4861 (N_4861,N_2621,N_3631);
xnor U4862 (N_4862,N_3720,N_3107);
or U4863 (N_4863,N_2450,N_3699);
and U4864 (N_4864,N_2696,N_2177);
nand U4865 (N_4865,N_2952,N_2579);
xor U4866 (N_4866,N_2730,N_3044);
nand U4867 (N_4867,N_2032,N_2914);
or U4868 (N_4868,N_3532,N_3908);
and U4869 (N_4869,N_3759,N_3975);
or U4870 (N_4870,N_3656,N_2777);
nor U4871 (N_4871,N_3898,N_2242);
or U4872 (N_4872,N_2968,N_3609);
xor U4873 (N_4873,N_3156,N_2921);
nor U4874 (N_4874,N_3335,N_2314);
and U4875 (N_4875,N_3758,N_2022);
nand U4876 (N_4876,N_2058,N_3719);
and U4877 (N_4877,N_3526,N_2402);
and U4878 (N_4878,N_3328,N_3630);
and U4879 (N_4879,N_3202,N_2917);
and U4880 (N_4880,N_2029,N_2006);
xor U4881 (N_4881,N_2418,N_3151);
nand U4882 (N_4882,N_2104,N_2950);
or U4883 (N_4883,N_2700,N_2536);
or U4884 (N_4884,N_3935,N_2617);
nor U4885 (N_4885,N_2732,N_3196);
or U4886 (N_4886,N_3557,N_3096);
and U4887 (N_4887,N_3002,N_3188);
and U4888 (N_4888,N_3996,N_2360);
nor U4889 (N_4889,N_2398,N_3778);
xor U4890 (N_4890,N_3853,N_2985);
or U4891 (N_4891,N_2157,N_2215);
and U4892 (N_4892,N_3842,N_3423);
xnor U4893 (N_4893,N_3820,N_3223);
xnor U4894 (N_4894,N_2880,N_3644);
nor U4895 (N_4895,N_3942,N_3622);
and U4896 (N_4896,N_3437,N_2448);
and U4897 (N_4897,N_3439,N_2183);
or U4898 (N_4898,N_3566,N_2082);
or U4899 (N_4899,N_2490,N_2502);
nand U4900 (N_4900,N_3770,N_3659);
or U4901 (N_4901,N_3104,N_2680);
nand U4902 (N_4902,N_3580,N_2367);
and U4903 (N_4903,N_3629,N_3229);
and U4904 (N_4904,N_2916,N_2525);
or U4905 (N_4905,N_2942,N_2576);
and U4906 (N_4906,N_2946,N_3618);
nand U4907 (N_4907,N_3208,N_2317);
xnor U4908 (N_4908,N_2685,N_2214);
or U4909 (N_4909,N_2651,N_3784);
or U4910 (N_4910,N_2827,N_3370);
nand U4911 (N_4911,N_2720,N_2233);
or U4912 (N_4912,N_2808,N_3624);
and U4913 (N_4913,N_2340,N_3155);
nand U4914 (N_4914,N_3375,N_2097);
nand U4915 (N_4915,N_2699,N_2212);
or U4916 (N_4916,N_3383,N_2687);
xnor U4917 (N_4917,N_3011,N_3320);
and U4918 (N_4918,N_2245,N_3382);
nor U4919 (N_4919,N_3191,N_2901);
or U4920 (N_4920,N_2300,N_3429);
nand U4921 (N_4921,N_3691,N_3257);
or U4922 (N_4922,N_3444,N_3118);
nand U4923 (N_4923,N_2427,N_2577);
nand U4924 (N_4924,N_2520,N_3401);
or U4925 (N_4925,N_2126,N_3822);
xor U4926 (N_4926,N_3015,N_2141);
nor U4927 (N_4927,N_3267,N_3990);
nand U4928 (N_4928,N_2835,N_3186);
and U4929 (N_4929,N_2019,N_3732);
nor U4930 (N_4930,N_2301,N_2016);
nor U4931 (N_4931,N_2585,N_2222);
xor U4932 (N_4932,N_3961,N_3122);
and U4933 (N_4933,N_3739,N_3888);
nor U4934 (N_4934,N_3089,N_3743);
and U4935 (N_4935,N_2176,N_2703);
xnor U4936 (N_4936,N_3902,N_3541);
or U4937 (N_4937,N_2311,N_3351);
xor U4938 (N_4938,N_3420,N_2883);
or U4939 (N_4939,N_2291,N_3366);
nor U4940 (N_4940,N_2822,N_3602);
xnor U4941 (N_4941,N_3080,N_3671);
nand U4942 (N_4942,N_3271,N_3230);
nor U4943 (N_4943,N_3073,N_2559);
and U4944 (N_4944,N_2983,N_3755);
nand U4945 (N_4945,N_3552,N_2303);
nand U4946 (N_4946,N_2875,N_3466);
and U4947 (N_4947,N_2187,N_3578);
nor U4948 (N_4948,N_3785,N_3998);
and U4949 (N_4949,N_3140,N_2549);
and U4950 (N_4950,N_2674,N_2715);
nand U4951 (N_4951,N_3029,N_2320);
xnor U4952 (N_4952,N_3854,N_2878);
or U4953 (N_4953,N_3330,N_2759);
xnor U4954 (N_4954,N_3455,N_2562);
xnor U4955 (N_4955,N_3369,N_3431);
nand U4956 (N_4956,N_2819,N_3960);
nand U4957 (N_4957,N_3530,N_3036);
and U4958 (N_4958,N_2403,N_2470);
nand U4959 (N_4959,N_3828,N_3454);
or U4960 (N_4960,N_2517,N_3980);
or U4961 (N_4961,N_3174,N_2451);
nand U4962 (N_4962,N_2953,N_2265);
and U4963 (N_4963,N_3891,N_3181);
nor U4964 (N_4964,N_2829,N_3984);
nand U4965 (N_4965,N_3091,N_2528);
nand U4966 (N_4966,N_2870,N_3354);
or U4967 (N_4967,N_2673,N_3227);
nor U4968 (N_4968,N_2115,N_2655);
xnor U4969 (N_4969,N_3457,N_2446);
or U4970 (N_4970,N_2609,N_2660);
nand U4971 (N_4971,N_3160,N_2874);
nand U4972 (N_4972,N_2308,N_2190);
or U4973 (N_4973,N_2996,N_2240);
or U4974 (N_4974,N_2787,N_3959);
and U4975 (N_4975,N_3295,N_2447);
or U4976 (N_4976,N_2879,N_3505);
and U4977 (N_4977,N_3035,N_3693);
nand U4978 (N_4978,N_2225,N_3554);
or U4979 (N_4979,N_3611,N_3912);
xor U4980 (N_4980,N_2786,N_2578);
nor U4981 (N_4981,N_2251,N_2027);
or U4982 (N_4982,N_2107,N_2745);
nor U4983 (N_4983,N_3944,N_3846);
nor U4984 (N_4984,N_3861,N_3177);
xor U4985 (N_4985,N_3129,N_2756);
xnor U4986 (N_4986,N_3730,N_3275);
or U4987 (N_4987,N_2821,N_2826);
nand U4988 (N_4988,N_2466,N_2876);
or U4989 (N_4989,N_3916,N_2932);
and U4990 (N_4990,N_3766,N_2449);
and U4991 (N_4991,N_3226,N_2172);
or U4992 (N_4992,N_2232,N_2719);
and U4993 (N_4993,N_3367,N_3300);
xor U4994 (N_4994,N_3517,N_3183);
and U4995 (N_4995,N_2479,N_3876);
nand U4996 (N_4996,N_2431,N_2843);
nor U4997 (N_4997,N_2463,N_3471);
or U4998 (N_4998,N_3921,N_3712);
nand U4999 (N_4999,N_2093,N_2394);
nor U5000 (N_5000,N_2238,N_3342);
and U5001 (N_5001,N_3855,N_3914);
or U5002 (N_5002,N_2528,N_3677);
and U5003 (N_5003,N_3253,N_3395);
and U5004 (N_5004,N_2850,N_3914);
xor U5005 (N_5005,N_3215,N_2982);
xnor U5006 (N_5006,N_3532,N_2980);
or U5007 (N_5007,N_2030,N_3146);
and U5008 (N_5008,N_3126,N_3845);
xor U5009 (N_5009,N_3920,N_2110);
and U5010 (N_5010,N_2166,N_2079);
nor U5011 (N_5011,N_3687,N_2150);
nor U5012 (N_5012,N_3413,N_2562);
nor U5013 (N_5013,N_3654,N_2531);
nor U5014 (N_5014,N_2101,N_2508);
nor U5015 (N_5015,N_3002,N_3310);
nor U5016 (N_5016,N_3544,N_3837);
or U5017 (N_5017,N_2116,N_2397);
and U5018 (N_5018,N_2835,N_2754);
nor U5019 (N_5019,N_2074,N_3891);
and U5020 (N_5020,N_3522,N_3732);
or U5021 (N_5021,N_2444,N_2987);
or U5022 (N_5022,N_2387,N_2148);
nand U5023 (N_5023,N_2172,N_3082);
and U5024 (N_5024,N_3551,N_2965);
and U5025 (N_5025,N_3272,N_2369);
xnor U5026 (N_5026,N_2206,N_2009);
or U5027 (N_5027,N_2899,N_2126);
nor U5028 (N_5028,N_3949,N_2749);
xor U5029 (N_5029,N_2373,N_2950);
nand U5030 (N_5030,N_3517,N_3864);
nand U5031 (N_5031,N_2555,N_2931);
nor U5032 (N_5032,N_2322,N_3709);
xnor U5033 (N_5033,N_2054,N_2109);
nor U5034 (N_5034,N_2618,N_3451);
nor U5035 (N_5035,N_3834,N_3305);
xor U5036 (N_5036,N_3399,N_3316);
nand U5037 (N_5037,N_2005,N_3785);
nor U5038 (N_5038,N_3497,N_2519);
or U5039 (N_5039,N_3474,N_2733);
nor U5040 (N_5040,N_2130,N_3284);
and U5041 (N_5041,N_2095,N_2626);
nor U5042 (N_5042,N_2827,N_2085);
nor U5043 (N_5043,N_2634,N_3870);
nand U5044 (N_5044,N_3576,N_3252);
nand U5045 (N_5045,N_3987,N_3008);
and U5046 (N_5046,N_3371,N_2856);
nand U5047 (N_5047,N_2795,N_2170);
nand U5048 (N_5048,N_3871,N_3302);
xnor U5049 (N_5049,N_2650,N_2136);
xnor U5050 (N_5050,N_3765,N_3764);
nor U5051 (N_5051,N_2441,N_3380);
or U5052 (N_5052,N_3869,N_3689);
and U5053 (N_5053,N_2891,N_2440);
nor U5054 (N_5054,N_3428,N_2234);
nor U5055 (N_5055,N_3360,N_3393);
and U5056 (N_5056,N_2849,N_3545);
nand U5057 (N_5057,N_3503,N_3219);
and U5058 (N_5058,N_3356,N_3192);
nand U5059 (N_5059,N_3484,N_3566);
nand U5060 (N_5060,N_3730,N_3859);
xor U5061 (N_5061,N_3962,N_2587);
and U5062 (N_5062,N_2344,N_2307);
and U5063 (N_5063,N_2935,N_2077);
or U5064 (N_5064,N_2430,N_3729);
or U5065 (N_5065,N_3569,N_2862);
nor U5066 (N_5066,N_2236,N_2306);
and U5067 (N_5067,N_2278,N_2921);
and U5068 (N_5068,N_2108,N_3994);
and U5069 (N_5069,N_2691,N_2235);
and U5070 (N_5070,N_2416,N_3603);
and U5071 (N_5071,N_2022,N_3660);
nand U5072 (N_5072,N_3261,N_3705);
or U5073 (N_5073,N_2905,N_2953);
xnor U5074 (N_5074,N_3316,N_3008);
and U5075 (N_5075,N_3706,N_3240);
or U5076 (N_5076,N_3170,N_3506);
xor U5077 (N_5077,N_2683,N_3663);
and U5078 (N_5078,N_2729,N_3910);
nand U5079 (N_5079,N_3706,N_3478);
nand U5080 (N_5080,N_3309,N_3784);
or U5081 (N_5081,N_2731,N_3713);
or U5082 (N_5082,N_2161,N_3062);
or U5083 (N_5083,N_3527,N_2038);
or U5084 (N_5084,N_3306,N_2211);
nand U5085 (N_5085,N_2082,N_2484);
nor U5086 (N_5086,N_2496,N_3967);
or U5087 (N_5087,N_3635,N_3232);
or U5088 (N_5088,N_3061,N_3220);
xnor U5089 (N_5089,N_3112,N_2235);
and U5090 (N_5090,N_2706,N_2861);
and U5091 (N_5091,N_2376,N_2461);
and U5092 (N_5092,N_2415,N_2088);
xor U5093 (N_5093,N_2474,N_3268);
nor U5094 (N_5094,N_2373,N_3721);
nor U5095 (N_5095,N_3383,N_3198);
xor U5096 (N_5096,N_2181,N_3472);
and U5097 (N_5097,N_3681,N_3176);
nand U5098 (N_5098,N_3360,N_3009);
and U5099 (N_5099,N_2348,N_2155);
nor U5100 (N_5100,N_3750,N_2097);
or U5101 (N_5101,N_3709,N_2198);
xnor U5102 (N_5102,N_2768,N_3734);
or U5103 (N_5103,N_3104,N_3809);
nand U5104 (N_5104,N_2055,N_2928);
nand U5105 (N_5105,N_2856,N_3751);
or U5106 (N_5106,N_3797,N_2936);
or U5107 (N_5107,N_3710,N_2529);
nor U5108 (N_5108,N_2852,N_2459);
xor U5109 (N_5109,N_2993,N_2493);
xnor U5110 (N_5110,N_3102,N_2233);
xnor U5111 (N_5111,N_2694,N_3634);
nor U5112 (N_5112,N_2136,N_2562);
nand U5113 (N_5113,N_2671,N_2962);
nand U5114 (N_5114,N_2569,N_2297);
nand U5115 (N_5115,N_3612,N_2168);
and U5116 (N_5116,N_2384,N_3381);
nor U5117 (N_5117,N_3018,N_2407);
nor U5118 (N_5118,N_3447,N_3370);
nand U5119 (N_5119,N_2371,N_3608);
and U5120 (N_5120,N_3141,N_2661);
nor U5121 (N_5121,N_2759,N_2896);
and U5122 (N_5122,N_3537,N_2498);
nor U5123 (N_5123,N_2145,N_3701);
nor U5124 (N_5124,N_3416,N_2968);
xnor U5125 (N_5125,N_2284,N_2773);
xnor U5126 (N_5126,N_2429,N_3351);
nand U5127 (N_5127,N_2910,N_2594);
xor U5128 (N_5128,N_2507,N_2757);
nor U5129 (N_5129,N_3400,N_2017);
xnor U5130 (N_5130,N_2392,N_2530);
and U5131 (N_5131,N_3417,N_2128);
nor U5132 (N_5132,N_3855,N_3412);
and U5133 (N_5133,N_3662,N_2505);
xnor U5134 (N_5134,N_2193,N_2129);
nand U5135 (N_5135,N_2440,N_2571);
nor U5136 (N_5136,N_3466,N_2626);
xnor U5137 (N_5137,N_2897,N_3866);
nor U5138 (N_5138,N_3339,N_2022);
nand U5139 (N_5139,N_3255,N_2840);
or U5140 (N_5140,N_2892,N_2290);
and U5141 (N_5141,N_3371,N_3846);
or U5142 (N_5142,N_3261,N_3971);
and U5143 (N_5143,N_3032,N_3540);
or U5144 (N_5144,N_3085,N_3302);
nand U5145 (N_5145,N_3373,N_2503);
xnor U5146 (N_5146,N_3957,N_3996);
or U5147 (N_5147,N_2408,N_3856);
and U5148 (N_5148,N_2459,N_3992);
nor U5149 (N_5149,N_3543,N_2181);
xnor U5150 (N_5150,N_3429,N_2843);
or U5151 (N_5151,N_3366,N_3270);
nor U5152 (N_5152,N_2692,N_2252);
nor U5153 (N_5153,N_3115,N_3959);
nor U5154 (N_5154,N_2963,N_2958);
or U5155 (N_5155,N_3786,N_3845);
or U5156 (N_5156,N_3279,N_3386);
nand U5157 (N_5157,N_2949,N_3435);
nor U5158 (N_5158,N_3797,N_2807);
nand U5159 (N_5159,N_3462,N_2031);
nand U5160 (N_5160,N_3519,N_2117);
or U5161 (N_5161,N_3839,N_3150);
nand U5162 (N_5162,N_3191,N_2917);
nor U5163 (N_5163,N_3070,N_3652);
xor U5164 (N_5164,N_2282,N_3159);
nor U5165 (N_5165,N_3274,N_3690);
and U5166 (N_5166,N_2517,N_2580);
and U5167 (N_5167,N_2187,N_2855);
nor U5168 (N_5168,N_2317,N_2793);
and U5169 (N_5169,N_3611,N_2334);
or U5170 (N_5170,N_3409,N_3764);
or U5171 (N_5171,N_3592,N_3902);
or U5172 (N_5172,N_2522,N_3100);
nand U5173 (N_5173,N_3836,N_3398);
or U5174 (N_5174,N_2380,N_3042);
nand U5175 (N_5175,N_2710,N_3751);
or U5176 (N_5176,N_2789,N_3403);
nor U5177 (N_5177,N_2352,N_2892);
and U5178 (N_5178,N_2522,N_3040);
xor U5179 (N_5179,N_3520,N_2579);
or U5180 (N_5180,N_3070,N_2882);
nor U5181 (N_5181,N_3368,N_2802);
xor U5182 (N_5182,N_3723,N_3366);
and U5183 (N_5183,N_2160,N_3794);
nor U5184 (N_5184,N_2473,N_3860);
nor U5185 (N_5185,N_2027,N_3297);
or U5186 (N_5186,N_2442,N_3049);
xor U5187 (N_5187,N_2323,N_2737);
or U5188 (N_5188,N_2827,N_2026);
nand U5189 (N_5189,N_3327,N_3153);
nor U5190 (N_5190,N_3471,N_3319);
nand U5191 (N_5191,N_2069,N_3799);
xnor U5192 (N_5192,N_3085,N_2588);
xor U5193 (N_5193,N_3668,N_3521);
xnor U5194 (N_5194,N_3104,N_2008);
nand U5195 (N_5195,N_3795,N_3829);
and U5196 (N_5196,N_3449,N_2096);
nand U5197 (N_5197,N_2516,N_2118);
or U5198 (N_5198,N_3534,N_3240);
nor U5199 (N_5199,N_2118,N_3774);
nor U5200 (N_5200,N_2091,N_2543);
and U5201 (N_5201,N_3013,N_3423);
xor U5202 (N_5202,N_3589,N_2236);
nor U5203 (N_5203,N_3265,N_3455);
xnor U5204 (N_5204,N_3300,N_3449);
or U5205 (N_5205,N_2448,N_2126);
nor U5206 (N_5206,N_3325,N_3585);
nor U5207 (N_5207,N_2792,N_2293);
nand U5208 (N_5208,N_3646,N_2978);
nand U5209 (N_5209,N_3188,N_3439);
nor U5210 (N_5210,N_2099,N_2360);
or U5211 (N_5211,N_3203,N_2465);
nand U5212 (N_5212,N_2401,N_3271);
or U5213 (N_5213,N_3809,N_3519);
or U5214 (N_5214,N_3706,N_3161);
or U5215 (N_5215,N_3078,N_2139);
or U5216 (N_5216,N_2755,N_2943);
xor U5217 (N_5217,N_3021,N_2941);
or U5218 (N_5218,N_3875,N_2497);
nand U5219 (N_5219,N_2268,N_2491);
nor U5220 (N_5220,N_2047,N_3126);
nand U5221 (N_5221,N_3321,N_3398);
xor U5222 (N_5222,N_2756,N_3622);
or U5223 (N_5223,N_2070,N_2453);
nand U5224 (N_5224,N_2958,N_3382);
nor U5225 (N_5225,N_3305,N_2391);
and U5226 (N_5226,N_3143,N_3602);
nand U5227 (N_5227,N_3057,N_3096);
and U5228 (N_5228,N_3629,N_2259);
xnor U5229 (N_5229,N_3551,N_3802);
or U5230 (N_5230,N_3777,N_2096);
nand U5231 (N_5231,N_3296,N_3192);
and U5232 (N_5232,N_2780,N_3084);
nor U5233 (N_5233,N_3425,N_2761);
or U5234 (N_5234,N_3309,N_2430);
or U5235 (N_5235,N_2160,N_3302);
or U5236 (N_5236,N_2960,N_2636);
nor U5237 (N_5237,N_2921,N_3353);
or U5238 (N_5238,N_3001,N_3114);
xor U5239 (N_5239,N_2260,N_2996);
and U5240 (N_5240,N_2375,N_3988);
or U5241 (N_5241,N_2029,N_3974);
or U5242 (N_5242,N_2766,N_3614);
and U5243 (N_5243,N_3386,N_2599);
and U5244 (N_5244,N_2929,N_3329);
nor U5245 (N_5245,N_3285,N_2423);
nor U5246 (N_5246,N_3583,N_2482);
nand U5247 (N_5247,N_3969,N_3285);
nand U5248 (N_5248,N_2688,N_3384);
nor U5249 (N_5249,N_3433,N_2548);
xor U5250 (N_5250,N_2621,N_3368);
xor U5251 (N_5251,N_3265,N_3994);
or U5252 (N_5252,N_3409,N_2508);
or U5253 (N_5253,N_3305,N_3872);
nand U5254 (N_5254,N_2705,N_3879);
nor U5255 (N_5255,N_2776,N_2886);
xnor U5256 (N_5256,N_2257,N_3769);
or U5257 (N_5257,N_3769,N_2557);
xor U5258 (N_5258,N_3104,N_3887);
nand U5259 (N_5259,N_2364,N_2470);
nor U5260 (N_5260,N_3387,N_2864);
nand U5261 (N_5261,N_3812,N_3082);
or U5262 (N_5262,N_2915,N_2574);
nand U5263 (N_5263,N_2247,N_2527);
and U5264 (N_5264,N_2734,N_2357);
nand U5265 (N_5265,N_2027,N_2692);
or U5266 (N_5266,N_3920,N_2059);
or U5267 (N_5267,N_2655,N_2044);
or U5268 (N_5268,N_3561,N_3849);
nand U5269 (N_5269,N_2758,N_3145);
nand U5270 (N_5270,N_2073,N_3072);
and U5271 (N_5271,N_2633,N_3927);
nand U5272 (N_5272,N_2455,N_2131);
nand U5273 (N_5273,N_3727,N_2650);
or U5274 (N_5274,N_3344,N_3306);
nor U5275 (N_5275,N_3468,N_3765);
or U5276 (N_5276,N_3515,N_2515);
or U5277 (N_5277,N_3645,N_2790);
nand U5278 (N_5278,N_3535,N_3906);
or U5279 (N_5279,N_3279,N_2062);
and U5280 (N_5280,N_2919,N_3106);
nand U5281 (N_5281,N_3132,N_2396);
or U5282 (N_5282,N_2061,N_3133);
or U5283 (N_5283,N_3209,N_2175);
nor U5284 (N_5284,N_2051,N_3584);
nor U5285 (N_5285,N_3333,N_2814);
and U5286 (N_5286,N_2578,N_3659);
and U5287 (N_5287,N_2242,N_2743);
nor U5288 (N_5288,N_2146,N_2752);
xnor U5289 (N_5289,N_2935,N_2036);
or U5290 (N_5290,N_2409,N_2186);
or U5291 (N_5291,N_2900,N_3524);
or U5292 (N_5292,N_2941,N_2970);
xnor U5293 (N_5293,N_2183,N_2361);
or U5294 (N_5294,N_3775,N_3439);
or U5295 (N_5295,N_2931,N_3253);
or U5296 (N_5296,N_2669,N_2331);
xnor U5297 (N_5297,N_2909,N_3708);
and U5298 (N_5298,N_2564,N_2065);
xor U5299 (N_5299,N_2170,N_3904);
or U5300 (N_5300,N_3982,N_3539);
nor U5301 (N_5301,N_3823,N_3599);
and U5302 (N_5302,N_3352,N_2981);
nor U5303 (N_5303,N_3932,N_2486);
nor U5304 (N_5304,N_2200,N_2962);
or U5305 (N_5305,N_3418,N_3019);
nand U5306 (N_5306,N_3964,N_2569);
nand U5307 (N_5307,N_3259,N_2532);
nor U5308 (N_5308,N_3508,N_3411);
nor U5309 (N_5309,N_2990,N_3672);
nor U5310 (N_5310,N_2621,N_2191);
or U5311 (N_5311,N_2348,N_2654);
nor U5312 (N_5312,N_3688,N_2026);
nand U5313 (N_5313,N_3575,N_3349);
nand U5314 (N_5314,N_3135,N_3010);
xor U5315 (N_5315,N_2421,N_2249);
xor U5316 (N_5316,N_3256,N_3647);
nor U5317 (N_5317,N_2560,N_2449);
nor U5318 (N_5318,N_3384,N_2482);
nand U5319 (N_5319,N_2962,N_3953);
or U5320 (N_5320,N_2183,N_2565);
nand U5321 (N_5321,N_3087,N_2006);
and U5322 (N_5322,N_3148,N_3709);
nor U5323 (N_5323,N_3918,N_2633);
xor U5324 (N_5324,N_2663,N_3762);
nand U5325 (N_5325,N_2202,N_2207);
xor U5326 (N_5326,N_2939,N_3060);
nand U5327 (N_5327,N_3936,N_2305);
xnor U5328 (N_5328,N_3782,N_2033);
nand U5329 (N_5329,N_2841,N_3088);
nand U5330 (N_5330,N_2682,N_3242);
and U5331 (N_5331,N_2924,N_2165);
or U5332 (N_5332,N_3441,N_2251);
nor U5333 (N_5333,N_3888,N_3938);
and U5334 (N_5334,N_3693,N_3174);
nand U5335 (N_5335,N_3045,N_2036);
xor U5336 (N_5336,N_2997,N_2831);
or U5337 (N_5337,N_3470,N_3814);
xor U5338 (N_5338,N_3728,N_3039);
xnor U5339 (N_5339,N_2247,N_3061);
or U5340 (N_5340,N_2746,N_2123);
and U5341 (N_5341,N_2457,N_2797);
nand U5342 (N_5342,N_2180,N_3612);
nor U5343 (N_5343,N_2691,N_2158);
nand U5344 (N_5344,N_3807,N_2666);
nand U5345 (N_5345,N_3488,N_2310);
nor U5346 (N_5346,N_3465,N_2937);
and U5347 (N_5347,N_2108,N_3233);
nor U5348 (N_5348,N_2263,N_2140);
xnor U5349 (N_5349,N_2179,N_3233);
or U5350 (N_5350,N_3107,N_2022);
or U5351 (N_5351,N_3104,N_3541);
nand U5352 (N_5352,N_2392,N_2995);
xor U5353 (N_5353,N_3873,N_3631);
xor U5354 (N_5354,N_2191,N_2643);
or U5355 (N_5355,N_3212,N_3983);
nor U5356 (N_5356,N_2691,N_3448);
and U5357 (N_5357,N_2081,N_3103);
xnor U5358 (N_5358,N_2275,N_3535);
and U5359 (N_5359,N_2847,N_2498);
nand U5360 (N_5360,N_3476,N_2961);
and U5361 (N_5361,N_3389,N_3512);
nand U5362 (N_5362,N_3083,N_2448);
xnor U5363 (N_5363,N_2937,N_3601);
or U5364 (N_5364,N_3939,N_2071);
and U5365 (N_5365,N_2873,N_3604);
nand U5366 (N_5366,N_2625,N_2665);
nand U5367 (N_5367,N_3417,N_3643);
xor U5368 (N_5368,N_2345,N_2451);
and U5369 (N_5369,N_2587,N_2384);
and U5370 (N_5370,N_3008,N_2967);
or U5371 (N_5371,N_2377,N_3252);
nand U5372 (N_5372,N_2926,N_3214);
and U5373 (N_5373,N_3962,N_3552);
xnor U5374 (N_5374,N_2396,N_3416);
nand U5375 (N_5375,N_3351,N_2155);
xor U5376 (N_5376,N_2668,N_2864);
xnor U5377 (N_5377,N_2243,N_2115);
xnor U5378 (N_5378,N_3286,N_2601);
and U5379 (N_5379,N_3804,N_3888);
nor U5380 (N_5380,N_3289,N_3062);
and U5381 (N_5381,N_2709,N_3816);
xnor U5382 (N_5382,N_3528,N_2766);
xor U5383 (N_5383,N_2406,N_2850);
or U5384 (N_5384,N_2130,N_3163);
xnor U5385 (N_5385,N_2569,N_3137);
and U5386 (N_5386,N_3477,N_3049);
nor U5387 (N_5387,N_2021,N_2603);
nand U5388 (N_5388,N_3567,N_2956);
and U5389 (N_5389,N_3254,N_2146);
nor U5390 (N_5390,N_3688,N_2531);
or U5391 (N_5391,N_3689,N_3972);
xor U5392 (N_5392,N_3512,N_2137);
nand U5393 (N_5393,N_3629,N_3094);
and U5394 (N_5394,N_2837,N_2282);
xor U5395 (N_5395,N_2472,N_3810);
xnor U5396 (N_5396,N_2238,N_3323);
xnor U5397 (N_5397,N_2431,N_3948);
and U5398 (N_5398,N_2567,N_2708);
and U5399 (N_5399,N_2336,N_3264);
nand U5400 (N_5400,N_2160,N_3099);
or U5401 (N_5401,N_3419,N_3350);
xnor U5402 (N_5402,N_2550,N_2619);
nor U5403 (N_5403,N_2730,N_2900);
or U5404 (N_5404,N_2346,N_3916);
and U5405 (N_5405,N_2444,N_3971);
or U5406 (N_5406,N_3803,N_2991);
xnor U5407 (N_5407,N_2960,N_2745);
or U5408 (N_5408,N_2213,N_3101);
nor U5409 (N_5409,N_2507,N_2927);
xor U5410 (N_5410,N_3614,N_3288);
or U5411 (N_5411,N_2141,N_3619);
nand U5412 (N_5412,N_3431,N_3012);
or U5413 (N_5413,N_3446,N_2955);
xnor U5414 (N_5414,N_2241,N_2301);
xor U5415 (N_5415,N_3312,N_3395);
nor U5416 (N_5416,N_2682,N_2325);
nor U5417 (N_5417,N_2209,N_3588);
or U5418 (N_5418,N_2387,N_2462);
and U5419 (N_5419,N_3694,N_2759);
nand U5420 (N_5420,N_2301,N_3759);
nor U5421 (N_5421,N_3306,N_3471);
xor U5422 (N_5422,N_3765,N_2067);
and U5423 (N_5423,N_2634,N_2645);
or U5424 (N_5424,N_2013,N_3326);
nor U5425 (N_5425,N_2411,N_3502);
and U5426 (N_5426,N_3564,N_3484);
xor U5427 (N_5427,N_2936,N_2055);
or U5428 (N_5428,N_3194,N_3767);
nor U5429 (N_5429,N_3496,N_3828);
xnor U5430 (N_5430,N_2985,N_2231);
nand U5431 (N_5431,N_2021,N_2322);
nand U5432 (N_5432,N_3463,N_2727);
and U5433 (N_5433,N_2380,N_2420);
or U5434 (N_5434,N_2951,N_3158);
xnor U5435 (N_5435,N_2407,N_2002);
nor U5436 (N_5436,N_2898,N_3569);
xor U5437 (N_5437,N_2216,N_3789);
or U5438 (N_5438,N_3806,N_3866);
xnor U5439 (N_5439,N_3390,N_2681);
nand U5440 (N_5440,N_3806,N_3526);
and U5441 (N_5441,N_2173,N_3199);
xor U5442 (N_5442,N_2449,N_2323);
nor U5443 (N_5443,N_3654,N_3727);
nand U5444 (N_5444,N_2005,N_2633);
and U5445 (N_5445,N_3998,N_3872);
nand U5446 (N_5446,N_3715,N_2548);
nand U5447 (N_5447,N_2197,N_3856);
xnor U5448 (N_5448,N_2470,N_3186);
nor U5449 (N_5449,N_2264,N_2346);
or U5450 (N_5450,N_2167,N_2861);
and U5451 (N_5451,N_3975,N_2388);
nand U5452 (N_5452,N_3862,N_3560);
xor U5453 (N_5453,N_2232,N_2457);
nand U5454 (N_5454,N_3564,N_2560);
nor U5455 (N_5455,N_3251,N_2310);
nor U5456 (N_5456,N_3554,N_2083);
nor U5457 (N_5457,N_3634,N_3373);
and U5458 (N_5458,N_2617,N_3002);
and U5459 (N_5459,N_2605,N_3994);
nor U5460 (N_5460,N_2397,N_3159);
and U5461 (N_5461,N_3141,N_3806);
xor U5462 (N_5462,N_2599,N_2939);
xnor U5463 (N_5463,N_3832,N_3646);
or U5464 (N_5464,N_2876,N_2281);
or U5465 (N_5465,N_3252,N_2400);
or U5466 (N_5466,N_3185,N_2577);
and U5467 (N_5467,N_2411,N_3909);
nor U5468 (N_5468,N_3953,N_3216);
xnor U5469 (N_5469,N_2457,N_3850);
nor U5470 (N_5470,N_2575,N_3446);
nor U5471 (N_5471,N_3659,N_3329);
nand U5472 (N_5472,N_2074,N_3792);
nor U5473 (N_5473,N_2291,N_3762);
and U5474 (N_5474,N_2379,N_2872);
xor U5475 (N_5475,N_3581,N_2337);
and U5476 (N_5476,N_2383,N_3474);
nor U5477 (N_5477,N_2661,N_2330);
xnor U5478 (N_5478,N_3868,N_3802);
and U5479 (N_5479,N_2038,N_3321);
nand U5480 (N_5480,N_2085,N_3695);
or U5481 (N_5481,N_2836,N_3154);
nor U5482 (N_5482,N_3099,N_2684);
or U5483 (N_5483,N_2252,N_3636);
xnor U5484 (N_5484,N_3082,N_3036);
nor U5485 (N_5485,N_3006,N_3800);
or U5486 (N_5486,N_2599,N_3916);
and U5487 (N_5487,N_2969,N_3431);
or U5488 (N_5488,N_3736,N_3687);
xor U5489 (N_5489,N_2563,N_3440);
xnor U5490 (N_5490,N_3939,N_2437);
or U5491 (N_5491,N_3187,N_2920);
nand U5492 (N_5492,N_3339,N_3096);
nand U5493 (N_5493,N_2488,N_2788);
and U5494 (N_5494,N_3787,N_2841);
or U5495 (N_5495,N_2975,N_3982);
xor U5496 (N_5496,N_2235,N_3720);
nand U5497 (N_5497,N_2942,N_2731);
xor U5498 (N_5498,N_3651,N_3977);
nand U5499 (N_5499,N_3390,N_2302);
nor U5500 (N_5500,N_3194,N_3970);
or U5501 (N_5501,N_2994,N_3275);
or U5502 (N_5502,N_2840,N_3218);
or U5503 (N_5503,N_3370,N_2016);
nor U5504 (N_5504,N_3293,N_2607);
or U5505 (N_5505,N_2950,N_3685);
or U5506 (N_5506,N_2752,N_2052);
and U5507 (N_5507,N_3782,N_3857);
xor U5508 (N_5508,N_3218,N_3104);
and U5509 (N_5509,N_2613,N_3553);
nand U5510 (N_5510,N_3463,N_3868);
or U5511 (N_5511,N_3244,N_2469);
and U5512 (N_5512,N_3775,N_2821);
and U5513 (N_5513,N_3458,N_3843);
nor U5514 (N_5514,N_2810,N_3240);
xor U5515 (N_5515,N_2808,N_2467);
and U5516 (N_5516,N_3950,N_3454);
nand U5517 (N_5517,N_2443,N_2387);
and U5518 (N_5518,N_3095,N_2557);
nand U5519 (N_5519,N_2956,N_3194);
or U5520 (N_5520,N_2853,N_3362);
nor U5521 (N_5521,N_2201,N_3095);
and U5522 (N_5522,N_2507,N_2485);
or U5523 (N_5523,N_3897,N_3804);
xnor U5524 (N_5524,N_3389,N_3838);
xnor U5525 (N_5525,N_2355,N_3136);
and U5526 (N_5526,N_2459,N_2456);
and U5527 (N_5527,N_2628,N_2877);
and U5528 (N_5528,N_2553,N_3792);
xor U5529 (N_5529,N_2855,N_2822);
xor U5530 (N_5530,N_2480,N_3321);
or U5531 (N_5531,N_3254,N_3645);
xnor U5532 (N_5532,N_3031,N_3113);
nand U5533 (N_5533,N_3418,N_3277);
nor U5534 (N_5534,N_3260,N_3952);
or U5535 (N_5535,N_2276,N_2574);
xor U5536 (N_5536,N_2824,N_2236);
xnor U5537 (N_5537,N_2805,N_2752);
nor U5538 (N_5538,N_3348,N_3924);
nand U5539 (N_5539,N_3583,N_3214);
and U5540 (N_5540,N_2884,N_2457);
or U5541 (N_5541,N_2249,N_2292);
and U5542 (N_5542,N_2782,N_2064);
or U5543 (N_5543,N_2238,N_3137);
nor U5544 (N_5544,N_3019,N_2818);
and U5545 (N_5545,N_2975,N_2041);
xor U5546 (N_5546,N_2096,N_3266);
nor U5547 (N_5547,N_3606,N_2726);
or U5548 (N_5548,N_3465,N_3928);
or U5549 (N_5549,N_3213,N_3605);
xor U5550 (N_5550,N_2200,N_2081);
nor U5551 (N_5551,N_2824,N_3722);
xnor U5552 (N_5552,N_2962,N_3587);
nand U5553 (N_5553,N_3230,N_2078);
and U5554 (N_5554,N_3895,N_3227);
and U5555 (N_5555,N_2437,N_2623);
xnor U5556 (N_5556,N_2943,N_2299);
xor U5557 (N_5557,N_2819,N_2136);
xnor U5558 (N_5558,N_3769,N_2646);
and U5559 (N_5559,N_3726,N_3110);
and U5560 (N_5560,N_2531,N_2909);
nand U5561 (N_5561,N_2359,N_3329);
or U5562 (N_5562,N_3223,N_2921);
nand U5563 (N_5563,N_2940,N_2526);
xnor U5564 (N_5564,N_3845,N_2836);
nor U5565 (N_5565,N_3303,N_3083);
and U5566 (N_5566,N_2836,N_3266);
and U5567 (N_5567,N_3926,N_2052);
and U5568 (N_5568,N_3054,N_3483);
or U5569 (N_5569,N_3920,N_3404);
nor U5570 (N_5570,N_3101,N_2509);
nor U5571 (N_5571,N_3709,N_3548);
or U5572 (N_5572,N_2948,N_3580);
xor U5573 (N_5573,N_2002,N_3801);
nor U5574 (N_5574,N_3085,N_2815);
or U5575 (N_5575,N_2109,N_3261);
nand U5576 (N_5576,N_3234,N_2059);
nand U5577 (N_5577,N_2855,N_3968);
xnor U5578 (N_5578,N_2623,N_2525);
or U5579 (N_5579,N_3206,N_3918);
xor U5580 (N_5580,N_3155,N_2516);
or U5581 (N_5581,N_3553,N_2288);
or U5582 (N_5582,N_3705,N_3502);
xor U5583 (N_5583,N_2348,N_2281);
and U5584 (N_5584,N_3620,N_3429);
or U5585 (N_5585,N_3101,N_2872);
xor U5586 (N_5586,N_2970,N_2364);
and U5587 (N_5587,N_3665,N_2735);
nor U5588 (N_5588,N_2077,N_3415);
nor U5589 (N_5589,N_2190,N_3361);
xor U5590 (N_5590,N_2990,N_2095);
and U5591 (N_5591,N_2674,N_2026);
nor U5592 (N_5592,N_3924,N_2098);
nand U5593 (N_5593,N_3974,N_3114);
or U5594 (N_5594,N_2999,N_2595);
nand U5595 (N_5595,N_3555,N_3156);
nor U5596 (N_5596,N_2915,N_2388);
or U5597 (N_5597,N_2828,N_2583);
nor U5598 (N_5598,N_2030,N_2316);
and U5599 (N_5599,N_3637,N_2978);
nor U5600 (N_5600,N_2139,N_3236);
or U5601 (N_5601,N_3979,N_2545);
or U5602 (N_5602,N_3104,N_3076);
nand U5603 (N_5603,N_2451,N_2915);
nor U5604 (N_5604,N_3393,N_2865);
and U5605 (N_5605,N_3063,N_3862);
xnor U5606 (N_5606,N_2836,N_2107);
and U5607 (N_5607,N_2591,N_3794);
nor U5608 (N_5608,N_2860,N_3355);
nand U5609 (N_5609,N_2383,N_3491);
xor U5610 (N_5610,N_3549,N_3913);
nor U5611 (N_5611,N_2235,N_2056);
nor U5612 (N_5612,N_2540,N_2262);
nand U5613 (N_5613,N_2305,N_3736);
xor U5614 (N_5614,N_3801,N_3926);
and U5615 (N_5615,N_3520,N_3637);
nand U5616 (N_5616,N_2275,N_3581);
or U5617 (N_5617,N_2415,N_3647);
or U5618 (N_5618,N_2899,N_3326);
or U5619 (N_5619,N_3203,N_2615);
nand U5620 (N_5620,N_3833,N_2805);
xnor U5621 (N_5621,N_2790,N_3425);
nand U5622 (N_5622,N_3558,N_3329);
nor U5623 (N_5623,N_2748,N_2941);
nand U5624 (N_5624,N_3124,N_3137);
nor U5625 (N_5625,N_3301,N_3565);
or U5626 (N_5626,N_3199,N_3441);
nor U5627 (N_5627,N_3607,N_3231);
or U5628 (N_5628,N_3080,N_2984);
nor U5629 (N_5629,N_2444,N_2310);
nor U5630 (N_5630,N_2454,N_2866);
nor U5631 (N_5631,N_2053,N_3442);
nor U5632 (N_5632,N_3164,N_2128);
xnor U5633 (N_5633,N_3382,N_2078);
and U5634 (N_5634,N_3656,N_3025);
nor U5635 (N_5635,N_3415,N_3919);
or U5636 (N_5636,N_3081,N_3313);
nand U5637 (N_5637,N_2622,N_3550);
nor U5638 (N_5638,N_3111,N_3417);
nor U5639 (N_5639,N_2489,N_2734);
nor U5640 (N_5640,N_2406,N_3805);
and U5641 (N_5641,N_3430,N_2610);
nand U5642 (N_5642,N_2235,N_2796);
or U5643 (N_5643,N_3346,N_3152);
nand U5644 (N_5644,N_2891,N_3834);
and U5645 (N_5645,N_3808,N_3390);
nor U5646 (N_5646,N_2049,N_2332);
or U5647 (N_5647,N_3162,N_3002);
or U5648 (N_5648,N_2715,N_3868);
nand U5649 (N_5649,N_2375,N_3812);
and U5650 (N_5650,N_2530,N_2666);
or U5651 (N_5651,N_3186,N_3498);
and U5652 (N_5652,N_3699,N_2240);
nand U5653 (N_5653,N_3812,N_2619);
and U5654 (N_5654,N_3153,N_2580);
nor U5655 (N_5655,N_3497,N_3345);
and U5656 (N_5656,N_2955,N_2336);
and U5657 (N_5657,N_3569,N_2140);
or U5658 (N_5658,N_2133,N_3939);
or U5659 (N_5659,N_2553,N_2949);
and U5660 (N_5660,N_3005,N_2730);
and U5661 (N_5661,N_2911,N_3223);
and U5662 (N_5662,N_3085,N_3458);
and U5663 (N_5663,N_2455,N_2102);
or U5664 (N_5664,N_3914,N_3694);
or U5665 (N_5665,N_3315,N_3359);
or U5666 (N_5666,N_2887,N_3359);
xor U5667 (N_5667,N_3535,N_3704);
nand U5668 (N_5668,N_3906,N_3419);
nand U5669 (N_5669,N_2724,N_3411);
nor U5670 (N_5670,N_3787,N_3508);
xor U5671 (N_5671,N_3354,N_2939);
nor U5672 (N_5672,N_2856,N_3962);
nor U5673 (N_5673,N_3899,N_3388);
nor U5674 (N_5674,N_3974,N_3970);
and U5675 (N_5675,N_3651,N_3110);
nor U5676 (N_5676,N_2880,N_3956);
nor U5677 (N_5677,N_2790,N_2670);
nor U5678 (N_5678,N_3454,N_2130);
or U5679 (N_5679,N_3765,N_2375);
nor U5680 (N_5680,N_2183,N_2980);
and U5681 (N_5681,N_2087,N_3842);
nand U5682 (N_5682,N_2412,N_3912);
xnor U5683 (N_5683,N_2690,N_2180);
nand U5684 (N_5684,N_2400,N_2578);
xnor U5685 (N_5685,N_2362,N_2263);
nor U5686 (N_5686,N_3480,N_2665);
nor U5687 (N_5687,N_2844,N_3416);
and U5688 (N_5688,N_2709,N_2160);
xnor U5689 (N_5689,N_3970,N_3883);
and U5690 (N_5690,N_2098,N_3715);
nor U5691 (N_5691,N_2325,N_2400);
nand U5692 (N_5692,N_3939,N_3977);
nand U5693 (N_5693,N_3046,N_3721);
nor U5694 (N_5694,N_3514,N_3415);
and U5695 (N_5695,N_2915,N_2753);
nand U5696 (N_5696,N_3193,N_2308);
nand U5697 (N_5697,N_2077,N_3926);
or U5698 (N_5698,N_2652,N_2361);
or U5699 (N_5699,N_3275,N_3939);
nor U5700 (N_5700,N_2042,N_2529);
or U5701 (N_5701,N_3367,N_3817);
nand U5702 (N_5702,N_3063,N_3140);
and U5703 (N_5703,N_3474,N_2778);
nor U5704 (N_5704,N_3270,N_3003);
nor U5705 (N_5705,N_2075,N_2097);
xnor U5706 (N_5706,N_2684,N_3910);
nand U5707 (N_5707,N_2742,N_3497);
nor U5708 (N_5708,N_2251,N_2156);
or U5709 (N_5709,N_3484,N_3833);
nand U5710 (N_5710,N_3816,N_2097);
xnor U5711 (N_5711,N_3190,N_2098);
nand U5712 (N_5712,N_3930,N_3971);
or U5713 (N_5713,N_2553,N_3181);
nor U5714 (N_5714,N_2612,N_3671);
nand U5715 (N_5715,N_2479,N_3202);
nand U5716 (N_5716,N_3407,N_2352);
and U5717 (N_5717,N_3928,N_3395);
and U5718 (N_5718,N_2662,N_2273);
xnor U5719 (N_5719,N_2809,N_3959);
xor U5720 (N_5720,N_3759,N_2858);
nor U5721 (N_5721,N_3233,N_3663);
nor U5722 (N_5722,N_2805,N_2027);
nand U5723 (N_5723,N_3452,N_2844);
and U5724 (N_5724,N_2144,N_2216);
or U5725 (N_5725,N_3785,N_2091);
and U5726 (N_5726,N_3484,N_2963);
nand U5727 (N_5727,N_3129,N_2045);
nand U5728 (N_5728,N_3408,N_3677);
nand U5729 (N_5729,N_2220,N_2984);
nand U5730 (N_5730,N_2047,N_3943);
nand U5731 (N_5731,N_2911,N_2346);
xor U5732 (N_5732,N_3571,N_3851);
xor U5733 (N_5733,N_2269,N_3996);
xnor U5734 (N_5734,N_3017,N_2434);
nand U5735 (N_5735,N_2068,N_3241);
nor U5736 (N_5736,N_2312,N_3979);
and U5737 (N_5737,N_3851,N_3176);
and U5738 (N_5738,N_2138,N_2224);
nor U5739 (N_5739,N_2564,N_3321);
xnor U5740 (N_5740,N_3595,N_3319);
nor U5741 (N_5741,N_3195,N_2748);
nand U5742 (N_5742,N_3157,N_3535);
xor U5743 (N_5743,N_3443,N_2086);
or U5744 (N_5744,N_3575,N_3420);
and U5745 (N_5745,N_3012,N_3318);
nor U5746 (N_5746,N_3302,N_3087);
and U5747 (N_5747,N_3184,N_2019);
or U5748 (N_5748,N_3178,N_3173);
xnor U5749 (N_5749,N_3410,N_2206);
and U5750 (N_5750,N_3011,N_3170);
or U5751 (N_5751,N_2929,N_3840);
nor U5752 (N_5752,N_3124,N_3946);
nand U5753 (N_5753,N_3999,N_2439);
nand U5754 (N_5754,N_2702,N_3192);
or U5755 (N_5755,N_2369,N_3385);
or U5756 (N_5756,N_3218,N_3912);
nor U5757 (N_5757,N_2090,N_2623);
or U5758 (N_5758,N_2728,N_3327);
xor U5759 (N_5759,N_2881,N_3687);
nor U5760 (N_5760,N_2830,N_3578);
nand U5761 (N_5761,N_2233,N_3895);
xor U5762 (N_5762,N_3082,N_2966);
nand U5763 (N_5763,N_2788,N_3331);
xnor U5764 (N_5764,N_2719,N_2812);
nor U5765 (N_5765,N_3103,N_2702);
xor U5766 (N_5766,N_2858,N_3215);
xor U5767 (N_5767,N_3724,N_2891);
xor U5768 (N_5768,N_3641,N_3407);
nor U5769 (N_5769,N_2697,N_2049);
or U5770 (N_5770,N_3439,N_2286);
nand U5771 (N_5771,N_3287,N_2467);
xnor U5772 (N_5772,N_2782,N_2488);
or U5773 (N_5773,N_2479,N_2939);
xnor U5774 (N_5774,N_2647,N_2048);
nor U5775 (N_5775,N_2332,N_3893);
or U5776 (N_5776,N_2406,N_2305);
or U5777 (N_5777,N_2625,N_3966);
nand U5778 (N_5778,N_3901,N_2508);
xor U5779 (N_5779,N_3215,N_2533);
xor U5780 (N_5780,N_3967,N_3327);
or U5781 (N_5781,N_3876,N_3234);
xnor U5782 (N_5782,N_2628,N_2239);
xor U5783 (N_5783,N_2848,N_2847);
xor U5784 (N_5784,N_3882,N_3586);
or U5785 (N_5785,N_3650,N_3675);
xnor U5786 (N_5786,N_3542,N_3631);
or U5787 (N_5787,N_2872,N_2646);
or U5788 (N_5788,N_3405,N_2769);
and U5789 (N_5789,N_2530,N_2600);
xnor U5790 (N_5790,N_3156,N_2816);
xor U5791 (N_5791,N_3389,N_2142);
and U5792 (N_5792,N_3313,N_2881);
nand U5793 (N_5793,N_2801,N_2594);
xor U5794 (N_5794,N_2431,N_3022);
xnor U5795 (N_5795,N_3926,N_3294);
xor U5796 (N_5796,N_2890,N_3786);
or U5797 (N_5797,N_3818,N_2612);
and U5798 (N_5798,N_3241,N_3269);
nand U5799 (N_5799,N_2892,N_2373);
nor U5800 (N_5800,N_3269,N_3866);
nand U5801 (N_5801,N_3832,N_2580);
nand U5802 (N_5802,N_2466,N_3515);
nor U5803 (N_5803,N_3718,N_3543);
nand U5804 (N_5804,N_3725,N_3045);
nor U5805 (N_5805,N_2270,N_3346);
or U5806 (N_5806,N_2090,N_2968);
xor U5807 (N_5807,N_3375,N_3746);
or U5808 (N_5808,N_3733,N_3079);
or U5809 (N_5809,N_3018,N_3039);
and U5810 (N_5810,N_2644,N_2621);
and U5811 (N_5811,N_2158,N_3172);
xor U5812 (N_5812,N_2952,N_2953);
xor U5813 (N_5813,N_3096,N_2700);
nor U5814 (N_5814,N_2351,N_3897);
xor U5815 (N_5815,N_3774,N_2579);
and U5816 (N_5816,N_2582,N_2011);
and U5817 (N_5817,N_2692,N_3786);
and U5818 (N_5818,N_3937,N_2050);
and U5819 (N_5819,N_2085,N_3831);
xnor U5820 (N_5820,N_2764,N_3110);
xor U5821 (N_5821,N_3924,N_3602);
nor U5822 (N_5822,N_3458,N_3307);
xnor U5823 (N_5823,N_2813,N_3748);
xor U5824 (N_5824,N_2398,N_2313);
or U5825 (N_5825,N_3462,N_3543);
nor U5826 (N_5826,N_3331,N_2672);
or U5827 (N_5827,N_2056,N_3891);
xor U5828 (N_5828,N_3903,N_2504);
xor U5829 (N_5829,N_2930,N_2061);
nand U5830 (N_5830,N_2773,N_3529);
xnor U5831 (N_5831,N_3737,N_2210);
nor U5832 (N_5832,N_2079,N_2576);
nor U5833 (N_5833,N_2092,N_3334);
and U5834 (N_5834,N_2512,N_3400);
xnor U5835 (N_5835,N_2283,N_2185);
nand U5836 (N_5836,N_3552,N_2930);
xnor U5837 (N_5837,N_2512,N_2368);
or U5838 (N_5838,N_2763,N_2182);
nand U5839 (N_5839,N_2392,N_2399);
and U5840 (N_5840,N_3506,N_2938);
or U5841 (N_5841,N_3549,N_2553);
or U5842 (N_5842,N_3026,N_2891);
nand U5843 (N_5843,N_2758,N_3020);
nor U5844 (N_5844,N_3100,N_2552);
xnor U5845 (N_5845,N_3234,N_2742);
nor U5846 (N_5846,N_2090,N_3259);
and U5847 (N_5847,N_3017,N_2145);
and U5848 (N_5848,N_3612,N_3121);
nor U5849 (N_5849,N_3141,N_2755);
nor U5850 (N_5850,N_3797,N_3626);
or U5851 (N_5851,N_2504,N_2676);
or U5852 (N_5852,N_2532,N_2057);
xnor U5853 (N_5853,N_3813,N_3175);
or U5854 (N_5854,N_2086,N_2093);
nand U5855 (N_5855,N_3286,N_2498);
xor U5856 (N_5856,N_2128,N_3055);
nand U5857 (N_5857,N_2401,N_3833);
and U5858 (N_5858,N_3476,N_3448);
and U5859 (N_5859,N_2418,N_2726);
or U5860 (N_5860,N_2227,N_2530);
nor U5861 (N_5861,N_3269,N_2095);
nand U5862 (N_5862,N_3407,N_3151);
and U5863 (N_5863,N_3011,N_2918);
nor U5864 (N_5864,N_2784,N_2617);
xnor U5865 (N_5865,N_3118,N_3730);
and U5866 (N_5866,N_3184,N_3456);
and U5867 (N_5867,N_2017,N_2470);
nand U5868 (N_5868,N_2643,N_3002);
nor U5869 (N_5869,N_3691,N_2018);
xor U5870 (N_5870,N_3889,N_3247);
xor U5871 (N_5871,N_3935,N_3409);
and U5872 (N_5872,N_2929,N_2682);
nor U5873 (N_5873,N_2274,N_3438);
xnor U5874 (N_5874,N_2644,N_3185);
xnor U5875 (N_5875,N_3550,N_3780);
and U5876 (N_5876,N_3502,N_2646);
nand U5877 (N_5877,N_2865,N_2751);
or U5878 (N_5878,N_3612,N_3011);
nor U5879 (N_5879,N_3236,N_3516);
or U5880 (N_5880,N_2808,N_2079);
nor U5881 (N_5881,N_3775,N_3803);
and U5882 (N_5882,N_3712,N_2539);
nand U5883 (N_5883,N_2033,N_3405);
nor U5884 (N_5884,N_3764,N_3938);
or U5885 (N_5885,N_3456,N_3350);
nand U5886 (N_5886,N_3105,N_2010);
or U5887 (N_5887,N_3341,N_2739);
nor U5888 (N_5888,N_3472,N_2214);
nor U5889 (N_5889,N_3400,N_3347);
or U5890 (N_5890,N_3782,N_3230);
or U5891 (N_5891,N_2184,N_3023);
and U5892 (N_5892,N_3402,N_2280);
xnor U5893 (N_5893,N_3917,N_2199);
xor U5894 (N_5894,N_2388,N_3856);
nor U5895 (N_5895,N_3094,N_2395);
and U5896 (N_5896,N_3799,N_3691);
nor U5897 (N_5897,N_2676,N_2546);
nor U5898 (N_5898,N_2931,N_2802);
xor U5899 (N_5899,N_2880,N_2891);
nor U5900 (N_5900,N_2067,N_3428);
xnor U5901 (N_5901,N_3681,N_3053);
and U5902 (N_5902,N_3029,N_2166);
or U5903 (N_5903,N_3464,N_3123);
and U5904 (N_5904,N_2182,N_2759);
xor U5905 (N_5905,N_2828,N_2822);
xor U5906 (N_5906,N_3096,N_2776);
or U5907 (N_5907,N_3036,N_3050);
nor U5908 (N_5908,N_2466,N_2214);
xnor U5909 (N_5909,N_3424,N_2735);
or U5910 (N_5910,N_2011,N_3056);
or U5911 (N_5911,N_2441,N_2009);
nor U5912 (N_5912,N_2369,N_2651);
or U5913 (N_5913,N_2274,N_3443);
or U5914 (N_5914,N_3246,N_3278);
nor U5915 (N_5915,N_2178,N_3989);
or U5916 (N_5916,N_3259,N_3884);
and U5917 (N_5917,N_2654,N_3702);
nor U5918 (N_5918,N_2429,N_2115);
nor U5919 (N_5919,N_3396,N_2164);
nand U5920 (N_5920,N_2362,N_2921);
nor U5921 (N_5921,N_3026,N_2573);
nand U5922 (N_5922,N_3609,N_2297);
nor U5923 (N_5923,N_3245,N_3539);
or U5924 (N_5924,N_2072,N_2234);
nor U5925 (N_5925,N_2809,N_2583);
nand U5926 (N_5926,N_3113,N_3956);
nand U5927 (N_5927,N_2093,N_2124);
and U5928 (N_5928,N_3467,N_3076);
and U5929 (N_5929,N_2421,N_3872);
and U5930 (N_5930,N_3970,N_3624);
and U5931 (N_5931,N_3988,N_3664);
nor U5932 (N_5932,N_2245,N_3889);
and U5933 (N_5933,N_3165,N_2584);
or U5934 (N_5934,N_2433,N_2602);
nand U5935 (N_5935,N_3092,N_2098);
nor U5936 (N_5936,N_2584,N_2349);
xor U5937 (N_5937,N_3327,N_2808);
and U5938 (N_5938,N_3904,N_3838);
and U5939 (N_5939,N_3180,N_3364);
xor U5940 (N_5940,N_2344,N_2068);
or U5941 (N_5941,N_2420,N_2688);
xor U5942 (N_5942,N_3036,N_2796);
and U5943 (N_5943,N_2079,N_3598);
xnor U5944 (N_5944,N_2253,N_2034);
and U5945 (N_5945,N_3378,N_2614);
xnor U5946 (N_5946,N_2595,N_3494);
and U5947 (N_5947,N_2796,N_3873);
or U5948 (N_5948,N_2085,N_2922);
xnor U5949 (N_5949,N_2267,N_2975);
and U5950 (N_5950,N_3462,N_2489);
nand U5951 (N_5951,N_2339,N_3214);
or U5952 (N_5952,N_3708,N_3556);
and U5953 (N_5953,N_2714,N_3575);
or U5954 (N_5954,N_3084,N_2481);
or U5955 (N_5955,N_3789,N_3517);
and U5956 (N_5956,N_2589,N_2677);
xor U5957 (N_5957,N_3109,N_2758);
nand U5958 (N_5958,N_3472,N_3357);
xor U5959 (N_5959,N_3502,N_2034);
or U5960 (N_5960,N_3263,N_2763);
xor U5961 (N_5961,N_3570,N_2476);
nor U5962 (N_5962,N_2718,N_2582);
or U5963 (N_5963,N_2597,N_2142);
nand U5964 (N_5964,N_3772,N_2601);
or U5965 (N_5965,N_2337,N_3669);
nand U5966 (N_5966,N_3862,N_3021);
and U5967 (N_5967,N_3996,N_2789);
or U5968 (N_5968,N_3634,N_2704);
nand U5969 (N_5969,N_3534,N_3243);
or U5970 (N_5970,N_3774,N_3782);
and U5971 (N_5971,N_3504,N_3831);
nand U5972 (N_5972,N_3492,N_3374);
xnor U5973 (N_5973,N_3872,N_2861);
nor U5974 (N_5974,N_2533,N_3838);
xor U5975 (N_5975,N_3476,N_2275);
nand U5976 (N_5976,N_3163,N_3875);
or U5977 (N_5977,N_3437,N_2685);
and U5978 (N_5978,N_2352,N_3308);
nand U5979 (N_5979,N_2578,N_2901);
nand U5980 (N_5980,N_3468,N_3868);
or U5981 (N_5981,N_3869,N_3450);
xor U5982 (N_5982,N_2382,N_3759);
xnor U5983 (N_5983,N_3938,N_2294);
xor U5984 (N_5984,N_2088,N_2673);
or U5985 (N_5985,N_2831,N_2317);
xor U5986 (N_5986,N_3691,N_2305);
nor U5987 (N_5987,N_2365,N_2966);
nor U5988 (N_5988,N_3559,N_3356);
nor U5989 (N_5989,N_3808,N_2782);
and U5990 (N_5990,N_2985,N_2646);
and U5991 (N_5991,N_2607,N_3100);
nor U5992 (N_5992,N_2899,N_2491);
or U5993 (N_5993,N_2577,N_2656);
or U5994 (N_5994,N_3739,N_2896);
nor U5995 (N_5995,N_2305,N_2528);
xor U5996 (N_5996,N_2318,N_3788);
or U5997 (N_5997,N_2817,N_2235);
nand U5998 (N_5998,N_2388,N_3499);
or U5999 (N_5999,N_2853,N_2817);
nand U6000 (N_6000,N_5224,N_4926);
nand U6001 (N_6001,N_5170,N_4592);
and U6002 (N_6002,N_5151,N_4953);
nor U6003 (N_6003,N_5734,N_5988);
nand U6004 (N_6004,N_5472,N_5764);
and U6005 (N_6005,N_5861,N_5521);
nand U6006 (N_6006,N_4754,N_5994);
and U6007 (N_6007,N_5034,N_5272);
and U6008 (N_6008,N_5337,N_5308);
nor U6009 (N_6009,N_4134,N_4076);
xnor U6010 (N_6010,N_5517,N_4129);
nand U6011 (N_6011,N_4061,N_4752);
and U6012 (N_6012,N_4983,N_4646);
nand U6013 (N_6013,N_5913,N_4197);
and U6014 (N_6014,N_4885,N_5992);
nor U6015 (N_6015,N_5356,N_5283);
xor U6016 (N_6016,N_5171,N_4711);
xor U6017 (N_6017,N_4620,N_4349);
or U6018 (N_6018,N_5225,N_5306);
nand U6019 (N_6019,N_5690,N_4180);
and U6020 (N_6020,N_4111,N_4788);
nor U6021 (N_6021,N_4471,N_4192);
xor U6022 (N_6022,N_4294,N_4618);
xnor U6023 (N_6023,N_4528,N_5282);
xnor U6024 (N_6024,N_4890,N_5009);
nor U6025 (N_6025,N_4574,N_5093);
xor U6026 (N_6026,N_4847,N_5546);
or U6027 (N_6027,N_4687,N_4059);
nor U6028 (N_6028,N_4946,N_5178);
nand U6029 (N_6029,N_4948,N_4087);
and U6030 (N_6030,N_4548,N_5120);
nor U6031 (N_6031,N_5500,N_5079);
nor U6032 (N_6032,N_5629,N_4727);
nand U6033 (N_6033,N_4625,N_5563);
xor U6034 (N_6034,N_5700,N_5425);
nand U6035 (N_6035,N_4793,N_4515);
xor U6036 (N_6036,N_5073,N_5376);
xor U6037 (N_6037,N_5245,N_4052);
nor U6038 (N_6038,N_5976,N_4122);
nor U6039 (N_6039,N_4614,N_4530);
and U6040 (N_6040,N_4317,N_5227);
nand U6041 (N_6041,N_5100,N_4585);
or U6042 (N_6042,N_5172,N_5681);
nor U6043 (N_6043,N_5366,N_4347);
xnor U6044 (N_6044,N_4132,N_4633);
and U6045 (N_6045,N_4673,N_5303);
and U6046 (N_6046,N_5555,N_4594);
or U6047 (N_6047,N_5378,N_5380);
or U6048 (N_6048,N_4274,N_5648);
or U6049 (N_6049,N_4504,N_4249);
and U6050 (N_6050,N_5561,N_4207);
and U6051 (N_6051,N_5132,N_5979);
nor U6052 (N_6052,N_5409,N_4360);
xor U6053 (N_6053,N_4522,N_4162);
and U6054 (N_6054,N_5639,N_4854);
and U6055 (N_6055,N_4586,N_5018);
and U6056 (N_6056,N_4467,N_4893);
or U6057 (N_6057,N_4193,N_5578);
nor U6058 (N_6058,N_5169,N_4863);
xnor U6059 (N_6059,N_4083,N_5019);
and U6060 (N_6060,N_4370,N_4767);
and U6061 (N_6061,N_4628,N_5857);
xnor U6062 (N_6062,N_5343,N_4278);
xnor U6063 (N_6063,N_5611,N_5523);
or U6064 (N_6064,N_4359,N_4035);
nand U6065 (N_6065,N_5756,N_5942);
or U6066 (N_6066,N_5781,N_5697);
xor U6067 (N_6067,N_5130,N_5256);
or U6068 (N_6068,N_5070,N_5569);
or U6069 (N_6069,N_5559,N_5807);
and U6070 (N_6070,N_5589,N_5035);
and U6071 (N_6071,N_4100,N_4679);
nand U6072 (N_6072,N_5436,N_5874);
xor U6073 (N_6073,N_5665,N_5250);
or U6074 (N_6074,N_5491,N_5760);
nand U6075 (N_6075,N_4588,N_5951);
or U6076 (N_6076,N_5742,N_5310);
nor U6077 (N_6077,N_5688,N_5428);
and U6078 (N_6078,N_5444,N_4627);
and U6079 (N_6079,N_4017,N_4984);
or U6080 (N_6080,N_5083,N_5934);
and U6081 (N_6081,N_5165,N_5751);
nand U6082 (N_6082,N_4730,N_4447);
nand U6083 (N_6083,N_4230,N_5887);
and U6084 (N_6084,N_5591,N_4326);
or U6085 (N_6085,N_5632,N_5512);
nor U6086 (N_6086,N_4365,N_5847);
nand U6087 (N_6087,N_5908,N_4526);
nand U6088 (N_6088,N_5138,N_4538);
and U6089 (N_6089,N_5363,N_4523);
nor U6090 (N_6090,N_5104,N_5040);
nand U6091 (N_6091,N_4891,N_4841);
xor U6092 (N_6092,N_5164,N_5274);
xor U6093 (N_6093,N_4986,N_4477);
or U6094 (N_6094,N_4080,N_4816);
nor U6095 (N_6095,N_5078,N_4099);
or U6096 (N_6096,N_5982,N_5362);
nand U6097 (N_6097,N_4559,N_4459);
and U6098 (N_6098,N_5647,N_5652);
or U6099 (N_6099,N_5486,N_5936);
nand U6100 (N_6100,N_5800,N_5066);
xnor U6101 (N_6101,N_5947,N_5309);
nor U6102 (N_6102,N_5268,N_4533);
xor U6103 (N_6103,N_5438,N_4838);
nand U6104 (N_6104,N_4290,N_4541);
or U6105 (N_6105,N_5174,N_4135);
and U6106 (N_6106,N_5177,N_5323);
xnor U6107 (N_6107,N_4635,N_5060);
xor U6108 (N_6108,N_4454,N_4884);
or U6109 (N_6109,N_5430,N_5207);
or U6110 (N_6110,N_4048,N_5048);
nor U6111 (N_6111,N_5968,N_5685);
nor U6112 (N_6112,N_4764,N_4051);
and U6113 (N_6113,N_4988,N_5014);
xor U6114 (N_6114,N_4581,N_4424);
and U6115 (N_6115,N_5289,N_4713);
or U6116 (N_6116,N_5889,N_4092);
nand U6117 (N_6117,N_4785,N_5106);
xor U6118 (N_6118,N_4272,N_5655);
nand U6119 (N_6119,N_5116,N_5520);
nor U6120 (N_6120,N_4259,N_5718);
nor U6121 (N_6121,N_5211,N_5941);
nor U6122 (N_6122,N_5881,N_5995);
nor U6123 (N_6123,N_4783,N_4546);
and U6124 (N_6124,N_5320,N_5198);
nor U6125 (N_6125,N_4794,N_4502);
xor U6126 (N_6126,N_4695,N_4248);
nand U6127 (N_6127,N_5352,N_5898);
xor U6128 (N_6128,N_4046,N_5902);
nor U6129 (N_6129,N_4503,N_4329);
xor U6130 (N_6130,N_5286,N_4762);
nor U6131 (N_6131,N_4246,N_5999);
nand U6132 (N_6132,N_4934,N_4185);
or U6133 (N_6133,N_5474,N_4427);
xor U6134 (N_6134,N_4166,N_4094);
or U6135 (N_6135,N_4889,N_5641);
xnor U6136 (N_6136,N_4066,N_4742);
nor U6137 (N_6137,N_4282,N_5181);
xnor U6138 (N_6138,N_4821,N_5131);
xor U6139 (N_6139,N_4340,N_5686);
and U6140 (N_6140,N_5072,N_5601);
nor U6141 (N_6141,N_4787,N_4173);
nor U6142 (N_6142,N_5209,N_5386);
nor U6143 (N_6143,N_4880,N_5485);
nand U6144 (N_6144,N_4848,N_5566);
xor U6145 (N_6145,N_5402,N_5571);
and U6146 (N_6146,N_4489,N_5406);
or U6147 (N_6147,N_4072,N_4086);
or U6148 (N_6148,N_4604,N_4426);
and U6149 (N_6149,N_5370,N_4989);
and U6150 (N_6150,N_4431,N_4461);
xnor U6151 (N_6151,N_5248,N_4577);
or U6152 (N_6152,N_4733,N_4853);
or U6153 (N_6153,N_5424,N_5064);
xor U6154 (N_6154,N_4911,N_5891);
and U6155 (N_6155,N_5417,N_5471);
xor U6156 (N_6156,N_5298,N_4795);
nand U6157 (N_6157,N_4043,N_4399);
or U6158 (N_6158,N_5126,N_5596);
nor U6159 (N_6159,N_4844,N_5278);
xnor U6160 (N_6160,N_5636,N_5670);
xnor U6161 (N_6161,N_4898,N_5918);
or U6162 (N_6162,N_4961,N_4070);
or U6163 (N_6163,N_5879,N_4299);
xor U6164 (N_6164,N_4959,N_4482);
nor U6165 (N_6165,N_5249,N_5706);
nand U6166 (N_6166,N_4830,N_5550);
xor U6167 (N_6167,N_5920,N_4746);
or U6168 (N_6168,N_4735,N_5324);
xor U6169 (N_6169,N_4544,N_5008);
nand U6170 (N_6170,N_5186,N_5082);
or U6171 (N_6171,N_4462,N_5032);
nand U6172 (N_6172,N_5345,N_5762);
nor U6173 (N_6173,N_5938,N_4313);
or U6174 (N_6174,N_4136,N_4700);
or U6175 (N_6175,N_5000,N_5831);
and U6176 (N_6176,N_5455,N_4979);
nor U6177 (N_6177,N_4393,N_5179);
nand U6178 (N_6178,N_4254,N_4146);
nand U6179 (N_6179,N_5206,N_5716);
or U6180 (N_6180,N_5758,N_4680);
or U6181 (N_6181,N_4743,N_4466);
nand U6182 (N_6182,N_5990,N_4808);
nand U6183 (N_6183,N_4545,N_5434);
nor U6184 (N_6184,N_5903,N_4827);
xnor U6185 (N_6185,N_4725,N_4167);
xor U6186 (N_6186,N_4148,N_5619);
xor U6187 (N_6187,N_4659,N_4600);
or U6188 (N_6188,N_4053,N_5787);
nand U6189 (N_6189,N_4772,N_5835);
and U6190 (N_6190,N_4138,N_4202);
or U6191 (N_6191,N_4837,N_4915);
nor U6192 (N_6192,N_4689,N_4539);
xnor U6193 (N_6193,N_4018,N_4974);
xor U6194 (N_6194,N_5433,N_4457);
and U6195 (N_6195,N_4331,N_4151);
nand U6196 (N_6196,N_5342,N_4871);
nor U6197 (N_6197,N_5400,N_4599);
nor U6198 (N_6198,N_4243,N_4570);
xor U6199 (N_6199,N_5574,N_4463);
and U6200 (N_6200,N_5545,N_5334);
xor U6201 (N_6201,N_5193,N_5943);
nor U6202 (N_6202,N_5316,N_4987);
nand U6203 (N_6203,N_4832,N_4710);
xor U6204 (N_6204,N_4267,N_4361);
or U6205 (N_6205,N_4064,N_5958);
or U6206 (N_6206,N_4745,N_4718);
or U6207 (N_6207,N_4114,N_5691);
nand U6208 (N_6208,N_4240,N_4956);
nand U6209 (N_6209,N_4496,N_5849);
nand U6210 (N_6210,N_5058,N_4560);
nand U6211 (N_6211,N_5625,N_4874);
nor U6212 (N_6212,N_5220,N_4971);
and U6213 (N_6213,N_4211,N_4917);
nor U6214 (N_6214,N_4210,N_5896);
and U6215 (N_6215,N_5488,N_5144);
or U6216 (N_6216,N_5226,N_4736);
xor U6217 (N_6217,N_5039,N_5701);
nand U6218 (N_6218,N_5877,N_5161);
nor U6219 (N_6219,N_4131,N_5530);
or U6220 (N_6220,N_5664,N_5257);
nor U6221 (N_6221,N_4065,N_4766);
and U6222 (N_6222,N_5931,N_4856);
xnor U6223 (N_6223,N_5797,N_4509);
nor U6224 (N_6224,N_4034,N_4943);
nor U6225 (N_6225,N_5522,N_5833);
nor U6226 (N_6226,N_5071,N_4201);
or U6227 (N_6227,N_5470,N_5870);
or U6228 (N_6228,N_5201,N_5585);
and U6229 (N_6229,N_5642,N_4090);
xnor U6230 (N_6230,N_4749,N_5203);
xnor U6231 (N_6231,N_5484,N_4801);
or U6232 (N_6232,N_4962,N_4147);
nand U6233 (N_6233,N_4784,N_4612);
nor U6234 (N_6234,N_5459,N_5302);
nor U6235 (N_6235,N_5348,N_5987);
nand U6236 (N_6236,N_5736,N_4098);
xnor U6237 (N_6237,N_5408,N_5615);
and U6238 (N_6238,N_5675,N_4770);
xor U6239 (N_6239,N_5969,N_5448);
nand U6240 (N_6240,N_5502,N_4261);
and U6241 (N_6241,N_4579,N_5710);
nand U6242 (N_6242,N_5937,N_5923);
nor U6243 (N_6243,N_5817,N_4158);
nor U6244 (N_6244,N_5330,N_4660);
xnor U6245 (N_6245,N_5962,N_4557);
or U6246 (N_6246,N_5163,N_5692);
nand U6247 (N_6247,N_5011,N_5509);
and U6248 (N_6248,N_4615,N_4605);
and U6249 (N_6249,N_4408,N_5059);
or U6250 (N_6250,N_4938,N_4106);
xnor U6251 (N_6251,N_5017,N_5483);
nand U6252 (N_6252,N_5614,N_4378);
xnor U6253 (N_6253,N_5075,N_5173);
or U6254 (N_6254,N_4460,N_4178);
nand U6255 (N_6255,N_4023,N_5441);
nor U6256 (N_6256,N_5863,N_4441);
xnor U6257 (N_6257,N_4491,N_5532);
and U6258 (N_6258,N_5111,N_5998);
nor U6259 (N_6259,N_4685,N_5640);
and U6260 (N_6260,N_5432,N_4701);
xor U6261 (N_6261,N_4144,N_4007);
and U6262 (N_6262,N_5883,N_4719);
and U6263 (N_6263,N_4343,N_5635);
and U6264 (N_6264,N_5195,N_4858);
and U6265 (N_6265,N_4047,N_5314);
xor U6266 (N_6266,N_5004,N_5809);
nor U6267 (N_6267,N_5341,N_4364);
nand U6268 (N_6268,N_5236,N_5057);
or U6269 (N_6269,N_5524,N_5715);
xnor U6270 (N_6270,N_4593,N_5020);
or U6271 (N_6271,N_4237,N_5077);
nand U6272 (N_6272,N_5346,N_4634);
and U6273 (N_6273,N_4597,N_4564);
and U6274 (N_6274,N_4995,N_4648);
and U6275 (N_6275,N_4927,N_5973);
xnor U6276 (N_6276,N_4892,N_5145);
nor U6277 (N_6277,N_5010,N_5733);
nor U6278 (N_6278,N_4654,N_5213);
and U6279 (N_6279,N_5147,N_5215);
or U6280 (N_6280,N_4667,N_4997);
and U6281 (N_6281,N_4169,N_5231);
or U6282 (N_6282,N_5354,N_5677);
nor U6283 (N_6283,N_4109,N_4354);
and U6284 (N_6284,N_4002,N_5719);
and U6285 (N_6285,N_5347,N_4110);
xor U6286 (N_6286,N_4866,N_4949);
or U6287 (N_6287,N_4705,N_5822);
nand U6288 (N_6288,N_4170,N_5105);
or U6289 (N_6289,N_4453,N_5288);
or U6290 (N_6290,N_5767,N_5492);
nand U6291 (N_6291,N_5910,N_5730);
nor U6292 (N_6292,N_5469,N_4403);
and U6293 (N_6293,N_5068,N_5924);
and U6294 (N_6294,N_4951,N_4717);
nand U6295 (N_6295,N_5155,N_4336);
and U6296 (N_6296,N_5698,N_5241);
xnor U6297 (N_6297,N_4493,N_4873);
nand U6298 (N_6298,N_4311,N_4353);
and U6299 (N_6299,N_5960,N_4590);
nand U6300 (N_6300,N_5727,N_5006);
and U6301 (N_6301,N_5813,N_4218);
nor U6302 (N_6302,N_4554,N_4476);
xor U6303 (N_6303,N_4498,N_4096);
xnor U6304 (N_6304,N_5600,N_5593);
nand U6305 (N_6305,N_4262,N_4511);
nor U6306 (N_6306,N_4985,N_5752);
or U6307 (N_6307,N_4865,N_4639);
or U6308 (N_6308,N_5875,N_4181);
nand U6309 (N_6309,N_5553,N_4228);
nand U6310 (N_6310,N_5127,N_4905);
nand U6311 (N_6311,N_4914,N_4081);
nor U6312 (N_6312,N_5694,N_4174);
nor U6313 (N_6313,N_5185,N_4287);
nor U6314 (N_6314,N_5045,N_4608);
nor U6315 (N_6315,N_4978,N_5737);
nand U6316 (N_6316,N_5832,N_5894);
nor U6317 (N_6317,N_4271,N_4696);
xor U6318 (N_6318,N_5305,N_4671);
nor U6319 (N_6319,N_5510,N_5328);
nor U6320 (N_6320,N_5156,N_5012);
xnor U6321 (N_6321,N_4652,N_4839);
nand U6322 (N_6322,N_4270,N_5930);
nand U6323 (N_6323,N_4789,N_4748);
or U6324 (N_6324,N_5412,N_4950);
xnor U6325 (N_6325,N_4179,N_4622);
xor U6326 (N_6326,N_4238,N_4833);
or U6327 (N_6327,N_5294,N_5663);
nor U6328 (N_6328,N_4478,N_4305);
and U6329 (N_6329,N_4401,N_4525);
and U6330 (N_6330,N_4485,N_4776);
nand U6331 (N_6331,N_4994,N_4348);
and U6332 (N_6332,N_4298,N_5056);
nor U6333 (N_6333,N_4391,N_5549);
or U6334 (N_6334,N_5872,N_5651);
or U6335 (N_6335,N_4596,N_4413);
nor U6336 (N_6336,N_5128,N_5047);
or U6337 (N_6337,N_4796,N_4536);
or U6338 (N_6338,N_4519,N_4714);
or U6339 (N_6339,N_4216,N_5229);
nand U6340 (N_6340,N_4647,N_4128);
or U6341 (N_6341,N_5753,N_5616);
xnor U6342 (N_6342,N_5714,N_4058);
or U6343 (N_6343,N_5580,N_4448);
xor U6344 (N_6344,N_5955,N_5301);
and U6345 (N_6345,N_5650,N_4433);
xnor U6346 (N_6346,N_5594,N_4321);
nand U6347 (N_6347,N_4982,N_4966);
nor U6348 (N_6348,N_5827,N_4550);
nand U6349 (N_6349,N_4507,N_4933);
xnor U6350 (N_6350,N_4606,N_5188);
nand U6351 (N_6351,N_5728,N_4993);
or U6352 (N_6352,N_5263,N_4610);
nor U6353 (N_6353,N_4814,N_4356);
nand U6354 (N_6354,N_5493,N_4418);
xor U6355 (N_6355,N_5199,N_4888);
and U6356 (N_6356,N_4130,N_5281);
and U6357 (N_6357,N_4834,N_4264);
nand U6358 (N_6358,N_5819,N_4750);
or U6359 (N_6359,N_4640,N_4442);
nand U6360 (N_6360,N_5460,N_4992);
and U6361 (N_6361,N_4119,N_4275);
and U6362 (N_6362,N_4535,N_4375);
nand U6363 (N_6363,N_5646,N_5013);
nor U6364 (N_6364,N_5842,N_5583);
or U6365 (N_6365,N_4825,N_5757);
nand U6366 (N_6366,N_5856,N_4224);
or U6367 (N_6367,N_4688,N_4583);
and U6368 (N_6368,N_4123,N_5738);
nor U6369 (N_6369,N_4177,N_4198);
nor U6370 (N_6370,N_5461,N_4775);
nor U6371 (N_6371,N_5411,N_5590);
nor U6372 (N_6372,N_4843,N_4422);
and U6373 (N_6373,N_5005,N_4464);
nand U6374 (N_6374,N_4383,N_4803);
nand U6375 (N_6375,N_5109,N_4663);
and U6376 (N_6376,N_4376,N_5573);
nor U6377 (N_6377,N_5622,N_4669);
or U6378 (N_6378,N_4603,N_5612);
nor U6379 (N_6379,N_5439,N_5296);
nor U6380 (N_6380,N_5971,N_4405);
nor U6381 (N_6381,N_5839,N_4682);
nor U6382 (N_6382,N_5627,N_4008);
or U6383 (N_6383,N_5026,N_5946);
and U6384 (N_6384,N_5036,N_4432);
xnor U6385 (N_6385,N_4397,N_5007);
nor U6386 (N_6386,N_5816,N_5266);
xor U6387 (N_6387,N_5854,N_4036);
nand U6388 (N_6388,N_5456,N_4371);
or U6389 (N_6389,N_5141,N_4763);
and U6390 (N_6390,N_4404,N_5251);
or U6391 (N_6391,N_4510,N_5030);
and U6392 (N_6392,N_4125,N_4251);
nor U6393 (N_6393,N_4859,N_5051);
or U6394 (N_6394,N_4344,N_4071);
nor U6395 (N_6395,N_5315,N_5041);
nor U6396 (N_6396,N_5605,N_4455);
or U6397 (N_6397,N_5292,N_5886);
and U6398 (N_6398,N_4565,N_4514);
and U6399 (N_6399,N_5933,N_4031);
xor U6400 (N_6400,N_4879,N_4555);
and U6401 (N_6401,N_4486,N_4021);
or U6402 (N_6402,N_5645,N_4760);
nand U6403 (N_6403,N_4222,N_4257);
and U6404 (N_6404,N_5450,N_4558);
or U6405 (N_6405,N_5961,N_4440);
and U6406 (N_6406,N_5223,N_4601);
nor U6407 (N_6407,N_4886,N_4004);
or U6408 (N_6408,N_4500,N_5233);
nand U6409 (N_6409,N_4105,N_4656);
nor U6410 (N_6410,N_5205,N_4578);
and U6411 (N_6411,N_5190,N_4683);
or U6412 (N_6412,N_5592,N_4395);
xor U6413 (N_6413,N_4300,N_4415);
or U6414 (N_6414,N_4255,N_4438);
nand U6415 (N_6415,N_4568,N_4410);
and U6416 (N_6416,N_4295,N_4650);
or U6417 (N_6417,N_5830,N_5487);
and U6418 (N_6418,N_5618,N_4723);
or U6419 (N_6419,N_4499,N_5094);
xnor U6420 (N_6420,N_4632,N_5925);
nand U6421 (N_6421,N_4030,N_5749);
nand U6422 (N_6422,N_5888,N_5214);
or U6423 (N_6423,N_4936,N_5575);
xnor U6424 (N_6424,N_4653,N_5811);
nand U6425 (N_6425,N_4269,N_5654);
and U6426 (N_6426,N_5383,N_5498);
and U6427 (N_6427,N_4293,N_4967);
xor U6428 (N_6428,N_5322,N_4469);
xnor U6429 (N_6429,N_5748,N_5741);
or U6430 (N_6430,N_4904,N_5465);
nor U6431 (N_6431,N_4420,N_5964);
nor U6432 (N_6432,N_4678,N_4041);
and U6433 (N_6433,N_5956,N_5778);
and U6434 (N_6434,N_5385,N_5890);
xor U6435 (N_6435,N_4731,N_4020);
nor U6436 (N_6436,N_5152,N_5382);
nand U6437 (N_6437,N_4027,N_5037);
nor U6438 (N_6438,N_5683,N_5836);
nor U6439 (N_6439,N_5295,N_4817);
or U6440 (N_6440,N_5708,N_4042);
nand U6441 (N_6441,N_4468,N_5750);
nor U6442 (N_6442,N_4707,N_5814);
nor U6443 (N_6443,N_4314,N_5723);
and U6444 (N_6444,N_5980,N_4268);
or U6445 (N_6445,N_5244,N_4323);
and U6446 (N_6446,N_5139,N_4739);
or U6447 (N_6447,N_5168,N_5519);
xor U6448 (N_6448,N_4195,N_4562);
xnor U6449 (N_6449,N_5381,N_4325);
xor U6450 (N_6450,N_4665,N_4483);
and U6451 (N_6451,N_5445,N_5506);
nor U6452 (N_6452,N_4690,N_4019);
and U6453 (N_6453,N_4363,N_4022);
and U6454 (N_6454,N_4587,N_5587);
or U6455 (N_6455,N_4931,N_4782);
nor U6456 (N_6456,N_5617,N_5759);
nor U6457 (N_6457,N_5709,N_5389);
or U6458 (N_6458,N_4219,N_4894);
or U6459 (N_6459,N_4172,N_4009);
nand U6460 (N_6460,N_4643,N_4728);
xor U6461 (N_6461,N_5997,N_4200);
xnor U6462 (N_6462,N_5954,N_4434);
nand U6463 (N_6463,N_5696,N_5135);
or U6464 (N_6464,N_4617,N_4233);
nor U6465 (N_6465,N_5092,N_4807);
xnor U6466 (N_6466,N_5538,N_4734);
and U6467 (N_6467,N_5419,N_5607);
and U6468 (N_6468,N_4975,N_4810);
nand U6469 (N_6469,N_5540,N_5541);
nand U6470 (N_6470,N_4223,N_4595);
or U6471 (N_6471,N_4897,N_5598);
xor U6472 (N_6472,N_4928,N_5582);
and U6473 (N_6473,N_5907,N_5350);
xnor U6474 (N_6474,N_5703,N_5410);
xnor U6475 (N_6475,N_5091,N_5016);
or U6476 (N_6476,N_4126,N_5893);
nand U6477 (N_6477,N_5399,N_5331);
xnor U6478 (N_6478,N_4553,N_4842);
xor U6479 (N_6479,N_5666,N_4316);
xnor U6480 (N_6480,N_5985,N_5791);
nor U6481 (N_6481,N_4531,N_5137);
and U6482 (N_6482,N_4802,N_5149);
or U6483 (N_6483,N_5801,N_4751);
nand U6484 (N_6484,N_5534,N_4747);
xor U6485 (N_6485,N_4909,N_5420);
nor U6486 (N_6486,N_5061,N_4277);
xor U6487 (N_6487,N_4077,N_4623);
or U6488 (N_6488,N_5312,N_4720);
nor U6489 (N_6489,N_4773,N_5452);
xnor U6490 (N_6490,N_4143,N_5446);
and U6491 (N_6491,N_4780,N_4252);
and U6492 (N_6492,N_4016,N_5786);
or U6493 (N_6493,N_5029,N_4804);
nor U6494 (N_6494,N_4616,N_5765);
nand U6495 (N_6495,N_4521,N_4025);
nand U6496 (N_6496,N_5098,N_4852);
nor U6497 (N_6497,N_4918,N_4155);
nor U6498 (N_6498,N_5815,N_5394);
and U6499 (N_6499,N_5595,N_4003);
nand U6500 (N_6500,N_5790,N_4923);
nand U6501 (N_6501,N_4845,N_4285);
and U6502 (N_6502,N_5200,N_5527);
nor U6503 (N_6503,N_5367,N_4245);
nor U6504 (N_6504,N_5562,N_5319);
or U6505 (N_6505,N_5153,N_5112);
or U6506 (N_6506,N_5533,N_5744);
nor U6507 (N_6507,N_5372,N_5481);
xor U6508 (N_6508,N_4755,N_4369);
or U6509 (N_6509,N_4188,N_5858);
or U6510 (N_6510,N_4176,N_4184);
or U6511 (N_6511,N_5572,N_4040);
or U6512 (N_6512,N_4495,N_5796);
and U6513 (N_6513,N_5069,N_4820);
or U6514 (N_6514,N_5628,N_5705);
or U6515 (N_6515,N_5768,N_5732);
or U6516 (N_6516,N_4014,N_4573);
nand U6517 (N_6517,N_4309,N_4542);
nor U6518 (N_6518,N_5917,N_4645);
nor U6519 (N_6519,N_5336,N_5610);
and U6520 (N_6520,N_4947,N_4142);
nand U6521 (N_6521,N_4304,N_5780);
xnor U6522 (N_6522,N_5280,N_5637);
nand U6523 (N_6523,N_4996,N_4039);
or U6524 (N_6524,N_4649,N_4910);
or U6525 (N_6525,N_5062,N_5495);
or U6526 (N_6526,N_4674,N_4001);
nor U6527 (N_6527,N_4149,N_5717);
nor U6528 (N_6528,N_4449,N_5119);
nor U6529 (N_6529,N_4085,N_4925);
nand U6530 (N_6530,N_4394,N_4338);
and U6531 (N_6531,N_5240,N_4549);
xnor U6532 (N_6532,N_4799,N_4345);
nand U6533 (N_6533,N_5901,N_5232);
or U6534 (N_6534,N_5621,N_4253);
nor U6535 (N_6535,N_4011,N_4276);
nor U6536 (N_6536,N_5353,N_5581);
xnor U6537 (N_6537,N_5860,N_5544);
nand U6538 (N_6538,N_4063,N_5739);
and U6539 (N_6539,N_4552,N_4227);
nand U6540 (N_6540,N_4302,N_5401);
xor U6541 (N_6541,N_4289,N_5876);
and U6542 (N_6542,N_4899,N_4942);
or U6543 (N_6543,N_5074,N_5991);
and U6544 (N_6544,N_4672,N_4883);
xor U6545 (N_6545,N_4341,N_4932);
nand U6546 (N_6546,N_5851,N_4075);
xnor U6547 (N_6547,N_5965,N_4818);
and U6548 (N_6548,N_5129,N_5371);
xor U6549 (N_6549,N_5333,N_5159);
nor U6550 (N_6550,N_5711,N_5258);
nand U6551 (N_6551,N_5914,N_5829);
nand U6552 (N_6552,N_4641,N_5584);
or U6553 (N_6553,N_5588,N_5187);
nor U6554 (N_6554,N_5443,N_5318);
nor U6555 (N_6555,N_5576,N_5067);
xor U6556 (N_6556,N_5437,N_4729);
and U6557 (N_6557,N_4806,N_5277);
nand U6558 (N_6558,N_5798,N_5497);
or U6559 (N_6559,N_5855,N_5375);
nand U6560 (N_6560,N_5508,N_5442);
xor U6561 (N_6561,N_5494,N_4470);
and U6562 (N_6562,N_5189,N_5560);
or U6563 (N_6563,N_5300,N_5359);
nor U6564 (N_6564,N_5848,N_4334);
and U6565 (N_6565,N_5055,N_5158);
and U6566 (N_6566,N_4582,N_5880);
nand U6567 (N_6567,N_5784,N_4901);
and U6568 (N_6568,N_4850,N_4697);
and U6569 (N_6569,N_4900,N_4792);
nand U6570 (N_6570,N_4703,N_4828);
xor U6571 (N_6571,N_4425,N_5291);
nor U6572 (N_6572,N_4416,N_5789);
or U6573 (N_6573,N_5543,N_4855);
nand U6574 (N_6574,N_4445,N_5451);
and U6575 (N_6575,N_4358,N_4339);
or U6576 (N_6576,N_5850,N_4609);
and U6577 (N_6577,N_5426,N_4217);
or U6578 (N_6578,N_4976,N_4791);
or U6579 (N_6579,N_5285,N_4676);
and U6580 (N_6580,N_4629,N_4037);
nor U6581 (N_6581,N_5395,N_5808);
nand U6582 (N_6582,N_5818,N_4937);
and U6583 (N_6583,N_5121,N_4516);
xor U6584 (N_6584,N_5482,N_5150);
and U6585 (N_6585,N_4320,N_4547);
and U6586 (N_6586,N_5110,N_5243);
nor U6587 (N_6587,N_5729,N_4512);
and U6588 (N_6588,N_5649,N_5338);
or U6589 (N_6589,N_5932,N_5271);
or U6590 (N_6590,N_5429,N_5770);
nor U6591 (N_6591,N_5124,N_4234);
and U6592 (N_6592,N_4777,N_4398);
xor U6593 (N_6593,N_5905,N_5118);
xnor U6594 (N_6594,N_4878,N_4912);
nor U6595 (N_6595,N_4774,N_4292);
xnor U6596 (N_6596,N_5099,N_5878);
xnor U6597 (N_6597,N_4458,N_5810);
xor U6598 (N_6598,N_4702,N_4258);
and U6599 (N_6599,N_5299,N_5953);
nand U6600 (N_6600,N_5398,N_5974);
and U6601 (N_6601,N_4757,N_5269);
and U6602 (N_6602,N_4187,N_4050);
nor U6603 (N_6603,N_4896,N_5940);
nand U6604 (N_6604,N_4273,N_5270);
xor U6605 (N_6605,N_5774,N_4919);
nor U6606 (N_6606,N_5754,N_5235);
nand U6607 (N_6607,N_5824,N_4465);
nand U6608 (N_6608,N_4157,N_5254);
and U6609 (N_6609,N_5490,N_4758);
and U6610 (N_6610,N_4242,N_5122);
nor U6611 (N_6611,N_5899,N_5396);
and U6612 (N_6612,N_4692,N_5570);
and U6613 (N_6613,N_4812,N_4153);
nor U6614 (N_6614,N_5977,N_4881);
or U6615 (N_6615,N_4517,N_4232);
or U6616 (N_6616,N_4337,N_4691);
or U6617 (N_6617,N_5489,N_4969);
nand U6618 (N_6618,N_5672,N_5449);
or U6619 (N_6619,N_4443,N_4813);
or U6620 (N_6620,N_5162,N_5115);
nand U6621 (N_6621,N_4849,N_5959);
or U6622 (N_6622,N_5024,N_4480);
nand U6623 (N_6623,N_5293,N_4532);
nor U6624 (N_6624,N_5031,N_5927);
xnor U6625 (N_6625,N_4366,N_5825);
nand U6626 (N_6626,N_4501,N_5046);
xnor U6627 (N_6627,N_5081,N_5273);
nand U6628 (N_6628,N_5844,N_4012);
nand U6629 (N_6629,N_5246,N_4286);
nand U6630 (N_6630,N_4955,N_4417);
xor U6631 (N_6631,N_4864,N_4877);
and U6632 (N_6632,N_4265,N_5001);
or U6633 (N_6633,N_4662,N_5511);
nand U6634 (N_6634,N_4472,N_4481);
or U6635 (N_6635,N_5504,N_5935);
nand U6636 (N_6636,N_4576,N_4999);
or U6637 (N_6637,N_4726,N_4284);
xor U6638 (N_6638,N_5679,N_4508);
or U6639 (N_6639,N_5421,N_4929);
and U6640 (N_6640,N_4226,N_4212);
and U6641 (N_6641,N_5658,N_4637);
xor U6642 (N_6642,N_4350,N_5921);
nor U6643 (N_6643,N_4049,N_5707);
nor U6644 (N_6644,N_5405,N_4824);
or U6645 (N_6645,N_5477,N_4666);
xor U6646 (N_6646,N_5025,N_5339);
or U6647 (N_6647,N_5657,N_4244);
nor U6648 (N_6648,N_5885,N_4263);
nand U6649 (N_6649,N_5539,N_4575);
nor U6650 (N_6650,N_5368,N_5297);
xnor U6651 (N_6651,N_5468,N_4124);
nor U6652 (N_6652,N_4698,N_4715);
or U6653 (N_6653,N_4797,N_5108);
nor U6654 (N_6654,N_5873,N_4400);
or U6655 (N_6655,N_5140,N_5699);
nor U6656 (N_6656,N_5332,N_4024);
nor U6657 (N_6657,N_4107,N_5552);
nand U6658 (N_6658,N_5196,N_4236);
nand U6659 (N_6659,N_4624,N_5023);
nand U6660 (N_6660,N_4161,N_5721);
and U6661 (N_6661,N_4291,N_4159);
and U6662 (N_6662,N_5803,N_5457);
nand U6663 (N_6663,N_5447,N_5357);
or U6664 (N_6664,N_5821,N_4903);
nand U6665 (N_6665,N_5422,N_4377);
and U6666 (N_6666,N_4352,N_4362);
nor U6667 (N_6667,N_5392,N_5166);
xnor U6668 (N_6668,N_5167,N_4186);
or U6669 (N_6669,N_5239,N_4805);
or U6670 (N_6670,N_5568,N_5678);
nor U6671 (N_6671,N_5080,N_5526);
or U6672 (N_6672,N_4657,N_5620);
xnor U6673 (N_6673,N_5745,N_4534);
nor U6674 (N_6674,N_5146,N_5464);
and U6675 (N_6675,N_5114,N_4346);
and U6676 (N_6676,N_4306,N_5052);
nor U6677 (N_6677,N_5247,N_5564);
xnor U6678 (N_6678,N_5782,N_4044);
or U6679 (N_6679,N_5828,N_5516);
or U6680 (N_6680,N_5626,N_4704);
nor U6681 (N_6681,N_4638,N_5053);
nand U6682 (N_6682,N_5957,N_4297);
and U6683 (N_6683,N_5972,N_4922);
xnor U6684 (N_6684,N_4235,N_4709);
nand U6685 (N_6685,N_5643,N_4851);
nor U6686 (N_6686,N_5993,N_5638);
nor U6687 (N_6687,N_5154,N_5769);
nand U6688 (N_6688,N_5556,N_5579);
or U6689 (N_6689,N_4699,N_4494);
and U6690 (N_6690,N_4811,N_4150);
xor U6691 (N_6691,N_5514,N_4963);
nand U6692 (N_6692,N_4189,N_4930);
xnor U6693 (N_6693,N_4939,N_4367);
nor U6694 (N_6694,N_4301,N_5535);
and U6695 (N_6695,N_5775,N_5027);
or U6696 (N_6696,N_4082,N_4205);
or U6697 (N_6697,N_5597,N_5391);
xor U6698 (N_6698,N_4831,N_4907);
and U6699 (N_6699,N_5157,N_4846);
nor U6700 (N_6700,N_4060,N_4407);
nor U6701 (N_6701,N_5785,N_4924);
xor U6702 (N_6702,N_5358,N_4038);
and U6703 (N_6703,N_4972,N_4229);
xor U6704 (N_6704,N_5003,N_5202);
xor U6705 (N_6705,N_5265,N_5440);
or U6706 (N_6706,N_4446,N_5788);
or U6707 (N_6707,N_4145,N_5397);
nand U6708 (N_6708,N_5702,N_4384);
nor U6709 (N_6709,N_5528,N_5868);
or U6710 (N_6710,N_5676,N_4869);
and U6711 (N_6711,N_4591,N_5415);
and U6712 (N_6712,N_4137,N_5922);
nand U6713 (N_6713,N_4256,N_5843);
or U6714 (N_6714,N_5661,N_5085);
xnor U6715 (N_6715,N_4412,N_4815);
nand U6716 (N_6716,N_4013,N_5966);
xnor U6717 (N_6717,N_4551,N_4823);
nand U6718 (N_6718,N_4479,N_4409);
xor U6719 (N_6719,N_4127,N_4373);
and U6720 (N_6720,N_5329,N_4613);
and U6721 (N_6721,N_4474,N_5284);
or U6722 (N_6722,N_4318,N_4074);
nor U6723 (N_6723,N_5480,N_5989);
or U6724 (N_6724,N_4069,N_4584);
nor U6725 (N_6725,N_4141,N_4706);
xnor U6726 (N_6726,N_5996,N_5712);
nand U6727 (N_6727,N_5379,N_4355);
and U6728 (N_6728,N_5325,N_4741);
xor U6729 (N_6729,N_4073,N_4567);
xnor U6730 (N_6730,N_4872,N_4308);
nand U6731 (N_6731,N_5667,N_5945);
nor U6732 (N_6732,N_5852,N_4968);
and U6733 (N_6733,N_5660,N_4221);
and U6734 (N_6734,N_5823,N_4475);
or U6735 (N_6735,N_5695,N_5028);
nor U6736 (N_6736,N_4160,N_5216);
and U6737 (N_6737,N_5393,N_5458);
nand U6738 (N_6738,N_5548,N_5909);
xor U6739 (N_6739,N_4740,N_4386);
nor U6740 (N_6740,N_4213,N_4944);
and U6741 (N_6741,N_5606,N_5313);
and U6742 (N_6742,N_4421,N_5735);
or U6743 (N_6743,N_5374,N_4154);
or U6744 (N_6744,N_4220,N_4857);
or U6745 (N_6745,N_5479,N_4380);
or U6746 (N_6746,N_4327,N_5558);
and U6747 (N_6747,N_4196,N_4759);
xnor U6748 (N_6748,N_5125,N_4451);
and U6749 (N_6749,N_4045,N_5264);
or U6750 (N_6750,N_4437,N_4097);
or U6751 (N_6751,N_5086,N_4115);
or U6752 (N_6752,N_5783,N_4152);
nor U6753 (N_6753,N_4388,N_5911);
or U6754 (N_6754,N_4561,N_5340);
or U6755 (N_6755,N_5912,N_5184);
xnor U6756 (N_6756,N_4089,N_4768);
or U6757 (N_6757,N_4619,N_5904);
nand U6758 (N_6758,N_4631,N_5634);
xor U6759 (N_6759,N_4283,N_5884);
and U6760 (N_6760,N_5926,N_4484);
nor U6761 (N_6761,N_4492,N_4389);
nand U6762 (N_6762,N_4139,N_5567);
and U6763 (N_6763,N_4684,N_4419);
or U6764 (N_6764,N_4487,N_4387);
and U6765 (N_6765,N_5143,N_4513);
nor U6766 (N_6766,N_4102,N_5720);
xnor U6767 (N_6767,N_4589,N_5970);
or U6768 (N_6768,N_4429,N_4328);
xor U6769 (N_6769,N_5713,N_4029);
xnor U6770 (N_6770,N_4829,N_4998);
xnor U6771 (N_6771,N_4781,N_5928);
xnor U6772 (N_6772,N_4920,N_4664);
nor U6773 (N_6773,N_5949,N_5939);
or U6774 (N_6774,N_4307,N_4537);
and U6775 (N_6775,N_4836,N_4055);
nor U6776 (N_6776,N_4957,N_5895);
nor U6777 (N_6777,N_5351,N_5344);
and U6778 (N_6778,N_4101,N_5097);
nor U6779 (N_6779,N_5388,N_4935);
nor U6780 (N_6780,N_4630,N_4168);
xnor U6781 (N_6781,N_4116,N_5210);
nand U6782 (N_6782,N_5687,N_5674);
nand U6783 (N_6783,N_4980,N_5529);
nand U6784 (N_6784,N_4140,N_5473);
xor U6785 (N_6785,N_4095,N_5191);
and U6786 (N_6786,N_5805,N_5794);
and U6787 (N_6787,N_5724,N_5287);
or U6788 (N_6788,N_5518,N_5102);
nor U6789 (N_6789,N_4406,N_5944);
and U6790 (N_6790,N_4693,N_4765);
and U6791 (N_6791,N_5586,N_4488);
or U6792 (N_6792,N_4093,N_4312);
nor U6793 (N_6793,N_5704,N_4163);
xnor U6794 (N_6794,N_5044,N_5671);
xnor U6795 (N_6795,N_4908,N_5865);
and U6796 (N_6796,N_5453,N_4655);
xnor U6797 (N_6797,N_5478,N_5840);
and U6798 (N_6798,N_4118,N_5123);
xor U6799 (N_6799,N_4241,N_4280);
nand U6800 (N_6800,N_4239,N_5262);
nor U6801 (N_6801,N_4895,N_5219);
and U6802 (N_6802,N_5531,N_4822);
or U6803 (N_6803,N_4250,N_4906);
or U6804 (N_6804,N_4744,N_4543);
or U6805 (N_6805,N_5002,N_4091);
nor U6806 (N_6806,N_5321,N_5722);
or U6807 (N_6807,N_5867,N_4724);
nand U6808 (N_6808,N_5043,N_5772);
or U6809 (N_6809,N_5793,N_4450);
nand U6810 (N_6810,N_4569,N_5820);
or U6811 (N_6811,N_5364,N_5307);
xnor U6812 (N_6812,N_4506,N_4032);
nand U6813 (N_6813,N_5689,N_4209);
or U6814 (N_6814,N_5565,N_5669);
nand U6815 (N_6815,N_4490,N_4973);
or U6816 (N_6816,N_4958,N_5462);
xor U6817 (N_6817,N_5763,N_4436);
nor U6818 (N_6818,N_5806,N_4771);
nor U6819 (N_6819,N_5662,N_4204);
nand U6820 (N_6820,N_5499,N_5630);
xnor U6821 (N_6821,N_4120,N_4524);
xor U6822 (N_6822,N_5653,N_4164);
and U6823 (N_6823,N_4214,N_5404);
nand U6824 (N_6824,N_5134,N_4786);
or U6825 (N_6825,N_4875,N_4079);
xor U6826 (N_6826,N_5551,N_4681);
xor U6827 (N_6827,N_4156,N_4977);
and U6828 (N_6828,N_5403,N_5197);
nor U6829 (N_6829,N_4712,N_4015);
nor U6830 (N_6830,N_4330,N_5349);
or U6831 (N_6831,N_4062,N_4737);
and U6832 (N_6832,N_5599,N_4721);
or U6833 (N_6833,N_4183,N_5656);
nor U6834 (N_6834,N_5609,N_5414);
xnor U6835 (N_6835,N_4006,N_4556);
xnor U6836 (N_6836,N_5360,N_5853);
nand U6837 (N_6837,N_5042,N_5311);
or U6838 (N_6838,N_5864,N_4310);
xnor U6839 (N_6839,N_4199,N_5743);
nand U6840 (N_6840,N_4991,N_5604);
or U6841 (N_6841,N_4026,N_4753);
and U6842 (N_6842,N_5369,N_4887);
or U6843 (N_6843,N_4000,N_5427);
or U6844 (N_6844,N_4940,N_5253);
xnor U6845 (N_6845,N_5373,N_4686);
xnor U6846 (N_6846,N_5475,N_4303);
nor U6847 (N_6847,N_5505,N_4602);
or U6848 (N_6848,N_4916,N_4182);
nand U6849 (N_6849,N_4868,N_4225);
nand U6850 (N_6850,N_4203,N_5217);
xor U6851 (N_6851,N_4374,N_4028);
nor U6852 (N_6852,N_4194,N_4372);
and U6853 (N_6853,N_5779,N_5608);
nand U6854 (N_6854,N_5228,N_4121);
and U6855 (N_6855,N_5826,N_4054);
nor U6856 (N_6856,N_5355,N_5435);
and U6857 (N_6857,N_5726,N_5117);
nor U6858 (N_6858,N_4322,N_5525);
xor U6859 (N_6859,N_4423,N_5407);
xnor U6860 (N_6860,N_5065,N_4809);
xnor U6861 (N_6861,N_5603,N_5978);
nand U6862 (N_6862,N_5260,N_5536);
nor U6863 (N_6863,N_5929,N_5252);
xor U6864 (N_6864,N_4921,N_4779);
xor U6865 (N_6865,N_4439,N_5845);
and U6866 (N_6866,N_5103,N_5113);
and U6867 (N_6867,N_5182,N_5838);
nor U6868 (N_6868,N_5613,N_4113);
nand U6869 (N_6869,N_4175,N_5021);
or U6870 (N_6870,N_5194,N_4260);
or U6871 (N_6871,N_4068,N_5466);
and U6872 (N_6872,N_4668,N_5327);
or U6873 (N_6873,N_4435,N_4658);
xnor U6874 (N_6874,N_5897,N_4819);
nand U6875 (N_6875,N_5513,N_4800);
and U6876 (N_6876,N_4190,N_4636);
nor U6877 (N_6877,N_5869,N_4279);
nand U6878 (N_6878,N_4206,N_4870);
and U6879 (N_6879,N_4769,N_4112);
nand U6880 (N_6880,N_5950,N_5101);
xor U6881 (N_6881,N_4563,N_5212);
nand U6882 (N_6882,N_5267,N_4621);
xnor U6883 (N_6883,N_5038,N_5862);
nor U6884 (N_6884,N_4191,N_5684);
and U6885 (N_6885,N_4288,N_5365);
or U6886 (N_6886,N_5834,N_4088);
xnor U6887 (N_6887,N_4945,N_4033);
nor U6888 (N_6888,N_4527,N_5326);
and U6889 (N_6889,N_5837,N_4351);
or U6890 (N_6890,N_4057,N_4732);
and U6891 (N_6891,N_4607,N_5503);
and U6892 (N_6892,N_4882,N_5777);
or U6893 (N_6893,N_4520,N_5088);
nand U6894 (N_6894,N_5919,N_5237);
and U6895 (N_6895,N_5984,N_4670);
and U6896 (N_6896,N_4722,N_4913);
nand U6897 (N_6897,N_4390,N_4611);
nor U6898 (N_6898,N_4861,N_5795);
nor U6899 (N_6899,N_5761,N_4385);
or U6900 (N_6900,N_4231,N_4902);
xor U6901 (N_6901,N_4661,N_5033);
xor U6902 (N_6902,N_5255,N_4964);
and U6903 (N_6903,N_4505,N_5631);
and U6904 (N_6904,N_5766,N_4860);
and U6905 (N_6905,N_4067,N_5802);
xnor U6906 (N_6906,N_5238,N_4078);
or U6907 (N_6907,N_5063,N_4761);
xnor U6908 (N_6908,N_4675,N_4010);
nand U6909 (N_6909,N_5602,N_5335);
or U6910 (N_6910,N_5846,N_5983);
and U6911 (N_6911,N_4215,N_4798);
or U6912 (N_6912,N_4315,N_5418);
or U6913 (N_6913,N_5680,N_4411);
nand U6914 (N_6914,N_5773,N_4965);
nand U6915 (N_6915,N_5275,N_4540);
nand U6916 (N_6916,N_4381,N_5384);
or U6917 (N_6917,N_5107,N_4005);
or U6918 (N_6918,N_5577,N_4790);
and U6919 (N_6919,N_5668,N_5467);
xor U6920 (N_6920,N_5892,N_5537);
xnor U6921 (N_6921,N_4876,N_5659);
and U6922 (N_6922,N_5986,N_4677);
and U6923 (N_6923,N_5871,N_4414);
or U6924 (N_6924,N_4642,N_4835);
nor U6925 (N_6925,N_4941,N_5682);
xnor U6926 (N_6926,N_5771,N_5133);
xnor U6927 (N_6927,N_5981,N_5948);
nand U6928 (N_6928,N_5454,N_4056);
and U6929 (N_6929,N_4990,N_5747);
and U6930 (N_6930,N_5142,N_5276);
xor U6931 (N_6931,N_5279,N_4319);
xor U6932 (N_6932,N_5192,N_4296);
and U6933 (N_6933,N_4981,N_5841);
or U6934 (N_6934,N_5222,N_4456);
nor U6935 (N_6935,N_4396,N_5740);
nor U6936 (N_6936,N_4452,N_5304);
nor U6937 (N_6937,N_5413,N_4247);
nand U6938 (N_6938,N_5054,N_4379);
xor U6939 (N_6939,N_5015,N_5136);
xor U6940 (N_6940,N_5431,N_4335);
and U6941 (N_6941,N_5644,N_5416);
nor U6942 (N_6942,N_5387,N_5208);
xor U6943 (N_6943,N_4862,N_4357);
or U6944 (N_6944,N_5087,N_5076);
nor U6945 (N_6945,N_4428,N_5673);
and U6946 (N_6946,N_5746,N_4084);
xor U6947 (N_6947,N_4104,N_4133);
xnor U6948 (N_6948,N_4444,N_4332);
nor U6949 (N_6949,N_5090,N_4368);
nor U6950 (N_6950,N_4392,N_5095);
nor U6951 (N_6951,N_4970,N_5377);
xor U6952 (N_6952,N_5554,N_5547);
and U6953 (N_6953,N_5792,N_4708);
nor U6954 (N_6954,N_4430,N_5804);
xor U6955 (N_6955,N_5259,N_5557);
and U6956 (N_6956,N_4826,N_4117);
nand U6957 (N_6957,N_4518,N_5776);
nor U6958 (N_6958,N_5221,N_4208);
nor U6959 (N_6959,N_5915,N_5975);
xnor U6960 (N_6960,N_5148,N_4626);
or U6961 (N_6961,N_5180,N_4651);
xnor U6962 (N_6962,N_4572,N_5160);
xor U6963 (N_6963,N_5633,N_4716);
nor U6964 (N_6964,N_4473,N_5290);
nor U6965 (N_6965,N_4497,N_5022);
and U6966 (N_6966,N_5866,N_5624);
nor U6967 (N_6967,N_4103,N_4960);
and U6968 (N_6968,N_4756,N_4694);
nor U6969 (N_6969,N_5725,N_5799);
xnor U6970 (N_6970,N_5900,N_4529);
nand U6971 (N_6971,N_4738,N_5967);
and U6972 (N_6972,N_5501,N_5496);
or U6973 (N_6973,N_5361,N_5882);
and U6974 (N_6974,N_5463,N_5089);
nand U6975 (N_6975,N_4266,N_5507);
nand U6976 (N_6976,N_4281,N_5176);
xnor U6977 (N_6977,N_5952,N_5242);
nor U6978 (N_6978,N_5963,N_4342);
nor U6979 (N_6979,N_5916,N_5515);
or U6980 (N_6980,N_5218,N_4324);
xnor U6981 (N_6981,N_5693,N_5261);
or U6982 (N_6982,N_4171,N_4598);
and U6983 (N_6983,N_4382,N_4867);
xnor U6984 (N_6984,N_4580,N_5234);
and U6985 (N_6985,N_4402,N_5476);
nor U6986 (N_6986,N_4778,N_5175);
nand U6987 (N_6987,N_5096,N_4644);
and U6988 (N_6988,N_5049,N_5183);
xor U6989 (N_6989,N_4954,N_4333);
xor U6990 (N_6990,N_5084,N_5812);
nand U6991 (N_6991,N_4108,N_4165);
nor U6992 (N_6992,N_4571,N_5050);
nand U6993 (N_6993,N_4840,N_5906);
and U6994 (N_6994,N_5731,N_5423);
nand U6995 (N_6995,N_5230,N_5755);
nor U6996 (N_6996,N_5317,N_4952);
xor U6997 (N_6997,N_5390,N_5542);
and U6998 (N_6998,N_4566,N_5859);
or U6999 (N_6999,N_5204,N_5623);
nand U7000 (N_7000,N_4276,N_4076);
and U7001 (N_7001,N_4273,N_5415);
nand U7002 (N_7002,N_4105,N_5568);
xnor U7003 (N_7003,N_5250,N_5434);
nand U7004 (N_7004,N_4249,N_5365);
nand U7005 (N_7005,N_5169,N_4513);
nand U7006 (N_7006,N_5470,N_4908);
and U7007 (N_7007,N_5984,N_4791);
xnor U7008 (N_7008,N_4232,N_5621);
nor U7009 (N_7009,N_4886,N_4698);
nand U7010 (N_7010,N_4448,N_4185);
and U7011 (N_7011,N_5789,N_4254);
xor U7012 (N_7012,N_5696,N_4965);
or U7013 (N_7013,N_4161,N_5234);
xor U7014 (N_7014,N_5039,N_4911);
or U7015 (N_7015,N_4961,N_5866);
nand U7016 (N_7016,N_4370,N_5864);
or U7017 (N_7017,N_4126,N_5008);
nand U7018 (N_7018,N_4911,N_4439);
or U7019 (N_7019,N_5737,N_4261);
or U7020 (N_7020,N_4395,N_5641);
or U7021 (N_7021,N_5316,N_5453);
nand U7022 (N_7022,N_4370,N_5699);
and U7023 (N_7023,N_4675,N_4242);
and U7024 (N_7024,N_5847,N_5235);
nor U7025 (N_7025,N_5220,N_5329);
or U7026 (N_7026,N_4005,N_5543);
or U7027 (N_7027,N_5558,N_5758);
nor U7028 (N_7028,N_4761,N_5563);
nor U7029 (N_7029,N_5507,N_4360);
xnor U7030 (N_7030,N_4473,N_4798);
xnor U7031 (N_7031,N_5072,N_5001);
nor U7032 (N_7032,N_4295,N_4644);
nor U7033 (N_7033,N_4597,N_5972);
or U7034 (N_7034,N_5019,N_5788);
and U7035 (N_7035,N_4693,N_5034);
nand U7036 (N_7036,N_5735,N_4393);
xor U7037 (N_7037,N_4034,N_5291);
nor U7038 (N_7038,N_5601,N_4100);
nand U7039 (N_7039,N_5404,N_5572);
nor U7040 (N_7040,N_5140,N_4619);
or U7041 (N_7041,N_5020,N_4374);
xor U7042 (N_7042,N_5362,N_5809);
and U7043 (N_7043,N_5829,N_4375);
and U7044 (N_7044,N_5235,N_4630);
or U7045 (N_7045,N_4480,N_5540);
xnor U7046 (N_7046,N_5281,N_5239);
nand U7047 (N_7047,N_4236,N_5375);
or U7048 (N_7048,N_4968,N_4282);
or U7049 (N_7049,N_5799,N_5528);
xnor U7050 (N_7050,N_5409,N_4500);
and U7051 (N_7051,N_4566,N_5903);
and U7052 (N_7052,N_5935,N_4635);
nand U7053 (N_7053,N_4869,N_4340);
or U7054 (N_7054,N_4953,N_4180);
or U7055 (N_7055,N_4055,N_5264);
and U7056 (N_7056,N_5799,N_4049);
nor U7057 (N_7057,N_5413,N_4110);
xor U7058 (N_7058,N_5723,N_5564);
or U7059 (N_7059,N_4352,N_5837);
nor U7060 (N_7060,N_4757,N_5525);
and U7061 (N_7061,N_5793,N_4072);
or U7062 (N_7062,N_5432,N_5428);
nand U7063 (N_7063,N_4497,N_5013);
and U7064 (N_7064,N_4603,N_5020);
nand U7065 (N_7065,N_5932,N_5697);
and U7066 (N_7066,N_5950,N_5680);
nand U7067 (N_7067,N_4956,N_4264);
nand U7068 (N_7068,N_4839,N_4581);
nand U7069 (N_7069,N_5202,N_5217);
or U7070 (N_7070,N_5626,N_5789);
and U7071 (N_7071,N_5057,N_5292);
and U7072 (N_7072,N_5774,N_4658);
and U7073 (N_7073,N_5905,N_4950);
xor U7074 (N_7074,N_5703,N_4212);
and U7075 (N_7075,N_5635,N_5388);
xor U7076 (N_7076,N_5724,N_4929);
nand U7077 (N_7077,N_4897,N_4548);
nand U7078 (N_7078,N_5104,N_5276);
or U7079 (N_7079,N_5012,N_5466);
nand U7080 (N_7080,N_5342,N_4154);
and U7081 (N_7081,N_4188,N_4104);
xnor U7082 (N_7082,N_5216,N_5820);
and U7083 (N_7083,N_5366,N_5152);
nand U7084 (N_7084,N_4758,N_4489);
xor U7085 (N_7085,N_4904,N_4278);
xor U7086 (N_7086,N_5345,N_4710);
xnor U7087 (N_7087,N_4095,N_4495);
or U7088 (N_7088,N_5233,N_4529);
or U7089 (N_7089,N_5558,N_4376);
nand U7090 (N_7090,N_4748,N_4138);
nand U7091 (N_7091,N_4541,N_4483);
nand U7092 (N_7092,N_5181,N_4716);
xnor U7093 (N_7093,N_4782,N_5742);
nor U7094 (N_7094,N_4505,N_4239);
or U7095 (N_7095,N_5607,N_4305);
nor U7096 (N_7096,N_5957,N_4128);
and U7097 (N_7097,N_4764,N_5040);
nand U7098 (N_7098,N_4695,N_5497);
nand U7099 (N_7099,N_5095,N_4876);
and U7100 (N_7100,N_5726,N_5416);
xnor U7101 (N_7101,N_5224,N_4958);
xnor U7102 (N_7102,N_4090,N_4380);
nand U7103 (N_7103,N_4048,N_5575);
and U7104 (N_7104,N_5250,N_4390);
or U7105 (N_7105,N_4913,N_5761);
nand U7106 (N_7106,N_4514,N_4685);
nand U7107 (N_7107,N_5913,N_5568);
nand U7108 (N_7108,N_5546,N_4875);
and U7109 (N_7109,N_4929,N_4091);
or U7110 (N_7110,N_4605,N_5683);
nand U7111 (N_7111,N_5081,N_5307);
or U7112 (N_7112,N_5815,N_5642);
xnor U7113 (N_7113,N_4861,N_4909);
or U7114 (N_7114,N_5105,N_4676);
or U7115 (N_7115,N_5382,N_5368);
xor U7116 (N_7116,N_4385,N_5129);
or U7117 (N_7117,N_5047,N_4648);
and U7118 (N_7118,N_5866,N_5428);
xor U7119 (N_7119,N_5762,N_5455);
xnor U7120 (N_7120,N_5569,N_4020);
nand U7121 (N_7121,N_4533,N_4319);
nor U7122 (N_7122,N_4689,N_4219);
or U7123 (N_7123,N_4037,N_5104);
nor U7124 (N_7124,N_5173,N_4471);
nor U7125 (N_7125,N_4448,N_4545);
xor U7126 (N_7126,N_5119,N_4666);
and U7127 (N_7127,N_5716,N_4176);
and U7128 (N_7128,N_4068,N_5127);
nand U7129 (N_7129,N_5633,N_5840);
xor U7130 (N_7130,N_5679,N_4251);
nand U7131 (N_7131,N_4940,N_4669);
nor U7132 (N_7132,N_5071,N_4073);
nand U7133 (N_7133,N_5990,N_4295);
or U7134 (N_7134,N_4232,N_4596);
xor U7135 (N_7135,N_5796,N_5080);
xor U7136 (N_7136,N_5356,N_4669);
or U7137 (N_7137,N_5848,N_4623);
and U7138 (N_7138,N_4683,N_5641);
nand U7139 (N_7139,N_4810,N_4688);
or U7140 (N_7140,N_5577,N_4035);
or U7141 (N_7141,N_5901,N_5663);
nand U7142 (N_7142,N_4827,N_4565);
nand U7143 (N_7143,N_5972,N_4966);
xnor U7144 (N_7144,N_5487,N_4726);
xnor U7145 (N_7145,N_4208,N_5537);
nand U7146 (N_7146,N_5960,N_5413);
nor U7147 (N_7147,N_5945,N_5414);
nor U7148 (N_7148,N_4410,N_4051);
and U7149 (N_7149,N_4991,N_4490);
and U7150 (N_7150,N_5659,N_5111);
nor U7151 (N_7151,N_5686,N_5791);
and U7152 (N_7152,N_4031,N_5383);
nor U7153 (N_7153,N_5002,N_5748);
nand U7154 (N_7154,N_5519,N_5080);
or U7155 (N_7155,N_4395,N_4055);
nand U7156 (N_7156,N_4193,N_5780);
nor U7157 (N_7157,N_5495,N_4066);
nor U7158 (N_7158,N_4087,N_5000);
xnor U7159 (N_7159,N_5635,N_5873);
nor U7160 (N_7160,N_4732,N_4099);
nand U7161 (N_7161,N_5230,N_4006);
nand U7162 (N_7162,N_5310,N_4478);
nand U7163 (N_7163,N_4323,N_4641);
xor U7164 (N_7164,N_5336,N_4945);
and U7165 (N_7165,N_5236,N_5400);
and U7166 (N_7166,N_4909,N_4120);
nor U7167 (N_7167,N_4285,N_5772);
or U7168 (N_7168,N_4019,N_5214);
and U7169 (N_7169,N_4793,N_5793);
and U7170 (N_7170,N_5778,N_4682);
and U7171 (N_7171,N_5357,N_4509);
and U7172 (N_7172,N_5577,N_4345);
or U7173 (N_7173,N_5583,N_4743);
or U7174 (N_7174,N_4689,N_4878);
or U7175 (N_7175,N_4994,N_5258);
and U7176 (N_7176,N_4965,N_4910);
and U7177 (N_7177,N_5728,N_4041);
and U7178 (N_7178,N_5919,N_4030);
nand U7179 (N_7179,N_5217,N_5618);
and U7180 (N_7180,N_5072,N_5721);
nor U7181 (N_7181,N_5268,N_5086);
or U7182 (N_7182,N_4042,N_5559);
and U7183 (N_7183,N_4095,N_5011);
and U7184 (N_7184,N_5199,N_5712);
nor U7185 (N_7185,N_4434,N_4539);
nand U7186 (N_7186,N_5149,N_4249);
xnor U7187 (N_7187,N_4629,N_4565);
nor U7188 (N_7188,N_5885,N_5153);
and U7189 (N_7189,N_4857,N_5824);
nand U7190 (N_7190,N_5935,N_4274);
and U7191 (N_7191,N_4461,N_4036);
xor U7192 (N_7192,N_4300,N_5437);
nor U7193 (N_7193,N_4825,N_4300);
or U7194 (N_7194,N_4434,N_5597);
nand U7195 (N_7195,N_5145,N_4701);
xnor U7196 (N_7196,N_4072,N_5925);
nand U7197 (N_7197,N_4719,N_5075);
xor U7198 (N_7198,N_5001,N_4817);
or U7199 (N_7199,N_5131,N_4101);
nor U7200 (N_7200,N_5418,N_4716);
or U7201 (N_7201,N_5454,N_4782);
and U7202 (N_7202,N_5855,N_5114);
or U7203 (N_7203,N_4761,N_5483);
nand U7204 (N_7204,N_5715,N_5662);
nor U7205 (N_7205,N_5348,N_4196);
nor U7206 (N_7206,N_5520,N_4772);
or U7207 (N_7207,N_4561,N_4659);
nor U7208 (N_7208,N_5530,N_5021);
nor U7209 (N_7209,N_4483,N_5021);
nor U7210 (N_7210,N_4579,N_4722);
nand U7211 (N_7211,N_5976,N_5543);
or U7212 (N_7212,N_5057,N_5808);
nor U7213 (N_7213,N_5746,N_4491);
or U7214 (N_7214,N_5830,N_5893);
nor U7215 (N_7215,N_5351,N_4885);
xnor U7216 (N_7216,N_4142,N_4793);
nand U7217 (N_7217,N_4987,N_5957);
nand U7218 (N_7218,N_5968,N_4140);
or U7219 (N_7219,N_4230,N_5276);
nor U7220 (N_7220,N_5008,N_4110);
xnor U7221 (N_7221,N_5497,N_4644);
and U7222 (N_7222,N_4919,N_4984);
nand U7223 (N_7223,N_4409,N_4262);
xor U7224 (N_7224,N_4795,N_4552);
or U7225 (N_7225,N_5460,N_4705);
xor U7226 (N_7226,N_4262,N_5938);
and U7227 (N_7227,N_5634,N_4911);
xor U7228 (N_7228,N_4006,N_4474);
or U7229 (N_7229,N_4786,N_5880);
and U7230 (N_7230,N_5977,N_4424);
xnor U7231 (N_7231,N_5687,N_4776);
xnor U7232 (N_7232,N_5083,N_5939);
or U7233 (N_7233,N_4504,N_5465);
and U7234 (N_7234,N_4267,N_5951);
or U7235 (N_7235,N_4475,N_4111);
or U7236 (N_7236,N_4271,N_5852);
or U7237 (N_7237,N_5533,N_5799);
nand U7238 (N_7238,N_5271,N_5668);
or U7239 (N_7239,N_4496,N_4005);
nand U7240 (N_7240,N_4669,N_5031);
nand U7241 (N_7241,N_4564,N_4237);
or U7242 (N_7242,N_5962,N_5184);
nand U7243 (N_7243,N_4360,N_5845);
nor U7244 (N_7244,N_4379,N_4194);
nand U7245 (N_7245,N_5771,N_4410);
and U7246 (N_7246,N_5588,N_4905);
and U7247 (N_7247,N_5400,N_5895);
or U7248 (N_7248,N_4664,N_4304);
xor U7249 (N_7249,N_5460,N_4025);
or U7250 (N_7250,N_4831,N_5828);
and U7251 (N_7251,N_4213,N_4136);
and U7252 (N_7252,N_5408,N_4467);
nor U7253 (N_7253,N_5135,N_4764);
xor U7254 (N_7254,N_4151,N_4184);
or U7255 (N_7255,N_5831,N_5893);
xnor U7256 (N_7256,N_5870,N_5799);
xnor U7257 (N_7257,N_5940,N_5675);
or U7258 (N_7258,N_4553,N_4507);
or U7259 (N_7259,N_4385,N_4742);
nand U7260 (N_7260,N_4665,N_4213);
nor U7261 (N_7261,N_5317,N_4200);
nand U7262 (N_7262,N_5298,N_4026);
nor U7263 (N_7263,N_4476,N_5299);
or U7264 (N_7264,N_5505,N_4491);
or U7265 (N_7265,N_4888,N_5298);
nand U7266 (N_7266,N_4578,N_5209);
nand U7267 (N_7267,N_5334,N_5095);
nand U7268 (N_7268,N_5718,N_4226);
nand U7269 (N_7269,N_5563,N_5861);
and U7270 (N_7270,N_4876,N_5163);
or U7271 (N_7271,N_4910,N_4498);
xor U7272 (N_7272,N_4954,N_5051);
xor U7273 (N_7273,N_5473,N_5537);
nor U7274 (N_7274,N_5394,N_4349);
xnor U7275 (N_7275,N_5967,N_5059);
or U7276 (N_7276,N_5837,N_4184);
nand U7277 (N_7277,N_4384,N_4842);
and U7278 (N_7278,N_5958,N_4516);
xor U7279 (N_7279,N_4182,N_5958);
and U7280 (N_7280,N_4945,N_4047);
nor U7281 (N_7281,N_5493,N_4439);
nand U7282 (N_7282,N_5116,N_4900);
and U7283 (N_7283,N_5461,N_4739);
nand U7284 (N_7284,N_4954,N_4314);
nor U7285 (N_7285,N_4032,N_4791);
nor U7286 (N_7286,N_4478,N_4386);
and U7287 (N_7287,N_5958,N_5822);
nand U7288 (N_7288,N_4303,N_4872);
and U7289 (N_7289,N_4356,N_4046);
or U7290 (N_7290,N_4093,N_5931);
or U7291 (N_7291,N_5165,N_5717);
nand U7292 (N_7292,N_5896,N_5058);
xor U7293 (N_7293,N_5001,N_4150);
or U7294 (N_7294,N_5550,N_4801);
and U7295 (N_7295,N_4561,N_4167);
or U7296 (N_7296,N_4040,N_4283);
xor U7297 (N_7297,N_5717,N_4900);
nand U7298 (N_7298,N_4133,N_5928);
or U7299 (N_7299,N_4361,N_4242);
nand U7300 (N_7300,N_4937,N_4174);
nor U7301 (N_7301,N_4307,N_4109);
nand U7302 (N_7302,N_5140,N_5432);
nor U7303 (N_7303,N_5887,N_5766);
nor U7304 (N_7304,N_4777,N_4015);
nor U7305 (N_7305,N_5458,N_4685);
nor U7306 (N_7306,N_4039,N_4648);
nor U7307 (N_7307,N_4469,N_4218);
xnor U7308 (N_7308,N_5119,N_5990);
or U7309 (N_7309,N_4016,N_4913);
or U7310 (N_7310,N_4040,N_5312);
nand U7311 (N_7311,N_4767,N_5676);
or U7312 (N_7312,N_5278,N_5190);
nand U7313 (N_7313,N_5018,N_5528);
xor U7314 (N_7314,N_5286,N_5306);
xor U7315 (N_7315,N_5362,N_4433);
and U7316 (N_7316,N_5245,N_5196);
and U7317 (N_7317,N_5211,N_5628);
and U7318 (N_7318,N_4924,N_5199);
or U7319 (N_7319,N_4188,N_4180);
xor U7320 (N_7320,N_4292,N_4233);
and U7321 (N_7321,N_4498,N_5349);
or U7322 (N_7322,N_4886,N_4867);
nand U7323 (N_7323,N_5614,N_5236);
xor U7324 (N_7324,N_4652,N_4088);
or U7325 (N_7325,N_5055,N_5705);
xnor U7326 (N_7326,N_5426,N_4172);
nand U7327 (N_7327,N_4457,N_4428);
nand U7328 (N_7328,N_4089,N_4851);
nor U7329 (N_7329,N_4681,N_4801);
nor U7330 (N_7330,N_4276,N_5138);
xor U7331 (N_7331,N_4503,N_4861);
nor U7332 (N_7332,N_5554,N_4433);
nand U7333 (N_7333,N_4082,N_4331);
or U7334 (N_7334,N_4070,N_4658);
xnor U7335 (N_7335,N_4313,N_4237);
nor U7336 (N_7336,N_5283,N_5583);
and U7337 (N_7337,N_5192,N_4393);
nor U7338 (N_7338,N_4998,N_5877);
and U7339 (N_7339,N_5968,N_4054);
xor U7340 (N_7340,N_4428,N_4476);
nor U7341 (N_7341,N_4520,N_4499);
xnor U7342 (N_7342,N_5571,N_4221);
nor U7343 (N_7343,N_4569,N_5003);
nand U7344 (N_7344,N_5430,N_4705);
xor U7345 (N_7345,N_4630,N_4260);
nor U7346 (N_7346,N_4764,N_5087);
and U7347 (N_7347,N_4307,N_5803);
xnor U7348 (N_7348,N_4626,N_5563);
xnor U7349 (N_7349,N_5877,N_4260);
or U7350 (N_7350,N_5944,N_5988);
xor U7351 (N_7351,N_4492,N_5826);
and U7352 (N_7352,N_4692,N_4507);
nand U7353 (N_7353,N_5871,N_4023);
xor U7354 (N_7354,N_4769,N_5972);
xor U7355 (N_7355,N_5943,N_4102);
nand U7356 (N_7356,N_5375,N_4208);
xor U7357 (N_7357,N_4470,N_4735);
nand U7358 (N_7358,N_5986,N_4099);
nor U7359 (N_7359,N_4521,N_5409);
nand U7360 (N_7360,N_4780,N_5201);
and U7361 (N_7361,N_4111,N_5443);
nor U7362 (N_7362,N_5503,N_4876);
or U7363 (N_7363,N_5260,N_4825);
and U7364 (N_7364,N_4303,N_5453);
or U7365 (N_7365,N_5374,N_5641);
or U7366 (N_7366,N_4690,N_5033);
xor U7367 (N_7367,N_4160,N_4575);
xnor U7368 (N_7368,N_5850,N_4555);
xnor U7369 (N_7369,N_4976,N_4574);
or U7370 (N_7370,N_5046,N_4807);
or U7371 (N_7371,N_4355,N_4845);
nor U7372 (N_7372,N_5128,N_5107);
nor U7373 (N_7373,N_5311,N_5510);
and U7374 (N_7374,N_4463,N_4039);
and U7375 (N_7375,N_5941,N_5165);
or U7376 (N_7376,N_5634,N_5474);
or U7377 (N_7377,N_4577,N_5907);
and U7378 (N_7378,N_4694,N_4125);
xor U7379 (N_7379,N_5288,N_4303);
or U7380 (N_7380,N_5236,N_4634);
and U7381 (N_7381,N_4204,N_5472);
nor U7382 (N_7382,N_4071,N_4431);
and U7383 (N_7383,N_5524,N_5693);
and U7384 (N_7384,N_4915,N_4285);
nand U7385 (N_7385,N_5798,N_4846);
or U7386 (N_7386,N_5895,N_4307);
and U7387 (N_7387,N_5532,N_4006);
xnor U7388 (N_7388,N_4928,N_4651);
or U7389 (N_7389,N_4481,N_5381);
nand U7390 (N_7390,N_4169,N_5347);
nor U7391 (N_7391,N_4360,N_5510);
nor U7392 (N_7392,N_4364,N_5641);
nor U7393 (N_7393,N_4466,N_4201);
or U7394 (N_7394,N_5443,N_5538);
or U7395 (N_7395,N_5835,N_5770);
nor U7396 (N_7396,N_4246,N_5030);
and U7397 (N_7397,N_4873,N_4425);
nand U7398 (N_7398,N_5026,N_5753);
and U7399 (N_7399,N_4905,N_5551);
nand U7400 (N_7400,N_4959,N_5596);
nor U7401 (N_7401,N_5138,N_4273);
or U7402 (N_7402,N_4017,N_5455);
xnor U7403 (N_7403,N_4757,N_5329);
nand U7404 (N_7404,N_5200,N_4226);
and U7405 (N_7405,N_4710,N_5474);
nand U7406 (N_7406,N_4271,N_4519);
and U7407 (N_7407,N_5229,N_5352);
xnor U7408 (N_7408,N_4215,N_4324);
and U7409 (N_7409,N_4376,N_5716);
nor U7410 (N_7410,N_5538,N_4692);
nand U7411 (N_7411,N_4487,N_4534);
nand U7412 (N_7412,N_4696,N_4118);
nand U7413 (N_7413,N_5193,N_5863);
and U7414 (N_7414,N_5828,N_5415);
and U7415 (N_7415,N_5907,N_5891);
nor U7416 (N_7416,N_4336,N_5028);
nor U7417 (N_7417,N_5484,N_4960);
xor U7418 (N_7418,N_5125,N_5463);
nor U7419 (N_7419,N_4424,N_4871);
nand U7420 (N_7420,N_5267,N_5331);
xor U7421 (N_7421,N_4367,N_4895);
or U7422 (N_7422,N_4069,N_4037);
nor U7423 (N_7423,N_5015,N_5944);
xor U7424 (N_7424,N_5039,N_4438);
or U7425 (N_7425,N_5132,N_5921);
and U7426 (N_7426,N_4895,N_4127);
or U7427 (N_7427,N_4553,N_5205);
or U7428 (N_7428,N_5156,N_4755);
nand U7429 (N_7429,N_5318,N_5998);
nand U7430 (N_7430,N_5295,N_4010);
xnor U7431 (N_7431,N_5418,N_4895);
nor U7432 (N_7432,N_4987,N_4123);
or U7433 (N_7433,N_5218,N_5660);
nor U7434 (N_7434,N_4644,N_5952);
nand U7435 (N_7435,N_4559,N_4723);
xor U7436 (N_7436,N_5054,N_5894);
nor U7437 (N_7437,N_5297,N_4392);
or U7438 (N_7438,N_5874,N_4119);
nor U7439 (N_7439,N_4095,N_5413);
nand U7440 (N_7440,N_4274,N_4622);
nor U7441 (N_7441,N_5602,N_5680);
nand U7442 (N_7442,N_5485,N_5622);
or U7443 (N_7443,N_4019,N_5677);
xor U7444 (N_7444,N_5374,N_4311);
or U7445 (N_7445,N_5957,N_5407);
and U7446 (N_7446,N_5516,N_5096);
or U7447 (N_7447,N_4205,N_4997);
nand U7448 (N_7448,N_4294,N_5862);
xor U7449 (N_7449,N_5339,N_5468);
and U7450 (N_7450,N_5046,N_4875);
nand U7451 (N_7451,N_4602,N_5889);
and U7452 (N_7452,N_4642,N_4142);
nand U7453 (N_7453,N_5147,N_4901);
nor U7454 (N_7454,N_5817,N_5391);
xor U7455 (N_7455,N_4301,N_5346);
xnor U7456 (N_7456,N_4438,N_4770);
nor U7457 (N_7457,N_5571,N_4343);
nor U7458 (N_7458,N_4053,N_5784);
nor U7459 (N_7459,N_4523,N_4419);
nand U7460 (N_7460,N_4563,N_4218);
or U7461 (N_7461,N_4327,N_4956);
nand U7462 (N_7462,N_4325,N_5769);
nor U7463 (N_7463,N_5006,N_4796);
nor U7464 (N_7464,N_5069,N_5149);
and U7465 (N_7465,N_5208,N_5876);
or U7466 (N_7466,N_5990,N_5611);
and U7467 (N_7467,N_4555,N_4531);
or U7468 (N_7468,N_4988,N_4764);
and U7469 (N_7469,N_4322,N_5393);
or U7470 (N_7470,N_5389,N_5841);
nor U7471 (N_7471,N_5257,N_5194);
and U7472 (N_7472,N_4167,N_5251);
nand U7473 (N_7473,N_5259,N_4331);
nor U7474 (N_7474,N_4187,N_4948);
nand U7475 (N_7475,N_4650,N_5998);
nor U7476 (N_7476,N_5098,N_5595);
and U7477 (N_7477,N_4325,N_5127);
and U7478 (N_7478,N_4242,N_5594);
or U7479 (N_7479,N_4246,N_4476);
nor U7480 (N_7480,N_5558,N_4574);
xnor U7481 (N_7481,N_4577,N_5268);
and U7482 (N_7482,N_4036,N_5832);
and U7483 (N_7483,N_4323,N_4151);
nand U7484 (N_7484,N_4855,N_5652);
and U7485 (N_7485,N_4642,N_4564);
or U7486 (N_7486,N_4188,N_4958);
xor U7487 (N_7487,N_4018,N_4821);
and U7488 (N_7488,N_5029,N_5544);
nand U7489 (N_7489,N_4095,N_5123);
or U7490 (N_7490,N_4419,N_5200);
nand U7491 (N_7491,N_4775,N_4444);
nor U7492 (N_7492,N_4798,N_5351);
or U7493 (N_7493,N_4951,N_4135);
and U7494 (N_7494,N_5547,N_4715);
or U7495 (N_7495,N_5768,N_4863);
xnor U7496 (N_7496,N_5238,N_4393);
nor U7497 (N_7497,N_4649,N_4681);
and U7498 (N_7498,N_4317,N_4323);
xor U7499 (N_7499,N_4563,N_4592);
or U7500 (N_7500,N_4171,N_5270);
xor U7501 (N_7501,N_4965,N_4571);
nor U7502 (N_7502,N_4222,N_4317);
or U7503 (N_7503,N_5236,N_5164);
nor U7504 (N_7504,N_4687,N_4550);
and U7505 (N_7505,N_5442,N_4658);
and U7506 (N_7506,N_5104,N_4345);
nand U7507 (N_7507,N_5349,N_5854);
nor U7508 (N_7508,N_5332,N_5038);
and U7509 (N_7509,N_4447,N_4629);
nand U7510 (N_7510,N_4657,N_4065);
nand U7511 (N_7511,N_5184,N_4040);
or U7512 (N_7512,N_4582,N_5377);
or U7513 (N_7513,N_5824,N_4643);
and U7514 (N_7514,N_5304,N_5320);
xor U7515 (N_7515,N_4671,N_5991);
nand U7516 (N_7516,N_4044,N_4836);
xnor U7517 (N_7517,N_4808,N_4414);
nand U7518 (N_7518,N_4550,N_4070);
nor U7519 (N_7519,N_5051,N_5930);
xnor U7520 (N_7520,N_4930,N_5746);
nor U7521 (N_7521,N_4930,N_4114);
nor U7522 (N_7522,N_4897,N_4504);
nand U7523 (N_7523,N_4400,N_4368);
and U7524 (N_7524,N_5343,N_5432);
and U7525 (N_7525,N_5419,N_4617);
and U7526 (N_7526,N_4921,N_5776);
nand U7527 (N_7527,N_4059,N_5320);
and U7528 (N_7528,N_5725,N_4602);
or U7529 (N_7529,N_5141,N_4107);
and U7530 (N_7530,N_5471,N_5468);
nand U7531 (N_7531,N_5459,N_5703);
nor U7532 (N_7532,N_4867,N_5785);
xor U7533 (N_7533,N_5330,N_5955);
nand U7534 (N_7534,N_4843,N_5344);
xnor U7535 (N_7535,N_5361,N_5960);
nor U7536 (N_7536,N_5210,N_5983);
xnor U7537 (N_7537,N_5396,N_5508);
nor U7538 (N_7538,N_4061,N_4569);
nand U7539 (N_7539,N_5972,N_4722);
and U7540 (N_7540,N_5381,N_5790);
or U7541 (N_7541,N_5966,N_4831);
or U7542 (N_7542,N_5395,N_4966);
nand U7543 (N_7543,N_5429,N_5606);
nor U7544 (N_7544,N_4876,N_4373);
and U7545 (N_7545,N_4451,N_5459);
nor U7546 (N_7546,N_5401,N_5722);
nor U7547 (N_7547,N_5504,N_5313);
and U7548 (N_7548,N_4224,N_4004);
nor U7549 (N_7549,N_4629,N_4479);
nand U7550 (N_7550,N_4372,N_4647);
nor U7551 (N_7551,N_4226,N_4935);
nand U7552 (N_7552,N_5104,N_4502);
nand U7553 (N_7553,N_5124,N_4733);
nand U7554 (N_7554,N_5123,N_4431);
nand U7555 (N_7555,N_5591,N_4813);
and U7556 (N_7556,N_4394,N_4101);
or U7557 (N_7557,N_5892,N_5361);
nor U7558 (N_7558,N_4651,N_5752);
nor U7559 (N_7559,N_5956,N_4408);
nor U7560 (N_7560,N_4488,N_5383);
or U7561 (N_7561,N_4396,N_5927);
nand U7562 (N_7562,N_4704,N_4841);
nor U7563 (N_7563,N_4023,N_5490);
xnor U7564 (N_7564,N_5666,N_4470);
nand U7565 (N_7565,N_5311,N_5172);
or U7566 (N_7566,N_4774,N_4203);
nor U7567 (N_7567,N_4601,N_4460);
xor U7568 (N_7568,N_5524,N_4571);
xnor U7569 (N_7569,N_5754,N_4314);
or U7570 (N_7570,N_4816,N_4046);
or U7571 (N_7571,N_5934,N_4881);
and U7572 (N_7572,N_4653,N_5077);
nor U7573 (N_7573,N_4641,N_5510);
xor U7574 (N_7574,N_5373,N_4657);
or U7575 (N_7575,N_4329,N_5514);
xor U7576 (N_7576,N_4413,N_5109);
or U7577 (N_7577,N_4453,N_5004);
and U7578 (N_7578,N_4107,N_5351);
nand U7579 (N_7579,N_4861,N_5324);
nand U7580 (N_7580,N_5466,N_5840);
or U7581 (N_7581,N_5728,N_4487);
or U7582 (N_7582,N_5767,N_5441);
xnor U7583 (N_7583,N_5219,N_4546);
xor U7584 (N_7584,N_4645,N_4423);
xor U7585 (N_7585,N_4086,N_5484);
or U7586 (N_7586,N_4030,N_5219);
or U7587 (N_7587,N_5702,N_4068);
nand U7588 (N_7588,N_4057,N_4747);
nand U7589 (N_7589,N_5666,N_5602);
xor U7590 (N_7590,N_4962,N_5816);
nor U7591 (N_7591,N_5708,N_4468);
or U7592 (N_7592,N_4689,N_4479);
xnor U7593 (N_7593,N_5715,N_4663);
or U7594 (N_7594,N_4487,N_5772);
nor U7595 (N_7595,N_4027,N_5301);
and U7596 (N_7596,N_4137,N_4982);
xor U7597 (N_7597,N_4871,N_5372);
xnor U7598 (N_7598,N_5732,N_5179);
nand U7599 (N_7599,N_5786,N_5699);
and U7600 (N_7600,N_4579,N_5205);
nor U7601 (N_7601,N_4064,N_5089);
nand U7602 (N_7602,N_5295,N_5753);
nor U7603 (N_7603,N_5615,N_4709);
and U7604 (N_7604,N_4433,N_4052);
and U7605 (N_7605,N_4472,N_5390);
nand U7606 (N_7606,N_5180,N_5148);
xor U7607 (N_7607,N_4283,N_5161);
nor U7608 (N_7608,N_4461,N_4202);
or U7609 (N_7609,N_4158,N_4250);
or U7610 (N_7610,N_4626,N_4242);
nand U7611 (N_7611,N_5821,N_4137);
or U7612 (N_7612,N_5992,N_5452);
nand U7613 (N_7613,N_5262,N_4368);
and U7614 (N_7614,N_5771,N_5212);
nor U7615 (N_7615,N_5039,N_4525);
nor U7616 (N_7616,N_5161,N_5946);
nor U7617 (N_7617,N_5196,N_5774);
nor U7618 (N_7618,N_4662,N_5301);
or U7619 (N_7619,N_4022,N_4509);
and U7620 (N_7620,N_4530,N_5693);
or U7621 (N_7621,N_4895,N_5922);
nor U7622 (N_7622,N_4597,N_5028);
and U7623 (N_7623,N_4666,N_4948);
nor U7624 (N_7624,N_5194,N_5153);
or U7625 (N_7625,N_5638,N_4049);
and U7626 (N_7626,N_5247,N_5323);
or U7627 (N_7627,N_5117,N_4225);
nand U7628 (N_7628,N_4734,N_5637);
and U7629 (N_7629,N_5060,N_4016);
and U7630 (N_7630,N_5676,N_5074);
nor U7631 (N_7631,N_5242,N_5899);
xnor U7632 (N_7632,N_5237,N_5281);
nand U7633 (N_7633,N_5230,N_5122);
xor U7634 (N_7634,N_5150,N_4083);
and U7635 (N_7635,N_4626,N_4176);
nand U7636 (N_7636,N_5593,N_5773);
xnor U7637 (N_7637,N_5524,N_5874);
or U7638 (N_7638,N_4083,N_5656);
and U7639 (N_7639,N_4262,N_5900);
and U7640 (N_7640,N_4125,N_5854);
and U7641 (N_7641,N_4349,N_4312);
nand U7642 (N_7642,N_4515,N_5737);
or U7643 (N_7643,N_4511,N_4316);
or U7644 (N_7644,N_4682,N_4912);
nand U7645 (N_7645,N_5263,N_5271);
and U7646 (N_7646,N_5946,N_5975);
nand U7647 (N_7647,N_4128,N_4817);
or U7648 (N_7648,N_5867,N_5909);
nand U7649 (N_7649,N_5400,N_5136);
xnor U7650 (N_7650,N_4750,N_5763);
xnor U7651 (N_7651,N_4056,N_5804);
xnor U7652 (N_7652,N_4760,N_4023);
xor U7653 (N_7653,N_4048,N_5276);
xor U7654 (N_7654,N_5762,N_5800);
nand U7655 (N_7655,N_5167,N_4853);
or U7656 (N_7656,N_4545,N_5541);
nor U7657 (N_7657,N_5246,N_4602);
xor U7658 (N_7658,N_4432,N_5014);
and U7659 (N_7659,N_4941,N_4070);
xnor U7660 (N_7660,N_4280,N_5350);
and U7661 (N_7661,N_5347,N_4046);
xor U7662 (N_7662,N_4707,N_5649);
nand U7663 (N_7663,N_5935,N_5459);
nor U7664 (N_7664,N_4644,N_5290);
or U7665 (N_7665,N_4733,N_5280);
xnor U7666 (N_7666,N_4663,N_4594);
xor U7667 (N_7667,N_4975,N_4626);
nand U7668 (N_7668,N_4064,N_4021);
and U7669 (N_7669,N_5485,N_5763);
xnor U7670 (N_7670,N_5873,N_4853);
and U7671 (N_7671,N_4371,N_5202);
xnor U7672 (N_7672,N_4264,N_5125);
nor U7673 (N_7673,N_4912,N_5275);
or U7674 (N_7674,N_4356,N_5742);
nor U7675 (N_7675,N_4411,N_5206);
nor U7676 (N_7676,N_4952,N_4583);
xor U7677 (N_7677,N_5201,N_4066);
or U7678 (N_7678,N_5733,N_4421);
or U7679 (N_7679,N_5861,N_4722);
nor U7680 (N_7680,N_5361,N_4453);
or U7681 (N_7681,N_4778,N_4097);
nand U7682 (N_7682,N_5025,N_5680);
or U7683 (N_7683,N_5053,N_5658);
nand U7684 (N_7684,N_4818,N_4953);
nand U7685 (N_7685,N_5961,N_4105);
or U7686 (N_7686,N_4351,N_4916);
xor U7687 (N_7687,N_4237,N_4178);
and U7688 (N_7688,N_4325,N_4450);
or U7689 (N_7689,N_5241,N_4700);
xor U7690 (N_7690,N_5609,N_4075);
nor U7691 (N_7691,N_5136,N_4448);
nor U7692 (N_7692,N_4187,N_5566);
xor U7693 (N_7693,N_4215,N_4997);
nor U7694 (N_7694,N_4119,N_4797);
nor U7695 (N_7695,N_4150,N_4849);
or U7696 (N_7696,N_4520,N_5483);
or U7697 (N_7697,N_4893,N_4299);
xnor U7698 (N_7698,N_4079,N_5750);
or U7699 (N_7699,N_4533,N_4390);
nand U7700 (N_7700,N_4647,N_4499);
or U7701 (N_7701,N_4969,N_4922);
xor U7702 (N_7702,N_4623,N_4697);
xnor U7703 (N_7703,N_4330,N_5010);
xnor U7704 (N_7704,N_5825,N_4737);
nor U7705 (N_7705,N_4798,N_5434);
xor U7706 (N_7706,N_5106,N_5163);
xor U7707 (N_7707,N_4017,N_4619);
or U7708 (N_7708,N_4971,N_4576);
xor U7709 (N_7709,N_5277,N_5695);
nand U7710 (N_7710,N_5327,N_4339);
nand U7711 (N_7711,N_4434,N_4927);
nor U7712 (N_7712,N_5728,N_5981);
nor U7713 (N_7713,N_4968,N_4511);
nor U7714 (N_7714,N_5171,N_4422);
nor U7715 (N_7715,N_4085,N_4562);
or U7716 (N_7716,N_5023,N_4082);
or U7717 (N_7717,N_4176,N_4008);
or U7718 (N_7718,N_5911,N_4485);
nor U7719 (N_7719,N_5470,N_5085);
xor U7720 (N_7720,N_5334,N_4710);
xor U7721 (N_7721,N_5417,N_5401);
nand U7722 (N_7722,N_4691,N_5358);
or U7723 (N_7723,N_4034,N_5833);
nor U7724 (N_7724,N_5953,N_4752);
nor U7725 (N_7725,N_4270,N_5045);
and U7726 (N_7726,N_4488,N_4791);
or U7727 (N_7727,N_4288,N_5791);
nor U7728 (N_7728,N_4330,N_5234);
nor U7729 (N_7729,N_5982,N_5351);
xnor U7730 (N_7730,N_5856,N_4642);
and U7731 (N_7731,N_4655,N_4315);
nor U7732 (N_7732,N_5133,N_5100);
nand U7733 (N_7733,N_5882,N_4116);
xnor U7734 (N_7734,N_4622,N_5381);
and U7735 (N_7735,N_4482,N_4724);
nand U7736 (N_7736,N_4801,N_4712);
nand U7737 (N_7737,N_5359,N_4766);
nand U7738 (N_7738,N_4504,N_5144);
and U7739 (N_7739,N_4741,N_4617);
xnor U7740 (N_7740,N_4074,N_5394);
nand U7741 (N_7741,N_5649,N_5111);
xor U7742 (N_7742,N_5117,N_5166);
nand U7743 (N_7743,N_5032,N_5373);
nor U7744 (N_7744,N_4187,N_5219);
or U7745 (N_7745,N_4165,N_5854);
xor U7746 (N_7746,N_5370,N_4035);
nor U7747 (N_7747,N_5024,N_4359);
nor U7748 (N_7748,N_4737,N_5352);
nand U7749 (N_7749,N_5534,N_5163);
or U7750 (N_7750,N_5209,N_5570);
nand U7751 (N_7751,N_5620,N_5579);
nand U7752 (N_7752,N_5607,N_4786);
nand U7753 (N_7753,N_5906,N_5804);
nor U7754 (N_7754,N_5046,N_5591);
and U7755 (N_7755,N_4917,N_4469);
nor U7756 (N_7756,N_4345,N_5564);
xor U7757 (N_7757,N_5332,N_4606);
or U7758 (N_7758,N_4009,N_4046);
or U7759 (N_7759,N_5323,N_4415);
or U7760 (N_7760,N_4621,N_5392);
nor U7761 (N_7761,N_4562,N_5185);
nand U7762 (N_7762,N_5644,N_5891);
nand U7763 (N_7763,N_4726,N_4590);
xnor U7764 (N_7764,N_4199,N_5654);
xnor U7765 (N_7765,N_4166,N_4061);
nand U7766 (N_7766,N_4565,N_5209);
nand U7767 (N_7767,N_4757,N_5787);
and U7768 (N_7768,N_4829,N_5114);
nand U7769 (N_7769,N_5558,N_5640);
nand U7770 (N_7770,N_4193,N_4930);
nor U7771 (N_7771,N_4113,N_5510);
or U7772 (N_7772,N_5085,N_5149);
and U7773 (N_7773,N_5213,N_4431);
and U7774 (N_7774,N_5205,N_5410);
and U7775 (N_7775,N_5096,N_4467);
nand U7776 (N_7776,N_5551,N_5838);
nor U7777 (N_7777,N_4406,N_5790);
and U7778 (N_7778,N_4091,N_4534);
xor U7779 (N_7779,N_4023,N_4110);
nand U7780 (N_7780,N_4857,N_4604);
nand U7781 (N_7781,N_5915,N_4880);
nand U7782 (N_7782,N_5786,N_4411);
or U7783 (N_7783,N_5264,N_5542);
or U7784 (N_7784,N_4027,N_5445);
or U7785 (N_7785,N_4852,N_4327);
and U7786 (N_7786,N_4714,N_4517);
or U7787 (N_7787,N_4821,N_4232);
or U7788 (N_7788,N_4832,N_5126);
or U7789 (N_7789,N_4377,N_4463);
nor U7790 (N_7790,N_5032,N_5657);
nor U7791 (N_7791,N_4541,N_4951);
nor U7792 (N_7792,N_5765,N_5088);
or U7793 (N_7793,N_5534,N_5462);
xor U7794 (N_7794,N_5869,N_5203);
and U7795 (N_7795,N_5750,N_5713);
nand U7796 (N_7796,N_5079,N_4826);
or U7797 (N_7797,N_4503,N_4837);
nand U7798 (N_7798,N_5599,N_5322);
and U7799 (N_7799,N_4105,N_5029);
xor U7800 (N_7800,N_5574,N_4801);
nor U7801 (N_7801,N_5829,N_5599);
nand U7802 (N_7802,N_4313,N_4752);
xnor U7803 (N_7803,N_5507,N_4372);
or U7804 (N_7804,N_4032,N_4570);
and U7805 (N_7805,N_4766,N_4387);
nor U7806 (N_7806,N_5502,N_5909);
nor U7807 (N_7807,N_4822,N_4698);
or U7808 (N_7808,N_4695,N_4765);
or U7809 (N_7809,N_5142,N_5493);
and U7810 (N_7810,N_5427,N_5175);
xnor U7811 (N_7811,N_5576,N_4509);
nand U7812 (N_7812,N_5421,N_5216);
or U7813 (N_7813,N_5693,N_4883);
or U7814 (N_7814,N_4756,N_5895);
and U7815 (N_7815,N_5674,N_4352);
nand U7816 (N_7816,N_4925,N_5455);
and U7817 (N_7817,N_4331,N_4411);
or U7818 (N_7818,N_4394,N_4571);
or U7819 (N_7819,N_4875,N_5650);
nor U7820 (N_7820,N_5730,N_5667);
and U7821 (N_7821,N_4932,N_4900);
nand U7822 (N_7822,N_5765,N_5331);
and U7823 (N_7823,N_5862,N_4013);
and U7824 (N_7824,N_5370,N_4897);
nor U7825 (N_7825,N_5792,N_4039);
xnor U7826 (N_7826,N_4743,N_5996);
xor U7827 (N_7827,N_5097,N_5733);
or U7828 (N_7828,N_5150,N_4229);
nand U7829 (N_7829,N_5067,N_4645);
nor U7830 (N_7830,N_4844,N_5906);
nor U7831 (N_7831,N_4663,N_5432);
nor U7832 (N_7832,N_4220,N_5987);
xnor U7833 (N_7833,N_4040,N_5425);
nand U7834 (N_7834,N_4580,N_5937);
xnor U7835 (N_7835,N_5977,N_5607);
nor U7836 (N_7836,N_4596,N_5127);
and U7837 (N_7837,N_5013,N_4147);
nor U7838 (N_7838,N_5571,N_4388);
and U7839 (N_7839,N_5546,N_5083);
and U7840 (N_7840,N_4908,N_5416);
nor U7841 (N_7841,N_5262,N_5399);
or U7842 (N_7842,N_4680,N_4410);
or U7843 (N_7843,N_4811,N_5038);
or U7844 (N_7844,N_4042,N_4907);
and U7845 (N_7845,N_4894,N_5180);
nor U7846 (N_7846,N_4586,N_4800);
or U7847 (N_7847,N_5997,N_4750);
nand U7848 (N_7848,N_5042,N_5152);
xnor U7849 (N_7849,N_4293,N_5926);
and U7850 (N_7850,N_5708,N_5377);
or U7851 (N_7851,N_4968,N_4452);
nor U7852 (N_7852,N_4652,N_5215);
xor U7853 (N_7853,N_5392,N_4803);
and U7854 (N_7854,N_4174,N_4612);
nand U7855 (N_7855,N_5781,N_5530);
or U7856 (N_7856,N_5285,N_4034);
xor U7857 (N_7857,N_5602,N_5605);
nor U7858 (N_7858,N_5242,N_4551);
and U7859 (N_7859,N_4573,N_4065);
nand U7860 (N_7860,N_4449,N_4511);
nand U7861 (N_7861,N_5249,N_4287);
nand U7862 (N_7862,N_5324,N_4766);
nor U7863 (N_7863,N_4284,N_4940);
or U7864 (N_7864,N_4400,N_5053);
nor U7865 (N_7865,N_5565,N_5620);
nor U7866 (N_7866,N_5738,N_5776);
or U7867 (N_7867,N_5651,N_4909);
and U7868 (N_7868,N_5578,N_4274);
or U7869 (N_7869,N_5161,N_4604);
nand U7870 (N_7870,N_5027,N_5657);
or U7871 (N_7871,N_4086,N_4158);
nor U7872 (N_7872,N_5955,N_4242);
nand U7873 (N_7873,N_5097,N_4266);
nor U7874 (N_7874,N_5469,N_5216);
and U7875 (N_7875,N_4955,N_4095);
and U7876 (N_7876,N_4022,N_4726);
xnor U7877 (N_7877,N_5189,N_4137);
and U7878 (N_7878,N_4089,N_4761);
and U7879 (N_7879,N_5849,N_4262);
xnor U7880 (N_7880,N_5762,N_5015);
nor U7881 (N_7881,N_5572,N_5866);
xor U7882 (N_7882,N_4017,N_4391);
nand U7883 (N_7883,N_5544,N_4744);
xnor U7884 (N_7884,N_4032,N_4601);
xnor U7885 (N_7885,N_4460,N_5849);
nand U7886 (N_7886,N_5005,N_4806);
xor U7887 (N_7887,N_5400,N_4508);
nand U7888 (N_7888,N_4123,N_4666);
nor U7889 (N_7889,N_4204,N_4805);
nor U7890 (N_7890,N_4868,N_4711);
xnor U7891 (N_7891,N_5768,N_5227);
and U7892 (N_7892,N_5346,N_4487);
and U7893 (N_7893,N_5292,N_4174);
xor U7894 (N_7894,N_5982,N_4025);
and U7895 (N_7895,N_5173,N_5812);
nand U7896 (N_7896,N_5151,N_4788);
and U7897 (N_7897,N_4580,N_5766);
nor U7898 (N_7898,N_5926,N_5744);
xor U7899 (N_7899,N_4173,N_5742);
nor U7900 (N_7900,N_5193,N_5287);
and U7901 (N_7901,N_4232,N_5636);
and U7902 (N_7902,N_5649,N_4694);
xor U7903 (N_7903,N_4420,N_5391);
and U7904 (N_7904,N_4878,N_5357);
or U7905 (N_7905,N_4829,N_4446);
nand U7906 (N_7906,N_4681,N_4013);
and U7907 (N_7907,N_4678,N_5174);
nor U7908 (N_7908,N_5196,N_4608);
nand U7909 (N_7909,N_4650,N_5887);
nand U7910 (N_7910,N_5528,N_4444);
or U7911 (N_7911,N_4188,N_4721);
or U7912 (N_7912,N_5430,N_5787);
nor U7913 (N_7913,N_4806,N_5776);
nand U7914 (N_7914,N_5019,N_5338);
and U7915 (N_7915,N_5422,N_4982);
and U7916 (N_7916,N_5085,N_5097);
and U7917 (N_7917,N_5305,N_4229);
and U7918 (N_7918,N_5328,N_4520);
nor U7919 (N_7919,N_4701,N_4250);
or U7920 (N_7920,N_4740,N_5993);
xor U7921 (N_7921,N_5939,N_5419);
and U7922 (N_7922,N_4442,N_5161);
nand U7923 (N_7923,N_4634,N_5661);
or U7924 (N_7924,N_5384,N_5271);
xnor U7925 (N_7925,N_5430,N_5616);
and U7926 (N_7926,N_5583,N_5261);
and U7927 (N_7927,N_5660,N_5982);
and U7928 (N_7928,N_4291,N_5175);
xnor U7929 (N_7929,N_4134,N_5035);
or U7930 (N_7930,N_5842,N_4057);
or U7931 (N_7931,N_4768,N_5829);
xor U7932 (N_7932,N_4672,N_5588);
xnor U7933 (N_7933,N_4178,N_4052);
xnor U7934 (N_7934,N_4059,N_5538);
nand U7935 (N_7935,N_4642,N_4092);
and U7936 (N_7936,N_4460,N_4134);
nand U7937 (N_7937,N_4141,N_4114);
nor U7938 (N_7938,N_5398,N_4713);
xnor U7939 (N_7939,N_5229,N_5566);
and U7940 (N_7940,N_5017,N_5140);
nand U7941 (N_7941,N_5692,N_5740);
and U7942 (N_7942,N_4944,N_4592);
nand U7943 (N_7943,N_5404,N_5655);
nand U7944 (N_7944,N_4587,N_5084);
or U7945 (N_7945,N_5685,N_5865);
nor U7946 (N_7946,N_5947,N_4115);
and U7947 (N_7947,N_5136,N_4101);
and U7948 (N_7948,N_5848,N_4127);
or U7949 (N_7949,N_5212,N_5138);
xnor U7950 (N_7950,N_4735,N_5366);
and U7951 (N_7951,N_4360,N_4396);
nor U7952 (N_7952,N_4667,N_4561);
and U7953 (N_7953,N_5980,N_4253);
nor U7954 (N_7954,N_5834,N_4316);
nand U7955 (N_7955,N_5759,N_4809);
or U7956 (N_7956,N_5244,N_4712);
or U7957 (N_7957,N_4768,N_5008);
or U7958 (N_7958,N_5779,N_5247);
and U7959 (N_7959,N_5913,N_4231);
or U7960 (N_7960,N_4073,N_5742);
xor U7961 (N_7961,N_4256,N_5822);
and U7962 (N_7962,N_4728,N_5879);
xor U7963 (N_7963,N_5007,N_4226);
or U7964 (N_7964,N_5003,N_4232);
xor U7965 (N_7965,N_5782,N_4539);
or U7966 (N_7966,N_5225,N_5966);
nor U7967 (N_7967,N_5659,N_5694);
nor U7968 (N_7968,N_5417,N_5377);
or U7969 (N_7969,N_4555,N_5442);
nand U7970 (N_7970,N_5931,N_5664);
nand U7971 (N_7971,N_4727,N_5530);
and U7972 (N_7972,N_4956,N_4587);
nand U7973 (N_7973,N_4946,N_4470);
and U7974 (N_7974,N_5307,N_5880);
or U7975 (N_7975,N_4376,N_5675);
nand U7976 (N_7976,N_4278,N_5482);
and U7977 (N_7977,N_5279,N_5837);
or U7978 (N_7978,N_5058,N_4530);
xor U7979 (N_7979,N_5522,N_4688);
nor U7980 (N_7980,N_4983,N_5991);
or U7981 (N_7981,N_4019,N_4374);
nor U7982 (N_7982,N_4073,N_5976);
nor U7983 (N_7983,N_4997,N_4149);
or U7984 (N_7984,N_4887,N_5190);
nand U7985 (N_7985,N_5125,N_5036);
nand U7986 (N_7986,N_5072,N_5203);
or U7987 (N_7987,N_4929,N_4467);
nor U7988 (N_7988,N_5615,N_4948);
xor U7989 (N_7989,N_4625,N_4977);
nor U7990 (N_7990,N_4498,N_4018);
nand U7991 (N_7991,N_5613,N_5501);
xor U7992 (N_7992,N_5754,N_5795);
nor U7993 (N_7993,N_5960,N_5576);
or U7994 (N_7994,N_4054,N_5141);
xor U7995 (N_7995,N_4274,N_4443);
nand U7996 (N_7996,N_5249,N_5307);
xor U7997 (N_7997,N_5787,N_5097);
or U7998 (N_7998,N_4992,N_4289);
xor U7999 (N_7999,N_5927,N_5077);
nor U8000 (N_8000,N_7948,N_7546);
and U8001 (N_8001,N_6910,N_6812);
or U8002 (N_8002,N_6636,N_7424);
xor U8003 (N_8003,N_7585,N_7276);
nand U8004 (N_8004,N_6359,N_6756);
or U8005 (N_8005,N_7639,N_7590);
xor U8006 (N_8006,N_6045,N_6343);
and U8007 (N_8007,N_6839,N_6856);
or U8008 (N_8008,N_6918,N_7441);
or U8009 (N_8009,N_6491,N_6282);
and U8010 (N_8010,N_7662,N_7569);
or U8011 (N_8011,N_7636,N_7248);
nor U8012 (N_8012,N_6390,N_7297);
and U8013 (N_8013,N_6240,N_6564);
and U8014 (N_8014,N_7182,N_6220);
or U8015 (N_8015,N_6297,N_7567);
xor U8016 (N_8016,N_6345,N_7169);
and U8017 (N_8017,N_7093,N_7750);
xor U8018 (N_8018,N_6973,N_7570);
xor U8019 (N_8019,N_7521,N_6960);
xor U8020 (N_8020,N_7753,N_6871);
nor U8021 (N_8021,N_7299,N_6201);
nor U8022 (N_8022,N_7392,N_6916);
and U8023 (N_8023,N_6843,N_6629);
nor U8024 (N_8024,N_6891,N_7519);
or U8025 (N_8025,N_7409,N_6801);
nor U8026 (N_8026,N_6167,N_6389);
or U8027 (N_8027,N_7732,N_6117);
or U8028 (N_8028,N_6983,N_7443);
nand U8029 (N_8029,N_6402,N_7418);
or U8030 (N_8030,N_7097,N_6293);
and U8031 (N_8031,N_7000,N_7808);
nor U8032 (N_8032,N_6006,N_7188);
nand U8033 (N_8033,N_6273,N_6506);
and U8034 (N_8034,N_7963,N_7795);
xnor U8035 (N_8035,N_6846,N_6906);
or U8036 (N_8036,N_7448,N_6138);
nand U8037 (N_8037,N_6952,N_7610);
nand U8038 (N_8038,N_6352,N_7246);
or U8039 (N_8039,N_6903,N_6662);
or U8040 (N_8040,N_6232,N_7778);
xor U8041 (N_8041,N_7178,N_6521);
nor U8042 (N_8042,N_7458,N_6575);
nor U8043 (N_8043,N_6294,N_6008);
and U8044 (N_8044,N_7369,N_7417);
and U8045 (N_8045,N_7958,N_6434);
nor U8046 (N_8046,N_7515,N_6866);
nor U8047 (N_8047,N_7062,N_6417);
nor U8048 (N_8048,N_7647,N_6333);
and U8049 (N_8049,N_7997,N_6030);
xor U8050 (N_8050,N_7875,N_6311);
and U8051 (N_8051,N_6925,N_7649);
nor U8052 (N_8052,N_6032,N_6215);
or U8053 (N_8053,N_6195,N_6815);
and U8054 (N_8054,N_6436,N_7942);
or U8055 (N_8055,N_6658,N_7333);
nand U8056 (N_8056,N_7588,N_7261);
and U8057 (N_8057,N_6139,N_6414);
xnor U8058 (N_8058,N_7586,N_6931);
and U8059 (N_8059,N_6994,N_6135);
or U8060 (N_8060,N_6487,N_6698);
and U8061 (N_8061,N_6314,N_7728);
xor U8062 (N_8062,N_7716,N_7596);
nor U8063 (N_8063,N_7275,N_6927);
xnor U8064 (N_8064,N_7819,N_7134);
nand U8065 (N_8065,N_7863,N_7425);
nand U8066 (N_8066,N_7430,N_6611);
nor U8067 (N_8067,N_6500,N_6486);
or U8068 (N_8068,N_7220,N_7108);
nand U8069 (N_8069,N_6111,N_6258);
nor U8070 (N_8070,N_7506,N_6723);
and U8071 (N_8071,N_7339,N_6589);
nor U8072 (N_8072,N_6554,N_7125);
or U8073 (N_8073,N_6078,N_6048);
or U8074 (N_8074,N_7051,N_6882);
and U8075 (N_8075,N_6769,N_6539);
nand U8076 (N_8076,N_6420,N_7995);
or U8077 (N_8077,N_6367,N_6504);
nor U8078 (N_8078,N_7208,N_7311);
or U8079 (N_8079,N_7754,N_6844);
nor U8080 (N_8080,N_7766,N_7207);
nor U8081 (N_8081,N_7849,N_7096);
and U8082 (N_8082,N_7526,N_6835);
nand U8083 (N_8083,N_7354,N_6895);
nand U8084 (N_8084,N_6216,N_6003);
xor U8085 (N_8085,N_7810,N_6643);
xor U8086 (N_8086,N_7440,N_7495);
nand U8087 (N_8087,N_7996,N_6696);
nor U8088 (N_8088,N_6922,N_7789);
and U8089 (N_8089,N_7070,N_7155);
xor U8090 (N_8090,N_6851,N_7676);
nor U8091 (N_8091,N_6919,N_7575);
nor U8092 (N_8092,N_6312,N_7666);
nand U8093 (N_8093,N_6509,N_7204);
or U8094 (N_8094,N_6650,N_6457);
xor U8095 (N_8095,N_7370,N_6710);
nand U8096 (N_8096,N_6369,N_7289);
or U8097 (N_8097,N_6630,N_6256);
and U8098 (N_8098,N_7288,N_6495);
and U8099 (N_8099,N_7039,N_7098);
nand U8100 (N_8100,N_7391,N_7340);
and U8101 (N_8101,N_6674,N_7637);
xor U8102 (N_8102,N_7697,N_6248);
nand U8103 (N_8103,N_6178,N_6870);
nand U8104 (N_8104,N_7386,N_7847);
xor U8105 (N_8105,N_7171,N_6415);
and U8106 (N_8106,N_7974,N_7233);
nand U8107 (N_8107,N_7555,N_7444);
nand U8108 (N_8108,N_7263,N_7041);
and U8109 (N_8109,N_6577,N_6641);
nor U8110 (N_8110,N_7293,N_7900);
nor U8111 (N_8111,N_6088,N_6704);
nand U8112 (N_8112,N_6626,N_6172);
or U8113 (N_8113,N_7490,N_6059);
and U8114 (N_8114,N_6091,N_6286);
or U8115 (N_8115,N_6096,N_6766);
xnor U8116 (N_8116,N_7027,N_6202);
xnor U8117 (N_8117,N_6174,N_6310);
and U8118 (N_8118,N_6515,N_7739);
xor U8119 (N_8119,N_6183,N_6671);
xor U8120 (N_8120,N_7497,N_6961);
or U8121 (N_8121,N_6763,N_7422);
or U8122 (N_8122,N_7015,N_7309);
or U8123 (N_8123,N_7326,N_7775);
nand U8124 (N_8124,N_7376,N_7320);
or U8125 (N_8125,N_7327,N_6627);
nor U8126 (N_8126,N_7267,N_7740);
or U8127 (N_8127,N_7230,N_6901);
nand U8128 (N_8128,N_6768,N_6560);
nor U8129 (N_8129,N_7707,N_7270);
nand U8130 (N_8130,N_7846,N_7988);
and U8131 (N_8131,N_6234,N_6301);
nor U8132 (N_8132,N_7659,N_6527);
nand U8133 (N_8133,N_7191,N_6298);
nand U8134 (N_8134,N_7231,N_7249);
and U8135 (N_8135,N_6609,N_7415);
or U8136 (N_8136,N_7640,N_7589);
xor U8137 (N_8137,N_7472,N_7932);
nand U8138 (N_8138,N_7989,N_7629);
xnor U8139 (N_8139,N_7608,N_7077);
and U8140 (N_8140,N_7264,N_7105);
nand U8141 (N_8141,N_7804,N_7269);
xnor U8142 (N_8142,N_6832,N_7964);
or U8143 (N_8143,N_6800,N_6413);
xnor U8144 (N_8144,N_6803,N_6092);
or U8145 (N_8145,N_6423,N_7111);
nor U8146 (N_8146,N_6099,N_7143);
xnor U8147 (N_8147,N_7262,N_7821);
and U8148 (N_8148,N_7818,N_6711);
and U8149 (N_8149,N_6709,N_6186);
nor U8150 (N_8150,N_6449,N_7186);
and U8151 (N_8151,N_7618,N_6245);
and U8152 (N_8152,N_6000,N_7813);
nor U8153 (N_8153,N_6373,N_6477);
nand U8154 (N_8154,N_6821,N_6653);
or U8155 (N_8155,N_7541,N_7967);
xnor U8156 (N_8156,N_7780,N_7198);
or U8157 (N_8157,N_6470,N_7765);
or U8158 (N_8158,N_7056,N_6401);
nand U8159 (N_8159,N_6638,N_6327);
and U8160 (N_8160,N_6141,N_6055);
nand U8161 (N_8161,N_6322,N_6037);
nand U8162 (N_8162,N_6244,N_6720);
nor U8163 (N_8163,N_7329,N_6208);
xor U8164 (N_8164,N_6446,N_6094);
or U8165 (N_8165,N_6073,N_7613);
and U8166 (N_8166,N_7350,N_6166);
nand U8167 (N_8167,N_6458,N_7302);
nand U8168 (N_8168,N_7985,N_6991);
xnor U8169 (N_8169,N_7152,N_7245);
nor U8170 (N_8170,N_7790,N_7987);
nor U8171 (N_8171,N_6180,N_7384);
nand U8172 (N_8172,N_6987,N_6580);
and U8173 (N_8173,N_6274,N_6015);
and U8174 (N_8174,N_7777,N_7014);
nand U8175 (N_8175,N_7805,N_7760);
nand U8176 (N_8176,N_7147,N_6881);
nor U8177 (N_8177,N_6363,N_7060);
xnor U8178 (N_8178,N_6308,N_6411);
nand U8179 (N_8179,N_6396,N_6972);
and U8180 (N_8180,N_6669,N_7265);
nor U8181 (N_8181,N_7710,N_7260);
or U8182 (N_8182,N_6614,N_7737);
nand U8183 (N_8183,N_6238,N_6950);
xnor U8184 (N_8184,N_7520,N_7724);
nand U8185 (N_8185,N_7970,N_6989);
nand U8186 (N_8186,N_6853,N_6805);
nand U8187 (N_8187,N_7976,N_6602);
or U8188 (N_8188,N_6061,N_6754);
and U8189 (N_8189,N_7650,N_6865);
nor U8190 (N_8190,N_7927,N_6271);
nand U8191 (N_8191,N_6321,N_6995);
nand U8192 (N_8192,N_7135,N_6316);
and U8193 (N_8193,N_6508,N_7825);
nor U8194 (N_8194,N_6198,N_7678);
and U8195 (N_8195,N_7310,N_7459);
and U8196 (N_8196,N_7530,N_6160);
nor U8197 (N_8197,N_7437,N_7190);
nor U8198 (N_8198,N_7571,N_6079);
or U8199 (N_8199,N_6632,N_6979);
nor U8200 (N_8200,N_6605,N_6749);
and U8201 (N_8201,N_6118,N_7901);
nor U8202 (N_8202,N_7447,N_7735);
and U8203 (N_8203,N_6574,N_6953);
nand U8204 (N_8204,N_6156,N_7903);
nand U8205 (N_8205,N_6075,N_7696);
or U8206 (N_8206,N_6767,N_6276);
nor U8207 (N_8207,N_6349,N_7324);
nand U8208 (N_8208,N_6691,N_7099);
and U8209 (N_8209,N_7500,N_6163);
nor U8210 (N_8210,N_7747,N_6999);
nand U8211 (N_8211,N_6666,N_6945);
xnor U8212 (N_8212,N_7061,N_6288);
xnor U8213 (N_8213,N_7252,N_7334);
and U8214 (N_8214,N_6200,N_6147);
nand U8215 (N_8215,N_7725,N_6937);
and U8216 (N_8216,N_7353,N_7219);
or U8217 (N_8217,N_7690,N_7057);
and U8218 (N_8218,N_6318,N_6811);
xnor U8219 (N_8219,N_7383,N_6142);
nand U8220 (N_8220,N_6440,N_6181);
nor U8221 (N_8221,N_7165,N_6012);
nand U8222 (N_8222,N_7212,N_7525);
xor U8223 (N_8223,N_7489,N_7655);
or U8224 (N_8224,N_6391,N_6228);
nor U8225 (N_8225,N_6703,N_6714);
or U8226 (N_8226,N_7451,N_6064);
xor U8227 (N_8227,N_6441,N_6455);
nand U8228 (N_8228,N_6513,N_6820);
or U8229 (N_8229,N_6468,N_7564);
nor U8230 (N_8230,N_6385,N_7749);
and U8231 (N_8231,N_7162,N_7476);
xnor U8232 (N_8232,N_6946,N_7416);
nand U8233 (N_8233,N_6510,N_7044);
nand U8234 (N_8234,N_6948,N_7318);
and U8235 (N_8235,N_6443,N_6320);
nor U8236 (N_8236,N_6409,N_6444);
or U8237 (N_8237,N_7524,N_6541);
xor U8238 (N_8238,N_7691,N_7870);
and U8239 (N_8239,N_7528,N_6695);
or U8240 (N_8240,N_6211,N_6520);
nand U8241 (N_8241,N_6606,N_7012);
xor U8242 (N_8242,N_7053,N_6375);
xor U8243 (N_8243,N_6159,N_7609);
nand U8244 (N_8244,N_6342,N_7960);
nor U8245 (N_8245,N_7812,N_6448);
nand U8246 (N_8246,N_7241,N_7411);
nand U8247 (N_8247,N_7468,N_7663);
xnor U8248 (N_8248,N_7362,N_7345);
and U8249 (N_8249,N_6255,N_7856);
nor U8250 (N_8250,N_6563,N_7251);
nor U8251 (N_8251,N_6553,N_7828);
nand U8252 (N_8252,N_7136,N_7718);
nor U8253 (N_8253,N_7313,N_6639);
nand U8254 (N_8254,N_6332,N_6133);
or U8255 (N_8255,N_6819,N_6601);
nand U8256 (N_8256,N_7692,N_7752);
and U8257 (N_8257,N_7535,N_7413);
nor U8258 (N_8258,N_7214,N_7034);
nand U8259 (N_8259,N_7154,N_7565);
nor U8260 (N_8260,N_7826,N_6374);
nor U8261 (N_8261,N_7047,N_7389);
xnor U8262 (N_8262,N_7806,N_7042);
and U8263 (N_8263,N_7599,N_6257);
xor U8264 (N_8264,N_6239,N_7715);
nand U8265 (N_8265,N_7457,N_6765);
or U8266 (N_8266,N_7868,N_7630);
nand U8267 (N_8267,N_7554,N_7414);
or U8268 (N_8268,N_6418,N_6898);
and U8269 (N_8269,N_7873,N_6108);
nand U8270 (N_8270,N_7914,N_7140);
xnor U8271 (N_8271,N_7355,N_7075);
and U8272 (N_8272,N_7092,N_7934);
nor U8273 (N_8273,N_7947,N_7978);
and U8274 (N_8274,N_7394,N_7453);
and U8275 (N_8275,N_7926,N_7877);
xor U8276 (N_8276,N_7084,N_7126);
nand U8277 (N_8277,N_7729,N_7065);
nand U8278 (N_8278,N_7367,N_6158);
and U8279 (N_8279,N_6528,N_6042);
xor U8280 (N_8280,N_7281,N_6975);
xor U8281 (N_8281,N_7180,N_7824);
xnor U8282 (N_8282,N_6493,N_6969);
nor U8283 (N_8283,N_6357,N_6031);
nand U8284 (N_8284,N_6090,N_6807);
nor U8285 (N_8285,N_6076,N_6600);
or U8286 (N_8286,N_7323,N_6543);
nor U8287 (N_8287,N_7938,N_7455);
xnor U8288 (N_8288,N_6066,N_6958);
and U8289 (N_8289,N_6779,N_6047);
and U8290 (N_8290,N_7247,N_6758);
and U8291 (N_8291,N_7073,N_7576);
or U8292 (N_8292,N_6708,N_7783);
nand U8293 (N_8293,N_6029,N_6573);
and U8294 (N_8294,N_7232,N_6532);
xnor U8295 (N_8295,N_6860,N_7894);
or U8296 (N_8296,N_6100,N_7712);
xnor U8297 (N_8297,N_7612,N_6472);
nand U8298 (N_8298,N_6850,N_7587);
nand U8299 (N_8299,N_7843,N_7036);
and U8300 (N_8300,N_7943,N_6517);
nand U8301 (N_8301,N_6206,N_7054);
xnor U8302 (N_8302,N_7660,N_6984);
and U8303 (N_8303,N_6334,N_6673);
nand U8304 (N_8304,N_7611,N_6362);
nor U8305 (N_8305,N_6814,N_7714);
or U8306 (N_8306,N_7562,N_7361);
and U8307 (N_8307,N_6584,N_7592);
nor U8308 (N_8308,N_6731,N_7142);
nand U8309 (N_8309,N_6962,N_7979);
and U8310 (N_8310,N_6259,N_7200);
nand U8311 (N_8311,N_7235,N_6599);
or U8312 (N_8312,N_7161,N_7001);
and U8313 (N_8313,N_7059,N_6336);
nor U8314 (N_8314,N_6161,N_7283);
and U8315 (N_8315,N_6397,N_6936);
nand U8316 (N_8316,N_7242,N_6876);
and U8317 (N_8317,N_6848,N_6102);
and U8318 (N_8318,N_7043,N_7201);
xnor U8319 (N_8319,N_7199,N_6595);
xnor U8320 (N_8320,N_7992,N_6942);
xor U8321 (N_8321,N_6624,N_7982);
nor U8322 (N_8322,N_6246,N_6547);
nor U8323 (N_8323,N_6944,N_6463);
xnor U8324 (N_8324,N_6529,N_7893);
xnor U8325 (N_8325,N_7454,N_7759);
and U8326 (N_8326,N_6247,N_6736);
nand U8327 (N_8327,N_7103,N_6124);
xnor U8328 (N_8328,N_7146,N_7481);
and U8329 (N_8329,N_7121,N_6346);
and U8330 (N_8330,N_7583,N_7138);
nand U8331 (N_8331,N_7237,N_6557);
xnor U8332 (N_8332,N_7531,N_7880);
nand U8333 (N_8333,N_7731,N_6616);
or U8334 (N_8334,N_6693,N_7965);
and U8335 (N_8335,N_7514,N_6738);
nand U8336 (N_8336,N_6127,N_6112);
xnor U8337 (N_8337,N_6537,N_6461);
nor U8338 (N_8338,N_7606,N_7347);
nand U8339 (N_8339,N_7924,N_6770);
xor U8340 (N_8340,N_6679,N_6561);
and U8341 (N_8341,N_7758,N_6262);
nand U8342 (N_8342,N_6777,N_6361);
or U8343 (N_8343,N_6149,N_7955);
xnor U8344 (N_8344,N_7072,N_7423);
and U8345 (N_8345,N_7920,N_7643);
and U8346 (N_8346,N_6677,N_6572);
or U8347 (N_8347,N_7645,N_6817);
or U8348 (N_8348,N_7642,N_7685);
nor U8349 (N_8349,N_6071,N_7284);
and U8350 (N_8350,N_7831,N_7533);
or U8351 (N_8351,N_6804,N_7827);
xnor U8352 (N_8352,N_6579,N_7717);
and U8353 (N_8353,N_6828,N_7025);
or U8354 (N_8354,N_6701,N_6466);
nor U8355 (N_8355,N_7131,N_7631);
nand U8356 (N_8356,N_6642,N_7835);
xnor U8357 (N_8357,N_7141,N_7446);
and U8358 (N_8358,N_6182,N_6210);
or U8359 (N_8359,N_7107,N_6852);
xor U8360 (N_8360,N_7603,N_7661);
or U8361 (N_8361,N_7787,N_7552);
or U8362 (N_8362,N_7498,N_6353);
nor U8363 (N_8363,N_7210,N_6660);
nor U8364 (N_8364,N_7348,N_7971);
or U8365 (N_8365,N_7445,N_6253);
xor U8366 (N_8366,N_6727,N_6039);
xor U8367 (N_8367,N_7052,N_7396);
or U8368 (N_8368,N_6407,N_6279);
nand U8369 (N_8369,N_7664,N_6284);
nand U8370 (N_8370,N_6207,N_6686);
and U8371 (N_8371,N_6717,N_6596);
xor U8372 (N_8372,N_7408,N_6364);
or U8373 (N_8373,N_6408,N_7442);
nand U8374 (N_8374,N_7887,N_6249);
and U8375 (N_8375,N_7933,N_7774);
xnor U8376 (N_8376,N_7584,N_6649);
xnor U8377 (N_8377,N_6663,N_7969);
nand U8378 (N_8378,N_7063,N_7879);
nor U8379 (N_8379,N_7365,N_7889);
and U8380 (N_8380,N_7022,N_6887);
and U8381 (N_8381,N_6416,N_7403);
nand U8382 (N_8382,N_6697,N_6292);
xor U8383 (N_8383,N_6546,N_6737);
or U8384 (N_8384,N_7918,N_6213);
and U8385 (N_8385,N_6475,N_6878);
or U8386 (N_8386,N_7658,N_6187);
or U8387 (N_8387,N_6990,N_6867);
and U8388 (N_8388,N_7523,N_6670);
and U8389 (N_8389,N_6035,N_7006);
and U8390 (N_8390,N_6864,N_6788);
nor U8391 (N_8391,N_6558,N_6780);
nand U8392 (N_8392,N_7322,N_7462);
nand U8393 (N_8393,N_6086,N_6725);
xor U8394 (N_8394,N_7399,N_7884);
and U8395 (N_8395,N_6330,N_7349);
nand U8396 (N_8396,N_6403,N_7109);
and U8397 (N_8397,N_6168,N_7503);
xor U8398 (N_8398,N_6219,N_6106);
nor U8399 (N_8399,N_7736,N_6753);
nand U8400 (N_8400,N_6268,N_6661);
or U8401 (N_8401,N_7296,N_6501);
or U8402 (N_8402,N_6806,N_6667);
and U8403 (N_8403,N_7174,N_6442);
nor U8404 (N_8404,N_7614,N_7751);
xnor U8405 (N_8405,N_6450,N_6145);
and U8406 (N_8406,N_6254,N_6426);
nor U8407 (N_8407,N_6746,N_7277);
and U8408 (N_8408,N_7534,N_6060);
nand U8409 (N_8409,N_6382,N_6706);
and U8410 (N_8410,N_7722,N_7474);
or U8411 (N_8411,N_7727,N_6741);
nand U8412 (N_8412,N_7360,N_6721);
xor U8413 (N_8413,N_7961,N_7866);
and U8414 (N_8414,N_6684,N_7286);
or U8415 (N_8415,N_6883,N_7159);
and U8416 (N_8416,N_6728,N_6307);
nand U8417 (N_8417,N_6760,N_7595);
or U8418 (N_8418,N_6956,N_7536);
xnor U8419 (N_8419,N_7285,N_7616);
and U8420 (N_8420,N_7292,N_7395);
xnor U8421 (N_8421,N_7838,N_6429);
xnor U8422 (N_8422,N_6184,N_6467);
xor U8423 (N_8423,N_6326,N_7194);
and U8424 (N_8424,N_6212,N_7907);
nand U8425 (N_8425,N_6179,N_7814);
nor U8426 (N_8426,N_6943,N_6103);
and U8427 (N_8427,N_6913,N_7719);
xor U8428 (N_8428,N_6251,N_6283);
or U8429 (N_8429,N_7461,N_6635);
and U8430 (N_8430,N_7460,N_6114);
nor U8431 (N_8431,N_7975,N_7380);
or U8432 (N_8432,N_6957,N_7545);
nor U8433 (N_8433,N_6772,N_6227);
or U8434 (N_8434,N_7702,N_6205);
and U8435 (N_8435,N_6433,N_6963);
and U8436 (N_8436,N_7465,N_7779);
nor U8437 (N_8437,N_7420,N_6452);
and U8438 (N_8438,N_6581,N_7953);
xor U8439 (N_8439,N_7641,N_6193);
nor U8440 (N_8440,N_7625,N_7484);
and U8441 (N_8441,N_7935,N_6915);
nor U8442 (N_8442,N_7703,N_7163);
and U8443 (N_8443,N_7486,N_6841);
xnor U8444 (N_8444,N_7864,N_6021);
nand U8445 (N_8445,N_7561,N_7325);
xor U8446 (N_8446,N_6365,N_6892);
xor U8447 (N_8447,N_6964,N_7351);
nor U8448 (N_8448,N_7836,N_7172);
and U8449 (N_8449,N_6136,N_7083);
xor U8450 (N_8450,N_7720,N_7013);
xnor U8451 (N_8451,N_7211,N_7952);
nor U8452 (N_8452,N_7910,N_7223);
and U8453 (N_8453,N_6976,N_7568);
or U8454 (N_8454,N_6132,N_6447);
or U8455 (N_8455,N_6038,N_6036);
nand U8456 (N_8456,N_7771,N_7929);
nand U8457 (N_8457,N_7745,N_6585);
or U8458 (N_8458,N_6836,N_6438);
or U8459 (N_8459,N_6926,N_6808);
nand U8460 (N_8460,N_6069,N_6016);
xor U8461 (N_8461,N_7221,N_6905);
nor U8462 (N_8462,N_6011,N_7999);
or U8463 (N_8463,N_6192,N_7106);
xor U8464 (N_8464,N_6104,N_6432);
nor U8465 (N_8465,N_6559,N_6313);
xnor U8466 (N_8466,N_7492,N_6516);
nand U8467 (N_8467,N_7830,N_6744);
xnor U8468 (N_8468,N_6387,N_7665);
and U8469 (N_8469,N_7761,N_6424);
nand U8470 (N_8470,N_7366,N_6694);
or U8471 (N_8471,N_6371,N_6017);
nor U8472 (N_8472,N_7607,N_7132);
nor U8473 (N_8473,N_7250,N_7509);
and U8474 (N_8474,N_7572,N_7139);
and U8475 (N_8475,N_7130,N_6109);
xnor U8476 (N_8476,N_7677,N_6538);
xnor U8477 (N_8477,N_7770,N_6459);
nor U8478 (N_8478,N_7031,N_6525);
nor U8479 (N_8479,N_6716,N_6033);
nand U8480 (N_8480,N_6465,N_7502);
or U8481 (N_8481,N_6608,N_6097);
and U8482 (N_8482,N_7434,N_6533);
xnor U8483 (N_8483,N_6985,N_7071);
nor U8484 (N_8484,N_6917,N_7002);
xor U8485 (N_8485,N_6378,N_6790);
xor U8486 (N_8486,N_6750,N_6462);
and U8487 (N_8487,N_6877,N_7786);
nor U8488 (N_8488,N_6439,N_6977);
xnor U8489 (N_8489,N_7195,N_6986);
and U8490 (N_8490,N_6290,N_7046);
nand U8491 (N_8491,N_7400,N_6840);
nand U8492 (N_8492,N_7145,N_6530);
and U8493 (N_8493,N_7372,N_7940);
xor U8494 (N_8494,N_7682,N_7398);
and U8495 (N_8495,N_7173,N_6291);
or U8496 (N_8496,N_7563,N_7508);
nor U8497 (N_8497,N_7738,N_7793);
or U8498 (N_8498,N_6226,N_7112);
or U8499 (N_8499,N_6778,N_6437);
or U8500 (N_8500,N_7449,N_6469);
or U8501 (N_8501,N_7473,N_7021);
nor U8502 (N_8502,N_6640,N_6802);
xnor U8503 (N_8503,N_7784,N_6194);
nand U8504 (N_8504,N_7343,N_7428);
nor U8505 (N_8505,N_6623,N_6296);
nor U8506 (N_8506,N_6394,N_7227);
xor U8507 (N_8507,N_7850,N_7419);
nand U8508 (N_8508,N_6089,N_7421);
xor U8509 (N_8509,N_7331,N_7913);
nand U8510 (N_8510,N_7491,N_7164);
nor U8511 (N_8511,N_7082,N_6914);
nand U8512 (N_8512,N_7872,N_6909);
and U8513 (N_8513,N_7518,N_7017);
and U8514 (N_8514,N_6063,N_7482);
nor U8515 (N_8515,N_7357,N_7944);
and U8516 (N_8516,N_7332,N_7257);
nand U8517 (N_8517,N_6932,N_7776);
xor U8518 (N_8518,N_7226,N_7091);
xor U8519 (N_8519,N_6384,N_6046);
xnor U8520 (N_8520,N_7090,N_6077);
nor U8521 (N_8521,N_7236,N_6997);
xnor U8522 (N_8522,N_6740,N_7433);
or U8523 (N_8523,N_6082,N_6855);
nand U8524 (N_8524,N_6875,N_7966);
and U8525 (N_8525,N_6070,N_6485);
nor U8526 (N_8526,N_6816,N_6847);
nand U8527 (N_8527,N_6360,N_6618);
xor U8528 (N_8528,N_7436,N_7763);
or U8529 (N_8529,N_7234,N_6941);
nand U8530 (N_8530,N_7591,N_6583);
nand U8531 (N_8531,N_7149,N_6849);
xnor U8532 (N_8532,N_7704,N_7859);
and U8533 (N_8533,N_6272,N_6043);
nand U8534 (N_8534,N_7791,N_7620);
or U8535 (N_8535,N_7216,N_6492);
nand U8536 (N_8536,N_7215,N_7410);
and U8537 (N_8537,N_6034,N_6366);
nand U8538 (N_8538,N_6218,N_7653);
and U8539 (N_8539,N_6565,N_7342);
nor U8540 (N_8540,N_7510,N_6065);
xnor U8541 (N_8541,N_7124,N_6988);
or U8542 (N_8542,N_7373,N_7405);
nand U8543 (N_8543,N_7928,N_7406);
xnor U8544 (N_8544,N_6083,N_6798);
and U8545 (N_8545,N_6499,N_6337);
nor U8546 (N_8546,N_7209,N_7213);
nor U8547 (N_8547,N_6791,N_7401);
xor U8548 (N_8548,N_7617,N_6269);
nand U8549 (N_8549,N_7679,N_6317);
nand U8550 (N_8550,N_7243,N_7921);
or U8551 (N_8551,N_7981,N_7954);
nand U8552 (N_8552,N_7429,N_6794);
nor U8553 (N_8553,N_6125,N_6464);
nand U8554 (N_8554,N_6729,N_6715);
or U8555 (N_8555,N_6542,N_6445);
nor U8556 (N_8556,N_6827,N_6351);
or U8557 (N_8557,N_6151,N_6518);
nand U8558 (N_8558,N_6339,N_7166);
nand U8559 (N_8559,N_6497,N_7597);
xor U8560 (N_8560,N_6123,N_6348);
xor U8561 (N_8561,N_6523,N_7379);
nor U8562 (N_8562,N_7956,N_7601);
nor U8563 (N_8563,N_6498,N_6863);
xnor U8564 (N_8564,N_7187,N_6938);
and U8565 (N_8565,N_6571,N_7621);
xor U8566 (N_8566,N_7892,N_6489);
xor U8567 (N_8567,N_6934,N_7882);
xnor U8568 (N_8568,N_6380,N_6911);
nor U8569 (N_8569,N_7346,N_6281);
nor U8570 (N_8570,N_7919,N_7193);
or U8571 (N_8571,N_7669,N_6949);
or U8572 (N_8572,N_7189,N_7110);
and U8573 (N_8573,N_7829,N_6224);
nand U8574 (N_8574,N_6275,N_6299);
xor U8575 (N_8575,N_7358,N_7282);
or U8576 (N_8576,N_7287,N_7438);
or U8577 (N_8577,N_6690,N_6395);
xor U8578 (N_8578,N_7950,N_7374);
nor U8579 (N_8579,N_7748,N_7431);
nor U8580 (N_8580,N_7713,N_7298);
nor U8581 (N_8581,N_7949,N_7116);
xnor U8582 (N_8582,N_6978,N_7593);
xor U8583 (N_8583,N_6095,N_7547);
xnor U8584 (N_8584,N_6502,N_7551);
nand U8585 (N_8585,N_6873,N_6354);
nor U8586 (N_8586,N_7317,N_7160);
and U8587 (N_8587,N_6897,N_6013);
nand U8588 (N_8588,N_7113,N_7390);
nand U8589 (N_8589,N_7815,N_7184);
and U8590 (N_8590,N_6908,N_7382);
or U8591 (N_8591,N_7951,N_6122);
xnor U8592 (N_8592,N_6933,N_7654);
xor U8593 (N_8593,N_6782,N_7811);
xor U8594 (N_8594,N_6110,N_6793);
xor U8595 (N_8595,N_7507,N_7023);
xor U8596 (N_8596,N_7917,N_7615);
nor U8597 (N_8597,N_7432,N_6594);
or U8598 (N_8598,N_6119,N_7513);
nand U8599 (N_8599,N_6243,N_6707);
xor U8600 (N_8600,N_6338,N_7010);
nor U8601 (N_8601,N_7028,N_7624);
and U8602 (N_8602,N_7798,N_7801);
xnor U8603 (N_8603,N_7377,N_7652);
nor U8604 (N_8604,N_6356,N_6164);
xor U8605 (N_8605,N_6597,N_7573);
and U8606 (N_8606,N_6087,N_7834);
nand U8607 (N_8607,N_6512,N_6372);
nand U8608 (N_8608,N_7123,N_6648);
and U8609 (N_8609,N_6896,N_6005);
nand U8610 (N_8610,N_7557,N_7170);
xnor U8611 (N_8611,N_6289,N_7656);
nor U8612 (N_8612,N_7011,N_7048);
or U8613 (N_8613,N_6884,N_6858);
xor U8614 (N_8614,N_7820,N_6787);
nand U8615 (N_8615,N_7254,N_6834);
nand U8616 (N_8616,N_6126,N_6004);
or U8617 (N_8617,N_7925,N_7266);
and U8618 (N_8618,N_7328,N_7680);
and U8619 (N_8619,N_7086,N_7381);
and U8620 (N_8620,N_7844,N_6761);
or U8621 (N_8621,N_6422,N_7833);
nand U8622 (N_8622,N_7537,N_7479);
or U8623 (N_8623,N_6456,N_6190);
nand U8624 (N_8624,N_7030,N_7202);
or U8625 (N_8625,N_7993,N_7667);
and U8626 (N_8626,N_6496,N_7908);
nand U8627 (N_8627,N_7407,N_7769);
nand U8628 (N_8628,N_6699,N_6612);
nor U8629 (N_8629,N_7144,N_7045);
or U8630 (N_8630,N_6566,N_7973);
and U8631 (N_8631,N_7634,N_6237);
or U8632 (N_8632,N_7319,N_7467);
nor U8633 (N_8633,N_6370,N_7579);
nand U8634 (N_8634,N_6067,N_6049);
nand U8635 (N_8635,N_6603,N_6900);
nor U8636 (N_8636,N_7582,N_6027);
nor U8637 (N_8637,N_6325,N_7529);
and U8638 (N_8638,N_6153,N_7878);
nand U8639 (N_8639,N_7773,N_6692);
nand U8640 (N_8640,N_6974,N_6923);
and U8641 (N_8641,N_7385,N_6586);
nor U8642 (N_8642,N_6024,N_7026);
or U8643 (N_8643,N_7852,N_7314);
and U8644 (N_8644,N_7633,N_6519);
and U8645 (N_8645,N_7253,N_6607);
xor U8646 (N_8646,N_7902,N_7794);
nor U8647 (N_8647,N_6453,N_7225);
nand U8648 (N_8648,N_7466,N_6924);
nand U8649 (N_8649,N_7295,N_7095);
xor U8650 (N_8650,N_6859,N_7566);
or U8651 (N_8651,N_6494,N_6762);
and U8652 (N_8652,N_7785,N_7371);
or U8653 (N_8653,N_7050,N_6368);
nand U8654 (N_8654,N_7553,N_7064);
and U8655 (N_8655,N_6622,N_6615);
or U8656 (N_8656,N_6148,N_7673);
nand U8657 (N_8657,N_7085,N_7464);
xor U8658 (N_8658,N_7550,N_7542);
or U8659 (N_8659,N_7364,N_7148);
or U8660 (N_8660,N_6971,N_6052);
or U8661 (N_8661,N_6885,N_6476);
xnor U8662 (N_8662,N_7842,N_7504);
and U8663 (N_8663,N_7671,N_7016);
or U8664 (N_8664,N_6774,N_7168);
nor U8665 (N_8665,N_7009,N_6678);
nand U8666 (N_8666,N_6146,N_7271);
nand U8667 (N_8667,N_6484,N_6734);
and U8668 (N_8668,N_7800,N_6732);
or U8669 (N_8669,N_7764,N_7336);
or U8670 (N_8670,N_7338,N_6549);
nand U8671 (N_8671,N_6633,N_7114);
xnor U8672 (N_8672,N_6028,N_7255);
or U8673 (N_8673,N_6018,N_7488);
xor U8674 (N_8674,N_7483,N_7899);
xor U8675 (N_8675,N_6764,N_6947);
and U8676 (N_8676,N_7559,N_7217);
nand U8677 (N_8677,N_7792,N_6098);
and U8678 (N_8678,N_6872,N_7196);
and U8679 (N_8679,N_7294,N_7726);
nand U8680 (N_8680,N_7356,N_7548);
nand U8681 (N_8681,N_7004,N_7274);
and U8682 (N_8682,N_7822,N_6526);
and U8683 (N_8683,N_7478,N_6524);
nand U8684 (N_8684,N_6672,N_7104);
nand U8685 (N_8685,N_6137,N_6637);
or U8686 (N_8686,N_7151,N_6818);
nor U8687 (N_8687,N_6451,N_6120);
and U8688 (N_8688,N_7038,N_7670);
xor U8689 (N_8689,N_7088,N_7743);
and U8690 (N_8690,N_7746,N_7694);
and U8691 (N_8691,N_6304,N_7699);
nor U8692 (N_8692,N_7206,N_7102);
or U8693 (N_8693,N_6540,N_7684);
nand U8694 (N_8694,N_7501,N_6482);
and U8695 (N_8695,N_7378,N_7303);
nor U8696 (N_8696,N_6970,N_6412);
nand U8697 (N_8697,N_6105,N_7066);
nand U8698 (N_8698,N_6019,N_6981);
or U8699 (N_8699,N_6072,N_7404);
or U8700 (N_8700,N_6959,N_7851);
or U8701 (N_8701,N_6792,N_6488);
xor U8702 (N_8702,N_6920,N_6645);
xor U8703 (N_8703,N_7916,N_7862);
nand U8704 (N_8704,N_6824,N_6260);
nor U8705 (N_8705,N_7876,N_7538);
and U8706 (N_8706,N_7915,N_6265);
nand U8707 (N_8707,N_6040,N_6335);
or U8708 (N_8708,N_6775,N_7977);
nand U8709 (N_8709,N_6203,N_6838);
or U8710 (N_8710,N_6022,N_7556);
or U8711 (N_8711,N_6280,N_6231);
xnor U8712 (N_8712,N_7397,N_6062);
xnor U8713 (N_8713,N_7622,N_7158);
and U8714 (N_8714,N_6252,N_6935);
nand U8715 (N_8715,N_7516,N_7359);
nor U8716 (N_8716,N_6893,N_6555);
xnor U8717 (N_8717,N_6115,N_7635);
nor U8718 (N_8718,N_6544,N_7604);
and U8719 (N_8719,N_6116,N_6874);
or U8720 (N_8720,N_7019,N_7450);
nand U8721 (N_8721,N_6285,N_6214);
and U8722 (N_8722,N_6204,N_7683);
xor U8723 (N_8723,N_7854,N_6845);
xor U8724 (N_8724,N_7594,N_6358);
and U8725 (N_8725,N_7522,N_7305);
nor U8726 (N_8726,N_6405,N_7544);
nor U8727 (N_8727,N_6675,N_6454);
nor U8728 (N_8728,N_7179,N_6980);
xnor U8729 (N_8729,N_6196,N_6665);
nand U8730 (N_8730,N_7674,N_6002);
nand U8731 (N_8731,N_6751,N_7990);
nor U8732 (N_8732,N_6305,N_7558);
and U8733 (N_8733,N_6588,N_7192);
or U8734 (N_8734,N_7788,N_6535);
and U8735 (N_8735,N_7681,N_7797);
and U8736 (N_8736,N_7883,N_7258);
and U8737 (N_8737,N_6295,N_6483);
nor U8738 (N_8738,N_6879,N_7602);
or U8739 (N_8739,N_6264,N_7968);
and U8740 (N_8740,N_7119,N_6562);
xor U8741 (N_8741,N_6236,N_6084);
nor U8742 (N_8742,N_7874,N_6652);
or U8743 (N_8743,N_7698,N_7923);
xor U8744 (N_8744,N_7906,N_7721);
nand U8745 (N_8745,N_7496,N_7845);
and U8746 (N_8746,N_7858,N_6300);
xnor U8747 (N_8747,N_7708,N_7991);
xor U8748 (N_8748,N_7307,N_7008);
xnor U8749 (N_8749,N_7705,N_6229);
and U8750 (N_8750,N_7772,N_6143);
or U8751 (N_8751,N_6303,N_7244);
nor U8752 (N_8752,N_6173,N_6628);
nand U8753 (N_8753,N_7912,N_7337);
or U8754 (N_8754,N_6503,N_6490);
xor U8755 (N_8755,N_6404,N_7439);
nand U8756 (N_8756,N_7427,N_6656);
xnor U8757 (N_8757,N_6014,N_7733);
or U8758 (N_8758,N_6869,N_6001);
and U8759 (N_8759,N_6996,N_6713);
nor U8760 (N_8760,N_6576,N_7560);
nand U8761 (N_8761,N_7628,N_6009);
nand U8762 (N_8762,N_6188,N_7352);
or U8763 (N_8763,N_6719,N_6217);
nor U8764 (N_8764,N_7581,N_6880);
nand U8765 (N_8765,N_7494,N_6393);
or U8766 (N_8766,N_6171,N_7129);
and U8767 (N_8767,N_6505,N_7128);
and U8768 (N_8768,N_7865,N_6733);
nand U8769 (N_8769,N_6722,N_6724);
and U8770 (N_8770,N_7580,N_7368);
and U8771 (N_8771,N_6702,N_6225);
nand U8772 (N_8772,N_7841,N_7853);
xor U8773 (N_8773,N_6209,N_7363);
and U8774 (N_8774,N_6053,N_6831);
xnor U8775 (N_8775,N_6427,N_7517);
nand U8776 (N_8776,N_7176,N_6421);
xnor U8777 (N_8777,N_6548,N_7632);
nand U8778 (N_8778,N_6197,N_7040);
and U8779 (N_8779,N_6329,N_7711);
nor U8780 (N_8780,N_7150,N_6169);
nor U8781 (N_8781,N_7018,N_6435);
nor U8782 (N_8782,N_7959,N_7623);
nand U8783 (N_8783,N_6861,N_6682);
xnor U8784 (N_8784,N_6051,N_6081);
nor U8785 (N_8785,N_7387,N_6154);
or U8786 (N_8786,N_6668,N_7768);
nor U8787 (N_8787,N_6743,N_7755);
nand U8788 (N_8788,N_7100,N_7074);
or U8789 (N_8789,N_6522,N_6930);
nand U8790 (N_8790,N_6068,N_6982);
or U8791 (N_8791,N_7799,N_7279);
or U8792 (N_8792,N_6056,N_6965);
xnor U8793 (N_8793,N_6823,N_6998);
and U8794 (N_8794,N_6735,N_6592);
nor U8795 (N_8795,N_7024,N_7972);
and U8796 (N_8796,N_7505,N_7888);
nand U8797 (N_8797,N_7306,N_6610);
or U8798 (N_8798,N_7598,N_6152);
xor U8799 (N_8799,N_6536,N_6189);
nor U8800 (N_8800,N_7832,N_6175);
xnor U8801 (N_8801,N_7700,N_6689);
nand U8802 (N_8802,N_6796,N_7945);
or U8803 (N_8803,N_6676,N_6129);
nor U8804 (N_8804,N_6657,N_6398);
nor U8805 (N_8805,N_6907,N_6425);
xor U8806 (N_8806,N_6748,N_7511);
nand U8807 (N_8807,N_7796,N_7133);
nand U8808 (N_8808,N_7756,N_6431);
or U8809 (N_8809,N_7268,N_7651);
xnor U8810 (N_8810,N_7321,N_6700);
and U8811 (N_8811,N_6376,N_7344);
or U8812 (N_8812,N_6726,N_7081);
nand U8813 (N_8813,N_7840,N_7493);
nand U8814 (N_8814,N_7316,N_6263);
or U8815 (N_8815,N_6955,N_7452);
nand U8816 (N_8816,N_7986,N_7701);
nor U8817 (N_8817,N_6306,N_7068);
nand U8818 (N_8818,N_7033,N_7003);
nand U8819 (N_8819,N_6888,N_7291);
and U8820 (N_8820,N_7686,N_7181);
and U8821 (N_8821,N_6854,N_6813);
nand U8822 (N_8822,N_6531,N_6587);
xor U8823 (N_8823,N_6328,N_6010);
xnor U8824 (N_8824,N_7067,N_7007);
or U8825 (N_8825,N_6223,N_6591);
xor U8826 (N_8826,N_7816,N_7456);
or U8827 (N_8827,N_6742,N_7885);
xnor U8828 (N_8828,N_6460,N_6319);
nand U8829 (N_8829,N_7512,N_7029);
nand U8830 (N_8830,N_7543,N_7304);
nor U8831 (N_8831,N_6842,N_7203);
nand U8832 (N_8832,N_6939,N_7983);
and U8833 (N_8833,N_7259,N_6221);
xnor U8834 (N_8834,N_6621,N_7341);
nor U8835 (N_8835,N_7475,N_6428);
xor U8836 (N_8836,N_7574,N_7646);
nor U8837 (N_8837,N_7807,N_7855);
nand U8838 (N_8838,N_7881,N_7049);
or U8839 (N_8839,N_6912,N_7222);
xor U8840 (N_8840,N_7706,N_6278);
xor U8841 (N_8841,N_6904,N_7080);
and U8842 (N_8842,N_7931,N_6085);
nor U8843 (N_8843,N_6822,N_7897);
nand U8844 (N_8844,N_6685,N_7402);
nand U8845 (N_8845,N_7239,N_6191);
or U8846 (N_8846,N_6617,N_7886);
nor U8847 (N_8847,N_6157,N_6688);
and U8848 (N_8848,N_7532,N_7375);
nand U8849 (N_8849,N_6593,N_6511);
or U8850 (N_8850,N_7477,N_7648);
and U8851 (N_8851,N_6619,N_6902);
and U8852 (N_8852,N_7734,N_6647);
xnor U8853 (N_8853,N_6659,N_7896);
nand U8854 (N_8854,N_6569,N_7930);
nor U8855 (N_8855,N_6705,N_7185);
or U8856 (N_8856,N_6514,N_7315);
xnor U8857 (N_8857,N_6131,N_6155);
nand U8858 (N_8858,N_7781,N_7137);
xnor U8859 (N_8859,N_7055,N_6177);
and U8860 (N_8860,N_6966,N_7848);
xor U8861 (N_8861,N_6250,N_7957);
or U8862 (N_8862,N_7898,N_7020);
and U8863 (N_8863,N_6739,N_6582);
or U8864 (N_8864,N_7480,N_7280);
or U8865 (N_8865,N_7936,N_6951);
or U8866 (N_8866,N_6406,N_6242);
nand U8867 (N_8867,N_6093,N_6222);
nand U8868 (N_8868,N_6759,N_6419);
nor U8869 (N_8869,N_6929,N_7122);
or U8870 (N_8870,N_6921,N_7984);
xor U8871 (N_8871,N_7463,N_7689);
nor U8872 (N_8872,N_6025,N_7087);
nor U8873 (N_8873,N_7600,N_7742);
nand U8874 (N_8874,N_7426,N_6940);
or U8875 (N_8875,N_7693,N_6007);
xor U8876 (N_8876,N_7802,N_6826);
nand U8877 (N_8877,N_7809,N_6752);
xor U8878 (N_8878,N_7939,N_6745);
or U8879 (N_8879,N_6776,N_6545);
nand U8880 (N_8880,N_7089,N_6057);
nand U8881 (N_8881,N_6054,N_7273);
xor U8882 (N_8882,N_7904,N_7312);
and U8883 (N_8883,N_6347,N_6241);
nor U8884 (N_8884,N_6185,N_6664);
nor U8885 (N_8885,N_6121,N_7946);
or U8886 (N_8886,N_7803,N_7330);
nand U8887 (N_8887,N_7224,N_6556);
nand U8888 (N_8888,N_6050,N_6130);
nand U8889 (N_8889,N_6113,N_6323);
xor U8890 (N_8890,N_6613,N_6379);
nor U8891 (N_8891,N_6578,N_7078);
nand U8892 (N_8892,N_6644,N_7308);
xor U8893 (N_8893,N_7817,N_6590);
nor U8894 (N_8894,N_7278,N_6150);
xnor U8895 (N_8895,N_6786,N_6781);
nand U8896 (N_8896,N_7994,N_6680);
nand U8897 (N_8897,N_7256,N_7300);
nand U8898 (N_8898,N_7120,N_7695);
xor U8899 (N_8899,N_6712,N_7741);
or U8900 (N_8900,N_7605,N_6400);
xnor U8901 (N_8901,N_6631,N_6430);
xor U8902 (N_8902,N_6381,N_7723);
or U8903 (N_8903,N_6134,N_7672);
xnor U8904 (N_8904,N_7857,N_7922);
and U8905 (N_8905,N_6967,N_7470);
xor U8906 (N_8906,N_7578,N_6862);
or U8907 (N_8907,N_6857,N_7980);
or U8908 (N_8908,N_6992,N_6473);
or U8909 (N_8909,N_7335,N_6080);
and U8910 (N_8910,N_7626,N_7911);
or U8911 (N_8911,N_6350,N_7941);
nand U8912 (N_8912,N_7861,N_6833);
and U8913 (N_8913,N_6233,N_6747);
and U8914 (N_8914,N_7005,N_6773);
or U8915 (N_8915,N_6481,N_7058);
and U8916 (N_8916,N_6789,N_6478);
and U8917 (N_8917,N_7839,N_7757);
xnor U8918 (N_8918,N_7871,N_7412);
xnor U8919 (N_8919,N_7668,N_7619);
or U8920 (N_8920,N_6534,N_7238);
nand U8921 (N_8921,N_6830,N_6474);
and U8922 (N_8922,N_6344,N_6176);
or U8923 (N_8923,N_6550,N_6266);
nor U8924 (N_8924,N_7962,N_6687);
and U8925 (N_8925,N_6471,N_6341);
xor U8926 (N_8926,N_6377,N_6783);
xnor U8927 (N_8927,N_6101,N_6809);
nor U8928 (N_8928,N_6567,N_6058);
nor U8929 (N_8929,N_7762,N_6718);
nand U8930 (N_8930,N_7079,N_7657);
xor U8931 (N_8931,N_7094,N_6886);
nand U8932 (N_8932,N_7627,N_6107);
nand U8933 (N_8933,N_6899,N_7709);
nor U8934 (N_8934,N_7183,N_7177);
or U8935 (N_8935,N_7895,N_7471);
nor U8936 (N_8936,N_6810,N_6261);
nand U8937 (N_8937,N_6165,N_7860);
and U8938 (N_8938,N_6507,N_7290);
nor U8939 (N_8939,N_6604,N_7156);
nand U8940 (N_8940,N_6928,N_7218);
nand U8941 (N_8941,N_6128,N_6331);
nor U8942 (N_8942,N_7032,N_6890);
and U8943 (N_8943,N_6795,N_6023);
and U8944 (N_8944,N_6620,N_7069);
and U8945 (N_8945,N_6162,N_6655);
and U8946 (N_8946,N_7205,N_6889);
xnor U8947 (N_8947,N_6270,N_6757);
nor U8948 (N_8948,N_6683,N_7435);
and U8949 (N_8949,N_7675,N_6399);
xor U8950 (N_8950,N_7240,N_7869);
xnor U8951 (N_8951,N_7035,N_6026);
xor U8952 (N_8952,N_6230,N_6287);
nor U8953 (N_8953,N_6386,N_6324);
nor U8954 (N_8954,N_7998,N_7037);
nor U8955 (N_8955,N_6551,N_6383);
xnor U8956 (N_8956,N_7539,N_7823);
and U8957 (N_8957,N_6634,N_7527);
nand U8958 (N_8958,N_7228,N_7117);
or U8959 (N_8959,N_6785,N_6392);
or U8960 (N_8960,N_6837,N_7076);
nor U8961 (N_8961,N_7301,N_6235);
or U8962 (N_8962,N_7890,N_7577);
nor U8963 (N_8963,N_7229,N_6868);
xnor U8964 (N_8964,N_6894,N_6277);
xor U8965 (N_8965,N_6654,N_6140);
or U8966 (N_8966,N_7485,N_6730);
and U8967 (N_8967,N_6755,N_6170);
xor U8968 (N_8968,N_6829,N_6388);
xor U8969 (N_8969,N_6954,N_7393);
or U8970 (N_8970,N_6797,N_6302);
or U8971 (N_8971,N_6315,N_7937);
and U8972 (N_8972,N_7638,N_6625);
nand U8973 (N_8973,N_7157,N_6799);
or U8974 (N_8974,N_6144,N_6480);
nand U8975 (N_8975,N_6598,N_6410);
or U8976 (N_8976,N_6771,N_6479);
and U8977 (N_8977,N_7905,N_7540);
nand U8978 (N_8978,N_6993,N_6309);
nor U8979 (N_8979,N_7167,N_6784);
xor U8980 (N_8980,N_6020,N_7687);
or U8981 (N_8981,N_7837,N_6681);
and U8982 (N_8982,N_7197,N_7782);
nor U8983 (N_8983,N_7127,N_7469);
nor U8984 (N_8984,N_6044,N_6825);
nand U8985 (N_8985,N_7688,N_6570);
or U8986 (N_8986,N_7115,N_6568);
nand U8987 (N_8987,N_7909,N_7388);
or U8988 (N_8988,N_7101,N_7867);
and U8989 (N_8989,N_6199,N_7487);
xnor U8990 (N_8990,N_7549,N_7153);
nand U8991 (N_8991,N_7118,N_6340);
or U8992 (N_8992,N_7644,N_7744);
nor U8993 (N_8993,N_6651,N_6968);
nand U8994 (N_8994,N_6646,N_6355);
or U8995 (N_8995,N_7175,N_7891);
nor U8996 (N_8996,N_7272,N_7730);
nor U8997 (N_8997,N_6267,N_6074);
xor U8998 (N_8998,N_7499,N_6552);
xor U8999 (N_8999,N_6041,N_7767);
or U9000 (N_9000,N_7847,N_6178);
nor U9001 (N_9001,N_7479,N_7399);
xor U9002 (N_9002,N_7849,N_6918);
nand U9003 (N_9003,N_7902,N_6628);
nand U9004 (N_9004,N_7808,N_7286);
xnor U9005 (N_9005,N_6643,N_7401);
or U9006 (N_9006,N_7251,N_6163);
xor U9007 (N_9007,N_7504,N_6957);
xnor U9008 (N_9008,N_6394,N_6796);
xor U9009 (N_9009,N_6060,N_7004);
nor U9010 (N_9010,N_7521,N_6625);
nand U9011 (N_9011,N_7990,N_7460);
or U9012 (N_9012,N_6591,N_7813);
nand U9013 (N_9013,N_6138,N_7644);
xnor U9014 (N_9014,N_7366,N_7537);
or U9015 (N_9015,N_7162,N_7572);
or U9016 (N_9016,N_7317,N_7580);
or U9017 (N_9017,N_7362,N_7411);
or U9018 (N_9018,N_7818,N_6797);
nand U9019 (N_9019,N_6792,N_6071);
xnor U9020 (N_9020,N_7641,N_7944);
nand U9021 (N_9021,N_6740,N_6168);
nor U9022 (N_9022,N_7195,N_7245);
or U9023 (N_9023,N_6976,N_7428);
nor U9024 (N_9024,N_7066,N_7126);
nand U9025 (N_9025,N_6826,N_7604);
nand U9026 (N_9026,N_7743,N_6522);
and U9027 (N_9027,N_6461,N_7226);
or U9028 (N_9028,N_6753,N_6636);
xnor U9029 (N_9029,N_6039,N_7701);
or U9030 (N_9030,N_7332,N_6064);
and U9031 (N_9031,N_7223,N_7081);
or U9032 (N_9032,N_7783,N_6197);
nor U9033 (N_9033,N_6997,N_7543);
nor U9034 (N_9034,N_7575,N_7762);
xnor U9035 (N_9035,N_6786,N_6427);
nor U9036 (N_9036,N_6777,N_6258);
and U9037 (N_9037,N_7749,N_7320);
nand U9038 (N_9038,N_7972,N_6607);
or U9039 (N_9039,N_6840,N_6964);
nand U9040 (N_9040,N_6694,N_7961);
nor U9041 (N_9041,N_7928,N_6241);
nor U9042 (N_9042,N_6330,N_6065);
xnor U9043 (N_9043,N_6488,N_6980);
and U9044 (N_9044,N_6780,N_6115);
or U9045 (N_9045,N_7453,N_6255);
xnor U9046 (N_9046,N_6081,N_7708);
or U9047 (N_9047,N_6124,N_6886);
nor U9048 (N_9048,N_6690,N_6997);
xor U9049 (N_9049,N_6756,N_6952);
and U9050 (N_9050,N_6705,N_7085);
nand U9051 (N_9051,N_6320,N_7597);
nand U9052 (N_9052,N_7465,N_7018);
xor U9053 (N_9053,N_6838,N_6554);
xnor U9054 (N_9054,N_7169,N_6553);
nor U9055 (N_9055,N_7485,N_7698);
and U9056 (N_9056,N_7994,N_6208);
nor U9057 (N_9057,N_6403,N_6584);
nor U9058 (N_9058,N_7015,N_6821);
nor U9059 (N_9059,N_7304,N_6570);
nand U9060 (N_9060,N_6394,N_7672);
xor U9061 (N_9061,N_6861,N_6705);
xor U9062 (N_9062,N_7845,N_6323);
nor U9063 (N_9063,N_7190,N_7441);
nor U9064 (N_9064,N_7236,N_7883);
nand U9065 (N_9065,N_7899,N_6674);
nor U9066 (N_9066,N_7692,N_6221);
and U9067 (N_9067,N_6117,N_6222);
nor U9068 (N_9068,N_6180,N_6265);
or U9069 (N_9069,N_7687,N_7034);
nor U9070 (N_9070,N_7549,N_6299);
nand U9071 (N_9071,N_7383,N_7250);
xnor U9072 (N_9072,N_6363,N_6535);
or U9073 (N_9073,N_6123,N_6037);
and U9074 (N_9074,N_6087,N_6274);
nor U9075 (N_9075,N_7097,N_7758);
nor U9076 (N_9076,N_7247,N_7938);
nor U9077 (N_9077,N_6402,N_6004);
nor U9078 (N_9078,N_7443,N_7081);
or U9079 (N_9079,N_7439,N_6226);
or U9080 (N_9080,N_7396,N_7172);
xnor U9081 (N_9081,N_7051,N_6498);
xnor U9082 (N_9082,N_6841,N_7354);
and U9083 (N_9083,N_7207,N_6312);
or U9084 (N_9084,N_7990,N_7388);
or U9085 (N_9085,N_7405,N_6326);
xnor U9086 (N_9086,N_6131,N_6729);
nor U9087 (N_9087,N_7818,N_6893);
nor U9088 (N_9088,N_6558,N_7005);
or U9089 (N_9089,N_6989,N_6269);
and U9090 (N_9090,N_6674,N_6388);
or U9091 (N_9091,N_6258,N_6676);
or U9092 (N_9092,N_6309,N_6779);
and U9093 (N_9093,N_7431,N_7150);
or U9094 (N_9094,N_6089,N_6035);
nand U9095 (N_9095,N_7983,N_6766);
nor U9096 (N_9096,N_7120,N_6134);
nand U9097 (N_9097,N_7320,N_6214);
nand U9098 (N_9098,N_6661,N_6353);
nand U9099 (N_9099,N_7989,N_7375);
and U9100 (N_9100,N_7010,N_7970);
nor U9101 (N_9101,N_6512,N_7558);
xor U9102 (N_9102,N_6774,N_7257);
and U9103 (N_9103,N_7511,N_6013);
nor U9104 (N_9104,N_7891,N_7004);
nor U9105 (N_9105,N_6821,N_6685);
and U9106 (N_9106,N_7170,N_7356);
xor U9107 (N_9107,N_7546,N_7957);
or U9108 (N_9108,N_6920,N_7306);
xnor U9109 (N_9109,N_7541,N_6169);
xor U9110 (N_9110,N_7386,N_6451);
and U9111 (N_9111,N_7478,N_7738);
nand U9112 (N_9112,N_7277,N_7436);
nand U9113 (N_9113,N_7992,N_6501);
and U9114 (N_9114,N_7219,N_7848);
nand U9115 (N_9115,N_7268,N_6703);
xnor U9116 (N_9116,N_6784,N_7624);
nand U9117 (N_9117,N_6161,N_7439);
or U9118 (N_9118,N_7227,N_7530);
nor U9119 (N_9119,N_7302,N_7057);
nor U9120 (N_9120,N_7499,N_7875);
xnor U9121 (N_9121,N_7965,N_6957);
nor U9122 (N_9122,N_6122,N_7433);
and U9123 (N_9123,N_7343,N_7306);
nand U9124 (N_9124,N_6740,N_6716);
nor U9125 (N_9125,N_6646,N_6305);
nand U9126 (N_9126,N_7344,N_7709);
nand U9127 (N_9127,N_7173,N_7121);
and U9128 (N_9128,N_6992,N_6381);
or U9129 (N_9129,N_6055,N_6201);
xor U9130 (N_9130,N_6077,N_6962);
xor U9131 (N_9131,N_6692,N_6853);
xor U9132 (N_9132,N_7208,N_7451);
or U9133 (N_9133,N_6988,N_7131);
xor U9134 (N_9134,N_6620,N_7074);
or U9135 (N_9135,N_6513,N_7344);
or U9136 (N_9136,N_7959,N_7452);
xnor U9137 (N_9137,N_7392,N_6129);
or U9138 (N_9138,N_6554,N_7586);
xnor U9139 (N_9139,N_6020,N_7625);
or U9140 (N_9140,N_6344,N_6925);
nand U9141 (N_9141,N_7117,N_6414);
nor U9142 (N_9142,N_7328,N_6910);
or U9143 (N_9143,N_7654,N_6662);
xor U9144 (N_9144,N_6057,N_7478);
nor U9145 (N_9145,N_6502,N_7201);
nand U9146 (N_9146,N_7135,N_7156);
nand U9147 (N_9147,N_6621,N_6685);
or U9148 (N_9148,N_6980,N_7323);
nor U9149 (N_9149,N_7675,N_6044);
or U9150 (N_9150,N_7323,N_6747);
or U9151 (N_9151,N_6663,N_6224);
nor U9152 (N_9152,N_6368,N_6893);
xor U9153 (N_9153,N_7129,N_6325);
or U9154 (N_9154,N_6865,N_7596);
xor U9155 (N_9155,N_6526,N_6821);
xnor U9156 (N_9156,N_7526,N_6627);
or U9157 (N_9157,N_6785,N_6305);
nand U9158 (N_9158,N_7358,N_7462);
or U9159 (N_9159,N_6137,N_7988);
xnor U9160 (N_9160,N_7019,N_7086);
nand U9161 (N_9161,N_6407,N_6840);
or U9162 (N_9162,N_7203,N_7779);
or U9163 (N_9163,N_6276,N_6770);
xnor U9164 (N_9164,N_6277,N_7101);
xnor U9165 (N_9165,N_6039,N_7462);
or U9166 (N_9166,N_6632,N_6676);
xor U9167 (N_9167,N_6516,N_7629);
xnor U9168 (N_9168,N_6889,N_6712);
xnor U9169 (N_9169,N_6288,N_7282);
nand U9170 (N_9170,N_6445,N_7203);
nand U9171 (N_9171,N_7804,N_6051);
nor U9172 (N_9172,N_7534,N_6652);
or U9173 (N_9173,N_7522,N_6912);
and U9174 (N_9174,N_7071,N_7689);
or U9175 (N_9175,N_6880,N_6413);
nand U9176 (N_9176,N_7511,N_6285);
and U9177 (N_9177,N_6902,N_6701);
xnor U9178 (N_9178,N_6601,N_7148);
xnor U9179 (N_9179,N_7128,N_7275);
nand U9180 (N_9180,N_7767,N_6969);
nand U9181 (N_9181,N_6331,N_7814);
xnor U9182 (N_9182,N_7845,N_7906);
nand U9183 (N_9183,N_6420,N_7612);
and U9184 (N_9184,N_6757,N_6402);
nand U9185 (N_9185,N_7146,N_6272);
nand U9186 (N_9186,N_6596,N_6038);
or U9187 (N_9187,N_6024,N_6173);
nor U9188 (N_9188,N_7793,N_7352);
nor U9189 (N_9189,N_7343,N_7442);
xnor U9190 (N_9190,N_7607,N_7024);
or U9191 (N_9191,N_7794,N_7455);
nor U9192 (N_9192,N_7055,N_7613);
nand U9193 (N_9193,N_6668,N_6309);
xor U9194 (N_9194,N_6852,N_7172);
xnor U9195 (N_9195,N_7863,N_6425);
or U9196 (N_9196,N_6268,N_7643);
and U9197 (N_9197,N_6422,N_6301);
and U9198 (N_9198,N_7862,N_7372);
and U9199 (N_9199,N_7074,N_7197);
nand U9200 (N_9200,N_7498,N_6611);
nand U9201 (N_9201,N_6562,N_6961);
xor U9202 (N_9202,N_7327,N_6971);
nor U9203 (N_9203,N_7520,N_6775);
nor U9204 (N_9204,N_6487,N_7454);
and U9205 (N_9205,N_6529,N_6321);
and U9206 (N_9206,N_7116,N_7043);
and U9207 (N_9207,N_7296,N_7565);
or U9208 (N_9208,N_7836,N_7410);
or U9209 (N_9209,N_6692,N_6691);
nor U9210 (N_9210,N_6984,N_7226);
nor U9211 (N_9211,N_6994,N_6150);
or U9212 (N_9212,N_6628,N_6903);
and U9213 (N_9213,N_6153,N_6693);
or U9214 (N_9214,N_7151,N_7495);
and U9215 (N_9215,N_6282,N_6122);
and U9216 (N_9216,N_7675,N_7751);
nand U9217 (N_9217,N_6924,N_6776);
nand U9218 (N_9218,N_6048,N_6390);
xor U9219 (N_9219,N_7182,N_7015);
or U9220 (N_9220,N_6379,N_7062);
or U9221 (N_9221,N_6044,N_7569);
xnor U9222 (N_9222,N_6164,N_7696);
nor U9223 (N_9223,N_7386,N_6829);
or U9224 (N_9224,N_6086,N_6118);
and U9225 (N_9225,N_6050,N_6671);
or U9226 (N_9226,N_6371,N_6887);
nand U9227 (N_9227,N_6932,N_6785);
xor U9228 (N_9228,N_6614,N_6503);
or U9229 (N_9229,N_7810,N_6760);
or U9230 (N_9230,N_6766,N_7401);
or U9231 (N_9231,N_6706,N_6551);
nand U9232 (N_9232,N_6457,N_7833);
and U9233 (N_9233,N_7513,N_7420);
and U9234 (N_9234,N_7137,N_7735);
or U9235 (N_9235,N_7636,N_6814);
and U9236 (N_9236,N_7995,N_7419);
nor U9237 (N_9237,N_7579,N_6846);
and U9238 (N_9238,N_7109,N_7840);
nor U9239 (N_9239,N_6771,N_6232);
or U9240 (N_9240,N_7084,N_6261);
or U9241 (N_9241,N_7272,N_7665);
or U9242 (N_9242,N_7705,N_6191);
nand U9243 (N_9243,N_6628,N_6864);
and U9244 (N_9244,N_6370,N_6633);
xnor U9245 (N_9245,N_6875,N_7181);
xnor U9246 (N_9246,N_7613,N_6344);
and U9247 (N_9247,N_7978,N_7652);
xor U9248 (N_9248,N_7839,N_6087);
and U9249 (N_9249,N_7595,N_6168);
or U9250 (N_9250,N_6792,N_7125);
xnor U9251 (N_9251,N_6340,N_7645);
nor U9252 (N_9252,N_6496,N_7666);
or U9253 (N_9253,N_6387,N_6225);
and U9254 (N_9254,N_7888,N_7319);
nor U9255 (N_9255,N_6233,N_7790);
nor U9256 (N_9256,N_7794,N_6109);
xor U9257 (N_9257,N_6700,N_6263);
xor U9258 (N_9258,N_7700,N_6387);
nor U9259 (N_9259,N_7465,N_6433);
or U9260 (N_9260,N_7873,N_6833);
or U9261 (N_9261,N_6572,N_6607);
nand U9262 (N_9262,N_7019,N_7863);
xor U9263 (N_9263,N_6922,N_6629);
or U9264 (N_9264,N_7331,N_6474);
nor U9265 (N_9265,N_7741,N_7033);
and U9266 (N_9266,N_7090,N_6674);
and U9267 (N_9267,N_6661,N_7890);
nand U9268 (N_9268,N_6397,N_6601);
nand U9269 (N_9269,N_7579,N_6251);
or U9270 (N_9270,N_7866,N_6039);
nand U9271 (N_9271,N_6596,N_7805);
nand U9272 (N_9272,N_6578,N_7675);
and U9273 (N_9273,N_7263,N_6743);
or U9274 (N_9274,N_7401,N_7083);
or U9275 (N_9275,N_6719,N_7621);
xnor U9276 (N_9276,N_7227,N_7894);
nor U9277 (N_9277,N_6379,N_7709);
nand U9278 (N_9278,N_7903,N_7857);
nor U9279 (N_9279,N_7194,N_7423);
or U9280 (N_9280,N_6494,N_7838);
nor U9281 (N_9281,N_7069,N_7730);
nand U9282 (N_9282,N_7816,N_6607);
and U9283 (N_9283,N_7276,N_6401);
nor U9284 (N_9284,N_7877,N_7329);
or U9285 (N_9285,N_7248,N_6323);
and U9286 (N_9286,N_6274,N_6562);
nand U9287 (N_9287,N_6414,N_7154);
and U9288 (N_9288,N_7365,N_7955);
nor U9289 (N_9289,N_6500,N_7665);
or U9290 (N_9290,N_6273,N_7491);
nor U9291 (N_9291,N_6889,N_6990);
nor U9292 (N_9292,N_6148,N_7725);
or U9293 (N_9293,N_7299,N_6882);
nor U9294 (N_9294,N_6381,N_6254);
nand U9295 (N_9295,N_7029,N_7985);
nor U9296 (N_9296,N_6579,N_6004);
nand U9297 (N_9297,N_6060,N_7423);
and U9298 (N_9298,N_7995,N_7001);
and U9299 (N_9299,N_7827,N_6181);
nor U9300 (N_9300,N_6743,N_6840);
or U9301 (N_9301,N_7312,N_6656);
nor U9302 (N_9302,N_6827,N_6591);
nor U9303 (N_9303,N_6257,N_6876);
nand U9304 (N_9304,N_6458,N_6735);
nor U9305 (N_9305,N_6450,N_6301);
or U9306 (N_9306,N_7528,N_7074);
or U9307 (N_9307,N_7902,N_6140);
or U9308 (N_9308,N_7379,N_7801);
or U9309 (N_9309,N_6106,N_6500);
nor U9310 (N_9310,N_6002,N_6380);
xnor U9311 (N_9311,N_6841,N_6248);
xnor U9312 (N_9312,N_6571,N_7727);
nor U9313 (N_9313,N_7815,N_7834);
and U9314 (N_9314,N_7653,N_7013);
nor U9315 (N_9315,N_7485,N_7067);
and U9316 (N_9316,N_7336,N_7186);
or U9317 (N_9317,N_6278,N_6968);
and U9318 (N_9318,N_7925,N_7244);
or U9319 (N_9319,N_6276,N_6546);
nand U9320 (N_9320,N_6288,N_7470);
nand U9321 (N_9321,N_7718,N_7748);
or U9322 (N_9322,N_7860,N_7467);
nand U9323 (N_9323,N_7203,N_7611);
xor U9324 (N_9324,N_7090,N_7097);
and U9325 (N_9325,N_7005,N_7399);
or U9326 (N_9326,N_7713,N_6813);
and U9327 (N_9327,N_7359,N_6116);
nand U9328 (N_9328,N_6343,N_6058);
nand U9329 (N_9329,N_6845,N_6502);
nor U9330 (N_9330,N_6384,N_6916);
nand U9331 (N_9331,N_6300,N_6079);
nand U9332 (N_9332,N_7142,N_6984);
and U9333 (N_9333,N_6631,N_6883);
nand U9334 (N_9334,N_7083,N_6438);
and U9335 (N_9335,N_7425,N_7738);
or U9336 (N_9336,N_6570,N_7857);
xor U9337 (N_9337,N_7977,N_7967);
xor U9338 (N_9338,N_6603,N_6638);
or U9339 (N_9339,N_7392,N_7123);
or U9340 (N_9340,N_7642,N_6866);
or U9341 (N_9341,N_6481,N_7382);
and U9342 (N_9342,N_6230,N_7997);
or U9343 (N_9343,N_7910,N_6585);
or U9344 (N_9344,N_7789,N_6570);
or U9345 (N_9345,N_7663,N_6240);
nand U9346 (N_9346,N_6007,N_6823);
nand U9347 (N_9347,N_7928,N_6690);
nor U9348 (N_9348,N_6248,N_7552);
and U9349 (N_9349,N_6545,N_6761);
nand U9350 (N_9350,N_6131,N_7688);
or U9351 (N_9351,N_6166,N_7451);
and U9352 (N_9352,N_7857,N_6146);
and U9353 (N_9353,N_7975,N_6651);
and U9354 (N_9354,N_6349,N_7225);
nor U9355 (N_9355,N_7894,N_7207);
nand U9356 (N_9356,N_6927,N_7415);
xnor U9357 (N_9357,N_6381,N_7061);
nor U9358 (N_9358,N_6563,N_7903);
or U9359 (N_9359,N_6100,N_7626);
or U9360 (N_9360,N_6511,N_6529);
nor U9361 (N_9361,N_6039,N_7153);
or U9362 (N_9362,N_6195,N_7900);
and U9363 (N_9363,N_7699,N_7048);
nor U9364 (N_9364,N_6028,N_6341);
nand U9365 (N_9365,N_7405,N_6129);
nand U9366 (N_9366,N_6226,N_7400);
and U9367 (N_9367,N_6687,N_6465);
nor U9368 (N_9368,N_6275,N_7916);
or U9369 (N_9369,N_7373,N_7034);
nand U9370 (N_9370,N_7466,N_7738);
or U9371 (N_9371,N_6474,N_6840);
or U9372 (N_9372,N_6241,N_6538);
or U9373 (N_9373,N_6815,N_7180);
or U9374 (N_9374,N_7779,N_6597);
or U9375 (N_9375,N_7209,N_6144);
and U9376 (N_9376,N_6604,N_7462);
xnor U9377 (N_9377,N_6426,N_7174);
nor U9378 (N_9378,N_7998,N_7731);
and U9379 (N_9379,N_6717,N_6428);
or U9380 (N_9380,N_7861,N_6027);
or U9381 (N_9381,N_7395,N_7184);
nor U9382 (N_9382,N_7635,N_7484);
or U9383 (N_9383,N_6984,N_6213);
and U9384 (N_9384,N_6992,N_7772);
xnor U9385 (N_9385,N_7185,N_6067);
nor U9386 (N_9386,N_6710,N_6630);
nand U9387 (N_9387,N_7912,N_6224);
and U9388 (N_9388,N_7680,N_6620);
and U9389 (N_9389,N_6551,N_6016);
xnor U9390 (N_9390,N_7549,N_6209);
nor U9391 (N_9391,N_7481,N_7935);
xnor U9392 (N_9392,N_7014,N_6418);
nor U9393 (N_9393,N_6157,N_6827);
nand U9394 (N_9394,N_6589,N_7694);
xnor U9395 (N_9395,N_7735,N_6648);
and U9396 (N_9396,N_7914,N_6127);
nor U9397 (N_9397,N_7139,N_7539);
xor U9398 (N_9398,N_7794,N_6494);
nand U9399 (N_9399,N_6872,N_7937);
and U9400 (N_9400,N_6849,N_6010);
xor U9401 (N_9401,N_7826,N_7354);
or U9402 (N_9402,N_6856,N_6322);
nor U9403 (N_9403,N_6978,N_7102);
or U9404 (N_9404,N_7595,N_6940);
xor U9405 (N_9405,N_6739,N_6328);
and U9406 (N_9406,N_6295,N_7302);
or U9407 (N_9407,N_6634,N_7693);
xor U9408 (N_9408,N_7500,N_6243);
or U9409 (N_9409,N_7515,N_7331);
nor U9410 (N_9410,N_6223,N_7295);
nor U9411 (N_9411,N_6739,N_6187);
nor U9412 (N_9412,N_7414,N_7810);
and U9413 (N_9413,N_7366,N_6124);
or U9414 (N_9414,N_6534,N_6771);
xnor U9415 (N_9415,N_6942,N_7528);
and U9416 (N_9416,N_7364,N_6890);
nor U9417 (N_9417,N_6014,N_6803);
xor U9418 (N_9418,N_7052,N_6923);
xor U9419 (N_9419,N_7529,N_6574);
xnor U9420 (N_9420,N_6056,N_7305);
nor U9421 (N_9421,N_6397,N_6912);
nor U9422 (N_9422,N_7230,N_7142);
nor U9423 (N_9423,N_7655,N_7194);
and U9424 (N_9424,N_7002,N_7474);
or U9425 (N_9425,N_7057,N_6596);
xor U9426 (N_9426,N_6220,N_6002);
or U9427 (N_9427,N_6189,N_7689);
xor U9428 (N_9428,N_6800,N_6608);
or U9429 (N_9429,N_6490,N_7829);
nor U9430 (N_9430,N_6212,N_7084);
or U9431 (N_9431,N_7121,N_6394);
or U9432 (N_9432,N_7570,N_7590);
xor U9433 (N_9433,N_6620,N_6721);
nand U9434 (N_9434,N_7149,N_6074);
and U9435 (N_9435,N_6339,N_6293);
and U9436 (N_9436,N_6997,N_7765);
nor U9437 (N_9437,N_7348,N_6771);
xor U9438 (N_9438,N_7119,N_7060);
or U9439 (N_9439,N_7774,N_6395);
nor U9440 (N_9440,N_7093,N_6585);
and U9441 (N_9441,N_6115,N_7158);
nand U9442 (N_9442,N_6776,N_7706);
nor U9443 (N_9443,N_6518,N_6192);
or U9444 (N_9444,N_6064,N_7663);
nand U9445 (N_9445,N_6774,N_7787);
nand U9446 (N_9446,N_7984,N_6998);
nor U9447 (N_9447,N_7979,N_6898);
or U9448 (N_9448,N_7222,N_6199);
xor U9449 (N_9449,N_7570,N_6214);
nand U9450 (N_9450,N_6591,N_7861);
and U9451 (N_9451,N_7755,N_6702);
nand U9452 (N_9452,N_7471,N_6647);
xnor U9453 (N_9453,N_7358,N_6646);
xnor U9454 (N_9454,N_7481,N_7066);
xor U9455 (N_9455,N_7957,N_6765);
and U9456 (N_9456,N_7814,N_6736);
xnor U9457 (N_9457,N_7802,N_6123);
and U9458 (N_9458,N_7387,N_6430);
nand U9459 (N_9459,N_7125,N_6185);
nand U9460 (N_9460,N_7056,N_7929);
xor U9461 (N_9461,N_7068,N_6091);
or U9462 (N_9462,N_6972,N_6527);
and U9463 (N_9463,N_6833,N_7201);
xor U9464 (N_9464,N_7199,N_7696);
nand U9465 (N_9465,N_6617,N_7520);
or U9466 (N_9466,N_6621,N_7501);
nor U9467 (N_9467,N_7597,N_6779);
xnor U9468 (N_9468,N_7415,N_7815);
xor U9469 (N_9469,N_7689,N_6487);
nor U9470 (N_9470,N_7988,N_6154);
xnor U9471 (N_9471,N_7373,N_7264);
or U9472 (N_9472,N_6153,N_6107);
nand U9473 (N_9473,N_7760,N_6853);
xnor U9474 (N_9474,N_6655,N_6545);
or U9475 (N_9475,N_6139,N_6274);
nor U9476 (N_9476,N_6542,N_7485);
or U9477 (N_9477,N_7553,N_6420);
nand U9478 (N_9478,N_7799,N_6109);
xor U9479 (N_9479,N_7533,N_6985);
or U9480 (N_9480,N_7053,N_6173);
nor U9481 (N_9481,N_6764,N_7752);
or U9482 (N_9482,N_7667,N_6838);
nor U9483 (N_9483,N_7529,N_7941);
nor U9484 (N_9484,N_6290,N_6203);
nand U9485 (N_9485,N_7702,N_6979);
or U9486 (N_9486,N_6997,N_6987);
or U9487 (N_9487,N_6374,N_6859);
xor U9488 (N_9488,N_7499,N_7824);
or U9489 (N_9489,N_6441,N_6626);
or U9490 (N_9490,N_6015,N_6858);
nand U9491 (N_9491,N_6556,N_6908);
and U9492 (N_9492,N_6915,N_7842);
nand U9493 (N_9493,N_6692,N_6423);
and U9494 (N_9494,N_7472,N_7689);
nor U9495 (N_9495,N_6532,N_6542);
nand U9496 (N_9496,N_7339,N_6675);
nand U9497 (N_9497,N_7083,N_6350);
xnor U9498 (N_9498,N_6461,N_6876);
and U9499 (N_9499,N_6409,N_6748);
xnor U9500 (N_9500,N_7742,N_7622);
nor U9501 (N_9501,N_7708,N_6798);
xor U9502 (N_9502,N_7730,N_7204);
and U9503 (N_9503,N_6529,N_7653);
nand U9504 (N_9504,N_6749,N_7230);
and U9505 (N_9505,N_7952,N_7638);
nand U9506 (N_9506,N_6564,N_7339);
nor U9507 (N_9507,N_6255,N_7804);
and U9508 (N_9508,N_7407,N_7240);
xor U9509 (N_9509,N_7738,N_6286);
nand U9510 (N_9510,N_7269,N_7716);
and U9511 (N_9511,N_6693,N_6791);
or U9512 (N_9512,N_7499,N_7944);
xor U9513 (N_9513,N_6110,N_6781);
or U9514 (N_9514,N_6324,N_6739);
and U9515 (N_9515,N_7234,N_7083);
nor U9516 (N_9516,N_7167,N_7305);
nor U9517 (N_9517,N_7737,N_6973);
nor U9518 (N_9518,N_6862,N_7149);
and U9519 (N_9519,N_7133,N_6928);
nor U9520 (N_9520,N_7328,N_7300);
xnor U9521 (N_9521,N_7697,N_7852);
nor U9522 (N_9522,N_6615,N_6694);
nor U9523 (N_9523,N_6943,N_6669);
xnor U9524 (N_9524,N_7666,N_7151);
and U9525 (N_9525,N_6623,N_6078);
nor U9526 (N_9526,N_7121,N_6040);
nand U9527 (N_9527,N_6635,N_6084);
or U9528 (N_9528,N_7988,N_6486);
xor U9529 (N_9529,N_7791,N_7398);
and U9530 (N_9530,N_6928,N_7361);
and U9531 (N_9531,N_6833,N_6270);
nand U9532 (N_9532,N_7965,N_6932);
and U9533 (N_9533,N_7749,N_7525);
xnor U9534 (N_9534,N_7340,N_7637);
xnor U9535 (N_9535,N_7209,N_6028);
or U9536 (N_9536,N_6920,N_6794);
xor U9537 (N_9537,N_7305,N_6908);
xor U9538 (N_9538,N_7790,N_7836);
nand U9539 (N_9539,N_6330,N_6076);
nor U9540 (N_9540,N_7422,N_6613);
nor U9541 (N_9541,N_6255,N_7633);
and U9542 (N_9542,N_7449,N_6357);
xor U9543 (N_9543,N_7184,N_6196);
or U9544 (N_9544,N_6131,N_7414);
xor U9545 (N_9545,N_6168,N_7105);
and U9546 (N_9546,N_6322,N_6248);
nor U9547 (N_9547,N_6694,N_7000);
nor U9548 (N_9548,N_6194,N_6825);
nand U9549 (N_9549,N_7979,N_6385);
and U9550 (N_9550,N_6759,N_7968);
and U9551 (N_9551,N_6745,N_6959);
or U9552 (N_9552,N_7897,N_7427);
xnor U9553 (N_9553,N_7107,N_6506);
xnor U9554 (N_9554,N_6210,N_6770);
nand U9555 (N_9555,N_7381,N_7510);
or U9556 (N_9556,N_7645,N_6164);
xor U9557 (N_9557,N_7968,N_7897);
or U9558 (N_9558,N_7808,N_7354);
or U9559 (N_9559,N_7633,N_6928);
xor U9560 (N_9560,N_7934,N_6060);
nor U9561 (N_9561,N_6240,N_6913);
nand U9562 (N_9562,N_7773,N_6380);
or U9563 (N_9563,N_6962,N_7010);
and U9564 (N_9564,N_6346,N_7133);
nand U9565 (N_9565,N_6997,N_6357);
nor U9566 (N_9566,N_7197,N_6206);
xor U9567 (N_9567,N_7257,N_7604);
or U9568 (N_9568,N_7390,N_6522);
and U9569 (N_9569,N_6219,N_6040);
and U9570 (N_9570,N_7415,N_7169);
or U9571 (N_9571,N_7218,N_6969);
and U9572 (N_9572,N_6075,N_7327);
or U9573 (N_9573,N_6341,N_7311);
xor U9574 (N_9574,N_6161,N_6645);
or U9575 (N_9575,N_6958,N_6935);
and U9576 (N_9576,N_7757,N_7020);
or U9577 (N_9577,N_6572,N_7042);
and U9578 (N_9578,N_6133,N_7960);
and U9579 (N_9579,N_6834,N_6493);
nand U9580 (N_9580,N_6318,N_6601);
nor U9581 (N_9581,N_7253,N_7496);
and U9582 (N_9582,N_7388,N_7103);
or U9583 (N_9583,N_6780,N_7286);
nand U9584 (N_9584,N_6093,N_6926);
nand U9585 (N_9585,N_7229,N_7969);
nand U9586 (N_9586,N_6760,N_7208);
or U9587 (N_9587,N_7638,N_7379);
nand U9588 (N_9588,N_6005,N_6640);
nor U9589 (N_9589,N_6684,N_6128);
and U9590 (N_9590,N_7048,N_6807);
or U9591 (N_9591,N_7408,N_7027);
and U9592 (N_9592,N_7347,N_7781);
and U9593 (N_9593,N_7269,N_6392);
and U9594 (N_9594,N_7315,N_7512);
or U9595 (N_9595,N_6136,N_7492);
nor U9596 (N_9596,N_7358,N_6200);
nand U9597 (N_9597,N_7902,N_6884);
and U9598 (N_9598,N_6030,N_7327);
nand U9599 (N_9599,N_6195,N_6473);
or U9600 (N_9600,N_7143,N_6056);
nor U9601 (N_9601,N_7114,N_7758);
nor U9602 (N_9602,N_6910,N_7918);
nor U9603 (N_9603,N_7150,N_7057);
nor U9604 (N_9604,N_7683,N_6372);
nand U9605 (N_9605,N_7436,N_6900);
nor U9606 (N_9606,N_6647,N_7112);
and U9607 (N_9607,N_6954,N_7773);
nor U9608 (N_9608,N_6746,N_7593);
xnor U9609 (N_9609,N_6197,N_6866);
xnor U9610 (N_9610,N_6575,N_6887);
or U9611 (N_9611,N_6703,N_7523);
nor U9612 (N_9612,N_6239,N_7902);
nor U9613 (N_9613,N_7515,N_7617);
and U9614 (N_9614,N_6719,N_6200);
xnor U9615 (N_9615,N_7810,N_6031);
or U9616 (N_9616,N_6553,N_7900);
xor U9617 (N_9617,N_6873,N_7577);
nor U9618 (N_9618,N_7331,N_6180);
xor U9619 (N_9619,N_7991,N_7731);
xnor U9620 (N_9620,N_6086,N_6810);
nand U9621 (N_9621,N_7322,N_6397);
nor U9622 (N_9622,N_7752,N_6521);
xnor U9623 (N_9623,N_6318,N_7509);
or U9624 (N_9624,N_6985,N_7884);
or U9625 (N_9625,N_7520,N_7451);
xnor U9626 (N_9626,N_6089,N_7238);
and U9627 (N_9627,N_7390,N_7699);
xor U9628 (N_9628,N_6069,N_6269);
or U9629 (N_9629,N_7640,N_6265);
nor U9630 (N_9630,N_7563,N_6550);
nor U9631 (N_9631,N_6757,N_6911);
nand U9632 (N_9632,N_7024,N_6381);
xor U9633 (N_9633,N_6655,N_6237);
nand U9634 (N_9634,N_7142,N_6282);
or U9635 (N_9635,N_7119,N_6729);
xnor U9636 (N_9636,N_6631,N_6922);
or U9637 (N_9637,N_6669,N_6696);
xor U9638 (N_9638,N_7506,N_7425);
or U9639 (N_9639,N_6630,N_6030);
xor U9640 (N_9640,N_6790,N_6956);
and U9641 (N_9641,N_6994,N_6874);
or U9642 (N_9642,N_7464,N_6811);
nor U9643 (N_9643,N_6860,N_7102);
or U9644 (N_9644,N_7745,N_7789);
nor U9645 (N_9645,N_6890,N_7003);
nand U9646 (N_9646,N_6768,N_6420);
xnor U9647 (N_9647,N_7106,N_6160);
nand U9648 (N_9648,N_7567,N_7051);
nor U9649 (N_9649,N_6138,N_7728);
nand U9650 (N_9650,N_6486,N_7141);
xor U9651 (N_9651,N_7623,N_6810);
nand U9652 (N_9652,N_7889,N_6601);
or U9653 (N_9653,N_6963,N_6321);
or U9654 (N_9654,N_6952,N_7458);
nor U9655 (N_9655,N_7108,N_7142);
nor U9656 (N_9656,N_6921,N_6844);
or U9657 (N_9657,N_6155,N_6498);
or U9658 (N_9658,N_6174,N_7538);
nor U9659 (N_9659,N_6190,N_6729);
nand U9660 (N_9660,N_7427,N_6754);
nand U9661 (N_9661,N_7430,N_6594);
nand U9662 (N_9662,N_7564,N_6036);
nor U9663 (N_9663,N_7151,N_7408);
nand U9664 (N_9664,N_7909,N_7294);
or U9665 (N_9665,N_7960,N_7367);
nor U9666 (N_9666,N_7992,N_6533);
xnor U9667 (N_9667,N_7412,N_7741);
nor U9668 (N_9668,N_6756,N_6159);
nor U9669 (N_9669,N_7822,N_7217);
or U9670 (N_9670,N_6699,N_7543);
or U9671 (N_9671,N_7302,N_6629);
nand U9672 (N_9672,N_7983,N_7637);
and U9673 (N_9673,N_7283,N_6167);
xor U9674 (N_9674,N_7384,N_7259);
nor U9675 (N_9675,N_7181,N_7122);
xor U9676 (N_9676,N_7473,N_6309);
and U9677 (N_9677,N_6951,N_6983);
and U9678 (N_9678,N_7225,N_6557);
or U9679 (N_9679,N_6236,N_7745);
and U9680 (N_9680,N_6464,N_7577);
xor U9681 (N_9681,N_6121,N_6938);
and U9682 (N_9682,N_6417,N_6198);
nor U9683 (N_9683,N_6965,N_7778);
nand U9684 (N_9684,N_6833,N_6507);
nor U9685 (N_9685,N_6293,N_7063);
or U9686 (N_9686,N_7632,N_7164);
and U9687 (N_9687,N_6767,N_7653);
xor U9688 (N_9688,N_6137,N_7172);
nor U9689 (N_9689,N_6933,N_6371);
nand U9690 (N_9690,N_7010,N_6940);
xor U9691 (N_9691,N_6629,N_7277);
or U9692 (N_9692,N_6775,N_7448);
xor U9693 (N_9693,N_7366,N_7055);
nor U9694 (N_9694,N_7923,N_6403);
nor U9695 (N_9695,N_7233,N_6210);
and U9696 (N_9696,N_6214,N_6556);
nand U9697 (N_9697,N_6005,N_7015);
nor U9698 (N_9698,N_6890,N_7297);
nand U9699 (N_9699,N_6822,N_6548);
nand U9700 (N_9700,N_6068,N_6981);
nand U9701 (N_9701,N_6626,N_7482);
xnor U9702 (N_9702,N_7142,N_7567);
nor U9703 (N_9703,N_6776,N_6762);
nand U9704 (N_9704,N_7804,N_7989);
and U9705 (N_9705,N_7951,N_7796);
xor U9706 (N_9706,N_6859,N_7298);
xor U9707 (N_9707,N_6798,N_7500);
or U9708 (N_9708,N_7649,N_7789);
and U9709 (N_9709,N_6478,N_6549);
and U9710 (N_9710,N_6247,N_6649);
nor U9711 (N_9711,N_7662,N_6018);
nand U9712 (N_9712,N_7994,N_6607);
nand U9713 (N_9713,N_6936,N_6123);
and U9714 (N_9714,N_7959,N_6145);
xor U9715 (N_9715,N_7678,N_7101);
nor U9716 (N_9716,N_7437,N_6126);
nand U9717 (N_9717,N_7276,N_6287);
xor U9718 (N_9718,N_6941,N_6858);
xnor U9719 (N_9719,N_7288,N_7897);
nor U9720 (N_9720,N_7738,N_7794);
nor U9721 (N_9721,N_6807,N_6319);
nor U9722 (N_9722,N_6746,N_7325);
nand U9723 (N_9723,N_7143,N_7658);
nand U9724 (N_9724,N_6400,N_6516);
xnor U9725 (N_9725,N_7132,N_7959);
nand U9726 (N_9726,N_6622,N_6852);
or U9727 (N_9727,N_7470,N_7427);
and U9728 (N_9728,N_7016,N_6461);
nand U9729 (N_9729,N_6301,N_6920);
or U9730 (N_9730,N_6924,N_6082);
or U9731 (N_9731,N_6931,N_7260);
and U9732 (N_9732,N_7540,N_6418);
or U9733 (N_9733,N_7795,N_6871);
nor U9734 (N_9734,N_7052,N_6357);
and U9735 (N_9735,N_7365,N_6185);
nor U9736 (N_9736,N_7655,N_6490);
nand U9737 (N_9737,N_7107,N_7597);
nand U9738 (N_9738,N_7736,N_7420);
and U9739 (N_9739,N_6055,N_7607);
or U9740 (N_9740,N_7003,N_7410);
nand U9741 (N_9741,N_6437,N_7838);
or U9742 (N_9742,N_6695,N_7520);
or U9743 (N_9743,N_6413,N_7203);
nand U9744 (N_9744,N_6788,N_6552);
or U9745 (N_9745,N_6658,N_6540);
xor U9746 (N_9746,N_7261,N_6606);
nand U9747 (N_9747,N_6639,N_6855);
nand U9748 (N_9748,N_7238,N_6232);
xor U9749 (N_9749,N_6435,N_6645);
nor U9750 (N_9750,N_7344,N_7959);
and U9751 (N_9751,N_6092,N_6316);
or U9752 (N_9752,N_7255,N_6032);
nand U9753 (N_9753,N_6276,N_7735);
and U9754 (N_9754,N_6132,N_6697);
nor U9755 (N_9755,N_7369,N_7698);
nor U9756 (N_9756,N_6700,N_6564);
nor U9757 (N_9757,N_7197,N_6051);
and U9758 (N_9758,N_7861,N_7352);
xnor U9759 (N_9759,N_7533,N_6111);
nand U9760 (N_9760,N_7869,N_6722);
nor U9761 (N_9761,N_7514,N_7151);
or U9762 (N_9762,N_6159,N_7555);
nand U9763 (N_9763,N_7250,N_6955);
nor U9764 (N_9764,N_6542,N_6014);
or U9765 (N_9765,N_7689,N_7648);
or U9766 (N_9766,N_7530,N_7355);
nand U9767 (N_9767,N_7290,N_7965);
xor U9768 (N_9768,N_6465,N_6965);
nand U9769 (N_9769,N_6666,N_7504);
xor U9770 (N_9770,N_7794,N_6761);
nor U9771 (N_9771,N_7452,N_6443);
nor U9772 (N_9772,N_7443,N_6001);
nand U9773 (N_9773,N_7267,N_6502);
or U9774 (N_9774,N_6233,N_7698);
nand U9775 (N_9775,N_7049,N_7420);
and U9776 (N_9776,N_6679,N_7284);
or U9777 (N_9777,N_6280,N_6909);
nand U9778 (N_9778,N_7493,N_6335);
nor U9779 (N_9779,N_6389,N_7516);
or U9780 (N_9780,N_7714,N_6234);
xnor U9781 (N_9781,N_6731,N_7013);
xnor U9782 (N_9782,N_7448,N_6023);
or U9783 (N_9783,N_6380,N_7193);
and U9784 (N_9784,N_7748,N_6650);
or U9785 (N_9785,N_7117,N_6978);
or U9786 (N_9786,N_7998,N_7062);
and U9787 (N_9787,N_6080,N_7532);
xor U9788 (N_9788,N_7219,N_7057);
or U9789 (N_9789,N_6050,N_6170);
nand U9790 (N_9790,N_7546,N_7625);
nand U9791 (N_9791,N_7670,N_7940);
nor U9792 (N_9792,N_7196,N_6373);
xor U9793 (N_9793,N_6045,N_7491);
nand U9794 (N_9794,N_6879,N_7147);
nand U9795 (N_9795,N_7860,N_6520);
and U9796 (N_9796,N_6383,N_7230);
xor U9797 (N_9797,N_7696,N_7974);
or U9798 (N_9798,N_6454,N_7083);
nand U9799 (N_9799,N_7569,N_7056);
or U9800 (N_9800,N_6428,N_6985);
or U9801 (N_9801,N_7271,N_7034);
nor U9802 (N_9802,N_7504,N_6626);
nor U9803 (N_9803,N_7517,N_6810);
nand U9804 (N_9804,N_6845,N_7944);
nand U9805 (N_9805,N_7389,N_7792);
nand U9806 (N_9806,N_7294,N_7445);
or U9807 (N_9807,N_7358,N_7397);
nand U9808 (N_9808,N_6954,N_7166);
xnor U9809 (N_9809,N_6568,N_7599);
and U9810 (N_9810,N_7049,N_6594);
nor U9811 (N_9811,N_6783,N_7816);
xnor U9812 (N_9812,N_6046,N_7453);
nor U9813 (N_9813,N_7746,N_6499);
and U9814 (N_9814,N_7658,N_6397);
and U9815 (N_9815,N_6733,N_7885);
nor U9816 (N_9816,N_7776,N_6626);
or U9817 (N_9817,N_7296,N_6593);
or U9818 (N_9818,N_6844,N_6609);
and U9819 (N_9819,N_7029,N_7675);
xor U9820 (N_9820,N_7685,N_6282);
nand U9821 (N_9821,N_6780,N_6778);
nand U9822 (N_9822,N_7538,N_6990);
xnor U9823 (N_9823,N_7248,N_7628);
xor U9824 (N_9824,N_7426,N_7406);
xor U9825 (N_9825,N_6582,N_6747);
nor U9826 (N_9826,N_6802,N_6755);
xnor U9827 (N_9827,N_7061,N_7120);
and U9828 (N_9828,N_6258,N_7542);
nand U9829 (N_9829,N_7705,N_7876);
nand U9830 (N_9830,N_6911,N_7607);
or U9831 (N_9831,N_7556,N_6336);
xnor U9832 (N_9832,N_7164,N_7673);
or U9833 (N_9833,N_6111,N_7084);
or U9834 (N_9834,N_6618,N_7442);
nand U9835 (N_9835,N_7700,N_7744);
nand U9836 (N_9836,N_7354,N_7223);
xor U9837 (N_9837,N_7331,N_7362);
xnor U9838 (N_9838,N_7800,N_7590);
or U9839 (N_9839,N_7311,N_7286);
nand U9840 (N_9840,N_6386,N_6005);
nand U9841 (N_9841,N_7898,N_7987);
and U9842 (N_9842,N_6659,N_7225);
nand U9843 (N_9843,N_6640,N_7965);
and U9844 (N_9844,N_6126,N_7782);
nand U9845 (N_9845,N_7194,N_6727);
and U9846 (N_9846,N_6584,N_6921);
and U9847 (N_9847,N_6100,N_7362);
or U9848 (N_9848,N_7553,N_6397);
xnor U9849 (N_9849,N_6893,N_7588);
nand U9850 (N_9850,N_6342,N_6099);
nand U9851 (N_9851,N_7071,N_7969);
or U9852 (N_9852,N_6636,N_6080);
nor U9853 (N_9853,N_6912,N_7085);
and U9854 (N_9854,N_6567,N_7554);
and U9855 (N_9855,N_7403,N_6384);
nor U9856 (N_9856,N_6210,N_7053);
xnor U9857 (N_9857,N_7980,N_7311);
nand U9858 (N_9858,N_7359,N_7556);
or U9859 (N_9859,N_7324,N_7178);
and U9860 (N_9860,N_7830,N_7088);
xor U9861 (N_9861,N_7034,N_6649);
or U9862 (N_9862,N_6598,N_6012);
or U9863 (N_9863,N_6974,N_6403);
or U9864 (N_9864,N_7807,N_6577);
nor U9865 (N_9865,N_6531,N_6865);
and U9866 (N_9866,N_6054,N_6970);
nor U9867 (N_9867,N_7496,N_7710);
xnor U9868 (N_9868,N_7700,N_7473);
xor U9869 (N_9869,N_6451,N_6095);
nor U9870 (N_9870,N_7482,N_6254);
or U9871 (N_9871,N_7180,N_7044);
xor U9872 (N_9872,N_7234,N_7181);
and U9873 (N_9873,N_7907,N_6366);
xnor U9874 (N_9874,N_6891,N_6177);
and U9875 (N_9875,N_6729,N_7674);
nand U9876 (N_9876,N_6310,N_6064);
or U9877 (N_9877,N_7935,N_7880);
or U9878 (N_9878,N_6293,N_7714);
or U9879 (N_9879,N_7327,N_6156);
or U9880 (N_9880,N_7875,N_7958);
nand U9881 (N_9881,N_6766,N_6179);
or U9882 (N_9882,N_7984,N_7498);
nor U9883 (N_9883,N_7160,N_7142);
and U9884 (N_9884,N_7335,N_7184);
and U9885 (N_9885,N_6043,N_7679);
nand U9886 (N_9886,N_7358,N_6456);
nor U9887 (N_9887,N_7855,N_7950);
nand U9888 (N_9888,N_6262,N_6916);
xnor U9889 (N_9889,N_7801,N_7138);
or U9890 (N_9890,N_7269,N_6886);
nor U9891 (N_9891,N_7046,N_7364);
nor U9892 (N_9892,N_6961,N_7875);
xnor U9893 (N_9893,N_7229,N_7373);
and U9894 (N_9894,N_6138,N_6147);
or U9895 (N_9895,N_6172,N_6968);
nor U9896 (N_9896,N_6011,N_6183);
or U9897 (N_9897,N_7765,N_7181);
or U9898 (N_9898,N_7718,N_7507);
xor U9899 (N_9899,N_7104,N_7712);
xor U9900 (N_9900,N_6407,N_7901);
nand U9901 (N_9901,N_6629,N_7470);
nor U9902 (N_9902,N_7234,N_6063);
and U9903 (N_9903,N_6168,N_7110);
nor U9904 (N_9904,N_6099,N_6593);
nand U9905 (N_9905,N_7399,N_6243);
and U9906 (N_9906,N_6602,N_7850);
or U9907 (N_9907,N_6858,N_7601);
nand U9908 (N_9908,N_7069,N_6241);
nand U9909 (N_9909,N_7733,N_7465);
and U9910 (N_9910,N_7807,N_7994);
nor U9911 (N_9911,N_6432,N_7745);
nand U9912 (N_9912,N_6659,N_7518);
and U9913 (N_9913,N_7790,N_6841);
or U9914 (N_9914,N_6062,N_7539);
and U9915 (N_9915,N_7683,N_6225);
xnor U9916 (N_9916,N_7627,N_7780);
or U9917 (N_9917,N_7539,N_6523);
nor U9918 (N_9918,N_7943,N_6542);
or U9919 (N_9919,N_7275,N_6316);
and U9920 (N_9920,N_7963,N_7981);
or U9921 (N_9921,N_6373,N_6485);
nand U9922 (N_9922,N_7400,N_6641);
or U9923 (N_9923,N_7247,N_6635);
or U9924 (N_9924,N_7208,N_6595);
and U9925 (N_9925,N_6333,N_6840);
xnor U9926 (N_9926,N_6348,N_6354);
and U9927 (N_9927,N_7194,N_6870);
nor U9928 (N_9928,N_7216,N_6857);
nor U9929 (N_9929,N_7432,N_6916);
or U9930 (N_9930,N_6779,N_6887);
and U9931 (N_9931,N_6606,N_6992);
nand U9932 (N_9932,N_7024,N_7079);
nand U9933 (N_9933,N_6387,N_6684);
xnor U9934 (N_9934,N_7633,N_7048);
nor U9935 (N_9935,N_6962,N_7315);
nand U9936 (N_9936,N_7858,N_7214);
xnor U9937 (N_9937,N_6539,N_6693);
nor U9938 (N_9938,N_7437,N_6933);
nor U9939 (N_9939,N_7849,N_6174);
or U9940 (N_9940,N_6834,N_6709);
and U9941 (N_9941,N_7946,N_7704);
or U9942 (N_9942,N_6026,N_6758);
and U9943 (N_9943,N_6259,N_6881);
nor U9944 (N_9944,N_7702,N_7142);
and U9945 (N_9945,N_7950,N_6786);
xor U9946 (N_9946,N_6699,N_6922);
or U9947 (N_9947,N_7491,N_6703);
nor U9948 (N_9948,N_7951,N_7242);
nor U9949 (N_9949,N_6700,N_6426);
xor U9950 (N_9950,N_7778,N_7745);
and U9951 (N_9951,N_6100,N_7710);
nand U9952 (N_9952,N_6245,N_6382);
nand U9953 (N_9953,N_6490,N_6790);
or U9954 (N_9954,N_7016,N_7493);
xnor U9955 (N_9955,N_6587,N_7558);
and U9956 (N_9956,N_7407,N_7469);
and U9957 (N_9957,N_7428,N_6564);
and U9958 (N_9958,N_6569,N_6050);
nor U9959 (N_9959,N_6771,N_6488);
nor U9960 (N_9960,N_6697,N_7397);
xor U9961 (N_9961,N_7124,N_7503);
nor U9962 (N_9962,N_6334,N_7617);
xnor U9963 (N_9963,N_7039,N_7762);
or U9964 (N_9964,N_6541,N_6107);
nor U9965 (N_9965,N_7983,N_7159);
nor U9966 (N_9966,N_7225,N_7086);
nor U9967 (N_9967,N_7223,N_7655);
xor U9968 (N_9968,N_6846,N_7049);
nand U9969 (N_9969,N_6064,N_7887);
xor U9970 (N_9970,N_6666,N_6048);
or U9971 (N_9971,N_7243,N_7765);
nand U9972 (N_9972,N_7519,N_7956);
xor U9973 (N_9973,N_7672,N_6809);
nand U9974 (N_9974,N_6902,N_6216);
xor U9975 (N_9975,N_7143,N_7886);
nand U9976 (N_9976,N_6598,N_7028);
or U9977 (N_9977,N_6545,N_7324);
nor U9978 (N_9978,N_7359,N_7099);
and U9979 (N_9979,N_6688,N_7766);
nor U9980 (N_9980,N_7195,N_6653);
nand U9981 (N_9981,N_7222,N_7386);
and U9982 (N_9982,N_7229,N_7319);
and U9983 (N_9983,N_6394,N_6767);
xnor U9984 (N_9984,N_7150,N_6268);
xor U9985 (N_9985,N_6334,N_7723);
nor U9986 (N_9986,N_7398,N_6553);
xnor U9987 (N_9987,N_6553,N_7884);
and U9988 (N_9988,N_7796,N_6599);
or U9989 (N_9989,N_7112,N_6723);
nand U9990 (N_9990,N_6385,N_6012);
xor U9991 (N_9991,N_7353,N_6142);
xor U9992 (N_9992,N_7623,N_6945);
nor U9993 (N_9993,N_7447,N_6536);
or U9994 (N_9994,N_6459,N_6738);
nor U9995 (N_9995,N_7662,N_7048);
nand U9996 (N_9996,N_6417,N_6080);
and U9997 (N_9997,N_7118,N_6419);
or U9998 (N_9998,N_7521,N_6434);
nand U9999 (N_9999,N_6486,N_7246);
nor U10000 (N_10000,N_9354,N_9351);
and U10001 (N_10001,N_9446,N_8139);
xnor U10002 (N_10002,N_9631,N_8847);
and U10003 (N_10003,N_9420,N_9416);
and U10004 (N_10004,N_8166,N_9261);
nor U10005 (N_10005,N_9089,N_8393);
and U10006 (N_10006,N_8553,N_8504);
xnor U10007 (N_10007,N_8782,N_8751);
xnor U10008 (N_10008,N_9186,N_9627);
xnor U10009 (N_10009,N_9174,N_8641);
and U10010 (N_10010,N_9094,N_9287);
nor U10011 (N_10011,N_9112,N_8586);
nor U10012 (N_10012,N_8060,N_8052);
xor U10013 (N_10013,N_8050,N_8106);
or U10014 (N_10014,N_8901,N_8981);
and U10015 (N_10015,N_8173,N_9408);
xnor U10016 (N_10016,N_9463,N_9377);
nand U10017 (N_10017,N_9756,N_9496);
and U10018 (N_10018,N_8008,N_8286);
xor U10019 (N_10019,N_8948,N_9888);
nor U10020 (N_10020,N_8792,N_9457);
nand U10021 (N_10021,N_9708,N_8328);
and U10022 (N_10022,N_8257,N_9647);
or U10023 (N_10023,N_9540,N_8157);
nor U10024 (N_10024,N_8491,N_9204);
nand U10025 (N_10025,N_9933,N_8089);
nor U10026 (N_10026,N_9221,N_9707);
or U10027 (N_10027,N_8592,N_9937);
nand U10028 (N_10028,N_8572,N_9476);
nand U10029 (N_10029,N_8868,N_8355);
xor U10030 (N_10030,N_9292,N_9034);
and U10031 (N_10031,N_9925,N_8450);
nand U10032 (N_10032,N_9431,N_8657);
nor U10033 (N_10033,N_9201,N_8967);
xor U10034 (N_10034,N_9171,N_8320);
and U10035 (N_10035,N_9185,N_8980);
xnor U10036 (N_10036,N_8266,N_8261);
or U10037 (N_10037,N_8447,N_9305);
xnor U10038 (N_10038,N_8585,N_8468);
and U10039 (N_10039,N_9447,N_8627);
xor U10040 (N_10040,N_9029,N_9227);
and U10041 (N_10041,N_9660,N_8741);
nand U10042 (N_10042,N_8777,N_9242);
and U10043 (N_10043,N_8081,N_8602);
or U10044 (N_10044,N_8875,N_8912);
nand U10045 (N_10045,N_9434,N_9704);
xnor U10046 (N_10046,N_9098,N_9720);
or U10047 (N_10047,N_9146,N_8839);
or U10048 (N_10048,N_9461,N_8742);
or U10049 (N_10049,N_9978,N_8323);
or U10050 (N_10050,N_8843,N_9914);
and U10051 (N_10051,N_9608,N_8453);
nand U10052 (N_10052,N_9999,N_8541);
nand U10053 (N_10053,N_9924,N_8509);
xnor U10054 (N_10054,N_8321,N_9423);
xnor U10055 (N_10055,N_9453,N_8965);
nand U10056 (N_10056,N_9963,N_8648);
nand U10057 (N_10057,N_9885,N_8047);
nor U10058 (N_10058,N_8814,N_9455);
or U10059 (N_10059,N_9593,N_8673);
nor U10060 (N_10060,N_9116,N_8217);
xnor U10061 (N_10061,N_9297,N_9003);
or U10062 (N_10062,N_9269,N_9807);
or U10063 (N_10063,N_9215,N_9679);
nor U10064 (N_10064,N_8688,N_8857);
and U10065 (N_10065,N_8154,N_9578);
nand U10066 (N_10066,N_8066,N_8189);
nand U10067 (N_10067,N_8376,N_9839);
nand U10068 (N_10068,N_9527,N_8512);
and U10069 (N_10069,N_8256,N_9726);
or U10070 (N_10070,N_8463,N_9570);
xnor U10071 (N_10071,N_9307,N_8579);
or U10072 (N_10072,N_9952,N_9485);
xnor U10073 (N_10073,N_8835,N_9219);
nor U10074 (N_10074,N_9024,N_8241);
and U10075 (N_10075,N_9896,N_9253);
or U10076 (N_10076,N_9109,N_9539);
nand U10077 (N_10077,N_9488,N_8822);
xor U10078 (N_10078,N_9993,N_8940);
nor U10079 (N_10079,N_8417,N_9519);
nand U10080 (N_10080,N_8097,N_8646);
xnor U10081 (N_10081,N_8775,N_8212);
nor U10082 (N_10082,N_8130,N_8853);
nor U10083 (N_10083,N_9267,N_8413);
or U10084 (N_10084,N_8730,N_9691);
nor U10085 (N_10085,N_8329,N_9622);
nor U10086 (N_10086,N_9567,N_8337);
nor U10087 (N_10087,N_9409,N_8921);
nor U10088 (N_10088,N_8536,N_9818);
nor U10089 (N_10089,N_8314,N_9370);
xor U10090 (N_10090,N_9609,N_9736);
xor U10091 (N_10091,N_8143,N_9342);
nor U10092 (N_10092,N_8976,N_9410);
xor U10093 (N_10093,N_8467,N_8045);
and U10094 (N_10094,N_9636,N_8518);
xor U10095 (N_10095,N_8435,N_9271);
and U10096 (N_10096,N_9779,N_8950);
or U10097 (N_10097,N_8736,N_9556);
and U10098 (N_10098,N_8459,N_9301);
and U10099 (N_10099,N_9376,N_8285);
nor U10100 (N_10100,N_8181,N_8497);
nor U10101 (N_10101,N_9421,N_9579);
nor U10102 (N_10102,N_8966,N_8169);
nor U10103 (N_10103,N_9590,N_9633);
nor U10104 (N_10104,N_9138,N_8483);
xor U10105 (N_10105,N_8599,N_9101);
xor U10106 (N_10106,N_9008,N_9440);
or U10107 (N_10107,N_8105,N_8327);
or U10108 (N_10108,N_9260,N_8028);
xnor U10109 (N_10109,N_9916,N_8119);
or U10110 (N_10110,N_8604,N_9365);
and U10111 (N_10111,N_9581,N_8872);
or U10112 (N_10112,N_9121,N_8810);
or U10113 (N_10113,N_9328,N_8942);
or U10114 (N_10114,N_9187,N_8394);
nor U10115 (N_10115,N_9536,N_8270);
nor U10116 (N_10116,N_8580,N_8725);
xnor U10117 (N_10117,N_9044,N_8564);
nand U10118 (N_10118,N_8003,N_9563);
nor U10119 (N_10119,N_8341,N_8218);
nand U10120 (N_10120,N_8142,N_9671);
nand U10121 (N_10121,N_8183,N_8860);
and U10122 (N_10122,N_9133,N_9306);
or U10123 (N_10123,N_9502,N_9213);
nor U10124 (N_10124,N_9787,N_8237);
nand U10125 (N_10125,N_8213,N_8044);
and U10126 (N_10126,N_8365,N_9979);
nor U10127 (N_10127,N_9758,N_9047);
nand U10128 (N_10128,N_8873,N_8684);
and U10129 (N_10129,N_9177,N_8158);
nand U10130 (N_10130,N_8554,N_8960);
or U10131 (N_10131,N_8722,N_9597);
and U10132 (N_10132,N_8914,N_8382);
nand U10133 (N_10133,N_9670,N_9415);
xnor U10134 (N_10134,N_9852,N_9768);
nor U10135 (N_10135,N_8910,N_9239);
and U10136 (N_10136,N_9694,N_8502);
or U10137 (N_10137,N_8350,N_9340);
nand U10138 (N_10138,N_9981,N_9676);
or U10139 (N_10139,N_9166,N_9036);
or U10140 (N_10140,N_8763,N_8631);
nand U10141 (N_10141,N_8523,N_8859);
and U10142 (N_10142,N_9811,N_8069);
and U10143 (N_10143,N_8304,N_9991);
and U10144 (N_10144,N_9737,N_8767);
xor U10145 (N_10145,N_9356,N_8471);
xor U10146 (N_10146,N_8973,N_8803);
and U10147 (N_10147,N_9533,N_9158);
or U10148 (N_10148,N_8771,N_9547);
or U10149 (N_10149,N_8390,N_9667);
nor U10150 (N_10150,N_9878,N_8146);
or U10151 (N_10151,N_9198,N_9445);
nor U10152 (N_10152,N_9890,N_8974);
nor U10153 (N_10153,N_8426,N_8824);
nand U10154 (N_10154,N_9809,N_8132);
or U10155 (N_10155,N_9231,N_8349);
or U10156 (N_10156,N_9551,N_8135);
or U10157 (N_10157,N_9998,N_9212);
or U10158 (N_10158,N_8208,N_8177);
nand U10159 (N_10159,N_8531,N_8882);
nand U10160 (N_10160,N_9110,N_8357);
or U10161 (N_10161,N_8419,N_8856);
or U10162 (N_10162,N_9197,N_9634);
xor U10163 (N_10163,N_8153,N_9398);
or U10164 (N_10164,N_8036,N_8443);
nor U10165 (N_10165,N_8638,N_9516);
or U10166 (N_10166,N_9841,N_8915);
or U10167 (N_10167,N_9135,N_8801);
nand U10168 (N_10168,N_9657,N_9915);
nand U10169 (N_10169,N_9908,N_8526);
or U10170 (N_10170,N_8225,N_9050);
nand U10171 (N_10171,N_9327,N_9065);
nand U10172 (N_10172,N_9318,N_8400);
or U10173 (N_10173,N_8291,N_9000);
nor U10174 (N_10174,N_9311,N_9298);
nor U10175 (N_10175,N_9395,N_9724);
xnor U10176 (N_10176,N_8269,N_8766);
or U10177 (N_10177,N_8494,N_9861);
nand U10178 (N_10178,N_9899,N_9299);
xor U10179 (N_10179,N_9247,N_8710);
and U10180 (N_10180,N_9483,N_9989);
nor U10181 (N_10181,N_9548,N_9823);
xor U10182 (N_10182,N_8529,N_8245);
or U10183 (N_10183,N_9680,N_9314);
nor U10184 (N_10184,N_8356,N_9601);
or U10185 (N_10185,N_9470,N_9644);
and U10186 (N_10186,N_9781,N_9450);
nand U10187 (N_10187,N_9437,N_8666);
nand U10188 (N_10188,N_9234,N_8378);
nor U10189 (N_10189,N_8031,N_8254);
nor U10190 (N_10190,N_8863,N_8652);
and U10191 (N_10191,N_8962,N_9595);
nand U10192 (N_10192,N_8242,N_9244);
xnor U10193 (N_10193,N_9586,N_8907);
or U10194 (N_10194,N_9405,N_9887);
nor U10195 (N_10195,N_8818,N_9430);
nand U10196 (N_10196,N_9514,N_8315);
and U10197 (N_10197,N_8834,N_9066);
and U10198 (N_10198,N_9172,N_8713);
or U10199 (N_10199,N_8452,N_8902);
nor U10200 (N_10200,N_8155,N_8439);
and U10201 (N_10201,N_8147,N_9790);
and U10202 (N_10202,N_8510,N_9134);
xor U10203 (N_10203,N_9873,N_8226);
or U10204 (N_10204,N_9294,N_9692);
nand U10205 (N_10205,N_8656,N_9725);
and U10206 (N_10206,N_8864,N_8959);
or U10207 (N_10207,N_9352,N_9642);
nor U10208 (N_10208,N_8540,N_9103);
nand U10209 (N_10209,N_8250,N_9557);
nor U10210 (N_10210,N_8401,N_9322);
nor U10211 (N_10211,N_9500,N_8871);
nand U10212 (N_10212,N_9009,N_9049);
nor U10213 (N_10213,N_9762,N_9976);
or U10214 (N_10214,N_8407,N_9684);
xnor U10215 (N_10215,N_9182,N_8065);
or U10216 (N_10216,N_9150,N_9569);
and U10217 (N_10217,N_8575,N_9111);
nand U10218 (N_10218,N_9958,N_8952);
and U10219 (N_10219,N_8107,N_9344);
xnor U10220 (N_10220,N_8140,N_9695);
nor U10221 (N_10221,N_8289,N_9599);
nand U10222 (N_10222,N_8555,N_9140);
nand U10223 (N_10223,N_8908,N_9630);
and U10224 (N_10224,N_9507,N_9895);
nor U10225 (N_10225,N_9286,N_8514);
nor U10226 (N_10226,N_9127,N_8787);
and U10227 (N_10227,N_9711,N_9025);
or U10228 (N_10228,N_8932,N_9700);
nor U10229 (N_10229,N_8519,N_8858);
or U10230 (N_10230,N_8612,N_8160);
xor U10231 (N_10231,N_8303,N_9960);
xor U10232 (N_10232,N_9490,N_8893);
and U10233 (N_10233,N_9938,N_9203);
nand U10234 (N_10234,N_8414,N_8903);
or U10235 (N_10235,N_8994,N_8347);
nand U10236 (N_10236,N_8373,N_9464);
xnor U10237 (N_10237,N_8535,N_9192);
or U10238 (N_10238,N_8570,N_8680);
and U10239 (N_10239,N_9100,N_8409);
nor U10240 (N_10240,N_8438,N_9153);
or U10241 (N_10241,N_9870,N_9503);
or U10242 (N_10242,N_8927,N_8802);
xor U10243 (N_10243,N_8682,N_9230);
nor U10244 (N_10244,N_9472,N_9478);
nor U10245 (N_10245,N_9857,N_9910);
nand U10246 (N_10246,N_8112,N_9649);
xnor U10247 (N_10247,N_8728,N_9773);
or U10248 (N_10248,N_8516,N_8849);
xnor U10249 (N_10249,N_9291,N_8668);
nor U10250 (N_10250,N_9739,N_8214);
nor U10251 (N_10251,N_8427,N_9308);
xnor U10252 (N_10252,N_9552,N_8551);
nor U10253 (N_10253,N_9295,N_9875);
xor U10254 (N_10254,N_9432,N_8622);
nand U10255 (N_10255,N_9935,N_9387);
and U10256 (N_10256,N_8170,N_9433);
nor U10257 (N_10257,N_9254,N_8244);
nand U10258 (N_10258,N_9335,N_9064);
nand U10259 (N_10259,N_8481,N_8358);
nor U10260 (N_10260,N_8636,N_8925);
nor U10261 (N_10261,N_8360,N_9836);
xor U10262 (N_10262,N_8005,N_8840);
or U10263 (N_10263,N_8505,N_9741);
or U10264 (N_10264,N_9619,N_9639);
or U10265 (N_10265,N_9929,N_8210);
or U10266 (N_10266,N_9575,N_8101);
nand U10267 (N_10267,N_8784,N_8207);
or U10268 (N_10268,N_9589,N_9235);
nor U10269 (N_10269,N_9827,N_8765);
nand U10270 (N_10270,N_9740,N_8808);
or U10271 (N_10271,N_8246,N_8986);
or U10272 (N_10272,N_8594,N_9079);
or U10273 (N_10273,N_9454,N_9296);
xnor U10274 (N_10274,N_8667,N_9822);
nor U10275 (N_10275,N_8593,N_9046);
nand U10276 (N_10276,N_9615,N_8030);
nor U10277 (N_10277,N_8404,N_8611);
nand U10278 (N_10278,N_8630,N_8054);
nand U10279 (N_10279,N_8022,N_9104);
xnor U10280 (N_10280,N_9374,N_9513);
and U10281 (N_10281,N_9394,N_8528);
and U10282 (N_10282,N_8440,N_8198);
or U10283 (N_10283,N_9414,N_9716);
xnor U10284 (N_10284,N_9643,N_9078);
nand U10285 (N_10285,N_9080,N_8361);
xnor U10286 (N_10286,N_8163,N_8807);
xnor U10287 (N_10287,N_9798,N_8074);
or U10288 (N_10288,N_8786,N_9777);
nor U10289 (N_10289,N_9444,N_8727);
and U10290 (N_10290,N_8862,N_9767);
and U10291 (N_10291,N_9002,N_8934);
xor U10292 (N_10292,N_8569,N_8281);
nor U10293 (N_10293,N_9661,N_9364);
nand U10294 (N_10294,N_8813,N_9091);
or U10295 (N_10295,N_9535,N_8283);
xor U10296 (N_10296,N_8869,N_9225);
and U10297 (N_10297,N_9710,N_9460);
xor U10298 (N_10298,N_9752,N_8928);
nand U10299 (N_10299,N_8778,N_8477);
or U10300 (N_10300,N_9125,N_8343);
nor U10301 (N_10301,N_8110,N_8661);
xor U10302 (N_10302,N_8263,N_9015);
nor U10303 (N_10303,N_9026,N_8092);
nand U10304 (N_10304,N_8423,N_9251);
and U10305 (N_10305,N_8574,N_9856);
or U10306 (N_10306,N_9031,N_8363);
nand U10307 (N_10307,N_8455,N_9126);
xor U10308 (N_10308,N_8756,N_8795);
and U10309 (N_10309,N_9392,N_8662);
or U10310 (N_10310,N_9013,N_8883);
nor U10311 (N_10311,N_8972,N_9648);
nand U10312 (N_10312,N_8821,N_8706);
nand U10313 (N_10313,N_8384,N_9977);
nor U10314 (N_10314,N_9092,N_9957);
xnor U10315 (N_10315,N_9577,N_8735);
nand U10316 (N_10316,N_8634,N_8276);
nor U10317 (N_10317,N_8560,N_9435);
nand U10318 (N_10318,N_9300,N_8220);
nand U10319 (N_10319,N_8456,N_9792);
xor U10320 (N_10320,N_8042,N_8164);
nand U10321 (N_10321,N_9738,N_9379);
and U10322 (N_10322,N_9764,N_8643);
nand U10323 (N_10323,N_9769,N_9391);
nand U10324 (N_10324,N_9288,N_9598);
nand U10325 (N_10325,N_9162,N_8041);
or U10326 (N_10326,N_8430,N_9477);
or U10327 (N_10327,N_9167,N_9161);
nor U10328 (N_10328,N_9638,N_9068);
nor U10329 (N_10329,N_9531,N_8156);
nor U10330 (N_10330,N_9129,N_9744);
xnor U10331 (N_10331,N_9393,N_8753);
xnor U10332 (N_10332,N_9947,N_8342);
xnor U10333 (N_10333,N_8024,N_8647);
nor U10334 (N_10334,N_9059,N_8332);
nand U10335 (N_10335,N_9232,N_9350);
nand U10336 (N_10336,N_9521,N_9316);
and U10337 (N_10337,N_8446,N_8597);
xor U10338 (N_10338,N_9217,N_9325);
and U10339 (N_10339,N_8654,N_9141);
nand U10340 (N_10340,N_9624,N_8739);
nand U10341 (N_10341,N_9629,N_8488);
nor U10342 (N_10342,N_9095,N_9165);
or U10343 (N_10343,N_8172,N_8239);
nor U10344 (N_10344,N_9336,N_9996);
or U10345 (N_10345,N_9677,N_8698);
xor U10346 (N_10346,N_9815,N_8374);
nand U10347 (N_10347,N_9117,N_8895);
and U10348 (N_10348,N_9688,N_9891);
xnor U10349 (N_10349,N_8761,N_9124);
nor U10350 (N_10350,N_9062,N_9346);
nor U10351 (N_10351,N_9210,N_9422);
nand U10352 (N_10352,N_9413,N_9195);
nand U10353 (N_10353,N_9149,N_9018);
nand U10354 (N_10354,N_8001,N_9179);
nand U10355 (N_10355,N_9632,N_8758);
nand U10356 (N_10356,N_9320,N_8268);
xnor U10357 (N_10357,N_8711,N_9900);
nand U10358 (N_10358,N_9946,N_9424);
nand U10359 (N_10359,N_8480,N_8705);
and U10360 (N_10360,N_9229,N_9984);
or U10361 (N_10361,N_9626,N_9438);
or U10362 (N_10362,N_8049,N_8415);
nor U10363 (N_10363,N_8434,N_8678);
nand U10364 (N_10364,N_8746,N_8364);
or U10365 (N_10365,N_9466,N_9714);
xor U10366 (N_10366,N_8136,N_8127);
nor U10367 (N_10367,N_9276,N_9971);
or U10368 (N_10368,N_9474,N_9867);
nand U10369 (N_10369,N_8262,N_9696);
nor U10370 (N_10370,N_8665,N_9682);
nor U10371 (N_10371,N_8428,N_8221);
nor U10372 (N_10372,N_9381,N_8436);
or U10373 (N_10373,N_8338,N_8398);
or U10374 (N_10374,N_9357,N_9911);
nand U10375 (N_10375,N_9909,N_8897);
nor U10376 (N_10376,N_8339,N_9982);
xor U10377 (N_10377,N_9537,N_9614);
xor U10378 (N_10378,N_9782,N_9193);
nor U10379 (N_10379,N_8577,N_9006);
and U10380 (N_10380,N_9530,N_9343);
and U10381 (N_10381,N_8125,N_8890);
and U10382 (N_10382,N_9600,N_8819);
nand U10383 (N_10383,N_9390,N_8836);
or U10384 (N_10384,N_9699,N_8197);
xnor U10385 (N_10385,N_9273,N_9238);
and U10386 (N_10386,N_9528,N_8995);
and U10387 (N_10387,N_8601,N_9526);
or U10388 (N_10388,N_9520,N_9169);
nand U10389 (N_10389,N_9456,N_9017);
nor U10390 (N_10390,N_9321,N_9718);
or U10391 (N_10391,N_8845,N_8124);
and U10392 (N_10392,N_9860,N_9067);
nand U10393 (N_10393,N_9912,N_9070);
nand U10394 (N_10394,N_8699,N_9128);
or U10395 (N_10395,N_8658,N_8708);
or U10396 (N_10396,N_9858,N_8492);
xnor U10397 (N_10397,N_9585,N_8876);
xnor U10398 (N_10398,N_8831,N_8410);
nand U10399 (N_10399,N_8230,N_8295);
nor U10400 (N_10400,N_9833,N_9345);
nor U10401 (N_10401,N_9021,N_9932);
or U10402 (N_10402,N_8877,N_9653);
and U10403 (N_10403,N_9214,N_9263);
xnor U10404 (N_10404,N_9156,N_8723);
and U10405 (N_10405,N_8366,N_8462);
nor U10406 (N_10406,N_9473,N_9208);
or U10407 (N_10407,N_8848,N_8993);
xnor U10408 (N_10408,N_8260,N_9917);
nand U10409 (N_10409,N_8754,N_9052);
nand U10410 (N_10410,N_8838,N_8117);
xnor U10411 (N_10411,N_9713,N_8053);
xor U10412 (N_10412,N_9705,N_8644);
and U10413 (N_10413,N_9130,N_9412);
or U10414 (N_10414,N_9250,N_9829);
or U10415 (N_10415,N_9039,N_9721);
and U10416 (N_10416,N_9850,N_8855);
nor U10417 (N_10417,N_8219,N_9505);
or U10418 (N_10418,N_8583,N_8991);
nor U10419 (N_10419,N_8354,N_8104);
nor U10420 (N_10420,N_9717,N_9011);
and U10421 (N_10421,N_9571,N_8947);
nor U10422 (N_10422,N_8305,N_9986);
nand U10423 (N_10423,N_9486,N_8996);
or U10424 (N_10424,N_9893,N_8206);
and U10425 (N_10425,N_8318,N_9765);
or U10426 (N_10426,N_8961,N_8576);
nor U10427 (N_10427,N_9555,N_9384);
xnor U10428 (N_10428,N_9702,N_9750);
nor U10429 (N_10429,N_9289,N_8812);
or U10430 (N_10430,N_9038,N_8825);
nand U10431 (N_10431,N_8501,N_8681);
or U10432 (N_10432,N_8930,N_8431);
nor U10433 (N_10433,N_9054,N_9236);
and U10434 (N_10434,N_9735,N_8016);
or U10435 (N_10435,N_9538,N_9151);
xor U10436 (N_10436,N_8773,N_9902);
xor U10437 (N_10437,N_8441,N_8204);
and U10438 (N_10438,N_9529,N_9517);
or U10439 (N_10439,N_8861,N_9800);
nand U10440 (N_10440,N_9821,N_8905);
or U10441 (N_10441,N_8396,N_8785);
xor U10442 (N_10442,N_9745,N_8618);
or U10443 (N_10443,N_9222,N_9259);
xnor U10444 (N_10444,N_8185,N_9831);
nor U10445 (N_10445,N_9027,N_8750);
and U10446 (N_10446,N_9030,N_9715);
nor U10447 (N_10447,N_8029,N_8235);
or U10448 (N_10448,N_9452,N_9617);
or U10449 (N_10449,N_8018,N_8793);
and U10450 (N_10450,N_9184,N_8120);
or U10451 (N_10451,N_8232,N_9766);
xnor U10452 (N_10452,N_9542,N_8815);
xor U10453 (N_10453,N_9220,N_8645);
xnor U10454 (N_10454,N_9774,N_8224);
nor U10455 (N_10455,N_8162,N_8700);
xnor U10456 (N_10456,N_8781,N_9180);
xnor U10457 (N_10457,N_9284,N_9939);
xor U10458 (N_10458,N_8889,N_9084);
and U10459 (N_10459,N_9894,N_9544);
nand U10460 (N_10460,N_9216,N_8625);
nor U10461 (N_10461,N_9931,N_9226);
nand U10462 (N_10462,N_8479,N_8258);
or U10463 (N_10463,N_8496,N_9077);
nand U10464 (N_10464,N_8402,N_9211);
or U10465 (N_10465,N_8628,N_9985);
nor U10466 (N_10466,N_8670,N_8999);
xor U10467 (N_10467,N_8885,N_8473);
nor U10468 (N_10468,N_8372,N_8669);
nand U10469 (N_10469,N_9572,N_9175);
and U10470 (N_10470,N_8179,N_8732);
xnor U10471 (N_10471,N_8223,N_8498);
or U10472 (N_10472,N_9145,N_9685);
and U10473 (N_10473,N_8465,N_9266);
nand U10474 (N_10474,N_9607,N_8685);
and U10475 (N_10475,N_8476,N_9990);
and U10476 (N_10476,N_9532,N_9341);
and U10477 (N_10477,N_8129,N_8904);
and U10478 (N_10478,N_8013,N_8038);
xor U10479 (N_10479,N_9451,N_8040);
xor U10480 (N_10480,N_8466,N_9268);
and U10481 (N_10481,N_9443,N_9338);
xor U10482 (N_10482,N_9975,N_9406);
xor U10483 (N_10483,N_8941,N_8264);
nand U10484 (N_10484,N_8701,N_8584);
nor U10485 (N_10485,N_8015,N_9603);
nor U10486 (N_10486,N_8368,N_8982);
and U10487 (N_10487,N_9869,N_8174);
nand U10488 (N_10488,N_9802,N_8037);
xor U10489 (N_10489,N_8547,N_9499);
nand U10490 (N_10490,N_8067,N_8137);
and U10491 (N_10491,N_9019,N_8333);
xor U10492 (N_10492,N_9275,N_9669);
xor U10493 (N_10493,N_8886,N_9360);
nor U10494 (N_10494,N_8588,N_8449);
nor U10495 (N_10495,N_8844,N_9348);
or U10496 (N_10496,N_9010,N_9848);
or U10497 (N_10497,N_9258,N_8093);
and U10498 (N_10498,N_9248,N_8236);
xor U10499 (N_10499,N_8126,N_9053);
and U10500 (N_10500,N_8086,N_8109);
nand U10501 (N_10501,N_8418,N_9930);
nand U10502 (N_10502,N_8587,N_9028);
nor U10503 (N_10503,N_8837,N_8716);
nand U10504 (N_10504,N_8403,N_8640);
and U10505 (N_10505,N_8425,N_8918);
or U10506 (N_10506,N_9160,N_9448);
nor U10507 (N_10507,N_8039,N_9865);
nand U10508 (N_10508,N_9223,N_8027);
nand U10509 (N_10509,N_9819,N_9202);
xnor U10510 (N_10510,N_9927,N_8433);
and U10511 (N_10511,N_8202,N_9339);
nand U10512 (N_10512,N_8820,N_8192);
nor U10513 (N_10513,N_9088,N_9131);
or U10514 (N_10514,N_9795,N_9518);
nand U10515 (N_10515,N_8805,N_8653);
xnor U10516 (N_10516,N_8809,N_8096);
nand U10517 (N_10517,N_8023,N_8309);
xor U10518 (N_10518,N_9945,N_8772);
and U10519 (N_10519,N_8788,N_8954);
and U10520 (N_10520,N_8544,N_8530);
or U10521 (N_10521,N_9954,N_8282);
xnor U10522 (N_10522,N_9206,N_8149);
xor U10523 (N_10523,N_9799,N_8387);
nor U10524 (N_10524,N_9972,N_9664);
and U10525 (N_10525,N_8935,N_8102);
or U10526 (N_10526,N_8098,N_8804);
nand U10527 (N_10527,N_9363,N_8629);
or U10528 (N_10528,N_9573,N_9749);
or U10529 (N_10529,N_8048,N_9561);
xnor U10530 (N_10530,N_8745,N_9805);
nand U10531 (N_10531,N_9083,N_8412);
nor U10532 (N_10532,N_9326,N_9879);
xor U10533 (N_10533,N_8478,N_9582);
or U10534 (N_10534,N_8308,N_9241);
and U10535 (N_10535,N_8300,N_8513);
and U10536 (N_10536,N_9734,N_8184);
xnor U10537 (N_10537,N_8073,N_8796);
xor U10538 (N_10538,N_8689,N_8987);
or U10539 (N_10539,N_8951,N_9386);
nand U10540 (N_10540,N_8021,N_8752);
or U10541 (N_10541,N_9042,N_9703);
nand U10542 (N_10542,N_8231,N_8764);
nand U10543 (N_10543,N_9099,N_8979);
nor U10544 (N_10544,N_8194,N_9918);
and U10545 (N_10545,N_8381,N_8297);
and U10546 (N_10546,N_9040,N_9761);
and U10547 (N_10547,N_9621,N_8159);
nor U10548 (N_10548,N_8850,N_8150);
xor U10549 (N_10549,N_9817,N_8963);
and U10550 (N_10550,N_8550,N_9257);
nand U10551 (N_10551,N_8284,N_8088);
nor U10552 (N_10552,N_9966,N_9706);
and U10553 (N_10553,N_9380,N_8058);
nor U10554 (N_10554,N_8542,N_8894);
nor U10555 (N_10555,N_9402,N_8377);
nor U10556 (N_10556,N_9233,N_9136);
nor U10557 (N_10557,N_9033,N_9304);
nand U10558 (N_10558,N_8080,N_9283);
nor U10559 (N_10559,N_9115,N_9093);
nor U10560 (N_10560,N_9139,N_9303);
and U10561 (N_10561,N_9584,N_9892);
xor U10562 (N_10562,N_9673,N_9007);
and U10563 (N_10563,N_9523,N_9546);
nand U10564 (N_10564,N_9602,N_9282);
xnor U10565 (N_10565,N_9388,N_9789);
nor U10566 (N_10566,N_9497,N_8919);
and U10567 (N_10567,N_9654,N_9926);
nand U10568 (N_10568,N_9674,N_8799);
nor U10569 (N_10569,N_9690,N_9375);
nor U10570 (N_10570,N_8079,N_8693);
or U10571 (N_10571,N_8552,N_9665);
xnor U10572 (N_10572,N_8664,N_8884);
and U10573 (N_10573,N_8019,N_8490);
or U10574 (N_10574,N_9190,N_8898);
nor U10575 (N_10575,N_8508,N_8249);
nand U10576 (N_10576,N_8511,N_9628);
or U10577 (N_10577,N_8051,N_9812);
nor U10578 (N_10578,N_9330,N_8193);
nand U10579 (N_10579,N_9425,N_8734);
xor U10580 (N_10580,N_9786,N_8589);
nor U10581 (N_10581,N_9479,N_9871);
or U10582 (N_10582,N_9032,N_8470);
nand U10583 (N_10583,N_8406,N_8559);
nor U10584 (N_10584,N_9090,N_8707);
nor U10585 (N_10585,N_9596,N_8116);
and U10586 (N_10586,N_9814,N_9237);
or U10587 (N_10587,N_8581,N_8989);
xor U10588 (N_10588,N_8687,N_9558);
nor U10589 (N_10589,N_9361,N_8527);
or U10590 (N_10590,N_9436,N_8141);
nand U10591 (N_10591,N_8046,N_8487);
nor U10592 (N_10592,N_9023,N_8953);
nor U10593 (N_10593,N_8334,N_9143);
xnor U10594 (N_10594,N_9606,N_9731);
or U10595 (N_10595,N_9278,N_9859);
nor U10596 (N_10596,N_9155,N_9041);
xnor U10597 (N_10597,N_8056,N_9515);
xor U10598 (N_10598,N_9057,N_9656);
xor U10599 (N_10599,N_8180,N_8774);
and U10600 (N_10600,N_9081,N_8100);
and U10601 (N_10601,N_9842,N_8026);
nor U10602 (N_10602,N_9323,N_9401);
or U10603 (N_10603,N_9411,N_9730);
nand U10604 (N_10604,N_8265,N_8720);
and U10605 (N_10605,N_9956,N_8442);
nand U10606 (N_10606,N_8151,N_8607);
nand U10607 (N_10607,N_9396,N_8448);
or U10608 (N_10608,N_9020,N_8211);
nand U10609 (N_10609,N_8798,N_9417);
or U10610 (N_10610,N_8424,N_8279);
nand U10611 (N_10611,N_8770,N_8562);
nor U10612 (N_10612,N_9613,N_8717);
xor U10613 (N_10613,N_8978,N_8168);
or U10614 (N_10614,N_8353,N_9672);
xor U10615 (N_10615,N_8486,N_8385);
nand U10616 (N_10616,N_9898,N_9449);
or U10617 (N_10617,N_8161,N_9844);
or U10618 (N_10618,N_9144,N_9564);
nor U10619 (N_10619,N_9906,N_9012);
nor U10620 (N_10620,N_9882,N_8128);
xnor U10621 (N_10621,N_8899,N_8134);
nand U10622 (N_10622,N_9426,N_8676);
nor U10623 (N_10623,N_9655,N_9541);
or U10624 (N_10624,N_8880,N_9853);
nand U10625 (N_10625,N_9096,N_9863);
xor U10626 (N_10626,N_9005,N_9701);
or U10627 (N_10627,N_9196,N_9534);
and U10628 (N_10628,N_8566,N_8521);
nor U10629 (N_10629,N_8233,N_9612);
nor U10630 (N_10630,N_9650,N_9968);
nand U10631 (N_10631,N_9407,N_9868);
nor U10632 (N_10632,N_9491,N_9492);
or U10633 (N_10633,N_8675,N_8990);
xnor U10634 (N_10634,N_8721,N_9319);
xnor U10635 (N_10635,N_8458,N_9880);
xor U10636 (N_10636,N_9512,N_8331);
and U10637 (N_10637,N_9825,N_9980);
or U10638 (N_10638,N_9776,N_9576);
nand U10639 (N_10639,N_8346,N_8167);
nand U10640 (N_10640,N_9838,N_9843);
or U10641 (N_10641,N_9389,N_8020);
nor U10642 (N_10642,N_9404,N_9970);
or U10643 (N_10643,N_8133,N_9524);
nor U10644 (N_10644,N_9194,N_9995);
xnor U10645 (N_10645,N_8697,N_9487);
and U10646 (N_10646,N_9783,N_8302);
nand U10647 (N_10647,N_9073,N_9329);
nor U10648 (N_10648,N_8114,N_8500);
and U10649 (N_10649,N_9205,N_8909);
xor U10650 (N_10650,N_8558,N_8937);
and U10651 (N_10651,N_8444,N_9748);
and U10652 (N_10652,N_9605,N_8534);
xnor U10653 (N_10653,N_8359,N_8275);
and U10654 (N_10654,N_9504,N_8288);
or U10655 (N_10655,N_8010,N_9493);
nand U10656 (N_10656,N_8617,N_8188);
nand U10657 (N_10657,N_8034,N_8548);
and U10658 (N_10658,N_9176,N_9562);
and U10659 (N_10659,N_9698,N_8499);
xnor U10660 (N_10660,N_9154,N_8964);
nor U10661 (N_10661,N_8896,N_9367);
or U10662 (N_10662,N_8916,N_9074);
nor U10663 (N_10663,N_8078,N_8827);
xnor U10664 (N_10664,N_8171,N_8520);
nor U10665 (N_10665,N_8823,N_8461);
nand U10666 (N_10666,N_9086,N_9191);
nor U10667 (N_10667,N_8842,N_9118);
nand U10668 (N_10668,N_9874,N_8059);
and U10669 (N_10669,N_9554,N_8391);
nor U10670 (N_10670,N_9723,N_9085);
xor U10671 (N_10671,N_8719,N_8123);
and U10672 (N_10672,N_9462,N_8420);
nor U10673 (N_10673,N_9102,N_8731);
nand U10674 (N_10674,N_9045,N_8878);
or U10675 (N_10675,N_9955,N_8780);
nor U10676 (N_10676,N_9359,N_8290);
or U10677 (N_10677,N_9919,N_8651);
or U10678 (N_10678,N_9123,N_9442);
nand U10679 (N_10679,N_8322,N_9592);
xor U10680 (N_10680,N_8639,N_8525);
nor U10681 (N_10681,N_9785,N_8014);
and U10682 (N_10682,N_9666,N_9886);
and U10683 (N_10683,N_9001,N_8603);
or U10684 (N_10684,N_9948,N_9157);
xnor U10685 (N_10685,N_9163,N_9742);
or U10686 (N_10686,N_8084,N_8879);
or U10687 (N_10687,N_8386,N_8271);
nand U10688 (N_10688,N_8561,N_8621);
xnor U10689 (N_10689,N_8399,N_9962);
xor U10690 (N_10690,N_8605,N_9663);
nand U10691 (N_10691,N_8062,N_9315);
and U10692 (N_10692,N_8362,N_9864);
nor U10693 (N_10693,N_9594,N_8324);
xor U10694 (N_10694,N_9243,N_9753);
nor U10695 (N_10695,N_8032,N_8165);
and U10696 (N_10696,N_9832,N_9913);
or U10697 (N_10697,N_9382,N_9553);
and U10698 (N_10698,N_9942,N_9903);
xnor U10699 (N_10699,N_8943,N_9934);
nor U10700 (N_10700,N_8316,N_9495);
or U10701 (N_10701,N_8929,N_8977);
nor U10702 (N_10702,N_8472,N_9759);
or U10703 (N_10703,N_9060,N_9964);
nand U10704 (N_10704,N_8379,N_8694);
nor U10705 (N_10705,N_8411,N_8199);
nor U10706 (N_10706,N_9907,N_9048);
xor U10707 (N_10707,N_9016,N_9760);
and U10708 (N_10708,N_9834,N_8931);
or U10709 (N_10709,N_8957,N_8351);
nor U10710 (N_10710,N_8335,N_8988);
nand U10711 (N_10711,N_8035,N_8243);
xor U10712 (N_10712,N_8319,N_9845);
nor U10713 (N_10713,N_9876,N_9652);
or U10714 (N_10714,N_9550,N_8642);
nand U10715 (N_10715,N_9113,N_9729);
xnor U10716 (N_10716,N_9358,N_8176);
xnor U10717 (N_10717,N_8108,N_8186);
xor U10718 (N_10718,N_8865,N_8222);
or U10719 (N_10719,N_9712,N_9837);
and U10720 (N_10720,N_8507,N_9988);
or U10721 (N_10721,N_8691,N_8388);
nand U10722 (N_10722,N_8025,N_8469);
or U10723 (N_10723,N_9122,N_8595);
or U10724 (N_10724,N_9828,N_8832);
nor U10725 (N_10725,N_8852,N_9522);
and U10726 (N_10726,N_9378,N_9944);
or U10727 (N_10727,N_9107,N_9418);
nand U10728 (N_10728,N_8637,N_9816);
xnor U10729 (N_10729,N_8655,N_8537);
or U10730 (N_10730,N_8674,N_8590);
nand U10731 (N_10731,N_8606,N_8301);
and U10732 (N_10732,N_9801,N_8913);
nor U10733 (N_10733,N_9114,N_9482);
or U10734 (N_10734,N_8416,N_9618);
xnor U10735 (N_10735,N_8624,N_9994);
or U10736 (N_10736,N_9987,N_8791);
xor U10737 (N_10737,N_8614,N_9240);
and U10738 (N_10738,N_8012,N_9588);
or U10739 (N_10739,N_8009,N_9849);
or U10740 (N_10740,N_8195,N_9559);
and U10741 (N_10741,N_8148,N_8524);
and U10742 (N_10742,N_8866,N_9992);
nand U10743 (N_10743,N_9568,N_9796);
nor U10744 (N_10744,N_9658,N_9897);
nand U10745 (N_10745,N_8779,N_9510);
and U10746 (N_10746,N_8063,N_8744);
and U10747 (N_10747,N_8881,N_9302);
or U10748 (N_10748,N_9285,N_8345);
and U10749 (N_10749,N_8070,N_9035);
nand U10750 (N_10750,N_9279,N_9277);
xor U10751 (N_10751,N_8094,N_8891);
nor U10752 (N_10752,N_9851,N_8600);
nand U10753 (N_10753,N_8099,N_8131);
nand U10754 (N_10754,N_8677,N_8609);
or U10755 (N_10755,N_8748,N_8789);
and U10756 (N_10756,N_8484,N_8545);
or U10757 (N_10757,N_8532,N_9246);
and U10758 (N_10758,N_8663,N_8200);
xor U10759 (N_10759,N_9545,N_8854);
or U10760 (N_10760,N_9427,N_8817);
and U10761 (N_10761,N_8255,N_8144);
or U10762 (N_10762,N_8482,N_8138);
and U10763 (N_10763,N_8299,N_8371);
and U10764 (N_10764,N_8671,N_9200);
or U10765 (N_10765,N_9262,N_8543);
nor U10766 (N_10766,N_8971,N_8082);
or U10767 (N_10767,N_8201,N_9403);
nor U10768 (N_10768,N_8267,N_8215);
nand U10769 (N_10769,N_9659,N_8975);
nand U10770 (N_10770,N_9465,N_8563);
nor U10771 (N_10771,N_9506,N_8460);
nand U10772 (N_10772,N_8057,N_8017);
and U10773 (N_10773,N_9508,N_9905);
xor U10774 (N_10774,N_8187,N_9108);
and U10775 (N_10775,N_9428,N_9862);
and U10776 (N_10776,N_8619,N_9983);
nor U10777 (N_10777,N_8326,N_8145);
or U10778 (N_10778,N_9368,N_9188);
nand U10779 (N_10779,N_9106,N_9178);
nor U10780 (N_10780,N_9662,N_9312);
or U10781 (N_10781,N_9668,N_8829);
nand U10782 (N_10782,N_8375,N_9400);
and U10783 (N_10783,N_8405,N_9142);
nand U10784 (N_10784,N_9611,N_9324);
or U10785 (N_10785,N_9399,N_8578);
and U10786 (N_10786,N_8464,N_8437);
and U10787 (N_10787,N_9936,N_8944);
and U10788 (N_10788,N_9763,N_9951);
or U10789 (N_10789,N_8997,N_8970);
nand U10790 (N_10790,N_8714,N_8278);
and U10791 (N_10791,N_8686,N_8608);
xor U10792 (N_10792,N_9884,N_9209);
nand U10793 (N_10793,N_8313,N_8917);
or U10794 (N_10794,N_8445,N_9471);
and U10795 (N_10795,N_9525,N_9061);
nand U10796 (N_10796,N_9604,N_9969);
xnor U10797 (N_10797,N_9069,N_8846);
xor U10798 (N_10798,N_9641,N_9310);
nor U10799 (N_10799,N_9719,N_9183);
nor U10800 (N_10800,N_9728,N_9199);
nor U10801 (N_10801,N_9543,N_9646);
nand U10802 (N_10802,N_8397,N_9159);
nor U10803 (N_10803,N_8421,N_8920);
or U10804 (N_10804,N_9640,N_8383);
nor U10805 (N_10805,N_8011,N_9943);
or U10806 (N_10806,N_9168,N_8649);
and U10807 (N_10807,N_9087,N_9772);
nand U10808 (N_10808,N_9591,N_9709);
or U10809 (N_10809,N_9249,N_8939);
nand U10810 (N_10810,N_9813,N_8533);
nor U10811 (N_10811,N_9637,N_9881);
nor U10812 (N_10812,N_8077,N_9920);
xor U10813 (N_10813,N_9511,N_9775);
nor U10814 (N_10814,N_9334,N_8317);
xor U10815 (N_10815,N_9872,N_9458);
nor U10816 (N_10816,N_8958,N_9678);
and U10817 (N_10817,N_9854,N_9004);
and U10818 (N_10818,N_8006,N_9475);
xor U10819 (N_10819,N_8475,N_9974);
and U10820 (N_10820,N_9043,N_8000);
xor U10821 (N_10821,N_9097,N_9132);
and U10822 (N_10822,N_9727,N_8826);
and U10823 (N_10823,N_8091,N_9797);
nand U10824 (N_10824,N_8620,N_9218);
xnor U10825 (N_10825,N_9693,N_8790);
and U10826 (N_10826,N_9056,N_9697);
nor U10827 (N_10827,N_8432,N_9137);
or U10828 (N_10828,N_9580,N_8272);
or U10829 (N_10829,N_9309,N_8887);
nor U10830 (N_10830,N_8352,N_9793);
or U10831 (N_10831,N_9755,N_9804);
or U10832 (N_10832,N_8007,N_8983);
nand U10833 (N_10833,N_9683,N_8522);
nand U10834 (N_10834,N_9509,N_9441);
nor U10835 (N_10835,N_8238,N_9468);
xor U10836 (N_10836,N_8659,N_9923);
or U10837 (N_10837,N_9771,N_9498);
xnor U10838 (N_10838,N_8076,N_8296);
or U10839 (N_10839,N_8298,N_8888);
and U10840 (N_10840,N_9397,N_9949);
or U10841 (N_10841,N_8064,N_9355);
or U10842 (N_10842,N_9620,N_8209);
nand U10843 (N_10843,N_9170,N_8068);
and U10844 (N_10844,N_9120,N_9058);
nand U10845 (N_10845,N_8247,N_9733);
nor U10846 (N_10846,N_9105,N_9973);
nand U10847 (N_10847,N_9651,N_8515);
and U10848 (N_10848,N_8938,N_9173);
and U10849 (N_10849,N_9353,N_9369);
or U10850 (N_10850,N_9877,N_8495);
and U10851 (N_10851,N_9921,N_8923);
nand U10852 (N_10852,N_8489,N_9501);
and U10853 (N_10853,N_9264,N_8205);
nor U10854 (N_10854,N_8075,N_9794);
nand U10855 (N_10855,N_9855,N_9732);
and U10856 (N_10856,N_8992,N_8936);
xor U10857 (N_10857,N_8841,N_8794);
xor U10858 (N_10858,N_9480,N_8729);
xor U10859 (N_10859,N_8924,N_8757);
nand U10860 (N_10860,N_9419,N_9997);
nand U10861 (N_10861,N_9383,N_8828);
nand U10862 (N_10862,N_8759,N_8395);
and U10863 (N_10863,N_8517,N_9959);
nor U10864 (N_10864,N_8287,N_8240);
nand U10865 (N_10865,N_8755,N_8259);
or U10866 (N_10866,N_9830,N_8274);
or U10867 (N_10867,N_9803,N_9928);
nor U10868 (N_10868,N_8152,N_9566);
or U10869 (N_10869,N_9883,N_8816);
xor U10870 (N_10870,N_9583,N_8111);
or U10871 (N_10871,N_9901,N_8945);
and U10872 (N_10872,N_9022,N_8061);
and U10873 (N_10873,N_9362,N_9076);
nand U10874 (N_10874,N_8367,N_8408);
or U10875 (N_10875,N_9181,N_8273);
nand U10876 (N_10876,N_8567,N_8280);
nor U10877 (N_10877,N_8203,N_8454);
nor U10878 (N_10878,N_9686,N_9317);
or U10879 (N_10879,N_9071,N_8392);
xnor U10880 (N_10880,N_8718,N_9549);
or U10881 (N_10881,N_8071,N_8633);
xor U10882 (N_10882,N_8002,N_8292);
and U10883 (N_10883,N_8085,N_8615);
nor U10884 (N_10884,N_8946,N_8429);
xor U10885 (N_10885,N_8797,N_8503);
and U10886 (N_10886,N_9560,N_9780);
and U10887 (N_10887,N_8055,N_8702);
or U10888 (N_10888,N_9587,N_8191);
and U10889 (N_10889,N_9616,N_9371);
nor U10890 (N_10890,N_8474,N_9072);
nor U10891 (N_10891,N_8874,N_8307);
nor U10892 (N_10892,N_8072,N_8087);
nand U10893 (N_10893,N_8253,N_8703);
and U10894 (N_10894,N_8998,N_8596);
and U10895 (N_10895,N_8178,N_8833);
nor U10896 (N_10896,N_9281,N_9846);
or U10897 (N_10897,N_9904,N_8546);
nand U10898 (N_10898,N_8083,N_8933);
nand U10899 (N_10899,N_9941,N_9866);
nand U10900 (N_10900,N_8369,N_8293);
or U10901 (N_10901,N_9051,N_8090);
nor U10902 (N_10902,N_9313,N_8216);
and U10903 (N_10903,N_8312,N_8582);
nor U10904 (N_10904,N_8672,N_8252);
nor U10905 (N_10905,N_8650,N_9922);
nor U10906 (N_10906,N_9459,N_8922);
or U10907 (N_10907,N_9228,N_9757);
nand U10908 (N_10908,N_8737,N_8591);
and U10909 (N_10909,N_9808,N_9840);
or U10910 (N_10910,N_8616,N_9961);
nor U10911 (N_10911,N_9293,N_9743);
nor U10912 (N_10912,N_8228,N_9751);
nand U10913 (N_10913,N_8115,N_8768);
nand U10914 (N_10914,N_8325,N_9245);
nor U10915 (N_10915,N_8043,N_8422);
and U10916 (N_10916,N_9826,N_8660);
nand U10917 (N_10917,N_8892,N_8493);
or U10918 (N_10918,N_8336,N_9164);
xor U10919 (N_10919,N_8248,N_8340);
nand U10920 (N_10920,N_8613,N_9967);
nand U10921 (N_10921,N_8506,N_8175);
and U10922 (N_10922,N_9481,N_8573);
and U10923 (N_10923,N_9625,N_9788);
and U10924 (N_10924,N_8549,N_9373);
xor U10925 (N_10925,N_9152,N_9489);
nor U10926 (N_10926,N_9347,N_8851);
xor U10927 (N_10927,N_8568,N_9385);
nand U10928 (N_10928,N_9681,N_8190);
or U10929 (N_10929,N_8738,N_8121);
or U10930 (N_10930,N_8565,N_9333);
xor U10931 (N_10931,N_9484,N_9675);
nand U10932 (N_10932,N_8196,N_9687);
and U10933 (N_10933,N_9207,N_8598);
nor U10934 (N_10934,N_8733,N_8769);
or U10935 (N_10935,N_9791,N_9255);
nor U10936 (N_10936,N_9252,N_9820);
and U10937 (N_10937,N_9950,N_8380);
and U10938 (N_10938,N_9224,N_8306);
or U10939 (N_10939,N_9349,N_9770);
and U10940 (N_10940,N_8968,N_9635);
or U10941 (N_10941,N_8294,N_8949);
nor U10942 (N_10942,N_8389,N_8806);
nor U10943 (N_10943,N_8539,N_8485);
and U10944 (N_10944,N_9366,N_8122);
and U10945 (N_10945,N_8900,N_8451);
xnor U10946 (N_10946,N_8556,N_8632);
or U10947 (N_10947,N_9784,N_8760);
and U10948 (N_10948,N_9778,N_9256);
nand U10949 (N_10949,N_8033,N_9280);
xor U10950 (N_10950,N_9055,N_9290);
xnor U10951 (N_10951,N_9746,N_9075);
nand U10952 (N_10952,N_8234,N_9824);
and U10953 (N_10953,N_8906,N_9272);
nand U10954 (N_10954,N_9565,N_8330);
and U10955 (N_10955,N_9439,N_8610);
xnor U10956 (N_10956,N_8370,N_8783);
nor U10957 (N_10957,N_8740,N_8724);
or U10958 (N_10958,N_9754,N_8626);
nand U10959 (N_10959,N_9953,N_8743);
nand U10960 (N_10960,N_9270,N_8118);
nor U10961 (N_10961,N_9265,N_9889);
nand U10962 (N_10962,N_8103,N_8095);
nand U10963 (N_10963,N_8344,N_8762);
nor U10964 (N_10964,N_9940,N_8955);
and U10965 (N_10965,N_8956,N_8695);
and U10966 (N_10966,N_9494,N_8251);
nand U10967 (N_10967,N_9722,N_8683);
nor U10968 (N_10968,N_8623,N_9689);
or U10969 (N_10969,N_8800,N_8830);
nor U10970 (N_10970,N_9469,N_8811);
nor U10971 (N_10971,N_9119,N_9467);
nor U10972 (N_10972,N_8726,N_8715);
or U10973 (N_10973,N_9331,N_8004);
or U10974 (N_10974,N_9610,N_8747);
nand U10975 (N_10975,N_8311,N_8704);
or U10976 (N_10976,N_9372,N_9063);
nand U10977 (N_10977,N_9747,N_8348);
and U10978 (N_10978,N_8985,N_9847);
and U10979 (N_10979,N_9274,N_8709);
nand U10980 (N_10980,N_9037,N_9147);
xor U10981 (N_10981,N_9337,N_8926);
xor U10982 (N_10982,N_9014,N_8635);
nand U10983 (N_10983,N_9082,N_8870);
xor U10984 (N_10984,N_8692,N_8113);
nand U10985 (N_10985,N_8867,N_8227);
nand U10986 (N_10986,N_8229,N_8679);
nand U10987 (N_10987,N_8776,N_9645);
nand U10988 (N_10988,N_8690,N_8310);
nor U10989 (N_10989,N_8712,N_9623);
and U10990 (N_10990,N_8557,N_8571);
xor U10991 (N_10991,N_8749,N_8969);
xor U10992 (N_10992,N_9965,N_9332);
xor U10993 (N_10993,N_8984,N_9835);
xor U10994 (N_10994,N_8696,N_8457);
nand U10995 (N_10995,N_8911,N_8182);
nor U10996 (N_10996,N_9148,N_9810);
nand U10997 (N_10997,N_8277,N_9189);
or U10998 (N_10998,N_9574,N_8538);
nor U10999 (N_10999,N_9429,N_9806);
or U11000 (N_11000,N_8499,N_8484);
nand U11001 (N_11001,N_8926,N_8922);
nor U11002 (N_11002,N_9435,N_9664);
nor U11003 (N_11003,N_9860,N_8411);
nor U11004 (N_11004,N_8054,N_8438);
or U11005 (N_11005,N_8387,N_9642);
or U11006 (N_11006,N_9427,N_9570);
nor U11007 (N_11007,N_8408,N_9853);
xnor U11008 (N_11008,N_8939,N_9609);
nand U11009 (N_11009,N_9098,N_8912);
nor U11010 (N_11010,N_9556,N_8168);
and U11011 (N_11011,N_8619,N_8769);
or U11012 (N_11012,N_9246,N_8741);
nand U11013 (N_11013,N_9487,N_8372);
nor U11014 (N_11014,N_8907,N_9732);
xor U11015 (N_11015,N_9438,N_9842);
xor U11016 (N_11016,N_9730,N_8634);
nor U11017 (N_11017,N_9329,N_9914);
and U11018 (N_11018,N_9225,N_9350);
and U11019 (N_11019,N_8650,N_9582);
or U11020 (N_11020,N_9256,N_8722);
xnor U11021 (N_11021,N_9742,N_8584);
nand U11022 (N_11022,N_8899,N_9550);
xnor U11023 (N_11023,N_8535,N_9592);
nand U11024 (N_11024,N_9708,N_8063);
or U11025 (N_11025,N_8180,N_8688);
or U11026 (N_11026,N_9274,N_8043);
nand U11027 (N_11027,N_8887,N_8481);
nor U11028 (N_11028,N_9632,N_9108);
xnor U11029 (N_11029,N_9167,N_8268);
nor U11030 (N_11030,N_9975,N_9234);
nor U11031 (N_11031,N_9474,N_8835);
xnor U11032 (N_11032,N_9012,N_9983);
and U11033 (N_11033,N_9927,N_9185);
and U11034 (N_11034,N_8359,N_8956);
xnor U11035 (N_11035,N_9618,N_8940);
and U11036 (N_11036,N_8267,N_8641);
or U11037 (N_11037,N_9615,N_9033);
xnor U11038 (N_11038,N_8457,N_8196);
xnor U11039 (N_11039,N_9854,N_9800);
nand U11040 (N_11040,N_8035,N_8422);
xor U11041 (N_11041,N_9023,N_8485);
nand U11042 (N_11042,N_8980,N_9158);
nor U11043 (N_11043,N_8850,N_9699);
nor U11044 (N_11044,N_9667,N_8851);
nand U11045 (N_11045,N_9578,N_8777);
xnor U11046 (N_11046,N_8391,N_8083);
xnor U11047 (N_11047,N_9287,N_8928);
and U11048 (N_11048,N_9748,N_9396);
xor U11049 (N_11049,N_9993,N_9165);
xnor U11050 (N_11050,N_8658,N_8288);
and U11051 (N_11051,N_9737,N_9620);
or U11052 (N_11052,N_8077,N_9654);
nor U11053 (N_11053,N_8715,N_9693);
nand U11054 (N_11054,N_9961,N_8148);
nand U11055 (N_11055,N_8637,N_9358);
and U11056 (N_11056,N_8400,N_8164);
or U11057 (N_11057,N_9311,N_9268);
and U11058 (N_11058,N_9594,N_8201);
nor U11059 (N_11059,N_8019,N_9713);
nand U11060 (N_11060,N_8044,N_9780);
and U11061 (N_11061,N_9729,N_8799);
and U11062 (N_11062,N_8738,N_9927);
nand U11063 (N_11063,N_9740,N_8755);
nor U11064 (N_11064,N_9680,N_9354);
nand U11065 (N_11065,N_9830,N_9504);
nor U11066 (N_11066,N_8185,N_8024);
or U11067 (N_11067,N_8595,N_8544);
and U11068 (N_11068,N_9203,N_8110);
nor U11069 (N_11069,N_8264,N_9387);
and U11070 (N_11070,N_8468,N_8133);
or U11071 (N_11071,N_9590,N_9106);
nand U11072 (N_11072,N_8305,N_8472);
xor U11073 (N_11073,N_9550,N_8857);
nand U11074 (N_11074,N_8637,N_9641);
or U11075 (N_11075,N_8545,N_9455);
or U11076 (N_11076,N_8150,N_8235);
nor U11077 (N_11077,N_9404,N_8207);
nor U11078 (N_11078,N_8019,N_8197);
nor U11079 (N_11079,N_8072,N_9694);
or U11080 (N_11080,N_9920,N_9272);
nand U11081 (N_11081,N_8716,N_8139);
nand U11082 (N_11082,N_8089,N_9198);
or U11083 (N_11083,N_9587,N_8411);
xnor U11084 (N_11084,N_9342,N_8158);
or U11085 (N_11085,N_9316,N_9325);
xnor U11086 (N_11086,N_8289,N_8167);
xnor U11087 (N_11087,N_8591,N_8892);
xnor U11088 (N_11088,N_8698,N_8285);
or U11089 (N_11089,N_8335,N_8703);
nand U11090 (N_11090,N_9601,N_8345);
nor U11091 (N_11091,N_8381,N_9346);
xor U11092 (N_11092,N_9830,N_9474);
and U11093 (N_11093,N_8673,N_9738);
or U11094 (N_11094,N_9861,N_9852);
or U11095 (N_11095,N_8282,N_8991);
and U11096 (N_11096,N_8765,N_9818);
or U11097 (N_11097,N_8983,N_8448);
xnor U11098 (N_11098,N_9261,N_9694);
xnor U11099 (N_11099,N_8150,N_8192);
nor U11100 (N_11100,N_9683,N_9934);
nand U11101 (N_11101,N_9325,N_9982);
nor U11102 (N_11102,N_9221,N_8805);
and U11103 (N_11103,N_8453,N_8236);
or U11104 (N_11104,N_8229,N_8028);
nand U11105 (N_11105,N_8553,N_9168);
and U11106 (N_11106,N_8543,N_9877);
nor U11107 (N_11107,N_8537,N_9473);
xnor U11108 (N_11108,N_8360,N_9357);
or U11109 (N_11109,N_9633,N_8613);
nor U11110 (N_11110,N_8339,N_9826);
or U11111 (N_11111,N_8897,N_9102);
nor U11112 (N_11112,N_8620,N_8419);
and U11113 (N_11113,N_8983,N_8705);
xor U11114 (N_11114,N_9393,N_9404);
nor U11115 (N_11115,N_9864,N_9466);
xor U11116 (N_11116,N_9048,N_8152);
xnor U11117 (N_11117,N_8837,N_8431);
and U11118 (N_11118,N_8025,N_9089);
or U11119 (N_11119,N_8764,N_8879);
and U11120 (N_11120,N_8222,N_9608);
or U11121 (N_11121,N_9391,N_9112);
and U11122 (N_11122,N_9605,N_9395);
xor U11123 (N_11123,N_8928,N_9368);
nor U11124 (N_11124,N_8926,N_8149);
nand U11125 (N_11125,N_9877,N_8122);
or U11126 (N_11126,N_9215,N_8228);
or U11127 (N_11127,N_8291,N_8964);
nand U11128 (N_11128,N_8943,N_9424);
and U11129 (N_11129,N_9028,N_8538);
and U11130 (N_11130,N_9278,N_8492);
nor U11131 (N_11131,N_8232,N_8017);
or U11132 (N_11132,N_8532,N_9005);
or U11133 (N_11133,N_8553,N_8157);
or U11134 (N_11134,N_8737,N_9132);
or U11135 (N_11135,N_9669,N_8294);
nor U11136 (N_11136,N_8515,N_8405);
or U11137 (N_11137,N_9413,N_8591);
nand U11138 (N_11138,N_9995,N_8759);
xor U11139 (N_11139,N_9704,N_8546);
xnor U11140 (N_11140,N_8850,N_8887);
and U11141 (N_11141,N_8919,N_9325);
or U11142 (N_11142,N_9806,N_9224);
xor U11143 (N_11143,N_9598,N_9861);
and U11144 (N_11144,N_9999,N_8783);
nand U11145 (N_11145,N_8499,N_9451);
xnor U11146 (N_11146,N_8181,N_9847);
and U11147 (N_11147,N_8507,N_8315);
or U11148 (N_11148,N_9291,N_8225);
nor U11149 (N_11149,N_9523,N_9548);
nor U11150 (N_11150,N_9533,N_8091);
xnor U11151 (N_11151,N_9601,N_8869);
and U11152 (N_11152,N_8211,N_9850);
or U11153 (N_11153,N_8910,N_9589);
and U11154 (N_11154,N_8855,N_9975);
and U11155 (N_11155,N_9560,N_9255);
or U11156 (N_11156,N_9278,N_8237);
or U11157 (N_11157,N_9532,N_8180);
nand U11158 (N_11158,N_8515,N_9373);
nand U11159 (N_11159,N_9269,N_8460);
nor U11160 (N_11160,N_8482,N_9655);
xor U11161 (N_11161,N_8209,N_9400);
nand U11162 (N_11162,N_8694,N_9523);
and U11163 (N_11163,N_9040,N_9513);
xor U11164 (N_11164,N_8255,N_8317);
and U11165 (N_11165,N_8954,N_8829);
xnor U11166 (N_11166,N_8872,N_8442);
nor U11167 (N_11167,N_8521,N_8441);
nor U11168 (N_11168,N_8817,N_8076);
xor U11169 (N_11169,N_8200,N_8391);
or U11170 (N_11170,N_8608,N_8865);
nor U11171 (N_11171,N_9081,N_9913);
nor U11172 (N_11172,N_8056,N_8994);
nand U11173 (N_11173,N_9840,N_8888);
or U11174 (N_11174,N_8485,N_8687);
nor U11175 (N_11175,N_8853,N_8781);
or U11176 (N_11176,N_9825,N_8566);
and U11177 (N_11177,N_8626,N_8466);
or U11178 (N_11178,N_8331,N_8815);
nor U11179 (N_11179,N_9111,N_8011);
and U11180 (N_11180,N_9226,N_9775);
and U11181 (N_11181,N_9144,N_8943);
and U11182 (N_11182,N_9729,N_9960);
xor U11183 (N_11183,N_8295,N_9121);
xnor U11184 (N_11184,N_9984,N_9216);
xor U11185 (N_11185,N_8445,N_9324);
xor U11186 (N_11186,N_9458,N_9295);
nand U11187 (N_11187,N_8364,N_8472);
xnor U11188 (N_11188,N_9520,N_8599);
nor U11189 (N_11189,N_9898,N_8910);
and U11190 (N_11190,N_8639,N_8954);
xor U11191 (N_11191,N_9568,N_9537);
nor U11192 (N_11192,N_8909,N_8765);
and U11193 (N_11193,N_9790,N_9230);
nand U11194 (N_11194,N_8789,N_9031);
or U11195 (N_11195,N_9145,N_8554);
and U11196 (N_11196,N_8938,N_9984);
and U11197 (N_11197,N_9769,N_8604);
and U11198 (N_11198,N_8424,N_8067);
or U11199 (N_11199,N_8282,N_9119);
xor U11200 (N_11200,N_9473,N_9507);
and U11201 (N_11201,N_8787,N_8272);
xnor U11202 (N_11202,N_8236,N_8450);
xor U11203 (N_11203,N_8436,N_8876);
or U11204 (N_11204,N_8984,N_9560);
nor U11205 (N_11205,N_8062,N_8513);
and U11206 (N_11206,N_9945,N_8400);
and U11207 (N_11207,N_8609,N_9449);
and U11208 (N_11208,N_9497,N_9717);
nor U11209 (N_11209,N_9569,N_9347);
nand U11210 (N_11210,N_8343,N_8788);
xor U11211 (N_11211,N_9539,N_9633);
xor U11212 (N_11212,N_8591,N_9598);
and U11213 (N_11213,N_9539,N_8908);
or U11214 (N_11214,N_9794,N_8039);
and U11215 (N_11215,N_8711,N_9010);
xor U11216 (N_11216,N_8834,N_8809);
and U11217 (N_11217,N_8669,N_8636);
nor U11218 (N_11218,N_9253,N_8468);
or U11219 (N_11219,N_8645,N_9728);
or U11220 (N_11220,N_9822,N_9744);
or U11221 (N_11221,N_8236,N_8944);
and U11222 (N_11222,N_8247,N_9017);
xor U11223 (N_11223,N_8833,N_8676);
and U11224 (N_11224,N_8701,N_8562);
or U11225 (N_11225,N_8989,N_9614);
or U11226 (N_11226,N_9036,N_8658);
and U11227 (N_11227,N_8856,N_9278);
and U11228 (N_11228,N_9797,N_9245);
xor U11229 (N_11229,N_9020,N_9226);
xnor U11230 (N_11230,N_8130,N_9295);
and U11231 (N_11231,N_8922,N_9015);
and U11232 (N_11232,N_8474,N_9065);
xnor U11233 (N_11233,N_9836,N_8028);
nand U11234 (N_11234,N_9088,N_9899);
nand U11235 (N_11235,N_9667,N_9459);
xnor U11236 (N_11236,N_9820,N_9817);
or U11237 (N_11237,N_8622,N_9856);
xor U11238 (N_11238,N_9483,N_9429);
or U11239 (N_11239,N_9451,N_8184);
nand U11240 (N_11240,N_8675,N_9599);
nor U11241 (N_11241,N_8096,N_8943);
nor U11242 (N_11242,N_8824,N_8328);
xor U11243 (N_11243,N_9252,N_9120);
and U11244 (N_11244,N_8091,N_9635);
xor U11245 (N_11245,N_8126,N_8782);
nand U11246 (N_11246,N_9934,N_8506);
nor U11247 (N_11247,N_8968,N_8579);
xor U11248 (N_11248,N_8344,N_9836);
or U11249 (N_11249,N_8350,N_9509);
and U11250 (N_11250,N_9069,N_8245);
xnor U11251 (N_11251,N_9215,N_8784);
nand U11252 (N_11252,N_8342,N_8306);
or U11253 (N_11253,N_8937,N_9439);
nor U11254 (N_11254,N_8897,N_9912);
nor U11255 (N_11255,N_8625,N_8389);
xnor U11256 (N_11256,N_9196,N_9289);
nor U11257 (N_11257,N_8890,N_8472);
xor U11258 (N_11258,N_9952,N_8944);
nor U11259 (N_11259,N_9611,N_9658);
xnor U11260 (N_11260,N_9693,N_8558);
nand U11261 (N_11261,N_9784,N_9945);
nor U11262 (N_11262,N_8770,N_9299);
and U11263 (N_11263,N_8364,N_9290);
nand U11264 (N_11264,N_9152,N_8947);
or U11265 (N_11265,N_9058,N_9923);
xnor U11266 (N_11266,N_8650,N_9077);
nor U11267 (N_11267,N_8101,N_9305);
nor U11268 (N_11268,N_9723,N_8406);
and U11269 (N_11269,N_8801,N_8912);
nand U11270 (N_11270,N_9816,N_9785);
nand U11271 (N_11271,N_8938,N_8970);
or U11272 (N_11272,N_9226,N_9677);
nor U11273 (N_11273,N_8339,N_8024);
xor U11274 (N_11274,N_8910,N_9488);
or U11275 (N_11275,N_8370,N_9297);
or U11276 (N_11276,N_9111,N_9198);
nor U11277 (N_11277,N_8634,N_9431);
xor U11278 (N_11278,N_9072,N_8324);
nand U11279 (N_11279,N_8128,N_8107);
nor U11280 (N_11280,N_9682,N_8837);
or U11281 (N_11281,N_9686,N_9460);
or U11282 (N_11282,N_8971,N_9798);
or U11283 (N_11283,N_8517,N_9525);
nor U11284 (N_11284,N_8317,N_9792);
nor U11285 (N_11285,N_9272,N_8239);
nand U11286 (N_11286,N_8041,N_8704);
nor U11287 (N_11287,N_8536,N_9231);
nor U11288 (N_11288,N_8297,N_9285);
nand U11289 (N_11289,N_9295,N_8581);
nand U11290 (N_11290,N_8006,N_8674);
or U11291 (N_11291,N_8657,N_8941);
nand U11292 (N_11292,N_9884,N_9335);
and U11293 (N_11293,N_8065,N_8209);
xor U11294 (N_11294,N_9593,N_8273);
nor U11295 (N_11295,N_9506,N_8983);
or U11296 (N_11296,N_8172,N_8744);
and U11297 (N_11297,N_8677,N_8994);
nand U11298 (N_11298,N_8676,N_9885);
and U11299 (N_11299,N_8900,N_8435);
and U11300 (N_11300,N_9610,N_8106);
xor U11301 (N_11301,N_9027,N_9496);
nand U11302 (N_11302,N_8561,N_8323);
nand U11303 (N_11303,N_8261,N_8834);
and U11304 (N_11304,N_9338,N_9154);
nand U11305 (N_11305,N_9326,N_9796);
nand U11306 (N_11306,N_8498,N_9290);
or U11307 (N_11307,N_9632,N_9356);
and U11308 (N_11308,N_9490,N_9321);
nand U11309 (N_11309,N_8528,N_9760);
or U11310 (N_11310,N_9956,N_9205);
and U11311 (N_11311,N_8940,N_8971);
nor U11312 (N_11312,N_9011,N_8470);
xor U11313 (N_11313,N_8289,N_8408);
and U11314 (N_11314,N_9805,N_8731);
and U11315 (N_11315,N_9525,N_9625);
nor U11316 (N_11316,N_9678,N_9987);
and U11317 (N_11317,N_8339,N_8566);
nand U11318 (N_11318,N_9975,N_9010);
nor U11319 (N_11319,N_9454,N_9035);
nor U11320 (N_11320,N_9196,N_8610);
or U11321 (N_11321,N_9951,N_9671);
and U11322 (N_11322,N_8171,N_8597);
xnor U11323 (N_11323,N_9833,N_8207);
or U11324 (N_11324,N_8294,N_8881);
xnor U11325 (N_11325,N_8833,N_9582);
nor U11326 (N_11326,N_8889,N_8829);
xor U11327 (N_11327,N_8810,N_8846);
nor U11328 (N_11328,N_8335,N_9271);
nor U11329 (N_11329,N_9822,N_8841);
xnor U11330 (N_11330,N_8255,N_8191);
or U11331 (N_11331,N_8935,N_9967);
and U11332 (N_11332,N_8778,N_9705);
or U11333 (N_11333,N_8157,N_8495);
and U11334 (N_11334,N_9077,N_9594);
or U11335 (N_11335,N_8453,N_8294);
xor U11336 (N_11336,N_9904,N_8486);
or U11337 (N_11337,N_8553,N_9294);
or U11338 (N_11338,N_8389,N_9862);
xor U11339 (N_11339,N_9961,N_9371);
and U11340 (N_11340,N_8164,N_8099);
xor U11341 (N_11341,N_9627,N_9712);
and U11342 (N_11342,N_8040,N_8454);
and U11343 (N_11343,N_8778,N_9057);
xor U11344 (N_11344,N_8480,N_9570);
nor U11345 (N_11345,N_8219,N_8046);
nor U11346 (N_11346,N_9197,N_8805);
and U11347 (N_11347,N_8410,N_9527);
nor U11348 (N_11348,N_8654,N_8854);
nand U11349 (N_11349,N_8011,N_8101);
xor U11350 (N_11350,N_9392,N_8512);
nand U11351 (N_11351,N_9292,N_8991);
and U11352 (N_11352,N_8169,N_8313);
or U11353 (N_11353,N_9846,N_9373);
nand U11354 (N_11354,N_8664,N_9190);
nand U11355 (N_11355,N_9465,N_9174);
nand U11356 (N_11356,N_8554,N_9294);
nand U11357 (N_11357,N_9187,N_8317);
nand U11358 (N_11358,N_8197,N_9624);
or U11359 (N_11359,N_8532,N_8517);
xnor U11360 (N_11360,N_9833,N_8281);
nand U11361 (N_11361,N_9790,N_8668);
nor U11362 (N_11362,N_8396,N_9249);
nor U11363 (N_11363,N_9679,N_9619);
nor U11364 (N_11364,N_9344,N_8340);
or U11365 (N_11365,N_8242,N_9548);
nor U11366 (N_11366,N_8249,N_9048);
nor U11367 (N_11367,N_8408,N_8180);
nor U11368 (N_11368,N_9259,N_8044);
and U11369 (N_11369,N_8634,N_8384);
or U11370 (N_11370,N_9034,N_8770);
nor U11371 (N_11371,N_9921,N_8335);
or U11372 (N_11372,N_9005,N_9361);
or U11373 (N_11373,N_9312,N_9886);
and U11374 (N_11374,N_8939,N_8868);
or U11375 (N_11375,N_8497,N_9880);
nand U11376 (N_11376,N_9047,N_8405);
and U11377 (N_11377,N_8774,N_9921);
or U11378 (N_11378,N_8276,N_9264);
and U11379 (N_11379,N_8572,N_8591);
and U11380 (N_11380,N_8016,N_9645);
nor U11381 (N_11381,N_9448,N_9554);
nand U11382 (N_11382,N_8772,N_8448);
or U11383 (N_11383,N_8461,N_8949);
or U11384 (N_11384,N_8314,N_9364);
xnor U11385 (N_11385,N_9183,N_8828);
or U11386 (N_11386,N_8646,N_9610);
and U11387 (N_11387,N_8217,N_8042);
and U11388 (N_11388,N_9256,N_8509);
and U11389 (N_11389,N_9038,N_9613);
nand U11390 (N_11390,N_9379,N_9857);
or U11391 (N_11391,N_8827,N_9443);
and U11392 (N_11392,N_8915,N_8467);
nor U11393 (N_11393,N_9372,N_8979);
nand U11394 (N_11394,N_8346,N_9629);
nand U11395 (N_11395,N_8842,N_9942);
or U11396 (N_11396,N_9184,N_9199);
or U11397 (N_11397,N_9235,N_8796);
nor U11398 (N_11398,N_8510,N_9456);
or U11399 (N_11399,N_9359,N_9871);
or U11400 (N_11400,N_8608,N_8044);
xor U11401 (N_11401,N_9449,N_9214);
nand U11402 (N_11402,N_9431,N_8025);
or U11403 (N_11403,N_9251,N_9750);
and U11404 (N_11404,N_9991,N_9387);
nand U11405 (N_11405,N_8726,N_9272);
or U11406 (N_11406,N_9489,N_8771);
nand U11407 (N_11407,N_8824,N_8224);
nor U11408 (N_11408,N_9048,N_8902);
nand U11409 (N_11409,N_8558,N_8191);
or U11410 (N_11410,N_8176,N_9936);
and U11411 (N_11411,N_9941,N_8780);
or U11412 (N_11412,N_8079,N_8715);
nor U11413 (N_11413,N_9882,N_8567);
xnor U11414 (N_11414,N_9179,N_8076);
or U11415 (N_11415,N_8448,N_8417);
nand U11416 (N_11416,N_9447,N_9966);
and U11417 (N_11417,N_9280,N_8415);
and U11418 (N_11418,N_8425,N_8954);
nand U11419 (N_11419,N_8888,N_9527);
nor U11420 (N_11420,N_9904,N_8652);
and U11421 (N_11421,N_9670,N_9081);
or U11422 (N_11422,N_9252,N_9603);
and U11423 (N_11423,N_9395,N_8418);
nand U11424 (N_11424,N_8117,N_9601);
nand U11425 (N_11425,N_8283,N_8465);
or U11426 (N_11426,N_9788,N_9884);
nor U11427 (N_11427,N_8845,N_9846);
or U11428 (N_11428,N_8389,N_8521);
and U11429 (N_11429,N_9922,N_8677);
nor U11430 (N_11430,N_9285,N_9733);
nor U11431 (N_11431,N_9671,N_9405);
or U11432 (N_11432,N_9953,N_8776);
nor U11433 (N_11433,N_9719,N_8524);
and U11434 (N_11434,N_8204,N_8996);
or U11435 (N_11435,N_9636,N_9076);
or U11436 (N_11436,N_8850,N_8576);
or U11437 (N_11437,N_9198,N_8929);
nor U11438 (N_11438,N_8338,N_9759);
nand U11439 (N_11439,N_8623,N_8239);
nor U11440 (N_11440,N_8053,N_8628);
nor U11441 (N_11441,N_9546,N_9885);
nand U11442 (N_11442,N_8017,N_9759);
and U11443 (N_11443,N_8896,N_8902);
or U11444 (N_11444,N_8323,N_8650);
nand U11445 (N_11445,N_9646,N_8143);
and U11446 (N_11446,N_8661,N_9300);
or U11447 (N_11447,N_8668,N_8671);
nand U11448 (N_11448,N_9186,N_9961);
nor U11449 (N_11449,N_8593,N_8975);
nand U11450 (N_11450,N_8542,N_9045);
nor U11451 (N_11451,N_9785,N_8634);
nand U11452 (N_11452,N_9292,N_9206);
nor U11453 (N_11453,N_8434,N_8019);
nor U11454 (N_11454,N_9979,N_8200);
and U11455 (N_11455,N_9297,N_8014);
xnor U11456 (N_11456,N_9545,N_8238);
nor U11457 (N_11457,N_8817,N_9988);
xnor U11458 (N_11458,N_8450,N_9060);
nand U11459 (N_11459,N_8863,N_8591);
nor U11460 (N_11460,N_9185,N_9705);
nor U11461 (N_11461,N_8353,N_8506);
nor U11462 (N_11462,N_8406,N_9221);
nand U11463 (N_11463,N_8480,N_9550);
and U11464 (N_11464,N_9580,N_9023);
nand U11465 (N_11465,N_9856,N_8837);
nand U11466 (N_11466,N_8403,N_8158);
and U11467 (N_11467,N_9040,N_9527);
and U11468 (N_11468,N_9017,N_8288);
xnor U11469 (N_11469,N_8460,N_9406);
or U11470 (N_11470,N_9626,N_8023);
nor U11471 (N_11471,N_8728,N_9058);
and U11472 (N_11472,N_9978,N_9727);
and U11473 (N_11473,N_9004,N_8615);
xor U11474 (N_11474,N_9656,N_8383);
and U11475 (N_11475,N_8777,N_8541);
nand U11476 (N_11476,N_9178,N_8582);
nor U11477 (N_11477,N_8449,N_9459);
nand U11478 (N_11478,N_9944,N_8719);
nor U11479 (N_11479,N_9819,N_9939);
xnor U11480 (N_11480,N_9011,N_8278);
or U11481 (N_11481,N_9514,N_8780);
nand U11482 (N_11482,N_9548,N_9345);
or U11483 (N_11483,N_8018,N_8557);
nor U11484 (N_11484,N_9461,N_8462);
nor U11485 (N_11485,N_9420,N_9861);
nor U11486 (N_11486,N_8505,N_8018);
nand U11487 (N_11487,N_9113,N_9649);
or U11488 (N_11488,N_8345,N_8918);
nand U11489 (N_11489,N_9384,N_8518);
nand U11490 (N_11490,N_9010,N_9232);
xnor U11491 (N_11491,N_8595,N_8790);
nor U11492 (N_11492,N_8733,N_8358);
and U11493 (N_11493,N_8178,N_9746);
or U11494 (N_11494,N_9243,N_9541);
nand U11495 (N_11495,N_9040,N_8397);
and U11496 (N_11496,N_9116,N_8735);
nor U11497 (N_11497,N_8141,N_9987);
or U11498 (N_11498,N_9560,N_8451);
or U11499 (N_11499,N_8671,N_9041);
nand U11500 (N_11500,N_9611,N_8016);
nor U11501 (N_11501,N_8066,N_8652);
and U11502 (N_11502,N_9169,N_8077);
xnor U11503 (N_11503,N_9400,N_9747);
xnor U11504 (N_11504,N_9902,N_8226);
nor U11505 (N_11505,N_8250,N_9910);
and U11506 (N_11506,N_9764,N_8165);
nand U11507 (N_11507,N_8457,N_8280);
nor U11508 (N_11508,N_9151,N_8519);
nor U11509 (N_11509,N_8632,N_9226);
or U11510 (N_11510,N_9536,N_8692);
nand U11511 (N_11511,N_9272,N_9571);
xnor U11512 (N_11512,N_9298,N_8261);
xor U11513 (N_11513,N_8251,N_8416);
xnor U11514 (N_11514,N_8844,N_8884);
xor U11515 (N_11515,N_8155,N_9599);
nand U11516 (N_11516,N_9365,N_8155);
nand U11517 (N_11517,N_8178,N_9211);
nor U11518 (N_11518,N_8640,N_9014);
and U11519 (N_11519,N_8394,N_9805);
and U11520 (N_11520,N_8327,N_8802);
nor U11521 (N_11521,N_8201,N_8109);
nor U11522 (N_11522,N_8568,N_9987);
xor U11523 (N_11523,N_9923,N_8790);
or U11524 (N_11524,N_8118,N_9766);
nor U11525 (N_11525,N_9715,N_8984);
nand U11526 (N_11526,N_9247,N_8550);
and U11527 (N_11527,N_9689,N_8669);
xor U11528 (N_11528,N_8148,N_9613);
nor U11529 (N_11529,N_9474,N_9217);
nor U11530 (N_11530,N_8638,N_9046);
nand U11531 (N_11531,N_9581,N_9095);
nand U11532 (N_11532,N_8150,N_9590);
or U11533 (N_11533,N_9269,N_8009);
xnor U11534 (N_11534,N_8035,N_9536);
or U11535 (N_11535,N_9301,N_8296);
nand U11536 (N_11536,N_8914,N_8245);
nor U11537 (N_11537,N_9536,N_9711);
nand U11538 (N_11538,N_9330,N_8882);
xnor U11539 (N_11539,N_9895,N_9741);
or U11540 (N_11540,N_9636,N_9864);
xor U11541 (N_11541,N_9333,N_8229);
xnor U11542 (N_11542,N_9886,N_9255);
nand U11543 (N_11543,N_9980,N_9907);
xor U11544 (N_11544,N_8752,N_9402);
nor U11545 (N_11545,N_9496,N_8405);
nor U11546 (N_11546,N_9504,N_8881);
or U11547 (N_11547,N_9129,N_9895);
nand U11548 (N_11548,N_9947,N_9185);
xor U11549 (N_11549,N_8134,N_9254);
nor U11550 (N_11550,N_8976,N_8122);
nor U11551 (N_11551,N_9775,N_9021);
xor U11552 (N_11552,N_8314,N_9972);
xor U11553 (N_11553,N_8019,N_8807);
or U11554 (N_11554,N_8366,N_9928);
or U11555 (N_11555,N_8300,N_8843);
nand U11556 (N_11556,N_8175,N_9577);
and U11557 (N_11557,N_9933,N_8411);
xor U11558 (N_11558,N_8787,N_9512);
nor U11559 (N_11559,N_9694,N_9616);
and U11560 (N_11560,N_8438,N_9168);
xor U11561 (N_11561,N_8854,N_9658);
nor U11562 (N_11562,N_9974,N_8022);
xnor U11563 (N_11563,N_9339,N_8591);
nand U11564 (N_11564,N_9840,N_8370);
and U11565 (N_11565,N_9420,N_8574);
and U11566 (N_11566,N_8896,N_9183);
or U11567 (N_11567,N_8172,N_8174);
nor U11568 (N_11568,N_8828,N_9973);
nand U11569 (N_11569,N_9760,N_9789);
nand U11570 (N_11570,N_8505,N_8487);
nand U11571 (N_11571,N_9953,N_8171);
or U11572 (N_11572,N_9430,N_9540);
or U11573 (N_11573,N_8100,N_8265);
nor U11574 (N_11574,N_9914,N_8095);
or U11575 (N_11575,N_9105,N_9722);
nand U11576 (N_11576,N_9755,N_9079);
or U11577 (N_11577,N_8660,N_9485);
nor U11578 (N_11578,N_8029,N_9507);
or U11579 (N_11579,N_9001,N_8055);
nor U11580 (N_11580,N_8127,N_9749);
and U11581 (N_11581,N_9996,N_9247);
or U11582 (N_11582,N_9467,N_9826);
xor U11583 (N_11583,N_8546,N_8024);
xor U11584 (N_11584,N_9813,N_9162);
or U11585 (N_11585,N_8201,N_9409);
nor U11586 (N_11586,N_8215,N_9129);
nor U11587 (N_11587,N_8954,N_8103);
or U11588 (N_11588,N_8068,N_9540);
xnor U11589 (N_11589,N_9899,N_8922);
nor U11590 (N_11590,N_9748,N_8833);
or U11591 (N_11591,N_9570,N_8634);
and U11592 (N_11592,N_9596,N_8639);
or U11593 (N_11593,N_8940,N_9541);
xor U11594 (N_11594,N_9675,N_9912);
or U11595 (N_11595,N_8310,N_8182);
xnor U11596 (N_11596,N_8468,N_9602);
or U11597 (N_11597,N_8453,N_8262);
nor U11598 (N_11598,N_8436,N_9880);
and U11599 (N_11599,N_8036,N_8312);
nor U11600 (N_11600,N_9763,N_8439);
nand U11601 (N_11601,N_8697,N_9971);
and U11602 (N_11602,N_9755,N_9631);
or U11603 (N_11603,N_8121,N_8511);
xnor U11604 (N_11604,N_9663,N_8509);
nand U11605 (N_11605,N_8498,N_9516);
nor U11606 (N_11606,N_8957,N_9522);
nand U11607 (N_11607,N_9291,N_8535);
and U11608 (N_11608,N_8775,N_9908);
and U11609 (N_11609,N_8671,N_9313);
nor U11610 (N_11610,N_8262,N_8490);
and U11611 (N_11611,N_9474,N_8108);
xnor U11612 (N_11612,N_9990,N_9400);
xnor U11613 (N_11613,N_8615,N_8394);
and U11614 (N_11614,N_8167,N_9892);
and U11615 (N_11615,N_8374,N_9610);
or U11616 (N_11616,N_9482,N_8843);
and U11617 (N_11617,N_9495,N_8707);
nor U11618 (N_11618,N_9710,N_8292);
nand U11619 (N_11619,N_8489,N_8259);
and U11620 (N_11620,N_9513,N_8982);
xor U11621 (N_11621,N_8038,N_9667);
nor U11622 (N_11622,N_8680,N_9200);
or U11623 (N_11623,N_9757,N_9537);
nand U11624 (N_11624,N_9130,N_9951);
nor U11625 (N_11625,N_8401,N_9196);
or U11626 (N_11626,N_9110,N_8200);
xor U11627 (N_11627,N_9794,N_9546);
nor U11628 (N_11628,N_8633,N_8854);
nor U11629 (N_11629,N_8677,N_8660);
nor U11630 (N_11630,N_9632,N_9113);
nand U11631 (N_11631,N_8757,N_9065);
nand U11632 (N_11632,N_8819,N_9320);
nor U11633 (N_11633,N_8359,N_9220);
and U11634 (N_11634,N_9531,N_9106);
xnor U11635 (N_11635,N_8601,N_8517);
nor U11636 (N_11636,N_8252,N_8777);
nor U11637 (N_11637,N_9660,N_8180);
nor U11638 (N_11638,N_8973,N_9016);
nand U11639 (N_11639,N_8975,N_8432);
or U11640 (N_11640,N_9805,N_9407);
or U11641 (N_11641,N_9036,N_9629);
and U11642 (N_11642,N_8615,N_9490);
or U11643 (N_11643,N_9175,N_9365);
nor U11644 (N_11644,N_9978,N_8329);
nor U11645 (N_11645,N_8054,N_8529);
nor U11646 (N_11646,N_8911,N_8019);
or U11647 (N_11647,N_9112,N_8067);
and U11648 (N_11648,N_9715,N_9328);
nor U11649 (N_11649,N_8681,N_8595);
xnor U11650 (N_11650,N_9961,N_9859);
nand U11651 (N_11651,N_8449,N_9217);
nand U11652 (N_11652,N_9247,N_9210);
and U11653 (N_11653,N_9762,N_9825);
nor U11654 (N_11654,N_8629,N_8979);
or U11655 (N_11655,N_8221,N_8192);
nand U11656 (N_11656,N_9210,N_8843);
nand U11657 (N_11657,N_9194,N_9815);
or U11658 (N_11658,N_8599,N_8921);
xor U11659 (N_11659,N_9564,N_9980);
nor U11660 (N_11660,N_9030,N_9701);
xor U11661 (N_11661,N_8858,N_8221);
and U11662 (N_11662,N_9062,N_8631);
nor U11663 (N_11663,N_9254,N_9423);
and U11664 (N_11664,N_8700,N_8110);
and U11665 (N_11665,N_9029,N_8085);
nand U11666 (N_11666,N_9875,N_9261);
nor U11667 (N_11667,N_9747,N_9349);
or U11668 (N_11668,N_9132,N_9251);
xor U11669 (N_11669,N_9405,N_8076);
xnor U11670 (N_11670,N_8203,N_8774);
nand U11671 (N_11671,N_9737,N_8508);
and U11672 (N_11672,N_9116,N_9216);
and U11673 (N_11673,N_9725,N_9388);
xnor U11674 (N_11674,N_8208,N_8322);
nand U11675 (N_11675,N_8781,N_9017);
and U11676 (N_11676,N_9543,N_8318);
xnor U11677 (N_11677,N_9952,N_9059);
xor U11678 (N_11678,N_8804,N_9629);
or U11679 (N_11679,N_8265,N_9134);
or U11680 (N_11680,N_8104,N_9269);
or U11681 (N_11681,N_8627,N_8280);
and U11682 (N_11682,N_8922,N_8967);
and U11683 (N_11683,N_8879,N_8813);
nand U11684 (N_11684,N_9190,N_8675);
xor U11685 (N_11685,N_9948,N_8168);
xor U11686 (N_11686,N_9949,N_9728);
nor U11687 (N_11687,N_8291,N_8683);
xor U11688 (N_11688,N_9082,N_9648);
nor U11689 (N_11689,N_9491,N_9197);
nand U11690 (N_11690,N_8950,N_9606);
or U11691 (N_11691,N_8117,N_9315);
or U11692 (N_11692,N_8382,N_9702);
and U11693 (N_11693,N_8060,N_8220);
or U11694 (N_11694,N_8814,N_8640);
nand U11695 (N_11695,N_8313,N_8816);
and U11696 (N_11696,N_9221,N_8875);
xnor U11697 (N_11697,N_8096,N_8200);
nor U11698 (N_11698,N_8533,N_8467);
or U11699 (N_11699,N_9161,N_8782);
and U11700 (N_11700,N_8653,N_8188);
xor U11701 (N_11701,N_9573,N_8332);
xor U11702 (N_11702,N_9429,N_8646);
or U11703 (N_11703,N_9174,N_8304);
and U11704 (N_11704,N_8789,N_9776);
or U11705 (N_11705,N_8372,N_8823);
xor U11706 (N_11706,N_8876,N_8523);
nand U11707 (N_11707,N_8887,N_8574);
nand U11708 (N_11708,N_9319,N_8287);
nand U11709 (N_11709,N_9554,N_8817);
xnor U11710 (N_11710,N_8291,N_9991);
nand U11711 (N_11711,N_9004,N_8981);
nand U11712 (N_11712,N_8346,N_8149);
nand U11713 (N_11713,N_8147,N_8708);
xor U11714 (N_11714,N_9774,N_9578);
xnor U11715 (N_11715,N_9684,N_9437);
or U11716 (N_11716,N_9370,N_8071);
or U11717 (N_11717,N_8089,N_8469);
nand U11718 (N_11718,N_8037,N_9295);
nor U11719 (N_11719,N_8965,N_9018);
and U11720 (N_11720,N_8632,N_8575);
nand U11721 (N_11721,N_9461,N_9436);
nand U11722 (N_11722,N_8132,N_8325);
nand U11723 (N_11723,N_9191,N_9516);
nand U11724 (N_11724,N_9724,N_8895);
and U11725 (N_11725,N_8150,N_8016);
nor U11726 (N_11726,N_9696,N_9303);
nand U11727 (N_11727,N_8773,N_8438);
and U11728 (N_11728,N_8064,N_8673);
nand U11729 (N_11729,N_9960,N_9317);
nand U11730 (N_11730,N_9854,N_9362);
or U11731 (N_11731,N_9378,N_8481);
nand U11732 (N_11732,N_9587,N_8703);
nand U11733 (N_11733,N_9925,N_8845);
xor U11734 (N_11734,N_9307,N_8376);
and U11735 (N_11735,N_8582,N_9163);
nand U11736 (N_11736,N_8771,N_9867);
or U11737 (N_11737,N_9967,N_9189);
and U11738 (N_11738,N_9863,N_9256);
and U11739 (N_11739,N_9508,N_9691);
or U11740 (N_11740,N_8281,N_8988);
nand U11741 (N_11741,N_9803,N_9321);
or U11742 (N_11742,N_9835,N_8172);
nand U11743 (N_11743,N_9953,N_8357);
xor U11744 (N_11744,N_8737,N_8134);
and U11745 (N_11745,N_8325,N_8408);
and U11746 (N_11746,N_8801,N_8948);
xor U11747 (N_11747,N_9319,N_9013);
nor U11748 (N_11748,N_9343,N_8434);
and U11749 (N_11749,N_9911,N_9228);
nor U11750 (N_11750,N_9874,N_9861);
or U11751 (N_11751,N_8260,N_8973);
and U11752 (N_11752,N_8411,N_8424);
nor U11753 (N_11753,N_9975,N_9737);
xor U11754 (N_11754,N_8513,N_9625);
xor U11755 (N_11755,N_8116,N_8171);
and U11756 (N_11756,N_9618,N_8971);
and U11757 (N_11757,N_8587,N_9652);
or U11758 (N_11758,N_8539,N_8965);
nor U11759 (N_11759,N_8655,N_9732);
and U11760 (N_11760,N_9362,N_8438);
xor U11761 (N_11761,N_9732,N_8595);
nand U11762 (N_11762,N_8224,N_9553);
or U11763 (N_11763,N_8215,N_8862);
or U11764 (N_11764,N_8650,N_9508);
or U11765 (N_11765,N_8175,N_9134);
nand U11766 (N_11766,N_9129,N_8216);
nand U11767 (N_11767,N_8878,N_9208);
nand U11768 (N_11768,N_9987,N_8561);
nand U11769 (N_11769,N_8463,N_9365);
and U11770 (N_11770,N_9002,N_9826);
nor U11771 (N_11771,N_8047,N_9802);
and U11772 (N_11772,N_8350,N_9525);
nand U11773 (N_11773,N_9934,N_9872);
nor U11774 (N_11774,N_8673,N_8328);
nor U11775 (N_11775,N_8768,N_8756);
and U11776 (N_11776,N_9140,N_8420);
xnor U11777 (N_11777,N_8844,N_8630);
and U11778 (N_11778,N_9223,N_8102);
nand U11779 (N_11779,N_8342,N_8366);
nor U11780 (N_11780,N_8267,N_8388);
and U11781 (N_11781,N_9756,N_9587);
xnor U11782 (N_11782,N_9420,N_8176);
nand U11783 (N_11783,N_8738,N_8158);
nor U11784 (N_11784,N_8661,N_9692);
xor U11785 (N_11785,N_9514,N_9361);
and U11786 (N_11786,N_8058,N_9373);
or U11787 (N_11787,N_8363,N_9943);
and U11788 (N_11788,N_8595,N_9015);
xnor U11789 (N_11789,N_8321,N_8764);
xor U11790 (N_11790,N_9073,N_8327);
and U11791 (N_11791,N_8879,N_8824);
and U11792 (N_11792,N_9788,N_9434);
xnor U11793 (N_11793,N_8244,N_8161);
nor U11794 (N_11794,N_9794,N_9058);
and U11795 (N_11795,N_8135,N_8743);
nor U11796 (N_11796,N_9625,N_8314);
xor U11797 (N_11797,N_8812,N_9247);
and U11798 (N_11798,N_9792,N_9021);
nor U11799 (N_11799,N_9821,N_9700);
and U11800 (N_11800,N_9081,N_9037);
nor U11801 (N_11801,N_9784,N_8708);
and U11802 (N_11802,N_8060,N_9252);
nand U11803 (N_11803,N_9129,N_8923);
and U11804 (N_11804,N_8412,N_8389);
nand U11805 (N_11805,N_8056,N_8755);
xnor U11806 (N_11806,N_9810,N_9167);
xor U11807 (N_11807,N_9726,N_9945);
xor U11808 (N_11808,N_9236,N_8915);
xor U11809 (N_11809,N_9856,N_9402);
nand U11810 (N_11810,N_8755,N_9661);
nand U11811 (N_11811,N_9739,N_8801);
and U11812 (N_11812,N_8402,N_8439);
nor U11813 (N_11813,N_9953,N_9932);
and U11814 (N_11814,N_9670,N_9276);
nor U11815 (N_11815,N_9386,N_8415);
xnor U11816 (N_11816,N_8760,N_9503);
nor U11817 (N_11817,N_8457,N_8020);
and U11818 (N_11818,N_9814,N_8867);
xor U11819 (N_11819,N_8144,N_8753);
nand U11820 (N_11820,N_8957,N_9683);
and U11821 (N_11821,N_9375,N_8323);
and U11822 (N_11822,N_8786,N_8126);
and U11823 (N_11823,N_8068,N_8974);
xnor U11824 (N_11824,N_9263,N_9792);
nand U11825 (N_11825,N_8732,N_9115);
or U11826 (N_11826,N_9056,N_9439);
or U11827 (N_11827,N_8907,N_9300);
xor U11828 (N_11828,N_9980,N_9592);
or U11829 (N_11829,N_8602,N_8768);
xnor U11830 (N_11830,N_9110,N_9824);
and U11831 (N_11831,N_9473,N_8266);
and U11832 (N_11832,N_9563,N_8260);
or U11833 (N_11833,N_8379,N_9781);
nand U11834 (N_11834,N_8911,N_9115);
nand U11835 (N_11835,N_9976,N_9749);
and U11836 (N_11836,N_8916,N_9318);
nor U11837 (N_11837,N_8611,N_8777);
nor U11838 (N_11838,N_8326,N_8098);
or U11839 (N_11839,N_9284,N_9582);
xnor U11840 (N_11840,N_9419,N_8017);
xor U11841 (N_11841,N_8388,N_9344);
nand U11842 (N_11842,N_9912,N_9698);
and U11843 (N_11843,N_8589,N_8756);
nand U11844 (N_11844,N_8045,N_9347);
or U11845 (N_11845,N_8254,N_8410);
nand U11846 (N_11846,N_8308,N_8153);
xor U11847 (N_11847,N_9230,N_8517);
xor U11848 (N_11848,N_8450,N_9461);
nor U11849 (N_11849,N_8449,N_8400);
nand U11850 (N_11850,N_8938,N_8281);
xor U11851 (N_11851,N_9620,N_9029);
or U11852 (N_11852,N_9451,N_9366);
and U11853 (N_11853,N_9730,N_9463);
xor U11854 (N_11854,N_9467,N_9680);
or U11855 (N_11855,N_8191,N_8157);
nand U11856 (N_11856,N_8049,N_9054);
nand U11857 (N_11857,N_8770,N_9076);
and U11858 (N_11858,N_9728,N_8731);
xnor U11859 (N_11859,N_9198,N_9552);
nand U11860 (N_11860,N_9094,N_8822);
and U11861 (N_11861,N_9901,N_9627);
nor U11862 (N_11862,N_9478,N_8637);
or U11863 (N_11863,N_9326,N_8721);
or U11864 (N_11864,N_8265,N_9509);
or U11865 (N_11865,N_9560,N_8219);
nand U11866 (N_11866,N_9451,N_9901);
xor U11867 (N_11867,N_8674,N_9388);
xor U11868 (N_11868,N_8971,N_9198);
nor U11869 (N_11869,N_8937,N_8562);
nand U11870 (N_11870,N_9265,N_9583);
or U11871 (N_11871,N_8561,N_9882);
and U11872 (N_11872,N_8718,N_8315);
and U11873 (N_11873,N_9246,N_9754);
nor U11874 (N_11874,N_8997,N_8183);
or U11875 (N_11875,N_9968,N_9452);
or U11876 (N_11876,N_8450,N_9919);
xor U11877 (N_11877,N_9698,N_8660);
xor U11878 (N_11878,N_9566,N_8775);
or U11879 (N_11879,N_9675,N_8562);
xnor U11880 (N_11880,N_8532,N_8244);
and U11881 (N_11881,N_8744,N_9152);
or U11882 (N_11882,N_8191,N_9129);
xnor U11883 (N_11883,N_9595,N_8201);
xnor U11884 (N_11884,N_9456,N_9712);
and U11885 (N_11885,N_9195,N_8998);
xor U11886 (N_11886,N_8364,N_9878);
nor U11887 (N_11887,N_8537,N_8626);
nand U11888 (N_11888,N_8978,N_8961);
or U11889 (N_11889,N_8881,N_9600);
xor U11890 (N_11890,N_8859,N_8298);
nand U11891 (N_11891,N_9717,N_8036);
xnor U11892 (N_11892,N_9472,N_8380);
and U11893 (N_11893,N_8529,N_9220);
nand U11894 (N_11894,N_9197,N_8752);
and U11895 (N_11895,N_9421,N_8273);
nand U11896 (N_11896,N_9188,N_8597);
nand U11897 (N_11897,N_8127,N_9962);
nand U11898 (N_11898,N_9398,N_8262);
and U11899 (N_11899,N_8396,N_8933);
nor U11900 (N_11900,N_8638,N_8360);
or U11901 (N_11901,N_8837,N_9059);
or U11902 (N_11902,N_8583,N_8304);
nor U11903 (N_11903,N_9039,N_8556);
or U11904 (N_11904,N_9023,N_8659);
xor U11905 (N_11905,N_9164,N_9577);
xor U11906 (N_11906,N_8807,N_8869);
nor U11907 (N_11907,N_8580,N_8643);
nor U11908 (N_11908,N_9126,N_8146);
xor U11909 (N_11909,N_8396,N_9348);
xor U11910 (N_11910,N_9228,N_8056);
nor U11911 (N_11911,N_9815,N_8372);
xnor U11912 (N_11912,N_8585,N_9605);
nor U11913 (N_11913,N_8972,N_9678);
and U11914 (N_11914,N_8897,N_8307);
xnor U11915 (N_11915,N_8851,N_9275);
xor U11916 (N_11916,N_9537,N_8187);
and U11917 (N_11917,N_9321,N_9829);
nand U11918 (N_11918,N_8467,N_8128);
or U11919 (N_11919,N_9448,N_8019);
and U11920 (N_11920,N_9364,N_8629);
and U11921 (N_11921,N_9373,N_8899);
or U11922 (N_11922,N_8400,N_9689);
nand U11923 (N_11923,N_8044,N_9300);
and U11924 (N_11924,N_9046,N_9548);
nand U11925 (N_11925,N_8964,N_9364);
xnor U11926 (N_11926,N_8440,N_8664);
nor U11927 (N_11927,N_8592,N_9477);
nor U11928 (N_11928,N_8372,N_8618);
and U11929 (N_11929,N_8501,N_9187);
xnor U11930 (N_11930,N_8071,N_9204);
xnor U11931 (N_11931,N_9240,N_9979);
nand U11932 (N_11932,N_8653,N_9504);
nand U11933 (N_11933,N_8932,N_8475);
nand U11934 (N_11934,N_8107,N_9501);
nand U11935 (N_11935,N_9138,N_8669);
or U11936 (N_11936,N_9256,N_9713);
and U11937 (N_11937,N_8623,N_9604);
xor U11938 (N_11938,N_9287,N_8041);
nor U11939 (N_11939,N_9896,N_8787);
nor U11940 (N_11940,N_9838,N_9867);
xnor U11941 (N_11941,N_8039,N_8482);
and U11942 (N_11942,N_9771,N_8954);
and U11943 (N_11943,N_8054,N_9310);
xor U11944 (N_11944,N_9428,N_9232);
nand U11945 (N_11945,N_8378,N_8561);
xnor U11946 (N_11946,N_8041,N_8475);
xor U11947 (N_11947,N_9941,N_8732);
nand U11948 (N_11948,N_8601,N_8342);
xor U11949 (N_11949,N_8843,N_8766);
xnor U11950 (N_11950,N_9239,N_9478);
and U11951 (N_11951,N_8964,N_9670);
and U11952 (N_11952,N_9366,N_9965);
nand U11953 (N_11953,N_8288,N_9443);
or U11954 (N_11954,N_8556,N_9936);
or U11955 (N_11955,N_9402,N_8942);
or U11956 (N_11956,N_8766,N_9852);
nand U11957 (N_11957,N_8049,N_8216);
or U11958 (N_11958,N_8821,N_9455);
and U11959 (N_11959,N_8699,N_9300);
nor U11960 (N_11960,N_8652,N_9496);
xor U11961 (N_11961,N_8289,N_9539);
nor U11962 (N_11962,N_9333,N_9219);
or U11963 (N_11963,N_8016,N_9756);
xor U11964 (N_11964,N_9984,N_9421);
nand U11965 (N_11965,N_8494,N_9357);
xor U11966 (N_11966,N_8704,N_8042);
or U11967 (N_11967,N_8978,N_9135);
nand U11968 (N_11968,N_9481,N_8199);
nand U11969 (N_11969,N_8279,N_8395);
or U11970 (N_11970,N_9627,N_9127);
or U11971 (N_11971,N_8803,N_8296);
xor U11972 (N_11972,N_8676,N_9127);
nand U11973 (N_11973,N_8531,N_8856);
and U11974 (N_11974,N_8794,N_8754);
xnor U11975 (N_11975,N_9742,N_9574);
or U11976 (N_11976,N_9451,N_9780);
xor U11977 (N_11977,N_8766,N_8297);
nor U11978 (N_11978,N_9708,N_9183);
nand U11979 (N_11979,N_8897,N_8848);
and U11980 (N_11980,N_9665,N_8869);
or U11981 (N_11981,N_9526,N_8390);
nor U11982 (N_11982,N_8382,N_9311);
nor U11983 (N_11983,N_9368,N_9308);
nand U11984 (N_11984,N_8862,N_9083);
nor U11985 (N_11985,N_9857,N_8433);
nor U11986 (N_11986,N_8219,N_9278);
or U11987 (N_11987,N_8609,N_9557);
or U11988 (N_11988,N_8375,N_8486);
and U11989 (N_11989,N_8947,N_9295);
nand U11990 (N_11990,N_9498,N_9083);
nand U11991 (N_11991,N_8283,N_8268);
xnor U11992 (N_11992,N_9506,N_8338);
nor U11993 (N_11993,N_9079,N_9500);
nor U11994 (N_11994,N_8791,N_8837);
or U11995 (N_11995,N_8826,N_9021);
xnor U11996 (N_11996,N_8356,N_8603);
nor U11997 (N_11997,N_8051,N_9730);
nor U11998 (N_11998,N_9184,N_9851);
or U11999 (N_11999,N_9673,N_9032);
nor U12000 (N_12000,N_11963,N_11055);
xnor U12001 (N_12001,N_10943,N_10548);
nor U12002 (N_12002,N_10065,N_10610);
nor U12003 (N_12003,N_11500,N_11159);
nor U12004 (N_12004,N_11077,N_10727);
nand U12005 (N_12005,N_10921,N_10929);
nand U12006 (N_12006,N_11929,N_11796);
nand U12007 (N_12007,N_11848,N_10939);
nor U12008 (N_12008,N_10718,N_11653);
nor U12009 (N_12009,N_10607,N_10177);
or U12010 (N_12010,N_10864,N_10379);
or U12011 (N_12011,N_11805,N_10699);
xnor U12012 (N_12012,N_10017,N_10170);
nand U12013 (N_12013,N_11187,N_11285);
nand U12014 (N_12014,N_11001,N_10638);
xor U12015 (N_12015,N_11383,N_11844);
nand U12016 (N_12016,N_11105,N_10658);
nand U12017 (N_12017,N_10028,N_11063);
nor U12018 (N_12018,N_11329,N_11302);
xnor U12019 (N_12019,N_10164,N_11817);
nor U12020 (N_12020,N_11346,N_10537);
nand U12021 (N_12021,N_11059,N_11238);
nor U12022 (N_12022,N_10119,N_11111);
xnor U12023 (N_12023,N_10267,N_10873);
nor U12024 (N_12024,N_10215,N_11171);
and U12025 (N_12025,N_11135,N_11969);
or U12026 (N_12026,N_10687,N_10226);
xnor U12027 (N_12027,N_10971,N_11153);
or U12028 (N_12028,N_11126,N_10994);
nand U12029 (N_12029,N_11470,N_10577);
xnor U12030 (N_12030,N_10905,N_10397);
xor U12031 (N_12031,N_11377,N_10644);
or U12032 (N_12032,N_11981,N_10214);
xor U12033 (N_12033,N_10458,N_10573);
xor U12034 (N_12034,N_10280,N_10269);
or U12035 (N_12035,N_11116,N_10315);
and U12036 (N_12036,N_11635,N_11403);
nand U12037 (N_12037,N_10796,N_10591);
or U12038 (N_12038,N_10098,N_11795);
nor U12039 (N_12039,N_11754,N_10775);
nand U12040 (N_12040,N_10179,N_10138);
nand U12041 (N_12041,N_11032,N_11737);
or U12042 (N_12042,N_11104,N_11511);
or U12043 (N_12043,N_11473,N_11599);
xnor U12044 (N_12044,N_11909,N_11519);
nand U12045 (N_12045,N_10886,N_10843);
xor U12046 (N_12046,N_11832,N_10750);
nor U12047 (N_12047,N_10744,N_11785);
nor U12048 (N_12048,N_10472,N_10195);
xnor U12049 (N_12049,N_11657,N_10307);
xnor U12050 (N_12050,N_11193,N_11529);
or U12051 (N_12051,N_11988,N_11647);
and U12052 (N_12052,N_11751,N_11531);
nor U12053 (N_12053,N_10211,N_10925);
nor U12054 (N_12054,N_10033,N_10813);
xor U12055 (N_12055,N_10163,N_10764);
or U12056 (N_12056,N_11348,N_10355);
xnor U12057 (N_12057,N_11043,N_11660);
or U12058 (N_12058,N_11125,N_11094);
and U12059 (N_12059,N_11337,N_10774);
and U12060 (N_12060,N_11025,N_11300);
and U12061 (N_12061,N_10575,N_11184);
nor U12062 (N_12062,N_10358,N_11971);
xor U12063 (N_12063,N_10451,N_10767);
nand U12064 (N_12064,N_11405,N_11062);
nand U12065 (N_12065,N_10833,N_11334);
nor U12066 (N_12066,N_10975,N_11281);
xnor U12067 (N_12067,N_10474,N_10229);
and U12068 (N_12068,N_10790,N_10456);
nor U12069 (N_12069,N_11974,N_10639);
xor U12070 (N_12070,N_11080,N_10159);
nand U12071 (N_12071,N_10869,N_11525);
nand U12072 (N_12072,N_10522,N_10538);
or U12073 (N_12073,N_11752,N_11290);
nand U12074 (N_12074,N_11219,N_10192);
nand U12075 (N_12075,N_10719,N_11609);
xnor U12076 (N_12076,N_10627,N_11864);
nand U12077 (N_12077,N_10129,N_11740);
nor U12078 (N_12078,N_10189,N_11940);
nand U12079 (N_12079,N_11052,N_11645);
nand U12080 (N_12080,N_11205,N_11937);
nor U12081 (N_12081,N_10212,N_11449);
nor U12082 (N_12082,N_11393,N_10361);
or U12083 (N_12083,N_11007,N_11333);
nand U12084 (N_12084,N_10983,N_11030);
nand U12085 (N_12085,N_10853,N_11252);
and U12086 (N_12086,N_11692,N_10672);
nand U12087 (N_12087,N_10679,N_11389);
xor U12088 (N_12088,N_10590,N_10419);
or U12089 (N_12089,N_11360,N_10623);
nor U12090 (N_12090,N_10407,N_10807);
nand U12091 (N_12091,N_10093,N_11150);
nand U12092 (N_12092,N_11227,N_11624);
xnor U12093 (N_12093,N_10025,N_10301);
nand U12094 (N_12094,N_10225,N_11666);
and U12095 (N_12095,N_11424,N_11565);
or U12096 (N_12096,N_10915,N_11115);
xor U12097 (N_12097,N_10231,N_11398);
or U12098 (N_12098,N_11671,N_11308);
nand U12099 (N_12099,N_11327,N_10675);
nor U12100 (N_12100,N_11190,N_10913);
nand U12101 (N_12101,N_11890,N_10768);
xor U12102 (N_12102,N_11761,N_11769);
nand U12103 (N_12103,N_11908,N_11201);
nand U12104 (N_12104,N_10064,N_11270);
xnor U12105 (N_12105,N_11841,N_10359);
and U12106 (N_12106,N_11092,N_10333);
xnor U12107 (N_12107,N_10842,N_10586);
and U12108 (N_12108,N_10297,N_10115);
and U12109 (N_12109,N_11467,N_11699);
nor U12110 (N_12110,N_11901,N_10081);
xor U12111 (N_12111,N_10092,N_11358);
xnor U12112 (N_12112,N_11408,N_10514);
nor U12113 (N_12113,N_10141,N_11475);
nand U12114 (N_12114,N_10977,N_11090);
and U12115 (N_12115,N_11873,N_10688);
and U12116 (N_12116,N_10665,N_10165);
nor U12117 (N_12117,N_10048,N_10637);
nor U12118 (N_12118,N_11233,N_10283);
nand U12119 (N_12119,N_10186,N_11605);
nor U12120 (N_12120,N_10726,N_10266);
nor U12121 (N_12121,N_10061,N_10636);
and U12122 (N_12122,N_10336,N_11556);
nand U12123 (N_12123,N_10659,N_11717);
nor U12124 (N_12124,N_10166,N_10128);
and U12125 (N_12125,N_10576,N_11416);
or U12126 (N_12126,N_10872,N_11222);
nor U12127 (N_12127,N_11324,N_10454);
nand U12128 (N_12128,N_11939,N_11876);
nand U12129 (N_12129,N_11048,N_10912);
nor U12130 (N_12130,N_11464,N_10888);
xnor U12131 (N_12131,N_11878,N_11382);
nand U12132 (N_12132,N_10695,N_10681);
xor U12133 (N_12133,N_11418,N_10715);
and U12134 (N_12134,N_10782,N_11808);
nand U12135 (N_12135,N_10376,N_10097);
nand U12136 (N_12136,N_10278,N_11573);
or U12137 (N_12137,N_10530,N_11085);
or U12138 (N_12138,N_11232,N_10292);
nor U12139 (N_12139,N_11916,N_11679);
nor U12140 (N_12140,N_10752,N_11102);
nand U12141 (N_12141,N_10019,N_11231);
and U12142 (N_12142,N_11894,N_10208);
and U12143 (N_12143,N_10470,N_11698);
nor U12144 (N_12144,N_11522,N_10222);
or U12145 (N_12145,N_10001,N_10331);
nand U12146 (N_12146,N_11654,N_10818);
xor U12147 (N_12147,N_11513,N_11203);
and U12148 (N_12148,N_10228,N_11774);
and U12149 (N_12149,N_11581,N_10550);
xnor U12150 (N_12150,N_10820,N_10467);
or U12151 (N_12151,N_10367,N_11716);
nand U12152 (N_12152,N_10256,N_11545);
and U12153 (N_12153,N_10452,N_11828);
xnor U12154 (N_12154,N_10776,N_11443);
xnor U12155 (N_12155,N_11613,N_10340);
nor U12156 (N_12156,N_10370,N_11258);
or U12157 (N_12157,N_10363,N_11496);
nand U12158 (N_12158,N_10520,N_11026);
xnor U12159 (N_12159,N_11093,N_10892);
nor U12160 (N_12160,N_11668,N_11306);
xor U12161 (N_12161,N_10007,N_11378);
xor U12162 (N_12162,N_11978,N_10196);
nor U12163 (N_12163,N_10809,N_10043);
and U12164 (N_12164,N_11180,N_10249);
nor U12165 (N_12165,N_11441,N_10987);
or U12166 (N_12166,N_11775,N_11476);
and U12167 (N_12167,N_10260,N_11049);
nand U12168 (N_12168,N_11585,N_11217);
and U12169 (N_12169,N_11975,N_10717);
nor U12170 (N_12170,N_10733,N_10923);
xnor U12171 (N_12171,N_11594,N_11409);
nand U12172 (N_12172,N_11835,N_10410);
nor U12173 (N_12173,N_10890,N_10594);
xor U12174 (N_12174,N_10974,N_11607);
nor U12175 (N_12175,N_10145,N_11355);
nor U12176 (N_12176,N_11788,N_10360);
xor U12177 (N_12177,N_11365,N_10383);
xor U12178 (N_12178,N_10124,N_11081);
and U12179 (N_12179,N_11945,N_11993);
or U12180 (N_12180,N_10626,N_10748);
nand U12181 (N_12181,N_11154,N_11315);
xor U12182 (N_12182,N_11215,N_10600);
nor U12183 (N_12183,N_11955,N_11784);
nand U12184 (N_12184,N_11938,N_10277);
and U12185 (N_12185,N_11492,N_11065);
nor U12186 (N_12186,N_10111,N_11206);
and U12187 (N_12187,N_11162,N_10499);
nor U12188 (N_12188,N_11709,N_10982);
and U12189 (N_12189,N_11713,N_10797);
xor U12190 (N_12190,N_11843,N_10227);
nand U12191 (N_12191,N_11028,N_11675);
xor U12192 (N_12192,N_11182,N_10749);
nand U12193 (N_12193,N_11818,N_11721);
nand U12194 (N_12194,N_10587,N_11568);
xnor U12195 (N_12195,N_10347,N_10692);
xor U12196 (N_12196,N_11626,N_10757);
or U12197 (N_12197,N_10123,N_10711);
or U12198 (N_12198,N_10099,N_11847);
and U12199 (N_12199,N_11319,N_10896);
nand U12200 (N_12200,N_10830,N_10992);
nand U12201 (N_12201,N_10816,N_10944);
or U12202 (N_12202,N_10691,N_10349);
nor U12203 (N_12203,N_10246,N_10544);
nand U12204 (N_12204,N_11623,N_10188);
and U12205 (N_12205,N_11794,N_10485);
nor U12206 (N_12206,N_10209,N_10435);
nor U12207 (N_12207,N_11046,N_10200);
nand U12208 (N_12208,N_10051,N_10369);
nand U12209 (N_12209,N_10673,N_10285);
xnor U12210 (N_12210,N_11905,N_10935);
nand U12211 (N_12211,N_11330,N_10684);
or U12212 (N_12212,N_10054,N_11875);
nor U12213 (N_12213,N_11619,N_10420);
nand U12214 (N_12214,N_10908,N_10066);
or U12215 (N_12215,N_10362,N_10385);
nor U12216 (N_12216,N_10042,N_11682);
xnor U12217 (N_12217,N_11935,N_11286);
nand U12218 (N_12218,N_11584,N_11830);
nor U12219 (N_12219,N_11447,N_10493);
and U12220 (N_12220,N_10318,N_11764);
and U12221 (N_12221,N_10402,N_11413);
or U12222 (N_12222,N_11574,N_10766);
or U12223 (N_12223,N_10022,N_10161);
and U12224 (N_12224,N_11865,N_11107);
or U12225 (N_12225,N_10941,N_10068);
nand U12226 (N_12226,N_10494,N_10745);
and U12227 (N_12227,N_10063,N_11851);
or U12228 (N_12228,N_11690,N_10965);
nand U12229 (N_12229,N_10381,N_11350);
and U12230 (N_12230,N_11820,N_10479);
and U12231 (N_12231,N_10605,N_10265);
xor U12232 (N_12232,N_10657,N_11490);
and U12233 (N_12233,N_11780,N_10069);
nor U12234 (N_12234,N_11601,N_11461);
and U12235 (N_12235,N_11806,N_10233);
nand U12236 (N_12236,N_10176,N_10505);
nor U12237 (N_12237,N_11108,N_11210);
nand U12238 (N_12238,N_10107,N_10940);
xor U12239 (N_12239,N_11741,N_11960);
xnor U12240 (N_12240,N_10549,N_10765);
or U12241 (N_12241,N_11271,N_11602);
and U12242 (N_12242,N_11349,N_10241);
xnor U12243 (N_12243,N_10497,N_10696);
or U12244 (N_12244,N_10339,N_11683);
or U12245 (N_12245,N_11731,N_10788);
nand U12246 (N_12246,N_10568,N_11175);
xor U12247 (N_12247,N_11606,N_11320);
nor U12248 (N_12248,N_10375,N_11711);
xor U12249 (N_12249,N_10565,N_11515);
nor U12250 (N_12250,N_11272,N_10094);
and U12251 (N_12251,N_11167,N_11417);
nand U12252 (N_12252,N_10117,N_10660);
xnor U12253 (N_12253,N_10802,N_10439);
or U12254 (N_12254,N_11379,N_11869);
xor U12255 (N_12255,N_10512,N_10323);
and U12256 (N_12256,N_10968,N_11002);
nor U12257 (N_12257,N_11042,N_11472);
nand U12258 (N_12258,N_10510,N_10720);
nor U12259 (N_12259,N_11497,N_10900);
xor U12260 (N_12260,N_10640,N_11211);
or U12261 (N_12261,N_11952,N_11956);
or U12262 (N_12262,N_10678,N_10706);
or U12263 (N_12263,N_11702,N_10149);
xor U12264 (N_12264,N_10299,N_10274);
and U12265 (N_12265,N_11127,N_11313);
and U12266 (N_12266,N_10422,N_11119);
or U12267 (N_12267,N_11712,N_11967);
or U12268 (N_12268,N_10822,N_10508);
or U12269 (N_12269,N_10263,N_11161);
or U12270 (N_12270,N_11555,N_11314);
nor U12271 (N_12271,N_11697,N_11163);
or U12272 (N_12272,N_11855,N_11837);
and U12273 (N_12273,N_11338,N_11392);
and U12274 (N_12274,N_11610,N_10846);
xnor U12275 (N_12275,N_11452,N_11380);
xor U12276 (N_12276,N_10536,N_11893);
xnor U12277 (N_12277,N_10158,N_11727);
or U12278 (N_12278,N_11036,N_10515);
nor U12279 (N_12279,N_11381,N_10516);
and U12280 (N_12280,N_10631,N_11106);
nor U12281 (N_12281,N_10578,N_10057);
or U12282 (N_12282,N_11518,N_10829);
nor U12283 (N_12283,N_11655,N_10534);
or U12284 (N_12284,N_10411,N_11246);
nor U12285 (N_12285,N_10449,N_10902);
nor U12286 (N_12286,N_10704,N_11577);
and U12287 (N_12287,N_11336,N_10210);
and U12288 (N_12288,N_11886,N_11240);
and U12289 (N_12289,N_10648,N_10909);
nor U12290 (N_12290,N_10795,N_11091);
nand U12291 (N_12291,N_11261,N_11451);
or U12292 (N_12292,N_11838,N_11693);
nor U12293 (N_12293,N_11342,N_11060);
xnor U12294 (N_12294,N_11031,N_10371);
and U12295 (N_12295,N_10106,N_10585);
nor U12296 (N_12296,N_10546,N_11444);
nor U12297 (N_12297,N_10374,N_11881);
nor U12298 (N_12298,N_10858,N_10304);
and U12299 (N_12299,N_10997,N_10473);
or U12300 (N_12300,N_11110,N_10386);
nand U12301 (N_12301,N_10781,N_11512);
nand U12302 (N_12302,N_10027,N_11402);
xor U12303 (N_12303,N_11816,N_10242);
and U12304 (N_12304,N_11014,N_10953);
nand U12305 (N_12305,N_10319,N_11165);
nand U12306 (N_12306,N_10014,N_11503);
nor U12307 (N_12307,N_11720,N_11351);
nor U12308 (N_12308,N_11648,N_10105);
and U12309 (N_12309,N_10310,N_10572);
nand U12310 (N_12310,N_10786,N_11612);
and U12311 (N_12311,N_10950,N_10824);
nor U12312 (N_12312,N_10770,N_10396);
or U12313 (N_12313,N_10552,N_11198);
and U12314 (N_12314,N_10352,N_10740);
and U12315 (N_12315,N_11598,N_11933);
nor U12316 (N_12316,N_11208,N_11782);
nor U12317 (N_12317,N_10172,N_10682);
xnor U12318 (N_12318,N_10959,N_11484);
or U12319 (N_12319,N_11684,N_11554);
xor U12320 (N_12320,N_11401,N_10198);
or U12321 (N_12321,N_11966,N_10555);
nor U12322 (N_12322,N_10366,N_10250);
xor U12323 (N_12323,N_11325,N_11688);
or U12324 (N_12324,N_11225,N_10838);
nor U12325 (N_12325,N_10826,N_11183);
nand U12326 (N_12326,N_11436,N_11725);
nor U12327 (N_12327,N_11109,N_10584);
and U12328 (N_12328,N_11652,N_10783);
or U12329 (N_12329,N_11501,N_10876);
or U12330 (N_12330,N_11756,N_11700);
xor U12331 (N_12331,N_10589,N_11385);
nor U12332 (N_12332,N_10700,N_11521);
xor U12333 (N_12333,N_11680,N_11221);
xor U12334 (N_12334,N_11207,N_11372);
xnor U12335 (N_12335,N_10251,N_10560);
nor U12336 (N_12336,N_11292,N_10963);
nand U12337 (N_12337,N_10104,N_10261);
nand U12338 (N_12338,N_10671,N_11113);
or U12339 (N_12339,N_10020,N_10810);
nor U12340 (N_12340,N_11061,N_11904);
and U12341 (N_12341,N_10523,N_10710);
xnor U12342 (N_12342,N_10697,N_11437);
nor U12343 (N_12343,N_10868,N_11734);
xnor U12344 (N_12344,N_10936,N_11291);
xnor U12345 (N_12345,N_10746,N_11996);
nor U12346 (N_12346,N_11214,N_10199);
or U12347 (N_12347,N_11039,N_10271);
and U12348 (N_12348,N_11138,N_11289);
nand U12349 (N_12349,N_11034,N_11722);
and U12350 (N_12350,N_10694,N_11442);
or U12351 (N_12351,N_10279,N_11957);
nor U12352 (N_12352,N_10085,N_10314);
or U12353 (N_12353,N_10074,N_10243);
or U12354 (N_12354,N_11199,N_10827);
nand U12355 (N_12355,N_11821,N_10597);
nor U12356 (N_12356,N_11508,N_11434);
nand U12357 (N_12357,N_10895,N_11457);
or U12358 (N_12358,N_10561,N_11854);
nor U12359 (N_12359,N_10961,N_11118);
or U12360 (N_12360,N_10095,N_10979);
xnor U12361 (N_12361,N_11811,N_10859);
xnor U12362 (N_12362,N_11414,N_11083);
and U12363 (N_12363,N_11757,N_10418);
or U12364 (N_12364,N_11133,N_10316);
nand U12365 (N_12365,N_10488,N_10747);
xor U12366 (N_12366,N_11140,N_10847);
xor U12367 (N_12367,N_10136,N_10254);
or U12368 (N_12368,N_11685,N_11248);
xnor U12369 (N_12369,N_10482,N_11148);
or U12370 (N_12370,N_10114,N_10993);
xor U12371 (N_12371,N_11262,N_10819);
or U12372 (N_12372,N_10815,N_10798);
and U12373 (N_12373,N_10026,N_10477);
and U12374 (N_12374,N_11387,N_11340);
nor U12375 (N_12375,N_11691,N_11235);
nor U12376 (N_12376,N_11024,N_10999);
nand U12377 (N_12377,N_10988,N_11396);
xor U12378 (N_12378,N_10155,N_11249);
nor U12379 (N_12379,N_10183,N_11840);
xor U12380 (N_12380,N_11860,N_11783);
or U12381 (N_12381,N_11883,N_10414);
nor U12382 (N_12382,N_11411,N_11216);
xor U12383 (N_12383,N_10529,N_10343);
and U12384 (N_12384,N_11990,N_10441);
and U12385 (N_12385,N_11275,N_10920);
nor U12386 (N_12386,N_11676,N_10991);
or U12387 (N_12387,N_10906,N_10690);
and U12388 (N_12388,N_11179,N_11259);
nor U12389 (N_12389,N_10220,N_10216);
xnor U12390 (N_12390,N_11339,N_11132);
nor U12391 (N_12391,N_10938,N_10791);
nor U12392 (N_12392,N_10357,N_11124);
or U12393 (N_12393,N_10312,N_10978);
nor U12394 (N_12394,N_11539,N_10047);
xor U12395 (N_12395,N_11128,N_10492);
xnor U12396 (N_12396,N_10884,N_10772);
nand U12397 (N_12397,N_10621,N_11825);
nor U12398 (N_12398,N_10330,N_11787);
xnor U12399 (N_12399,N_11446,N_11614);
nor U12400 (N_12400,N_10739,N_10634);
nand U12401 (N_12401,N_11245,N_11569);
or U12402 (N_12402,N_10990,N_10702);
xnor U12403 (N_12403,N_11178,N_10413);
and U12404 (N_12404,N_11800,N_10511);
xor U12405 (N_12405,N_11812,N_11256);
and U12406 (N_12406,N_10320,N_10799);
or U12407 (N_12407,N_10335,N_11678);
nand U12408 (N_12408,N_10364,N_11071);
and U12409 (N_12409,N_10519,N_11099);
nor U12410 (N_12410,N_10554,N_10882);
nand U12411 (N_12411,N_11778,N_11041);
or U12412 (N_12412,N_10429,N_10592);
and U12413 (N_12413,N_11200,N_11265);
xnor U12414 (N_12414,N_10234,N_11510);
or U12415 (N_12415,N_11559,N_10685);
nand U12416 (N_12416,N_11897,N_10601);
nor U12417 (N_12417,N_10259,N_11600);
xor U12418 (N_12418,N_10855,N_10409);
xnor U12419 (N_12419,N_10469,N_10351);
nand U12420 (N_12420,N_10405,N_10622);
xor U12421 (N_12421,N_11482,N_11891);
nor U12422 (N_12422,N_11771,N_11538);
nand U12423 (N_12423,N_10253,N_10354);
nor U12424 (N_12424,N_11912,N_11181);
or U12425 (N_12425,N_11516,N_11715);
xnor U12426 (N_12426,N_10823,N_10431);
nor U12427 (N_12427,N_10291,N_10611);
or U12428 (N_12428,N_10683,N_10599);
nand U12429 (N_12429,N_10539,N_10629);
or U12430 (N_12430,N_11595,N_11638);
or U12431 (N_12431,N_10503,N_10021);
or U12432 (N_12432,N_10147,N_11564);
and U12433 (N_12433,N_10338,N_10760);
or U12434 (N_12434,N_11913,N_10447);
and U12435 (N_12435,N_11474,N_10604);
nand U12436 (N_12436,N_11618,N_10836);
xor U12437 (N_12437,N_11629,N_10769);
or U12438 (N_12438,N_10023,N_11807);
and U12439 (N_12439,N_11493,N_10077);
xnor U12440 (N_12440,N_11122,N_10168);
xnor U12441 (N_12441,N_11662,N_11212);
nor U12442 (N_12442,N_10295,N_10879);
nand U12443 (N_12443,N_10005,N_11504);
xor U12444 (N_12444,N_11871,N_11866);
nor U12445 (N_12445,N_10735,N_10016);
nor U12446 (N_12446,N_11964,N_11485);
or U12447 (N_12447,N_10930,N_11000);
or U12448 (N_12448,N_10705,N_11829);
or U12449 (N_12449,N_11432,N_11058);
nand U12450 (N_12450,N_11176,N_11551);
nor U12451 (N_12451,N_10777,N_11266);
nand U12452 (N_12452,N_11984,N_10875);
nand U12453 (N_12453,N_10924,N_11868);
nor U12454 (N_12454,N_10500,N_10154);
xnor U12455 (N_12455,N_10230,N_11799);
nand U12456 (N_12456,N_11765,N_10787);
nor U12457 (N_12457,N_11834,N_11204);
xnor U12458 (N_12458,N_11019,N_11045);
xor U12459 (N_12459,N_10040,N_10353);
nor U12460 (N_12460,N_10532,N_10756);
and U12461 (N_12461,N_11137,N_10952);
nand U12462 (N_12462,N_10203,N_11611);
nand U12463 (N_12463,N_10430,N_11621);
and U12464 (N_12464,N_10423,N_11879);
and U12465 (N_12465,N_10845,N_10185);
xnor U12466 (N_12466,N_11910,N_11022);
and U12467 (N_12467,N_11400,N_10862);
or U12468 (N_12468,N_10916,N_11907);
nand U12469 (N_12469,N_10543,N_10219);
nand U12470 (N_12470,N_11750,N_11420);
xnor U12471 (N_12471,N_11149,N_10793);
or U12472 (N_12472,N_10571,N_11278);
and U12473 (N_12473,N_10495,N_10004);
nand U12474 (N_12474,N_11035,N_11874);
nor U12475 (N_12475,N_11220,N_10643);
nand U12476 (N_12476,N_10137,N_11057);
and U12477 (N_12477,N_11846,N_11524);
xnor U12478 (N_12478,N_10390,N_11882);
xnor U12479 (N_12479,N_10287,N_11117);
nand U12480 (N_12480,N_11591,N_11543);
nand U12481 (N_12481,N_10667,N_11714);
and U12482 (N_12482,N_11950,N_11995);
xor U12483 (N_12483,N_11930,N_11823);
nand U12484 (N_12484,N_10541,N_11656);
nand U12485 (N_12485,N_10966,N_10403);
nand U12486 (N_12486,N_11746,N_11029);
nor U12487 (N_12487,N_10670,N_11985);
and U12488 (N_12488,N_10303,N_11361);
and U12489 (N_12489,N_10334,N_10808);
and U12490 (N_12490,N_11435,N_10135);
nor U12491 (N_12491,N_11726,N_10645);
nand U12492 (N_12492,N_10664,N_10417);
nand U12493 (N_12493,N_10871,N_10100);
xor U12494 (N_12494,N_10736,N_10937);
and U12495 (N_12495,N_11670,N_11013);
xnor U12496 (N_12496,N_11718,N_10433);
xor U12497 (N_12497,N_10917,N_10928);
nand U12498 (N_12498,N_11951,N_10981);
or U12499 (N_12499,N_10190,N_10273);
or U12500 (N_12500,N_11896,N_11658);
nor U12501 (N_12501,N_11419,N_11644);
xnor U12502 (N_12502,N_10524,N_10642);
xnor U12503 (N_12503,N_11431,N_11228);
nand U12504 (N_12504,N_10197,N_11130);
xnor U12505 (N_12505,N_10089,N_10998);
nor U12506 (N_12506,N_11553,N_10309);
and U12507 (N_12507,N_10526,N_10486);
or U12508 (N_12508,N_11344,N_10248);
nor U12509 (N_12509,N_11363,N_11226);
nand U12510 (N_12510,N_10202,N_11288);
xnor U12511 (N_12511,N_11236,N_11357);
or U12512 (N_12512,N_10121,N_10244);
and U12513 (N_12513,N_10406,N_10588);
or U12514 (N_12514,N_11477,N_11833);
or U12515 (N_12515,N_10551,N_10432);
or U12516 (N_12516,N_11051,N_10453);
or U12517 (N_12517,N_10547,N_11064);
nand U12518 (N_12518,N_11465,N_10960);
nand U12519 (N_12519,N_11853,N_11753);
or U12520 (N_12520,N_11706,N_11998);
or U12521 (N_12521,N_10828,N_11895);
nand U12522 (N_12522,N_11250,N_11287);
nand U12523 (N_12523,N_10581,N_10080);
nor U12524 (N_12524,N_11637,N_11983);
or U12525 (N_12525,N_11677,N_11151);
xor U12526 (N_12526,N_10160,N_10109);
or U12527 (N_12527,N_10139,N_10901);
nand U12528 (N_12528,N_11747,N_11095);
or U12529 (N_12529,N_11738,N_10954);
xnor U12530 (N_12530,N_10156,N_10707);
nor U12531 (N_12531,N_10071,N_11244);
xor U12532 (N_12532,N_10465,N_11947);
nand U12533 (N_12533,N_11488,N_10459);
xnor U12534 (N_12534,N_11428,N_11931);
xor U12535 (N_12535,N_10031,N_10011);
nand U12536 (N_12536,N_11570,N_10052);
nor U12537 (N_12537,N_11050,N_11247);
xor U12538 (N_12538,N_11312,N_10970);
nor U12539 (N_12539,N_11824,N_10595);
and U12540 (N_12540,N_10206,N_10743);
or U12541 (N_12541,N_10722,N_11604);
xnor U12542 (N_12542,N_11914,N_11136);
nand U12543 (N_12543,N_10528,N_10471);
nor U12544 (N_12544,N_10995,N_10771);
or U12545 (N_12545,N_10801,N_11427);
or U12546 (N_12546,N_11197,N_10009);
nand U12547 (N_12547,N_10045,N_11364);
nand U12548 (N_12548,N_11798,N_11517);
nand U12549 (N_12549,N_10837,N_11088);
nor U12550 (N_12550,N_10703,N_11056);
nand U12551 (N_12551,N_10108,N_10053);
and U12552 (N_12552,N_10264,N_11341);
nor U12553 (N_12553,N_10800,N_11260);
xor U12554 (N_12554,N_11494,N_11375);
and U12555 (N_12555,N_10780,N_10003);
or U12556 (N_12556,N_11953,N_10288);
or U12557 (N_12557,N_11536,N_10899);
or U12558 (N_12558,N_10945,N_10035);
xor U12559 (N_12559,N_11580,N_10932);
and U12560 (N_12560,N_10624,N_11112);
nor U12561 (N_12561,N_10655,N_11777);
or U12562 (N_12562,N_11852,N_11997);
or U12563 (N_12563,N_10984,N_11576);
or U12564 (N_12564,N_11970,N_11918);
and U12565 (N_12565,N_11528,N_11972);
nand U12566 (N_12566,N_10468,N_11254);
nand U12567 (N_12567,N_11663,N_10817);
nor U12568 (N_12568,N_10217,N_11968);
xnor U12569 (N_12569,N_11487,N_10464);
nand U12570 (N_12570,N_11760,N_11172);
nand U12571 (N_12571,N_10763,N_10268);
xnor U12572 (N_12572,N_10270,N_10373);
or U12573 (N_12573,N_10445,N_10325);
xnor U12574 (N_12574,N_11965,N_11766);
xnor U12575 (N_12575,N_11462,N_10326);
nor U12576 (N_12576,N_10348,N_11237);
or U12577 (N_12577,N_10504,N_11548);
xor U12578 (N_12578,N_11188,N_10002);
nand U12579 (N_12579,N_11949,N_10891);
or U12580 (N_12580,N_10907,N_10341);
nor U12581 (N_12581,N_10792,N_10118);
nand U12582 (N_12582,N_11368,N_11020);
xnor U12583 (N_12583,N_11857,N_11946);
or U12584 (N_12584,N_10041,N_10753);
nand U12585 (N_12585,N_11903,N_10450);
or U12586 (N_12586,N_10296,N_11547);
and U12587 (N_12587,N_10455,N_10531);
and U12588 (N_12588,N_11066,N_11646);
nor U12589 (N_12589,N_11297,N_11044);
nor U12590 (N_12590,N_10785,N_10305);
or U12591 (N_12591,N_11628,N_11526);
or U12592 (N_12592,N_10213,N_11541);
xor U12593 (N_12593,N_10088,N_10321);
and U12594 (N_12594,N_11922,N_10852);
xnor U12595 (N_12595,N_11450,N_11719);
nor U12596 (N_12596,N_10521,N_11386);
nor U12597 (N_12597,N_11098,N_10221);
xor U12598 (N_12598,N_11072,N_11463);
nand U12599 (N_12599,N_11027,N_11779);
xnor U12600 (N_12600,N_11310,N_11103);
nand U12601 (N_12601,N_10731,N_11962);
or U12602 (N_12602,N_10223,N_11762);
and U12603 (N_12603,N_11369,N_10603);
nor U12604 (N_12604,N_10487,N_10039);
xnor U12605 (N_12605,N_10608,N_10894);
nand U12606 (N_12606,N_10773,N_10394);
nand U12607 (N_12607,N_11772,N_10517);
nor U12608 (N_12608,N_10507,N_10728);
or U12609 (N_12609,N_10583,N_11481);
and U12610 (N_12610,N_10723,N_11466);
xor U12611 (N_12611,N_10300,N_11067);
nor U12612 (N_12612,N_11243,N_11924);
xnor U12613 (N_12613,N_10475,N_11146);
or U12614 (N_12614,N_10641,N_11471);
nor U12615 (N_12615,N_10814,N_10102);
nand U12616 (N_12616,N_10778,N_11872);
and U12617 (N_12617,N_10491,N_11453);
nor U12618 (N_12618,N_10805,N_10666);
nor U12619 (N_12619,N_11944,N_11633);
and U12620 (N_12620,N_11742,N_11005);
xnor U12621 (N_12621,N_10290,N_11366);
nand U12622 (N_12622,N_11069,N_11575);
xnor U12623 (N_12623,N_11264,N_10036);
or U12624 (N_12624,N_10562,N_10425);
xor U12625 (N_12625,N_11023,N_11705);
xnor U12626 (N_12626,N_10582,N_10967);
xnor U12627 (N_12627,N_11622,N_11669);
xnor U12628 (N_12628,N_11651,N_11755);
nand U12629 (N_12629,N_11100,N_11303);
and U12630 (N_12630,N_11730,N_10388);
nor U12631 (N_12631,N_10880,N_10980);
nand U12632 (N_12632,N_11445,N_11708);
or U12633 (N_12633,N_10395,N_10317);
and U12634 (N_12634,N_11804,N_10618);
xor U12635 (N_12635,N_10840,N_11276);
or U12636 (N_12636,N_10257,N_10481);
or U12637 (N_12637,N_11343,N_11101);
nand U12638 (N_12638,N_10931,N_11404);
nand U12639 (N_12639,N_11793,N_11406);
or U12640 (N_12640,N_11169,N_11977);
and U12641 (N_12641,N_11701,N_11296);
and U12642 (N_12642,N_10910,N_11021);
or U12643 (N_12643,N_11160,N_11571);
nand U12644 (N_12644,N_10286,N_10457);
nand U12645 (N_12645,N_11791,N_10730);
nand U12646 (N_12646,N_11495,N_11822);
or U12647 (N_12647,N_10973,N_10958);
and U12648 (N_12648,N_11759,N_11439);
or U12649 (N_12649,N_11850,N_11919);
and U12650 (N_12650,N_10918,N_10157);
nand U12651 (N_12651,N_11625,N_10133);
nand U12652 (N_12652,N_10346,N_10421);
and U12653 (N_12653,N_11925,N_11535);
xnor U12654 (N_12654,N_11813,N_10755);
nor U12655 (N_12655,N_10751,N_10446);
nand U12656 (N_12656,N_11478,N_11121);
and U12657 (N_12657,N_10380,N_10324);
xnor U12658 (N_12658,N_10060,N_10806);
and U12659 (N_12659,N_10985,N_11650);
xnor U12660 (N_12660,N_10496,N_11926);
and U12661 (N_12661,N_11616,N_11311);
and U12662 (N_12662,N_10151,N_10887);
or U12663 (N_12663,N_10237,N_11317);
or U12664 (N_12664,N_11145,N_10926);
or U12665 (N_12665,N_10518,N_10377);
xnor U12666 (N_12666,N_10686,N_10498);
nor U12667 (N_12667,N_10885,N_11994);
nand U12668 (N_12668,N_11959,N_10689);
and U12669 (N_12669,N_10327,N_10898);
or U12670 (N_12670,N_10553,N_11819);
and U12671 (N_12671,N_11885,N_11695);
nor U12672 (N_12672,N_11732,N_11141);
and U12673 (N_12673,N_11295,N_11627);
xor U12674 (N_12674,N_11376,N_11620);
or U12675 (N_12675,N_10350,N_10839);
nor U12676 (N_12676,N_11590,N_11196);
nor U12677 (N_12677,N_10442,N_10024);
nor U12678 (N_12678,N_11073,N_10525);
xor U12679 (N_12679,N_11560,N_10152);
nand U12680 (N_12680,N_10078,N_10628);
or U12681 (N_12681,N_11152,N_11597);
and U12682 (N_12682,N_10252,N_10056);
nor U12683 (N_12683,N_10947,N_11430);
and U12684 (N_12684,N_10870,N_11563);
xnor U12685 (N_12685,N_10877,N_10120);
xnor U12686 (N_12686,N_10615,N_11158);
xor U12687 (N_12687,N_10272,N_11086);
xnor U12688 (N_12688,N_10122,N_10191);
xnor U12689 (N_12689,N_10598,N_10193);
nor U12690 (N_12690,N_11142,N_11507);
nand U12691 (N_12691,N_11371,N_11649);
nand U12692 (N_12692,N_11948,N_11640);
xnor U12693 (N_12693,N_10676,N_11729);
nand U12694 (N_12694,N_10478,N_10079);
and U12695 (N_12695,N_10044,N_11194);
and U12696 (N_12696,N_11686,N_11898);
and U12697 (N_12697,N_11976,N_10101);
nor U12698 (N_12698,N_10556,N_10962);
nand U12699 (N_12699,N_11241,N_11412);
xor U12700 (N_12700,N_11583,N_10018);
or U12701 (N_12701,N_11631,N_11502);
nand U12702 (N_12702,N_10946,N_10904);
and U12703 (N_12703,N_11744,N_10434);
xor U12704 (N_12704,N_11407,N_11394);
nor U12705 (N_12705,N_11724,N_11615);
xor U12706 (N_12706,N_11084,N_10509);
xnor U12707 (N_12707,N_10825,N_11870);
xor U12708 (N_12708,N_11438,N_10861);
nor U12709 (N_12709,N_11703,N_11572);
nand U12710 (N_12710,N_11251,N_10835);
nor U12711 (N_12711,N_11592,N_11982);
and U12712 (N_12712,N_10540,N_11307);
nand U12713 (N_12713,N_10742,N_11562);
nand U12714 (N_12714,N_10398,N_11810);
and U12715 (N_12715,N_10662,N_11074);
and U12716 (N_12716,N_10754,N_11332);
nor U12717 (N_12717,N_11177,N_11911);
nor U12718 (N_12718,N_11704,N_11009);
and U12719 (N_12719,N_11748,N_11301);
nor U12720 (N_12720,N_11263,N_11189);
xor U12721 (N_12721,N_11293,N_10964);
nand U12722 (N_12722,N_11097,N_10090);
or U12723 (N_12723,N_10874,N_10734);
and U12724 (N_12724,N_10038,N_10708);
xnor U12725 (N_12725,N_10384,N_10976);
nor U12726 (N_12726,N_10382,N_11667);
xnor U12727 (N_12727,N_11425,N_11054);
and U12728 (N_12728,N_10144,N_10564);
xnor U12729 (N_12729,N_11053,N_11877);
or U12730 (N_12730,N_10236,N_11017);
nand U12731 (N_12731,N_11674,N_10574);
or U12732 (N_12732,N_10289,N_11739);
or U12733 (N_12733,N_10668,N_11578);
and U12734 (N_12734,N_11267,N_11639);
xnor U12735 (N_12735,N_10207,N_10850);
or U12736 (N_12736,N_11792,N_10356);
and U12737 (N_12737,N_11234,N_10328);
nor U12738 (N_12738,N_10724,N_11603);
or U12739 (N_12739,N_11856,N_10050);
and U12740 (N_12740,N_10461,N_11421);
xor U12741 (N_12741,N_11936,N_10545);
xor U12742 (N_12742,N_10255,N_10393);
nand U12743 (N_12743,N_10391,N_11123);
xnor U12744 (N_12744,N_10049,N_11542);
nand U12745 (N_12745,N_10181,N_10721);
or U12746 (N_12746,N_11586,N_10951);
or U12747 (N_12747,N_10501,N_11318);
nor U12748 (N_12748,N_10239,N_11015);
nor U12749 (N_12749,N_11134,N_11155);
or U12750 (N_12750,N_10758,N_11075);
nor U12751 (N_12751,N_11588,N_11468);
nand U12752 (N_12752,N_11305,N_10831);
and U12753 (N_12753,N_10867,N_10942);
nor U12754 (N_12754,N_11863,N_10663);
nand U12755 (N_12755,N_11980,N_10633);
and U12756 (N_12756,N_11989,N_11749);
nand U12757 (N_12757,N_10972,N_10566);
nand U12758 (N_12758,N_10329,N_10713);
nand U12759 (N_12759,N_11168,N_10013);
nor U12760 (N_12760,N_10012,N_10344);
nor U12761 (N_12761,N_11803,N_10649);
and U12762 (N_12762,N_10653,N_10083);
or U12763 (N_12763,N_11801,N_10476);
or U12764 (N_12764,N_11505,N_11257);
nor U12765 (N_12765,N_11523,N_11689);
or U12766 (N_12766,N_10059,N_10076);
nand U12767 (N_12767,N_11809,N_10709);
nor U12768 (N_12768,N_10378,N_11229);
or U12769 (N_12769,N_11038,N_11328);
xor U12770 (N_12770,N_11218,N_11902);
and U12771 (N_12771,N_10000,N_11277);
or U12772 (N_12772,N_11082,N_11797);
nand U12773 (N_12773,N_11770,N_10620);
nand U12774 (N_12774,N_10062,N_11632);
or U12775 (N_12775,N_11316,N_10558);
nor U12776 (N_12776,N_11887,N_11040);
and U12777 (N_12777,N_11279,N_10460);
nand U12778 (N_12778,N_10651,N_10652);
and U12779 (N_12779,N_10030,N_10948);
nand U12780 (N_12780,N_10070,N_10204);
xnor U12781 (N_12781,N_10258,N_11397);
or U12782 (N_12782,N_11173,N_11239);
nand U12783 (N_12783,N_10428,N_10881);
or U12784 (N_12784,N_11373,N_10856);
nor U12785 (N_12785,N_11617,N_11230);
nand U12786 (N_12786,N_11353,N_11096);
xor U12787 (N_12787,N_10883,N_11634);
xor U12788 (N_12788,N_10613,N_10143);
or U12789 (N_12789,N_10400,N_10440);
nand U12790 (N_12790,N_10175,N_10399);
nand U12791 (N_12791,N_11710,N_10617);
xor U12792 (N_12792,N_10794,N_10436);
or U12793 (N_12793,N_11326,N_10848);
nand U12794 (N_12794,N_11582,N_11992);
xnor U12795 (N_12795,N_11532,N_11681);
nor U12796 (N_12796,N_11489,N_10878);
nand U12797 (N_12797,N_10437,N_11942);
nor U12798 (N_12798,N_10178,N_10632);
and U12799 (N_12799,N_10919,N_10484);
xnor U12800 (N_12800,N_11673,N_10201);
or U12801 (N_12801,N_11561,N_11460);
nand U12802 (N_12802,N_11356,N_10113);
or U12803 (N_12803,N_11129,N_10412);
nor U12804 (N_12804,N_11943,N_11773);
xor U12805 (N_12805,N_10606,N_10116);
xnor U12806 (N_12806,N_11839,N_11185);
and U12807 (N_12807,N_10580,N_11954);
nor U12808 (N_12808,N_11899,N_10311);
nor U12809 (N_12809,N_11426,N_10125);
nand U12810 (N_12810,N_11758,N_10342);
nand U12811 (N_12811,N_10596,N_11694);
nand U12812 (N_12812,N_11986,N_10087);
nor U12813 (N_12813,N_10126,N_10073);
or U12814 (N_12814,N_11867,N_10131);
or U12815 (N_12815,N_11987,N_11223);
and U12816 (N_12816,N_10184,N_11934);
xnor U12817 (N_12817,N_11423,N_10298);
or U12818 (N_12818,N_11550,N_10654);
nor U12819 (N_12819,N_11790,N_10527);
and U12820 (N_12820,N_11932,N_11011);
nand U12821 (N_12821,N_11078,N_11354);
and U12822 (N_12822,N_11008,N_11696);
nor U12823 (N_12823,N_11268,N_10332);
nand U12824 (N_12824,N_11143,N_10674);
nand U12825 (N_12825,N_10927,N_10759);
nor U12826 (N_12826,N_10112,N_11004);
or U12827 (N_12827,N_11849,N_11567);
xnor U12828 (N_12828,N_10365,N_10712);
or U12829 (N_12829,N_10779,N_10058);
xor U12830 (N_12830,N_11156,N_10032);
and U12831 (N_12831,N_10466,N_11608);
nor U12832 (N_12832,N_11242,N_10996);
or U12833 (N_12833,N_11991,N_10865);
xnor U12834 (N_12834,N_10282,N_10656);
nand U12835 (N_12835,N_11367,N_10716);
and U12836 (N_12836,N_10345,N_10863);
nand U12837 (N_12837,N_10153,N_10567);
or U12838 (N_12838,N_11294,N_10408);
xnor U12839 (N_12839,N_11520,N_10293);
nand U12840 (N_12840,N_10557,N_11858);
or U12841 (N_12841,N_10194,N_11776);
and U12842 (N_12842,N_11499,N_11395);
xnor U12843 (N_12843,N_10903,N_11087);
xor U12844 (N_12844,N_10008,N_10955);
and U12845 (N_12845,N_10034,N_11641);
nand U12846 (N_12846,N_10854,N_10281);
xnor U12847 (N_12847,N_10046,N_10180);
and U12848 (N_12848,N_11139,N_11076);
nand U12849 (N_12849,N_11537,N_11814);
nor U12850 (N_12850,N_10130,N_11456);
or U12851 (N_12851,N_11587,N_10103);
xnor U12852 (N_12852,N_11596,N_10563);
xnor U12853 (N_12853,N_11789,N_11391);
and U12854 (N_12854,N_10029,N_10132);
or U12855 (N_12855,N_11831,N_11440);
nor U12856 (N_12856,N_10075,N_11549);
or U12857 (N_12857,N_10187,N_11335);
xnor U12858 (N_12858,N_11664,N_11273);
xor U12859 (N_12859,N_10669,N_11999);
and U12860 (N_12860,N_10741,N_11815);
nor U12861 (N_12861,N_11923,N_11958);
and U12862 (N_12862,N_11579,N_10693);
or U12863 (N_12863,N_10146,N_11410);
xnor U12864 (N_12864,N_10593,N_11224);
nand U12865 (N_12865,N_10714,N_11253);
and U12866 (N_12866,N_11665,N_10322);
nor U12867 (N_12867,N_10857,N_11707);
and U12868 (N_12868,N_11322,N_11506);
nand U12869 (N_12869,N_10737,N_10415);
nor U12870 (N_12870,N_10490,N_10372);
or U12871 (N_12871,N_10934,N_11767);
xnor U12872 (N_12872,N_11213,N_11540);
xor U12873 (N_12873,N_10205,N_11979);
nor U12874 (N_12874,N_11917,N_10275);
nand U12875 (N_12875,N_10173,N_11010);
nor U12876 (N_12876,N_11388,N_10392);
and U12877 (N_12877,N_11195,N_11636);
xnor U12878 (N_12878,N_11514,N_10803);
or U12879 (N_12879,N_11166,N_11915);
xor U12880 (N_12880,N_11845,N_10762);
or U12881 (N_12881,N_11530,N_10037);
xor U12882 (N_12882,N_10462,N_10502);
or U12883 (N_12883,N_11479,N_10015);
or U12884 (N_12884,N_10480,N_10933);
and U12885 (N_12885,N_10569,N_11842);
nor U12886 (N_12886,N_10162,N_11209);
nand U12887 (N_12887,N_10804,N_11003);
xor U12888 (N_12888,N_10306,N_11458);
nand U12889 (N_12889,N_10082,N_11557);
or U12890 (N_12890,N_10625,N_10677);
xnor U12891 (N_12891,N_10218,N_11889);
or U12892 (N_12892,N_10922,N_10276);
and U12893 (N_12893,N_10489,N_11491);
and U12894 (N_12894,N_11202,N_10969);
xnor U12895 (N_12895,N_10559,N_11486);
and U12896 (N_12896,N_11589,N_11037);
or U12897 (N_12897,N_11321,N_11068);
nor U12898 (N_12898,N_10055,N_11384);
and U12899 (N_12899,N_10084,N_10368);
nor U12900 (N_12900,N_10401,N_10424);
or U12901 (N_12901,N_10448,N_10789);
xnor U12902 (N_12902,N_10602,N_11544);
xnor U12903 (N_12903,N_10416,N_11880);
xor U12904 (N_12904,N_11661,N_10483);
nand U12905 (N_12905,N_11642,N_11131);
nand U12906 (N_12906,N_11144,N_10127);
xor U12907 (N_12907,N_11283,N_10067);
xor U12908 (N_12908,N_10091,N_10232);
nor U12909 (N_12909,N_10337,N_10240);
nand U12910 (N_12910,N_10646,N_10150);
and U12911 (N_12911,N_10614,N_11928);
and U12912 (N_12912,N_11016,N_11347);
or U12913 (N_12913,N_11298,N_10247);
and U12914 (N_12914,N_11735,N_11399);
or U12915 (N_12915,N_11630,N_11961);
and U12916 (N_12916,N_10893,N_10072);
xor U12917 (N_12917,N_10387,N_10860);
nand U12918 (N_12918,N_10262,N_10911);
nand U12919 (N_12919,N_10086,N_10701);
or U12920 (N_12920,N_10619,N_11941);
or U12921 (N_12921,N_11345,N_10832);
nand U12922 (N_12922,N_11012,N_10010);
and U12923 (N_12923,N_10635,N_10834);
xor U12924 (N_12924,N_10579,N_11157);
nor U12925 (N_12925,N_11455,N_11280);
or U12926 (N_12926,N_11826,N_11659);
xnor U12927 (N_12927,N_11483,N_11921);
xor U12928 (N_12928,N_11033,N_11309);
and U12929 (N_12929,N_10302,N_11186);
nor U12930 (N_12930,N_10986,N_11174);
nand U12931 (N_12931,N_10729,N_11566);
nor U12932 (N_12932,N_11070,N_11299);
or U12933 (N_12933,N_10844,N_10889);
or U12934 (N_12934,N_11359,N_10506);
nand U12935 (N_12935,N_11802,N_10443);
nand U12936 (N_12936,N_10914,N_10235);
xor U12937 (N_12937,N_11459,N_11147);
and U12938 (N_12938,N_10535,N_10647);
xor U12939 (N_12939,N_10542,N_10096);
and U12940 (N_12940,N_11672,N_10956);
nor U12941 (N_12941,N_11255,N_11888);
or U12942 (N_12942,N_11892,N_11884);
xnor U12943 (N_12943,N_10224,N_11448);
and U12944 (N_12944,N_10426,N_10389);
xor U12945 (N_12945,N_11900,N_11533);
xor U12946 (N_12946,N_11527,N_10444);
and U12947 (N_12947,N_10732,N_10006);
xor U12948 (N_12948,N_11733,N_11352);
xnor U12949 (N_12949,N_10612,N_10738);
xnor U12950 (N_12950,N_11927,N_11552);
xor U12951 (N_12951,N_11164,N_10134);
or U12952 (N_12952,N_10140,N_11433);
and U12953 (N_12953,N_10821,N_11920);
or U12954 (N_12954,N_11836,N_11859);
nand U12955 (N_12955,N_10513,N_10284);
and U12956 (N_12956,N_10811,N_11973);
nand U12957 (N_12957,N_10142,N_11079);
nor U12958 (N_12958,N_10630,N_11018);
xor U12959 (N_12959,N_10989,N_11274);
nand U12960 (N_12960,N_11370,N_10438);
or U12961 (N_12961,N_10725,N_10463);
and U12962 (N_12962,N_11469,N_11480);
nand U12963 (N_12963,N_10957,N_11786);
xnor U12964 (N_12964,N_10851,N_11861);
nand U12965 (N_12965,N_10897,N_10169);
nand U12966 (N_12966,N_11498,N_11546);
and U12967 (N_12967,N_10294,N_10167);
or U12968 (N_12968,N_11284,N_10849);
nor U12969 (N_12969,N_11192,N_11089);
nand U12970 (N_12970,N_11390,N_10313);
nand U12971 (N_12971,N_11827,N_11593);
nor U12972 (N_12972,N_11429,N_10784);
nor U12973 (N_12973,N_10698,N_11763);
nand U12974 (N_12974,N_11454,N_10866);
or U12975 (N_12975,N_11006,N_11509);
nand U12976 (N_12976,N_10650,N_11728);
nand U12977 (N_12977,N_11534,N_11114);
nand U12978 (N_12978,N_10609,N_10404);
xor U12979 (N_12979,N_10171,N_10308);
and U12980 (N_12980,N_10427,N_11781);
and U12981 (N_12981,N_11191,N_11745);
nand U12982 (N_12982,N_10533,N_11269);
xnor U12983 (N_12983,N_11282,N_10570);
nor U12984 (N_12984,N_10182,N_11768);
xnor U12985 (N_12985,N_10110,N_11862);
nand U12986 (N_12986,N_10661,N_10238);
and U12987 (N_12987,N_10174,N_11723);
or U12988 (N_12988,N_11047,N_10680);
nand U12989 (N_12989,N_11743,N_11331);
and U12990 (N_12990,N_10841,N_11422);
nand U12991 (N_12991,N_11415,N_11906);
nor U12992 (N_12992,N_11736,N_10245);
xnor U12993 (N_12993,N_11687,N_10148);
nor U12994 (N_12994,N_10761,N_11120);
nor U12995 (N_12995,N_10616,N_11374);
or U12996 (N_12996,N_11643,N_11170);
and U12997 (N_12997,N_10812,N_11558);
nand U12998 (N_12998,N_11304,N_11362);
and U12999 (N_12999,N_10949,N_11323);
nand U13000 (N_13000,N_10316,N_11998);
nor U13001 (N_13001,N_11734,N_11241);
and U13002 (N_13002,N_10807,N_10459);
or U13003 (N_13003,N_11475,N_11103);
nor U13004 (N_13004,N_10104,N_11844);
nor U13005 (N_13005,N_11539,N_11841);
nand U13006 (N_13006,N_10695,N_10766);
and U13007 (N_13007,N_11943,N_10741);
nor U13008 (N_13008,N_10056,N_10610);
nor U13009 (N_13009,N_11839,N_10725);
xnor U13010 (N_13010,N_11631,N_11948);
nand U13011 (N_13011,N_10303,N_11369);
nor U13012 (N_13012,N_11705,N_11601);
or U13013 (N_13013,N_11616,N_10323);
or U13014 (N_13014,N_10643,N_11928);
nor U13015 (N_13015,N_11440,N_10503);
and U13016 (N_13016,N_11256,N_10619);
nand U13017 (N_13017,N_10117,N_11647);
nand U13018 (N_13018,N_10611,N_10659);
xnor U13019 (N_13019,N_11656,N_11954);
and U13020 (N_13020,N_11552,N_11889);
nor U13021 (N_13021,N_10101,N_10967);
or U13022 (N_13022,N_10281,N_11055);
or U13023 (N_13023,N_10850,N_10315);
and U13024 (N_13024,N_11590,N_10258);
nand U13025 (N_13025,N_11332,N_11281);
xor U13026 (N_13026,N_11597,N_10951);
or U13027 (N_13027,N_10751,N_11621);
nor U13028 (N_13028,N_10045,N_10052);
and U13029 (N_13029,N_10892,N_10352);
xnor U13030 (N_13030,N_10297,N_10380);
nand U13031 (N_13031,N_11517,N_10618);
nand U13032 (N_13032,N_10035,N_10188);
nand U13033 (N_13033,N_11786,N_10353);
xnor U13034 (N_13034,N_11881,N_11528);
nor U13035 (N_13035,N_10354,N_10900);
nand U13036 (N_13036,N_10076,N_11154);
or U13037 (N_13037,N_10211,N_10952);
or U13038 (N_13038,N_10745,N_11441);
xnor U13039 (N_13039,N_11549,N_10910);
nor U13040 (N_13040,N_10824,N_10210);
xor U13041 (N_13041,N_10658,N_10224);
or U13042 (N_13042,N_10585,N_10059);
xor U13043 (N_13043,N_10956,N_11071);
or U13044 (N_13044,N_10137,N_11155);
xor U13045 (N_13045,N_10807,N_11163);
or U13046 (N_13046,N_11779,N_11392);
nor U13047 (N_13047,N_11883,N_11102);
nor U13048 (N_13048,N_10496,N_11403);
or U13049 (N_13049,N_11945,N_10031);
nand U13050 (N_13050,N_10664,N_11060);
nand U13051 (N_13051,N_10597,N_10862);
nor U13052 (N_13052,N_11417,N_11883);
and U13053 (N_13053,N_10551,N_10242);
or U13054 (N_13054,N_11128,N_10170);
xor U13055 (N_13055,N_11023,N_10674);
nand U13056 (N_13056,N_11990,N_10092);
nand U13057 (N_13057,N_11193,N_10216);
and U13058 (N_13058,N_10552,N_10526);
and U13059 (N_13059,N_10798,N_10391);
xnor U13060 (N_13060,N_10865,N_10671);
nand U13061 (N_13061,N_11410,N_10335);
and U13062 (N_13062,N_11919,N_10730);
xor U13063 (N_13063,N_11036,N_10692);
or U13064 (N_13064,N_11008,N_10729);
nand U13065 (N_13065,N_10301,N_10458);
nor U13066 (N_13066,N_11940,N_10044);
nor U13067 (N_13067,N_11968,N_10977);
or U13068 (N_13068,N_10090,N_11942);
or U13069 (N_13069,N_11366,N_10425);
nand U13070 (N_13070,N_10962,N_10135);
nor U13071 (N_13071,N_11023,N_10128);
or U13072 (N_13072,N_10493,N_11578);
and U13073 (N_13073,N_10906,N_10274);
or U13074 (N_13074,N_10358,N_10215);
xor U13075 (N_13075,N_11037,N_10854);
nor U13076 (N_13076,N_11909,N_10687);
nand U13077 (N_13077,N_11294,N_11066);
nor U13078 (N_13078,N_11054,N_11141);
nand U13079 (N_13079,N_10932,N_11489);
or U13080 (N_13080,N_10847,N_10458);
or U13081 (N_13081,N_11814,N_10930);
nand U13082 (N_13082,N_10196,N_10895);
or U13083 (N_13083,N_10310,N_10752);
nand U13084 (N_13084,N_10243,N_10090);
nand U13085 (N_13085,N_11439,N_11311);
xor U13086 (N_13086,N_11122,N_11259);
or U13087 (N_13087,N_11112,N_11888);
xor U13088 (N_13088,N_10048,N_11355);
xor U13089 (N_13089,N_11271,N_10061);
or U13090 (N_13090,N_10188,N_10013);
xnor U13091 (N_13091,N_11407,N_11870);
or U13092 (N_13092,N_10700,N_11715);
nand U13093 (N_13093,N_10262,N_11577);
or U13094 (N_13094,N_11600,N_11581);
or U13095 (N_13095,N_10447,N_11443);
or U13096 (N_13096,N_11246,N_11112);
or U13097 (N_13097,N_10328,N_10553);
xnor U13098 (N_13098,N_11686,N_11467);
xnor U13099 (N_13099,N_10202,N_11972);
nand U13100 (N_13100,N_10399,N_10875);
or U13101 (N_13101,N_10368,N_10394);
and U13102 (N_13102,N_11407,N_11157);
or U13103 (N_13103,N_10016,N_10597);
or U13104 (N_13104,N_10135,N_10817);
xnor U13105 (N_13105,N_10828,N_10434);
or U13106 (N_13106,N_11399,N_11189);
xor U13107 (N_13107,N_11582,N_11848);
xor U13108 (N_13108,N_10184,N_11693);
nor U13109 (N_13109,N_10048,N_10959);
nand U13110 (N_13110,N_10115,N_10981);
nor U13111 (N_13111,N_10333,N_10931);
and U13112 (N_13112,N_11928,N_11688);
nor U13113 (N_13113,N_11104,N_10676);
xnor U13114 (N_13114,N_10002,N_10209);
nor U13115 (N_13115,N_11913,N_10318);
and U13116 (N_13116,N_10334,N_11246);
or U13117 (N_13117,N_10794,N_10309);
nand U13118 (N_13118,N_11805,N_11254);
or U13119 (N_13119,N_10937,N_10979);
xnor U13120 (N_13120,N_10738,N_10656);
nand U13121 (N_13121,N_10622,N_11404);
and U13122 (N_13122,N_11899,N_11715);
nand U13123 (N_13123,N_11923,N_11421);
xnor U13124 (N_13124,N_10656,N_11297);
nand U13125 (N_13125,N_10873,N_11761);
xnor U13126 (N_13126,N_10360,N_11200);
nand U13127 (N_13127,N_10933,N_10352);
or U13128 (N_13128,N_10605,N_11546);
nor U13129 (N_13129,N_11662,N_10622);
nor U13130 (N_13130,N_10758,N_10265);
xnor U13131 (N_13131,N_11186,N_11353);
or U13132 (N_13132,N_11306,N_10150);
or U13133 (N_13133,N_11283,N_10960);
nand U13134 (N_13134,N_11719,N_11586);
nand U13135 (N_13135,N_11699,N_10898);
or U13136 (N_13136,N_11680,N_11784);
and U13137 (N_13137,N_11340,N_11019);
xnor U13138 (N_13138,N_11592,N_10880);
nand U13139 (N_13139,N_11104,N_10387);
and U13140 (N_13140,N_11331,N_11847);
xnor U13141 (N_13141,N_10112,N_11510);
xor U13142 (N_13142,N_10142,N_10916);
and U13143 (N_13143,N_10826,N_10910);
xnor U13144 (N_13144,N_11812,N_11539);
or U13145 (N_13145,N_10352,N_10720);
nor U13146 (N_13146,N_10349,N_10526);
xor U13147 (N_13147,N_10177,N_11884);
and U13148 (N_13148,N_11520,N_10253);
xnor U13149 (N_13149,N_11944,N_11002);
nand U13150 (N_13150,N_10337,N_11174);
xor U13151 (N_13151,N_10207,N_10602);
and U13152 (N_13152,N_11179,N_11775);
xor U13153 (N_13153,N_10460,N_10444);
nor U13154 (N_13154,N_11015,N_10988);
or U13155 (N_13155,N_11912,N_10616);
and U13156 (N_13156,N_11104,N_11841);
and U13157 (N_13157,N_11791,N_11112);
nand U13158 (N_13158,N_10427,N_11536);
nand U13159 (N_13159,N_10200,N_11881);
nor U13160 (N_13160,N_11635,N_10498);
nor U13161 (N_13161,N_11553,N_11515);
xnor U13162 (N_13162,N_10593,N_10597);
xnor U13163 (N_13163,N_11764,N_11682);
nor U13164 (N_13164,N_11381,N_11786);
nor U13165 (N_13165,N_10392,N_10156);
nor U13166 (N_13166,N_10000,N_10604);
xor U13167 (N_13167,N_10517,N_11277);
nor U13168 (N_13168,N_10654,N_11017);
nand U13169 (N_13169,N_11525,N_11269);
nor U13170 (N_13170,N_10366,N_10571);
xor U13171 (N_13171,N_10028,N_10375);
xnor U13172 (N_13172,N_10469,N_10028);
and U13173 (N_13173,N_11231,N_10655);
and U13174 (N_13174,N_11964,N_10538);
nor U13175 (N_13175,N_10012,N_10909);
nand U13176 (N_13176,N_10464,N_11248);
xor U13177 (N_13177,N_10490,N_10311);
nand U13178 (N_13178,N_10004,N_10450);
or U13179 (N_13179,N_11537,N_10415);
and U13180 (N_13180,N_11768,N_11602);
nor U13181 (N_13181,N_11337,N_11676);
and U13182 (N_13182,N_10444,N_10125);
and U13183 (N_13183,N_11745,N_10051);
and U13184 (N_13184,N_11662,N_10290);
or U13185 (N_13185,N_10142,N_10392);
nand U13186 (N_13186,N_10984,N_11177);
nor U13187 (N_13187,N_11596,N_11738);
nor U13188 (N_13188,N_11230,N_10075);
nor U13189 (N_13189,N_11098,N_10229);
nor U13190 (N_13190,N_10473,N_11697);
and U13191 (N_13191,N_11785,N_11538);
nand U13192 (N_13192,N_10174,N_10551);
nor U13193 (N_13193,N_11185,N_11026);
or U13194 (N_13194,N_11268,N_10810);
nand U13195 (N_13195,N_10612,N_11880);
nand U13196 (N_13196,N_11764,N_10425);
and U13197 (N_13197,N_11021,N_11720);
xnor U13198 (N_13198,N_11989,N_11736);
or U13199 (N_13199,N_11617,N_10837);
xnor U13200 (N_13200,N_10308,N_10838);
nor U13201 (N_13201,N_11939,N_10457);
xor U13202 (N_13202,N_11902,N_10252);
xnor U13203 (N_13203,N_10424,N_10016);
xnor U13204 (N_13204,N_10582,N_11874);
and U13205 (N_13205,N_11652,N_11161);
nor U13206 (N_13206,N_11486,N_11071);
xnor U13207 (N_13207,N_10743,N_10928);
nor U13208 (N_13208,N_11158,N_11895);
or U13209 (N_13209,N_11207,N_11109);
nor U13210 (N_13210,N_11261,N_11039);
xor U13211 (N_13211,N_10948,N_11853);
and U13212 (N_13212,N_10922,N_11789);
or U13213 (N_13213,N_10148,N_10293);
and U13214 (N_13214,N_11998,N_11369);
nor U13215 (N_13215,N_11997,N_11249);
nand U13216 (N_13216,N_11498,N_11383);
or U13217 (N_13217,N_10185,N_10002);
and U13218 (N_13218,N_10855,N_11913);
nor U13219 (N_13219,N_11365,N_10873);
xnor U13220 (N_13220,N_10989,N_10673);
or U13221 (N_13221,N_10365,N_10581);
or U13222 (N_13222,N_11427,N_10677);
and U13223 (N_13223,N_10191,N_10447);
or U13224 (N_13224,N_11483,N_10891);
xor U13225 (N_13225,N_11862,N_10023);
and U13226 (N_13226,N_10065,N_11189);
nor U13227 (N_13227,N_11494,N_11188);
xor U13228 (N_13228,N_10582,N_11183);
or U13229 (N_13229,N_11772,N_11776);
nand U13230 (N_13230,N_11034,N_11791);
xnor U13231 (N_13231,N_10780,N_11835);
nand U13232 (N_13232,N_10007,N_10312);
nand U13233 (N_13233,N_11594,N_11093);
xor U13234 (N_13234,N_11060,N_10720);
xor U13235 (N_13235,N_10914,N_10808);
or U13236 (N_13236,N_10470,N_10302);
and U13237 (N_13237,N_10673,N_11547);
nand U13238 (N_13238,N_11493,N_11473);
or U13239 (N_13239,N_11134,N_11634);
nand U13240 (N_13240,N_10628,N_11793);
xor U13241 (N_13241,N_10494,N_10629);
and U13242 (N_13242,N_10498,N_10025);
nand U13243 (N_13243,N_11060,N_10407);
and U13244 (N_13244,N_11345,N_11455);
xnor U13245 (N_13245,N_11981,N_10707);
xnor U13246 (N_13246,N_11948,N_10947);
nand U13247 (N_13247,N_10776,N_11784);
nand U13248 (N_13248,N_10348,N_11724);
xor U13249 (N_13249,N_10105,N_11082);
nand U13250 (N_13250,N_10341,N_11011);
xor U13251 (N_13251,N_10404,N_11079);
xnor U13252 (N_13252,N_11282,N_11595);
xor U13253 (N_13253,N_10313,N_11183);
and U13254 (N_13254,N_10527,N_11023);
xor U13255 (N_13255,N_10825,N_10228);
nand U13256 (N_13256,N_10329,N_10459);
nor U13257 (N_13257,N_11096,N_10210);
or U13258 (N_13258,N_11005,N_10811);
nand U13259 (N_13259,N_11229,N_10698);
and U13260 (N_13260,N_11488,N_10244);
or U13261 (N_13261,N_10987,N_10677);
and U13262 (N_13262,N_11144,N_11397);
and U13263 (N_13263,N_11769,N_10780);
and U13264 (N_13264,N_11970,N_10820);
nand U13265 (N_13265,N_10692,N_11192);
and U13266 (N_13266,N_11347,N_11426);
nor U13267 (N_13267,N_10983,N_11824);
and U13268 (N_13268,N_11195,N_10094);
nor U13269 (N_13269,N_10157,N_11816);
or U13270 (N_13270,N_11875,N_11259);
nor U13271 (N_13271,N_10933,N_10115);
and U13272 (N_13272,N_11179,N_10427);
or U13273 (N_13273,N_10756,N_11567);
xor U13274 (N_13274,N_10544,N_11232);
nand U13275 (N_13275,N_10808,N_10807);
or U13276 (N_13276,N_10876,N_11895);
nor U13277 (N_13277,N_10425,N_10630);
nor U13278 (N_13278,N_11960,N_11959);
and U13279 (N_13279,N_10677,N_11738);
and U13280 (N_13280,N_11836,N_10311);
nor U13281 (N_13281,N_10139,N_11539);
or U13282 (N_13282,N_11413,N_11869);
nand U13283 (N_13283,N_11328,N_11317);
and U13284 (N_13284,N_10835,N_10266);
nor U13285 (N_13285,N_10527,N_10624);
xor U13286 (N_13286,N_11602,N_11537);
or U13287 (N_13287,N_11365,N_10664);
and U13288 (N_13288,N_11238,N_11047);
nor U13289 (N_13289,N_10974,N_10756);
or U13290 (N_13290,N_11024,N_11446);
xor U13291 (N_13291,N_11881,N_10632);
and U13292 (N_13292,N_11786,N_11182);
or U13293 (N_13293,N_11985,N_10977);
nor U13294 (N_13294,N_10155,N_10898);
xnor U13295 (N_13295,N_10640,N_10118);
nor U13296 (N_13296,N_11526,N_10355);
or U13297 (N_13297,N_11145,N_11180);
and U13298 (N_13298,N_11112,N_10629);
nor U13299 (N_13299,N_11943,N_10674);
or U13300 (N_13300,N_11382,N_11617);
nor U13301 (N_13301,N_10143,N_10638);
xnor U13302 (N_13302,N_11113,N_11565);
nor U13303 (N_13303,N_10975,N_10065);
xor U13304 (N_13304,N_10963,N_10282);
or U13305 (N_13305,N_10911,N_10279);
or U13306 (N_13306,N_10518,N_10945);
nor U13307 (N_13307,N_10813,N_10774);
nand U13308 (N_13308,N_11601,N_10639);
nor U13309 (N_13309,N_11008,N_11525);
nand U13310 (N_13310,N_11360,N_10604);
nand U13311 (N_13311,N_10717,N_10967);
nor U13312 (N_13312,N_11771,N_11188);
xnor U13313 (N_13313,N_11936,N_10822);
nand U13314 (N_13314,N_11099,N_10852);
or U13315 (N_13315,N_10448,N_10062);
and U13316 (N_13316,N_10098,N_10537);
xor U13317 (N_13317,N_11701,N_11227);
nor U13318 (N_13318,N_11403,N_10175);
nand U13319 (N_13319,N_11155,N_10268);
xor U13320 (N_13320,N_10139,N_10874);
nor U13321 (N_13321,N_11455,N_10298);
nor U13322 (N_13322,N_10846,N_10494);
xor U13323 (N_13323,N_11073,N_10685);
xor U13324 (N_13324,N_10024,N_10145);
nand U13325 (N_13325,N_10530,N_11422);
or U13326 (N_13326,N_11372,N_11458);
nand U13327 (N_13327,N_11511,N_10809);
nand U13328 (N_13328,N_10625,N_11846);
or U13329 (N_13329,N_11649,N_11358);
and U13330 (N_13330,N_11463,N_11737);
xor U13331 (N_13331,N_11948,N_11089);
or U13332 (N_13332,N_11230,N_10919);
and U13333 (N_13333,N_11944,N_11205);
or U13334 (N_13334,N_11637,N_10367);
nor U13335 (N_13335,N_11011,N_10591);
nor U13336 (N_13336,N_11441,N_11523);
nand U13337 (N_13337,N_10196,N_10436);
nand U13338 (N_13338,N_11099,N_10162);
or U13339 (N_13339,N_10270,N_10934);
nor U13340 (N_13340,N_10287,N_10030);
nor U13341 (N_13341,N_11831,N_11165);
nand U13342 (N_13342,N_10461,N_11082);
nor U13343 (N_13343,N_10200,N_11364);
or U13344 (N_13344,N_10108,N_10874);
nand U13345 (N_13345,N_11846,N_10601);
xor U13346 (N_13346,N_11886,N_11925);
or U13347 (N_13347,N_11706,N_10299);
nor U13348 (N_13348,N_10629,N_10076);
or U13349 (N_13349,N_10207,N_10296);
and U13350 (N_13350,N_10417,N_10961);
nor U13351 (N_13351,N_11917,N_11611);
and U13352 (N_13352,N_11250,N_10243);
nor U13353 (N_13353,N_10651,N_11109);
xor U13354 (N_13354,N_10895,N_10524);
nor U13355 (N_13355,N_11645,N_11361);
or U13356 (N_13356,N_11902,N_10167);
nor U13357 (N_13357,N_10106,N_11677);
and U13358 (N_13358,N_10273,N_11947);
nor U13359 (N_13359,N_11395,N_11871);
and U13360 (N_13360,N_11252,N_11067);
xnor U13361 (N_13361,N_10038,N_11433);
and U13362 (N_13362,N_11652,N_11050);
and U13363 (N_13363,N_10069,N_11394);
or U13364 (N_13364,N_11956,N_10981);
xnor U13365 (N_13365,N_11671,N_10453);
xor U13366 (N_13366,N_10822,N_11864);
nor U13367 (N_13367,N_10619,N_10752);
and U13368 (N_13368,N_10630,N_11534);
or U13369 (N_13369,N_10551,N_10305);
and U13370 (N_13370,N_11643,N_10836);
nand U13371 (N_13371,N_11829,N_11551);
and U13372 (N_13372,N_10100,N_11259);
and U13373 (N_13373,N_10569,N_10859);
xnor U13374 (N_13374,N_11051,N_11301);
xor U13375 (N_13375,N_10761,N_11386);
or U13376 (N_13376,N_10783,N_11186);
nor U13377 (N_13377,N_10149,N_11002);
nor U13378 (N_13378,N_10334,N_10574);
or U13379 (N_13379,N_10722,N_11211);
and U13380 (N_13380,N_11993,N_10128);
nor U13381 (N_13381,N_10713,N_11703);
and U13382 (N_13382,N_10680,N_10820);
nor U13383 (N_13383,N_11824,N_11182);
nand U13384 (N_13384,N_11453,N_10702);
nand U13385 (N_13385,N_11134,N_10436);
or U13386 (N_13386,N_10867,N_11943);
nor U13387 (N_13387,N_10212,N_10381);
xor U13388 (N_13388,N_11640,N_10584);
or U13389 (N_13389,N_11376,N_10943);
xor U13390 (N_13390,N_11283,N_10204);
or U13391 (N_13391,N_11879,N_10327);
or U13392 (N_13392,N_11254,N_10588);
nand U13393 (N_13393,N_10114,N_11688);
nand U13394 (N_13394,N_10195,N_11178);
and U13395 (N_13395,N_11185,N_11084);
xor U13396 (N_13396,N_10155,N_10311);
and U13397 (N_13397,N_11993,N_11809);
nand U13398 (N_13398,N_11873,N_11442);
and U13399 (N_13399,N_11609,N_11638);
xnor U13400 (N_13400,N_10915,N_10793);
nand U13401 (N_13401,N_11145,N_10673);
nand U13402 (N_13402,N_11374,N_11202);
and U13403 (N_13403,N_10064,N_10615);
and U13404 (N_13404,N_11865,N_11823);
or U13405 (N_13405,N_10361,N_11537);
and U13406 (N_13406,N_10389,N_11052);
xnor U13407 (N_13407,N_11732,N_10728);
or U13408 (N_13408,N_11304,N_10973);
or U13409 (N_13409,N_11513,N_10381);
nand U13410 (N_13410,N_10396,N_10623);
and U13411 (N_13411,N_10244,N_11504);
and U13412 (N_13412,N_10938,N_10050);
nand U13413 (N_13413,N_11417,N_10116);
nand U13414 (N_13414,N_10935,N_10338);
nand U13415 (N_13415,N_10214,N_11816);
or U13416 (N_13416,N_11961,N_10675);
nand U13417 (N_13417,N_11382,N_10293);
nand U13418 (N_13418,N_11360,N_10265);
nor U13419 (N_13419,N_11419,N_11544);
or U13420 (N_13420,N_10660,N_10301);
nand U13421 (N_13421,N_11301,N_11180);
nand U13422 (N_13422,N_10617,N_10107);
nand U13423 (N_13423,N_11203,N_10959);
nor U13424 (N_13424,N_11120,N_11152);
and U13425 (N_13425,N_10266,N_10071);
nand U13426 (N_13426,N_10974,N_11874);
nor U13427 (N_13427,N_11644,N_11998);
or U13428 (N_13428,N_11470,N_10362);
and U13429 (N_13429,N_11471,N_11988);
nand U13430 (N_13430,N_10793,N_10847);
nand U13431 (N_13431,N_10716,N_10128);
xnor U13432 (N_13432,N_10598,N_10497);
xor U13433 (N_13433,N_11923,N_11825);
and U13434 (N_13434,N_11562,N_11181);
xor U13435 (N_13435,N_11167,N_11570);
nor U13436 (N_13436,N_10409,N_10265);
nor U13437 (N_13437,N_10914,N_11979);
nor U13438 (N_13438,N_10200,N_10198);
nand U13439 (N_13439,N_10887,N_11026);
nand U13440 (N_13440,N_11014,N_10002);
or U13441 (N_13441,N_10938,N_11412);
or U13442 (N_13442,N_10021,N_11946);
xnor U13443 (N_13443,N_11424,N_10265);
nor U13444 (N_13444,N_10712,N_10865);
and U13445 (N_13445,N_10537,N_11113);
or U13446 (N_13446,N_10423,N_11655);
and U13447 (N_13447,N_10381,N_10416);
nand U13448 (N_13448,N_11336,N_11005);
nand U13449 (N_13449,N_11114,N_10133);
xnor U13450 (N_13450,N_10700,N_11391);
and U13451 (N_13451,N_10848,N_11137);
nor U13452 (N_13452,N_10011,N_11518);
nor U13453 (N_13453,N_10844,N_10223);
and U13454 (N_13454,N_10629,N_11323);
nor U13455 (N_13455,N_10963,N_11504);
nor U13456 (N_13456,N_11576,N_10681);
or U13457 (N_13457,N_10629,N_11817);
and U13458 (N_13458,N_11099,N_11946);
and U13459 (N_13459,N_10226,N_10257);
and U13460 (N_13460,N_11528,N_10452);
nand U13461 (N_13461,N_10509,N_11593);
nand U13462 (N_13462,N_11721,N_10719);
nand U13463 (N_13463,N_10762,N_10081);
and U13464 (N_13464,N_10118,N_11827);
nand U13465 (N_13465,N_11562,N_10577);
xor U13466 (N_13466,N_10304,N_10563);
nand U13467 (N_13467,N_10649,N_10433);
or U13468 (N_13468,N_11133,N_10690);
nor U13469 (N_13469,N_10651,N_10661);
xnor U13470 (N_13470,N_11985,N_10167);
nand U13471 (N_13471,N_10680,N_11028);
or U13472 (N_13472,N_10493,N_11151);
nand U13473 (N_13473,N_10484,N_11709);
or U13474 (N_13474,N_10783,N_10518);
nand U13475 (N_13475,N_10942,N_11920);
or U13476 (N_13476,N_11903,N_10298);
nand U13477 (N_13477,N_11330,N_10659);
or U13478 (N_13478,N_10472,N_11276);
and U13479 (N_13479,N_10037,N_11359);
and U13480 (N_13480,N_10180,N_11183);
or U13481 (N_13481,N_10006,N_10966);
or U13482 (N_13482,N_11206,N_11778);
nor U13483 (N_13483,N_11666,N_10477);
xor U13484 (N_13484,N_10202,N_11977);
xor U13485 (N_13485,N_10203,N_11254);
and U13486 (N_13486,N_11093,N_10059);
and U13487 (N_13487,N_10249,N_11029);
nor U13488 (N_13488,N_10970,N_11396);
and U13489 (N_13489,N_11887,N_11993);
nand U13490 (N_13490,N_10765,N_10177);
or U13491 (N_13491,N_10416,N_11608);
nor U13492 (N_13492,N_11647,N_10151);
nand U13493 (N_13493,N_11070,N_11451);
nand U13494 (N_13494,N_11242,N_11045);
or U13495 (N_13495,N_10565,N_11312);
nor U13496 (N_13496,N_10003,N_11092);
nor U13497 (N_13497,N_10605,N_10829);
nor U13498 (N_13498,N_11564,N_10977);
nor U13499 (N_13499,N_11156,N_10434);
and U13500 (N_13500,N_11903,N_11301);
nand U13501 (N_13501,N_10672,N_11407);
nand U13502 (N_13502,N_10449,N_10843);
xor U13503 (N_13503,N_10997,N_10938);
and U13504 (N_13504,N_11886,N_10317);
and U13505 (N_13505,N_10226,N_11516);
and U13506 (N_13506,N_10718,N_11289);
nand U13507 (N_13507,N_11431,N_11752);
nand U13508 (N_13508,N_11288,N_11108);
xnor U13509 (N_13509,N_10955,N_11386);
and U13510 (N_13510,N_10280,N_10888);
nand U13511 (N_13511,N_10237,N_10594);
or U13512 (N_13512,N_10308,N_11033);
and U13513 (N_13513,N_11639,N_10392);
and U13514 (N_13514,N_10625,N_10730);
nand U13515 (N_13515,N_11722,N_10800);
or U13516 (N_13516,N_10924,N_11121);
and U13517 (N_13517,N_10221,N_10342);
or U13518 (N_13518,N_10314,N_10032);
or U13519 (N_13519,N_10891,N_11901);
nand U13520 (N_13520,N_10624,N_10517);
or U13521 (N_13521,N_11977,N_10099);
nor U13522 (N_13522,N_11203,N_10821);
nor U13523 (N_13523,N_11202,N_11395);
or U13524 (N_13524,N_11844,N_10302);
xor U13525 (N_13525,N_11872,N_10114);
and U13526 (N_13526,N_10092,N_10331);
nand U13527 (N_13527,N_11408,N_11880);
nand U13528 (N_13528,N_10978,N_10334);
and U13529 (N_13529,N_11827,N_10187);
xor U13530 (N_13530,N_10880,N_10095);
and U13531 (N_13531,N_10694,N_10589);
and U13532 (N_13532,N_11588,N_11783);
or U13533 (N_13533,N_10569,N_11629);
xnor U13534 (N_13534,N_10041,N_10477);
nand U13535 (N_13535,N_11223,N_11731);
and U13536 (N_13536,N_11985,N_10658);
xor U13537 (N_13537,N_11234,N_10232);
nor U13538 (N_13538,N_10233,N_11192);
nor U13539 (N_13539,N_11526,N_11518);
nor U13540 (N_13540,N_10746,N_11458);
or U13541 (N_13541,N_11808,N_11398);
and U13542 (N_13542,N_11094,N_11904);
xnor U13543 (N_13543,N_11198,N_11407);
or U13544 (N_13544,N_11678,N_10309);
nor U13545 (N_13545,N_10753,N_10583);
nor U13546 (N_13546,N_11137,N_10068);
nor U13547 (N_13547,N_10345,N_10608);
xnor U13548 (N_13548,N_11710,N_10512);
nor U13549 (N_13549,N_11249,N_11386);
or U13550 (N_13550,N_10985,N_10876);
xor U13551 (N_13551,N_11628,N_10129);
xnor U13552 (N_13552,N_11831,N_11843);
nand U13553 (N_13553,N_10443,N_10765);
xnor U13554 (N_13554,N_10906,N_10363);
xnor U13555 (N_13555,N_10830,N_10102);
or U13556 (N_13556,N_10181,N_10362);
nand U13557 (N_13557,N_10632,N_11625);
xor U13558 (N_13558,N_11091,N_10253);
nand U13559 (N_13559,N_10803,N_10743);
and U13560 (N_13560,N_11703,N_10749);
nor U13561 (N_13561,N_10059,N_10823);
nor U13562 (N_13562,N_10929,N_11290);
or U13563 (N_13563,N_10272,N_11382);
xnor U13564 (N_13564,N_11619,N_11599);
nand U13565 (N_13565,N_11812,N_11567);
nand U13566 (N_13566,N_11978,N_10205);
xor U13567 (N_13567,N_11183,N_10709);
nand U13568 (N_13568,N_10631,N_10948);
nor U13569 (N_13569,N_10044,N_11128);
nor U13570 (N_13570,N_11104,N_11131);
or U13571 (N_13571,N_10891,N_10267);
or U13572 (N_13572,N_11197,N_10690);
and U13573 (N_13573,N_11290,N_11344);
or U13574 (N_13574,N_10530,N_11620);
nand U13575 (N_13575,N_10788,N_10582);
nand U13576 (N_13576,N_10625,N_10796);
or U13577 (N_13577,N_11778,N_11789);
or U13578 (N_13578,N_11936,N_11594);
nor U13579 (N_13579,N_10652,N_11563);
and U13580 (N_13580,N_10299,N_11898);
xnor U13581 (N_13581,N_11110,N_10282);
nor U13582 (N_13582,N_10486,N_11137);
nor U13583 (N_13583,N_11986,N_10390);
or U13584 (N_13584,N_10567,N_10289);
xnor U13585 (N_13585,N_11134,N_11750);
and U13586 (N_13586,N_10786,N_11534);
xor U13587 (N_13587,N_11655,N_11850);
nor U13588 (N_13588,N_10808,N_11788);
and U13589 (N_13589,N_11733,N_11303);
nor U13590 (N_13590,N_10360,N_10730);
and U13591 (N_13591,N_11423,N_10725);
nor U13592 (N_13592,N_11508,N_11541);
nand U13593 (N_13593,N_11639,N_11545);
nor U13594 (N_13594,N_10957,N_10649);
nand U13595 (N_13595,N_11245,N_11384);
nand U13596 (N_13596,N_10071,N_11960);
and U13597 (N_13597,N_10179,N_10998);
xor U13598 (N_13598,N_10769,N_10316);
nand U13599 (N_13599,N_11592,N_11237);
xnor U13600 (N_13600,N_11488,N_10902);
xnor U13601 (N_13601,N_10362,N_11416);
or U13602 (N_13602,N_11895,N_10941);
nor U13603 (N_13603,N_10174,N_10796);
nand U13604 (N_13604,N_10839,N_11450);
or U13605 (N_13605,N_11526,N_10797);
nand U13606 (N_13606,N_11258,N_11215);
nor U13607 (N_13607,N_11681,N_11444);
xnor U13608 (N_13608,N_10884,N_11643);
nand U13609 (N_13609,N_11305,N_11089);
nor U13610 (N_13610,N_11129,N_11739);
nand U13611 (N_13611,N_10785,N_11571);
nand U13612 (N_13612,N_10098,N_11524);
nand U13613 (N_13613,N_10617,N_11382);
nand U13614 (N_13614,N_11674,N_11256);
xnor U13615 (N_13615,N_10669,N_11300);
or U13616 (N_13616,N_11726,N_11718);
nor U13617 (N_13617,N_11413,N_10635);
and U13618 (N_13618,N_10661,N_11404);
or U13619 (N_13619,N_10930,N_10157);
nor U13620 (N_13620,N_11081,N_10035);
and U13621 (N_13621,N_11705,N_11589);
xor U13622 (N_13622,N_11751,N_10521);
xnor U13623 (N_13623,N_11450,N_11116);
and U13624 (N_13624,N_11140,N_11069);
and U13625 (N_13625,N_11319,N_11504);
nor U13626 (N_13626,N_11104,N_10116);
or U13627 (N_13627,N_11116,N_10214);
or U13628 (N_13628,N_10244,N_10744);
xor U13629 (N_13629,N_11926,N_11067);
or U13630 (N_13630,N_10627,N_10530);
nor U13631 (N_13631,N_10251,N_11878);
nand U13632 (N_13632,N_10359,N_10111);
and U13633 (N_13633,N_11923,N_10683);
xor U13634 (N_13634,N_10296,N_11936);
or U13635 (N_13635,N_10108,N_11844);
nand U13636 (N_13636,N_11739,N_11341);
nand U13637 (N_13637,N_11494,N_11116);
nand U13638 (N_13638,N_11606,N_11009);
and U13639 (N_13639,N_10728,N_11451);
and U13640 (N_13640,N_10805,N_10972);
xnor U13641 (N_13641,N_10043,N_10757);
or U13642 (N_13642,N_11217,N_11787);
nand U13643 (N_13643,N_11790,N_11591);
or U13644 (N_13644,N_11746,N_10497);
and U13645 (N_13645,N_10914,N_11538);
nor U13646 (N_13646,N_11247,N_10937);
nand U13647 (N_13647,N_10455,N_11023);
nor U13648 (N_13648,N_10048,N_11339);
or U13649 (N_13649,N_10541,N_11306);
nand U13650 (N_13650,N_10891,N_10508);
or U13651 (N_13651,N_10385,N_10836);
or U13652 (N_13652,N_10517,N_10989);
xnor U13653 (N_13653,N_10494,N_11573);
xnor U13654 (N_13654,N_10899,N_10192);
and U13655 (N_13655,N_10363,N_10837);
xnor U13656 (N_13656,N_11999,N_11980);
xor U13657 (N_13657,N_10151,N_10558);
nor U13658 (N_13658,N_11839,N_10195);
xor U13659 (N_13659,N_11674,N_10810);
or U13660 (N_13660,N_11825,N_10532);
nor U13661 (N_13661,N_11154,N_10163);
nand U13662 (N_13662,N_10765,N_11021);
xnor U13663 (N_13663,N_10738,N_11186);
and U13664 (N_13664,N_10711,N_10780);
or U13665 (N_13665,N_11244,N_11755);
xor U13666 (N_13666,N_10918,N_10089);
or U13667 (N_13667,N_11052,N_11925);
nand U13668 (N_13668,N_10515,N_11907);
xnor U13669 (N_13669,N_11659,N_10212);
and U13670 (N_13670,N_11813,N_11423);
nand U13671 (N_13671,N_11771,N_10768);
xnor U13672 (N_13672,N_10370,N_10043);
xnor U13673 (N_13673,N_10062,N_11732);
xnor U13674 (N_13674,N_10270,N_11842);
or U13675 (N_13675,N_11834,N_10673);
xor U13676 (N_13676,N_10954,N_10475);
xnor U13677 (N_13677,N_11497,N_11243);
xnor U13678 (N_13678,N_11916,N_11732);
xnor U13679 (N_13679,N_11949,N_10686);
and U13680 (N_13680,N_11693,N_11677);
and U13681 (N_13681,N_10083,N_10992);
or U13682 (N_13682,N_10844,N_11080);
and U13683 (N_13683,N_11583,N_10220);
or U13684 (N_13684,N_11686,N_10676);
nand U13685 (N_13685,N_10512,N_10734);
or U13686 (N_13686,N_11695,N_10268);
nor U13687 (N_13687,N_10079,N_11497);
nor U13688 (N_13688,N_10810,N_10152);
nand U13689 (N_13689,N_10656,N_11925);
and U13690 (N_13690,N_11788,N_11878);
and U13691 (N_13691,N_11918,N_10213);
xnor U13692 (N_13692,N_11958,N_11687);
nor U13693 (N_13693,N_10340,N_11779);
nor U13694 (N_13694,N_11666,N_11162);
nor U13695 (N_13695,N_10862,N_10814);
and U13696 (N_13696,N_11579,N_10431);
xnor U13697 (N_13697,N_10590,N_11460);
nor U13698 (N_13698,N_10855,N_10390);
xnor U13699 (N_13699,N_10112,N_10133);
nand U13700 (N_13700,N_10905,N_11184);
nand U13701 (N_13701,N_11052,N_10744);
nor U13702 (N_13702,N_10625,N_10005);
nor U13703 (N_13703,N_10204,N_11862);
and U13704 (N_13704,N_11682,N_10539);
or U13705 (N_13705,N_11918,N_11913);
nand U13706 (N_13706,N_11066,N_11344);
nand U13707 (N_13707,N_11647,N_11484);
and U13708 (N_13708,N_10323,N_10099);
nor U13709 (N_13709,N_11739,N_10931);
xor U13710 (N_13710,N_11603,N_10402);
or U13711 (N_13711,N_10747,N_11801);
nor U13712 (N_13712,N_10727,N_11133);
xnor U13713 (N_13713,N_10724,N_11356);
and U13714 (N_13714,N_10095,N_11803);
nor U13715 (N_13715,N_11757,N_11736);
or U13716 (N_13716,N_10857,N_11468);
and U13717 (N_13717,N_11509,N_11552);
nor U13718 (N_13718,N_10585,N_11900);
and U13719 (N_13719,N_11045,N_11067);
and U13720 (N_13720,N_11117,N_10127);
and U13721 (N_13721,N_11592,N_11961);
xor U13722 (N_13722,N_10902,N_10968);
xor U13723 (N_13723,N_11956,N_10029);
nand U13724 (N_13724,N_11297,N_10749);
nand U13725 (N_13725,N_10251,N_11005);
nand U13726 (N_13726,N_11370,N_10615);
and U13727 (N_13727,N_10174,N_11530);
nor U13728 (N_13728,N_10818,N_10837);
and U13729 (N_13729,N_11598,N_11765);
xor U13730 (N_13730,N_11341,N_10721);
xnor U13731 (N_13731,N_10016,N_10136);
and U13732 (N_13732,N_10291,N_10443);
xnor U13733 (N_13733,N_11749,N_11042);
nor U13734 (N_13734,N_10925,N_11018);
and U13735 (N_13735,N_11242,N_11955);
nand U13736 (N_13736,N_11123,N_11578);
nor U13737 (N_13737,N_11969,N_10637);
nand U13738 (N_13738,N_11226,N_11180);
nor U13739 (N_13739,N_10379,N_11941);
nand U13740 (N_13740,N_11519,N_11370);
nor U13741 (N_13741,N_10277,N_11508);
and U13742 (N_13742,N_11513,N_10729);
or U13743 (N_13743,N_11045,N_11130);
nor U13744 (N_13744,N_11912,N_11467);
nand U13745 (N_13745,N_11286,N_11501);
nor U13746 (N_13746,N_11308,N_11798);
nor U13747 (N_13747,N_10693,N_10528);
xor U13748 (N_13748,N_10945,N_11761);
nand U13749 (N_13749,N_11786,N_11524);
or U13750 (N_13750,N_11521,N_11003);
nand U13751 (N_13751,N_11829,N_10692);
xnor U13752 (N_13752,N_11972,N_11363);
and U13753 (N_13753,N_11800,N_11338);
xnor U13754 (N_13754,N_10000,N_10979);
nand U13755 (N_13755,N_10701,N_11881);
and U13756 (N_13756,N_11794,N_11219);
nor U13757 (N_13757,N_10656,N_11121);
and U13758 (N_13758,N_11845,N_10512);
or U13759 (N_13759,N_11775,N_10091);
nor U13760 (N_13760,N_11785,N_11701);
nand U13761 (N_13761,N_11639,N_11753);
xor U13762 (N_13762,N_10256,N_11846);
and U13763 (N_13763,N_11664,N_10646);
nand U13764 (N_13764,N_11697,N_11495);
nand U13765 (N_13765,N_11312,N_11911);
nor U13766 (N_13766,N_10468,N_11225);
xnor U13767 (N_13767,N_10889,N_10822);
nand U13768 (N_13768,N_10954,N_10316);
or U13769 (N_13769,N_11456,N_11863);
or U13770 (N_13770,N_11948,N_10135);
or U13771 (N_13771,N_11618,N_10078);
and U13772 (N_13772,N_10337,N_11905);
xor U13773 (N_13773,N_11206,N_10809);
xnor U13774 (N_13774,N_11857,N_11424);
or U13775 (N_13775,N_11168,N_11967);
or U13776 (N_13776,N_11755,N_10548);
nand U13777 (N_13777,N_10763,N_10433);
or U13778 (N_13778,N_11166,N_11890);
or U13779 (N_13779,N_10712,N_10052);
nor U13780 (N_13780,N_10523,N_11566);
nand U13781 (N_13781,N_11933,N_10352);
nand U13782 (N_13782,N_10216,N_11781);
and U13783 (N_13783,N_11567,N_10617);
xnor U13784 (N_13784,N_11038,N_10902);
nor U13785 (N_13785,N_10835,N_10224);
nor U13786 (N_13786,N_11837,N_11416);
and U13787 (N_13787,N_11074,N_11634);
xor U13788 (N_13788,N_11007,N_11951);
xnor U13789 (N_13789,N_10098,N_11697);
and U13790 (N_13790,N_11943,N_10541);
xnor U13791 (N_13791,N_10379,N_10617);
nand U13792 (N_13792,N_10155,N_10810);
or U13793 (N_13793,N_10514,N_11139);
xor U13794 (N_13794,N_11794,N_10561);
or U13795 (N_13795,N_11064,N_11091);
nor U13796 (N_13796,N_10892,N_10818);
nand U13797 (N_13797,N_10504,N_10554);
xnor U13798 (N_13798,N_10639,N_11524);
or U13799 (N_13799,N_11902,N_10064);
or U13800 (N_13800,N_11147,N_10258);
and U13801 (N_13801,N_11021,N_10486);
nor U13802 (N_13802,N_10515,N_10609);
or U13803 (N_13803,N_11881,N_11924);
nand U13804 (N_13804,N_11813,N_11290);
and U13805 (N_13805,N_10201,N_10618);
nor U13806 (N_13806,N_10997,N_10485);
and U13807 (N_13807,N_11868,N_10460);
xor U13808 (N_13808,N_10181,N_11025);
or U13809 (N_13809,N_11710,N_10343);
or U13810 (N_13810,N_11795,N_11242);
or U13811 (N_13811,N_10928,N_11816);
nor U13812 (N_13812,N_11311,N_11151);
nor U13813 (N_13813,N_10266,N_10503);
or U13814 (N_13814,N_11168,N_11676);
xnor U13815 (N_13815,N_11555,N_10526);
nor U13816 (N_13816,N_10485,N_11898);
or U13817 (N_13817,N_10122,N_10698);
xnor U13818 (N_13818,N_10374,N_10565);
nand U13819 (N_13819,N_10052,N_11567);
nor U13820 (N_13820,N_11942,N_11512);
or U13821 (N_13821,N_10417,N_11543);
nand U13822 (N_13822,N_10121,N_11496);
xnor U13823 (N_13823,N_10259,N_11629);
nand U13824 (N_13824,N_11004,N_11953);
xnor U13825 (N_13825,N_10421,N_11313);
xor U13826 (N_13826,N_10698,N_10996);
and U13827 (N_13827,N_11030,N_11764);
xor U13828 (N_13828,N_10022,N_10754);
and U13829 (N_13829,N_11842,N_11426);
or U13830 (N_13830,N_11020,N_10452);
and U13831 (N_13831,N_11815,N_11703);
xnor U13832 (N_13832,N_10507,N_11003);
nor U13833 (N_13833,N_10167,N_10054);
xor U13834 (N_13834,N_10406,N_10308);
nor U13835 (N_13835,N_11504,N_11515);
nand U13836 (N_13836,N_10059,N_10220);
nor U13837 (N_13837,N_11822,N_11133);
and U13838 (N_13838,N_11915,N_10223);
nor U13839 (N_13839,N_11691,N_11374);
nor U13840 (N_13840,N_11824,N_11115);
nor U13841 (N_13841,N_10833,N_11474);
xnor U13842 (N_13842,N_11661,N_11234);
xnor U13843 (N_13843,N_11969,N_11993);
nor U13844 (N_13844,N_10766,N_10045);
or U13845 (N_13845,N_10602,N_11188);
nand U13846 (N_13846,N_10685,N_10086);
nand U13847 (N_13847,N_11690,N_10099);
xnor U13848 (N_13848,N_11928,N_11713);
xor U13849 (N_13849,N_10761,N_11147);
and U13850 (N_13850,N_11043,N_11671);
xnor U13851 (N_13851,N_10278,N_11591);
or U13852 (N_13852,N_10267,N_10626);
xnor U13853 (N_13853,N_10568,N_11321);
or U13854 (N_13854,N_10357,N_10106);
or U13855 (N_13855,N_10807,N_10912);
and U13856 (N_13856,N_11655,N_11064);
nor U13857 (N_13857,N_10624,N_10057);
nor U13858 (N_13858,N_10501,N_11426);
and U13859 (N_13859,N_11518,N_10682);
nor U13860 (N_13860,N_11017,N_11587);
or U13861 (N_13861,N_10517,N_10691);
xnor U13862 (N_13862,N_10024,N_11226);
and U13863 (N_13863,N_10226,N_10569);
and U13864 (N_13864,N_11189,N_11571);
nand U13865 (N_13865,N_10081,N_11506);
and U13866 (N_13866,N_10070,N_11470);
nand U13867 (N_13867,N_10766,N_11440);
nor U13868 (N_13868,N_10739,N_10227);
nand U13869 (N_13869,N_11847,N_11051);
or U13870 (N_13870,N_11441,N_11557);
xor U13871 (N_13871,N_10848,N_11064);
and U13872 (N_13872,N_10543,N_11422);
nand U13873 (N_13873,N_11346,N_11467);
or U13874 (N_13874,N_11708,N_10002);
xor U13875 (N_13875,N_10106,N_10576);
and U13876 (N_13876,N_11966,N_10538);
nor U13877 (N_13877,N_11006,N_10369);
nand U13878 (N_13878,N_11815,N_11768);
and U13879 (N_13879,N_11798,N_11092);
nand U13880 (N_13880,N_11655,N_11071);
nand U13881 (N_13881,N_11888,N_10092);
nand U13882 (N_13882,N_11740,N_10842);
and U13883 (N_13883,N_10609,N_11827);
or U13884 (N_13884,N_10176,N_11414);
and U13885 (N_13885,N_10694,N_11940);
and U13886 (N_13886,N_10847,N_10632);
nor U13887 (N_13887,N_10143,N_11056);
nand U13888 (N_13888,N_10146,N_11419);
or U13889 (N_13889,N_11203,N_10711);
or U13890 (N_13890,N_11190,N_11595);
and U13891 (N_13891,N_11578,N_11472);
or U13892 (N_13892,N_10417,N_11562);
nand U13893 (N_13893,N_10685,N_11706);
xor U13894 (N_13894,N_11197,N_11394);
xor U13895 (N_13895,N_11387,N_11445);
xor U13896 (N_13896,N_10072,N_10329);
and U13897 (N_13897,N_10065,N_11434);
and U13898 (N_13898,N_10348,N_10947);
nand U13899 (N_13899,N_11448,N_11500);
nand U13900 (N_13900,N_10265,N_10318);
and U13901 (N_13901,N_10483,N_10103);
xor U13902 (N_13902,N_10296,N_10323);
nor U13903 (N_13903,N_10160,N_10369);
or U13904 (N_13904,N_10520,N_10889);
nor U13905 (N_13905,N_11447,N_11767);
xor U13906 (N_13906,N_11563,N_11452);
xnor U13907 (N_13907,N_10182,N_11031);
nand U13908 (N_13908,N_10114,N_11572);
xor U13909 (N_13909,N_11100,N_11607);
nor U13910 (N_13910,N_11467,N_11473);
nand U13911 (N_13911,N_10394,N_10738);
nand U13912 (N_13912,N_10020,N_10760);
nand U13913 (N_13913,N_11876,N_10380);
nand U13914 (N_13914,N_10184,N_10765);
nand U13915 (N_13915,N_11469,N_11188);
nor U13916 (N_13916,N_11362,N_10241);
or U13917 (N_13917,N_11934,N_11912);
nand U13918 (N_13918,N_11079,N_10845);
or U13919 (N_13919,N_11361,N_10966);
nor U13920 (N_13920,N_11128,N_11654);
xnor U13921 (N_13921,N_11421,N_10449);
xnor U13922 (N_13922,N_11297,N_10679);
and U13923 (N_13923,N_10489,N_10545);
nand U13924 (N_13924,N_11977,N_11359);
nand U13925 (N_13925,N_10839,N_11571);
nand U13926 (N_13926,N_11832,N_11663);
or U13927 (N_13927,N_11001,N_10447);
and U13928 (N_13928,N_10591,N_10310);
or U13929 (N_13929,N_11415,N_11851);
nand U13930 (N_13930,N_10950,N_11244);
or U13931 (N_13931,N_10256,N_11690);
xnor U13932 (N_13932,N_11328,N_11285);
and U13933 (N_13933,N_11421,N_10814);
xnor U13934 (N_13934,N_10334,N_11468);
xor U13935 (N_13935,N_11263,N_11417);
xor U13936 (N_13936,N_10912,N_11206);
xor U13937 (N_13937,N_10118,N_11610);
xnor U13938 (N_13938,N_10855,N_10083);
or U13939 (N_13939,N_10133,N_10755);
nand U13940 (N_13940,N_11945,N_10133);
xnor U13941 (N_13941,N_10814,N_11803);
nand U13942 (N_13942,N_11480,N_10903);
nand U13943 (N_13943,N_11078,N_10607);
nand U13944 (N_13944,N_10867,N_11244);
nor U13945 (N_13945,N_11124,N_10182);
xnor U13946 (N_13946,N_11213,N_11081);
or U13947 (N_13947,N_10191,N_10378);
or U13948 (N_13948,N_11235,N_10657);
or U13949 (N_13949,N_11226,N_11918);
xnor U13950 (N_13950,N_10981,N_11519);
nand U13951 (N_13951,N_11025,N_10939);
or U13952 (N_13952,N_11010,N_11213);
and U13953 (N_13953,N_10318,N_11746);
or U13954 (N_13954,N_10942,N_11283);
nor U13955 (N_13955,N_10306,N_11607);
or U13956 (N_13956,N_11900,N_10618);
nand U13957 (N_13957,N_11489,N_10018);
and U13958 (N_13958,N_10245,N_10418);
xnor U13959 (N_13959,N_10715,N_10570);
nor U13960 (N_13960,N_11256,N_10929);
nor U13961 (N_13961,N_10268,N_11409);
and U13962 (N_13962,N_11960,N_10226);
nor U13963 (N_13963,N_11298,N_11066);
nor U13964 (N_13964,N_11820,N_11313);
xnor U13965 (N_13965,N_10004,N_11002);
or U13966 (N_13966,N_10432,N_10711);
and U13967 (N_13967,N_11196,N_11917);
nand U13968 (N_13968,N_10230,N_10521);
nor U13969 (N_13969,N_11691,N_11701);
nand U13970 (N_13970,N_10471,N_10900);
xor U13971 (N_13971,N_10655,N_10158);
and U13972 (N_13972,N_11904,N_10349);
or U13973 (N_13973,N_10991,N_10457);
and U13974 (N_13974,N_10054,N_10588);
and U13975 (N_13975,N_10524,N_10043);
nor U13976 (N_13976,N_11358,N_11122);
nor U13977 (N_13977,N_10878,N_10268);
nand U13978 (N_13978,N_11899,N_10267);
or U13979 (N_13979,N_11364,N_11083);
xor U13980 (N_13980,N_11852,N_10151);
and U13981 (N_13981,N_10759,N_10496);
or U13982 (N_13982,N_10855,N_10253);
or U13983 (N_13983,N_11482,N_10384);
nor U13984 (N_13984,N_10048,N_11695);
or U13985 (N_13985,N_10434,N_10713);
nand U13986 (N_13986,N_11043,N_10404);
and U13987 (N_13987,N_10924,N_10123);
nand U13988 (N_13988,N_10348,N_11256);
nor U13989 (N_13989,N_10643,N_11011);
nand U13990 (N_13990,N_11989,N_11888);
nor U13991 (N_13991,N_11511,N_10210);
nor U13992 (N_13992,N_11364,N_10636);
or U13993 (N_13993,N_11099,N_10052);
nor U13994 (N_13994,N_11819,N_10683);
and U13995 (N_13995,N_11365,N_10206);
and U13996 (N_13996,N_10202,N_11504);
nand U13997 (N_13997,N_10418,N_10539);
nand U13998 (N_13998,N_10217,N_11769);
nor U13999 (N_13999,N_11641,N_11976);
or U14000 (N_14000,N_13515,N_12782);
and U14001 (N_14001,N_13634,N_12889);
and U14002 (N_14002,N_13955,N_13494);
nor U14003 (N_14003,N_12699,N_13421);
nand U14004 (N_14004,N_13207,N_12125);
nor U14005 (N_14005,N_13740,N_13474);
nor U14006 (N_14006,N_13298,N_13963);
or U14007 (N_14007,N_12233,N_13813);
nand U14008 (N_14008,N_12498,N_13423);
and U14009 (N_14009,N_13417,N_12179);
nand U14010 (N_14010,N_13310,N_12249);
xor U14011 (N_14011,N_13028,N_12718);
or U14012 (N_14012,N_13873,N_12381);
or U14013 (N_14013,N_13777,N_13383);
and U14014 (N_14014,N_12823,N_12982);
or U14015 (N_14015,N_12645,N_13610);
and U14016 (N_14016,N_12225,N_12892);
or U14017 (N_14017,N_13734,N_13859);
and U14018 (N_14018,N_13018,N_13342);
and U14019 (N_14019,N_13010,N_13198);
or U14020 (N_14020,N_13825,N_12956);
or U14021 (N_14021,N_13792,N_13576);
nand U14022 (N_14022,N_12988,N_13228);
nand U14023 (N_14023,N_13640,N_12829);
nand U14024 (N_14024,N_12993,N_12375);
nor U14025 (N_14025,N_13560,N_12084);
and U14026 (N_14026,N_12634,N_12974);
and U14027 (N_14027,N_13573,N_12041);
nand U14028 (N_14028,N_12262,N_13622);
and U14029 (N_14029,N_12131,N_13781);
or U14030 (N_14030,N_13375,N_13350);
and U14031 (N_14031,N_13492,N_13993);
and U14032 (N_14032,N_13325,N_13346);
xor U14033 (N_14033,N_12414,N_13916);
and U14034 (N_14034,N_13655,N_12399);
xnor U14035 (N_14035,N_13169,N_13946);
or U14036 (N_14036,N_13901,N_13518);
or U14037 (N_14037,N_12261,N_13351);
nor U14038 (N_14038,N_13508,N_12919);
and U14039 (N_14039,N_13312,N_12208);
nor U14040 (N_14040,N_12203,N_13378);
or U14041 (N_14041,N_12296,N_13373);
or U14042 (N_14042,N_12390,N_12006);
nand U14043 (N_14043,N_12142,N_13763);
or U14044 (N_14044,N_13087,N_12001);
nand U14045 (N_14045,N_13209,N_12424);
nor U14046 (N_14046,N_13776,N_13539);
nor U14047 (N_14047,N_12873,N_12469);
or U14048 (N_14048,N_12692,N_13775);
nor U14049 (N_14049,N_13224,N_12513);
xnor U14050 (N_14050,N_13270,N_12326);
nor U14051 (N_14051,N_13819,N_12547);
and U14052 (N_14052,N_13858,N_12644);
nor U14053 (N_14053,N_13554,N_12015);
xnor U14054 (N_14054,N_13773,N_12906);
or U14055 (N_14055,N_12039,N_13048);
or U14056 (N_14056,N_13960,N_13358);
xnor U14057 (N_14057,N_12525,N_13709);
or U14058 (N_14058,N_13550,N_13355);
and U14059 (N_14059,N_12031,N_13000);
nand U14060 (N_14060,N_13121,N_13448);
or U14061 (N_14061,N_12394,N_13532);
or U14062 (N_14062,N_12463,N_13432);
and U14063 (N_14063,N_13076,N_12653);
nand U14064 (N_14064,N_13103,N_12351);
nor U14065 (N_14065,N_12839,N_13670);
xnor U14066 (N_14066,N_13957,N_13142);
nand U14067 (N_14067,N_12675,N_13931);
nor U14068 (N_14068,N_12279,N_12449);
nor U14069 (N_14069,N_12247,N_12470);
and U14070 (N_14070,N_13976,N_13639);
and U14071 (N_14071,N_13745,N_13045);
and U14072 (N_14072,N_12447,N_12794);
or U14073 (N_14073,N_12013,N_12243);
and U14074 (N_14074,N_13463,N_13767);
nand U14075 (N_14075,N_12908,N_12552);
xor U14076 (N_14076,N_13766,N_12206);
nand U14077 (N_14077,N_13537,N_13031);
nor U14078 (N_14078,N_12884,N_13185);
nor U14079 (N_14079,N_12132,N_13132);
nor U14080 (N_14080,N_12940,N_13923);
xnor U14081 (N_14081,N_13283,N_12727);
nor U14082 (N_14082,N_12722,N_13687);
nor U14083 (N_14083,N_13362,N_13799);
nor U14084 (N_14084,N_12489,N_12978);
xor U14085 (N_14085,N_12454,N_12952);
or U14086 (N_14086,N_12866,N_12253);
xor U14087 (N_14087,N_12932,N_13036);
nand U14088 (N_14088,N_12330,N_12274);
nor U14089 (N_14089,N_12056,N_12746);
and U14090 (N_14090,N_12964,N_12744);
xnor U14091 (N_14091,N_12711,N_12098);
and U14092 (N_14092,N_12314,N_12539);
nand U14093 (N_14093,N_13762,N_12079);
and U14094 (N_14094,N_12044,N_12849);
and U14095 (N_14095,N_13262,N_13829);
nand U14096 (N_14096,N_12370,N_13951);
and U14097 (N_14097,N_12104,N_13144);
and U14098 (N_14098,N_13961,N_13703);
nor U14099 (N_14099,N_12604,N_12648);
nor U14100 (N_14100,N_12074,N_12704);
nand U14101 (N_14101,N_13086,N_13305);
nand U14102 (N_14102,N_13319,N_12875);
or U14103 (N_14103,N_12112,N_12834);
nand U14104 (N_14104,N_13197,N_13252);
xnor U14105 (N_14105,N_13027,N_13435);
nand U14106 (N_14106,N_12021,N_13221);
and U14107 (N_14107,N_13941,N_12459);
and U14108 (N_14108,N_13746,N_13314);
xor U14109 (N_14109,N_13327,N_13743);
and U14110 (N_14110,N_13807,N_12462);
and U14111 (N_14111,N_12676,N_13187);
nor U14112 (N_14112,N_13764,N_12628);
xor U14113 (N_14113,N_13876,N_12357);
nor U14114 (N_14114,N_12791,N_12569);
xor U14115 (N_14115,N_13968,N_12743);
nor U14116 (N_14116,N_12771,N_12780);
nor U14117 (N_14117,N_12979,N_13316);
xor U14118 (N_14118,N_13279,N_12384);
xor U14119 (N_14119,N_13893,N_12555);
xnor U14120 (N_14120,N_13973,N_12936);
xnor U14121 (N_14121,N_13296,N_12923);
xor U14122 (N_14122,N_12290,N_12788);
or U14123 (N_14123,N_13101,N_12587);
xnor U14124 (N_14124,N_13694,N_13225);
and U14125 (N_14125,N_12511,N_13013);
and U14126 (N_14126,N_12325,N_13587);
or U14127 (N_14127,N_13604,N_13301);
nor U14128 (N_14128,N_13927,N_12848);
and U14129 (N_14129,N_13843,N_12717);
nor U14130 (N_14130,N_12755,N_12003);
nand U14131 (N_14131,N_12761,N_12741);
xor U14132 (N_14132,N_13393,N_12052);
xnor U14133 (N_14133,N_12911,N_13870);
nand U14134 (N_14134,N_12629,N_12081);
and U14135 (N_14135,N_12561,N_13970);
nand U14136 (N_14136,N_13281,N_12825);
nand U14137 (N_14137,N_12205,N_12775);
nand U14138 (N_14138,N_13735,N_13832);
and U14139 (N_14139,N_13713,N_12655);
nor U14140 (N_14140,N_12385,N_13881);
nor U14141 (N_14141,N_13966,N_12963);
xnor U14142 (N_14142,N_13820,N_12302);
xor U14143 (N_14143,N_12422,N_12673);
xor U14144 (N_14144,N_13452,N_13880);
nor U14145 (N_14145,N_13102,N_13693);
xnor U14146 (N_14146,N_12211,N_13878);
or U14147 (N_14147,N_12267,N_12011);
nor U14148 (N_14148,N_12452,N_12163);
nor U14149 (N_14149,N_13758,N_12999);
or U14150 (N_14150,N_13612,N_13804);
nand U14151 (N_14151,N_12986,N_12538);
nand U14152 (N_14152,N_13530,N_13778);
nor U14153 (N_14153,N_12182,N_13736);
nor U14154 (N_14154,N_12637,N_12027);
xnor U14155 (N_14155,N_12801,N_12624);
nor U14156 (N_14156,N_13456,N_12859);
and U14157 (N_14157,N_13645,N_13158);
and U14158 (N_14158,N_13996,N_13078);
and U14159 (N_14159,N_13487,N_13480);
nor U14160 (N_14160,N_12881,N_13007);
and U14161 (N_14161,N_12591,N_13715);
and U14162 (N_14162,N_12234,N_12969);
nor U14163 (N_14163,N_13979,N_13302);
or U14164 (N_14164,N_13995,N_12338);
and U14165 (N_14165,N_12951,N_12888);
or U14166 (N_14166,N_13377,N_12689);
nor U14167 (N_14167,N_12925,N_12900);
and U14168 (N_14168,N_12705,N_13410);
and U14169 (N_14169,N_12541,N_13149);
xnor U14170 (N_14170,N_13110,N_12260);
xnor U14171 (N_14171,N_12603,N_13629);
and U14172 (N_14172,N_13871,N_12273);
nand U14173 (N_14173,N_12481,N_13181);
and U14174 (N_14174,N_13192,N_12912);
or U14175 (N_14175,N_13691,N_13161);
or U14176 (N_14176,N_13058,N_12852);
and U14177 (N_14177,N_13277,N_13379);
nor U14178 (N_14178,N_12440,N_12441);
or U14179 (N_14179,N_12492,N_12301);
xor U14180 (N_14180,N_13730,N_12148);
and U14181 (N_14181,N_13724,N_12058);
or U14182 (N_14182,N_12739,N_12686);
and U14183 (N_14183,N_13193,N_12147);
or U14184 (N_14184,N_12363,N_12677);
and U14185 (N_14185,N_12651,N_13572);
nor U14186 (N_14186,N_12070,N_12501);
nand U14187 (N_14187,N_12124,N_13287);
xnor U14188 (N_14188,N_12347,N_12299);
or U14189 (N_14189,N_12169,N_13864);
nor U14190 (N_14190,N_12472,N_13324);
or U14191 (N_14191,N_13106,N_13910);
nor U14192 (N_14192,N_13822,N_12137);
nand U14193 (N_14193,N_13326,N_13601);
xor U14194 (N_14194,N_13415,N_12512);
or U14195 (N_14195,N_13397,N_12922);
and U14196 (N_14196,N_12568,N_13399);
or U14197 (N_14197,N_12855,N_13543);
and U14198 (N_14198,N_12187,N_13190);
nor U14199 (N_14199,N_13582,N_12909);
xnor U14200 (N_14200,N_13363,N_13846);
xnor U14201 (N_14201,N_13615,N_12983);
nand U14202 (N_14202,N_13244,N_13912);
or U14203 (N_14203,N_13567,N_13426);
xnor U14204 (N_14204,N_13117,N_12890);
and U14205 (N_14205,N_12941,N_12703);
and U14206 (N_14206,N_12130,N_12120);
xor U14207 (N_14207,N_13549,N_12893);
nor U14208 (N_14208,N_12596,N_13584);
and U14209 (N_14209,N_13131,N_12397);
and U14210 (N_14210,N_13280,N_13411);
or U14211 (N_14211,N_12954,N_13268);
and U14212 (N_14212,N_12799,N_13129);
and U14213 (N_14213,N_13684,N_12141);
nand U14214 (N_14214,N_13844,N_12110);
or U14215 (N_14215,N_13588,N_13321);
and U14216 (N_14216,N_12362,N_13605);
nand U14217 (N_14217,N_12544,N_13717);
and U14218 (N_14218,N_13359,N_13438);
and U14219 (N_14219,N_12753,N_12431);
xnor U14220 (N_14220,N_12631,N_13726);
and U14221 (N_14221,N_12766,N_13728);
nor U14222 (N_14222,N_13558,N_13356);
or U14223 (N_14223,N_13412,N_13761);
nor U14224 (N_14224,N_12996,N_12804);
nor U14225 (N_14225,N_12085,N_13786);
or U14226 (N_14226,N_12204,N_13056);
and U14227 (N_14227,N_13008,N_12806);
xor U14228 (N_14228,N_12507,N_13096);
nor U14229 (N_14229,N_12574,N_13145);
nand U14230 (N_14230,N_12281,N_12992);
nand U14231 (N_14231,N_13266,N_12641);
or U14232 (N_14232,N_12265,N_12480);
nor U14233 (N_14233,N_13511,N_13066);
nand U14234 (N_14234,N_13330,N_13365);
or U14235 (N_14235,N_13063,N_12336);
or U14236 (N_14236,N_12256,N_13959);
xor U14237 (N_14237,N_13372,N_12836);
xor U14238 (N_14238,N_12691,N_12763);
xor U14239 (N_14239,N_13139,N_13124);
and U14240 (N_14240,N_12479,N_13428);
nor U14241 (N_14241,N_12672,N_13339);
nor U14242 (N_14242,N_13542,N_12343);
and U14243 (N_14243,N_12311,N_12961);
or U14244 (N_14244,N_12847,N_12537);
or U14245 (N_14245,N_12231,N_12597);
and U14246 (N_14246,N_12623,N_12474);
nand U14247 (N_14247,N_12049,N_13742);
xnor U14248 (N_14248,N_13552,N_12412);
or U14249 (N_14249,N_13241,N_13455);
xnor U14250 (N_14250,N_12712,N_12904);
nor U14251 (N_14251,N_13442,N_13757);
nand U14252 (N_14252,N_13566,N_13320);
or U14253 (N_14253,N_13984,N_12613);
nor U14254 (N_14254,N_12860,N_13935);
nor U14255 (N_14255,N_13579,N_13636);
nor U14256 (N_14256,N_12043,N_13528);
xnor U14257 (N_14257,N_12019,N_13205);
nand U14258 (N_14258,N_13134,N_12051);
nand U14259 (N_14259,N_12361,N_13202);
nand U14260 (N_14260,N_13065,N_12706);
or U14261 (N_14261,N_13665,N_13104);
nand U14262 (N_14262,N_13210,N_13422);
and U14263 (N_14263,N_13395,N_13936);
nand U14264 (N_14264,N_13578,N_13830);
xnor U14265 (N_14265,N_13125,N_12482);
and U14266 (N_14266,N_12895,N_12191);
nor U14267 (N_14267,N_12713,N_12497);
nand U14268 (N_14268,N_12443,N_12948);
nor U14269 (N_14269,N_13476,N_12005);
nor U14270 (N_14270,N_13685,N_12500);
nor U14271 (N_14271,N_12867,N_13035);
xnor U14272 (N_14272,N_13877,N_12171);
xor U14273 (N_14273,N_13213,N_12776);
nand U14274 (N_14274,N_13328,N_13540);
and U14275 (N_14275,N_12113,N_12294);
xnor U14276 (N_14276,N_13484,N_13214);
and U14277 (N_14277,N_13470,N_12103);
or U14278 (N_14278,N_13535,N_13188);
or U14279 (N_14279,N_13904,N_12646);
xor U14280 (N_14280,N_12874,N_12149);
or U14281 (N_14281,N_13416,N_12478);
xnor U14282 (N_14282,N_13340,N_13440);
or U14283 (N_14283,N_13220,N_12310);
xor U14284 (N_14284,N_12349,N_12610);
xor U14285 (N_14285,N_13991,N_12838);
xnor U14286 (N_14286,N_13998,N_12876);
and U14287 (N_14287,N_13364,N_13978);
nand U14288 (N_14288,N_12076,N_12812);
nand U14289 (N_14289,N_12707,N_12615);
xor U14290 (N_14290,N_12793,N_12972);
xor U14291 (N_14291,N_12626,N_12393);
nor U14292 (N_14292,N_13044,N_12698);
and U14293 (N_14293,N_12575,N_13186);
xnor U14294 (N_14294,N_13520,N_13595);
and U14295 (N_14295,N_13444,N_12078);
and U14296 (N_14296,N_13183,N_13711);
nor U14297 (N_14297,N_13299,N_13025);
xnor U14298 (N_14298,N_13392,N_13309);
nor U14299 (N_14299,N_13021,N_13817);
and U14300 (N_14300,N_13907,N_12377);
nor U14301 (N_14301,N_13128,N_12292);
xnor U14302 (N_14302,N_12089,N_13654);
xor U14303 (N_14303,N_13648,N_12102);
nor U14304 (N_14304,N_12458,N_13632);
and U14305 (N_14305,N_13700,N_12467);
and U14306 (N_14306,N_13387,N_12298);
xnor U14307 (N_14307,N_12026,N_13704);
nor U14308 (N_14308,N_12400,N_12854);
nand U14309 (N_14309,N_13919,N_12549);
and U14310 (N_14310,N_12731,N_13585);
nand U14311 (N_14311,N_12288,N_12259);
xor U14312 (N_14312,N_12061,N_12185);
xor U14313 (N_14313,N_12505,N_13522);
or U14314 (N_14314,N_12223,N_12272);
and U14315 (N_14315,N_12708,N_12416);
nor U14316 (N_14316,N_13173,N_12977);
nand U14317 (N_14317,N_12355,N_13721);
or U14318 (N_14318,N_13338,N_12025);
or U14319 (N_14319,N_13928,N_12177);
xor U14320 (N_14320,N_12329,N_12570);
nor U14321 (N_14321,N_13023,N_12144);
or U14322 (N_14322,N_12046,N_13093);
and U14323 (N_14323,N_13014,N_12319);
nor U14324 (N_14324,N_13929,N_13551);
nor U14325 (N_14325,N_13831,N_13627);
and U14326 (N_14326,N_12869,N_13800);
and U14327 (N_14327,N_12803,N_12668);
nor U14328 (N_14328,N_13219,N_12002);
xor U14329 (N_14329,N_12030,N_12960);
xnor U14330 (N_14330,N_12495,N_12680);
nor U14331 (N_14331,N_12636,N_12468);
xor U14332 (N_14332,N_12087,N_13234);
and U14333 (N_14333,N_13771,N_12664);
or U14334 (N_14334,N_13490,N_13942);
nand U14335 (N_14335,N_12899,N_13940);
nand U14336 (N_14336,N_12465,N_12134);
or U14337 (N_14337,N_12333,N_12732);
or U14338 (N_14338,N_13111,N_12910);
or U14339 (N_14339,N_12401,N_12945);
nand U14340 (N_14340,N_12216,N_13815);
nand U14341 (N_14341,N_13656,N_12226);
nor U14342 (N_14342,N_13896,N_12145);
nand U14343 (N_14343,N_13238,N_12251);
and U14344 (N_14344,N_13872,N_12679);
and U14345 (N_14345,N_12832,N_13565);
nand U14346 (N_14346,N_12307,N_13630);
or U14347 (N_14347,N_13123,N_13801);
nand U14348 (N_14348,N_13289,N_12433);
and U14349 (N_14349,N_13047,N_13345);
and U14350 (N_14350,N_13853,N_12840);
xor U14351 (N_14351,N_12588,N_12594);
xnor U14352 (N_14352,N_13517,N_12725);
nor U14353 (N_14353,N_12324,N_12075);
or U14354 (N_14354,N_13980,N_13180);
xnor U14355 (N_14355,N_12252,N_12487);
xnor U14356 (N_14356,N_12638,N_12749);
nand U14357 (N_14357,N_13406,N_12627);
xor U14358 (N_14358,N_12862,N_12493);
nand U14359 (N_14359,N_12166,N_13855);
and U14360 (N_14360,N_12554,N_12815);
nor U14361 (N_14361,N_13500,N_13033);
nand U14362 (N_14362,N_13425,N_13918);
nor U14363 (N_14363,N_12295,N_12451);
or U14364 (N_14364,N_13137,N_12740);
and U14365 (N_14365,N_13571,N_12991);
nor U14366 (N_14366,N_12576,N_12444);
and U14367 (N_14367,N_12657,N_13466);
and U14368 (N_14368,N_12682,N_13114);
xor U14369 (N_14369,N_12022,N_13529);
and U14370 (N_14370,N_13596,N_12990);
and U14371 (N_14371,N_12536,N_12477);
and U14372 (N_14372,N_13006,N_13638);
xor U14373 (N_14373,N_13159,N_13401);
nand U14374 (N_14374,N_13300,N_12916);
or U14375 (N_14375,N_12426,N_13203);
nand U14376 (N_14376,N_12716,N_13559);
nor U14377 (N_14377,N_12460,N_12116);
nand U14378 (N_14378,N_13646,N_12632);
nand U14379 (N_14379,N_13127,N_12304);
nor U14380 (N_14380,N_12800,N_13780);
and U14381 (N_14381,N_12222,N_13677);
nor U14382 (N_14382,N_12697,N_12580);
and U14383 (N_14383,N_13155,N_13669);
or U14384 (N_14384,N_13754,N_12366);
xor U14385 (N_14385,N_12129,N_13344);
xor U14386 (N_14386,N_12957,N_12567);
and U14387 (N_14387,N_12097,N_12318);
xnor U14388 (N_14388,N_12358,N_12432);
or U14389 (N_14389,N_12618,N_12198);
xnor U14390 (N_14390,N_13336,N_13095);
nor U14391 (N_14391,N_12499,N_13436);
xor U14392 (N_14392,N_13624,N_12475);
xnor U14393 (N_14393,N_12028,N_13739);
nand U14394 (N_14394,N_13897,N_12870);
and U14395 (N_14395,N_13826,N_12783);
nor U14396 (N_14396,N_12315,N_12271);
xnor U14397 (N_14397,N_12640,N_13510);
nor U14398 (N_14398,N_13660,N_13212);
and U14399 (N_14399,N_13286,N_12313);
xnor U14400 (N_14400,N_13865,N_13649);
and U14401 (N_14401,N_13337,N_12528);
and U14402 (N_14402,N_12425,N_12778);
xor U14403 (N_14403,N_13652,N_12781);
or U14404 (N_14404,N_13390,N_13174);
and U14405 (N_14405,N_13230,N_13163);
nand U14406 (N_14406,N_13441,N_12872);
and U14407 (N_14407,N_12647,N_12785);
nor U14408 (N_14408,N_13080,N_13501);
nor U14409 (N_14409,N_13544,N_12398);
nand U14410 (N_14410,N_13489,N_13729);
and U14411 (N_14411,N_12072,N_13577);
nand U14412 (N_14412,N_12524,N_13950);
nand U14413 (N_14413,N_12843,N_12949);
nor U14414 (N_14414,N_12335,N_13697);
nand U14415 (N_14415,N_13040,N_13026);
and U14416 (N_14416,N_13409,N_12887);
nor U14417 (N_14417,N_12192,N_13388);
and U14418 (N_14418,N_12200,N_13661);
nand U14419 (N_14419,N_12723,N_13211);
xnor U14420 (N_14420,N_13148,N_13386);
nand U14421 (N_14421,N_13598,N_13019);
and U14422 (N_14422,N_12735,N_13308);
xnor U14423 (N_14423,N_13564,N_13206);
nand U14424 (N_14424,N_13414,N_12614);
nand U14425 (N_14425,N_13472,N_12715);
nor U14426 (N_14426,N_12109,N_12833);
and U14427 (N_14427,N_13852,N_12820);
nor U14428 (N_14428,N_13315,N_12040);
nor U14429 (N_14429,N_13043,N_13905);
or U14430 (N_14430,N_12082,N_13814);
nand U14431 (N_14431,N_13130,N_13097);
or U14432 (N_14432,N_12428,N_12818);
nand U14433 (N_14433,N_13143,N_12935);
and U14434 (N_14434,N_13886,N_13863);
xnor U14435 (N_14435,N_12898,N_12207);
and U14436 (N_14436,N_12967,N_12540);
xor U14437 (N_14437,N_13461,N_13067);
or U14438 (N_14438,N_12209,N_12819);
or U14439 (N_14439,N_12920,N_12880);
and U14440 (N_14440,N_13545,N_13705);
or U14441 (N_14441,N_12543,N_13591);
nor U14442 (N_14442,N_13256,N_13841);
xnor U14443 (N_14443,N_12365,N_12188);
nor U14444 (N_14444,N_13505,N_13177);
xor U14445 (N_14445,N_13295,N_13851);
nor U14446 (N_14446,N_12578,N_13182);
nor U14447 (N_14447,N_12054,N_13682);
xor U14448 (N_14448,N_12106,N_12584);
nand U14449 (N_14449,N_12710,N_13431);
xnor U14450 (N_14450,N_13274,N_12514);
nor U14451 (N_14451,N_13171,N_12558);
xnor U14452 (N_14452,N_12736,N_12622);
nor U14453 (N_14453,N_13790,N_12371);
and U14454 (N_14454,N_13062,N_13663);
nor U14455 (N_14455,N_12321,N_13447);
xor U14456 (N_14456,N_12257,N_13921);
nand U14457 (N_14457,N_13609,N_13460);
or U14458 (N_14458,N_13267,N_13874);
and U14459 (N_14459,N_12828,N_13176);
nand U14460 (N_14460,N_13623,N_12404);
and U14461 (N_14461,N_12572,N_13657);
or U14462 (N_14462,N_12434,N_13394);
nand U14463 (N_14463,N_12417,N_13385);
nor U14464 (N_14464,N_12563,N_12720);
or U14465 (N_14465,N_12306,N_12345);
nand U14466 (N_14466,N_13361,N_12456);
nand U14467 (N_14467,N_13418,N_13334);
nor U14468 (N_14468,N_12611,N_12268);
and U14469 (N_14469,N_12408,N_12418);
nor U14470 (N_14470,N_12665,N_13429);
nor U14471 (N_14471,N_12504,N_13022);
and U14472 (N_14472,N_12060,N_13223);
or U14473 (N_14473,N_13348,N_13765);
xnor U14474 (N_14474,N_12938,N_13404);
nor U14475 (N_14475,N_13568,N_13553);
and U14476 (N_14476,N_13304,N_12856);
nand U14477 (N_14477,N_13818,N_13900);
or U14478 (N_14478,N_13029,N_13502);
xnor U14479 (N_14479,N_12787,N_12118);
xnor U14480 (N_14480,N_13686,N_12024);
and U14481 (N_14481,N_12602,N_13306);
or U14482 (N_14482,N_12915,N_13094);
and U14483 (N_14483,N_12905,N_12521);
xor U14484 (N_14484,N_12559,N_12660);
nor U14485 (N_14485,N_13323,N_12903);
nor U14486 (N_14486,N_13424,N_13034);
nor U14487 (N_14487,N_12926,N_13459);
or U14488 (N_14488,N_13191,N_12745);
or U14489 (N_14489,N_13498,N_12530);
xnor U14490 (N_14490,N_12968,N_13602);
xor U14491 (N_14491,N_12156,N_12656);
nor U14492 (N_14492,N_12891,N_13891);
nor U14493 (N_14493,N_12018,N_12190);
and U14494 (N_14494,N_13811,N_12639);
nor U14495 (N_14495,N_13109,N_13059);
nand U14496 (N_14496,N_13621,N_12527);
nor U14497 (N_14497,N_13945,N_12159);
xor U14498 (N_14498,N_12368,N_12795);
and U14499 (N_14499,N_12410,N_13606);
and U14500 (N_14500,N_13257,N_13888);
nor U14501 (N_14501,N_12411,N_12535);
and U14502 (N_14502,N_12976,N_12817);
xor U14503 (N_14503,N_12842,N_13407);
or U14504 (N_14504,N_12045,N_12092);
nand U14505 (N_14505,N_13278,N_12327);
nor U14506 (N_14506,N_13254,N_12896);
and U14507 (N_14507,N_13548,N_12067);
nor U14508 (N_14508,N_12844,N_12386);
nand U14509 (N_14509,N_12050,N_12143);
and U14510 (N_14510,N_12369,N_12714);
nor U14511 (N_14511,N_13074,N_13408);
or U14512 (N_14512,N_13987,N_12606);
nor U14513 (N_14513,N_13294,N_12387);
and U14514 (N_14514,N_12409,N_12966);
or U14515 (N_14515,N_13495,N_13037);
nor U14516 (N_14516,N_12937,N_12733);
xor U14517 (N_14517,N_12033,N_13994);
and U14518 (N_14518,N_13643,N_13091);
and U14519 (N_14519,N_13710,N_12532);
and U14520 (N_14520,N_13136,N_12308);
nor U14521 (N_14521,N_13293,N_13531);
nor U14522 (N_14522,N_12764,N_12219);
nor U14523 (N_14523,N_12189,N_12681);
or U14524 (N_14524,N_13297,N_12217);
or U14525 (N_14525,N_13948,N_12429);
xnor U14526 (N_14526,N_13162,N_12760);
nor U14527 (N_14527,N_13264,N_13737);
nand U14528 (N_14528,N_13892,N_13722);
or U14529 (N_14529,N_13982,N_13450);
xor U14530 (N_14530,N_12167,N_13869);
or U14531 (N_14531,N_13030,N_12035);
or U14532 (N_14532,N_13678,N_12342);
and U14533 (N_14533,N_12608,N_12747);
or U14534 (N_14534,N_13366,N_13357);
or U14535 (N_14535,N_13154,N_12297);
nor U14536 (N_14536,N_12748,N_12091);
nand U14537 (N_14537,N_12805,N_13611);
and U14538 (N_14538,N_13335,N_13708);
and U14539 (N_14539,N_13885,N_12997);
xnor U14540 (N_14540,N_13702,N_13467);
and U14541 (N_14541,N_13823,N_12670);
xnor U14542 (N_14542,N_13172,N_12503);
nand U14543 (N_14543,N_13369,N_12621);
xnor U14544 (N_14544,N_13454,N_12663);
or U14545 (N_14545,N_12201,N_12678);
nand U14546 (N_14546,N_12062,N_12285);
nand U14547 (N_14547,N_13347,N_13647);
nand U14548 (N_14548,N_12918,N_12269);
xnor U14549 (N_14549,N_12824,N_12438);
and U14550 (N_14550,N_12121,N_13860);
nand U14551 (N_14551,N_12322,N_13322);
nand U14552 (N_14552,N_12822,N_13857);
or U14553 (N_14553,N_13288,N_13068);
nand U14554 (N_14554,N_12305,N_13462);
xnor U14555 (N_14555,N_12215,N_12625);
and U14556 (N_14556,N_12248,N_13626);
nor U14557 (N_14557,N_12245,N_12119);
nor U14558 (N_14558,N_12696,N_13313);
xnor U14559 (N_14559,N_13593,N_12186);
or U14560 (N_14560,N_13748,N_13133);
xor U14561 (N_14561,N_12518,N_12556);
nor U14562 (N_14562,N_12790,N_13046);
or U14563 (N_14563,N_13990,N_13525);
and U14564 (N_14564,N_13538,N_13894);
nand U14565 (N_14565,N_13402,N_12865);
nor U14566 (N_14566,N_13516,N_12879);
or U14567 (N_14567,N_12032,N_12055);
and U14568 (N_14568,N_12439,N_13439);
nand U14569 (N_14569,N_12894,N_13583);
or U14570 (N_14570,N_12218,N_13911);
or U14571 (N_14571,N_13261,N_12980);
xnor U14572 (N_14572,N_13196,N_12984);
or U14573 (N_14573,N_13002,N_13135);
nor U14574 (N_14574,N_12436,N_13473);
nand U14575 (N_14575,N_13752,N_13445);
xor U14576 (N_14576,N_13974,N_12970);
and U14577 (N_14577,N_12300,N_13534);
or U14578 (N_14578,N_13833,N_13464);
xnor U14579 (N_14579,N_12826,N_12921);
nand U14580 (N_14580,N_13914,N_13635);
or U14581 (N_14581,N_12229,N_13837);
nor U14582 (N_14582,N_13150,N_12173);
and U14583 (N_14583,N_13793,N_13255);
nor U14584 (N_14584,N_13011,N_13437);
nor U14585 (N_14585,N_12729,N_12571);
nor U14586 (N_14586,N_12088,N_12389);
nand U14587 (N_14587,N_13231,N_12642);
nand U14588 (N_14588,N_12210,N_12153);
nand U14589 (N_14589,N_12671,N_13233);
nand U14590 (N_14590,N_13903,N_13506);
or U14591 (N_14591,N_13497,N_12476);
nor U14592 (N_14592,N_13152,N_12709);
or U14593 (N_14593,N_12415,N_13856);
xor U14594 (N_14594,N_12593,N_12565);
xnor U14595 (N_14595,N_12768,N_13164);
and U14596 (N_14596,N_13967,N_12789);
nor U14597 (N_14597,N_12170,N_12582);
and U14598 (N_14598,N_12901,N_13156);
xor U14599 (N_14599,N_13533,N_13053);
and U14600 (N_14600,N_12573,N_12373);
nand U14601 (N_14601,N_12255,N_13245);
nor U14602 (N_14602,N_12551,N_13250);
xor U14603 (N_14603,N_12762,N_13756);
or U14604 (N_14604,N_13235,N_12965);
nand U14605 (N_14605,N_13938,N_12086);
or U14606 (N_14606,N_13920,N_13718);
nor U14607 (N_14607,N_12437,N_13229);
nor U14608 (N_14608,N_13240,N_13695);
nand U14609 (N_14609,N_12490,N_13194);
nand U14610 (N_14610,N_12312,N_13712);
nor U14611 (N_14611,N_12367,N_12374);
or U14612 (N_14612,N_13039,N_13933);
nor U14613 (N_14613,N_13491,N_13719);
nand U14614 (N_14614,N_12531,N_13042);
and U14615 (N_14615,N_13070,N_13430);
and U14616 (N_14616,N_12380,N_13992);
nor U14617 (N_14617,N_12927,N_13953);
nor U14618 (N_14618,N_13689,N_13977);
nor U14619 (N_14619,N_12466,N_13118);
xor U14620 (N_14620,N_13204,N_12564);
xnor U14621 (N_14621,N_12464,N_12289);
and U14622 (N_14622,N_13465,N_13318);
or U14623 (N_14623,N_13696,N_13969);
xor U14624 (N_14624,N_12542,N_12172);
and U14625 (N_14625,N_13380,N_12309);
or U14626 (N_14626,N_12270,N_13064);
xor U14627 (N_14627,N_12816,N_12693);
nand U14628 (N_14628,N_13075,N_12010);
nand U14629 (N_14629,N_12792,N_12929);
xnor U14630 (N_14630,N_12772,N_13924);
nand U14631 (N_14631,N_13083,N_12017);
nor U14632 (N_14632,N_13733,N_13482);
nor U14633 (N_14633,N_12099,N_13488);
and U14634 (N_14634,N_13962,N_13253);
or U14635 (N_14635,N_12254,N_12101);
nor U14636 (N_14636,N_12423,N_12446);
nand U14637 (N_14637,N_12105,N_13716);
nand U14638 (N_14638,N_12633,N_12934);
nand U14639 (N_14639,N_13675,N_12947);
nand U14640 (N_14640,N_12958,N_12094);
nand U14641 (N_14641,N_13389,N_12376);
xnor U14642 (N_14642,N_12917,N_13051);
nand U14643 (N_14643,N_13839,N_13753);
nor U14644 (N_14644,N_13838,N_12830);
or U14645 (N_14645,N_13769,N_12093);
nor U14646 (N_14646,N_13667,N_12320);
and U14647 (N_14647,N_13796,N_13569);
xnor U14648 (N_14648,N_13055,N_12545);
xor U14649 (N_14649,N_12246,N_12012);
or U14650 (N_14650,N_13847,N_12034);
nand U14651 (N_14651,N_12635,N_12738);
or U14652 (N_14652,N_12115,N_12123);
and U14653 (N_14653,N_13504,N_12240);
nand U14654 (N_14654,N_12837,N_13536);
nand U14655 (N_14655,N_12291,N_13273);
nand U14656 (N_14656,N_12726,N_12029);
and U14657 (N_14657,N_13659,N_13750);
and U14658 (N_14658,N_12846,N_13845);
xor U14659 (N_14659,N_12346,N_12827);
nor U14660 (N_14660,N_13247,N_13072);
xor U14661 (N_14661,N_12071,N_13971);
and U14662 (N_14662,N_13802,N_13513);
nor U14663 (N_14663,N_13311,N_12517);
nor U14664 (N_14664,N_12734,N_13650);
nor U14665 (N_14665,N_12858,N_13727);
nand U14666 (N_14666,N_12821,N_13009);
nand U14667 (N_14667,N_13616,N_12353);
and U14668 (N_14668,N_13666,N_12688);
xnor U14669 (N_14669,N_12009,N_12453);
nor U14670 (N_14670,N_12004,N_12491);
nand U14671 (N_14671,N_12600,N_12759);
and U14672 (N_14672,N_13787,N_13483);
or U14673 (N_14673,N_13561,N_12548);
or U14674 (N_14674,N_13908,N_13681);
and U14675 (N_14675,N_13824,N_12339);
xnor U14676 (N_14676,N_12508,N_13242);
nor U14677 (N_14677,N_12550,N_12114);
nor U14678 (N_14678,N_12212,N_13875);
and U14679 (N_14679,N_12777,N_13307);
nor U14680 (N_14680,N_12784,N_12841);
and U14681 (N_14681,N_13282,N_13884);
nor U14682 (N_14682,N_13332,N_13570);
nand U14683 (N_14683,N_12811,N_13057);
and U14684 (N_14684,N_13089,N_12155);
nor U14685 (N_14685,N_13597,N_12328);
xor U14686 (N_14686,N_12224,N_12649);
or U14687 (N_14687,N_13507,N_13600);
or U14688 (N_14688,N_12981,N_12807);
nand U14689 (N_14689,N_13079,N_12403);
xor U14690 (N_14690,N_12612,N_12150);
and U14691 (N_14691,N_13798,N_12973);
or U14692 (N_14692,N_13384,N_13343);
and U14693 (N_14693,N_13810,N_13449);
and U14694 (N_14694,N_13720,N_12348);
or U14695 (N_14695,N_13836,N_13653);
xor U14696 (N_14696,N_13768,N_13862);
or U14697 (N_14697,N_13419,N_12221);
xor U14698 (N_14698,N_12752,N_13272);
nor U14699 (N_14699,N_12194,N_12430);
nand U14700 (N_14700,N_12146,N_13222);
nor U14701 (N_14701,N_12902,N_13433);
xor U14702 (N_14702,N_12195,N_12683);
xnor U14703 (N_14703,N_12379,N_13956);
and U14704 (N_14704,N_13090,N_13509);
xnor U14705 (N_14705,N_13981,N_13732);
xor U14706 (N_14706,N_12442,N_12165);
and U14707 (N_14707,N_12258,N_13012);
xnor U14708 (N_14708,N_13119,N_13382);
nand U14709 (N_14709,N_13285,N_13707);
nor U14710 (N_14710,N_13519,N_13749);
nor U14711 (N_14711,N_12038,N_12360);
nand U14712 (N_14712,N_13599,N_13975);
or U14713 (N_14713,N_12331,N_13706);
or U14714 (N_14714,N_13641,N_13922);
xor U14715 (N_14715,N_13867,N_13251);
xnor U14716 (N_14716,N_13842,N_13292);
or U14717 (N_14717,N_12998,N_13524);
xor U14718 (N_14718,N_13794,N_13496);
xor U14719 (N_14719,N_13747,N_13122);
xnor U14720 (N_14720,N_12340,N_13403);
xor U14721 (N_14721,N_12077,N_13291);
xnor U14722 (N_14722,N_12962,N_12364);
xor U14723 (N_14723,N_12420,N_13575);
or U14724 (N_14724,N_12863,N_12845);
or U14725 (N_14725,N_13360,N_13614);
and U14726 (N_14726,N_13917,N_13038);
or U14727 (N_14727,N_12486,N_13644);
nand U14728 (N_14728,N_13899,N_12620);
xor U14729 (N_14729,N_12769,N_12341);
or U14730 (N_14730,N_13503,N_13642);
nor U14731 (N_14731,N_13349,N_13054);
nor U14732 (N_14732,N_12939,N_12601);
xnor U14733 (N_14733,N_13633,N_13115);
nor U14734 (N_14734,N_12864,N_12914);
xnor U14735 (N_14735,N_13608,N_13527);
and U14736 (N_14736,N_13116,N_12523);
xnor U14737 (N_14737,N_13265,N_12157);
xnor U14738 (N_14738,N_13485,N_12694);
and U14739 (N_14739,N_13099,N_12154);
or U14740 (N_14740,N_12196,N_13592);
and U14741 (N_14741,N_12036,N_13200);
nor U14742 (N_14742,N_13809,N_13887);
xnor U14743 (N_14743,N_13806,N_12213);
nand U14744 (N_14744,N_13168,N_12080);
nor U14745 (N_14745,N_13069,N_12522);
nand U14746 (N_14746,N_13049,N_13759);
and U14747 (N_14747,N_12199,N_12151);
xnor U14748 (N_14748,N_12502,N_13698);
nor U14749 (N_14749,N_12122,N_13679);
xnor U14750 (N_14750,N_12850,N_13284);
and U14751 (N_14751,N_12687,N_13353);
nand U14752 (N_14752,N_12955,N_12402);
or U14753 (N_14753,N_12546,N_12053);
nor U14754 (N_14754,N_13989,N_12419);
nor U14755 (N_14755,N_13586,N_12303);
xor U14756 (N_14756,N_13619,N_13671);
and U14757 (N_14757,N_12228,N_12765);
or U14758 (N_14758,N_12174,N_13160);
nor U14759 (N_14759,N_12930,N_12421);
nand U14760 (N_14760,N_13555,N_13175);
and U14761 (N_14761,N_13848,N_12690);
nor U14762 (N_14762,N_13521,N_13248);
nor U14763 (N_14763,N_12607,N_12994);
and U14764 (N_14764,N_12354,N_12737);
or U14765 (N_14765,N_13783,N_12232);
nor U14766 (N_14766,N_12037,N_12184);
and U14767 (N_14767,N_12164,N_12515);
nand U14768 (N_14768,N_13631,N_12359);
or U14769 (N_14769,N_12770,N_13523);
and U14770 (N_14770,N_13236,N_13258);
nand U14771 (N_14771,N_12111,N_13170);
xnor U14772 (N_14772,N_12654,N_13547);
or U14773 (N_14773,N_13499,N_13071);
or U14774 (N_14774,N_12277,N_13107);
and U14775 (N_14775,N_12589,N_13041);
nor U14776 (N_14776,N_12178,N_13714);
or U14777 (N_14777,N_13479,N_13208);
or U14778 (N_14778,N_13821,N_13988);
nor U14779 (N_14779,N_12461,N_12519);
nor U14780 (N_14780,N_12168,N_12214);
or U14781 (N_14781,N_12382,N_12700);
and U14782 (N_14782,N_12244,N_12971);
and U14783 (N_14783,N_13249,N_13672);
nor U14784 (N_14784,N_12238,N_12250);
xor U14785 (N_14785,N_13795,N_13563);
nand U14786 (N_14786,N_13937,N_12662);
xor U14787 (N_14787,N_12616,N_13883);
or U14788 (N_14788,N_13594,N_12406);
xor U14789 (N_14789,N_13081,N_12924);
or U14790 (N_14790,N_13902,N_12853);
nor U14791 (N_14791,N_13791,N_13882);
or U14792 (N_14792,N_12813,N_13458);
nand U14793 (N_14793,N_13077,N_12509);
nand U14794 (N_14794,N_13997,N_13774);
xor U14795 (N_14795,N_13189,N_12450);
and U14796 (N_14796,N_12352,N_12193);
nand U14797 (N_14797,N_13405,N_12488);
or U14798 (N_14798,N_13964,N_12652);
or U14799 (N_14799,N_12928,N_12396);
nand U14800 (N_14800,N_13471,N_13179);
and U14801 (N_14801,N_13468,N_12831);
or U14802 (N_14802,N_13751,N_13772);
xor U14803 (N_14803,N_12350,N_13889);
or U14804 (N_14804,N_13239,N_12263);
or U14805 (N_14805,N_13965,N_13004);
or U14806 (N_14806,N_12230,N_13017);
nand U14807 (N_14807,N_12617,N_12181);
nor U14808 (N_14808,N_13243,N_12197);
and U14809 (N_14809,N_12378,N_12797);
nand U14810 (N_14810,N_12042,N_12933);
nand U14811 (N_14811,N_13723,N_12774);
xor U14812 (N_14812,N_13932,N_13589);
nand U14813 (N_14813,N_12133,N_13986);
or U14814 (N_14814,N_13581,N_13620);
or U14815 (N_14815,N_13178,N_12128);
xor U14816 (N_14816,N_13371,N_12445);
or U14817 (N_14817,N_12598,N_13784);
nand U14818 (N_14818,N_13827,N_13789);
nor U14819 (N_14819,N_12278,N_12592);
nand U14820 (N_14820,N_13603,N_13303);
or U14821 (N_14821,N_13105,N_12630);
nand U14822 (N_14822,N_12241,N_13061);
and U14823 (N_14823,N_12877,N_13890);
and U14824 (N_14824,N_13909,N_13275);
or U14825 (N_14825,N_13699,N_12069);
or U14826 (N_14826,N_13259,N_12266);
nand U14827 (N_14827,N_13376,N_12014);
nand U14828 (N_14828,N_13331,N_12595);
xnor U14829 (N_14829,N_12562,N_13797);
and U14830 (N_14830,N_12395,N_13317);
and U14831 (N_14831,N_12758,N_13100);
xnor U14832 (N_14832,N_12510,N_13617);
xor U14833 (N_14833,N_13840,N_13451);
nand U14834 (N_14834,N_13341,N_13201);
or U14835 (N_14835,N_13060,N_13618);
or U14836 (N_14836,N_13983,N_12483);
xnor U14837 (N_14837,N_12455,N_13374);
or U14838 (N_14838,N_13944,N_13263);
xor U14839 (N_14839,N_12435,N_13092);
nand U14840 (N_14840,N_13915,N_12287);
xor U14841 (N_14841,N_12599,N_13805);
xnor U14842 (N_14842,N_13868,N_13731);
or U14843 (N_14843,N_13688,N_12773);
or U14844 (N_14844,N_12237,N_12096);
xnor U14845 (N_14845,N_13260,N_12851);
and U14846 (N_14846,N_13082,N_13381);
xor U14847 (N_14847,N_13165,N_12586);
and U14848 (N_14848,N_12946,N_12560);
nor U14849 (N_14849,N_12083,N_12985);
nand U14850 (N_14850,N_13861,N_12950);
xnor U14851 (N_14851,N_12886,N_13664);
nand U14852 (N_14852,N_12066,N_13779);
and U14853 (N_14853,N_12427,N_13141);
nor U14854 (N_14854,N_12334,N_13140);
nand U14855 (N_14855,N_13808,N_12619);
nand U14856 (N_14856,N_13673,N_13333);
nand U14857 (N_14857,N_12283,N_12264);
nand U14858 (N_14858,N_13269,N_12581);
nand U14859 (N_14859,N_13658,N_13613);
nand U14860 (N_14860,N_12057,N_13690);
nand U14861 (N_14861,N_13541,N_13926);
nor U14862 (N_14862,N_12868,N_13427);
and U14863 (N_14863,N_13590,N_13367);
and U14864 (N_14864,N_13434,N_13199);
nand U14865 (N_14865,N_12064,N_12883);
xor U14866 (N_14866,N_13741,N_13226);
or U14867 (N_14867,N_12007,N_12605);
or U14868 (N_14868,N_13512,N_12882);
xor U14869 (N_14869,N_12577,N_12020);
nand U14870 (N_14870,N_13157,N_12457);
or U14871 (N_14871,N_13925,N_13084);
and U14872 (N_14872,N_13271,N_13113);
and U14873 (N_14873,N_12227,N_12754);
or U14874 (N_14874,N_13849,N_13001);
nand U14875 (N_14875,N_12317,N_13352);
and U14876 (N_14876,N_13692,N_12666);
or U14877 (N_14877,N_13760,N_12885);
and U14878 (N_14878,N_13866,N_13913);
and U14879 (N_14879,N_12484,N_12534);
nand U14880 (N_14880,N_13785,N_13216);
and U14881 (N_14881,N_12073,N_13812);
nor U14882 (N_14882,N_12809,N_12405);
nand U14883 (N_14883,N_13580,N_13290);
nor U14884 (N_14884,N_13943,N_12063);
nor U14885 (N_14885,N_13370,N_13195);
and U14886 (N_14886,N_13952,N_12730);
and U14887 (N_14887,N_12407,N_13985);
xnor U14888 (N_14888,N_12579,N_12658);
or U14889 (N_14889,N_12135,N_12332);
nand U14890 (N_14890,N_12953,N_12861);
xor U14891 (N_14891,N_13972,N_12810);
or U14892 (N_14892,N_13215,N_12701);
xor U14893 (N_14893,N_12496,N_12659);
nor U14894 (N_14894,N_13329,N_13052);
nand U14895 (N_14895,N_13481,N_12108);
nand U14896 (N_14896,N_13738,N_12107);
and U14897 (N_14897,N_13788,N_13217);
or U14898 (N_14898,N_12286,N_12650);
xor U14899 (N_14899,N_13396,N_13701);
nand U14900 (N_14900,N_12392,N_12117);
xnor U14901 (N_14901,N_12494,N_13147);
xor U14902 (N_14902,N_13574,N_12065);
xnor U14903 (N_14903,N_13674,N_13167);
and U14904 (N_14904,N_12202,N_12702);
xnor U14905 (N_14905,N_12337,N_12583);
nand U14906 (N_14906,N_12391,N_12100);
nand U14907 (N_14907,N_12280,N_12127);
and U14908 (N_14908,N_13050,N_12684);
and U14909 (N_14909,N_12236,N_12520);
and U14910 (N_14910,N_12931,N_12975);
nand U14911 (N_14911,N_13151,N_12750);
and U14912 (N_14912,N_12987,N_12000);
nand U14913 (N_14913,N_12344,N_12674);
or U14914 (N_14914,N_12786,N_12767);
nand U14915 (N_14915,N_13088,N_12136);
xor U14916 (N_14916,N_12943,N_12048);
nor U14917 (N_14917,N_13651,N_12995);
xor U14918 (N_14918,N_13015,N_12695);
nand U14919 (N_14919,N_12284,N_12242);
nand U14920 (N_14920,N_13227,N_12721);
xnor U14921 (N_14921,N_12140,N_12239);
nor U14922 (N_14922,N_12293,N_13166);
xor U14923 (N_14923,N_13098,N_12796);
nor U14924 (N_14924,N_13237,N_13120);
or U14925 (N_14925,N_13443,N_13400);
nor U14926 (N_14926,N_12942,N_13628);
xnor U14927 (N_14927,N_12802,N_12323);
nand U14928 (N_14928,N_12643,N_13354);
and U14929 (N_14929,N_13457,N_12383);
and U14930 (N_14930,N_13954,N_12047);
or U14931 (N_14931,N_12090,N_12529);
and U14932 (N_14932,N_13493,N_12126);
or U14933 (N_14933,N_13755,N_13477);
or U14934 (N_14934,N_12944,N_12176);
xnor U14935 (N_14935,N_13024,N_13005);
or U14936 (N_14936,N_12158,N_13546);
and U14937 (N_14937,N_13246,N_13683);
nor U14938 (N_14938,N_13835,N_13557);
xor U14939 (N_14939,N_13625,N_13906);
nand U14940 (N_14940,N_13391,N_12751);
or U14941 (N_14941,N_13453,N_12798);
nor U14942 (N_14942,N_12068,N_12533);
nor U14943 (N_14943,N_12023,N_13073);
xnor U14944 (N_14944,N_13879,N_12756);
or U14945 (N_14945,N_12448,N_13828);
or U14946 (N_14946,N_12316,N_13668);
nor U14947 (N_14947,N_12506,N_12516);
or U14948 (N_14948,N_13398,N_12139);
xor U14949 (N_14949,N_12016,N_13368);
or U14950 (N_14950,N_12388,N_12235);
and U14951 (N_14951,N_12471,N_13930);
or U14952 (N_14952,N_12871,N_12835);
nand U14953 (N_14953,N_13854,N_12276);
xor U14954 (N_14954,N_12008,N_12413);
nand U14955 (N_14955,N_13803,N_12356);
xor U14956 (N_14956,N_12526,N_13232);
xnor U14957 (N_14957,N_13949,N_12175);
nor U14958 (N_14958,N_12485,N_13276);
or U14959 (N_14959,N_13138,N_12814);
and U14960 (N_14960,N_12183,N_12989);
and U14961 (N_14961,N_13469,N_12959);
xnor U14962 (N_14962,N_12808,N_12553);
xor U14963 (N_14963,N_13526,N_13218);
and U14964 (N_14964,N_12857,N_13446);
nand U14965 (N_14965,N_13744,N_12685);
nor U14966 (N_14966,N_12724,N_12667);
nor U14967 (N_14967,N_13486,N_13680);
nor U14968 (N_14968,N_12095,N_12138);
xnor U14969 (N_14969,N_13085,N_12779);
nand U14970 (N_14970,N_12162,N_12669);
nor U14971 (N_14971,N_13895,N_13676);
and U14972 (N_14972,N_13958,N_13834);
xnor U14973 (N_14973,N_12742,N_12282);
nand U14974 (N_14974,N_12913,N_13947);
xor U14975 (N_14975,N_13478,N_12585);
nand U14976 (N_14976,N_12473,N_12220);
nor U14977 (N_14977,N_12160,N_13003);
or U14978 (N_14978,N_13032,N_13556);
nand U14979 (N_14979,N_12275,N_12728);
nor U14980 (N_14980,N_12372,N_12161);
and U14981 (N_14981,N_13662,N_12661);
and U14982 (N_14982,N_12757,N_13898);
xnor U14983 (N_14983,N_13016,N_13934);
xnor U14984 (N_14984,N_13562,N_13770);
nand U14985 (N_14985,N_13939,N_13637);
and U14986 (N_14986,N_13153,N_13420);
or U14987 (N_14987,N_13413,N_13020);
xnor U14988 (N_14988,N_12719,N_12180);
or U14989 (N_14989,N_13725,N_12059);
nor U14990 (N_14990,N_12907,N_13607);
and U14991 (N_14991,N_13816,N_12566);
xnor U14992 (N_14992,N_13475,N_13999);
and U14993 (N_14993,N_13184,N_12557);
or U14994 (N_14994,N_13126,N_12609);
nand U14995 (N_14995,N_13108,N_12152);
nand U14996 (N_14996,N_13146,N_13514);
or U14997 (N_14997,N_12878,N_12590);
and U14998 (N_14998,N_13850,N_13112);
nor U14999 (N_14999,N_13782,N_12897);
nand U15000 (N_15000,N_13352,N_12182);
xor U15001 (N_15001,N_13305,N_12500);
nor U15002 (N_15002,N_13928,N_12147);
nand U15003 (N_15003,N_12115,N_13178);
or U15004 (N_15004,N_12044,N_12621);
or U15005 (N_15005,N_13212,N_13311);
xnor U15006 (N_15006,N_12864,N_13113);
nand U15007 (N_15007,N_13982,N_12930);
xor U15008 (N_15008,N_12618,N_12356);
xnor U15009 (N_15009,N_12357,N_12858);
or U15010 (N_15010,N_13805,N_12453);
or U15011 (N_15011,N_13350,N_12539);
or U15012 (N_15012,N_12573,N_13241);
nand U15013 (N_15013,N_13576,N_13457);
xnor U15014 (N_15014,N_13160,N_13121);
xnor U15015 (N_15015,N_12211,N_13056);
or U15016 (N_15016,N_13106,N_13838);
xor U15017 (N_15017,N_13285,N_13367);
nand U15018 (N_15018,N_13878,N_13620);
xnor U15019 (N_15019,N_13918,N_13835);
and U15020 (N_15020,N_13310,N_13140);
nand U15021 (N_15021,N_13985,N_12876);
or U15022 (N_15022,N_13485,N_12801);
and U15023 (N_15023,N_12427,N_13992);
nand U15024 (N_15024,N_12850,N_12764);
or U15025 (N_15025,N_13470,N_13769);
or U15026 (N_15026,N_12062,N_13055);
xnor U15027 (N_15027,N_12881,N_13399);
nor U15028 (N_15028,N_12669,N_13142);
and U15029 (N_15029,N_13773,N_12104);
nand U15030 (N_15030,N_13586,N_13798);
or U15031 (N_15031,N_12735,N_13388);
nor U15032 (N_15032,N_12684,N_12797);
or U15033 (N_15033,N_13221,N_13298);
nand U15034 (N_15034,N_12533,N_13627);
or U15035 (N_15035,N_13290,N_13442);
xor U15036 (N_15036,N_13832,N_13760);
or U15037 (N_15037,N_12392,N_13835);
nor U15038 (N_15038,N_13330,N_13238);
xnor U15039 (N_15039,N_12555,N_13993);
nor U15040 (N_15040,N_12327,N_12921);
nand U15041 (N_15041,N_13941,N_12252);
or U15042 (N_15042,N_12450,N_12302);
or U15043 (N_15043,N_12065,N_13336);
xnor U15044 (N_15044,N_12388,N_12253);
and U15045 (N_15045,N_12348,N_12272);
and U15046 (N_15046,N_13988,N_13230);
nor U15047 (N_15047,N_13710,N_12902);
nor U15048 (N_15048,N_13963,N_13408);
or U15049 (N_15049,N_13623,N_13947);
nand U15050 (N_15050,N_12417,N_13396);
nor U15051 (N_15051,N_13908,N_13497);
or U15052 (N_15052,N_12969,N_13376);
xor U15053 (N_15053,N_13483,N_13591);
or U15054 (N_15054,N_13492,N_13771);
xnor U15055 (N_15055,N_13343,N_12553);
xnor U15056 (N_15056,N_12412,N_13627);
and U15057 (N_15057,N_12238,N_12542);
nor U15058 (N_15058,N_13246,N_13324);
xnor U15059 (N_15059,N_13140,N_12711);
xnor U15060 (N_15060,N_12531,N_13374);
nor U15061 (N_15061,N_12786,N_12229);
and U15062 (N_15062,N_12340,N_12587);
nor U15063 (N_15063,N_12065,N_12924);
xor U15064 (N_15064,N_12247,N_12522);
nand U15065 (N_15065,N_12606,N_12768);
nor U15066 (N_15066,N_13403,N_12058);
or U15067 (N_15067,N_12676,N_12891);
xnor U15068 (N_15068,N_12106,N_13013);
nor U15069 (N_15069,N_13439,N_13409);
nand U15070 (N_15070,N_13665,N_13819);
xor U15071 (N_15071,N_13147,N_12961);
nor U15072 (N_15072,N_12185,N_13976);
or U15073 (N_15073,N_13655,N_13183);
or U15074 (N_15074,N_12238,N_13479);
nand U15075 (N_15075,N_12847,N_13713);
nor U15076 (N_15076,N_13337,N_12614);
xor U15077 (N_15077,N_12837,N_13599);
xnor U15078 (N_15078,N_13227,N_12934);
nand U15079 (N_15079,N_12754,N_12164);
xor U15080 (N_15080,N_12419,N_12631);
nor U15081 (N_15081,N_13464,N_13946);
xor U15082 (N_15082,N_13094,N_13592);
and U15083 (N_15083,N_12516,N_13076);
nand U15084 (N_15084,N_12302,N_12934);
xor U15085 (N_15085,N_13703,N_12450);
or U15086 (N_15086,N_12980,N_13242);
and U15087 (N_15087,N_12245,N_12005);
nor U15088 (N_15088,N_12948,N_12320);
or U15089 (N_15089,N_12484,N_12578);
nor U15090 (N_15090,N_12766,N_13614);
or U15091 (N_15091,N_12420,N_13410);
or U15092 (N_15092,N_12241,N_12756);
xnor U15093 (N_15093,N_12524,N_12500);
xnor U15094 (N_15094,N_13397,N_13470);
nor U15095 (N_15095,N_12130,N_13907);
xor U15096 (N_15096,N_13574,N_13530);
nor U15097 (N_15097,N_12664,N_12874);
nor U15098 (N_15098,N_12938,N_13134);
and U15099 (N_15099,N_13955,N_13344);
and U15100 (N_15100,N_12265,N_13267);
xor U15101 (N_15101,N_13054,N_12867);
and U15102 (N_15102,N_13910,N_13705);
or U15103 (N_15103,N_12718,N_13768);
xnor U15104 (N_15104,N_12718,N_13052);
nor U15105 (N_15105,N_13073,N_13257);
nor U15106 (N_15106,N_13507,N_12635);
or U15107 (N_15107,N_12015,N_13657);
nand U15108 (N_15108,N_12195,N_13973);
and U15109 (N_15109,N_12703,N_12831);
nand U15110 (N_15110,N_12686,N_13640);
and U15111 (N_15111,N_12017,N_13597);
nor U15112 (N_15112,N_13776,N_12328);
nand U15113 (N_15113,N_12975,N_12348);
nor U15114 (N_15114,N_13363,N_12394);
nor U15115 (N_15115,N_12727,N_12557);
and U15116 (N_15116,N_13659,N_12280);
nor U15117 (N_15117,N_12672,N_13723);
and U15118 (N_15118,N_12502,N_12907);
xor U15119 (N_15119,N_12559,N_13003);
nand U15120 (N_15120,N_12263,N_13469);
xnor U15121 (N_15121,N_13465,N_12693);
or U15122 (N_15122,N_12187,N_13552);
xnor U15123 (N_15123,N_13852,N_13020);
nand U15124 (N_15124,N_12613,N_12305);
or U15125 (N_15125,N_12628,N_12833);
or U15126 (N_15126,N_12806,N_12425);
or U15127 (N_15127,N_13393,N_12273);
nand U15128 (N_15128,N_12072,N_13209);
nor U15129 (N_15129,N_13040,N_12960);
or U15130 (N_15130,N_12354,N_13060);
and U15131 (N_15131,N_12653,N_13166);
nand U15132 (N_15132,N_13670,N_13167);
nand U15133 (N_15133,N_12172,N_13341);
nand U15134 (N_15134,N_12790,N_12556);
and U15135 (N_15135,N_12287,N_13524);
nand U15136 (N_15136,N_12779,N_13152);
nand U15137 (N_15137,N_12356,N_12979);
nand U15138 (N_15138,N_13453,N_12773);
nor U15139 (N_15139,N_12606,N_12835);
or U15140 (N_15140,N_12043,N_13693);
or U15141 (N_15141,N_12306,N_12735);
or U15142 (N_15142,N_13978,N_13073);
and U15143 (N_15143,N_13473,N_13945);
nand U15144 (N_15144,N_12770,N_13812);
and U15145 (N_15145,N_13510,N_13883);
xor U15146 (N_15146,N_12536,N_13621);
xnor U15147 (N_15147,N_13080,N_13066);
xor U15148 (N_15148,N_12002,N_12578);
nor U15149 (N_15149,N_12523,N_12922);
nand U15150 (N_15150,N_13761,N_12761);
nand U15151 (N_15151,N_13408,N_12302);
nor U15152 (N_15152,N_13470,N_13392);
nand U15153 (N_15153,N_13650,N_13070);
nor U15154 (N_15154,N_13801,N_12163);
and U15155 (N_15155,N_12352,N_13921);
nor U15156 (N_15156,N_13272,N_12412);
nor U15157 (N_15157,N_12518,N_12109);
or U15158 (N_15158,N_13996,N_13165);
nor U15159 (N_15159,N_12037,N_13075);
nor U15160 (N_15160,N_13766,N_12735);
xnor U15161 (N_15161,N_13522,N_12367);
nand U15162 (N_15162,N_13284,N_12977);
nand U15163 (N_15163,N_12329,N_12114);
and U15164 (N_15164,N_13638,N_12961);
nor U15165 (N_15165,N_13858,N_12827);
and U15166 (N_15166,N_12002,N_12219);
nand U15167 (N_15167,N_12476,N_13924);
xor U15168 (N_15168,N_13235,N_13517);
nand U15169 (N_15169,N_13911,N_12674);
and U15170 (N_15170,N_13167,N_13036);
nor U15171 (N_15171,N_13171,N_12837);
or U15172 (N_15172,N_12272,N_12778);
nor U15173 (N_15173,N_12971,N_12488);
nand U15174 (N_15174,N_12833,N_12565);
and U15175 (N_15175,N_13753,N_13312);
nand U15176 (N_15176,N_13230,N_13094);
nor U15177 (N_15177,N_12041,N_12481);
xor U15178 (N_15178,N_13762,N_13226);
or U15179 (N_15179,N_12729,N_13395);
nor U15180 (N_15180,N_13189,N_12867);
nand U15181 (N_15181,N_12264,N_13472);
and U15182 (N_15182,N_13597,N_13842);
xor U15183 (N_15183,N_13177,N_12268);
xnor U15184 (N_15184,N_13889,N_13865);
nor U15185 (N_15185,N_12735,N_13220);
or U15186 (N_15186,N_13882,N_12821);
nand U15187 (N_15187,N_13523,N_12314);
or U15188 (N_15188,N_13395,N_13695);
nand U15189 (N_15189,N_12219,N_13864);
nand U15190 (N_15190,N_12743,N_13610);
xor U15191 (N_15191,N_12008,N_13180);
and U15192 (N_15192,N_13645,N_12542);
nand U15193 (N_15193,N_12898,N_12769);
and U15194 (N_15194,N_13416,N_13578);
or U15195 (N_15195,N_13001,N_13521);
or U15196 (N_15196,N_12415,N_13827);
nand U15197 (N_15197,N_12463,N_13136);
nand U15198 (N_15198,N_13207,N_12194);
or U15199 (N_15199,N_12110,N_13035);
nor U15200 (N_15200,N_12648,N_12921);
or U15201 (N_15201,N_12987,N_13154);
nand U15202 (N_15202,N_12940,N_13812);
xnor U15203 (N_15203,N_13244,N_12075);
and U15204 (N_15204,N_13743,N_13233);
and U15205 (N_15205,N_13081,N_12585);
or U15206 (N_15206,N_13203,N_13161);
or U15207 (N_15207,N_12805,N_12076);
xor U15208 (N_15208,N_12540,N_13196);
xnor U15209 (N_15209,N_13203,N_13603);
nor U15210 (N_15210,N_13231,N_13119);
and U15211 (N_15211,N_13401,N_13179);
and U15212 (N_15212,N_13790,N_12187);
nor U15213 (N_15213,N_13320,N_12198);
xnor U15214 (N_15214,N_12076,N_13724);
and U15215 (N_15215,N_12391,N_13077);
and U15216 (N_15216,N_13070,N_12278);
or U15217 (N_15217,N_12729,N_13464);
or U15218 (N_15218,N_13548,N_12095);
or U15219 (N_15219,N_13692,N_13165);
or U15220 (N_15220,N_12858,N_12578);
xnor U15221 (N_15221,N_13945,N_13276);
nand U15222 (N_15222,N_12463,N_13313);
and U15223 (N_15223,N_13294,N_13819);
nand U15224 (N_15224,N_13385,N_12881);
nand U15225 (N_15225,N_12516,N_13211);
nor U15226 (N_15226,N_12240,N_13759);
or U15227 (N_15227,N_12720,N_13348);
or U15228 (N_15228,N_13932,N_13285);
and U15229 (N_15229,N_13205,N_12359);
nor U15230 (N_15230,N_12803,N_12042);
or U15231 (N_15231,N_13802,N_12672);
and U15232 (N_15232,N_13763,N_13413);
nor U15233 (N_15233,N_13360,N_12849);
and U15234 (N_15234,N_12019,N_13181);
nand U15235 (N_15235,N_13630,N_12551);
nand U15236 (N_15236,N_13561,N_12843);
nor U15237 (N_15237,N_13004,N_12389);
or U15238 (N_15238,N_12420,N_13747);
nand U15239 (N_15239,N_13558,N_12681);
nor U15240 (N_15240,N_12028,N_12437);
and U15241 (N_15241,N_13381,N_13261);
or U15242 (N_15242,N_12162,N_13019);
nor U15243 (N_15243,N_12567,N_12832);
and U15244 (N_15244,N_12733,N_12666);
nand U15245 (N_15245,N_13669,N_13861);
and U15246 (N_15246,N_12970,N_12062);
nor U15247 (N_15247,N_13972,N_13718);
nand U15248 (N_15248,N_13765,N_12324);
xnor U15249 (N_15249,N_13585,N_13411);
and U15250 (N_15250,N_13235,N_13275);
nand U15251 (N_15251,N_12531,N_12820);
nor U15252 (N_15252,N_13726,N_13047);
nor U15253 (N_15253,N_13061,N_13109);
nor U15254 (N_15254,N_12724,N_13373);
and U15255 (N_15255,N_12574,N_12034);
nor U15256 (N_15256,N_13678,N_13095);
and U15257 (N_15257,N_13506,N_13563);
nor U15258 (N_15258,N_12469,N_12415);
nor U15259 (N_15259,N_13912,N_12183);
nor U15260 (N_15260,N_12125,N_12208);
or U15261 (N_15261,N_13792,N_13965);
nor U15262 (N_15262,N_13636,N_13115);
xnor U15263 (N_15263,N_12431,N_12749);
and U15264 (N_15264,N_13155,N_12029);
xnor U15265 (N_15265,N_13957,N_13970);
or U15266 (N_15266,N_12099,N_12094);
nor U15267 (N_15267,N_12481,N_13628);
xor U15268 (N_15268,N_12780,N_13915);
xnor U15269 (N_15269,N_12340,N_13063);
nor U15270 (N_15270,N_13112,N_12608);
nand U15271 (N_15271,N_13779,N_12830);
and U15272 (N_15272,N_13865,N_12480);
nand U15273 (N_15273,N_12987,N_13307);
and U15274 (N_15274,N_13602,N_12219);
xnor U15275 (N_15275,N_13217,N_12715);
xor U15276 (N_15276,N_13392,N_12198);
and U15277 (N_15277,N_12611,N_12982);
nand U15278 (N_15278,N_12544,N_12913);
nand U15279 (N_15279,N_13955,N_12551);
or U15280 (N_15280,N_13594,N_12058);
and U15281 (N_15281,N_13440,N_12918);
nor U15282 (N_15282,N_13512,N_12981);
or U15283 (N_15283,N_13695,N_13767);
nor U15284 (N_15284,N_12891,N_12224);
nor U15285 (N_15285,N_13001,N_12315);
nand U15286 (N_15286,N_13032,N_13898);
nand U15287 (N_15287,N_13677,N_12630);
nor U15288 (N_15288,N_12830,N_13933);
xnor U15289 (N_15289,N_13870,N_13676);
nand U15290 (N_15290,N_13605,N_12575);
xnor U15291 (N_15291,N_13068,N_12909);
nand U15292 (N_15292,N_13459,N_12900);
xnor U15293 (N_15293,N_13245,N_12485);
or U15294 (N_15294,N_12682,N_13345);
nand U15295 (N_15295,N_12590,N_12337);
nor U15296 (N_15296,N_12880,N_13804);
xnor U15297 (N_15297,N_12605,N_12915);
nor U15298 (N_15298,N_13301,N_12481);
nand U15299 (N_15299,N_13896,N_13997);
nor U15300 (N_15300,N_13932,N_13594);
xor U15301 (N_15301,N_12195,N_13571);
and U15302 (N_15302,N_13981,N_12344);
nand U15303 (N_15303,N_13246,N_12205);
and U15304 (N_15304,N_13625,N_12012);
nor U15305 (N_15305,N_13814,N_12024);
xor U15306 (N_15306,N_13366,N_12584);
nand U15307 (N_15307,N_12063,N_13971);
and U15308 (N_15308,N_12309,N_12067);
and U15309 (N_15309,N_12411,N_12632);
and U15310 (N_15310,N_13584,N_13422);
nand U15311 (N_15311,N_12997,N_12081);
and U15312 (N_15312,N_12240,N_13545);
and U15313 (N_15313,N_12373,N_13534);
nor U15314 (N_15314,N_13103,N_12584);
nor U15315 (N_15315,N_13757,N_12196);
or U15316 (N_15316,N_12751,N_12335);
or U15317 (N_15317,N_12050,N_12428);
and U15318 (N_15318,N_13716,N_12874);
nor U15319 (N_15319,N_13601,N_12260);
nand U15320 (N_15320,N_12137,N_12309);
or U15321 (N_15321,N_12594,N_13340);
and U15322 (N_15322,N_13295,N_12891);
and U15323 (N_15323,N_13887,N_12698);
nor U15324 (N_15324,N_13228,N_13812);
xnor U15325 (N_15325,N_12032,N_13525);
or U15326 (N_15326,N_12137,N_13371);
and U15327 (N_15327,N_12003,N_12439);
nand U15328 (N_15328,N_13026,N_12188);
nand U15329 (N_15329,N_13791,N_12814);
and U15330 (N_15330,N_13332,N_13935);
nor U15331 (N_15331,N_12764,N_13283);
nand U15332 (N_15332,N_13872,N_12972);
xor U15333 (N_15333,N_12215,N_12405);
xnor U15334 (N_15334,N_12813,N_12166);
and U15335 (N_15335,N_12553,N_13269);
xor U15336 (N_15336,N_12443,N_13681);
and U15337 (N_15337,N_13352,N_13960);
nand U15338 (N_15338,N_12926,N_13131);
xnor U15339 (N_15339,N_12199,N_12534);
nand U15340 (N_15340,N_12620,N_12126);
xor U15341 (N_15341,N_12437,N_13405);
or U15342 (N_15342,N_12355,N_13665);
nand U15343 (N_15343,N_13201,N_12283);
and U15344 (N_15344,N_13696,N_13666);
xor U15345 (N_15345,N_13305,N_12865);
and U15346 (N_15346,N_13765,N_13777);
nor U15347 (N_15347,N_13034,N_13269);
and U15348 (N_15348,N_13987,N_12975);
or U15349 (N_15349,N_13349,N_13139);
nand U15350 (N_15350,N_12052,N_12605);
nand U15351 (N_15351,N_13714,N_13378);
nand U15352 (N_15352,N_13731,N_13325);
and U15353 (N_15353,N_12920,N_13468);
nor U15354 (N_15354,N_12501,N_13105);
and U15355 (N_15355,N_13223,N_12293);
or U15356 (N_15356,N_13228,N_13959);
and U15357 (N_15357,N_13154,N_13930);
xnor U15358 (N_15358,N_13493,N_12912);
xor U15359 (N_15359,N_13249,N_12453);
nand U15360 (N_15360,N_13226,N_13562);
and U15361 (N_15361,N_13796,N_13877);
and U15362 (N_15362,N_13128,N_13475);
or U15363 (N_15363,N_13769,N_12695);
xnor U15364 (N_15364,N_12556,N_12485);
xnor U15365 (N_15365,N_12776,N_13090);
or U15366 (N_15366,N_13674,N_13864);
and U15367 (N_15367,N_13455,N_12380);
and U15368 (N_15368,N_12451,N_13981);
xor U15369 (N_15369,N_13075,N_13807);
nor U15370 (N_15370,N_12811,N_13175);
and U15371 (N_15371,N_13614,N_13162);
nand U15372 (N_15372,N_13743,N_13037);
nor U15373 (N_15373,N_12810,N_12360);
xor U15374 (N_15374,N_13400,N_13435);
xnor U15375 (N_15375,N_12139,N_13254);
or U15376 (N_15376,N_13603,N_12092);
and U15377 (N_15377,N_12740,N_13034);
nor U15378 (N_15378,N_12513,N_12815);
or U15379 (N_15379,N_12469,N_12377);
nand U15380 (N_15380,N_13261,N_13333);
nor U15381 (N_15381,N_13755,N_12332);
xor U15382 (N_15382,N_12225,N_13493);
or U15383 (N_15383,N_12845,N_13904);
xor U15384 (N_15384,N_13206,N_12752);
and U15385 (N_15385,N_12618,N_13113);
and U15386 (N_15386,N_12508,N_12165);
nand U15387 (N_15387,N_13805,N_13207);
xor U15388 (N_15388,N_12116,N_12125);
and U15389 (N_15389,N_13159,N_12970);
xor U15390 (N_15390,N_12034,N_12057);
nand U15391 (N_15391,N_13588,N_12583);
nor U15392 (N_15392,N_13734,N_13541);
nor U15393 (N_15393,N_12881,N_12575);
nand U15394 (N_15394,N_12120,N_13374);
xor U15395 (N_15395,N_13427,N_13337);
and U15396 (N_15396,N_13459,N_13849);
or U15397 (N_15397,N_13702,N_12227);
nand U15398 (N_15398,N_13019,N_13393);
and U15399 (N_15399,N_13882,N_13227);
nor U15400 (N_15400,N_13753,N_13386);
nor U15401 (N_15401,N_12727,N_12171);
nand U15402 (N_15402,N_13606,N_13476);
and U15403 (N_15403,N_12659,N_13880);
xnor U15404 (N_15404,N_12546,N_13454);
nor U15405 (N_15405,N_12224,N_13913);
xnor U15406 (N_15406,N_13941,N_12369);
nor U15407 (N_15407,N_12626,N_13877);
or U15408 (N_15408,N_13698,N_13323);
nor U15409 (N_15409,N_13861,N_12453);
xnor U15410 (N_15410,N_13223,N_12416);
nand U15411 (N_15411,N_13599,N_13292);
xor U15412 (N_15412,N_12817,N_13198);
xnor U15413 (N_15413,N_13417,N_12266);
nand U15414 (N_15414,N_12554,N_12650);
nor U15415 (N_15415,N_12080,N_13954);
and U15416 (N_15416,N_13331,N_12891);
xnor U15417 (N_15417,N_12535,N_12249);
and U15418 (N_15418,N_12808,N_12195);
and U15419 (N_15419,N_13611,N_13846);
xnor U15420 (N_15420,N_13357,N_13049);
and U15421 (N_15421,N_13161,N_12190);
nor U15422 (N_15422,N_13369,N_12305);
xor U15423 (N_15423,N_13941,N_13913);
or U15424 (N_15424,N_12133,N_12381);
xnor U15425 (N_15425,N_12034,N_13939);
nor U15426 (N_15426,N_13845,N_12370);
and U15427 (N_15427,N_12665,N_12479);
nand U15428 (N_15428,N_12294,N_12020);
nand U15429 (N_15429,N_13065,N_12448);
nand U15430 (N_15430,N_12455,N_12018);
nor U15431 (N_15431,N_13217,N_12449);
nand U15432 (N_15432,N_12423,N_13605);
or U15433 (N_15433,N_13393,N_13060);
nor U15434 (N_15434,N_12029,N_13325);
or U15435 (N_15435,N_12087,N_12273);
or U15436 (N_15436,N_12919,N_12535);
and U15437 (N_15437,N_12698,N_13480);
or U15438 (N_15438,N_13299,N_12928);
nand U15439 (N_15439,N_13090,N_13704);
nand U15440 (N_15440,N_13972,N_12636);
and U15441 (N_15441,N_12858,N_12344);
or U15442 (N_15442,N_13513,N_13481);
nor U15443 (N_15443,N_12841,N_12676);
xor U15444 (N_15444,N_13538,N_13630);
nor U15445 (N_15445,N_12461,N_13531);
nor U15446 (N_15446,N_13010,N_12916);
nor U15447 (N_15447,N_13852,N_12742);
nand U15448 (N_15448,N_12759,N_13486);
and U15449 (N_15449,N_13863,N_12117);
and U15450 (N_15450,N_12460,N_12718);
nor U15451 (N_15451,N_12767,N_12426);
xnor U15452 (N_15452,N_12523,N_12131);
and U15453 (N_15453,N_13757,N_12726);
nor U15454 (N_15454,N_13490,N_12237);
and U15455 (N_15455,N_12877,N_12854);
nor U15456 (N_15456,N_12862,N_12187);
or U15457 (N_15457,N_13985,N_12993);
nor U15458 (N_15458,N_13412,N_13636);
xnor U15459 (N_15459,N_13014,N_12170);
or U15460 (N_15460,N_13761,N_12956);
or U15461 (N_15461,N_13609,N_13522);
or U15462 (N_15462,N_12714,N_13433);
nor U15463 (N_15463,N_13458,N_13790);
nand U15464 (N_15464,N_12826,N_13135);
or U15465 (N_15465,N_13431,N_13123);
nor U15466 (N_15466,N_12819,N_13669);
nor U15467 (N_15467,N_13238,N_13590);
xor U15468 (N_15468,N_13016,N_13852);
or U15469 (N_15469,N_12450,N_12191);
and U15470 (N_15470,N_13234,N_13500);
and U15471 (N_15471,N_12616,N_12217);
nand U15472 (N_15472,N_12743,N_13179);
or U15473 (N_15473,N_13482,N_13261);
nand U15474 (N_15474,N_13390,N_12947);
xor U15475 (N_15475,N_13161,N_12139);
or U15476 (N_15476,N_13817,N_13094);
nand U15477 (N_15477,N_13420,N_13643);
or U15478 (N_15478,N_12399,N_12635);
or U15479 (N_15479,N_12321,N_12043);
nor U15480 (N_15480,N_12442,N_13469);
and U15481 (N_15481,N_12291,N_13764);
nor U15482 (N_15482,N_13090,N_12321);
or U15483 (N_15483,N_12304,N_13610);
nand U15484 (N_15484,N_13458,N_13198);
or U15485 (N_15485,N_13806,N_13873);
nor U15486 (N_15486,N_12326,N_13227);
nor U15487 (N_15487,N_13644,N_13746);
and U15488 (N_15488,N_12245,N_12214);
nor U15489 (N_15489,N_13378,N_12242);
xor U15490 (N_15490,N_12816,N_12438);
and U15491 (N_15491,N_13741,N_12955);
nand U15492 (N_15492,N_12427,N_13205);
or U15493 (N_15493,N_13617,N_13161);
nand U15494 (N_15494,N_13355,N_12977);
xor U15495 (N_15495,N_13823,N_12340);
xnor U15496 (N_15496,N_13435,N_13653);
nand U15497 (N_15497,N_12337,N_13526);
nand U15498 (N_15498,N_13163,N_13527);
nand U15499 (N_15499,N_12115,N_13865);
and U15500 (N_15500,N_12702,N_12435);
xor U15501 (N_15501,N_13903,N_12565);
xor U15502 (N_15502,N_13258,N_13397);
and U15503 (N_15503,N_12255,N_12066);
or U15504 (N_15504,N_13481,N_13740);
and U15505 (N_15505,N_12134,N_12779);
and U15506 (N_15506,N_12334,N_12277);
nor U15507 (N_15507,N_12000,N_12271);
or U15508 (N_15508,N_13656,N_13193);
nor U15509 (N_15509,N_12417,N_13093);
nor U15510 (N_15510,N_13350,N_13704);
or U15511 (N_15511,N_13565,N_13064);
and U15512 (N_15512,N_13365,N_13539);
xnor U15513 (N_15513,N_12799,N_12106);
xor U15514 (N_15514,N_12655,N_12566);
xnor U15515 (N_15515,N_13533,N_13842);
and U15516 (N_15516,N_12910,N_12848);
xnor U15517 (N_15517,N_12525,N_12502);
xor U15518 (N_15518,N_12778,N_13402);
or U15519 (N_15519,N_13055,N_12615);
or U15520 (N_15520,N_12203,N_13831);
and U15521 (N_15521,N_13126,N_13498);
xnor U15522 (N_15522,N_12094,N_12548);
nand U15523 (N_15523,N_12940,N_12699);
or U15524 (N_15524,N_13024,N_13577);
nand U15525 (N_15525,N_13611,N_13055);
and U15526 (N_15526,N_12768,N_12230);
or U15527 (N_15527,N_13352,N_12690);
nor U15528 (N_15528,N_12071,N_13025);
nor U15529 (N_15529,N_13296,N_13981);
nor U15530 (N_15530,N_12046,N_13033);
and U15531 (N_15531,N_13916,N_13917);
nand U15532 (N_15532,N_13043,N_12054);
or U15533 (N_15533,N_13214,N_13181);
nand U15534 (N_15534,N_12247,N_12947);
nor U15535 (N_15535,N_13870,N_13401);
or U15536 (N_15536,N_12819,N_12133);
and U15537 (N_15537,N_13328,N_12256);
nor U15538 (N_15538,N_12547,N_12022);
or U15539 (N_15539,N_13671,N_13008);
nor U15540 (N_15540,N_12357,N_12733);
or U15541 (N_15541,N_13185,N_12499);
or U15542 (N_15542,N_13271,N_13819);
nand U15543 (N_15543,N_12876,N_13699);
xor U15544 (N_15544,N_12421,N_13389);
and U15545 (N_15545,N_13402,N_12924);
or U15546 (N_15546,N_13414,N_12965);
xor U15547 (N_15547,N_12938,N_13680);
nand U15548 (N_15548,N_13660,N_13382);
nand U15549 (N_15549,N_12503,N_13608);
nand U15550 (N_15550,N_12467,N_13195);
or U15551 (N_15551,N_13945,N_13347);
and U15552 (N_15552,N_12540,N_12929);
xor U15553 (N_15553,N_12477,N_12867);
and U15554 (N_15554,N_13678,N_13518);
nor U15555 (N_15555,N_13768,N_13764);
xor U15556 (N_15556,N_13492,N_12866);
xor U15557 (N_15557,N_13465,N_13663);
xor U15558 (N_15558,N_12238,N_13469);
and U15559 (N_15559,N_12246,N_12975);
nor U15560 (N_15560,N_12627,N_12978);
nor U15561 (N_15561,N_13563,N_13252);
nor U15562 (N_15562,N_13623,N_13860);
or U15563 (N_15563,N_12340,N_12703);
nand U15564 (N_15564,N_13815,N_12904);
nand U15565 (N_15565,N_12172,N_13154);
or U15566 (N_15566,N_12729,N_13276);
nand U15567 (N_15567,N_13389,N_13657);
and U15568 (N_15568,N_12285,N_13483);
and U15569 (N_15569,N_13974,N_12550);
xor U15570 (N_15570,N_13196,N_12663);
nor U15571 (N_15571,N_12253,N_12613);
xnor U15572 (N_15572,N_12565,N_13668);
xor U15573 (N_15573,N_13328,N_13336);
and U15574 (N_15574,N_13523,N_12869);
and U15575 (N_15575,N_13516,N_12517);
nor U15576 (N_15576,N_13662,N_13104);
nand U15577 (N_15577,N_12611,N_13934);
nor U15578 (N_15578,N_12261,N_12411);
nand U15579 (N_15579,N_12577,N_12713);
nor U15580 (N_15580,N_13780,N_13711);
or U15581 (N_15581,N_13427,N_13714);
xor U15582 (N_15582,N_13208,N_12808);
nand U15583 (N_15583,N_12574,N_13750);
xor U15584 (N_15584,N_13143,N_12171);
or U15585 (N_15585,N_13071,N_12651);
or U15586 (N_15586,N_13317,N_12615);
nand U15587 (N_15587,N_13239,N_13928);
and U15588 (N_15588,N_12779,N_12675);
nand U15589 (N_15589,N_13842,N_12654);
nand U15590 (N_15590,N_12348,N_12130);
and U15591 (N_15591,N_12442,N_12709);
and U15592 (N_15592,N_12251,N_12743);
and U15593 (N_15593,N_13840,N_13428);
nor U15594 (N_15594,N_12575,N_13347);
and U15595 (N_15595,N_13826,N_13222);
or U15596 (N_15596,N_13858,N_12117);
or U15597 (N_15597,N_12767,N_13503);
nor U15598 (N_15598,N_12396,N_12708);
nand U15599 (N_15599,N_13578,N_12938);
xor U15600 (N_15600,N_13994,N_13251);
nand U15601 (N_15601,N_12549,N_13888);
nand U15602 (N_15602,N_12335,N_12911);
xnor U15603 (N_15603,N_12582,N_12276);
or U15604 (N_15604,N_13798,N_13829);
nand U15605 (N_15605,N_12583,N_13052);
and U15606 (N_15606,N_12859,N_13382);
nor U15607 (N_15607,N_13239,N_13461);
nor U15608 (N_15608,N_13334,N_13582);
xnor U15609 (N_15609,N_13074,N_12637);
nand U15610 (N_15610,N_12152,N_13001);
nand U15611 (N_15611,N_12582,N_13314);
xnor U15612 (N_15612,N_12064,N_12502);
xor U15613 (N_15613,N_13798,N_13312);
xnor U15614 (N_15614,N_13261,N_12417);
nand U15615 (N_15615,N_13598,N_13917);
or U15616 (N_15616,N_13499,N_13437);
and U15617 (N_15617,N_12333,N_12284);
nand U15618 (N_15618,N_12408,N_13102);
xor U15619 (N_15619,N_12863,N_12402);
and U15620 (N_15620,N_13787,N_12368);
nor U15621 (N_15621,N_12127,N_13105);
and U15622 (N_15622,N_13828,N_13858);
or U15623 (N_15623,N_12702,N_13642);
nor U15624 (N_15624,N_13541,N_13071);
and U15625 (N_15625,N_12727,N_12683);
nand U15626 (N_15626,N_12645,N_12630);
nand U15627 (N_15627,N_13513,N_13673);
xnor U15628 (N_15628,N_13655,N_12797);
xnor U15629 (N_15629,N_13440,N_12859);
nand U15630 (N_15630,N_12107,N_13299);
and U15631 (N_15631,N_13921,N_13018);
or U15632 (N_15632,N_13009,N_13167);
nor U15633 (N_15633,N_12894,N_13585);
xor U15634 (N_15634,N_13932,N_13491);
or U15635 (N_15635,N_13922,N_13137);
and U15636 (N_15636,N_12173,N_12678);
nor U15637 (N_15637,N_12997,N_13602);
xnor U15638 (N_15638,N_12806,N_13469);
and U15639 (N_15639,N_12655,N_13542);
or U15640 (N_15640,N_13042,N_12535);
nand U15641 (N_15641,N_13137,N_13721);
nand U15642 (N_15642,N_13798,N_13597);
nor U15643 (N_15643,N_13022,N_13072);
xnor U15644 (N_15644,N_12290,N_12112);
nor U15645 (N_15645,N_12273,N_13657);
xor U15646 (N_15646,N_12887,N_13506);
or U15647 (N_15647,N_13297,N_13344);
nand U15648 (N_15648,N_13607,N_12438);
nand U15649 (N_15649,N_12583,N_13180);
or U15650 (N_15650,N_12936,N_13549);
and U15651 (N_15651,N_12675,N_12493);
nand U15652 (N_15652,N_12280,N_13019);
nand U15653 (N_15653,N_13149,N_12260);
nor U15654 (N_15654,N_13017,N_12699);
xor U15655 (N_15655,N_12464,N_12255);
nor U15656 (N_15656,N_13760,N_13663);
nand U15657 (N_15657,N_13080,N_12274);
nor U15658 (N_15658,N_12772,N_12018);
and U15659 (N_15659,N_13239,N_13269);
xor U15660 (N_15660,N_13697,N_13073);
xor U15661 (N_15661,N_13731,N_12792);
and U15662 (N_15662,N_12471,N_12558);
and U15663 (N_15663,N_12490,N_12464);
and U15664 (N_15664,N_12092,N_13063);
nand U15665 (N_15665,N_13626,N_12332);
nand U15666 (N_15666,N_12086,N_12577);
nand U15667 (N_15667,N_12113,N_13947);
or U15668 (N_15668,N_13528,N_12217);
or U15669 (N_15669,N_12033,N_12247);
nand U15670 (N_15670,N_12629,N_13555);
and U15671 (N_15671,N_12021,N_13581);
or U15672 (N_15672,N_12787,N_13581);
nand U15673 (N_15673,N_12370,N_12588);
xor U15674 (N_15674,N_12000,N_12966);
and U15675 (N_15675,N_13696,N_13306);
nor U15676 (N_15676,N_13912,N_12229);
xnor U15677 (N_15677,N_13572,N_12995);
and U15678 (N_15678,N_13110,N_12954);
nor U15679 (N_15679,N_12516,N_12253);
nand U15680 (N_15680,N_12207,N_12333);
nor U15681 (N_15681,N_12147,N_12985);
and U15682 (N_15682,N_13776,N_12878);
or U15683 (N_15683,N_13972,N_13595);
and U15684 (N_15684,N_13256,N_13974);
or U15685 (N_15685,N_13036,N_12386);
xor U15686 (N_15686,N_12342,N_12920);
or U15687 (N_15687,N_12164,N_12705);
and U15688 (N_15688,N_13449,N_13978);
xor U15689 (N_15689,N_12819,N_13875);
nor U15690 (N_15690,N_13405,N_12560);
nor U15691 (N_15691,N_13908,N_12111);
nor U15692 (N_15692,N_13521,N_12983);
nor U15693 (N_15693,N_12678,N_13039);
nand U15694 (N_15694,N_12709,N_13531);
nor U15695 (N_15695,N_12247,N_13147);
nand U15696 (N_15696,N_13314,N_12772);
and U15697 (N_15697,N_13085,N_12463);
nor U15698 (N_15698,N_12255,N_12456);
and U15699 (N_15699,N_12682,N_13111);
xnor U15700 (N_15700,N_13138,N_12784);
nor U15701 (N_15701,N_12693,N_13507);
xnor U15702 (N_15702,N_13343,N_12956);
nor U15703 (N_15703,N_12818,N_12462);
nand U15704 (N_15704,N_12635,N_12508);
or U15705 (N_15705,N_13145,N_12768);
nand U15706 (N_15706,N_12588,N_13132);
nand U15707 (N_15707,N_12726,N_13527);
nand U15708 (N_15708,N_13715,N_13489);
and U15709 (N_15709,N_13791,N_12011);
and U15710 (N_15710,N_12483,N_13499);
nand U15711 (N_15711,N_12491,N_13855);
nor U15712 (N_15712,N_13956,N_13524);
or U15713 (N_15713,N_12733,N_12600);
or U15714 (N_15714,N_12798,N_12097);
or U15715 (N_15715,N_12592,N_12821);
xor U15716 (N_15716,N_12405,N_13006);
xnor U15717 (N_15717,N_12094,N_12043);
nand U15718 (N_15718,N_12245,N_12921);
or U15719 (N_15719,N_13070,N_13876);
nor U15720 (N_15720,N_13210,N_12997);
and U15721 (N_15721,N_12346,N_12989);
xor U15722 (N_15722,N_12957,N_12854);
or U15723 (N_15723,N_12959,N_12616);
or U15724 (N_15724,N_12117,N_13081);
nor U15725 (N_15725,N_13565,N_13805);
and U15726 (N_15726,N_12011,N_12145);
or U15727 (N_15727,N_12354,N_13252);
nand U15728 (N_15728,N_13371,N_13601);
nand U15729 (N_15729,N_12896,N_12056);
xor U15730 (N_15730,N_13382,N_13568);
or U15731 (N_15731,N_13739,N_13233);
xor U15732 (N_15732,N_13078,N_13209);
and U15733 (N_15733,N_13974,N_13670);
nor U15734 (N_15734,N_13769,N_12686);
and U15735 (N_15735,N_12979,N_13600);
or U15736 (N_15736,N_12300,N_12867);
nor U15737 (N_15737,N_13849,N_13442);
xor U15738 (N_15738,N_12289,N_13077);
or U15739 (N_15739,N_12150,N_12544);
xor U15740 (N_15740,N_12649,N_13612);
xor U15741 (N_15741,N_12522,N_12385);
nor U15742 (N_15742,N_12183,N_13714);
nor U15743 (N_15743,N_13627,N_13186);
or U15744 (N_15744,N_13523,N_13796);
and U15745 (N_15745,N_13108,N_12092);
and U15746 (N_15746,N_12245,N_12270);
xor U15747 (N_15747,N_12927,N_13255);
or U15748 (N_15748,N_13262,N_12787);
nor U15749 (N_15749,N_12945,N_12848);
nand U15750 (N_15750,N_13832,N_12463);
xor U15751 (N_15751,N_12316,N_12286);
xnor U15752 (N_15752,N_13698,N_12836);
nor U15753 (N_15753,N_13524,N_12590);
nand U15754 (N_15754,N_12594,N_13640);
and U15755 (N_15755,N_13300,N_13560);
and U15756 (N_15756,N_12442,N_13085);
or U15757 (N_15757,N_12026,N_13506);
and U15758 (N_15758,N_13527,N_12996);
and U15759 (N_15759,N_12658,N_13747);
xor U15760 (N_15760,N_13955,N_13567);
nor U15761 (N_15761,N_13046,N_12982);
and U15762 (N_15762,N_13291,N_12202);
nor U15763 (N_15763,N_12254,N_13480);
xnor U15764 (N_15764,N_13473,N_13762);
and U15765 (N_15765,N_13422,N_13141);
or U15766 (N_15766,N_12828,N_13732);
or U15767 (N_15767,N_13134,N_12544);
or U15768 (N_15768,N_12974,N_12921);
nand U15769 (N_15769,N_13329,N_12464);
xnor U15770 (N_15770,N_13910,N_13726);
xnor U15771 (N_15771,N_13276,N_13427);
nand U15772 (N_15772,N_13958,N_13243);
xnor U15773 (N_15773,N_12243,N_13450);
and U15774 (N_15774,N_13361,N_13490);
or U15775 (N_15775,N_12833,N_13166);
nand U15776 (N_15776,N_13269,N_13152);
xnor U15777 (N_15777,N_12467,N_13245);
and U15778 (N_15778,N_12662,N_13979);
or U15779 (N_15779,N_12370,N_13831);
nand U15780 (N_15780,N_13280,N_13785);
nand U15781 (N_15781,N_12405,N_13482);
nor U15782 (N_15782,N_12736,N_13618);
nand U15783 (N_15783,N_13001,N_12272);
or U15784 (N_15784,N_12122,N_12416);
or U15785 (N_15785,N_12632,N_13399);
and U15786 (N_15786,N_13181,N_12293);
nor U15787 (N_15787,N_13312,N_12687);
nand U15788 (N_15788,N_12261,N_13515);
nor U15789 (N_15789,N_12409,N_13657);
and U15790 (N_15790,N_12837,N_13557);
nand U15791 (N_15791,N_12803,N_12824);
xor U15792 (N_15792,N_12683,N_13758);
or U15793 (N_15793,N_13632,N_12920);
or U15794 (N_15794,N_13740,N_12122);
nand U15795 (N_15795,N_12187,N_13537);
and U15796 (N_15796,N_12858,N_12882);
nand U15797 (N_15797,N_13717,N_13099);
nand U15798 (N_15798,N_13663,N_13190);
nand U15799 (N_15799,N_12792,N_13109);
nand U15800 (N_15800,N_13056,N_13176);
and U15801 (N_15801,N_12557,N_12804);
xor U15802 (N_15802,N_12712,N_12694);
and U15803 (N_15803,N_13189,N_13546);
or U15804 (N_15804,N_13227,N_12879);
or U15805 (N_15805,N_12619,N_13803);
xor U15806 (N_15806,N_13361,N_13718);
nand U15807 (N_15807,N_12217,N_13854);
and U15808 (N_15808,N_13630,N_13740);
nor U15809 (N_15809,N_12195,N_12547);
or U15810 (N_15810,N_12610,N_13653);
nor U15811 (N_15811,N_13517,N_12674);
and U15812 (N_15812,N_12523,N_12429);
nor U15813 (N_15813,N_13266,N_13746);
nor U15814 (N_15814,N_12142,N_13294);
nor U15815 (N_15815,N_12569,N_13639);
xnor U15816 (N_15816,N_12023,N_12877);
nand U15817 (N_15817,N_12631,N_13029);
and U15818 (N_15818,N_12812,N_13414);
and U15819 (N_15819,N_12767,N_13338);
xnor U15820 (N_15820,N_13703,N_12273);
or U15821 (N_15821,N_13705,N_13336);
or U15822 (N_15822,N_13195,N_13240);
nor U15823 (N_15823,N_13856,N_13369);
xnor U15824 (N_15824,N_13362,N_13624);
xor U15825 (N_15825,N_12571,N_13818);
nor U15826 (N_15826,N_12121,N_13632);
nor U15827 (N_15827,N_12198,N_13381);
nor U15828 (N_15828,N_13025,N_13490);
nor U15829 (N_15829,N_12246,N_12653);
nand U15830 (N_15830,N_13561,N_12890);
nand U15831 (N_15831,N_12867,N_12833);
nand U15832 (N_15832,N_13651,N_12256);
nor U15833 (N_15833,N_12578,N_12793);
nor U15834 (N_15834,N_12348,N_12730);
xnor U15835 (N_15835,N_12315,N_13728);
nand U15836 (N_15836,N_12057,N_13028);
xor U15837 (N_15837,N_13404,N_12657);
or U15838 (N_15838,N_13152,N_13084);
nand U15839 (N_15839,N_12527,N_13900);
nor U15840 (N_15840,N_13354,N_12672);
or U15841 (N_15841,N_13651,N_12842);
nor U15842 (N_15842,N_12025,N_13685);
nand U15843 (N_15843,N_12497,N_13543);
xnor U15844 (N_15844,N_13085,N_12004);
nand U15845 (N_15845,N_13556,N_12503);
or U15846 (N_15846,N_13755,N_13846);
nand U15847 (N_15847,N_12302,N_13304);
nand U15848 (N_15848,N_13871,N_12515);
nor U15849 (N_15849,N_13774,N_12823);
and U15850 (N_15850,N_13945,N_12070);
nand U15851 (N_15851,N_13922,N_12792);
and U15852 (N_15852,N_12898,N_13541);
or U15853 (N_15853,N_13719,N_12998);
xnor U15854 (N_15854,N_13206,N_13629);
nand U15855 (N_15855,N_13578,N_13291);
or U15856 (N_15856,N_13803,N_12090);
nor U15857 (N_15857,N_12000,N_12977);
and U15858 (N_15858,N_13631,N_13877);
nand U15859 (N_15859,N_12638,N_12608);
and U15860 (N_15860,N_13831,N_13695);
nor U15861 (N_15861,N_12023,N_13365);
xor U15862 (N_15862,N_12433,N_13918);
and U15863 (N_15863,N_12855,N_13871);
nor U15864 (N_15864,N_12855,N_12188);
or U15865 (N_15865,N_13045,N_12450);
nand U15866 (N_15866,N_12281,N_12830);
nand U15867 (N_15867,N_13400,N_12831);
and U15868 (N_15868,N_13795,N_12427);
xnor U15869 (N_15869,N_13863,N_12626);
nand U15870 (N_15870,N_12053,N_12846);
and U15871 (N_15871,N_12418,N_12573);
nor U15872 (N_15872,N_12749,N_12315);
and U15873 (N_15873,N_12662,N_13251);
and U15874 (N_15874,N_13077,N_13149);
xnor U15875 (N_15875,N_12288,N_12986);
xnor U15876 (N_15876,N_13226,N_12058);
xnor U15877 (N_15877,N_13578,N_13009);
nand U15878 (N_15878,N_12267,N_12000);
nor U15879 (N_15879,N_12791,N_12173);
nand U15880 (N_15880,N_13566,N_13397);
nor U15881 (N_15881,N_12081,N_12972);
nor U15882 (N_15882,N_13861,N_12496);
nand U15883 (N_15883,N_13075,N_13631);
nor U15884 (N_15884,N_12001,N_13105);
nand U15885 (N_15885,N_12835,N_13638);
nand U15886 (N_15886,N_12282,N_13264);
xnor U15887 (N_15887,N_12646,N_13082);
or U15888 (N_15888,N_13226,N_13468);
nor U15889 (N_15889,N_13607,N_12533);
or U15890 (N_15890,N_13673,N_13443);
nor U15891 (N_15891,N_12218,N_12794);
nand U15892 (N_15892,N_12306,N_12324);
or U15893 (N_15893,N_12705,N_13967);
nand U15894 (N_15894,N_13929,N_13237);
nor U15895 (N_15895,N_12422,N_13287);
xnor U15896 (N_15896,N_12066,N_12285);
or U15897 (N_15897,N_13986,N_13199);
xor U15898 (N_15898,N_13259,N_13718);
nor U15899 (N_15899,N_13641,N_12623);
nand U15900 (N_15900,N_12116,N_13141);
nor U15901 (N_15901,N_12653,N_12843);
xor U15902 (N_15902,N_12108,N_13146);
nand U15903 (N_15903,N_13218,N_12825);
nand U15904 (N_15904,N_12783,N_12776);
or U15905 (N_15905,N_13797,N_13308);
xnor U15906 (N_15906,N_12100,N_12140);
xor U15907 (N_15907,N_12842,N_13162);
nand U15908 (N_15908,N_13352,N_13935);
nand U15909 (N_15909,N_13650,N_13325);
xnor U15910 (N_15910,N_12140,N_13141);
or U15911 (N_15911,N_13665,N_13532);
xnor U15912 (N_15912,N_12351,N_13071);
nand U15913 (N_15913,N_12516,N_13713);
nand U15914 (N_15914,N_12583,N_12657);
nand U15915 (N_15915,N_13192,N_12248);
and U15916 (N_15916,N_13955,N_13543);
nor U15917 (N_15917,N_13564,N_13800);
and U15918 (N_15918,N_13687,N_12499);
nand U15919 (N_15919,N_13010,N_13804);
or U15920 (N_15920,N_12821,N_12373);
and U15921 (N_15921,N_12431,N_13033);
and U15922 (N_15922,N_12013,N_12204);
nand U15923 (N_15923,N_12559,N_12754);
nor U15924 (N_15924,N_12047,N_12754);
nand U15925 (N_15925,N_12820,N_12957);
nand U15926 (N_15926,N_13488,N_13520);
xor U15927 (N_15927,N_13906,N_13291);
or U15928 (N_15928,N_12396,N_12863);
nor U15929 (N_15929,N_12424,N_12150);
or U15930 (N_15930,N_13383,N_12502);
and U15931 (N_15931,N_12459,N_12940);
nand U15932 (N_15932,N_12374,N_13876);
or U15933 (N_15933,N_13508,N_12170);
xor U15934 (N_15934,N_12687,N_13953);
xnor U15935 (N_15935,N_12893,N_12916);
or U15936 (N_15936,N_13252,N_12342);
xor U15937 (N_15937,N_13835,N_13236);
nor U15938 (N_15938,N_12111,N_13129);
or U15939 (N_15939,N_12214,N_13598);
and U15940 (N_15940,N_13341,N_12833);
xnor U15941 (N_15941,N_13996,N_13942);
nor U15942 (N_15942,N_13391,N_13923);
and U15943 (N_15943,N_13119,N_13854);
or U15944 (N_15944,N_13096,N_13439);
or U15945 (N_15945,N_13414,N_12998);
nand U15946 (N_15946,N_13576,N_13548);
xor U15947 (N_15947,N_12794,N_12520);
and U15948 (N_15948,N_13883,N_13297);
or U15949 (N_15949,N_13711,N_13122);
and U15950 (N_15950,N_13083,N_13959);
xor U15951 (N_15951,N_12150,N_12732);
nor U15952 (N_15952,N_12274,N_12203);
or U15953 (N_15953,N_12174,N_13661);
nand U15954 (N_15954,N_13726,N_12033);
nand U15955 (N_15955,N_13373,N_13374);
or U15956 (N_15956,N_13809,N_12292);
or U15957 (N_15957,N_12723,N_12249);
and U15958 (N_15958,N_12348,N_13367);
or U15959 (N_15959,N_12637,N_12154);
or U15960 (N_15960,N_13709,N_13758);
and U15961 (N_15961,N_13135,N_13173);
xor U15962 (N_15962,N_13796,N_13243);
nor U15963 (N_15963,N_12761,N_12164);
and U15964 (N_15964,N_12961,N_13788);
or U15965 (N_15965,N_13499,N_13728);
nor U15966 (N_15966,N_12103,N_12446);
nand U15967 (N_15967,N_12846,N_12221);
nor U15968 (N_15968,N_13478,N_13532);
xor U15969 (N_15969,N_13434,N_13107);
or U15970 (N_15970,N_12646,N_13485);
nand U15971 (N_15971,N_12277,N_13732);
nor U15972 (N_15972,N_12412,N_13264);
nand U15973 (N_15973,N_13378,N_13000);
nor U15974 (N_15974,N_12160,N_13937);
and U15975 (N_15975,N_13537,N_13581);
xor U15976 (N_15976,N_13422,N_12515);
xnor U15977 (N_15977,N_13288,N_13188);
or U15978 (N_15978,N_12349,N_13394);
nor U15979 (N_15979,N_12458,N_12463);
nand U15980 (N_15980,N_12038,N_13380);
and U15981 (N_15981,N_13640,N_12890);
and U15982 (N_15982,N_13731,N_12604);
nor U15983 (N_15983,N_12731,N_12963);
nor U15984 (N_15984,N_13251,N_13756);
xnor U15985 (N_15985,N_13342,N_13605);
nor U15986 (N_15986,N_12663,N_13829);
and U15987 (N_15987,N_13146,N_12748);
or U15988 (N_15988,N_12189,N_13102);
or U15989 (N_15989,N_13614,N_13870);
nor U15990 (N_15990,N_13196,N_12576);
and U15991 (N_15991,N_12053,N_12774);
nor U15992 (N_15992,N_13250,N_13931);
and U15993 (N_15993,N_12876,N_12778);
or U15994 (N_15994,N_13434,N_13296);
nand U15995 (N_15995,N_13440,N_12572);
nand U15996 (N_15996,N_12765,N_13832);
and U15997 (N_15997,N_13014,N_13129);
xor U15998 (N_15998,N_12196,N_13924);
nand U15999 (N_15999,N_12595,N_12859);
xor U16000 (N_16000,N_14065,N_14954);
and U16001 (N_16001,N_14183,N_14940);
xnor U16002 (N_16002,N_15872,N_15032);
nand U16003 (N_16003,N_14621,N_15820);
or U16004 (N_16004,N_15294,N_14222);
nand U16005 (N_16005,N_15363,N_15585);
or U16006 (N_16006,N_14857,N_14879);
and U16007 (N_16007,N_14055,N_14289);
or U16008 (N_16008,N_14429,N_14081);
or U16009 (N_16009,N_15384,N_14618);
or U16010 (N_16010,N_15853,N_14273);
nor U16011 (N_16011,N_15062,N_15277);
xnor U16012 (N_16012,N_14852,N_14450);
and U16013 (N_16013,N_15567,N_14258);
and U16014 (N_16014,N_15347,N_15008);
xnor U16015 (N_16015,N_15026,N_15058);
xnor U16016 (N_16016,N_15126,N_14474);
or U16017 (N_16017,N_15275,N_14306);
nor U16018 (N_16018,N_14607,N_14752);
nand U16019 (N_16019,N_15782,N_15159);
or U16020 (N_16020,N_15776,N_14919);
nand U16021 (N_16021,N_15387,N_15768);
or U16022 (N_16022,N_14294,N_14272);
or U16023 (N_16023,N_15259,N_14430);
xnor U16024 (N_16024,N_14234,N_14800);
and U16025 (N_16025,N_15166,N_14604);
nand U16026 (N_16026,N_14275,N_14544);
and U16027 (N_16027,N_15681,N_15167);
and U16028 (N_16028,N_14851,N_15056);
nand U16029 (N_16029,N_14768,N_14286);
nand U16030 (N_16030,N_15508,N_14652);
or U16031 (N_16031,N_14682,N_14391);
nand U16032 (N_16032,N_14401,N_14611);
nor U16033 (N_16033,N_15688,N_14263);
xnor U16034 (N_16034,N_14021,N_15727);
or U16035 (N_16035,N_15705,N_14188);
nor U16036 (N_16036,N_14063,N_14714);
nand U16037 (N_16037,N_15466,N_14190);
and U16038 (N_16038,N_14358,N_15946);
and U16039 (N_16039,N_15541,N_14482);
and U16040 (N_16040,N_14526,N_15002);
or U16041 (N_16041,N_15645,N_14127);
and U16042 (N_16042,N_15865,N_14601);
nand U16043 (N_16043,N_15579,N_15182);
or U16044 (N_16044,N_14157,N_15692);
xor U16045 (N_16045,N_15754,N_15119);
and U16046 (N_16046,N_14005,N_15391);
nor U16047 (N_16047,N_14584,N_14766);
xnor U16048 (N_16048,N_14783,N_15813);
nor U16049 (N_16049,N_15817,N_14855);
nand U16050 (N_16050,N_15532,N_15918);
or U16051 (N_16051,N_14916,N_15818);
or U16052 (N_16052,N_15824,N_14168);
nand U16053 (N_16053,N_14507,N_14269);
and U16054 (N_16054,N_15805,N_15267);
and U16055 (N_16055,N_15691,N_14962);
and U16056 (N_16056,N_15891,N_15697);
and U16057 (N_16057,N_14945,N_15402);
or U16058 (N_16058,N_14773,N_14200);
nor U16059 (N_16059,N_14000,N_14178);
nand U16060 (N_16060,N_14895,N_14575);
and U16061 (N_16061,N_14339,N_15673);
nand U16062 (N_16062,N_14463,N_14672);
and U16063 (N_16063,N_14284,N_14461);
nor U16064 (N_16064,N_14525,N_14560);
nand U16065 (N_16065,N_15979,N_15368);
xnor U16066 (N_16066,N_15765,N_14785);
xnor U16067 (N_16067,N_15665,N_14078);
nor U16068 (N_16068,N_15897,N_14161);
and U16069 (N_16069,N_15844,N_14769);
nor U16070 (N_16070,N_14442,N_15354);
xor U16071 (N_16071,N_15662,N_14781);
nand U16072 (N_16072,N_15473,N_14405);
nand U16073 (N_16073,N_15395,N_15380);
nor U16074 (N_16074,N_14208,N_14014);
nand U16075 (N_16075,N_15509,N_15537);
xnor U16076 (N_16076,N_14641,N_15235);
and U16077 (N_16077,N_15086,N_14364);
nand U16078 (N_16078,N_15792,N_14943);
and U16079 (N_16079,N_14343,N_15256);
and U16080 (N_16080,N_14197,N_14661);
and U16081 (N_16081,N_15147,N_15513);
or U16082 (N_16082,N_15006,N_14225);
and U16083 (N_16083,N_15299,N_15366);
or U16084 (N_16084,N_15201,N_15666);
xnor U16085 (N_16085,N_14288,N_14293);
nor U16086 (N_16086,N_14932,N_14624);
xor U16087 (N_16087,N_15869,N_14907);
and U16088 (N_16088,N_15791,N_15411);
nand U16089 (N_16089,N_15640,N_15877);
nand U16090 (N_16090,N_15131,N_14828);
and U16091 (N_16091,N_14236,N_15452);
nand U16092 (N_16092,N_14988,N_15515);
and U16093 (N_16093,N_14230,N_14912);
nor U16094 (N_16094,N_15485,N_15359);
and U16095 (N_16095,N_15575,N_15652);
or U16096 (N_16096,N_14131,N_15752);
or U16097 (N_16097,N_14497,N_15350);
xnor U16098 (N_16098,N_14321,N_14169);
and U16099 (N_16099,N_14698,N_15399);
xor U16100 (N_16100,N_15732,N_15634);
or U16101 (N_16101,N_15507,N_14252);
and U16102 (N_16102,N_14172,N_15178);
nand U16103 (N_16103,N_14092,N_15322);
nand U16104 (N_16104,N_14586,N_15572);
or U16105 (N_16105,N_15557,N_14413);
nand U16106 (N_16106,N_14559,N_14136);
nor U16107 (N_16107,N_15139,N_15687);
or U16108 (N_16108,N_14244,N_14340);
nand U16109 (N_16109,N_14040,N_14483);
and U16110 (N_16110,N_15238,N_15472);
xnor U16111 (N_16111,N_14490,N_15834);
and U16112 (N_16112,N_15065,N_15904);
xor U16113 (N_16113,N_15079,N_14439);
or U16114 (N_16114,N_15686,N_14823);
xor U16115 (N_16115,N_14900,N_14326);
nand U16116 (N_16116,N_15760,N_14148);
or U16117 (N_16117,N_14342,N_14026);
xnor U16118 (N_16118,N_15084,N_15262);
nor U16119 (N_16119,N_15096,N_15200);
xor U16120 (N_16120,N_14281,N_14674);
nand U16121 (N_16121,N_14170,N_15733);
or U16122 (N_16122,N_14129,N_15106);
xor U16123 (N_16123,N_15528,N_15312);
xnor U16124 (N_16124,N_15048,N_15220);
nor U16125 (N_16125,N_14084,N_15708);
nor U16126 (N_16126,N_15954,N_15955);
or U16127 (N_16127,N_15713,N_14826);
xnor U16128 (N_16128,N_14995,N_15751);
or U16129 (N_16129,N_15598,N_14735);
and U16130 (N_16130,N_14382,N_15854);
or U16131 (N_16131,N_15264,N_15371);
xor U16132 (N_16132,N_15790,N_15547);
nand U16133 (N_16133,N_15160,N_15231);
and U16134 (N_16134,N_14632,N_14726);
nor U16135 (N_16135,N_15801,N_14285);
nand U16136 (N_16136,N_15292,N_14181);
nand U16137 (N_16137,N_14419,N_15555);
and U16138 (N_16138,N_15203,N_14082);
xor U16139 (N_16139,N_15566,N_14761);
xnor U16140 (N_16140,N_14502,N_15629);
nand U16141 (N_16141,N_15544,N_14791);
and U16142 (N_16142,N_14212,N_14116);
and U16143 (N_16143,N_15110,N_15206);
nand U16144 (N_16144,N_15621,N_15460);
and U16145 (N_16145,N_15306,N_15193);
nand U16146 (N_16146,N_15367,N_15280);
nand U16147 (N_16147,N_15356,N_15029);
nand U16148 (N_16148,N_14570,N_15448);
xor U16149 (N_16149,N_15632,N_14716);
and U16150 (N_16150,N_14941,N_14509);
nor U16151 (N_16151,N_14989,N_15064);
nor U16152 (N_16152,N_14410,N_14144);
nor U16153 (N_16153,N_14378,N_15775);
or U16154 (N_16154,N_15578,N_14087);
nand U16155 (N_16155,N_15385,N_15156);
or U16156 (N_16156,N_15827,N_15923);
nor U16157 (N_16157,N_14747,N_15145);
nor U16158 (N_16158,N_15802,N_15573);
and U16159 (N_16159,N_14369,N_14274);
nand U16160 (N_16160,N_14512,N_14639);
xor U16161 (N_16161,N_14583,N_15531);
nand U16162 (N_16162,N_14438,N_15471);
xnor U16163 (N_16163,N_15021,N_14444);
and U16164 (N_16164,N_15533,N_14185);
xor U16165 (N_16165,N_14673,N_15761);
xor U16166 (N_16166,N_15878,N_15043);
xnor U16167 (N_16167,N_14891,N_15137);
or U16168 (N_16168,N_14859,N_14786);
and U16169 (N_16169,N_14540,N_15462);
and U16170 (N_16170,N_15100,N_14455);
xnor U16171 (N_16171,N_15511,N_14911);
or U16172 (N_16172,N_15720,N_14204);
or U16173 (N_16173,N_15153,N_15631);
nand U16174 (N_16174,N_15922,N_15187);
or U16175 (N_16175,N_15024,N_14479);
nor U16176 (N_16176,N_15896,N_15653);
xor U16177 (N_16177,N_15647,N_14612);
nor U16178 (N_16178,N_14635,N_15022);
xor U16179 (N_16179,N_15154,N_14390);
and U16180 (N_16180,N_15076,N_14523);
xor U16181 (N_16181,N_14018,N_14603);
nor U16182 (N_16182,N_15659,N_14447);
and U16183 (N_16183,N_14189,N_14901);
or U16184 (N_16184,N_15469,N_14904);
and U16185 (N_16185,N_15669,N_14112);
nand U16186 (N_16186,N_15317,N_15826);
nand U16187 (N_16187,N_15444,N_14022);
nor U16188 (N_16188,N_14742,N_14610);
and U16189 (N_16189,N_14443,N_15906);
nor U16190 (N_16190,N_15502,N_15229);
nand U16191 (N_16191,N_15626,N_15221);
xnor U16192 (N_16192,N_15650,N_15376);
or U16193 (N_16193,N_15935,N_14505);
nor U16194 (N_16194,N_14515,N_14840);
and U16195 (N_16195,N_15672,N_14566);
nor U16196 (N_16196,N_14558,N_15773);
nor U16197 (N_16197,N_15983,N_15516);
nand U16198 (N_16198,N_15842,N_15630);
xnor U16199 (N_16199,N_15902,N_15493);
or U16200 (N_16200,N_15287,N_15044);
and U16201 (N_16201,N_15253,N_14744);
nand U16202 (N_16202,N_14062,N_14134);
nor U16203 (N_16203,N_15789,N_15974);
nand U16204 (N_16204,N_15345,N_15426);
nor U16205 (N_16205,N_14992,N_14520);
or U16206 (N_16206,N_14167,N_14676);
xor U16207 (N_16207,N_14217,N_14915);
or U16208 (N_16208,N_14867,N_15702);
xnor U16209 (N_16209,N_14478,N_14693);
nand U16210 (N_16210,N_14871,N_15241);
and U16211 (N_16211,N_15192,N_15348);
xor U16212 (N_16212,N_15216,N_14598);
and U16213 (N_16213,N_14008,N_14500);
and U16214 (N_16214,N_15975,N_15524);
or U16215 (N_16215,N_15604,N_15726);
or U16216 (N_16216,N_15198,N_14657);
nor U16217 (N_16217,N_14597,N_15082);
and U16218 (N_16218,N_15454,N_15795);
and U16219 (N_16219,N_14395,N_14346);
xnor U16220 (N_16220,N_15181,N_15311);
and U16221 (N_16221,N_15693,N_14875);
xnor U16222 (N_16222,N_14171,N_15793);
nand U16223 (N_16223,N_14383,N_14532);
nand U16224 (N_16224,N_14671,N_15675);
or U16225 (N_16225,N_14408,N_15457);
nand U16226 (N_16226,N_14060,N_15398);
or U16227 (N_16227,N_15085,N_15859);
xnor U16228 (N_16228,N_15849,N_14513);
and U16229 (N_16229,N_14663,N_14357);
or U16230 (N_16230,N_14414,N_14554);
and U16231 (N_16231,N_14832,N_14743);
nand U16232 (N_16232,N_14910,N_14514);
nor U16233 (N_16233,N_15617,N_14812);
and U16234 (N_16234,N_14240,N_15487);
and U16235 (N_16235,N_15329,N_15179);
nor U16236 (N_16236,N_14261,N_14649);
or U16237 (N_16237,N_14978,N_14277);
and U16238 (N_16238,N_15199,N_15577);
nand U16239 (N_16239,N_14035,N_14276);
xor U16240 (N_16240,N_14638,N_14563);
nand U16241 (N_16241,N_15595,N_15397);
xnor U16242 (N_16242,N_14806,N_15717);
or U16243 (N_16243,N_15207,N_15046);
and U16244 (N_16244,N_15816,N_14206);
xnor U16245 (N_16245,N_15736,N_15871);
xor U16246 (N_16246,N_14790,N_14530);
or U16247 (N_16247,N_14211,N_14475);
nor U16248 (N_16248,N_14874,N_14847);
xnor U16249 (N_16249,N_14881,N_14980);
nand U16250 (N_16250,N_14352,N_14938);
nor U16251 (N_16251,N_14917,N_14268);
nor U16252 (N_16252,N_15459,N_15352);
xnor U16253 (N_16253,N_14366,N_15386);
or U16254 (N_16254,N_15711,N_15165);
nor U16255 (N_16255,N_14986,N_14634);
nor U16256 (N_16256,N_14887,N_15441);
nand U16257 (N_16257,N_14436,N_14156);
and U16258 (N_16258,N_14220,N_14906);
xnor U16259 (N_16259,N_14587,N_14377);
xor U16260 (N_16260,N_15176,N_15962);
and U16261 (N_16261,N_14754,N_14445);
and U16262 (N_16262,N_14098,N_14905);
and U16263 (N_16263,N_14424,N_14247);
nor U16264 (N_16264,N_15186,N_14020);
or U16265 (N_16265,N_14555,N_14884);
nor U16266 (N_16266,N_15045,N_14025);
nand U16267 (N_16267,N_15781,N_14224);
nand U16268 (N_16268,N_14071,N_14259);
or U16269 (N_16269,N_14701,N_15445);
nor U16270 (N_16270,N_14070,N_14088);
or U16271 (N_16271,N_14792,N_15494);
and U16272 (N_16272,N_14334,N_15224);
nand U16273 (N_16273,N_14402,N_14933);
nand U16274 (N_16274,N_15033,N_15934);
nor U16275 (N_16275,N_15476,N_14468);
nand U16276 (N_16276,N_15568,N_14922);
nor U16277 (N_16277,N_14925,N_14044);
and U16278 (N_16278,N_14556,N_14101);
nand U16279 (N_16279,N_14573,N_15234);
and U16280 (N_16280,N_15608,N_14564);
xor U16281 (N_16281,N_15310,N_15778);
or U16282 (N_16282,N_14042,N_15680);
and U16283 (N_16283,N_14964,N_14238);
nor U16284 (N_16284,N_15709,N_14582);
nand U16285 (N_16285,N_15339,N_14015);
xnor U16286 (N_16286,N_15796,N_15050);
and U16287 (N_16287,N_15288,N_14903);
or U16288 (N_16288,N_15836,N_14282);
nor U16289 (N_16289,N_15808,N_14458);
xor U16290 (N_16290,N_15439,N_14074);
and U16291 (N_16291,N_14311,N_15609);
xnor U16292 (N_16292,N_15077,N_14387);
nand U16293 (N_16293,N_15349,N_14797);
or U16294 (N_16294,N_15747,N_15093);
or U16295 (N_16295,N_15941,N_14868);
nand U16296 (N_16296,N_14361,N_14972);
nor U16297 (N_16297,N_15880,N_15148);
xnor U16298 (N_16298,N_15898,N_14923);
xnor U16299 (N_16299,N_15542,N_15116);
or U16300 (N_16300,N_14307,N_15840);
or U16301 (N_16301,N_14034,N_14692);
and U16302 (N_16302,N_14707,N_14122);
or U16303 (N_16303,N_15641,N_14368);
and U16304 (N_16304,N_14163,N_15970);
xnor U16305 (N_16305,N_15060,N_14699);
nor U16306 (N_16306,N_15307,N_14232);
xor U16307 (N_16307,N_14898,N_15945);
nor U16308 (N_16308,N_15111,N_14821);
nor U16309 (N_16309,N_15581,N_15510);
nand U16310 (N_16310,N_15741,N_15453);
nand U16311 (N_16311,N_14741,N_14386);
nand U16312 (N_16312,N_15197,N_15185);
or U16313 (N_16313,N_14837,N_14600);
nor U16314 (N_16314,N_14375,N_14623);
or U16315 (N_16315,N_15240,N_15416);
and U16316 (N_16316,N_15276,N_15924);
and U16317 (N_16317,N_14524,N_14608);
nor U16318 (N_16318,N_14985,N_15657);
xnor U16319 (N_16319,N_14976,N_15314);
xor U16320 (N_16320,N_14213,N_14918);
and U16321 (N_16321,N_14757,N_14924);
nand U16322 (N_16322,N_15097,N_15562);
and U16323 (N_16323,N_14813,N_14158);
nor U16324 (N_16324,N_15500,N_15987);
or U16325 (N_16325,N_15155,N_14054);
or U16326 (N_16326,N_14333,N_14684);
nor U16327 (N_16327,N_15249,N_14409);
or U16328 (N_16328,N_14899,N_15740);
and U16329 (N_16329,N_15461,N_15829);
and U16330 (N_16330,N_15195,N_15035);
nor U16331 (N_16331,N_14567,N_15489);
xor U16332 (N_16332,N_14728,N_15638);
and U16333 (N_16333,N_15936,N_15841);
and U16334 (N_16334,N_14207,N_15788);
nor U16335 (N_16335,N_15422,N_15756);
xor U16336 (N_16336,N_15564,N_15921);
nand U16337 (N_16337,N_14376,N_14725);
nor U16338 (N_16338,N_14271,N_15215);
and U16339 (N_16339,N_14001,N_15889);
nor U16340 (N_16340,N_14815,N_14324);
and U16341 (N_16341,N_15973,N_15695);
xor U16342 (N_16342,N_14680,N_15858);
and U16343 (N_16343,N_15677,N_14820);
nor U16344 (N_16344,N_15978,N_14384);
or U16345 (N_16345,N_15619,N_15755);
and U16346 (N_16346,N_15625,N_14968);
nand U16347 (N_16347,N_14605,N_15302);
nor U16348 (N_16348,N_14838,N_15690);
and U16349 (N_16349,N_15830,N_14648);
nor U16350 (N_16350,N_15353,N_14498);
nand U16351 (N_16351,N_15143,N_14090);
nor U16352 (N_16352,N_15714,N_15944);
xnor U16353 (N_16353,N_14546,N_14998);
nand U16354 (N_16354,N_14495,N_15016);
nor U16355 (N_16355,N_14446,N_14394);
nand U16356 (N_16356,N_15558,N_14591);
nand U16357 (N_16357,N_14727,N_15117);
xnor U16358 (N_16358,N_15614,N_15260);
xnor U16359 (N_16359,N_14825,N_14441);
xor U16360 (N_16360,N_15696,N_15540);
or U16361 (N_16361,N_15456,N_15912);
or U16362 (N_16362,N_15012,N_14568);
nor U16363 (N_16363,N_14314,N_15539);
xor U16364 (N_16364,N_15316,N_15226);
or U16365 (N_16365,N_14338,N_15990);
nor U16366 (N_16366,N_15779,N_14335);
or U16367 (N_16367,N_14109,N_15698);
and U16368 (N_16368,N_14733,N_15301);
nand U16369 (N_16369,N_14543,N_14897);
nand U16370 (N_16370,N_15730,N_15451);
nor U16371 (N_16371,N_15455,N_14107);
xnor U16372 (N_16372,N_15501,N_15560);
and U16373 (N_16373,N_14929,N_14243);
nor U16374 (N_16374,N_14609,N_15414);
xnor U16375 (N_16375,N_15679,N_14336);
nand U16376 (N_16376,N_14047,N_15704);
or U16377 (N_16377,N_14731,N_15027);
or U16378 (N_16378,N_14266,N_15815);
nor U16379 (N_16379,N_15994,N_14713);
nor U16380 (N_16380,N_14287,N_15053);
and U16381 (N_16381,N_14774,N_15724);
or U16382 (N_16382,N_15429,N_14075);
nand U16383 (N_16383,N_15170,N_14669);
nand U16384 (N_16384,N_15248,N_14719);
nand U16385 (N_16385,N_15092,N_14872);
or U16386 (N_16386,N_15832,N_14404);
xor U16387 (N_16387,N_15895,N_15252);
nor U16388 (N_16388,N_15406,N_14691);
or U16389 (N_16389,N_15437,N_15289);
nand U16390 (N_16390,N_14440,N_15000);
nand U16391 (N_16391,N_15383,N_15098);
xor U16392 (N_16392,N_15342,N_14646);
nand U16393 (N_16393,N_14734,N_15504);
nor U16394 (N_16394,N_15019,N_15886);
or U16395 (N_16395,N_15965,N_15514);
and U16396 (N_16396,N_15599,N_14072);
xor U16397 (N_16397,N_14279,N_14961);
nor U16398 (N_16398,N_14548,N_15548);
nor U16399 (N_16399,N_14779,N_14640);
xnor U16400 (N_16400,N_14508,N_15482);
or U16401 (N_16401,N_15369,N_14689);
and U16402 (N_16402,N_15081,N_14374);
nand U16403 (N_16403,N_14969,N_14466);
and U16404 (N_16404,N_14533,N_14202);
nor U16405 (N_16405,N_14953,N_15318);
nor U16406 (N_16406,N_15588,N_14347);
nand U16407 (N_16407,N_14795,N_14192);
or U16408 (N_16408,N_15863,N_14705);
or U16409 (N_16409,N_15569,N_15723);
nor U16410 (N_16410,N_14085,N_15674);
nor U16411 (N_16411,N_15018,N_15963);
xor U16412 (N_16412,N_15209,N_15194);
or U16413 (N_16413,N_15900,N_14841);
and U16414 (N_16414,N_14073,N_15956);
xor U16415 (N_16415,N_14348,N_15251);
or U16416 (N_16416,N_15236,N_15710);
nand U16417 (N_16417,N_15338,N_15649);
xnor U16418 (N_16418,N_15377,N_15467);
or U16419 (N_16419,N_14330,N_15728);
or U16420 (N_16420,N_14146,N_14510);
or U16421 (N_16421,N_14746,N_15327);
or U16422 (N_16422,N_14367,N_15474);
nor U16423 (N_16423,N_15633,N_15150);
or U16424 (N_16424,N_14798,N_15556);
or U16425 (N_16425,N_14089,N_15561);
and U16426 (N_16426,N_14765,N_14951);
or U16427 (N_16427,N_14993,N_14878);
xor U16428 (N_16428,N_14118,N_14173);
or U16429 (N_16429,N_15703,N_15358);
nand U16430 (N_16430,N_15670,N_15757);
xnor U16431 (N_16431,N_14086,N_15847);
or U16432 (N_16432,N_14239,N_15133);
and U16433 (N_16433,N_14095,N_15188);
nor U16434 (N_16434,N_15623,N_14531);
and U16435 (N_16435,N_15417,N_14740);
or U16436 (N_16436,N_14249,N_15925);
nand U16437 (N_16437,N_14133,N_14010);
xnor U16438 (N_16438,N_15042,N_15225);
nand U16439 (N_16439,N_15161,N_14602);
nor U16440 (N_16440,N_15828,N_15146);
nand U16441 (N_16441,N_14755,N_15518);
nor U16442 (N_16442,N_15169,N_15468);
or U16443 (N_16443,N_15798,N_15587);
nor U16444 (N_16444,N_15066,N_14066);
nand U16445 (N_16445,N_15269,N_14399);
xnor U16446 (N_16446,N_15475,N_14542);
xor U16447 (N_16447,N_14406,N_14304);
nand U16448 (N_16448,N_14425,N_14106);
nor U16449 (N_16449,N_14103,N_14145);
nor U16450 (N_16450,N_14793,N_14198);
nor U16451 (N_16451,N_14827,N_14049);
or U16452 (N_16452,N_15010,N_14147);
nand U16453 (N_16453,N_15997,N_14599);
nor U16454 (N_16454,N_14117,N_14037);
and U16455 (N_16455,N_15597,N_14142);
or U16456 (N_16456,N_14308,N_15244);
or U16457 (N_16457,N_14350,N_14935);
nor U16458 (N_16458,N_15063,N_14028);
or U16459 (N_16459,N_15308,N_15857);
xor U16460 (N_16460,N_15694,N_14553);
or U16461 (N_16461,N_14778,N_15712);
and U16462 (N_16462,N_14873,N_14831);
nor U16463 (N_16463,N_14521,N_14331);
nor U16464 (N_16464,N_14569,N_15142);
xor U16465 (N_16465,N_15839,N_14050);
and U16466 (N_16466,N_14844,N_15202);
or U16467 (N_16467,N_15286,N_14996);
nor U16468 (N_16468,N_14416,N_15041);
nor U16469 (N_16469,N_15434,N_15603);
nor U16470 (N_16470,N_15162,N_15685);
and U16471 (N_16471,N_15953,N_14298);
nor U16472 (N_16472,N_14226,N_14856);
nand U16473 (N_16473,N_15636,N_14736);
nor U16474 (N_16474,N_14574,N_14004);
xor U16475 (N_16475,N_14228,N_15981);
nand U16476 (N_16476,N_14077,N_15243);
and U16477 (N_16477,N_14720,N_15001);
nand U16478 (N_16478,N_15479,N_14027);
and U16479 (N_16479,N_15804,N_15210);
xnor U16480 (N_16480,N_15109,N_14914);
and U16481 (N_16481,N_14114,N_15409);
xor U16482 (N_16482,N_15663,N_15438);
nor U16483 (N_16483,N_15774,N_15862);
and U16484 (N_16484,N_15919,N_14889);
or U16485 (N_16485,N_14162,N_15586);
and U16486 (N_16486,N_14024,N_15094);
and U16487 (N_16487,N_14760,N_14459);
or U16488 (N_16488,N_14472,N_14470);
xnor U16489 (N_16489,N_15876,N_14660);
nand U16490 (N_16490,N_14571,N_14987);
or U16491 (N_16491,N_14195,N_14315);
xnor U16492 (N_16492,N_15341,N_14764);
and U16493 (N_16493,N_15340,N_14477);
nand U16494 (N_16494,N_15388,N_14242);
nor U16495 (N_16495,N_14928,N_15103);
or U16496 (N_16496,N_14869,N_15622);
or U16497 (N_16497,N_14246,N_14184);
xnor U16498 (N_16498,N_14397,N_15591);
xor U16499 (N_16499,N_14448,N_15803);
nor U16500 (N_16500,N_14149,N_14164);
nor U16501 (N_16501,N_15957,N_14400);
nor U16502 (N_16502,N_15431,N_15204);
nand U16503 (N_16503,N_14006,N_15057);
nor U16504 (N_16504,N_15405,N_14865);
xnor U16505 (N_16505,N_15419,N_15725);
or U16506 (N_16506,N_14979,N_15393);
or U16507 (N_16507,N_14749,N_15282);
nor U16508 (N_16508,N_14141,N_14411);
and U16509 (N_16509,N_15932,N_14854);
nand U16510 (N_16510,N_14536,N_15122);
xnor U16511 (N_16511,N_14894,N_14694);
xor U16512 (N_16512,N_14363,N_14180);
nor U16513 (N_16513,N_14934,N_14829);
or U16514 (N_16514,N_14013,N_14418);
or U16515 (N_16515,N_14080,N_15447);
nor U16516 (N_16516,N_15620,N_15637);
or U16517 (N_16517,N_14876,N_15071);
and U16518 (N_16518,N_15257,N_14214);
and U16519 (N_16519,N_15554,N_15051);
nand U16520 (N_16520,N_15365,N_14805);
nor U16521 (N_16521,N_15835,N_15343);
nor U16522 (N_16522,N_15390,N_15279);
or U16523 (N_16523,N_15303,N_14313);
nor U16524 (N_16524,N_14633,N_14469);
or U16525 (N_16525,N_15324,N_15034);
nor U16526 (N_16526,N_14862,N_14808);
and U16527 (N_16527,N_14864,N_14944);
or U16528 (N_16528,N_15149,N_14102);
nor U16529 (N_16529,N_15361,N_15903);
and U16530 (N_16530,N_14007,N_14819);
nor U16531 (N_16531,N_14362,N_15731);
xor U16532 (N_16532,N_14830,N_15389);
nor U16533 (N_16533,N_15336,N_14329);
or U16534 (N_16534,N_15894,N_15966);
and U16535 (N_16535,N_14846,N_14627);
xnor U16536 (N_16536,N_14203,N_15007);
nor U16537 (N_16537,N_14538,N_14029);
nand U16538 (N_16538,N_14380,N_14892);
and U16539 (N_16539,N_14896,N_15960);
and U16540 (N_16540,N_14596,N_15770);
nor U16541 (N_16541,N_14836,N_15360);
and U16542 (N_16542,N_14654,N_14219);
and U16543 (N_16543,N_14166,N_14046);
xnor U16544 (N_16544,N_14299,N_15683);
nand U16545 (N_16545,N_15410,N_15700);
nor U16546 (N_16546,N_15769,N_14069);
or U16547 (N_16547,N_15580,N_15141);
xnor U16548 (N_16548,N_14421,N_15415);
or U16549 (N_16549,N_15090,N_15261);
nor U16550 (N_16550,N_14341,N_15744);
nor U16551 (N_16551,N_14955,N_14317);
xnor U16552 (N_16552,N_15223,N_15346);
or U16553 (N_16553,N_14465,N_14328);
and U16554 (N_16554,N_15615,N_14250);
and U16555 (N_16555,N_15701,N_15408);
and U16556 (N_16556,N_15285,N_14578);
and U16557 (N_16557,N_14360,N_15184);
or U16558 (N_16558,N_14799,N_15606);
or U16559 (N_16559,N_14686,N_15927);
nand U16560 (N_16560,N_14345,N_15811);
nand U16561 (N_16561,N_15601,N_14803);
xor U16562 (N_16562,N_15091,N_14517);
nor U16563 (N_16563,N_15247,N_14139);
nor U16564 (N_16564,N_14927,N_14677);
nand U16565 (N_16565,N_15047,N_15413);
and U16566 (N_16566,N_15483,N_15656);
nor U16567 (N_16567,N_15684,N_14312);
and U16568 (N_16568,N_15848,N_15861);
xor U16569 (N_16569,N_15913,N_14422);
nand U16570 (N_16570,N_14453,N_15646);
nand U16571 (N_16571,N_15233,N_14437);
nor U16572 (N_16572,N_15901,N_14093);
and U16573 (N_16573,N_14292,N_15884);
nor U16574 (N_16574,N_14280,N_15864);
xnor U16575 (N_16575,N_15982,N_14999);
or U16576 (N_16576,N_15470,N_14886);
nand U16577 (N_16577,N_15613,N_15612);
and U16578 (N_16578,N_14784,N_14143);
or U16579 (N_16579,N_15070,N_14950);
or U16580 (N_16580,N_15721,N_15078);
xnor U16581 (N_16581,N_15331,N_15095);
nor U16582 (N_16582,N_15173,N_15909);
xor U16583 (N_16583,N_15394,N_14460);
or U16584 (N_16584,N_14948,N_15738);
nor U16585 (N_16585,N_14511,N_15205);
and U16586 (N_16586,N_15976,N_14708);
or U16587 (N_16587,N_15964,N_14254);
and U16588 (N_16588,N_15984,N_15605);
nand U16589 (N_16589,N_15538,N_14971);
nor U16590 (N_16590,N_14858,N_15265);
nand U16591 (N_16591,N_14058,N_15425);
nor U16592 (N_16592,N_14751,N_15196);
and U16593 (N_16593,N_14381,N_15887);
or U16594 (N_16594,N_15490,N_14817);
xnor U16595 (N_16595,N_15972,N_15628);
and U16596 (N_16596,N_14264,N_14435);
xor U16597 (N_16597,N_15576,N_14123);
nand U16598 (N_16598,N_14534,N_14002);
or U16599 (N_16599,N_14154,N_14845);
nor U16600 (N_16600,N_14257,N_14908);
xnor U16601 (N_16601,N_15758,N_14849);
or U16602 (N_16602,N_15105,N_14128);
or U16603 (N_16603,N_14351,N_14788);
and U16604 (N_16604,N_15183,N_15929);
and U16605 (N_16605,N_14100,N_14967);
nand U16606 (N_16606,N_14237,N_15512);
and U16607 (N_16607,N_15971,N_14659);
nor U16608 (N_16608,N_14581,N_14415);
or U16609 (N_16609,N_15521,N_15219);
and U16610 (N_16610,N_15565,N_14059);
nor U16611 (N_16611,N_14494,N_15883);
and U16612 (N_16612,N_15734,N_14732);
xnor U16613 (N_16613,N_14956,N_14290);
xnor U16614 (N_16614,N_15495,N_15998);
and U16615 (N_16615,N_15379,N_14427);
xor U16616 (N_16616,N_14843,N_14032);
and U16617 (N_16617,N_14121,N_15545);
and U16618 (N_16618,N_14965,N_15013);
nand U16619 (N_16619,N_15682,N_15917);
nor U16620 (N_16620,N_15856,N_15328);
nand U16621 (N_16621,N_14175,N_15295);
or U16622 (N_16622,N_15763,N_14223);
or U16623 (N_16623,N_15266,N_15028);
nand U16624 (N_16624,N_14650,N_14990);
xor U16625 (N_16625,N_14631,N_15072);
nand U16626 (N_16626,N_14695,N_14681);
nand U16627 (N_16627,N_15823,N_15873);
xnor U16628 (N_16628,N_15879,N_14977);
xnor U16629 (N_16629,N_14125,N_15237);
nor U16630 (N_16630,N_14947,N_15175);
or U16631 (N_16631,N_15748,N_14758);
or U16632 (N_16632,N_15313,N_14667);
xnor U16633 (N_16633,N_14433,N_14706);
or U16634 (N_16634,N_14325,N_15440);
nand U16635 (N_16635,N_15481,N_15716);
nor U16636 (N_16636,N_15926,N_15333);
nor U16637 (N_16637,N_15552,N_14303);
xor U16638 (N_16638,N_14942,N_14113);
nand U16639 (N_16639,N_14711,N_15144);
or U16640 (N_16640,N_14789,N_15938);
xor U16641 (N_16641,N_14613,N_14572);
nor U16642 (N_16642,N_14337,N_14255);
xor U16643 (N_16643,N_14305,N_14160);
and U16644 (N_16644,N_15290,N_15843);
or U16645 (N_16645,N_15089,N_15888);
or U16646 (N_16646,N_15446,N_14355);
or U16647 (N_16647,N_15916,N_15450);
or U16648 (N_16648,N_14626,N_15812);
xnor U16649 (N_16649,N_15332,N_15940);
xor U16650 (N_16650,N_15968,N_15404);
and U16651 (N_16651,N_15610,N_15937);
xor U16652 (N_16652,N_14519,N_14697);
nand U16653 (N_16653,N_15163,N_14539);
or U16654 (N_16654,N_15191,N_15893);
or U16655 (N_16655,N_14883,N_15668);
xor U16656 (N_16656,N_14637,N_14017);
and U16657 (N_16657,N_14165,N_15517);
nand U16658 (N_16658,N_14412,N_15522);
xnor U16659 (N_16659,N_14655,N_14577);
xnor U16660 (N_16660,N_14431,N_15263);
nor U16661 (N_16661,N_14193,N_15102);
nand U16662 (N_16662,N_14651,N_14428);
xor U16663 (N_16663,N_15039,N_15718);
nor U16664 (N_16664,N_14094,N_15118);
and U16665 (N_16665,N_14551,N_15351);
xnor U16666 (N_16666,N_14748,N_15967);
and U16667 (N_16667,N_14423,N_15794);
or U16668 (N_16668,N_14480,N_15996);
nor U16669 (N_16669,N_14763,N_14670);
nor U16670 (N_16670,N_15499,N_14199);
and U16671 (N_16671,N_15309,N_14629);
xnor U16672 (N_16672,N_14931,N_14816);
or U16673 (N_16673,N_14982,N_15036);
nand U16674 (N_16674,N_15268,N_14678);
nand U16675 (N_16675,N_15831,N_15910);
nand U16676 (N_16676,N_15378,N_14496);
and U16677 (N_16677,N_14019,N_15930);
xor U16678 (N_16678,N_14012,N_15486);
nor U16679 (N_16679,N_14818,N_14484);
xor U16680 (N_16680,N_15214,N_15372);
xnor U16681 (N_16681,N_15315,N_14780);
xor U16682 (N_16682,N_14201,N_14426);
and U16683 (N_16683,N_14593,N_14703);
nand U16684 (N_16684,N_14580,N_15874);
and U16685 (N_16685,N_14679,N_15074);
and U16686 (N_16686,N_14061,N_14589);
nor U16687 (N_16687,N_14504,N_14579);
and U16688 (N_16688,N_14052,N_15958);
or U16689 (N_16689,N_15911,N_14260);
xor U16690 (N_16690,N_15616,N_15014);
nor U16691 (N_16691,N_14870,N_15059);
and U16692 (N_16692,N_14636,N_14913);
or U16693 (N_16693,N_15928,N_15535);
and U16694 (N_16694,N_14486,N_14690);
or U16695 (N_16695,N_15574,N_15948);
and U16696 (N_16696,N_15382,N_14552);
nand U16697 (N_16697,N_14619,N_15177);
nor U16698 (N_16698,N_14323,N_14888);
or U16699 (N_16699,N_15882,N_14730);
nand U16700 (N_16700,N_15950,N_15040);
xnor U16701 (N_16701,N_14270,N_15977);
xor U16702 (N_16702,N_14151,N_15484);
nand U16703 (N_16703,N_14245,N_15401);
nor U16704 (N_16704,N_15809,N_14712);
xor U16705 (N_16705,N_15742,N_14622);
xnor U16706 (N_16706,N_15180,N_15592);
and U16707 (N_16707,N_14316,N_15771);
and U16708 (N_16708,N_14215,N_15297);
nand U16709 (N_16709,N_15766,N_14527);
nor U16710 (N_16710,N_15722,N_15326);
xor U16711 (N_16711,N_15892,N_14135);
xor U16712 (N_16712,N_15273,N_15664);
nor U16713 (N_16713,N_15739,N_15651);
and U16714 (N_16714,N_15190,N_15885);
and U16715 (N_16715,N_14759,N_15465);
or U16716 (N_16716,N_15325,N_15819);
and U16717 (N_16717,N_14770,N_14011);
xor U16718 (N_16718,N_14283,N_14664);
or U16719 (N_16719,N_14991,N_14091);
nor U16720 (N_16720,N_14709,N_14332);
nor U16721 (N_16721,N_15134,N_14687);
and U16722 (N_16722,N_15777,N_14048);
and U16723 (N_16723,N_15523,N_15584);
and U16724 (N_16724,N_15988,N_14153);
nand U16725 (N_16725,N_15321,N_14882);
xnor U16726 (N_16726,N_15797,N_14349);
nand U16727 (N_16727,N_15432,N_14880);
xnor U16728 (N_16728,N_15152,N_15020);
nor U16729 (N_16729,N_15129,N_14615);
or U16730 (N_16730,N_14715,N_14205);
nor U16731 (N_16731,N_15520,N_15989);
and U16732 (N_16732,N_15492,N_14702);
xnor U16733 (N_16733,N_15255,N_15083);
or U16734 (N_16734,N_14737,N_15270);
xnor U16735 (N_16735,N_14807,N_14432);
or U16736 (N_16736,N_15037,N_15232);
nor U16737 (N_16737,N_14301,N_15553);
nor U16738 (N_16738,N_14009,N_14710);
and U16739 (N_16739,N_14140,N_15753);
nor U16740 (N_16740,N_15624,N_14750);
and U16741 (N_16741,N_15868,N_15952);
xor U16742 (N_16742,N_15745,N_14057);
or U16743 (N_16743,N_14233,N_15534);
or U16744 (N_16744,N_15947,N_14138);
and U16745 (N_16745,N_15890,N_14372);
nor U16746 (N_16746,N_14617,N_15846);
nor U16747 (N_16747,N_14036,N_14467);
xnor U16748 (N_16748,N_15049,N_14541);
nand U16749 (N_16749,N_15355,N_15870);
and U16750 (N_16750,N_14159,N_14491);
xor U16751 (N_16751,N_14392,N_15136);
xor U16752 (N_16752,N_14456,N_15130);
and U16753 (N_16753,N_14772,N_14248);
xnor U16754 (N_16754,N_14322,N_14388);
nor U16755 (N_16755,N_14724,N_15767);
or U16756 (N_16756,N_14485,N_15442);
nor U16757 (N_16757,N_15648,N_15806);
nor U16758 (N_16758,N_14229,N_14811);
and U16759 (N_16759,N_15855,N_14628);
and U16760 (N_16760,N_15420,N_15506);
or U16761 (N_16761,N_15135,N_14179);
xor U16762 (N_16762,N_14866,N_15498);
or U16763 (N_16763,N_14963,N_14970);
xnor U16764 (N_16764,N_15583,N_14493);
nor U16765 (N_16765,N_14119,N_15785);
nand U16766 (N_16766,N_15627,N_15344);
or U16767 (N_16767,N_15428,N_15644);
nor U16768 (N_16768,N_14814,N_15525);
nor U16769 (N_16769,N_14371,N_15931);
nand U16770 (N_16770,N_15464,N_15172);
and U16771 (N_16771,N_15213,N_14937);
xnor U16772 (N_16772,N_14417,N_15396);
nor U16773 (N_16773,N_14030,N_14834);
nand U16774 (N_16774,N_14473,N_15334);
nand U16775 (N_16775,N_15222,N_14662);
and U16776 (N_16776,N_14191,N_14949);
xnor U16777 (N_16777,N_14665,N_14187);
nor U16778 (N_16778,N_15600,N_15463);
nor U16779 (N_16779,N_14488,N_14174);
nand U16780 (N_16780,N_14489,N_15719);
xnor U16781 (N_16781,N_14594,N_14777);
nor U16782 (N_16782,N_14842,N_15436);
and U16783 (N_16783,N_15850,N_14522);
nor U16784 (N_16784,N_15113,N_14616);
nand U16785 (N_16785,N_14518,N_15330);
or U16786 (N_16786,N_15661,N_14096);
or U16787 (N_16787,N_15140,N_14981);
or U16788 (N_16788,N_14885,N_14457);
or U16789 (N_16789,N_15852,N_15563);
and U16790 (N_16790,N_15618,N_14003);
xor U16791 (N_16791,N_14810,N_14099);
or U16792 (N_16792,N_15030,N_14738);
nor U16793 (N_16793,N_14535,N_15799);
nand U16794 (N_16794,N_14562,N_14385);
and U16795 (N_16795,N_15611,N_15715);
and U16796 (N_16796,N_15054,N_14861);
xnor U16797 (N_16797,N_15374,N_15867);
xor U16798 (N_16798,N_14723,N_14318);
xor U16799 (N_16799,N_14105,N_15009);
xor U16800 (N_16800,N_14300,N_15069);
and U16801 (N_16801,N_15477,N_15939);
nor U16802 (N_16802,N_14302,N_14420);
or U16803 (N_16803,N_15699,N_14794);
or U16804 (N_16804,N_15899,N_15772);
or U16805 (N_16805,N_14210,N_15108);
xor U16806 (N_16806,N_15080,N_14804);
and U16807 (N_16807,N_14241,N_14557);
and U16808 (N_16808,N_14356,N_14396);
or U16809 (N_16809,N_15212,N_14824);
xnor U16810 (N_16810,N_15593,N_14393);
and U16811 (N_16811,N_14960,N_15132);
nand U16812 (N_16812,N_15005,N_15845);
nand U16813 (N_16813,N_15860,N_14319);
nand U16814 (N_16814,N_15654,N_14877);
xnor U16815 (N_16815,N_15038,N_15550);
and U16816 (N_16816,N_15025,N_14291);
or U16817 (N_16817,N_14471,N_15549);
and U16818 (N_16818,N_15571,N_15519);
and U16819 (N_16819,N_14860,N_15412);
nor U16820 (N_16820,N_15157,N_14549);
nand U16821 (N_16821,N_15607,N_14344);
or U16822 (N_16822,N_15914,N_14053);
xnor U16823 (N_16823,N_15115,N_15004);
and U16824 (N_16824,N_14499,N_15875);
and U16825 (N_16825,N_14909,N_14056);
and U16826 (N_16826,N_14256,N_14354);
nor U16827 (N_16827,N_14958,N_15959);
and U16828 (N_16828,N_15281,N_14043);
nand U16829 (N_16829,N_14630,N_15227);
or U16830 (N_16830,N_15424,N_14625);
or U16831 (N_16831,N_15821,N_15107);
and U16832 (N_16832,N_14051,N_15559);
nor U16833 (N_16833,N_14451,N_14688);
nor U16834 (N_16834,N_15211,N_14097);
nor U16835 (N_16835,N_14802,N_15061);
nand U16836 (N_16836,N_15735,N_15443);
and U16837 (N_16837,N_14481,N_14890);
xnor U16838 (N_16838,N_15101,N_14997);
nand U16839 (N_16839,N_15254,N_15920);
and U16840 (N_16840,N_15392,N_14666);
nor U16841 (N_16841,N_15969,N_14186);
xnor U16842 (N_16842,N_15138,N_14606);
nor U16843 (N_16843,N_15642,N_15278);
nand U16844 (N_16844,N_15570,N_15530);
xnor U16845 (N_16845,N_15786,N_14939);
and U16846 (N_16846,N_14595,N_15017);
xnor U16847 (N_16847,N_15643,N_14920);
nor U16848 (N_16848,N_14529,N_14561);
xnor U16849 (N_16849,N_15635,N_15589);
and U16850 (N_16850,N_15003,N_14115);
nor U16851 (N_16851,N_15293,N_15915);
or U16852 (N_16852,N_15364,N_15536);
xnor U16853 (N_16853,N_14398,N_15905);
and U16854 (N_16854,N_14984,N_14718);
xor U16855 (N_16855,N_14721,N_14216);
and U16856 (N_16856,N_15123,N_15729);
nor U16857 (N_16857,N_14930,N_14124);
nand U16858 (N_16858,N_14959,N_15749);
nand U16859 (N_16859,N_14454,N_15992);
and U16860 (N_16860,N_15458,N_14403);
nand U16861 (N_16861,N_15011,N_14550);
and U16862 (N_16862,N_15762,N_15228);
nor U16863 (N_16863,N_14645,N_14130);
nor U16864 (N_16864,N_15337,N_15421);
nand U16865 (N_16865,N_15907,N_15319);
or U16866 (N_16866,N_14994,N_15239);
or U16867 (N_16867,N_15480,N_15951);
xnor U16868 (N_16868,N_15283,N_15127);
xor U16869 (N_16869,N_14359,N_14647);
nor U16870 (N_16870,N_14196,N_15284);
xor U16871 (N_16871,N_14137,N_14104);
or U16872 (N_16872,N_14016,N_15943);
nor U16873 (N_16873,N_14492,N_15073);
nor U16874 (N_16874,N_14120,N_15750);
nand U16875 (N_16875,N_14476,N_15546);
or U16876 (N_16876,N_15689,N_15189);
nor U16877 (N_16877,N_15375,N_15602);
and U16878 (N_16878,N_14155,N_15296);
xnor U16879 (N_16879,N_14176,N_15551);
nand U16880 (N_16880,N_14067,N_15218);
xnor U16881 (N_16881,N_15015,N_14506);
and U16882 (N_16882,N_14685,N_15737);
xnor U16883 (N_16883,N_15423,N_14407);
or U16884 (N_16884,N_15357,N_15400);
or U16885 (N_16885,N_15543,N_14653);
and U16886 (N_16886,N_14045,N_15582);
and U16887 (N_16887,N_15171,N_15660);
nor U16888 (N_16888,N_15335,N_15031);
nand U16889 (N_16889,N_14320,N_14722);
or U16890 (N_16890,N_14064,N_14209);
or U16891 (N_16891,N_14262,N_14353);
nor U16892 (N_16892,N_15529,N_14771);
xor U16893 (N_16893,N_14177,N_14739);
nor U16894 (N_16894,N_14310,N_14218);
xnor U16895 (N_16895,N_15851,N_15961);
nor U16896 (N_16896,N_14565,N_15023);
or U16897 (N_16897,N_14452,N_15151);
and U16898 (N_16898,N_15488,N_15881);
nor U16899 (N_16899,N_15503,N_14983);
or U16900 (N_16900,N_14110,N_15250);
nor U16901 (N_16901,N_15418,N_15121);
xor U16902 (N_16902,N_15838,N_14973);
xor U16903 (N_16903,N_15271,N_15676);
or U16904 (N_16904,N_15272,N_14449);
nor U16905 (N_16905,N_14464,N_14182);
or U16906 (N_16906,N_14031,N_14296);
and U16907 (N_16907,N_15128,N_14952);
xor U16908 (N_16908,N_14150,N_14936);
nand U16909 (N_16909,N_14863,N_15746);
nand U16910 (N_16910,N_14809,N_14327);
nand U16911 (N_16911,N_14833,N_14516);
or U16912 (N_16912,N_15174,N_14853);
nand U16913 (N_16913,N_14083,N_14265);
xor U16914 (N_16914,N_14822,N_14309);
and U16915 (N_16915,N_15158,N_14033);
nand U16916 (N_16916,N_15430,N_14975);
nand U16917 (N_16917,N_15433,N_15291);
xor U16918 (N_16918,N_15168,N_15655);
xnor U16919 (N_16919,N_14585,N_15764);
and U16920 (N_16920,N_15596,N_15814);
xnor U16921 (N_16921,N_15230,N_14231);
and U16922 (N_16922,N_14957,N_14767);
or U16923 (N_16923,N_14696,N_14796);
and U16924 (N_16924,N_14642,N_14379);
or U16925 (N_16925,N_14221,N_15949);
nor U16926 (N_16926,N_15833,N_15991);
nor U16927 (N_16927,N_15995,N_14801);
nor U16928 (N_16928,N_15055,N_14462);
xnor U16929 (N_16929,N_14267,N_15807);
nor U16930 (N_16930,N_15678,N_14946);
nor U16931 (N_16931,N_15993,N_14227);
or U16932 (N_16932,N_15068,N_14038);
nor U16933 (N_16933,N_15743,N_15304);
or U16934 (N_16934,N_15403,N_14787);
or U16935 (N_16935,N_15787,N_15639);
nand U16936 (N_16936,N_15381,N_14921);
nor U16937 (N_16937,N_14278,N_14839);
or U16938 (N_16938,N_15435,N_15822);
and U16939 (N_16939,N_14588,N_14295);
nor U16940 (N_16940,N_15164,N_15594);
nor U16941 (N_16941,N_15114,N_15759);
xnor U16942 (N_16942,N_14576,N_15125);
xnor U16943 (N_16943,N_14111,N_15497);
or U16944 (N_16944,N_14537,N_15274);
or U16945 (N_16945,N_14365,N_14503);
xnor U16946 (N_16946,N_14389,N_15104);
xnor U16947 (N_16947,N_15305,N_14756);
nor U16948 (N_16948,N_14194,N_14126);
and U16949 (N_16949,N_14297,N_15478);
nand U16950 (N_16950,N_15258,N_14076);
nand U16951 (N_16951,N_14528,N_15671);
nor U16952 (N_16952,N_15780,N_14717);
nand U16953 (N_16953,N_15075,N_15496);
nand U16954 (N_16954,N_14675,N_15908);
and U16955 (N_16955,N_15067,N_15837);
xnor U16956 (N_16956,N_14068,N_15088);
or U16957 (N_16957,N_15099,N_14926);
xor U16958 (N_16958,N_15370,N_15942);
and U16959 (N_16959,N_14235,N_14590);
nand U16960 (N_16960,N_14658,N_15800);
xnor U16961 (N_16961,N_14039,N_14974);
or U16962 (N_16962,N_14656,N_14782);
nor U16963 (N_16963,N_15985,N_15087);
xor U16964 (N_16964,N_14434,N_15980);
nand U16965 (N_16965,N_14592,N_15320);
or U16966 (N_16966,N_14152,N_14614);
nor U16967 (N_16967,N_15120,N_15505);
nand U16968 (N_16968,N_14850,N_15323);
or U16969 (N_16969,N_14644,N_14643);
xnor U16970 (N_16970,N_14775,N_15112);
and U16971 (N_16971,N_14547,N_15590);
and U16972 (N_16972,N_15784,N_15933);
nand U16973 (N_16973,N_15124,N_15706);
xnor U16974 (N_16974,N_14729,N_14373);
or U16975 (N_16975,N_14620,N_15373);
xor U16976 (N_16976,N_14132,N_14966);
xor U16977 (N_16977,N_14745,N_15298);
and U16978 (N_16978,N_15783,N_14762);
nor U16979 (N_16979,N_15825,N_14041);
nand U16980 (N_16980,N_15449,N_14487);
nand U16981 (N_16981,N_15242,N_15407);
nor U16982 (N_16982,N_15427,N_15245);
or U16983 (N_16983,N_14108,N_14753);
or U16984 (N_16984,N_14704,N_14668);
nor U16985 (N_16985,N_14835,N_14253);
or U16986 (N_16986,N_15667,N_14848);
and U16987 (N_16987,N_15986,N_15707);
nor U16988 (N_16988,N_15362,N_15246);
xor U16989 (N_16989,N_15658,N_14079);
nor U16990 (N_16990,N_15527,N_14023);
and U16991 (N_16991,N_14902,N_15052);
or U16992 (N_16992,N_15208,N_15217);
nand U16993 (N_16993,N_14893,N_15491);
xor U16994 (N_16994,N_14370,N_14700);
and U16995 (N_16995,N_14776,N_15866);
nor U16996 (N_16996,N_15526,N_15300);
nor U16997 (N_16997,N_14501,N_14251);
xor U16998 (N_16998,N_14683,N_15810);
and U16999 (N_16999,N_15999,N_14545);
nand U17000 (N_17000,N_15442,N_14707);
nand U17001 (N_17001,N_14235,N_14384);
nor U17002 (N_17002,N_15563,N_14869);
nand U17003 (N_17003,N_14281,N_15682);
xor U17004 (N_17004,N_14588,N_14763);
or U17005 (N_17005,N_14415,N_15836);
xor U17006 (N_17006,N_14950,N_15339);
and U17007 (N_17007,N_15348,N_15519);
and U17008 (N_17008,N_14938,N_14313);
and U17009 (N_17009,N_15641,N_15328);
nand U17010 (N_17010,N_14410,N_14516);
nand U17011 (N_17011,N_15846,N_14919);
nand U17012 (N_17012,N_15860,N_15368);
and U17013 (N_17013,N_14168,N_15061);
or U17014 (N_17014,N_14018,N_15299);
nor U17015 (N_17015,N_15765,N_14933);
xor U17016 (N_17016,N_14081,N_14109);
nor U17017 (N_17017,N_14630,N_14307);
and U17018 (N_17018,N_15282,N_15303);
nor U17019 (N_17019,N_14784,N_14801);
nor U17020 (N_17020,N_15641,N_15939);
or U17021 (N_17021,N_15475,N_15484);
nor U17022 (N_17022,N_14711,N_14605);
nor U17023 (N_17023,N_15658,N_15214);
nor U17024 (N_17024,N_15932,N_14262);
and U17025 (N_17025,N_14646,N_15917);
nor U17026 (N_17026,N_15608,N_14003);
or U17027 (N_17027,N_14745,N_14722);
or U17028 (N_17028,N_15522,N_14216);
and U17029 (N_17029,N_14839,N_14595);
xnor U17030 (N_17030,N_14681,N_14730);
and U17031 (N_17031,N_14519,N_15979);
and U17032 (N_17032,N_15150,N_15216);
xnor U17033 (N_17033,N_14718,N_15399);
nor U17034 (N_17034,N_15160,N_14018);
nand U17035 (N_17035,N_14048,N_14125);
or U17036 (N_17036,N_14958,N_14885);
nor U17037 (N_17037,N_14684,N_14004);
and U17038 (N_17038,N_15588,N_15878);
and U17039 (N_17039,N_15672,N_15586);
nand U17040 (N_17040,N_14708,N_15010);
and U17041 (N_17041,N_15028,N_14612);
or U17042 (N_17042,N_15039,N_15589);
and U17043 (N_17043,N_15976,N_14845);
xnor U17044 (N_17044,N_14318,N_15328);
nor U17045 (N_17045,N_14172,N_14361);
or U17046 (N_17046,N_14622,N_14388);
nor U17047 (N_17047,N_15836,N_14696);
xnor U17048 (N_17048,N_15615,N_15023);
nand U17049 (N_17049,N_15826,N_14677);
and U17050 (N_17050,N_14067,N_14044);
or U17051 (N_17051,N_14955,N_15055);
or U17052 (N_17052,N_14899,N_15272);
nand U17053 (N_17053,N_14881,N_14263);
nand U17054 (N_17054,N_15403,N_15872);
xor U17055 (N_17055,N_14718,N_14708);
nand U17056 (N_17056,N_15382,N_14955);
or U17057 (N_17057,N_14491,N_15088);
xnor U17058 (N_17058,N_15960,N_15151);
nor U17059 (N_17059,N_15331,N_14724);
nor U17060 (N_17060,N_15447,N_15251);
and U17061 (N_17061,N_15937,N_15739);
xor U17062 (N_17062,N_15094,N_15474);
or U17063 (N_17063,N_15835,N_15050);
or U17064 (N_17064,N_15048,N_15887);
and U17065 (N_17065,N_14435,N_14407);
nand U17066 (N_17066,N_14725,N_15266);
nor U17067 (N_17067,N_15729,N_14181);
or U17068 (N_17068,N_15844,N_15788);
and U17069 (N_17069,N_14474,N_15416);
xor U17070 (N_17070,N_15418,N_14764);
and U17071 (N_17071,N_15642,N_14965);
or U17072 (N_17072,N_15250,N_14392);
and U17073 (N_17073,N_15841,N_14457);
or U17074 (N_17074,N_15087,N_14107);
nand U17075 (N_17075,N_14311,N_15151);
and U17076 (N_17076,N_14633,N_15717);
xor U17077 (N_17077,N_15316,N_15726);
or U17078 (N_17078,N_15606,N_15148);
nand U17079 (N_17079,N_15746,N_15890);
nand U17080 (N_17080,N_15286,N_15717);
nor U17081 (N_17081,N_14153,N_14232);
nor U17082 (N_17082,N_15705,N_15258);
xnor U17083 (N_17083,N_14008,N_14469);
xnor U17084 (N_17084,N_15263,N_15159);
xnor U17085 (N_17085,N_14372,N_15539);
xor U17086 (N_17086,N_14130,N_15974);
or U17087 (N_17087,N_14293,N_14363);
and U17088 (N_17088,N_15233,N_14680);
and U17089 (N_17089,N_15741,N_15582);
or U17090 (N_17090,N_14740,N_15678);
xor U17091 (N_17091,N_15995,N_15298);
and U17092 (N_17092,N_14701,N_15228);
nor U17093 (N_17093,N_14962,N_14378);
or U17094 (N_17094,N_15679,N_15445);
and U17095 (N_17095,N_14710,N_15998);
and U17096 (N_17096,N_15466,N_14550);
nand U17097 (N_17097,N_14170,N_15274);
and U17098 (N_17098,N_15679,N_14086);
xor U17099 (N_17099,N_15929,N_15030);
or U17100 (N_17100,N_14996,N_14634);
and U17101 (N_17101,N_14251,N_15140);
xnor U17102 (N_17102,N_14416,N_15933);
xnor U17103 (N_17103,N_14124,N_15875);
nor U17104 (N_17104,N_15333,N_14333);
nand U17105 (N_17105,N_14729,N_15442);
xor U17106 (N_17106,N_14396,N_15312);
nor U17107 (N_17107,N_14759,N_14225);
xnor U17108 (N_17108,N_15512,N_14856);
nor U17109 (N_17109,N_15951,N_15025);
nand U17110 (N_17110,N_14017,N_15402);
and U17111 (N_17111,N_15903,N_15004);
nand U17112 (N_17112,N_15108,N_14216);
or U17113 (N_17113,N_14317,N_15402);
xnor U17114 (N_17114,N_14621,N_15158);
nor U17115 (N_17115,N_15383,N_14942);
xnor U17116 (N_17116,N_15139,N_15158);
nand U17117 (N_17117,N_14085,N_14115);
xor U17118 (N_17118,N_14177,N_15727);
nand U17119 (N_17119,N_15115,N_14790);
nand U17120 (N_17120,N_15173,N_14172);
or U17121 (N_17121,N_15205,N_15766);
or U17122 (N_17122,N_15508,N_14254);
nand U17123 (N_17123,N_14579,N_14099);
or U17124 (N_17124,N_14446,N_15853);
xnor U17125 (N_17125,N_15167,N_14033);
xor U17126 (N_17126,N_15695,N_14364);
xnor U17127 (N_17127,N_14483,N_14764);
and U17128 (N_17128,N_15842,N_14376);
nand U17129 (N_17129,N_14118,N_14922);
and U17130 (N_17130,N_15080,N_14665);
nor U17131 (N_17131,N_14587,N_15404);
xnor U17132 (N_17132,N_14485,N_14277);
nor U17133 (N_17133,N_15019,N_14884);
nand U17134 (N_17134,N_14455,N_14965);
nor U17135 (N_17135,N_15874,N_14747);
nand U17136 (N_17136,N_15511,N_14793);
nand U17137 (N_17137,N_15604,N_14828);
nand U17138 (N_17138,N_14963,N_15328);
nand U17139 (N_17139,N_15259,N_15281);
nand U17140 (N_17140,N_14615,N_14107);
and U17141 (N_17141,N_15923,N_15506);
or U17142 (N_17142,N_15903,N_14421);
and U17143 (N_17143,N_15941,N_15074);
or U17144 (N_17144,N_14983,N_14142);
or U17145 (N_17145,N_14928,N_14684);
xnor U17146 (N_17146,N_15126,N_15470);
and U17147 (N_17147,N_15423,N_15466);
nand U17148 (N_17148,N_14494,N_15382);
nand U17149 (N_17149,N_15078,N_15643);
and U17150 (N_17150,N_14024,N_15515);
and U17151 (N_17151,N_15997,N_14627);
nor U17152 (N_17152,N_14231,N_15002);
xnor U17153 (N_17153,N_15937,N_15086);
xnor U17154 (N_17154,N_14245,N_15711);
and U17155 (N_17155,N_15910,N_14597);
xnor U17156 (N_17156,N_15340,N_14065);
and U17157 (N_17157,N_15498,N_14648);
and U17158 (N_17158,N_15556,N_15977);
or U17159 (N_17159,N_15388,N_14125);
nand U17160 (N_17160,N_14467,N_15909);
or U17161 (N_17161,N_14948,N_15343);
nor U17162 (N_17162,N_14021,N_14862);
or U17163 (N_17163,N_15542,N_15454);
or U17164 (N_17164,N_14634,N_14204);
or U17165 (N_17165,N_14773,N_15848);
nor U17166 (N_17166,N_14155,N_14182);
nand U17167 (N_17167,N_15737,N_14590);
nor U17168 (N_17168,N_14558,N_14462);
and U17169 (N_17169,N_15991,N_15434);
or U17170 (N_17170,N_14591,N_14703);
nand U17171 (N_17171,N_14194,N_15343);
nand U17172 (N_17172,N_15353,N_14181);
and U17173 (N_17173,N_14363,N_14114);
and U17174 (N_17174,N_14549,N_15748);
xnor U17175 (N_17175,N_14897,N_15273);
or U17176 (N_17176,N_14709,N_15118);
nand U17177 (N_17177,N_15501,N_15864);
or U17178 (N_17178,N_15375,N_15381);
nand U17179 (N_17179,N_14944,N_15351);
xnor U17180 (N_17180,N_14857,N_15501);
nor U17181 (N_17181,N_15545,N_14524);
nor U17182 (N_17182,N_14864,N_14211);
or U17183 (N_17183,N_14041,N_15953);
xnor U17184 (N_17184,N_14859,N_14484);
nand U17185 (N_17185,N_14489,N_15189);
nand U17186 (N_17186,N_15753,N_14600);
xor U17187 (N_17187,N_15854,N_14213);
xnor U17188 (N_17188,N_14308,N_14223);
xnor U17189 (N_17189,N_14145,N_15112);
or U17190 (N_17190,N_14532,N_14679);
and U17191 (N_17191,N_15225,N_15417);
nand U17192 (N_17192,N_14767,N_14766);
nor U17193 (N_17193,N_15665,N_15418);
nand U17194 (N_17194,N_14477,N_14999);
nor U17195 (N_17195,N_14144,N_15800);
xnor U17196 (N_17196,N_14443,N_14256);
or U17197 (N_17197,N_14803,N_14127);
nand U17198 (N_17198,N_14599,N_14070);
nor U17199 (N_17199,N_15322,N_14938);
and U17200 (N_17200,N_15447,N_14428);
or U17201 (N_17201,N_15986,N_15886);
nand U17202 (N_17202,N_15872,N_15803);
or U17203 (N_17203,N_14477,N_15955);
nand U17204 (N_17204,N_14340,N_15901);
nor U17205 (N_17205,N_14919,N_15333);
and U17206 (N_17206,N_15780,N_14068);
xnor U17207 (N_17207,N_15192,N_14543);
and U17208 (N_17208,N_14475,N_14698);
or U17209 (N_17209,N_15268,N_14142);
nand U17210 (N_17210,N_14283,N_14730);
nand U17211 (N_17211,N_15433,N_15747);
and U17212 (N_17212,N_15775,N_15652);
nand U17213 (N_17213,N_15837,N_14763);
nand U17214 (N_17214,N_14862,N_15050);
and U17215 (N_17215,N_14989,N_14940);
and U17216 (N_17216,N_15289,N_15318);
xor U17217 (N_17217,N_14140,N_15399);
and U17218 (N_17218,N_14385,N_14604);
nand U17219 (N_17219,N_15520,N_15702);
or U17220 (N_17220,N_15242,N_14653);
xor U17221 (N_17221,N_14971,N_14103);
xnor U17222 (N_17222,N_15620,N_14557);
or U17223 (N_17223,N_14504,N_14152);
or U17224 (N_17224,N_15911,N_15407);
xor U17225 (N_17225,N_15955,N_15173);
nand U17226 (N_17226,N_15574,N_14364);
or U17227 (N_17227,N_15289,N_15507);
xnor U17228 (N_17228,N_15979,N_14124);
nor U17229 (N_17229,N_14435,N_15095);
and U17230 (N_17230,N_15650,N_15147);
or U17231 (N_17231,N_15215,N_15556);
xor U17232 (N_17232,N_15192,N_15076);
xor U17233 (N_17233,N_14239,N_15454);
or U17234 (N_17234,N_14826,N_14500);
xnor U17235 (N_17235,N_14619,N_14505);
or U17236 (N_17236,N_15011,N_14747);
nand U17237 (N_17237,N_15805,N_14997);
and U17238 (N_17238,N_15805,N_14062);
and U17239 (N_17239,N_14115,N_14402);
nor U17240 (N_17240,N_14939,N_14597);
and U17241 (N_17241,N_14790,N_15220);
nand U17242 (N_17242,N_14945,N_14828);
and U17243 (N_17243,N_14532,N_14588);
nand U17244 (N_17244,N_15968,N_14277);
and U17245 (N_17245,N_14090,N_15194);
nor U17246 (N_17246,N_14722,N_14086);
xor U17247 (N_17247,N_15135,N_14003);
nor U17248 (N_17248,N_14012,N_15574);
nand U17249 (N_17249,N_14266,N_14196);
nand U17250 (N_17250,N_14719,N_15906);
nand U17251 (N_17251,N_14123,N_15037);
and U17252 (N_17252,N_15202,N_15831);
or U17253 (N_17253,N_15674,N_14355);
or U17254 (N_17254,N_15104,N_15911);
nor U17255 (N_17255,N_15518,N_15321);
xnor U17256 (N_17256,N_15487,N_15301);
xor U17257 (N_17257,N_15446,N_15561);
or U17258 (N_17258,N_14309,N_14239);
nand U17259 (N_17259,N_15515,N_14846);
or U17260 (N_17260,N_15150,N_15894);
or U17261 (N_17261,N_15617,N_15670);
nand U17262 (N_17262,N_15336,N_14396);
nor U17263 (N_17263,N_14332,N_15886);
xor U17264 (N_17264,N_14079,N_15669);
xnor U17265 (N_17265,N_15982,N_15520);
nand U17266 (N_17266,N_15988,N_15718);
and U17267 (N_17267,N_14042,N_14850);
or U17268 (N_17268,N_15481,N_14063);
xor U17269 (N_17269,N_15344,N_14002);
nor U17270 (N_17270,N_15390,N_15979);
xor U17271 (N_17271,N_15319,N_14822);
nor U17272 (N_17272,N_14647,N_14242);
and U17273 (N_17273,N_15417,N_15380);
nand U17274 (N_17274,N_15208,N_14775);
nand U17275 (N_17275,N_14791,N_14659);
nor U17276 (N_17276,N_14456,N_14581);
nor U17277 (N_17277,N_15975,N_14896);
and U17278 (N_17278,N_14058,N_15897);
nand U17279 (N_17279,N_14187,N_15750);
nor U17280 (N_17280,N_14127,N_15792);
or U17281 (N_17281,N_14006,N_14749);
nand U17282 (N_17282,N_15621,N_14853);
xor U17283 (N_17283,N_15646,N_15419);
or U17284 (N_17284,N_14974,N_15789);
nor U17285 (N_17285,N_15400,N_15653);
nor U17286 (N_17286,N_15324,N_14296);
nand U17287 (N_17287,N_14256,N_15977);
and U17288 (N_17288,N_14298,N_14066);
nand U17289 (N_17289,N_15855,N_15570);
xor U17290 (N_17290,N_14762,N_14949);
xor U17291 (N_17291,N_14365,N_15966);
nor U17292 (N_17292,N_15841,N_14014);
nand U17293 (N_17293,N_15916,N_14967);
nor U17294 (N_17294,N_14708,N_14201);
nand U17295 (N_17295,N_14905,N_15054);
nand U17296 (N_17296,N_14852,N_14659);
nand U17297 (N_17297,N_14395,N_14408);
nor U17298 (N_17298,N_14842,N_14548);
xor U17299 (N_17299,N_15919,N_14256);
nand U17300 (N_17300,N_15496,N_15925);
or U17301 (N_17301,N_14708,N_15909);
or U17302 (N_17302,N_14813,N_14935);
nor U17303 (N_17303,N_14989,N_15177);
nand U17304 (N_17304,N_15179,N_14574);
nand U17305 (N_17305,N_14295,N_14107);
nand U17306 (N_17306,N_14281,N_14904);
xor U17307 (N_17307,N_14979,N_15081);
nor U17308 (N_17308,N_15056,N_14494);
nand U17309 (N_17309,N_14446,N_14069);
nor U17310 (N_17310,N_15378,N_15343);
and U17311 (N_17311,N_15883,N_15506);
and U17312 (N_17312,N_15395,N_15217);
nor U17313 (N_17313,N_14727,N_15087);
nor U17314 (N_17314,N_15699,N_14813);
xor U17315 (N_17315,N_15249,N_14631);
nand U17316 (N_17316,N_14155,N_15038);
xnor U17317 (N_17317,N_15123,N_15997);
or U17318 (N_17318,N_15236,N_14242);
and U17319 (N_17319,N_14991,N_14335);
nand U17320 (N_17320,N_15257,N_15927);
and U17321 (N_17321,N_15483,N_15345);
nor U17322 (N_17322,N_15353,N_15403);
xnor U17323 (N_17323,N_15217,N_15450);
and U17324 (N_17324,N_15703,N_15622);
or U17325 (N_17325,N_14239,N_14403);
nor U17326 (N_17326,N_15030,N_14237);
nor U17327 (N_17327,N_14856,N_15473);
or U17328 (N_17328,N_14260,N_14087);
and U17329 (N_17329,N_14752,N_15149);
nand U17330 (N_17330,N_14963,N_15452);
or U17331 (N_17331,N_14453,N_14365);
nor U17332 (N_17332,N_15981,N_15432);
nand U17333 (N_17333,N_15883,N_14234);
nand U17334 (N_17334,N_14239,N_14356);
and U17335 (N_17335,N_15675,N_14181);
nand U17336 (N_17336,N_15168,N_15091);
nor U17337 (N_17337,N_15999,N_14282);
nor U17338 (N_17338,N_14403,N_14809);
nand U17339 (N_17339,N_14273,N_14914);
or U17340 (N_17340,N_15409,N_15610);
nor U17341 (N_17341,N_14131,N_15653);
or U17342 (N_17342,N_15567,N_15327);
nand U17343 (N_17343,N_14722,N_14270);
nand U17344 (N_17344,N_15754,N_14572);
and U17345 (N_17345,N_14669,N_14176);
and U17346 (N_17346,N_14835,N_15199);
xor U17347 (N_17347,N_15339,N_14346);
xnor U17348 (N_17348,N_14243,N_15591);
nand U17349 (N_17349,N_15323,N_14117);
and U17350 (N_17350,N_15370,N_15751);
xnor U17351 (N_17351,N_15739,N_15901);
and U17352 (N_17352,N_14167,N_15799);
or U17353 (N_17353,N_14443,N_14906);
or U17354 (N_17354,N_15408,N_15762);
and U17355 (N_17355,N_15861,N_15785);
and U17356 (N_17356,N_14294,N_15266);
or U17357 (N_17357,N_14658,N_14931);
xnor U17358 (N_17358,N_14556,N_15905);
nand U17359 (N_17359,N_15153,N_15969);
and U17360 (N_17360,N_14289,N_15466);
nand U17361 (N_17361,N_15577,N_15165);
or U17362 (N_17362,N_14067,N_14141);
and U17363 (N_17363,N_14194,N_15721);
xor U17364 (N_17364,N_15585,N_15194);
and U17365 (N_17365,N_15685,N_15420);
or U17366 (N_17366,N_15162,N_15956);
nor U17367 (N_17367,N_15289,N_15922);
nand U17368 (N_17368,N_15701,N_15882);
xor U17369 (N_17369,N_15272,N_15351);
xnor U17370 (N_17370,N_15806,N_15169);
nand U17371 (N_17371,N_15696,N_15054);
nand U17372 (N_17372,N_14536,N_15910);
nor U17373 (N_17373,N_15364,N_15326);
and U17374 (N_17374,N_15024,N_14285);
xnor U17375 (N_17375,N_15989,N_14827);
nand U17376 (N_17376,N_14200,N_14559);
or U17377 (N_17377,N_14852,N_15499);
or U17378 (N_17378,N_14387,N_14571);
xor U17379 (N_17379,N_14505,N_14003);
xnor U17380 (N_17380,N_15226,N_15966);
or U17381 (N_17381,N_15386,N_14943);
nand U17382 (N_17382,N_15652,N_14874);
nand U17383 (N_17383,N_14521,N_14626);
nor U17384 (N_17384,N_15373,N_15019);
nor U17385 (N_17385,N_14753,N_14429);
xnor U17386 (N_17386,N_14366,N_15839);
or U17387 (N_17387,N_15473,N_14463);
nand U17388 (N_17388,N_14534,N_15392);
and U17389 (N_17389,N_14337,N_14682);
nor U17390 (N_17390,N_15324,N_15126);
nand U17391 (N_17391,N_14813,N_14480);
xor U17392 (N_17392,N_14158,N_15584);
nor U17393 (N_17393,N_14183,N_15482);
xnor U17394 (N_17394,N_15701,N_15513);
or U17395 (N_17395,N_14021,N_14658);
and U17396 (N_17396,N_14382,N_15461);
nor U17397 (N_17397,N_15978,N_15004);
nand U17398 (N_17398,N_15220,N_15961);
nor U17399 (N_17399,N_14505,N_14823);
xnor U17400 (N_17400,N_14161,N_14923);
or U17401 (N_17401,N_14314,N_15938);
nor U17402 (N_17402,N_15661,N_15928);
nor U17403 (N_17403,N_15154,N_15298);
xnor U17404 (N_17404,N_14517,N_15680);
and U17405 (N_17405,N_14316,N_15210);
xnor U17406 (N_17406,N_15419,N_15192);
and U17407 (N_17407,N_14965,N_15686);
nor U17408 (N_17408,N_15519,N_15848);
xor U17409 (N_17409,N_15909,N_15914);
or U17410 (N_17410,N_15366,N_14057);
nand U17411 (N_17411,N_14523,N_15913);
or U17412 (N_17412,N_14730,N_14438);
and U17413 (N_17413,N_15417,N_14229);
and U17414 (N_17414,N_15212,N_14577);
or U17415 (N_17415,N_14589,N_14147);
or U17416 (N_17416,N_15934,N_15444);
or U17417 (N_17417,N_15213,N_14835);
xor U17418 (N_17418,N_15919,N_14991);
nor U17419 (N_17419,N_15023,N_14331);
and U17420 (N_17420,N_14115,N_15894);
nor U17421 (N_17421,N_14847,N_15705);
nand U17422 (N_17422,N_15065,N_15742);
nor U17423 (N_17423,N_14135,N_15445);
or U17424 (N_17424,N_14057,N_14059);
nor U17425 (N_17425,N_14417,N_14015);
nand U17426 (N_17426,N_15355,N_15976);
nand U17427 (N_17427,N_14179,N_15492);
or U17428 (N_17428,N_14038,N_14307);
nand U17429 (N_17429,N_15842,N_15953);
or U17430 (N_17430,N_15032,N_14805);
and U17431 (N_17431,N_14774,N_14275);
or U17432 (N_17432,N_15496,N_15243);
and U17433 (N_17433,N_14657,N_14357);
nand U17434 (N_17434,N_15137,N_14246);
xor U17435 (N_17435,N_14228,N_14792);
and U17436 (N_17436,N_14690,N_14926);
and U17437 (N_17437,N_15930,N_15015);
nor U17438 (N_17438,N_15884,N_15980);
or U17439 (N_17439,N_14934,N_15330);
nor U17440 (N_17440,N_15105,N_15773);
or U17441 (N_17441,N_14984,N_14321);
and U17442 (N_17442,N_15912,N_14962);
xor U17443 (N_17443,N_14998,N_15112);
or U17444 (N_17444,N_15613,N_15012);
and U17445 (N_17445,N_15686,N_14852);
or U17446 (N_17446,N_15041,N_14829);
and U17447 (N_17447,N_15788,N_15506);
nor U17448 (N_17448,N_15190,N_15558);
nor U17449 (N_17449,N_15923,N_15576);
xor U17450 (N_17450,N_14838,N_15323);
nor U17451 (N_17451,N_15431,N_15560);
nor U17452 (N_17452,N_15957,N_14362);
xor U17453 (N_17453,N_15925,N_15631);
xor U17454 (N_17454,N_14263,N_14534);
xnor U17455 (N_17455,N_15563,N_14006);
nand U17456 (N_17456,N_15839,N_14960);
nor U17457 (N_17457,N_15673,N_15917);
or U17458 (N_17458,N_15002,N_14360);
nand U17459 (N_17459,N_14159,N_15572);
xor U17460 (N_17460,N_14433,N_15109);
and U17461 (N_17461,N_14725,N_15273);
and U17462 (N_17462,N_14190,N_14933);
nand U17463 (N_17463,N_14715,N_14233);
nand U17464 (N_17464,N_14765,N_15971);
and U17465 (N_17465,N_15449,N_14418);
nand U17466 (N_17466,N_14256,N_14169);
or U17467 (N_17467,N_15707,N_14464);
nor U17468 (N_17468,N_15899,N_14575);
xor U17469 (N_17469,N_15898,N_14022);
xnor U17470 (N_17470,N_14753,N_14308);
xnor U17471 (N_17471,N_15409,N_15300);
xor U17472 (N_17472,N_14291,N_15418);
nand U17473 (N_17473,N_14988,N_14763);
and U17474 (N_17474,N_14407,N_14066);
xnor U17475 (N_17475,N_15190,N_14564);
or U17476 (N_17476,N_14186,N_14784);
and U17477 (N_17477,N_15897,N_15221);
nand U17478 (N_17478,N_14556,N_14919);
or U17479 (N_17479,N_15356,N_15491);
xor U17480 (N_17480,N_15943,N_15989);
and U17481 (N_17481,N_14577,N_15125);
and U17482 (N_17482,N_14230,N_14709);
nor U17483 (N_17483,N_15018,N_14703);
nor U17484 (N_17484,N_15874,N_14159);
or U17485 (N_17485,N_15026,N_14884);
and U17486 (N_17486,N_14979,N_15432);
nand U17487 (N_17487,N_15614,N_14049);
nor U17488 (N_17488,N_14223,N_14764);
nand U17489 (N_17489,N_15884,N_15215);
nor U17490 (N_17490,N_15250,N_15784);
or U17491 (N_17491,N_14434,N_15425);
xnor U17492 (N_17492,N_14606,N_14980);
nor U17493 (N_17493,N_14953,N_14020);
xnor U17494 (N_17494,N_14619,N_15057);
nor U17495 (N_17495,N_14362,N_15656);
or U17496 (N_17496,N_15057,N_14471);
nor U17497 (N_17497,N_15317,N_14284);
xnor U17498 (N_17498,N_14547,N_14960);
or U17499 (N_17499,N_14462,N_15999);
nor U17500 (N_17500,N_14377,N_15127);
nor U17501 (N_17501,N_15232,N_15114);
or U17502 (N_17502,N_15434,N_14964);
xnor U17503 (N_17503,N_14473,N_14093);
nand U17504 (N_17504,N_15889,N_15942);
and U17505 (N_17505,N_14415,N_15933);
or U17506 (N_17506,N_14229,N_15701);
xor U17507 (N_17507,N_14546,N_14665);
nand U17508 (N_17508,N_14978,N_15515);
nor U17509 (N_17509,N_15929,N_14877);
nand U17510 (N_17510,N_15910,N_14946);
and U17511 (N_17511,N_14632,N_14086);
xor U17512 (N_17512,N_14649,N_14506);
and U17513 (N_17513,N_14172,N_14490);
and U17514 (N_17514,N_14476,N_15695);
xnor U17515 (N_17515,N_14077,N_15781);
nand U17516 (N_17516,N_14531,N_14105);
xnor U17517 (N_17517,N_15118,N_15539);
or U17518 (N_17518,N_15607,N_14508);
nand U17519 (N_17519,N_14009,N_14770);
nand U17520 (N_17520,N_14252,N_15302);
and U17521 (N_17521,N_15734,N_14784);
nor U17522 (N_17522,N_15409,N_15905);
xnor U17523 (N_17523,N_14035,N_15693);
nor U17524 (N_17524,N_15543,N_15448);
nand U17525 (N_17525,N_15986,N_15770);
nor U17526 (N_17526,N_15987,N_15749);
or U17527 (N_17527,N_15264,N_15706);
or U17528 (N_17528,N_15507,N_15362);
xnor U17529 (N_17529,N_15039,N_15349);
and U17530 (N_17530,N_15236,N_15383);
xor U17531 (N_17531,N_15085,N_15936);
and U17532 (N_17532,N_14085,N_14088);
xnor U17533 (N_17533,N_15716,N_15996);
nor U17534 (N_17534,N_15394,N_15729);
nor U17535 (N_17535,N_15972,N_15954);
nor U17536 (N_17536,N_15773,N_14347);
and U17537 (N_17537,N_14217,N_14468);
or U17538 (N_17538,N_14274,N_15717);
xnor U17539 (N_17539,N_14415,N_15370);
nand U17540 (N_17540,N_15154,N_14812);
nor U17541 (N_17541,N_14416,N_15395);
xor U17542 (N_17542,N_15195,N_15635);
nor U17543 (N_17543,N_15440,N_14238);
nor U17544 (N_17544,N_15582,N_14769);
nand U17545 (N_17545,N_15984,N_15247);
and U17546 (N_17546,N_14251,N_15886);
nand U17547 (N_17547,N_15670,N_14592);
nor U17548 (N_17548,N_15376,N_15513);
or U17549 (N_17549,N_15155,N_15728);
xor U17550 (N_17550,N_14434,N_14415);
nand U17551 (N_17551,N_15325,N_15835);
nand U17552 (N_17552,N_15952,N_15118);
nor U17553 (N_17553,N_15567,N_15250);
nand U17554 (N_17554,N_15374,N_15736);
and U17555 (N_17555,N_15650,N_14678);
or U17556 (N_17556,N_14251,N_15364);
xnor U17557 (N_17557,N_14479,N_15161);
or U17558 (N_17558,N_15579,N_14004);
nand U17559 (N_17559,N_15719,N_15916);
nor U17560 (N_17560,N_15828,N_14764);
nor U17561 (N_17561,N_14593,N_14813);
or U17562 (N_17562,N_14977,N_14285);
or U17563 (N_17563,N_14552,N_15513);
nand U17564 (N_17564,N_15724,N_14167);
xnor U17565 (N_17565,N_15204,N_15906);
nor U17566 (N_17566,N_15575,N_15133);
and U17567 (N_17567,N_14161,N_15379);
nand U17568 (N_17568,N_15648,N_14941);
nand U17569 (N_17569,N_14173,N_14520);
and U17570 (N_17570,N_15227,N_15383);
or U17571 (N_17571,N_15238,N_14970);
xor U17572 (N_17572,N_15925,N_15973);
nand U17573 (N_17573,N_15390,N_14930);
nand U17574 (N_17574,N_15573,N_15214);
xor U17575 (N_17575,N_14624,N_14312);
nand U17576 (N_17576,N_15227,N_15818);
and U17577 (N_17577,N_15091,N_15892);
and U17578 (N_17578,N_14869,N_15864);
and U17579 (N_17579,N_14652,N_14135);
nand U17580 (N_17580,N_15699,N_14167);
or U17581 (N_17581,N_15898,N_14045);
and U17582 (N_17582,N_15512,N_15824);
xor U17583 (N_17583,N_15944,N_14147);
and U17584 (N_17584,N_14123,N_14108);
nor U17585 (N_17585,N_15113,N_14780);
xnor U17586 (N_17586,N_14877,N_15557);
nor U17587 (N_17587,N_15389,N_15609);
nor U17588 (N_17588,N_14952,N_14156);
nor U17589 (N_17589,N_14782,N_15409);
nand U17590 (N_17590,N_14180,N_15390);
and U17591 (N_17591,N_15011,N_15567);
or U17592 (N_17592,N_15293,N_15150);
nand U17593 (N_17593,N_15448,N_14533);
and U17594 (N_17594,N_15883,N_14635);
nand U17595 (N_17595,N_15427,N_15122);
nor U17596 (N_17596,N_15448,N_14276);
xor U17597 (N_17597,N_14184,N_14473);
nor U17598 (N_17598,N_15452,N_15666);
and U17599 (N_17599,N_14271,N_15086);
xor U17600 (N_17600,N_15744,N_14271);
nor U17601 (N_17601,N_14931,N_15471);
or U17602 (N_17602,N_15054,N_15169);
or U17603 (N_17603,N_15782,N_15689);
or U17604 (N_17604,N_15989,N_14710);
nand U17605 (N_17605,N_15406,N_14572);
or U17606 (N_17606,N_14881,N_14578);
xnor U17607 (N_17607,N_14624,N_14471);
xor U17608 (N_17608,N_14498,N_15775);
nor U17609 (N_17609,N_15265,N_14758);
and U17610 (N_17610,N_15546,N_15772);
or U17611 (N_17611,N_14212,N_14485);
nand U17612 (N_17612,N_14514,N_15456);
or U17613 (N_17613,N_14549,N_14986);
nor U17614 (N_17614,N_15121,N_15758);
or U17615 (N_17615,N_15738,N_14342);
nor U17616 (N_17616,N_15295,N_14212);
nand U17617 (N_17617,N_14878,N_14485);
nand U17618 (N_17618,N_14086,N_15809);
or U17619 (N_17619,N_15532,N_14960);
and U17620 (N_17620,N_14044,N_14855);
or U17621 (N_17621,N_14458,N_15346);
nor U17622 (N_17622,N_15978,N_14370);
xnor U17623 (N_17623,N_14485,N_15016);
and U17624 (N_17624,N_14090,N_14938);
or U17625 (N_17625,N_15841,N_15166);
or U17626 (N_17626,N_15524,N_14063);
nand U17627 (N_17627,N_14028,N_15562);
xor U17628 (N_17628,N_15921,N_14803);
or U17629 (N_17629,N_14101,N_15438);
xor U17630 (N_17630,N_15779,N_14123);
nand U17631 (N_17631,N_14418,N_14810);
xor U17632 (N_17632,N_14146,N_15816);
and U17633 (N_17633,N_14128,N_14632);
nand U17634 (N_17634,N_15012,N_15078);
and U17635 (N_17635,N_14548,N_14396);
xnor U17636 (N_17636,N_15502,N_14217);
nand U17637 (N_17637,N_15090,N_15301);
nor U17638 (N_17638,N_15402,N_14791);
nor U17639 (N_17639,N_14811,N_14074);
nor U17640 (N_17640,N_14245,N_15223);
and U17641 (N_17641,N_15201,N_14180);
xor U17642 (N_17642,N_15115,N_14872);
or U17643 (N_17643,N_14698,N_14074);
and U17644 (N_17644,N_14860,N_14962);
nor U17645 (N_17645,N_15009,N_14364);
nor U17646 (N_17646,N_15804,N_14907);
or U17647 (N_17647,N_14464,N_14105);
xor U17648 (N_17648,N_14506,N_15668);
xnor U17649 (N_17649,N_15990,N_15567);
xnor U17650 (N_17650,N_14627,N_14619);
and U17651 (N_17651,N_14615,N_15886);
or U17652 (N_17652,N_14020,N_14150);
nor U17653 (N_17653,N_14337,N_15667);
nand U17654 (N_17654,N_14564,N_14361);
or U17655 (N_17655,N_14574,N_14227);
nand U17656 (N_17656,N_15759,N_14018);
nand U17657 (N_17657,N_15949,N_15333);
xor U17658 (N_17658,N_15267,N_14228);
nor U17659 (N_17659,N_15791,N_15564);
or U17660 (N_17660,N_14482,N_14070);
or U17661 (N_17661,N_15115,N_15663);
nand U17662 (N_17662,N_15032,N_15684);
xnor U17663 (N_17663,N_14909,N_14654);
nor U17664 (N_17664,N_15775,N_15865);
xor U17665 (N_17665,N_14724,N_15320);
or U17666 (N_17666,N_14384,N_14255);
or U17667 (N_17667,N_15653,N_14342);
and U17668 (N_17668,N_15898,N_14347);
and U17669 (N_17669,N_14766,N_14768);
or U17670 (N_17670,N_14528,N_15910);
and U17671 (N_17671,N_15886,N_14943);
or U17672 (N_17672,N_14562,N_15608);
nand U17673 (N_17673,N_14541,N_15451);
or U17674 (N_17674,N_14549,N_14421);
nor U17675 (N_17675,N_14886,N_14297);
and U17676 (N_17676,N_15729,N_14335);
and U17677 (N_17677,N_14398,N_14793);
nor U17678 (N_17678,N_14635,N_15238);
xor U17679 (N_17679,N_15154,N_14572);
nand U17680 (N_17680,N_14387,N_15550);
nand U17681 (N_17681,N_15545,N_14191);
nand U17682 (N_17682,N_14748,N_15844);
and U17683 (N_17683,N_15246,N_15857);
nor U17684 (N_17684,N_14210,N_15265);
nor U17685 (N_17685,N_15547,N_15930);
xnor U17686 (N_17686,N_15019,N_14017);
and U17687 (N_17687,N_15226,N_14962);
nor U17688 (N_17688,N_15665,N_14528);
xor U17689 (N_17689,N_15073,N_15967);
or U17690 (N_17690,N_14377,N_15118);
or U17691 (N_17691,N_15529,N_14947);
and U17692 (N_17692,N_14361,N_15861);
nand U17693 (N_17693,N_15544,N_14059);
or U17694 (N_17694,N_15036,N_15472);
xor U17695 (N_17695,N_15782,N_14032);
nand U17696 (N_17696,N_14253,N_14965);
xor U17697 (N_17697,N_15959,N_15893);
xor U17698 (N_17698,N_15975,N_15917);
nand U17699 (N_17699,N_15640,N_14435);
xnor U17700 (N_17700,N_14108,N_15957);
xor U17701 (N_17701,N_14415,N_14401);
or U17702 (N_17702,N_14032,N_14772);
xor U17703 (N_17703,N_15805,N_14454);
xnor U17704 (N_17704,N_15618,N_15325);
xor U17705 (N_17705,N_15603,N_15863);
nand U17706 (N_17706,N_15949,N_14469);
nor U17707 (N_17707,N_15775,N_14853);
or U17708 (N_17708,N_14571,N_14493);
xnor U17709 (N_17709,N_14743,N_15787);
nor U17710 (N_17710,N_15569,N_15313);
nand U17711 (N_17711,N_14473,N_15842);
and U17712 (N_17712,N_14790,N_15995);
nand U17713 (N_17713,N_14908,N_14535);
nand U17714 (N_17714,N_14650,N_14410);
and U17715 (N_17715,N_15244,N_14383);
nand U17716 (N_17716,N_14710,N_14068);
xnor U17717 (N_17717,N_14666,N_15650);
nor U17718 (N_17718,N_14923,N_15813);
and U17719 (N_17719,N_15026,N_15984);
or U17720 (N_17720,N_14787,N_14751);
xor U17721 (N_17721,N_14789,N_14769);
and U17722 (N_17722,N_14300,N_15631);
nand U17723 (N_17723,N_15060,N_15500);
nor U17724 (N_17724,N_15420,N_15322);
nand U17725 (N_17725,N_14840,N_15812);
nand U17726 (N_17726,N_14127,N_15677);
or U17727 (N_17727,N_14267,N_15056);
xnor U17728 (N_17728,N_14713,N_15020);
nor U17729 (N_17729,N_14150,N_14054);
or U17730 (N_17730,N_14959,N_15044);
or U17731 (N_17731,N_15882,N_15694);
or U17732 (N_17732,N_15473,N_15132);
xor U17733 (N_17733,N_14187,N_15627);
xnor U17734 (N_17734,N_14897,N_15195);
and U17735 (N_17735,N_15906,N_14816);
or U17736 (N_17736,N_15572,N_14122);
nand U17737 (N_17737,N_15530,N_14994);
and U17738 (N_17738,N_15181,N_15865);
or U17739 (N_17739,N_15518,N_15196);
xnor U17740 (N_17740,N_14054,N_14181);
and U17741 (N_17741,N_14517,N_14658);
nor U17742 (N_17742,N_14747,N_14710);
and U17743 (N_17743,N_15818,N_14207);
and U17744 (N_17744,N_15577,N_14966);
or U17745 (N_17745,N_14071,N_14730);
and U17746 (N_17746,N_14090,N_14625);
and U17747 (N_17747,N_14715,N_14681);
xnor U17748 (N_17748,N_15195,N_15498);
or U17749 (N_17749,N_15020,N_14026);
and U17750 (N_17750,N_14650,N_14982);
nor U17751 (N_17751,N_14032,N_15048);
and U17752 (N_17752,N_15540,N_15971);
xor U17753 (N_17753,N_14052,N_14321);
or U17754 (N_17754,N_15239,N_14135);
and U17755 (N_17755,N_15999,N_15644);
nand U17756 (N_17756,N_14454,N_14117);
xnor U17757 (N_17757,N_15916,N_15798);
xnor U17758 (N_17758,N_14188,N_15907);
nor U17759 (N_17759,N_15876,N_14316);
nor U17760 (N_17760,N_14039,N_15977);
xnor U17761 (N_17761,N_15817,N_14223);
nand U17762 (N_17762,N_15617,N_14468);
and U17763 (N_17763,N_14192,N_14945);
xor U17764 (N_17764,N_14754,N_15626);
xnor U17765 (N_17765,N_14967,N_15156);
and U17766 (N_17766,N_15836,N_14048);
or U17767 (N_17767,N_15147,N_15179);
nand U17768 (N_17768,N_14686,N_15495);
nor U17769 (N_17769,N_14836,N_14464);
or U17770 (N_17770,N_14495,N_14064);
or U17771 (N_17771,N_15498,N_15124);
and U17772 (N_17772,N_14560,N_14220);
nor U17773 (N_17773,N_14070,N_14870);
xnor U17774 (N_17774,N_15040,N_15570);
or U17775 (N_17775,N_14219,N_14606);
nand U17776 (N_17776,N_15807,N_15073);
nor U17777 (N_17777,N_14784,N_14726);
xnor U17778 (N_17778,N_14440,N_15366);
xor U17779 (N_17779,N_14365,N_15817);
xnor U17780 (N_17780,N_14193,N_15663);
and U17781 (N_17781,N_14795,N_14288);
xor U17782 (N_17782,N_15727,N_15200);
and U17783 (N_17783,N_14339,N_15157);
nor U17784 (N_17784,N_14053,N_14264);
or U17785 (N_17785,N_14169,N_14368);
xor U17786 (N_17786,N_15639,N_15421);
xnor U17787 (N_17787,N_14387,N_14599);
xor U17788 (N_17788,N_15847,N_14788);
nand U17789 (N_17789,N_15382,N_15644);
or U17790 (N_17790,N_14715,N_15024);
nand U17791 (N_17791,N_15774,N_14536);
and U17792 (N_17792,N_15653,N_14550);
and U17793 (N_17793,N_15216,N_15438);
and U17794 (N_17794,N_14416,N_15719);
nand U17795 (N_17795,N_14779,N_15774);
or U17796 (N_17796,N_15228,N_14380);
or U17797 (N_17797,N_15461,N_15965);
and U17798 (N_17798,N_15567,N_14386);
or U17799 (N_17799,N_15107,N_14487);
nand U17800 (N_17800,N_14855,N_14120);
and U17801 (N_17801,N_15278,N_15157);
and U17802 (N_17802,N_14786,N_15608);
xor U17803 (N_17803,N_14123,N_14242);
and U17804 (N_17804,N_14513,N_14595);
xnor U17805 (N_17805,N_14354,N_14592);
nor U17806 (N_17806,N_14061,N_14232);
nand U17807 (N_17807,N_14486,N_14811);
xnor U17808 (N_17808,N_15089,N_15068);
nor U17809 (N_17809,N_14854,N_15985);
nor U17810 (N_17810,N_14261,N_15973);
and U17811 (N_17811,N_14705,N_14266);
nor U17812 (N_17812,N_14050,N_15768);
nand U17813 (N_17813,N_14124,N_14879);
nand U17814 (N_17814,N_14193,N_14469);
or U17815 (N_17815,N_15024,N_15669);
or U17816 (N_17816,N_14037,N_14256);
or U17817 (N_17817,N_15491,N_14491);
and U17818 (N_17818,N_14415,N_14685);
or U17819 (N_17819,N_15376,N_15810);
nand U17820 (N_17820,N_15323,N_15784);
and U17821 (N_17821,N_15119,N_15254);
xor U17822 (N_17822,N_14145,N_15343);
and U17823 (N_17823,N_14071,N_15505);
and U17824 (N_17824,N_15038,N_15668);
or U17825 (N_17825,N_15672,N_14996);
nand U17826 (N_17826,N_15626,N_15336);
and U17827 (N_17827,N_15123,N_14960);
or U17828 (N_17828,N_14856,N_14651);
nor U17829 (N_17829,N_14887,N_15639);
nor U17830 (N_17830,N_14502,N_14541);
nor U17831 (N_17831,N_15090,N_15001);
or U17832 (N_17832,N_15738,N_14119);
xnor U17833 (N_17833,N_14299,N_14073);
or U17834 (N_17834,N_14593,N_14581);
or U17835 (N_17835,N_14618,N_14139);
nor U17836 (N_17836,N_15170,N_15826);
nand U17837 (N_17837,N_15091,N_15496);
nand U17838 (N_17838,N_14415,N_15746);
xor U17839 (N_17839,N_15255,N_15780);
nand U17840 (N_17840,N_15599,N_14450);
nand U17841 (N_17841,N_14582,N_14979);
xnor U17842 (N_17842,N_14099,N_15748);
xor U17843 (N_17843,N_15734,N_15433);
nor U17844 (N_17844,N_14765,N_14364);
xor U17845 (N_17845,N_15318,N_15166);
xor U17846 (N_17846,N_15269,N_15905);
xnor U17847 (N_17847,N_15160,N_15320);
or U17848 (N_17848,N_15475,N_15894);
xnor U17849 (N_17849,N_15232,N_15253);
or U17850 (N_17850,N_14204,N_14102);
xor U17851 (N_17851,N_14654,N_14353);
nand U17852 (N_17852,N_14372,N_14419);
nand U17853 (N_17853,N_15576,N_15616);
and U17854 (N_17854,N_14457,N_14514);
xor U17855 (N_17855,N_15390,N_14953);
nand U17856 (N_17856,N_14465,N_15750);
and U17857 (N_17857,N_15538,N_14549);
xnor U17858 (N_17858,N_15505,N_15818);
nand U17859 (N_17859,N_15820,N_15330);
and U17860 (N_17860,N_15695,N_14204);
and U17861 (N_17861,N_14561,N_15186);
xor U17862 (N_17862,N_14661,N_15171);
and U17863 (N_17863,N_14051,N_15117);
or U17864 (N_17864,N_14071,N_15897);
or U17865 (N_17865,N_15340,N_15785);
and U17866 (N_17866,N_15978,N_14547);
or U17867 (N_17867,N_14957,N_15269);
nor U17868 (N_17868,N_15674,N_14418);
nor U17869 (N_17869,N_15915,N_14329);
nand U17870 (N_17870,N_14818,N_14837);
nor U17871 (N_17871,N_15842,N_14515);
and U17872 (N_17872,N_14108,N_15414);
or U17873 (N_17873,N_14296,N_14413);
or U17874 (N_17874,N_15387,N_15650);
nand U17875 (N_17875,N_14169,N_15049);
or U17876 (N_17876,N_14501,N_14988);
and U17877 (N_17877,N_14394,N_15560);
and U17878 (N_17878,N_15818,N_15604);
or U17879 (N_17879,N_14268,N_14521);
nor U17880 (N_17880,N_15985,N_15980);
nor U17881 (N_17881,N_14716,N_15400);
xor U17882 (N_17882,N_15910,N_14686);
or U17883 (N_17883,N_15502,N_15040);
nor U17884 (N_17884,N_14694,N_14828);
xnor U17885 (N_17885,N_15402,N_14878);
and U17886 (N_17886,N_14520,N_15066);
or U17887 (N_17887,N_15674,N_14664);
nor U17888 (N_17888,N_14423,N_14890);
nor U17889 (N_17889,N_15091,N_14552);
nand U17890 (N_17890,N_14944,N_14886);
or U17891 (N_17891,N_14225,N_14431);
nand U17892 (N_17892,N_15987,N_14906);
or U17893 (N_17893,N_15161,N_15223);
nand U17894 (N_17894,N_15811,N_14298);
and U17895 (N_17895,N_14612,N_14518);
and U17896 (N_17896,N_15123,N_15017);
nand U17897 (N_17897,N_14896,N_15693);
or U17898 (N_17898,N_14796,N_15136);
nand U17899 (N_17899,N_15707,N_15098);
and U17900 (N_17900,N_15199,N_15753);
nand U17901 (N_17901,N_15521,N_14994);
or U17902 (N_17902,N_15801,N_15020);
xnor U17903 (N_17903,N_15180,N_15228);
and U17904 (N_17904,N_14196,N_14106);
xor U17905 (N_17905,N_15201,N_15766);
xor U17906 (N_17906,N_15758,N_14841);
or U17907 (N_17907,N_14991,N_15882);
xnor U17908 (N_17908,N_15329,N_14913);
or U17909 (N_17909,N_14159,N_15662);
and U17910 (N_17910,N_14975,N_15132);
nor U17911 (N_17911,N_14900,N_15558);
or U17912 (N_17912,N_15438,N_14953);
xor U17913 (N_17913,N_15918,N_15682);
or U17914 (N_17914,N_15841,N_15561);
xnor U17915 (N_17915,N_15694,N_15007);
and U17916 (N_17916,N_14861,N_15475);
nand U17917 (N_17917,N_14657,N_15586);
xor U17918 (N_17918,N_14716,N_15448);
nor U17919 (N_17919,N_14692,N_15299);
xnor U17920 (N_17920,N_15267,N_14443);
and U17921 (N_17921,N_14877,N_15676);
or U17922 (N_17922,N_14163,N_14953);
nor U17923 (N_17923,N_15308,N_14885);
nor U17924 (N_17924,N_14140,N_15759);
or U17925 (N_17925,N_14553,N_14192);
nor U17926 (N_17926,N_15440,N_14800);
or U17927 (N_17927,N_14132,N_14001);
xnor U17928 (N_17928,N_15165,N_14064);
xor U17929 (N_17929,N_15042,N_14370);
nor U17930 (N_17930,N_15634,N_14850);
and U17931 (N_17931,N_15197,N_15569);
nand U17932 (N_17932,N_14279,N_14657);
nand U17933 (N_17933,N_15645,N_14175);
xnor U17934 (N_17934,N_14414,N_15956);
nand U17935 (N_17935,N_14254,N_15860);
nand U17936 (N_17936,N_14891,N_14628);
or U17937 (N_17937,N_15252,N_14207);
or U17938 (N_17938,N_14852,N_15996);
xnor U17939 (N_17939,N_14845,N_14079);
or U17940 (N_17940,N_15112,N_14158);
and U17941 (N_17941,N_15737,N_15823);
nor U17942 (N_17942,N_14428,N_15129);
xor U17943 (N_17943,N_14179,N_15122);
nand U17944 (N_17944,N_14213,N_14081);
and U17945 (N_17945,N_14421,N_15519);
nor U17946 (N_17946,N_14897,N_15471);
nor U17947 (N_17947,N_15389,N_15180);
xor U17948 (N_17948,N_14383,N_14913);
nor U17949 (N_17949,N_14310,N_15485);
xnor U17950 (N_17950,N_15513,N_15375);
xnor U17951 (N_17951,N_15937,N_14599);
or U17952 (N_17952,N_14301,N_15381);
xor U17953 (N_17953,N_14021,N_14397);
and U17954 (N_17954,N_14653,N_15013);
nand U17955 (N_17955,N_15162,N_15599);
nand U17956 (N_17956,N_14530,N_14286);
xnor U17957 (N_17957,N_14078,N_15195);
nor U17958 (N_17958,N_14272,N_14785);
nand U17959 (N_17959,N_14300,N_15084);
nor U17960 (N_17960,N_15740,N_14230);
nor U17961 (N_17961,N_15001,N_14703);
and U17962 (N_17962,N_14882,N_15182);
or U17963 (N_17963,N_14656,N_15398);
or U17964 (N_17964,N_14101,N_14150);
or U17965 (N_17965,N_14448,N_14804);
nor U17966 (N_17966,N_14814,N_14741);
xor U17967 (N_17967,N_14833,N_14969);
and U17968 (N_17968,N_15775,N_15093);
nor U17969 (N_17969,N_15437,N_14278);
nor U17970 (N_17970,N_14091,N_15444);
and U17971 (N_17971,N_15711,N_15522);
xnor U17972 (N_17972,N_15473,N_15333);
xnor U17973 (N_17973,N_14583,N_15168);
or U17974 (N_17974,N_15167,N_14280);
xnor U17975 (N_17975,N_15045,N_15771);
xnor U17976 (N_17976,N_15981,N_15099);
xnor U17977 (N_17977,N_14182,N_14989);
and U17978 (N_17978,N_14148,N_15452);
or U17979 (N_17979,N_14770,N_15150);
xnor U17980 (N_17980,N_15839,N_15389);
xnor U17981 (N_17981,N_14012,N_15917);
and U17982 (N_17982,N_15853,N_15774);
nand U17983 (N_17983,N_14829,N_14537);
nand U17984 (N_17984,N_15820,N_15231);
or U17985 (N_17985,N_15199,N_15656);
and U17986 (N_17986,N_15116,N_14698);
nor U17987 (N_17987,N_15250,N_15041);
nor U17988 (N_17988,N_15123,N_14963);
and U17989 (N_17989,N_14953,N_14820);
nor U17990 (N_17990,N_15874,N_15758);
nand U17991 (N_17991,N_15935,N_14080);
xnor U17992 (N_17992,N_15450,N_15340);
xor U17993 (N_17993,N_14448,N_15510);
xnor U17994 (N_17994,N_15847,N_14562);
xor U17995 (N_17995,N_15830,N_15726);
or U17996 (N_17996,N_15557,N_15696);
or U17997 (N_17997,N_14512,N_14131);
or U17998 (N_17998,N_14983,N_14829);
xnor U17999 (N_17999,N_15404,N_14447);
xor U18000 (N_18000,N_16860,N_17786);
nor U18001 (N_18001,N_17554,N_17410);
and U18002 (N_18002,N_16065,N_17220);
nor U18003 (N_18003,N_16851,N_16003);
nand U18004 (N_18004,N_16630,N_16534);
and U18005 (N_18005,N_16089,N_16456);
or U18006 (N_18006,N_16505,N_16041);
xor U18007 (N_18007,N_17474,N_16569);
nor U18008 (N_18008,N_17773,N_16932);
nor U18009 (N_18009,N_16028,N_16220);
or U18010 (N_18010,N_17562,N_17144);
nand U18011 (N_18011,N_16733,N_16146);
xor U18012 (N_18012,N_16381,N_16032);
nand U18013 (N_18013,N_17039,N_16196);
xnor U18014 (N_18014,N_17394,N_16725);
nand U18015 (N_18015,N_17884,N_16378);
or U18016 (N_18016,N_16948,N_17865);
nor U18017 (N_18017,N_17150,N_16424);
xor U18018 (N_18018,N_17119,N_17856);
nor U18019 (N_18019,N_17137,N_17698);
nand U18020 (N_18020,N_16844,N_17518);
nor U18021 (N_18021,N_17836,N_17250);
nand U18022 (N_18022,N_17659,N_16788);
or U18023 (N_18023,N_17519,N_17702);
nor U18024 (N_18024,N_17524,N_16467);
nand U18025 (N_18025,N_16856,N_16596);
and U18026 (N_18026,N_16887,N_16421);
nand U18027 (N_18027,N_17335,N_16077);
or U18028 (N_18028,N_17556,N_16328);
nand U18029 (N_18029,N_16434,N_16473);
or U18030 (N_18030,N_17405,N_16379);
nand U18031 (N_18031,N_16965,N_16585);
xor U18032 (N_18032,N_17569,N_17767);
or U18033 (N_18033,N_16440,N_16064);
and U18034 (N_18034,N_16261,N_17254);
or U18035 (N_18035,N_16121,N_17579);
and U18036 (N_18036,N_17857,N_17322);
or U18037 (N_18037,N_16855,N_17789);
or U18038 (N_18038,N_17074,N_16275);
nand U18039 (N_18039,N_17950,N_17291);
nor U18040 (N_18040,N_16242,N_16773);
nand U18041 (N_18041,N_17872,N_16590);
nor U18042 (N_18042,N_17034,N_17852);
nor U18043 (N_18043,N_17647,N_16971);
or U18044 (N_18044,N_16067,N_16057);
nor U18045 (N_18045,N_17149,N_17957);
xnor U18046 (N_18046,N_16136,N_16869);
xnor U18047 (N_18047,N_16129,N_16076);
xor U18048 (N_18048,N_16222,N_16293);
nand U18049 (N_18049,N_17969,N_17009);
and U18050 (N_18050,N_17365,N_17289);
xnor U18051 (N_18051,N_17192,N_16576);
nor U18052 (N_18052,N_17985,N_17143);
nor U18053 (N_18053,N_16812,N_16289);
nor U18054 (N_18054,N_17833,N_17926);
nor U18055 (N_18055,N_17649,N_17928);
and U18056 (N_18056,N_16472,N_17910);
or U18057 (N_18057,N_17771,N_16124);
nor U18058 (N_18058,N_17333,N_17815);
and U18059 (N_18059,N_17976,N_17453);
nor U18060 (N_18060,N_16911,N_17401);
or U18061 (N_18061,N_17779,N_16995);
nor U18062 (N_18062,N_16853,N_16270);
nor U18063 (N_18063,N_16607,N_17433);
or U18064 (N_18064,N_17099,N_16168);
nand U18065 (N_18065,N_17670,N_17349);
xnor U18066 (N_18066,N_16142,N_17834);
nand U18067 (N_18067,N_16800,N_17613);
or U18068 (N_18068,N_16419,N_16690);
nand U18069 (N_18069,N_16039,N_16563);
and U18070 (N_18070,N_16503,N_16359);
and U18071 (N_18071,N_16046,N_16801);
nor U18072 (N_18072,N_16891,N_16380);
xor U18073 (N_18073,N_16483,N_16075);
nor U18074 (N_18074,N_17196,N_17687);
nor U18075 (N_18075,N_16859,N_16166);
xor U18076 (N_18076,N_17752,N_16970);
or U18077 (N_18077,N_16682,N_16582);
xor U18078 (N_18078,N_16088,N_17310);
and U18079 (N_18079,N_16763,N_17213);
xor U18080 (N_18080,N_16258,N_17078);
and U18081 (N_18081,N_16287,N_17368);
nor U18082 (N_18082,N_17530,N_17995);
or U18083 (N_18083,N_16194,N_16054);
and U18084 (N_18084,N_16882,N_17774);
nand U18085 (N_18085,N_17071,N_17471);
or U18086 (N_18086,N_17768,N_16179);
nand U18087 (N_18087,N_16488,N_16538);
or U18088 (N_18088,N_17100,N_17545);
nand U18089 (N_18089,N_17712,N_16881);
or U18090 (N_18090,N_17998,N_16349);
xnor U18091 (N_18091,N_17124,N_16524);
and U18092 (N_18092,N_16916,N_16464);
nor U18093 (N_18093,N_17205,N_17323);
nand U18094 (N_18094,N_17520,N_17006);
nor U18095 (N_18095,N_16436,N_16414);
and U18096 (N_18096,N_16370,N_16192);
nand U18097 (N_18097,N_17001,N_17364);
and U18098 (N_18098,N_17352,N_16500);
or U18099 (N_18099,N_16539,N_17480);
nand U18100 (N_18100,N_16390,N_16454);
and U18101 (N_18101,N_17302,N_16197);
nor U18102 (N_18102,N_16762,N_17182);
nand U18103 (N_18103,N_16227,N_17876);
or U18104 (N_18104,N_17750,N_16308);
nor U18105 (N_18105,N_17542,N_17044);
and U18106 (N_18106,N_16479,N_16968);
xor U18107 (N_18107,N_16314,N_17790);
xnor U18108 (N_18108,N_16274,N_16363);
and U18109 (N_18109,N_16672,N_16988);
or U18110 (N_18110,N_16727,N_17744);
nor U18111 (N_18111,N_17120,N_16110);
and U18112 (N_18112,N_17499,N_16498);
or U18113 (N_18113,N_16496,N_16409);
nand U18114 (N_18114,N_17369,N_16876);
xor U18115 (N_18115,N_17027,N_17716);
xnor U18116 (N_18116,N_17296,N_16508);
nor U18117 (N_18117,N_17327,N_16953);
nand U18118 (N_18118,N_17076,N_16893);
and U18119 (N_18119,N_17958,N_17746);
nand U18120 (N_18120,N_16748,N_16160);
nand U18121 (N_18121,N_17840,N_17970);
nand U18122 (N_18122,N_17913,N_17724);
nor U18123 (N_18123,N_16779,N_17465);
and U18124 (N_18124,N_16085,N_17458);
and U18125 (N_18125,N_16109,N_16332);
or U18126 (N_18126,N_17088,N_17717);
or U18127 (N_18127,N_17838,N_17235);
or U18128 (N_18128,N_16214,N_16273);
and U18129 (N_18129,N_16907,N_16246);
nand U18130 (N_18130,N_17096,N_16329);
xor U18131 (N_18131,N_17892,N_16566);
or U18132 (N_18132,N_17475,N_16427);
and U18133 (N_18133,N_16969,N_17468);
xnor U18134 (N_18134,N_17018,N_17202);
xor U18135 (N_18135,N_17396,N_16511);
xor U18136 (N_18136,N_17328,N_16551);
xor U18137 (N_18137,N_17125,N_16444);
or U18138 (N_18138,N_17491,N_17282);
nor U18139 (N_18139,N_17563,N_16647);
nand U18140 (N_18140,N_17811,N_17440);
xor U18141 (N_18141,N_17211,N_17986);
xnor U18142 (N_18142,N_17005,N_17741);
xor U18143 (N_18143,N_16260,N_17300);
nand U18144 (N_18144,N_16894,N_16589);
and U18145 (N_18145,N_17206,N_16072);
xnor U18146 (N_18146,N_17760,N_17156);
or U18147 (N_18147,N_16661,N_16778);
nor U18148 (N_18148,N_17821,N_16134);
nand U18149 (N_18149,N_17638,N_17904);
or U18150 (N_18150,N_16803,N_16754);
nor U18151 (N_18151,N_17759,N_16143);
xor U18152 (N_18152,N_17439,N_17230);
and U18153 (N_18153,N_16845,N_16943);
nand U18154 (N_18154,N_16398,N_17690);
or U18155 (N_18155,N_16158,N_17607);
and U18156 (N_18156,N_16297,N_17932);
xor U18157 (N_18157,N_16835,N_17867);
and U18158 (N_18158,N_17146,N_17336);
or U18159 (N_18159,N_16183,N_17377);
or U18160 (N_18160,N_17047,N_17631);
xor U18161 (N_18161,N_17916,N_16412);
and U18162 (N_18162,N_16716,N_16397);
and U18163 (N_18163,N_17123,N_17278);
and U18164 (N_18164,N_16252,N_16862);
nand U18165 (N_18165,N_16857,N_16335);
nor U18166 (N_18166,N_16818,N_16651);
nor U18167 (N_18167,N_16235,N_16700);
nor U18168 (N_18168,N_17829,N_17466);
nor U18169 (N_18169,N_16573,N_16091);
or U18170 (N_18170,N_17981,N_16249);
or U18171 (N_18171,N_17451,N_17595);
xor U18172 (N_18172,N_16055,N_16896);
nor U18173 (N_18173,N_16577,N_16974);
xor U18174 (N_18174,N_16611,N_16317);
nor U18175 (N_18175,N_16755,N_16321);
and U18176 (N_18176,N_17019,N_16086);
nand U18177 (N_18177,N_16164,N_16541);
nand U18178 (N_18178,N_17265,N_17195);
and U18179 (N_18179,N_17705,N_16336);
xor U18180 (N_18180,N_16805,N_17955);
xor U18181 (N_18181,N_17081,N_16912);
xnor U18182 (N_18182,N_17093,N_16777);
nand U18183 (N_18183,N_17589,N_16120);
and U18184 (N_18184,N_17126,N_17184);
nand U18185 (N_18185,N_17267,N_17948);
xnor U18186 (N_18186,N_16375,N_17016);
xor U18187 (N_18187,N_17387,N_17485);
nand U18188 (N_18188,N_16394,N_17279);
or U18189 (N_18189,N_17729,N_17070);
or U18190 (N_18190,N_17669,N_17148);
nor U18191 (N_18191,N_17656,N_16083);
and U18192 (N_18192,N_16504,N_17843);
nor U18193 (N_18193,N_16344,N_17260);
nor U18194 (N_18194,N_16646,N_16090);
nand U18195 (N_18195,N_16059,N_17371);
nand U18196 (N_18196,N_17618,N_16231);
and U18197 (N_18197,N_16338,N_17536);
nor U18198 (N_18198,N_17888,N_17984);
nand U18199 (N_18199,N_16527,N_17809);
or U18200 (N_18200,N_16127,N_17527);
or U18201 (N_18201,N_17747,N_16206);
and U18202 (N_18202,N_16334,N_16309);
nand U18203 (N_18203,N_17403,N_16849);
nor U18204 (N_18204,N_16832,N_17068);
nor U18205 (N_18205,N_16357,N_16914);
xor U18206 (N_18206,N_17544,N_16395);
nand U18207 (N_18207,N_17919,N_16316);
and U18208 (N_18208,N_17543,N_17197);
and U18209 (N_18209,N_16229,N_16765);
nand U18210 (N_18210,N_17325,N_17210);
and U18211 (N_18211,N_17208,N_16518);
and U18212 (N_18212,N_17003,N_17108);
xor U18213 (N_18213,N_16886,N_16996);
xor U18214 (N_18214,N_17469,N_17055);
nor U18215 (N_18215,N_16128,N_17105);
xnor U18216 (N_18216,N_17592,N_16437);
and U18217 (N_18217,N_17341,N_16068);
nor U18218 (N_18218,N_16311,N_16903);
and U18219 (N_18219,N_16707,N_17923);
nor U18220 (N_18220,N_17602,N_16556);
nand U18221 (N_18221,N_16023,N_17868);
nor U18222 (N_18222,N_17306,N_16808);
or U18223 (N_18223,N_17939,N_16792);
or U18224 (N_18224,N_17112,N_17848);
and U18225 (N_18225,N_16787,N_16108);
nor U18226 (N_18226,N_17577,N_17431);
or U18227 (N_18227,N_16485,N_17338);
or U18228 (N_18228,N_17229,N_17882);
or U18229 (N_18229,N_16111,N_16025);
nor U18230 (N_18230,N_16678,N_17813);
nand U18231 (N_18231,N_16071,N_16098);
xor U18232 (N_18232,N_16985,N_17639);
xnor U18233 (N_18233,N_17715,N_17135);
xnor U18234 (N_18234,N_17007,N_17351);
and U18235 (N_18235,N_16705,N_16695);
nor U18236 (N_18236,N_16040,N_17564);
nor U18237 (N_18237,N_17781,N_16899);
or U18238 (N_18238,N_17617,N_17091);
and U18239 (N_18239,N_16366,N_16752);
and U18240 (N_18240,N_17608,N_16213);
nand U18241 (N_18241,N_17029,N_17785);
and U18242 (N_18242,N_17632,N_17812);
xnor U18243 (N_18243,N_16669,N_16720);
or U18244 (N_18244,N_17136,N_17145);
or U18245 (N_18245,N_17477,N_17641);
xnor U18246 (N_18246,N_17929,N_17064);
xnor U18247 (N_18247,N_17329,N_17688);
or U18248 (N_18248,N_17181,N_16081);
or U18249 (N_18249,N_17972,N_17620);
nand U18250 (N_18250,N_16704,N_17011);
xnor U18251 (N_18251,N_17508,N_16509);
nand U18252 (N_18252,N_17997,N_17728);
or U18253 (N_18253,N_16063,N_16847);
or U18254 (N_18254,N_16936,N_17676);
xor U18255 (N_18255,N_16416,N_16313);
or U18256 (N_18256,N_16178,N_16623);
nand U18257 (N_18257,N_17793,N_16941);
nand U18258 (N_18258,N_17594,N_17959);
xnor U18259 (N_18259,N_16187,N_16211);
and U18260 (N_18260,N_16676,N_17452);
and U18261 (N_18261,N_17917,N_16605);
or U18262 (N_18262,N_16614,N_17438);
nand U18263 (N_18263,N_16404,N_16712);
nand U18264 (N_18264,N_17521,N_17069);
xor U18265 (N_18265,N_17622,N_16299);
xor U18266 (N_18266,N_16536,N_17885);
nor U18267 (N_18267,N_16738,N_17286);
nor U18268 (N_18268,N_17416,N_17427);
nor U18269 (N_18269,N_17419,N_17117);
and U18270 (N_18270,N_16680,N_17207);
xnor U18271 (N_18271,N_17274,N_16771);
nor U18272 (N_18272,N_16243,N_16612);
nand U18273 (N_18273,N_17045,N_16692);
nand U18274 (N_18274,N_16986,N_16296);
xnor U18275 (N_18275,N_17931,N_16867);
nor U18276 (N_18276,N_16926,N_17493);
and U18277 (N_18277,N_17719,N_16952);
nand U18278 (N_18278,N_17893,N_17938);
nand U18279 (N_18279,N_17924,N_16544);
or U18280 (N_18280,N_17215,N_17245);
nor U18281 (N_18281,N_17691,N_16162);
and U18282 (N_18282,N_16460,N_16766);
or U18283 (N_18283,N_16245,N_16772);
and U18284 (N_18284,N_17353,N_16056);
nor U18285 (N_18285,N_17386,N_17253);
nor U18286 (N_18286,N_17106,N_17354);
xnor U18287 (N_18287,N_17996,N_16240);
nand U18288 (N_18288,N_16925,N_16864);
xnor U18289 (N_18289,N_16639,N_16342);
nor U18290 (N_18290,N_16422,N_16852);
nand U18291 (N_18291,N_16491,N_16718);
and U18292 (N_18292,N_17337,N_17102);
nor U18293 (N_18293,N_17481,N_16571);
nor U18294 (N_18294,N_17823,N_17324);
and U18295 (N_18295,N_16307,N_17583);
and U18296 (N_18296,N_16392,N_17171);
and U18297 (N_18297,N_16927,N_16880);
nor U18298 (N_18298,N_16224,N_16837);
xor U18299 (N_18299,N_16262,N_17457);
nor U18300 (N_18300,N_17978,N_17512);
or U18301 (N_18301,N_17227,N_17604);
nor U18302 (N_18302,N_17478,N_16199);
or U18303 (N_18303,N_16084,N_17308);
or U18304 (N_18304,N_17566,N_17163);
nand U18305 (N_18305,N_17418,N_17412);
and U18306 (N_18306,N_16685,N_17915);
nor U18307 (N_18307,N_17721,N_17990);
nor U18308 (N_18308,N_17601,N_17361);
nor U18309 (N_18309,N_17678,N_16151);
or U18310 (N_18310,N_17551,N_17083);
xor U18311 (N_18311,N_16592,N_16874);
or U18312 (N_18312,N_16815,N_17444);
xor U18313 (N_18313,N_17129,N_17385);
nor U18314 (N_18314,N_17733,N_16346);
or U18315 (N_18315,N_16185,N_16665);
and U18316 (N_18316,N_17933,N_17303);
nor U18317 (N_18317,N_16070,N_16537);
nand U18318 (N_18318,N_17851,N_16044);
nand U18319 (N_18319,N_16030,N_17487);
xor U18320 (N_18320,N_16784,N_17072);
nor U18321 (N_18321,N_17894,N_17671);
xnor U18322 (N_18322,N_17526,N_16450);
nand U18323 (N_18323,N_16466,N_17186);
nor U18324 (N_18324,N_17307,N_16648);
and U18325 (N_18325,N_17672,N_16946);
nand U18326 (N_18326,N_16931,N_17581);
nand U18327 (N_18327,N_17586,N_16182);
xnor U18328 (N_18328,N_16546,N_16204);
or U18329 (N_18329,N_17248,N_17549);
nor U18330 (N_18330,N_17086,N_16218);
nand U18331 (N_18331,N_16940,N_16497);
and U18332 (N_18332,N_16846,N_16355);
nor U18333 (N_18333,N_16137,N_16999);
nor U18334 (N_18334,N_16833,N_16303);
xor U18335 (N_18335,N_17753,N_16652);
nor U18336 (N_18336,N_16934,N_16561);
nand U18337 (N_18337,N_16283,N_17225);
or U18338 (N_18338,N_17391,N_17379);
nor U18339 (N_18339,N_16734,N_16586);
nor U18340 (N_18340,N_16257,N_17804);
or U18341 (N_18341,N_17905,N_16732);
nor U18342 (N_18342,N_17187,N_16186);
or U18343 (N_18343,N_17918,N_16458);
and U18344 (N_18344,N_16244,N_17402);
or U18345 (N_18345,N_16318,N_17292);
and U18346 (N_18346,N_16002,N_16300);
nand U18347 (N_18347,N_17936,N_17486);
nand U18348 (N_18348,N_17326,N_17898);
nand U18349 (N_18349,N_17050,N_16606);
and U18350 (N_18350,N_16163,N_17151);
nand U18351 (N_18351,N_16722,N_16324);
nand U18352 (N_18352,N_16820,N_17021);
or U18353 (N_18353,N_16209,N_17845);
nand U18354 (N_18354,N_16074,N_17272);
nand U18355 (N_18355,N_17515,N_16601);
nor U18356 (N_18356,N_17121,N_16291);
and U18357 (N_18357,N_17841,N_17194);
nor U18358 (N_18358,N_17020,N_16060);
nand U18359 (N_18359,N_16499,N_17141);
xor U18360 (N_18360,N_17165,N_17965);
and U18361 (N_18361,N_17535,N_17233);
nand U18362 (N_18362,N_17008,N_16470);
and U18363 (N_18363,N_17339,N_17650);
nor U18364 (N_18364,N_16572,N_17190);
or U18365 (N_18365,N_16583,N_16660);
xnor U18366 (N_18366,N_16385,N_17128);
and U18367 (N_18367,N_17805,N_16012);
or U18368 (N_18368,N_17334,N_17413);
nand U18369 (N_18369,N_16810,N_16776);
nor U18370 (N_18370,N_17111,N_17209);
nor U18371 (N_18371,N_17243,N_16489);
xor U18372 (N_18372,N_16451,N_17658);
nor U18373 (N_18373,N_16482,N_16963);
xor U18374 (N_18374,N_16565,N_16521);
or U18375 (N_18375,N_16821,N_16383);
xor U18376 (N_18376,N_16027,N_16447);
nand U18377 (N_18377,N_16957,N_16011);
or U18378 (N_18378,N_16052,N_17052);
and U18379 (N_18379,N_16928,N_16751);
or U18380 (N_18380,N_16868,N_17598);
nor U18381 (N_18381,N_17828,N_17046);
or U18382 (N_18382,N_17152,N_16683);
xor U18383 (N_18383,N_17503,N_17257);
xor U18384 (N_18384,N_17320,N_17643);
xor U18385 (N_18385,N_17830,N_16983);
nor U18386 (N_18386,N_17974,N_17814);
xor U18387 (N_18387,N_17921,N_17153);
xor U18388 (N_18388,N_16465,N_16339);
nor U18389 (N_18389,N_16304,N_17426);
or U18390 (N_18390,N_17674,N_17450);
and U18391 (N_18391,N_16118,N_17802);
and U18392 (N_18392,N_16594,N_17384);
or U18393 (N_18393,N_16510,N_17492);
nor U18394 (N_18394,N_16761,N_16717);
or U18395 (N_18395,N_16939,N_17820);
xnor U18396 (N_18396,N_16062,N_16147);
xnor U18397 (N_18397,N_17345,N_17689);
or U18398 (N_18398,N_16133,N_17599);
nand U18399 (N_18399,N_17695,N_17037);
nor U18400 (N_18400,N_16453,N_16350);
nand U18401 (N_18401,N_17509,N_16205);
and U18402 (N_18402,N_17134,N_17373);
nand U18403 (N_18403,N_16923,N_17222);
and U18404 (N_18404,N_17590,N_16892);
nand U18405 (N_18405,N_16426,N_16955);
nand U18406 (N_18406,N_17550,N_16517);
nand U18407 (N_18407,N_17701,N_17621);
and U18408 (N_18408,N_17999,N_16616);
nor U18409 (N_18409,N_17496,N_16533);
and U18410 (N_18410,N_16740,N_17548);
and U18411 (N_18411,N_16615,N_17014);
or U18412 (N_18412,N_16037,N_17818);
nor U18413 (N_18413,N_16232,N_16320);
nand U18414 (N_18414,N_17428,N_17778);
nor U18415 (N_18415,N_16391,N_16123);
xnor U18416 (N_18416,N_16719,N_16883);
and U18417 (N_18417,N_17682,N_16446);
xnor U18418 (N_18418,N_16687,N_17359);
xnor U18419 (N_18419,N_17501,N_17318);
and U18420 (N_18420,N_16640,N_16557);
or U18421 (N_18421,N_16984,N_16008);
xnor U18422 (N_18422,N_16728,N_16938);
or U18423 (N_18423,N_16066,N_17528);
and U18424 (N_18424,N_16026,N_17538);
xnor U18425 (N_18425,N_17627,N_17367);
xnor U18426 (N_18426,N_16688,N_16139);
and U18427 (N_18427,N_17546,N_17902);
or U18428 (N_18428,N_16530,N_17425);
xnor U18429 (N_18429,N_17640,N_16302);
and U18430 (N_18430,N_16947,N_16170);
and U18431 (N_18431,N_17281,N_16670);
nand U18432 (N_18432,N_17288,N_16420);
nand U18433 (N_18433,N_16325,N_17920);
nor U18434 (N_18434,N_16714,N_16050);
nor U18435 (N_18435,N_17201,N_16140);
xnor U18436 (N_18436,N_17023,N_17662);
xnor U18437 (N_18437,N_17139,N_17858);
xor U18438 (N_18438,N_16267,N_16699);
nand U18439 (N_18439,N_16345,N_17539);
and U18440 (N_18440,N_17988,N_16095);
xor U18441 (N_18441,N_16958,N_17683);
xnor U18442 (N_18442,N_16861,N_16119);
nand U18443 (N_18443,N_17395,N_16905);
or U18444 (N_18444,N_17934,N_17162);
or U18445 (N_18445,N_16587,N_17537);
and U18446 (N_18446,N_17606,N_17226);
nor U18447 (N_18447,N_16884,N_17935);
and U18448 (N_18448,N_16184,N_17945);
nand U18449 (N_18449,N_16389,N_16522);
and U18450 (N_18450,N_16742,N_16295);
nor U18451 (N_18451,N_16047,N_17489);
nor U18452 (N_18452,N_17982,N_17635);
and U18453 (N_18453,N_17525,N_17249);
and U18454 (N_18454,N_17889,N_17827);
and U18455 (N_18455,N_16341,N_17073);
nand U18456 (N_18456,N_17616,N_17456);
nand U18457 (N_18457,N_16992,N_16545);
nor U18458 (N_18458,N_17285,N_17944);
or U18459 (N_18459,N_17553,N_17953);
nand U18460 (N_18460,N_17189,N_16264);
nand U18461 (N_18461,N_16658,N_17490);
xor U18462 (N_18462,N_17284,N_17090);
nor U18463 (N_18463,N_17652,N_17943);
xnor U18464 (N_18464,N_17315,N_16981);
or U18465 (N_18465,N_17404,N_16749);
xnor U18466 (N_18466,N_16212,N_16286);
or U18467 (N_18467,N_17342,N_17449);
nor U18468 (N_18468,N_16276,N_16730);
nand U18469 (N_18469,N_16701,N_17113);
xor U18470 (N_18470,N_16322,N_16966);
or U18471 (N_18471,N_17287,N_17596);
nand U18472 (N_18472,N_17203,N_16092);
or U18473 (N_18473,N_16004,N_16824);
nor U18474 (N_18474,N_16282,N_16410);
nor U18475 (N_18475,N_16455,N_16481);
nand U18476 (N_18476,N_17762,N_16609);
and U18477 (N_18477,N_17178,N_16005);
nor U18478 (N_18478,N_16376,N_16181);
nor U18479 (N_18479,N_16367,N_17173);
nor U18480 (N_18480,N_17199,N_16642);
nor U18481 (N_18481,N_17757,N_16442);
and U18482 (N_18482,N_17247,N_17277);
or U18483 (N_18483,N_16144,N_17314);
xnor U18484 (N_18484,N_16620,N_16711);
and U18485 (N_18485,N_17883,N_17879);
nand U18486 (N_18486,N_17890,N_16809);
nand U18487 (N_18487,N_17435,N_16272);
nor U18488 (N_18488,N_16105,N_16049);
nor U18489 (N_18489,N_17605,N_17010);
nand U18490 (N_18490,N_17684,N_17723);
nor U18491 (N_18491,N_16831,N_16764);
and U18492 (N_18492,N_16841,N_16584);
nand U18493 (N_18493,N_16850,N_17573);
nor U18494 (N_18494,N_16908,N_16369);
nor U18495 (N_18495,N_16333,N_17505);
and U18496 (N_18496,N_17217,N_16666);
and U18497 (N_18497,N_17927,N_17488);
or U18498 (N_18498,N_17507,N_17079);
nor U18499 (N_18499,N_17587,N_16155);
nor U18500 (N_18500,N_16649,N_17855);
or U18501 (N_18501,N_16169,N_16097);
or U18502 (N_18502,N_17735,N_17236);
xnor U18503 (N_18503,N_17792,N_16082);
xor U18504 (N_18504,N_17447,N_17362);
nor U18505 (N_18505,N_16560,N_16625);
and U18506 (N_18506,N_16250,N_16671);
xnor U18507 (N_18507,N_17764,N_17615);
nand U18508 (N_18508,N_17675,N_16753);
nand U18509 (N_18509,N_17644,N_17147);
xor U18510 (N_18510,N_17619,N_17132);
or U18511 (N_18511,N_17956,N_17873);
and U18512 (N_18512,N_17041,N_16053);
nor U18513 (N_18513,N_17624,N_16326);
and U18514 (N_18514,N_16208,N_16290);
and U18515 (N_18515,N_17035,N_17231);
nor U18516 (N_18516,N_17381,N_17738);
nand U18517 (N_18517,N_16698,N_16167);
nor U18518 (N_18518,N_16621,N_17941);
nand U18519 (N_18519,N_16840,N_17399);
nand U18520 (N_18520,N_17628,N_17473);
or U18521 (N_18521,N_17761,N_17441);
or U18522 (N_18522,N_17448,N_16193);
and U18523 (N_18523,N_16469,N_17708);
or U18524 (N_18524,N_17271,N_17633);
nor U18525 (N_18525,N_17370,N_17751);
xnor U18526 (N_18526,N_16207,N_16675);
nand U18527 (N_18527,N_16774,N_17383);
nand U18528 (N_18528,N_17963,N_16474);
nand U18529 (N_18529,N_16663,N_16429);
nand U18530 (N_18530,N_16622,N_16870);
nand U18531 (N_18531,N_16811,N_17321);
nand U18532 (N_18532,N_17565,N_17642);
and U18533 (N_18533,N_16356,N_17214);
and U18534 (N_18534,N_16487,N_16013);
xor U18535 (N_18535,N_16130,N_17040);
and U18536 (N_18536,N_16828,N_16009);
xor U18537 (N_18537,N_16094,N_17740);
and U18538 (N_18538,N_16288,N_16445);
and U18539 (N_18539,N_17022,N_17912);
nand U18540 (N_18540,N_17863,N_16400);
xor U18541 (N_18541,N_16048,N_17500);
nor U18542 (N_18542,N_16608,N_16662);
and U18543 (N_18543,N_16529,N_16371);
xnor U18544 (N_18544,N_16735,N_17028);
xor U18545 (N_18545,N_16478,N_17726);
xnor U18546 (N_18546,N_16782,N_17309);
nor U18547 (N_18547,N_17510,N_16760);
and U18548 (N_18548,N_16960,N_17026);
nand U18549 (N_18549,N_16918,N_16574);
nor U18550 (N_18550,N_17597,N_16523);
nor U18551 (N_18551,N_17609,N_17860);
xnor U18552 (N_18552,N_16348,N_17360);
and U18553 (N_18553,N_16593,N_17311);
xnor U18554 (N_18554,N_17736,N_17555);
and U18555 (N_18555,N_17718,N_17591);
xor U18556 (N_18556,N_17446,N_16816);
xor U18557 (N_18557,N_16921,N_16602);
or U18558 (N_18558,N_17677,N_17299);
nor U18559 (N_18559,N_16343,N_17560);
nor U18560 (N_18560,N_17552,N_16148);
nand U18561 (N_18561,N_17237,N_17193);
and U18562 (N_18562,N_16677,N_16654);
or U18563 (N_18563,N_16531,N_16058);
nor U18564 (N_18564,N_16975,N_16567);
or U18565 (N_18565,N_17694,N_16746);
nor U18566 (N_18566,N_16998,N_16830);
xor U18567 (N_18567,N_16578,N_17907);
nand U18568 (N_18568,N_16659,N_17696);
xor U18569 (N_18569,N_16631,N_17084);
nor U18570 (N_18570,N_16976,N_16433);
xor U18571 (N_18571,N_17363,N_17067);
xnor U18572 (N_18572,N_16189,N_17409);
or U18573 (N_18573,N_16635,N_17380);
or U18574 (N_18574,N_17048,N_16506);
or U18575 (N_18575,N_16156,N_16964);
and U18576 (N_18576,N_16228,N_16829);
and U18577 (N_18577,N_17523,N_17414);
nor U18578 (N_18578,N_17947,N_16396);
nor U18579 (N_18579,N_16744,N_16399);
nor U18580 (N_18580,N_17024,N_16713);
nand U18581 (N_18581,N_16402,N_16361);
nor U18582 (N_18582,N_16736,N_16132);
and U18583 (N_18583,N_17513,N_17664);
and U18584 (N_18584,N_16171,N_16637);
xnor U18585 (N_18585,N_17030,N_16997);
xor U18586 (N_18586,N_16269,N_16248);
nor U18587 (N_18587,N_17937,N_17584);
and U18588 (N_18588,N_17704,N_16930);
nand U18589 (N_18589,N_16900,N_17442);
and U18590 (N_18590,N_17946,N_16978);
xnor U18591 (N_18591,N_17138,N_16785);
xor U18592 (N_18592,N_17842,N_16917);
and U18593 (N_18593,N_16679,N_17588);
nor U18594 (N_18594,N_17470,N_17637);
or U18595 (N_18595,N_17216,N_16579);
xnor U18596 (N_18596,N_16644,N_17517);
nor U18597 (N_18597,N_17476,N_16967);
xor U18598 (N_18598,N_17130,N_16595);
nor U18599 (N_18599,N_16405,N_17133);
nor U18600 (N_18600,N_17940,N_16285);
and U18601 (N_18601,N_17255,N_16842);
or U18602 (N_18602,N_16922,N_16709);
nand U18603 (N_18603,N_16138,N_16558);
nor U18604 (N_18604,N_16268,N_16909);
nor U18605 (N_18605,N_17506,N_17975);
or U18606 (N_18606,N_16520,N_16180);
xor U18607 (N_18607,N_16364,N_16035);
nor U18608 (N_18608,N_16598,N_16775);
nand U18609 (N_18609,N_16668,N_17375);
or U18610 (N_18610,N_16216,N_17317);
and U18611 (N_18611,N_17095,N_17049);
nor U18612 (N_18612,N_16241,N_17808);
or U18613 (N_18613,N_16007,N_17241);
nand U18614 (N_18614,N_17174,N_17796);
or U18615 (N_18615,N_17340,N_17777);
nor U18616 (N_18616,N_16347,N_17654);
or U18617 (N_18617,N_17259,N_16484);
and U18618 (N_18618,N_16016,N_16633);
or U18619 (N_18619,N_17280,N_16036);
or U18620 (N_18620,N_16650,N_17901);
nor U18621 (N_18621,N_17408,N_16238);
or U18622 (N_18622,N_16875,N_16786);
xnor U18623 (N_18623,N_17967,N_17421);
nand U18624 (N_18624,N_17204,N_16327);
or U18625 (N_18625,N_16301,N_17854);
xnor U18626 (N_18626,N_17058,N_17484);
nand U18627 (N_18627,N_16247,N_17784);
or U18628 (N_18628,N_17900,N_16407);
nand U18629 (N_18629,N_16555,N_16234);
nand U18630 (N_18630,N_17713,N_16629);
and U18631 (N_18631,N_17378,N_16315);
nor U18632 (N_18632,N_17077,N_17060);
or U18633 (N_18633,N_17629,N_16106);
or U18634 (N_18634,N_17700,N_16982);
xor U18635 (N_18635,N_16362,N_16459);
nand U18636 (N_18636,N_17033,N_17534);
and U18637 (N_18637,N_17109,N_17803);
and U18638 (N_18638,N_17168,N_16959);
nand U18639 (N_18639,N_17454,N_16490);
and U18640 (N_18640,N_16116,N_17951);
nor U18641 (N_18641,N_17817,N_16358);
or U18642 (N_18642,N_17004,N_17623);
or U18643 (N_18643,N_16721,N_17801);
nor U18644 (N_18644,N_16382,N_16873);
and U18645 (N_18645,N_17732,N_17720);
nand U18646 (N_18646,N_17514,N_17343);
nand U18647 (N_18647,N_17406,N_16933);
xnor U18648 (N_18648,N_17561,N_16929);
and U18649 (N_18649,N_17131,N_16225);
and U18650 (N_18650,N_17874,N_16581);
and U18651 (N_18651,N_16096,N_16159);
or U18652 (N_18652,N_16073,N_17822);
nor U18653 (N_18653,N_16443,N_17063);
nand U18654 (N_18654,N_16475,N_17832);
nor U18655 (N_18655,N_17826,N_16126);
or U18656 (N_18656,N_16502,N_17925);
or U18657 (N_18657,N_17429,N_16408);
and U18658 (N_18658,N_17603,N_16354);
nand U18659 (N_18659,N_16131,N_17107);
xnor U18660 (N_18660,N_17332,N_17392);
nor U18661 (N_18661,N_16463,N_17331);
nand U18662 (N_18662,N_17903,N_17780);
xnor U18663 (N_18663,N_16767,N_16655);
and U18664 (N_18664,N_16337,N_16031);
and U18665 (N_18665,N_16681,N_16991);
or U18666 (N_18666,N_17798,N_17042);
nand U18667 (N_18667,N_17887,N_16256);
nand U18668 (N_18668,N_16980,N_16277);
xor U18669 (N_18669,N_17175,N_17625);
or U18670 (N_18670,N_17422,N_16877);
or U18671 (N_18671,N_17680,N_16854);
and U18672 (N_18672,N_17949,N_16449);
nand U18673 (N_18673,N_17293,N_17166);
xnor U18674 (N_18674,N_16029,N_17870);
xnor U18675 (N_18675,N_17062,N_17961);
or U18676 (N_18676,N_16703,N_16653);
nor U18677 (N_18677,N_17118,N_16069);
and U18678 (N_18678,N_16493,N_17859);
or U18679 (N_18679,N_16312,N_17770);
nor U18680 (N_18680,N_17571,N_17578);
or U18681 (N_18681,N_17612,N_16384);
xor U18682 (N_18682,N_17749,N_17794);
nor U18683 (N_18683,N_16798,N_16330);
nor U18684 (N_18684,N_17661,N_17013);
nand U18685 (N_18685,N_16457,N_16913);
or U18686 (N_18686,N_17731,N_16667);
nand U18687 (N_18687,N_17745,N_16797);
or U18688 (N_18688,N_16950,N_17266);
or U18689 (N_18689,N_17994,N_16254);
nor U18690 (N_18690,N_16554,N_17263);
xor U18691 (N_18691,N_17223,N_16697);
nor U18692 (N_18692,N_16122,N_16769);
xor U18693 (N_18693,N_16514,N_17585);
and U18694 (N_18694,N_16203,N_17455);
and U18695 (N_18695,N_17799,N_16024);
and U18696 (N_18696,N_17319,N_17283);
and U18697 (N_18697,N_17098,N_17769);
or U18698 (N_18698,N_17415,N_16863);
xnor U18699 (N_18699,N_16627,N_17347);
nor U18700 (N_18700,N_16745,N_17835);
nor U18701 (N_18701,N_17568,N_17238);
nor U18702 (N_18702,N_17930,N_17057);
nor U18703 (N_18703,N_16657,N_16271);
and U18704 (N_18704,N_16468,N_17630);
or U18705 (N_18705,N_17906,N_17183);
and U18706 (N_18706,N_17398,N_16417);
nor U18707 (N_18707,N_16154,N_16610);
nor U18708 (N_18708,N_16588,N_16791);
and U18709 (N_18709,N_17663,N_17909);
nand U18710 (N_18710,N_16462,N_17116);
and U18711 (N_18711,N_17031,N_17464);
and U18712 (N_18712,N_16480,N_16942);
xor U18713 (N_18713,N_16726,N_17390);
or U18714 (N_18714,N_16516,N_16141);
and U18715 (N_18715,N_16949,N_16708);
xnor U18716 (N_18716,N_17660,N_16080);
nand U18717 (N_18717,N_17810,N_16051);
xor U18718 (N_18718,N_16872,N_17572);
or U18719 (N_18719,N_16535,N_16888);
and U18720 (N_18720,N_17002,N_17258);
or U18721 (N_18721,N_17097,N_16438);
nand U18722 (N_18722,N_16153,N_17610);
and U18723 (N_18723,N_16802,N_16737);
or U18724 (N_18724,N_17142,N_16353);
and U18725 (N_18725,N_16619,N_17765);
or U18726 (N_18726,N_17877,N_17908);
nand U18727 (N_18727,N_16239,N_16919);
and U18728 (N_18728,N_17012,N_17847);
nand U18729 (N_18729,N_17191,N_17101);
or U18730 (N_18730,N_16897,N_16174);
xnor U18731 (N_18731,N_16042,N_17389);
or U18732 (N_18732,N_17754,N_17025);
nand U18733 (N_18733,N_17157,N_17582);
nand U18734 (N_18734,N_17304,N_17532);
xor U18735 (N_18735,N_17103,N_17968);
and U18736 (N_18736,N_17160,N_16406);
nor U18737 (N_18737,N_16014,N_16340);
or U18738 (N_18738,N_17653,N_16817);
or U18739 (N_18739,N_16360,N_17000);
and U18740 (N_18740,N_17580,N_17198);
nand U18741 (N_18741,N_17417,N_16580);
or U18742 (N_18742,N_16599,N_17611);
and U18743 (N_18743,N_17256,N_17991);
and U18744 (N_18744,N_16177,N_16401);
xor U18745 (N_18745,N_17993,N_16799);
nand U18746 (N_18746,N_17710,N_16994);
nor U18747 (N_18747,N_16298,N_17540);
nor U18748 (N_18748,N_16553,N_17871);
nor U18749 (N_18749,N_16255,N_17697);
and U18750 (N_18750,N_17897,N_16937);
xor U18751 (N_18751,N_16236,N_17158);
nor U18752 (N_18752,N_16306,N_17170);
and U18753 (N_18753,N_17316,N_17053);
nor U18754 (N_18754,N_17758,N_17983);
and U18755 (N_18755,N_16201,N_16838);
nor U18756 (N_18756,N_16781,N_17837);
and U18757 (N_18757,N_17707,N_16706);
nor U18758 (N_18758,N_17397,N_17853);
nor U18759 (N_18759,N_17964,N_17437);
nand U18760 (N_18760,N_17472,N_17734);
or U18761 (N_18761,N_16562,N_16547);
and U18762 (N_18762,N_17032,N_17461);
or U18763 (N_18763,N_16101,N_17356);
and U18764 (N_18764,N_17382,N_17372);
and U18765 (N_18765,N_17176,N_17164);
and U18766 (N_18766,N_16018,N_17559);
xnor U18767 (N_18767,N_16265,N_16281);
and U18768 (N_18768,N_16176,N_17531);
and U18769 (N_18769,N_17240,N_16471);
or U18770 (N_18770,N_17511,N_17866);
or U18771 (N_18771,N_17791,N_16528);
xor U18772 (N_18772,N_17992,N_17558);
nand U18773 (N_18773,N_17766,N_16822);
xnor U18774 (N_18774,N_16724,N_17600);
or U18775 (N_18775,N_17221,N_17942);
and U18776 (N_18776,N_16632,N_16439);
or U18777 (N_18777,N_17301,N_17634);
nor U18778 (N_18778,N_17849,N_17483);
xor U18779 (N_18779,N_17756,N_17570);
or U18780 (N_18780,N_16759,N_17896);
nor U18781 (N_18781,N_17977,N_16756);
and U18782 (N_18782,N_16694,N_16351);
nand U18783 (N_18783,N_17636,N_17085);
or U18784 (N_18784,N_17411,N_16100);
xnor U18785 (N_18785,N_16895,N_16898);
or U18786 (N_18786,N_16804,N_17593);
or U18787 (N_18787,N_17312,N_17576);
xnor U18788 (N_18788,N_17224,N_17775);
nand U18789 (N_18789,N_16368,N_17330);
and U18790 (N_18790,N_16430,N_17420);
xor U18791 (N_18791,N_16022,N_17092);
nand U18792 (N_18792,N_16796,N_17966);
xnor U18793 (N_18793,N_16495,N_17059);
and U18794 (N_18794,N_17772,N_17344);
xnor U18795 (N_18795,N_16954,N_16188);
nand U18796 (N_18796,N_16702,N_16202);
xor U18797 (N_18797,N_17816,N_17651);
nand U18798 (N_18798,N_16836,N_16435);
xor U18799 (N_18799,N_17479,N_17797);
or U18800 (N_18800,N_16603,N_17987);
nand U18801 (N_18801,N_16924,N_16890);
or U18802 (N_18802,N_16645,N_16226);
and U18803 (N_18803,N_16425,N_17722);
or U18804 (N_18804,N_16175,N_16871);
nor U18805 (N_18805,N_16834,N_16078);
nand U18806 (N_18806,N_16195,N_17645);
nand U18807 (N_18807,N_16848,N_16806);
or U18808 (N_18808,N_16045,N_16944);
or U18809 (N_18809,N_16878,N_17706);
nand U18810 (N_18810,N_17298,N_16813);
nand U18811 (N_18811,N_16033,N_16600);
or U18812 (N_18812,N_17831,N_16492);
and U18813 (N_18813,N_16559,N_16476);
or U18814 (N_18814,N_16741,N_16656);
xnor U18815 (N_18815,N_17443,N_16161);
xor U18816 (N_18816,N_16428,N_16758);
or U18817 (N_18817,N_17668,N_17374);
nor U18818 (N_18818,N_17755,N_17054);
nand U18819 (N_18819,N_16945,N_16448);
and U18820 (N_18820,N_16061,N_17881);
nand U18821 (N_18821,N_16021,N_17911);
or U18822 (N_18822,N_17262,N_17922);
nor U18823 (N_18823,N_17665,N_16618);
or U18824 (N_18824,N_16512,N_16020);
xor U18825 (N_18825,N_16198,N_16613);
nor U18826 (N_18826,N_16904,N_17541);
or U18827 (N_18827,N_17357,N_16902);
xor U18828 (N_18828,N_17080,N_17498);
or U18829 (N_18829,N_16575,N_17686);
nor U18830 (N_18830,N_17504,N_17679);
or U18831 (N_18831,N_16865,N_16278);
xor U18832 (N_18832,N_17376,N_16323);
nand U18833 (N_18833,N_17219,N_16843);
nor U18834 (N_18834,N_16624,N_17557);
and U18835 (N_18835,N_16961,N_16501);
nand U18836 (N_18836,N_17748,N_17709);
xnor U18837 (N_18837,N_17358,N_16415);
xor U18838 (N_18838,N_16173,N_16564);
xnor U18839 (N_18839,N_17782,N_16641);
and U18840 (N_18840,N_17159,N_17743);
nor U18841 (N_18841,N_17122,N_16826);
nand U18842 (N_18842,N_16452,N_16015);
xnor U18843 (N_18843,N_16789,N_17891);
or U18844 (N_18844,N_16634,N_16839);
xor U18845 (N_18845,N_16626,N_17297);
and U18846 (N_18846,N_17954,N_16568);
or U18847 (N_18847,N_16263,N_17355);
or U18848 (N_18848,N_17270,N_17393);
nor U18849 (N_18849,N_16117,N_17714);
xnor U18850 (N_18850,N_16387,N_16973);
nand U18851 (N_18851,N_16217,N_17275);
nand U18852 (N_18852,N_17348,N_16825);
nor U18853 (N_18853,N_17971,N_16548);
xnor U18854 (N_18854,N_16221,N_17869);
and U18855 (N_18855,N_17140,N_16628);
and U18856 (N_18856,N_16150,N_16374);
nand U18857 (N_18857,N_17115,N_16001);
xor U18858 (N_18858,N_17574,N_16223);
xor U18859 (N_18859,N_16200,N_17273);
and U18860 (N_18860,N_17878,N_17015);
xor U18861 (N_18861,N_16866,N_16135);
xnor U18862 (N_18862,N_16388,N_17423);
nor U18863 (N_18863,N_16691,N_16879);
nand U18864 (N_18864,N_17529,N_17850);
nand U18865 (N_18865,N_17788,N_16962);
and U18866 (N_18866,N_17839,N_17276);
and U18867 (N_18867,N_16418,N_16319);
nor U18868 (N_18868,N_17114,N_16259);
xnor U18869 (N_18869,N_17864,N_16977);
nor U18870 (N_18870,N_17844,N_16386);
nand U18871 (N_18871,N_17730,N_16885);
or U18872 (N_18872,N_16365,N_16757);
or U18873 (N_18873,N_16827,N_17979);
or U18874 (N_18874,N_17127,N_17305);
nand U18875 (N_18875,N_17261,N_16794);
nand U18876 (N_18876,N_16006,N_17655);
nand U18877 (N_18877,N_16664,N_16519);
nand U18878 (N_18878,N_16780,N_17776);
nor U18879 (N_18879,N_16783,N_16043);
and U18880 (N_18880,N_17463,N_17110);
nand U18881 (N_18881,N_17350,N_16393);
nor U18882 (N_18882,N_17252,N_17495);
nor U18883 (N_18883,N_16543,N_17646);
nand U18884 (N_18884,N_17212,N_16920);
and U18885 (N_18885,N_17846,N_16693);
nor U18886 (N_18886,N_16532,N_17290);
nand U18887 (N_18887,N_17989,N_16038);
nand U18888 (N_18888,N_17180,N_17807);
and U18889 (N_18889,N_16310,N_16525);
nor U18890 (N_18890,N_17685,N_16377);
nand U18891 (N_18891,N_16251,N_16591);
nand U18892 (N_18892,N_16715,N_16987);
xnor U18893 (N_18893,N_17200,N_16079);
xnor U18894 (N_18894,N_16858,N_17737);
or U18895 (N_18895,N_16570,N_17269);
and U18896 (N_18896,N_16747,N_17727);
and U18897 (N_18897,N_17094,N_16372);
nand U18898 (N_18898,N_16604,N_16552);
xor U18899 (N_18899,N_17742,N_16423);
or U18900 (N_18900,N_16104,N_17516);
xor U18901 (N_18901,N_17075,N_16739);
nor U18902 (N_18902,N_17244,N_17366);
nand U18903 (N_18903,N_16597,N_16093);
or U18904 (N_18904,N_17783,N_16515);
or U18905 (N_18905,N_16233,N_17154);
or U18906 (N_18906,N_16750,N_16411);
nand U18907 (N_18907,N_17313,N_16172);
xnor U18908 (N_18908,N_17434,N_16731);
nand U18909 (N_18909,N_16099,N_16352);
xor U18910 (N_18910,N_17104,N_17188);
nand U18911 (N_18911,N_17824,N_17980);
nor U18912 (N_18912,N_17725,N_17875);
or U18913 (N_18913,N_16507,N_16673);
nand U18914 (N_18914,N_17962,N_17739);
and U18915 (N_18915,N_17800,N_16280);
or U18916 (N_18916,N_17268,N_17056);
nor U18917 (N_18917,N_16403,N_17407);
nor U18918 (N_18918,N_16107,N_17082);
xnor U18919 (N_18919,N_17043,N_17960);
or U18920 (N_18920,N_17522,N_17861);
nand U18921 (N_18921,N_16215,N_16431);
xnor U18922 (N_18922,N_17065,N_16461);
or U18923 (N_18923,N_17673,N_16686);
nand U18924 (N_18924,N_16115,N_16915);
nand U18925 (N_18925,N_16814,N_16889);
xnor U18926 (N_18926,N_16413,N_17061);
nand U18927 (N_18927,N_16793,N_16034);
nand U18928 (N_18928,N_17795,N_16000);
nor U18929 (N_18929,N_16901,N_16770);
and U18930 (N_18930,N_16689,N_16819);
nand U18931 (N_18931,N_16972,N_17703);
or U18932 (N_18932,N_16989,N_17234);
or U18933 (N_18933,N_17400,N_17952);
and U18934 (N_18934,N_16191,N_17251);
nor U18935 (N_18935,N_17699,N_16087);
or U18936 (N_18936,N_17087,N_16165);
nor U18937 (N_18937,N_17692,N_17467);
xnor U18938 (N_18938,N_17218,N_16638);
xnor U18939 (N_18939,N_16795,N_17899);
or U18940 (N_18940,N_17819,N_17172);
xnor U18941 (N_18941,N_17895,N_16152);
or U18942 (N_18942,N_16696,N_17533);
or U18943 (N_18943,N_16145,N_16149);
xnor U18944 (N_18944,N_16210,N_17167);
or U18945 (N_18945,N_17482,N_17614);
and U18946 (N_18946,N_16114,N_16549);
or U18947 (N_18947,N_16294,N_17575);
nand U18948 (N_18948,N_16768,N_16526);
nand U18949 (N_18949,N_16253,N_16477);
nand U18950 (N_18950,N_16674,N_16990);
or U18951 (N_18951,N_17462,N_16550);
xor U18952 (N_18952,N_16112,N_17430);
nand U18953 (N_18953,N_16125,N_17806);
nand U18954 (N_18954,N_16723,N_17264);
nand U18955 (N_18955,N_17066,N_16102);
xnor U18956 (N_18956,N_16729,N_17177);
nand U18957 (N_18957,N_17346,N_16636);
and U18958 (N_18958,N_16292,N_17502);
or U18959 (N_18959,N_17295,N_16103);
nand U18960 (N_18960,N_16019,N_17185);
and U18961 (N_18961,N_16494,N_17494);
and U18962 (N_18962,N_16935,N_17667);
xor U18963 (N_18963,N_16542,N_17246);
and U18964 (N_18964,N_17161,N_17169);
nand U18965 (N_18965,N_17036,N_16993);
nand U18966 (N_18966,N_16710,N_16010);
nor U18967 (N_18967,N_17155,N_16432);
and U18968 (N_18968,N_17294,N_16486);
or U18969 (N_18969,N_17432,N_17232);
nand U18970 (N_18970,N_16230,N_16157);
nor U18971 (N_18971,N_16743,N_17763);
xor U18972 (N_18972,N_17424,N_17038);
nand U18973 (N_18973,N_17051,N_16684);
nor U18974 (N_18974,N_17825,N_17017);
xnor U18975 (N_18975,N_16807,N_16906);
nor U18976 (N_18976,N_17693,N_17787);
nand U18977 (N_18977,N_17711,N_17089);
nand U18978 (N_18978,N_17657,N_16956);
nor U18979 (N_18979,N_17648,N_17460);
and U18980 (N_18980,N_17497,N_17626);
or U18981 (N_18981,N_17459,N_17228);
or U18982 (N_18982,N_16951,N_17547);
xor U18983 (N_18983,N_17436,N_17973);
nor U18984 (N_18984,N_16910,N_17179);
nor U18985 (N_18985,N_17914,N_17880);
nor U18986 (N_18986,N_17886,N_16284);
or U18987 (N_18987,N_17567,N_17681);
or U18988 (N_18988,N_17445,N_16113);
or U18989 (N_18989,N_16266,N_16237);
nor U18990 (N_18990,N_17388,N_16017);
or U18991 (N_18991,N_16441,N_16617);
nand U18992 (N_18992,N_16219,N_17666);
nor U18993 (N_18993,N_16513,N_16305);
or U18994 (N_18994,N_17239,N_16979);
or U18995 (N_18995,N_16643,N_16279);
xor U18996 (N_18996,N_16790,N_16823);
xor U18997 (N_18997,N_16331,N_17862);
or U18998 (N_18998,N_16373,N_16190);
or U18999 (N_18999,N_17242,N_16540);
or U19000 (N_19000,N_16713,N_17802);
nor U19001 (N_19001,N_17896,N_16823);
xor U19002 (N_19002,N_17983,N_17617);
or U19003 (N_19003,N_17733,N_17858);
or U19004 (N_19004,N_17961,N_17868);
xnor U19005 (N_19005,N_17985,N_17769);
and U19006 (N_19006,N_16335,N_17603);
xor U19007 (N_19007,N_16450,N_16984);
nand U19008 (N_19008,N_17366,N_17909);
or U19009 (N_19009,N_16778,N_17867);
nor U19010 (N_19010,N_17585,N_17701);
xor U19011 (N_19011,N_17947,N_17253);
or U19012 (N_19012,N_16837,N_16943);
and U19013 (N_19013,N_16673,N_17814);
nor U19014 (N_19014,N_17879,N_16468);
nor U19015 (N_19015,N_17501,N_17548);
nor U19016 (N_19016,N_16078,N_17916);
nand U19017 (N_19017,N_17605,N_16903);
or U19018 (N_19018,N_17394,N_17669);
nor U19019 (N_19019,N_17484,N_17882);
nor U19020 (N_19020,N_17440,N_16574);
and U19021 (N_19021,N_16436,N_16157);
nor U19022 (N_19022,N_16572,N_17399);
and U19023 (N_19023,N_16017,N_17085);
nor U19024 (N_19024,N_17072,N_17919);
and U19025 (N_19025,N_16685,N_16809);
nor U19026 (N_19026,N_16605,N_16838);
nand U19027 (N_19027,N_17423,N_16878);
xnor U19028 (N_19028,N_17058,N_16689);
nand U19029 (N_19029,N_16640,N_17908);
or U19030 (N_19030,N_16110,N_17256);
nor U19031 (N_19031,N_16103,N_17682);
and U19032 (N_19032,N_16134,N_16245);
nand U19033 (N_19033,N_17093,N_17176);
and U19034 (N_19034,N_17327,N_16535);
nand U19035 (N_19035,N_16865,N_16209);
xnor U19036 (N_19036,N_17804,N_17708);
nand U19037 (N_19037,N_17643,N_16348);
xnor U19038 (N_19038,N_17690,N_17219);
xor U19039 (N_19039,N_17032,N_17650);
xor U19040 (N_19040,N_16520,N_16089);
xor U19041 (N_19041,N_17419,N_17600);
or U19042 (N_19042,N_16812,N_17774);
or U19043 (N_19043,N_17605,N_16644);
nand U19044 (N_19044,N_16159,N_17167);
nor U19045 (N_19045,N_17410,N_16983);
nor U19046 (N_19046,N_17187,N_16586);
nand U19047 (N_19047,N_16061,N_17024);
nor U19048 (N_19048,N_17188,N_16145);
nand U19049 (N_19049,N_16709,N_16253);
nor U19050 (N_19050,N_17919,N_16793);
or U19051 (N_19051,N_16852,N_16011);
xor U19052 (N_19052,N_16977,N_17800);
xor U19053 (N_19053,N_16523,N_16148);
xor U19054 (N_19054,N_17023,N_16953);
nand U19055 (N_19055,N_16129,N_17702);
nor U19056 (N_19056,N_17690,N_16833);
and U19057 (N_19057,N_16762,N_17575);
nor U19058 (N_19058,N_17719,N_16267);
or U19059 (N_19059,N_17476,N_16991);
nor U19060 (N_19060,N_16267,N_16919);
or U19061 (N_19061,N_17446,N_17222);
xor U19062 (N_19062,N_17058,N_16347);
nor U19063 (N_19063,N_17513,N_17810);
nor U19064 (N_19064,N_17618,N_17509);
or U19065 (N_19065,N_16061,N_17453);
and U19066 (N_19066,N_17642,N_17417);
or U19067 (N_19067,N_16970,N_16195);
or U19068 (N_19068,N_17071,N_17366);
or U19069 (N_19069,N_17791,N_17674);
xor U19070 (N_19070,N_16901,N_17956);
and U19071 (N_19071,N_17984,N_17778);
or U19072 (N_19072,N_16835,N_17719);
or U19073 (N_19073,N_17551,N_17571);
nor U19074 (N_19074,N_17313,N_17092);
or U19075 (N_19075,N_16936,N_17219);
xnor U19076 (N_19076,N_16377,N_16384);
and U19077 (N_19077,N_16198,N_17517);
nand U19078 (N_19078,N_16463,N_16858);
or U19079 (N_19079,N_16695,N_16073);
nor U19080 (N_19080,N_17931,N_17589);
nand U19081 (N_19081,N_16503,N_17429);
or U19082 (N_19082,N_16252,N_17007);
nand U19083 (N_19083,N_16321,N_16462);
xor U19084 (N_19084,N_16070,N_17101);
nor U19085 (N_19085,N_17890,N_17898);
xor U19086 (N_19086,N_17965,N_16572);
nand U19087 (N_19087,N_17029,N_17955);
and U19088 (N_19088,N_16805,N_17786);
and U19089 (N_19089,N_17270,N_16228);
nor U19090 (N_19090,N_16330,N_16859);
or U19091 (N_19091,N_16240,N_17094);
and U19092 (N_19092,N_17300,N_17326);
xor U19093 (N_19093,N_17333,N_16455);
xnor U19094 (N_19094,N_17414,N_16526);
nand U19095 (N_19095,N_16404,N_16238);
or U19096 (N_19096,N_17141,N_16210);
nor U19097 (N_19097,N_16074,N_17779);
and U19098 (N_19098,N_17891,N_16754);
and U19099 (N_19099,N_16699,N_17912);
nand U19100 (N_19100,N_16669,N_17699);
and U19101 (N_19101,N_17134,N_16741);
xor U19102 (N_19102,N_16802,N_17468);
xnor U19103 (N_19103,N_16085,N_16315);
xnor U19104 (N_19104,N_17236,N_17341);
or U19105 (N_19105,N_16499,N_16840);
or U19106 (N_19106,N_16692,N_17977);
xnor U19107 (N_19107,N_16740,N_17562);
nor U19108 (N_19108,N_17948,N_17275);
or U19109 (N_19109,N_16342,N_17090);
and U19110 (N_19110,N_16688,N_17977);
xnor U19111 (N_19111,N_17174,N_17193);
xnor U19112 (N_19112,N_16076,N_16835);
xor U19113 (N_19113,N_16330,N_17621);
and U19114 (N_19114,N_16794,N_16390);
and U19115 (N_19115,N_17574,N_17487);
or U19116 (N_19116,N_16978,N_16789);
xor U19117 (N_19117,N_16841,N_16294);
nor U19118 (N_19118,N_16155,N_16494);
and U19119 (N_19119,N_16826,N_16569);
or U19120 (N_19120,N_16928,N_16675);
and U19121 (N_19121,N_16760,N_17912);
nand U19122 (N_19122,N_17400,N_16538);
nand U19123 (N_19123,N_17460,N_16234);
nor U19124 (N_19124,N_17280,N_17323);
and U19125 (N_19125,N_17724,N_16667);
nor U19126 (N_19126,N_17882,N_17160);
nand U19127 (N_19127,N_16353,N_16070);
or U19128 (N_19128,N_17827,N_17201);
or U19129 (N_19129,N_16437,N_16722);
nor U19130 (N_19130,N_16809,N_16910);
nor U19131 (N_19131,N_16603,N_16343);
or U19132 (N_19132,N_16711,N_17969);
and U19133 (N_19133,N_16749,N_16175);
xnor U19134 (N_19134,N_16147,N_17480);
nor U19135 (N_19135,N_17101,N_17640);
nor U19136 (N_19136,N_16725,N_16355);
xor U19137 (N_19137,N_16668,N_17846);
xor U19138 (N_19138,N_17092,N_17083);
nand U19139 (N_19139,N_16835,N_17112);
nor U19140 (N_19140,N_16164,N_17721);
nand U19141 (N_19141,N_17818,N_17290);
nor U19142 (N_19142,N_16662,N_16896);
or U19143 (N_19143,N_16257,N_16412);
or U19144 (N_19144,N_17519,N_17787);
and U19145 (N_19145,N_17472,N_17971);
and U19146 (N_19146,N_17407,N_16385);
nand U19147 (N_19147,N_17910,N_17175);
or U19148 (N_19148,N_17992,N_17581);
xor U19149 (N_19149,N_16863,N_17040);
xor U19150 (N_19150,N_17751,N_16895);
nand U19151 (N_19151,N_16495,N_17413);
nor U19152 (N_19152,N_16812,N_16634);
and U19153 (N_19153,N_16425,N_17781);
nand U19154 (N_19154,N_16109,N_16927);
xnor U19155 (N_19155,N_17808,N_17546);
nor U19156 (N_19156,N_17459,N_17638);
xor U19157 (N_19157,N_16853,N_17629);
nand U19158 (N_19158,N_17045,N_16937);
nor U19159 (N_19159,N_16197,N_17206);
and U19160 (N_19160,N_17119,N_16792);
xor U19161 (N_19161,N_16961,N_16779);
nor U19162 (N_19162,N_16757,N_17492);
or U19163 (N_19163,N_16547,N_17899);
nor U19164 (N_19164,N_17955,N_17484);
xnor U19165 (N_19165,N_17866,N_16609);
xor U19166 (N_19166,N_16213,N_16353);
or U19167 (N_19167,N_17068,N_17389);
xor U19168 (N_19168,N_16939,N_17287);
xnor U19169 (N_19169,N_16050,N_17352);
nand U19170 (N_19170,N_17441,N_16795);
or U19171 (N_19171,N_16820,N_17115);
xor U19172 (N_19172,N_16908,N_16933);
or U19173 (N_19173,N_17802,N_17955);
nor U19174 (N_19174,N_16295,N_16801);
or U19175 (N_19175,N_17967,N_16789);
xor U19176 (N_19176,N_16435,N_17723);
nor U19177 (N_19177,N_16529,N_17586);
nor U19178 (N_19178,N_17580,N_16342);
or U19179 (N_19179,N_16184,N_16835);
or U19180 (N_19180,N_17616,N_17601);
and U19181 (N_19181,N_17091,N_17705);
nand U19182 (N_19182,N_17132,N_16280);
nand U19183 (N_19183,N_16795,N_16426);
nand U19184 (N_19184,N_16032,N_17809);
nor U19185 (N_19185,N_16491,N_16542);
xnor U19186 (N_19186,N_17105,N_17424);
or U19187 (N_19187,N_16721,N_17956);
and U19188 (N_19188,N_16244,N_17009);
or U19189 (N_19189,N_16298,N_16897);
or U19190 (N_19190,N_17023,N_17310);
or U19191 (N_19191,N_16048,N_16528);
nor U19192 (N_19192,N_16194,N_16461);
xnor U19193 (N_19193,N_16237,N_17821);
or U19194 (N_19194,N_17927,N_16928);
or U19195 (N_19195,N_17225,N_17852);
and U19196 (N_19196,N_17202,N_16559);
xor U19197 (N_19197,N_17347,N_16721);
nand U19198 (N_19198,N_16722,N_16097);
nor U19199 (N_19199,N_17896,N_16100);
nor U19200 (N_19200,N_16627,N_17874);
and U19201 (N_19201,N_17422,N_17901);
nand U19202 (N_19202,N_16518,N_16142);
nand U19203 (N_19203,N_17702,N_17073);
nor U19204 (N_19204,N_16625,N_17370);
and U19205 (N_19205,N_16470,N_16858);
nor U19206 (N_19206,N_16310,N_17258);
xnor U19207 (N_19207,N_17694,N_17190);
xor U19208 (N_19208,N_17230,N_16032);
xnor U19209 (N_19209,N_17596,N_17190);
nor U19210 (N_19210,N_16813,N_17637);
and U19211 (N_19211,N_16772,N_17330);
nand U19212 (N_19212,N_16102,N_17012);
or U19213 (N_19213,N_16261,N_16606);
and U19214 (N_19214,N_17074,N_17187);
or U19215 (N_19215,N_17352,N_17093);
nand U19216 (N_19216,N_17302,N_17123);
nand U19217 (N_19217,N_16305,N_17853);
nor U19218 (N_19218,N_17836,N_17289);
and U19219 (N_19219,N_17070,N_17278);
nand U19220 (N_19220,N_17905,N_17576);
and U19221 (N_19221,N_16479,N_17032);
and U19222 (N_19222,N_16035,N_16042);
xnor U19223 (N_19223,N_17848,N_16937);
nor U19224 (N_19224,N_16084,N_16746);
xnor U19225 (N_19225,N_16105,N_16728);
nand U19226 (N_19226,N_16442,N_16450);
nand U19227 (N_19227,N_16442,N_17400);
nand U19228 (N_19228,N_16279,N_17553);
nand U19229 (N_19229,N_17793,N_16635);
and U19230 (N_19230,N_17687,N_17668);
nor U19231 (N_19231,N_16503,N_16976);
nand U19232 (N_19232,N_17229,N_16907);
xnor U19233 (N_19233,N_17674,N_17762);
nor U19234 (N_19234,N_17630,N_17922);
and U19235 (N_19235,N_16608,N_17857);
or U19236 (N_19236,N_16300,N_17583);
xnor U19237 (N_19237,N_16596,N_16618);
xnor U19238 (N_19238,N_17151,N_16066);
or U19239 (N_19239,N_17945,N_16101);
xnor U19240 (N_19240,N_16243,N_16967);
xor U19241 (N_19241,N_16098,N_17903);
xnor U19242 (N_19242,N_17964,N_16726);
xnor U19243 (N_19243,N_17384,N_17054);
nand U19244 (N_19244,N_17263,N_16932);
or U19245 (N_19245,N_17640,N_17253);
nand U19246 (N_19246,N_16937,N_17618);
and U19247 (N_19247,N_16345,N_17057);
xor U19248 (N_19248,N_16799,N_16872);
nand U19249 (N_19249,N_16634,N_17465);
and U19250 (N_19250,N_16131,N_17639);
xnor U19251 (N_19251,N_17966,N_16426);
or U19252 (N_19252,N_17135,N_16992);
or U19253 (N_19253,N_16675,N_17765);
nor U19254 (N_19254,N_17574,N_16184);
nor U19255 (N_19255,N_17680,N_17409);
and U19256 (N_19256,N_17305,N_17692);
nor U19257 (N_19257,N_16714,N_17840);
and U19258 (N_19258,N_16461,N_17750);
or U19259 (N_19259,N_17355,N_17610);
nor U19260 (N_19260,N_16060,N_16759);
nor U19261 (N_19261,N_17300,N_16331);
and U19262 (N_19262,N_16168,N_17435);
or U19263 (N_19263,N_16424,N_17808);
or U19264 (N_19264,N_17123,N_17962);
xnor U19265 (N_19265,N_17254,N_17344);
and U19266 (N_19266,N_16848,N_17152);
and U19267 (N_19267,N_17840,N_17682);
or U19268 (N_19268,N_17931,N_17640);
or U19269 (N_19269,N_17259,N_16057);
xor U19270 (N_19270,N_17892,N_17287);
or U19271 (N_19271,N_16461,N_17872);
or U19272 (N_19272,N_16390,N_17373);
xor U19273 (N_19273,N_17557,N_17908);
and U19274 (N_19274,N_16824,N_16411);
nand U19275 (N_19275,N_17523,N_16514);
nor U19276 (N_19276,N_16864,N_16741);
xnor U19277 (N_19277,N_17445,N_16181);
and U19278 (N_19278,N_17624,N_16554);
nor U19279 (N_19279,N_16957,N_16455);
or U19280 (N_19280,N_16415,N_17466);
nor U19281 (N_19281,N_16631,N_17519);
nor U19282 (N_19282,N_17197,N_16471);
xnor U19283 (N_19283,N_17164,N_17355);
xnor U19284 (N_19284,N_16803,N_16878);
xor U19285 (N_19285,N_16495,N_16576);
or U19286 (N_19286,N_16323,N_16707);
or U19287 (N_19287,N_17854,N_17461);
or U19288 (N_19288,N_17537,N_17615);
or U19289 (N_19289,N_16777,N_17046);
nor U19290 (N_19290,N_16532,N_17177);
and U19291 (N_19291,N_17666,N_17394);
and U19292 (N_19292,N_17011,N_17392);
and U19293 (N_19293,N_17672,N_17980);
nor U19294 (N_19294,N_17135,N_16873);
xnor U19295 (N_19295,N_17879,N_17054);
xor U19296 (N_19296,N_16095,N_16416);
or U19297 (N_19297,N_16543,N_16838);
nand U19298 (N_19298,N_17710,N_17190);
nand U19299 (N_19299,N_16809,N_16610);
nand U19300 (N_19300,N_17815,N_16838);
xnor U19301 (N_19301,N_16587,N_17868);
and U19302 (N_19302,N_17775,N_16264);
or U19303 (N_19303,N_17917,N_16330);
and U19304 (N_19304,N_16278,N_17421);
and U19305 (N_19305,N_17338,N_17746);
or U19306 (N_19306,N_16813,N_17961);
and U19307 (N_19307,N_16457,N_17527);
and U19308 (N_19308,N_16747,N_16901);
nand U19309 (N_19309,N_17263,N_17884);
xor U19310 (N_19310,N_17706,N_16149);
nand U19311 (N_19311,N_17504,N_16890);
and U19312 (N_19312,N_16283,N_16929);
or U19313 (N_19313,N_17134,N_16710);
and U19314 (N_19314,N_16071,N_17649);
or U19315 (N_19315,N_16287,N_16627);
nor U19316 (N_19316,N_16544,N_17809);
nand U19317 (N_19317,N_17224,N_17155);
nor U19318 (N_19318,N_16158,N_17404);
and U19319 (N_19319,N_16196,N_17434);
nor U19320 (N_19320,N_16186,N_16195);
and U19321 (N_19321,N_16095,N_16324);
and U19322 (N_19322,N_16517,N_17378);
and U19323 (N_19323,N_16301,N_17807);
xor U19324 (N_19324,N_16252,N_17899);
xor U19325 (N_19325,N_17036,N_17248);
and U19326 (N_19326,N_16700,N_16533);
nor U19327 (N_19327,N_17841,N_17682);
or U19328 (N_19328,N_16024,N_17713);
and U19329 (N_19329,N_17544,N_17502);
nand U19330 (N_19330,N_17665,N_17861);
or U19331 (N_19331,N_16374,N_16422);
xnor U19332 (N_19332,N_17393,N_17206);
xnor U19333 (N_19333,N_17437,N_16080);
and U19334 (N_19334,N_16034,N_16633);
and U19335 (N_19335,N_17424,N_17922);
and U19336 (N_19336,N_17270,N_16994);
or U19337 (N_19337,N_16030,N_16205);
nand U19338 (N_19338,N_17520,N_16236);
nand U19339 (N_19339,N_17985,N_17206);
nand U19340 (N_19340,N_17166,N_16848);
nand U19341 (N_19341,N_17235,N_16779);
or U19342 (N_19342,N_16940,N_16310);
or U19343 (N_19343,N_17387,N_17728);
nand U19344 (N_19344,N_16225,N_16683);
or U19345 (N_19345,N_16737,N_16872);
nor U19346 (N_19346,N_17700,N_17681);
and U19347 (N_19347,N_17946,N_16983);
nand U19348 (N_19348,N_17053,N_16999);
or U19349 (N_19349,N_16922,N_16975);
nand U19350 (N_19350,N_16917,N_17434);
or U19351 (N_19351,N_16342,N_17198);
and U19352 (N_19352,N_16672,N_17585);
nor U19353 (N_19353,N_17710,N_17012);
and U19354 (N_19354,N_17918,N_16721);
or U19355 (N_19355,N_16648,N_17240);
or U19356 (N_19356,N_17150,N_16680);
and U19357 (N_19357,N_17277,N_17051);
xor U19358 (N_19358,N_17055,N_17971);
and U19359 (N_19359,N_16499,N_16728);
xnor U19360 (N_19360,N_17977,N_16257);
nor U19361 (N_19361,N_17760,N_17908);
xor U19362 (N_19362,N_16762,N_16766);
or U19363 (N_19363,N_17996,N_17649);
nor U19364 (N_19364,N_17536,N_16584);
or U19365 (N_19365,N_17154,N_16277);
xor U19366 (N_19366,N_17107,N_16611);
or U19367 (N_19367,N_16285,N_16995);
nand U19368 (N_19368,N_17416,N_16504);
nor U19369 (N_19369,N_17127,N_16427);
nand U19370 (N_19370,N_16739,N_16779);
or U19371 (N_19371,N_16473,N_16011);
and U19372 (N_19372,N_17781,N_16202);
nand U19373 (N_19373,N_17267,N_17758);
nor U19374 (N_19374,N_16805,N_17667);
nor U19375 (N_19375,N_16073,N_16897);
nand U19376 (N_19376,N_17579,N_16723);
xor U19377 (N_19377,N_16584,N_16429);
and U19378 (N_19378,N_16972,N_17830);
nand U19379 (N_19379,N_16201,N_17421);
and U19380 (N_19380,N_17877,N_17854);
xor U19381 (N_19381,N_16568,N_16902);
nor U19382 (N_19382,N_17680,N_17277);
xnor U19383 (N_19383,N_17793,N_17204);
or U19384 (N_19384,N_16490,N_17753);
nand U19385 (N_19385,N_16118,N_17247);
xor U19386 (N_19386,N_17587,N_17473);
and U19387 (N_19387,N_17198,N_16695);
nor U19388 (N_19388,N_17649,N_17345);
and U19389 (N_19389,N_16532,N_17506);
or U19390 (N_19390,N_17383,N_17438);
nor U19391 (N_19391,N_16591,N_17585);
or U19392 (N_19392,N_16532,N_16365);
and U19393 (N_19393,N_16649,N_16118);
xnor U19394 (N_19394,N_17712,N_16616);
nor U19395 (N_19395,N_17036,N_17210);
nor U19396 (N_19396,N_16982,N_16097);
and U19397 (N_19397,N_16255,N_16450);
nand U19398 (N_19398,N_17358,N_17233);
or U19399 (N_19399,N_16710,N_16928);
nor U19400 (N_19400,N_16288,N_17776);
and U19401 (N_19401,N_17306,N_17998);
nand U19402 (N_19402,N_17759,N_17146);
and U19403 (N_19403,N_17265,N_16734);
or U19404 (N_19404,N_16089,N_17505);
nand U19405 (N_19405,N_16594,N_17382);
nor U19406 (N_19406,N_17177,N_17091);
and U19407 (N_19407,N_16675,N_16007);
or U19408 (N_19408,N_17121,N_17626);
nor U19409 (N_19409,N_16219,N_16140);
or U19410 (N_19410,N_17778,N_17081);
xnor U19411 (N_19411,N_16481,N_16405);
xor U19412 (N_19412,N_16443,N_16322);
nand U19413 (N_19413,N_17004,N_16778);
nor U19414 (N_19414,N_16834,N_16369);
xnor U19415 (N_19415,N_16149,N_16121);
nand U19416 (N_19416,N_17147,N_17778);
nor U19417 (N_19417,N_17945,N_16874);
nor U19418 (N_19418,N_16336,N_17702);
nor U19419 (N_19419,N_16828,N_17004);
and U19420 (N_19420,N_16631,N_16241);
nor U19421 (N_19421,N_17157,N_17802);
nor U19422 (N_19422,N_16790,N_16760);
or U19423 (N_19423,N_17187,N_16176);
and U19424 (N_19424,N_17003,N_17307);
xor U19425 (N_19425,N_17744,N_17106);
nand U19426 (N_19426,N_17193,N_16098);
and U19427 (N_19427,N_16319,N_17441);
and U19428 (N_19428,N_17827,N_16151);
or U19429 (N_19429,N_16849,N_16688);
and U19430 (N_19430,N_17445,N_17779);
xor U19431 (N_19431,N_16287,N_17145);
xor U19432 (N_19432,N_16295,N_17280);
and U19433 (N_19433,N_16260,N_16033);
or U19434 (N_19434,N_17019,N_16569);
or U19435 (N_19435,N_16291,N_16358);
nand U19436 (N_19436,N_17829,N_17705);
nor U19437 (N_19437,N_16438,N_16385);
and U19438 (N_19438,N_16473,N_16165);
nor U19439 (N_19439,N_17184,N_16167);
and U19440 (N_19440,N_17911,N_16332);
nand U19441 (N_19441,N_16017,N_16653);
or U19442 (N_19442,N_16222,N_17285);
and U19443 (N_19443,N_16765,N_17822);
or U19444 (N_19444,N_17638,N_17007);
and U19445 (N_19445,N_16730,N_16107);
xnor U19446 (N_19446,N_17244,N_16599);
or U19447 (N_19447,N_16555,N_16504);
xnor U19448 (N_19448,N_16190,N_16429);
nor U19449 (N_19449,N_17592,N_17348);
xor U19450 (N_19450,N_16397,N_16524);
nor U19451 (N_19451,N_17823,N_16375);
and U19452 (N_19452,N_17059,N_17601);
nor U19453 (N_19453,N_17600,N_16530);
nor U19454 (N_19454,N_16079,N_17746);
nor U19455 (N_19455,N_17750,N_16373);
and U19456 (N_19456,N_17929,N_16987);
and U19457 (N_19457,N_16065,N_17150);
and U19458 (N_19458,N_16805,N_16737);
and U19459 (N_19459,N_16289,N_16377);
or U19460 (N_19460,N_16028,N_16904);
nor U19461 (N_19461,N_16545,N_17288);
nand U19462 (N_19462,N_17122,N_17518);
and U19463 (N_19463,N_17862,N_17985);
and U19464 (N_19464,N_16106,N_17544);
and U19465 (N_19465,N_17391,N_17129);
nor U19466 (N_19466,N_16116,N_17243);
nor U19467 (N_19467,N_17113,N_16807);
and U19468 (N_19468,N_16587,N_16981);
nor U19469 (N_19469,N_16751,N_17839);
nand U19470 (N_19470,N_17357,N_16406);
nand U19471 (N_19471,N_16787,N_17179);
xor U19472 (N_19472,N_17348,N_17426);
or U19473 (N_19473,N_17629,N_16482);
or U19474 (N_19474,N_17034,N_17423);
nor U19475 (N_19475,N_16525,N_17121);
or U19476 (N_19476,N_16133,N_16668);
or U19477 (N_19477,N_16904,N_16983);
or U19478 (N_19478,N_17807,N_17589);
xor U19479 (N_19479,N_16823,N_17271);
nor U19480 (N_19480,N_16907,N_17473);
and U19481 (N_19481,N_16283,N_17208);
xor U19482 (N_19482,N_17514,N_16393);
nor U19483 (N_19483,N_17408,N_16911);
xnor U19484 (N_19484,N_16813,N_17144);
and U19485 (N_19485,N_17355,N_16788);
xnor U19486 (N_19486,N_16242,N_16375);
nand U19487 (N_19487,N_16480,N_16152);
nand U19488 (N_19488,N_16105,N_16975);
nor U19489 (N_19489,N_16610,N_17710);
xor U19490 (N_19490,N_16087,N_17252);
xnor U19491 (N_19491,N_17331,N_17149);
nor U19492 (N_19492,N_17653,N_16794);
or U19493 (N_19493,N_17606,N_16969);
and U19494 (N_19494,N_17304,N_16004);
xnor U19495 (N_19495,N_16106,N_16142);
xor U19496 (N_19496,N_17561,N_16207);
nand U19497 (N_19497,N_16794,N_17773);
nand U19498 (N_19498,N_16604,N_16797);
and U19499 (N_19499,N_16459,N_17167);
nor U19500 (N_19500,N_17283,N_16966);
and U19501 (N_19501,N_16758,N_16118);
or U19502 (N_19502,N_16907,N_16557);
and U19503 (N_19503,N_16860,N_17581);
nand U19504 (N_19504,N_17447,N_17135);
nor U19505 (N_19505,N_17049,N_16085);
or U19506 (N_19506,N_16494,N_17792);
and U19507 (N_19507,N_17903,N_16760);
and U19508 (N_19508,N_17689,N_16768);
nor U19509 (N_19509,N_16594,N_16771);
nor U19510 (N_19510,N_17392,N_16106);
or U19511 (N_19511,N_17269,N_16856);
xor U19512 (N_19512,N_17338,N_16799);
xnor U19513 (N_19513,N_16440,N_17487);
or U19514 (N_19514,N_16934,N_16362);
nand U19515 (N_19515,N_16521,N_16601);
xor U19516 (N_19516,N_17047,N_16023);
and U19517 (N_19517,N_16976,N_16379);
xnor U19518 (N_19518,N_16347,N_17729);
nor U19519 (N_19519,N_17182,N_16090);
nand U19520 (N_19520,N_17763,N_16537);
or U19521 (N_19521,N_16948,N_17718);
nand U19522 (N_19522,N_17742,N_16633);
nand U19523 (N_19523,N_17349,N_16265);
or U19524 (N_19524,N_16694,N_16539);
nand U19525 (N_19525,N_17604,N_17664);
nand U19526 (N_19526,N_16094,N_17341);
and U19527 (N_19527,N_16735,N_16541);
and U19528 (N_19528,N_17114,N_17424);
nand U19529 (N_19529,N_16047,N_16314);
xor U19530 (N_19530,N_17326,N_17206);
xor U19531 (N_19531,N_17981,N_17968);
xnor U19532 (N_19532,N_17921,N_16721);
nand U19533 (N_19533,N_16045,N_16366);
xor U19534 (N_19534,N_16598,N_17669);
and U19535 (N_19535,N_17310,N_16151);
nand U19536 (N_19536,N_17186,N_16133);
and U19537 (N_19537,N_16898,N_17086);
nor U19538 (N_19538,N_17494,N_16129);
nor U19539 (N_19539,N_16971,N_16911);
nor U19540 (N_19540,N_16108,N_16322);
nor U19541 (N_19541,N_16800,N_17321);
xnor U19542 (N_19542,N_16326,N_16026);
or U19543 (N_19543,N_17045,N_16274);
nand U19544 (N_19544,N_16768,N_17064);
xor U19545 (N_19545,N_16721,N_17098);
or U19546 (N_19546,N_16605,N_16461);
or U19547 (N_19547,N_17767,N_16566);
and U19548 (N_19548,N_17308,N_16588);
nor U19549 (N_19549,N_17282,N_17212);
nand U19550 (N_19550,N_16953,N_17582);
nand U19551 (N_19551,N_17575,N_16969);
nand U19552 (N_19552,N_16959,N_16990);
nor U19553 (N_19553,N_17936,N_17451);
and U19554 (N_19554,N_17637,N_17551);
and U19555 (N_19555,N_16034,N_16172);
and U19556 (N_19556,N_17622,N_17317);
nand U19557 (N_19557,N_16657,N_16859);
nor U19558 (N_19558,N_16310,N_16472);
nor U19559 (N_19559,N_17183,N_17799);
nor U19560 (N_19560,N_16976,N_16763);
and U19561 (N_19561,N_17277,N_16901);
and U19562 (N_19562,N_16420,N_17518);
and U19563 (N_19563,N_16905,N_17921);
or U19564 (N_19564,N_16556,N_17922);
nor U19565 (N_19565,N_17575,N_17649);
xnor U19566 (N_19566,N_17313,N_17938);
nand U19567 (N_19567,N_17390,N_17191);
nand U19568 (N_19568,N_17789,N_16219);
nor U19569 (N_19569,N_16183,N_17397);
and U19570 (N_19570,N_16467,N_17695);
nand U19571 (N_19571,N_17665,N_16468);
xnor U19572 (N_19572,N_16827,N_16396);
nor U19573 (N_19573,N_16048,N_16913);
and U19574 (N_19574,N_17262,N_16015);
xnor U19575 (N_19575,N_16902,N_16347);
or U19576 (N_19576,N_16740,N_17228);
nand U19577 (N_19577,N_17268,N_16744);
or U19578 (N_19578,N_17512,N_16864);
or U19579 (N_19579,N_17091,N_17310);
nor U19580 (N_19580,N_17646,N_16195);
nor U19581 (N_19581,N_17987,N_17453);
and U19582 (N_19582,N_16543,N_17066);
or U19583 (N_19583,N_16526,N_16362);
nor U19584 (N_19584,N_17341,N_17471);
nor U19585 (N_19585,N_17852,N_16811);
nand U19586 (N_19586,N_16272,N_17780);
and U19587 (N_19587,N_17646,N_16519);
nand U19588 (N_19588,N_16509,N_17004);
nand U19589 (N_19589,N_17098,N_17979);
xor U19590 (N_19590,N_17720,N_16833);
and U19591 (N_19591,N_16158,N_16537);
nand U19592 (N_19592,N_16943,N_16871);
nor U19593 (N_19593,N_17815,N_17494);
xnor U19594 (N_19594,N_17694,N_16254);
nand U19595 (N_19595,N_17934,N_16511);
and U19596 (N_19596,N_16563,N_16424);
nand U19597 (N_19597,N_16418,N_16460);
nand U19598 (N_19598,N_17363,N_16046);
nor U19599 (N_19599,N_16626,N_17314);
and U19600 (N_19600,N_16211,N_17328);
and U19601 (N_19601,N_16200,N_17491);
xor U19602 (N_19602,N_17961,N_17753);
nor U19603 (N_19603,N_17091,N_16087);
xnor U19604 (N_19604,N_17642,N_16189);
and U19605 (N_19605,N_16547,N_17112);
or U19606 (N_19606,N_17368,N_17887);
or U19607 (N_19607,N_17389,N_16359);
xnor U19608 (N_19608,N_17045,N_17886);
nor U19609 (N_19609,N_16922,N_16052);
nor U19610 (N_19610,N_17240,N_17060);
and U19611 (N_19611,N_16240,N_16498);
xor U19612 (N_19612,N_17330,N_17076);
xor U19613 (N_19613,N_17878,N_17947);
or U19614 (N_19614,N_16083,N_17928);
and U19615 (N_19615,N_17999,N_16973);
nor U19616 (N_19616,N_16056,N_16641);
nor U19617 (N_19617,N_17909,N_17820);
or U19618 (N_19618,N_16513,N_17957);
nand U19619 (N_19619,N_17514,N_16526);
nand U19620 (N_19620,N_16594,N_16994);
xor U19621 (N_19621,N_16111,N_16206);
nor U19622 (N_19622,N_16317,N_17296);
xnor U19623 (N_19623,N_16408,N_16905);
and U19624 (N_19624,N_17432,N_17326);
or U19625 (N_19625,N_17908,N_16395);
nand U19626 (N_19626,N_16779,N_16999);
and U19627 (N_19627,N_17225,N_17367);
and U19628 (N_19628,N_16912,N_16581);
or U19629 (N_19629,N_16469,N_17734);
or U19630 (N_19630,N_17381,N_17984);
nand U19631 (N_19631,N_17014,N_17986);
or U19632 (N_19632,N_17369,N_17318);
or U19633 (N_19633,N_17490,N_17823);
or U19634 (N_19634,N_16540,N_16313);
xor U19635 (N_19635,N_17890,N_16463);
or U19636 (N_19636,N_17855,N_16838);
xnor U19637 (N_19637,N_16736,N_17899);
or U19638 (N_19638,N_16664,N_16833);
xor U19639 (N_19639,N_16801,N_16994);
or U19640 (N_19640,N_17986,N_16895);
nand U19641 (N_19641,N_16778,N_17094);
and U19642 (N_19642,N_16743,N_17583);
nor U19643 (N_19643,N_17066,N_17433);
nand U19644 (N_19644,N_16518,N_17518);
xnor U19645 (N_19645,N_17065,N_17077);
nand U19646 (N_19646,N_17997,N_17738);
nand U19647 (N_19647,N_17163,N_16193);
nand U19648 (N_19648,N_17724,N_17130);
or U19649 (N_19649,N_16386,N_17547);
nor U19650 (N_19650,N_16187,N_17272);
xor U19651 (N_19651,N_17354,N_17309);
nand U19652 (N_19652,N_16140,N_17798);
nor U19653 (N_19653,N_16615,N_17375);
and U19654 (N_19654,N_16994,N_17608);
xor U19655 (N_19655,N_17894,N_16745);
or U19656 (N_19656,N_17224,N_16129);
and U19657 (N_19657,N_16548,N_16772);
nand U19658 (N_19658,N_16310,N_16661);
xor U19659 (N_19659,N_16294,N_16798);
nor U19660 (N_19660,N_16444,N_16916);
xnor U19661 (N_19661,N_16606,N_16984);
nand U19662 (N_19662,N_16440,N_17359);
xor U19663 (N_19663,N_16694,N_17098);
nor U19664 (N_19664,N_16651,N_17486);
and U19665 (N_19665,N_17325,N_17938);
nor U19666 (N_19666,N_17760,N_16330);
nand U19667 (N_19667,N_17062,N_17856);
nor U19668 (N_19668,N_17586,N_16416);
nand U19669 (N_19669,N_16253,N_17520);
and U19670 (N_19670,N_17362,N_17469);
xor U19671 (N_19671,N_16566,N_16979);
and U19672 (N_19672,N_17134,N_16972);
nand U19673 (N_19673,N_17615,N_17029);
nor U19674 (N_19674,N_17282,N_16948);
nand U19675 (N_19675,N_16912,N_17435);
nand U19676 (N_19676,N_17774,N_17254);
nand U19677 (N_19677,N_16133,N_17417);
xnor U19678 (N_19678,N_17979,N_16285);
nand U19679 (N_19679,N_17084,N_16467);
nor U19680 (N_19680,N_16531,N_16231);
nand U19681 (N_19681,N_17937,N_16676);
and U19682 (N_19682,N_17192,N_17584);
xnor U19683 (N_19683,N_17473,N_17171);
nand U19684 (N_19684,N_17173,N_17276);
nor U19685 (N_19685,N_16874,N_17977);
and U19686 (N_19686,N_17053,N_17365);
xnor U19687 (N_19687,N_16832,N_17909);
nand U19688 (N_19688,N_16160,N_17250);
and U19689 (N_19689,N_16665,N_16331);
nor U19690 (N_19690,N_17108,N_17688);
xnor U19691 (N_19691,N_17333,N_17298);
nor U19692 (N_19692,N_16025,N_16125);
nand U19693 (N_19693,N_17102,N_17203);
or U19694 (N_19694,N_17953,N_16962);
xnor U19695 (N_19695,N_17455,N_16772);
nand U19696 (N_19696,N_16046,N_16438);
nand U19697 (N_19697,N_17483,N_17184);
and U19698 (N_19698,N_17934,N_17379);
nand U19699 (N_19699,N_17418,N_16415);
nand U19700 (N_19700,N_16002,N_16562);
nor U19701 (N_19701,N_17079,N_16005);
nand U19702 (N_19702,N_16054,N_17579);
xnor U19703 (N_19703,N_16402,N_16484);
nand U19704 (N_19704,N_16935,N_16623);
and U19705 (N_19705,N_16102,N_17545);
or U19706 (N_19706,N_17533,N_16434);
and U19707 (N_19707,N_17408,N_16062);
nand U19708 (N_19708,N_17277,N_17884);
xnor U19709 (N_19709,N_17270,N_16112);
and U19710 (N_19710,N_16144,N_16356);
or U19711 (N_19711,N_16630,N_16299);
nor U19712 (N_19712,N_17486,N_16448);
or U19713 (N_19713,N_16053,N_16544);
or U19714 (N_19714,N_17238,N_17003);
xor U19715 (N_19715,N_16725,N_17357);
xor U19716 (N_19716,N_17670,N_17646);
or U19717 (N_19717,N_16921,N_17881);
xnor U19718 (N_19718,N_17288,N_17055);
nor U19719 (N_19719,N_17979,N_17677);
and U19720 (N_19720,N_17711,N_16286);
and U19721 (N_19721,N_17094,N_17757);
and U19722 (N_19722,N_16236,N_16171);
nor U19723 (N_19723,N_16974,N_17766);
xnor U19724 (N_19724,N_16539,N_17328);
or U19725 (N_19725,N_17391,N_16873);
or U19726 (N_19726,N_16736,N_17943);
xnor U19727 (N_19727,N_17691,N_16881);
nor U19728 (N_19728,N_17525,N_16486);
xor U19729 (N_19729,N_16966,N_17247);
xnor U19730 (N_19730,N_16736,N_17654);
xor U19731 (N_19731,N_17796,N_16475);
or U19732 (N_19732,N_16422,N_17487);
nor U19733 (N_19733,N_17157,N_17906);
nor U19734 (N_19734,N_16450,N_17295);
or U19735 (N_19735,N_17994,N_17360);
xor U19736 (N_19736,N_16066,N_17907);
and U19737 (N_19737,N_17278,N_16741);
and U19738 (N_19738,N_17688,N_16184);
or U19739 (N_19739,N_16048,N_17456);
nand U19740 (N_19740,N_16040,N_17534);
nor U19741 (N_19741,N_16153,N_16722);
and U19742 (N_19742,N_17251,N_17554);
nor U19743 (N_19743,N_16650,N_16620);
nand U19744 (N_19744,N_16995,N_17214);
or U19745 (N_19745,N_17216,N_16826);
and U19746 (N_19746,N_16379,N_16604);
xor U19747 (N_19747,N_16135,N_16510);
nand U19748 (N_19748,N_17829,N_16501);
nand U19749 (N_19749,N_16177,N_16302);
or U19750 (N_19750,N_16702,N_16170);
xnor U19751 (N_19751,N_17229,N_16339);
or U19752 (N_19752,N_17339,N_16546);
nand U19753 (N_19753,N_17778,N_16356);
and U19754 (N_19754,N_17459,N_16827);
nand U19755 (N_19755,N_17744,N_16080);
xor U19756 (N_19756,N_17435,N_17265);
xor U19757 (N_19757,N_17827,N_17400);
xor U19758 (N_19758,N_17325,N_17301);
nor U19759 (N_19759,N_16974,N_17825);
xor U19760 (N_19760,N_16770,N_16557);
or U19761 (N_19761,N_16596,N_17168);
xor U19762 (N_19762,N_17926,N_17989);
xor U19763 (N_19763,N_17594,N_17393);
nand U19764 (N_19764,N_16563,N_16929);
xor U19765 (N_19765,N_16460,N_16924);
and U19766 (N_19766,N_16351,N_16359);
nand U19767 (N_19767,N_16665,N_16856);
or U19768 (N_19768,N_17217,N_17781);
and U19769 (N_19769,N_17319,N_16407);
nor U19770 (N_19770,N_17849,N_17441);
nand U19771 (N_19771,N_16354,N_16651);
or U19772 (N_19772,N_17895,N_17396);
and U19773 (N_19773,N_17129,N_16962);
nand U19774 (N_19774,N_17651,N_16520);
xor U19775 (N_19775,N_17653,N_16613);
xor U19776 (N_19776,N_16622,N_16850);
nor U19777 (N_19777,N_16140,N_17239);
or U19778 (N_19778,N_16127,N_16803);
and U19779 (N_19779,N_16624,N_16839);
xnor U19780 (N_19780,N_16061,N_16761);
nor U19781 (N_19781,N_16709,N_16433);
xor U19782 (N_19782,N_17856,N_16753);
and U19783 (N_19783,N_16439,N_16074);
nand U19784 (N_19784,N_16298,N_17372);
nor U19785 (N_19785,N_16046,N_17360);
nand U19786 (N_19786,N_16256,N_16853);
and U19787 (N_19787,N_16031,N_17393);
nand U19788 (N_19788,N_16022,N_17014);
and U19789 (N_19789,N_17858,N_17276);
nand U19790 (N_19790,N_16576,N_17117);
or U19791 (N_19791,N_17980,N_17804);
nand U19792 (N_19792,N_16522,N_16026);
nand U19793 (N_19793,N_16421,N_17645);
nor U19794 (N_19794,N_16185,N_17150);
nor U19795 (N_19795,N_17903,N_17487);
and U19796 (N_19796,N_16718,N_16999);
nor U19797 (N_19797,N_17136,N_17405);
or U19798 (N_19798,N_17600,N_17995);
nor U19799 (N_19799,N_16636,N_16261);
nand U19800 (N_19800,N_17471,N_17855);
or U19801 (N_19801,N_16710,N_16355);
or U19802 (N_19802,N_16546,N_16126);
nor U19803 (N_19803,N_17333,N_16125);
xnor U19804 (N_19804,N_16243,N_17967);
or U19805 (N_19805,N_16523,N_17974);
and U19806 (N_19806,N_17607,N_17505);
nand U19807 (N_19807,N_16447,N_16813);
xor U19808 (N_19808,N_16054,N_17054);
and U19809 (N_19809,N_17141,N_16173);
or U19810 (N_19810,N_16787,N_17189);
xor U19811 (N_19811,N_17683,N_16250);
or U19812 (N_19812,N_16612,N_16849);
nand U19813 (N_19813,N_17130,N_17892);
nand U19814 (N_19814,N_17551,N_16675);
or U19815 (N_19815,N_16019,N_16705);
or U19816 (N_19816,N_17861,N_16678);
xor U19817 (N_19817,N_16818,N_16383);
or U19818 (N_19818,N_16030,N_17249);
and U19819 (N_19819,N_16265,N_17275);
nor U19820 (N_19820,N_16536,N_16015);
and U19821 (N_19821,N_17682,N_17052);
or U19822 (N_19822,N_17826,N_16749);
and U19823 (N_19823,N_17116,N_17638);
and U19824 (N_19824,N_16601,N_16737);
xor U19825 (N_19825,N_16930,N_16740);
or U19826 (N_19826,N_16524,N_17313);
or U19827 (N_19827,N_17644,N_16313);
xor U19828 (N_19828,N_17605,N_17381);
xor U19829 (N_19829,N_17280,N_16716);
xor U19830 (N_19830,N_16361,N_17305);
nand U19831 (N_19831,N_16385,N_16681);
nand U19832 (N_19832,N_17110,N_17932);
or U19833 (N_19833,N_16870,N_17388);
nand U19834 (N_19834,N_17015,N_16423);
nand U19835 (N_19835,N_16334,N_16899);
nand U19836 (N_19836,N_16421,N_16903);
and U19837 (N_19837,N_17983,N_17403);
or U19838 (N_19838,N_16479,N_16142);
xor U19839 (N_19839,N_17316,N_16049);
and U19840 (N_19840,N_17434,N_16542);
nand U19841 (N_19841,N_16994,N_17027);
nor U19842 (N_19842,N_16251,N_16214);
nand U19843 (N_19843,N_17183,N_17561);
xnor U19844 (N_19844,N_16657,N_17991);
and U19845 (N_19845,N_17838,N_17772);
nand U19846 (N_19846,N_17914,N_17777);
nor U19847 (N_19847,N_16581,N_16946);
nor U19848 (N_19848,N_17560,N_16114);
or U19849 (N_19849,N_16207,N_17973);
xnor U19850 (N_19850,N_16765,N_17623);
nand U19851 (N_19851,N_17032,N_17827);
nor U19852 (N_19852,N_16208,N_16868);
xor U19853 (N_19853,N_16105,N_16058);
or U19854 (N_19854,N_17873,N_17091);
nand U19855 (N_19855,N_17444,N_16744);
xor U19856 (N_19856,N_17277,N_16883);
nor U19857 (N_19857,N_17733,N_17041);
nand U19858 (N_19858,N_17160,N_16751);
and U19859 (N_19859,N_16702,N_17140);
and U19860 (N_19860,N_16546,N_17193);
xor U19861 (N_19861,N_16362,N_17727);
nand U19862 (N_19862,N_17271,N_16074);
nand U19863 (N_19863,N_16943,N_17236);
or U19864 (N_19864,N_16153,N_16837);
xor U19865 (N_19865,N_17148,N_17704);
nand U19866 (N_19866,N_17307,N_16343);
nand U19867 (N_19867,N_16944,N_17435);
nand U19868 (N_19868,N_16838,N_16356);
nand U19869 (N_19869,N_16615,N_17628);
xnor U19870 (N_19870,N_17471,N_17281);
nor U19871 (N_19871,N_16809,N_16178);
and U19872 (N_19872,N_17784,N_16389);
and U19873 (N_19873,N_16690,N_17522);
nor U19874 (N_19874,N_17614,N_16501);
xnor U19875 (N_19875,N_16224,N_17968);
or U19876 (N_19876,N_16946,N_16854);
or U19877 (N_19877,N_17286,N_16251);
nand U19878 (N_19878,N_17558,N_16757);
nand U19879 (N_19879,N_16691,N_17001);
nand U19880 (N_19880,N_16898,N_17265);
nor U19881 (N_19881,N_17410,N_16288);
nand U19882 (N_19882,N_17803,N_17382);
xor U19883 (N_19883,N_17463,N_17731);
nor U19884 (N_19884,N_16815,N_17988);
or U19885 (N_19885,N_17661,N_16511);
xor U19886 (N_19886,N_17882,N_16859);
and U19887 (N_19887,N_16475,N_17060);
and U19888 (N_19888,N_16541,N_16738);
xnor U19889 (N_19889,N_16984,N_16291);
and U19890 (N_19890,N_16037,N_17255);
nor U19891 (N_19891,N_16333,N_16858);
nor U19892 (N_19892,N_16947,N_16470);
and U19893 (N_19893,N_16264,N_17730);
or U19894 (N_19894,N_17933,N_17651);
xor U19895 (N_19895,N_17398,N_17150);
and U19896 (N_19896,N_16011,N_16005);
or U19897 (N_19897,N_16145,N_17633);
xor U19898 (N_19898,N_17661,N_16398);
nor U19899 (N_19899,N_17413,N_17601);
nand U19900 (N_19900,N_17625,N_16203);
nor U19901 (N_19901,N_16131,N_17193);
nor U19902 (N_19902,N_16149,N_17168);
or U19903 (N_19903,N_16920,N_17290);
nand U19904 (N_19904,N_17461,N_16973);
and U19905 (N_19905,N_17809,N_16359);
xor U19906 (N_19906,N_17971,N_16247);
xor U19907 (N_19907,N_16512,N_17785);
nor U19908 (N_19908,N_17652,N_17437);
or U19909 (N_19909,N_16461,N_17030);
xnor U19910 (N_19910,N_16622,N_17839);
nand U19911 (N_19911,N_17246,N_16160);
nand U19912 (N_19912,N_17825,N_17118);
and U19913 (N_19913,N_17559,N_17469);
xnor U19914 (N_19914,N_17499,N_17424);
xnor U19915 (N_19915,N_16246,N_17547);
or U19916 (N_19916,N_16812,N_16034);
nor U19917 (N_19917,N_16184,N_17371);
xnor U19918 (N_19918,N_16189,N_16415);
nor U19919 (N_19919,N_16064,N_16620);
nor U19920 (N_19920,N_17503,N_17370);
xor U19921 (N_19921,N_16862,N_16567);
nand U19922 (N_19922,N_17874,N_16535);
and U19923 (N_19923,N_17861,N_16247);
or U19924 (N_19924,N_17338,N_16767);
nor U19925 (N_19925,N_16211,N_17280);
nor U19926 (N_19926,N_17977,N_16767);
nor U19927 (N_19927,N_16034,N_16960);
or U19928 (N_19928,N_17790,N_16271);
nor U19929 (N_19929,N_17175,N_16870);
nor U19930 (N_19930,N_16306,N_16348);
nor U19931 (N_19931,N_17869,N_16553);
and U19932 (N_19932,N_16567,N_16067);
nor U19933 (N_19933,N_17453,N_16184);
nor U19934 (N_19934,N_16799,N_17344);
nand U19935 (N_19935,N_16426,N_17850);
xor U19936 (N_19936,N_17645,N_16410);
or U19937 (N_19937,N_17374,N_17160);
and U19938 (N_19938,N_17747,N_17866);
nand U19939 (N_19939,N_16185,N_16641);
or U19940 (N_19940,N_17568,N_16069);
nor U19941 (N_19941,N_16676,N_16349);
nor U19942 (N_19942,N_17257,N_17796);
nor U19943 (N_19943,N_17093,N_17673);
or U19944 (N_19944,N_16756,N_16889);
or U19945 (N_19945,N_17828,N_16801);
and U19946 (N_19946,N_17898,N_16660);
nand U19947 (N_19947,N_17945,N_16970);
nand U19948 (N_19948,N_17207,N_17646);
or U19949 (N_19949,N_16091,N_16110);
nand U19950 (N_19950,N_16806,N_16828);
or U19951 (N_19951,N_16803,N_17718);
nand U19952 (N_19952,N_16952,N_16999);
nand U19953 (N_19953,N_17426,N_17621);
or U19954 (N_19954,N_16476,N_16285);
nor U19955 (N_19955,N_17019,N_16978);
xor U19956 (N_19956,N_16225,N_16106);
or U19957 (N_19957,N_17553,N_17411);
or U19958 (N_19958,N_17036,N_16709);
and U19959 (N_19959,N_17828,N_16645);
nor U19960 (N_19960,N_16553,N_17527);
and U19961 (N_19961,N_16065,N_16993);
or U19962 (N_19962,N_17951,N_16329);
xor U19963 (N_19963,N_16627,N_17537);
xor U19964 (N_19964,N_17703,N_16818);
nor U19965 (N_19965,N_16700,N_17041);
nand U19966 (N_19966,N_17507,N_16305);
and U19967 (N_19967,N_17696,N_16950);
xnor U19968 (N_19968,N_17816,N_16539);
or U19969 (N_19969,N_16505,N_16647);
xor U19970 (N_19970,N_17881,N_17308);
xnor U19971 (N_19971,N_16629,N_17310);
xor U19972 (N_19972,N_17694,N_17506);
nor U19973 (N_19973,N_17531,N_17503);
nor U19974 (N_19974,N_16229,N_16177);
xor U19975 (N_19975,N_16555,N_16197);
xnor U19976 (N_19976,N_16212,N_17748);
nand U19977 (N_19977,N_16861,N_16224);
nand U19978 (N_19978,N_16140,N_17992);
xnor U19979 (N_19979,N_17850,N_16660);
nor U19980 (N_19980,N_17078,N_17593);
or U19981 (N_19981,N_17376,N_16430);
xor U19982 (N_19982,N_17364,N_17938);
xnor U19983 (N_19983,N_16251,N_16722);
or U19984 (N_19984,N_16700,N_16007);
nor U19985 (N_19985,N_17529,N_17685);
nand U19986 (N_19986,N_16656,N_16121);
nor U19987 (N_19987,N_16178,N_17772);
nand U19988 (N_19988,N_16893,N_17733);
xor U19989 (N_19989,N_16379,N_16046);
nor U19990 (N_19990,N_16672,N_17693);
or U19991 (N_19991,N_17552,N_17220);
nor U19992 (N_19992,N_16187,N_16164);
nor U19993 (N_19993,N_16119,N_17227);
and U19994 (N_19994,N_16678,N_16321);
or U19995 (N_19995,N_16765,N_17494);
nor U19996 (N_19996,N_17599,N_17665);
nor U19997 (N_19997,N_17781,N_17807);
xor U19998 (N_19998,N_16562,N_16835);
nor U19999 (N_19999,N_16665,N_17410);
nand UO_0 (O_0,N_19742,N_19896);
nand UO_1 (O_1,N_18585,N_19280);
or UO_2 (O_2,N_18021,N_18869);
nor UO_3 (O_3,N_18969,N_19974);
nor UO_4 (O_4,N_18277,N_19435);
nand UO_5 (O_5,N_19258,N_18828);
nand UO_6 (O_6,N_18194,N_18750);
nor UO_7 (O_7,N_19074,N_18690);
nor UO_8 (O_8,N_18444,N_19334);
nor UO_9 (O_9,N_18874,N_18863);
and UO_10 (O_10,N_18739,N_19541);
or UO_11 (O_11,N_18349,N_19807);
and UO_12 (O_12,N_18531,N_19458);
nor UO_13 (O_13,N_18421,N_18800);
nor UO_14 (O_14,N_19487,N_19219);
nand UO_15 (O_15,N_18077,N_18814);
or UO_16 (O_16,N_18078,N_18144);
xnor UO_17 (O_17,N_18150,N_19493);
nor UO_18 (O_18,N_18573,N_18908);
xnor UO_19 (O_19,N_19937,N_19430);
nor UO_20 (O_20,N_18528,N_19038);
xor UO_21 (O_21,N_19838,N_18075);
xor UO_22 (O_22,N_19893,N_19980);
nand UO_23 (O_23,N_19819,N_19369);
xor UO_24 (O_24,N_18061,N_18326);
or UO_25 (O_25,N_18020,N_18072);
nor UO_26 (O_26,N_18027,N_19264);
xor UO_27 (O_27,N_19717,N_18148);
or UO_28 (O_28,N_19946,N_19221);
and UO_29 (O_29,N_18871,N_19461);
or UO_30 (O_30,N_19877,N_18972);
or UO_31 (O_31,N_18909,N_19087);
and UO_32 (O_32,N_19216,N_18426);
nor UO_33 (O_33,N_18420,N_19993);
nand UO_34 (O_34,N_19881,N_19408);
or UO_35 (O_35,N_19339,N_18703);
nor UO_36 (O_36,N_18660,N_18847);
and UO_37 (O_37,N_19543,N_18130);
nand UO_38 (O_38,N_18255,N_19026);
and UO_39 (O_39,N_18396,N_18861);
nor UO_40 (O_40,N_19525,N_19640);
or UO_41 (O_41,N_19698,N_18720);
xnor UO_42 (O_42,N_18544,N_18032);
and UO_43 (O_43,N_19923,N_18128);
xnor UO_44 (O_44,N_19257,N_18285);
nand UO_45 (O_45,N_19224,N_18329);
nor UO_46 (O_46,N_18623,N_19996);
and UO_47 (O_47,N_19664,N_19758);
xor UO_48 (O_48,N_19020,N_19860);
xor UO_49 (O_49,N_18256,N_19774);
nand UO_50 (O_50,N_18701,N_18224);
and UO_51 (O_51,N_19791,N_18533);
or UO_52 (O_52,N_18133,N_18944);
nor UO_53 (O_53,N_18007,N_19126);
and UO_54 (O_54,N_19093,N_19494);
or UO_55 (O_55,N_18577,N_18580);
nand UO_56 (O_56,N_18024,N_18629);
nor UO_57 (O_57,N_19009,N_19704);
nor UO_58 (O_58,N_18473,N_19943);
nor UO_59 (O_59,N_19713,N_18292);
nor UO_60 (O_60,N_18608,N_18073);
or UO_61 (O_61,N_19315,N_19155);
and UO_62 (O_62,N_18672,N_18220);
or UO_63 (O_63,N_18671,N_18803);
or UO_64 (O_64,N_18272,N_18715);
or UO_65 (O_65,N_18118,N_18653);
or UO_66 (O_66,N_18113,N_18914);
nand UO_67 (O_67,N_18764,N_18813);
nand UO_68 (O_68,N_19086,N_19331);
and UO_69 (O_69,N_19184,N_18700);
xnor UO_70 (O_70,N_19965,N_18460);
nand UO_71 (O_71,N_19231,N_19612);
nor UO_72 (O_72,N_19687,N_19410);
xnor UO_73 (O_73,N_19803,N_19659);
and UO_74 (O_74,N_19981,N_19969);
xnor UO_75 (O_75,N_18947,N_19622);
xnor UO_76 (O_76,N_19646,N_18534);
xor UO_77 (O_77,N_19685,N_19380);
nand UO_78 (O_78,N_19457,N_18584);
and UO_79 (O_79,N_19507,N_19144);
xnor UO_80 (O_80,N_18393,N_19871);
and UO_81 (O_81,N_18778,N_19284);
or UO_82 (O_82,N_19736,N_19043);
and UO_83 (O_83,N_18797,N_19962);
nand UO_84 (O_84,N_19729,N_18890);
or UO_85 (O_85,N_18465,N_19347);
nand UO_86 (O_86,N_18180,N_18645);
xor UO_87 (O_87,N_19689,N_18003);
or UO_88 (O_88,N_18517,N_19474);
or UO_89 (O_89,N_19952,N_18755);
or UO_90 (O_90,N_18789,N_18074);
or UO_91 (O_91,N_18265,N_19185);
and UO_92 (O_92,N_18012,N_19137);
nor UO_93 (O_93,N_19630,N_19957);
or UO_94 (O_94,N_18605,N_19773);
or UO_95 (O_95,N_18897,N_18681);
xor UO_96 (O_96,N_18160,N_19124);
nand UO_97 (O_97,N_19683,N_19175);
xnor UO_98 (O_98,N_19145,N_19915);
nor UO_99 (O_99,N_18390,N_19436);
nor UO_100 (O_100,N_19480,N_19628);
nand UO_101 (O_101,N_18793,N_19478);
or UO_102 (O_102,N_18397,N_18450);
and UO_103 (O_103,N_19608,N_19207);
or UO_104 (O_104,N_18731,N_19629);
or UO_105 (O_105,N_19186,N_18938);
nand UO_106 (O_106,N_18615,N_18518);
and UO_107 (O_107,N_18056,N_18172);
nand UO_108 (O_108,N_19036,N_19739);
and UO_109 (O_109,N_18999,N_19007);
nand UO_110 (O_110,N_18772,N_18419);
nor UO_111 (O_111,N_18880,N_18208);
nor UO_112 (O_112,N_19463,N_19577);
nor UO_113 (O_113,N_18744,N_19308);
xnor UO_114 (O_114,N_19741,N_19572);
xnor UO_115 (O_115,N_18187,N_18207);
or UO_116 (O_116,N_19076,N_19547);
nand UO_117 (O_117,N_19336,N_18347);
nor UO_118 (O_118,N_18722,N_18483);
and UO_119 (O_119,N_19085,N_19502);
nand UO_120 (O_120,N_18066,N_18173);
and UO_121 (O_121,N_18181,N_19989);
or UO_122 (O_122,N_19808,N_18447);
xor UO_123 (O_123,N_18787,N_18891);
nand UO_124 (O_124,N_18649,N_19508);
and UO_125 (O_125,N_19010,N_18721);
xor UO_126 (O_126,N_18964,N_18399);
xor UO_127 (O_127,N_19355,N_18226);
and UO_128 (O_128,N_19288,N_18348);
nor UO_129 (O_129,N_19305,N_18037);
or UO_130 (O_130,N_19912,N_19814);
or UO_131 (O_131,N_18009,N_18284);
nand UO_132 (O_132,N_19266,N_19101);
nand UO_133 (O_133,N_18433,N_18994);
or UO_134 (O_134,N_18484,N_18271);
nor UO_135 (O_135,N_18067,N_19829);
or UO_136 (O_136,N_18951,N_18146);
nand UO_137 (O_137,N_19413,N_19575);
and UO_138 (O_138,N_18586,N_19559);
nand UO_139 (O_139,N_18087,N_19156);
or UO_140 (O_140,N_18238,N_19617);
xor UO_141 (O_141,N_19850,N_18109);
and UO_142 (O_142,N_18103,N_19165);
and UO_143 (O_143,N_19634,N_18136);
nand UO_144 (O_144,N_19290,N_18634);
xnor UO_145 (O_145,N_18263,N_19389);
and UO_146 (O_146,N_19166,N_18598);
xor UO_147 (O_147,N_19187,N_19585);
xor UO_148 (O_148,N_19821,N_18082);
and UO_149 (O_149,N_19652,N_18134);
nand UO_150 (O_150,N_18051,N_19695);
nor UO_151 (O_151,N_18918,N_18990);
and UO_152 (O_152,N_18788,N_19482);
nand UO_153 (O_153,N_18572,N_18495);
xor UO_154 (O_154,N_18449,N_19747);
and UO_155 (O_155,N_19274,N_18817);
xor UO_156 (O_156,N_18478,N_18986);
nand UO_157 (O_157,N_18221,N_18808);
nand UO_158 (O_158,N_18178,N_19263);
nor UO_159 (O_159,N_19265,N_19591);
nand UO_160 (O_160,N_19568,N_18727);
and UO_161 (O_161,N_18291,N_18795);
nor UO_162 (O_162,N_18818,N_18462);
xor UO_163 (O_163,N_19095,N_18406);
xor UO_164 (O_164,N_19599,N_18838);
or UO_165 (O_165,N_19040,N_19109);
or UO_166 (O_166,N_19498,N_19826);
nor UO_167 (O_167,N_19781,N_19812);
nor UO_168 (O_168,N_18378,N_18699);
and UO_169 (O_169,N_19354,N_19914);
xor UO_170 (O_170,N_18163,N_18697);
or UO_171 (O_171,N_19986,N_19909);
or UO_172 (O_172,N_19611,N_19842);
xor UO_173 (O_173,N_18153,N_19365);
xnor UO_174 (O_174,N_19471,N_19540);
nor UO_175 (O_175,N_19327,N_18923);
and UO_176 (O_176,N_18568,N_18843);
and UO_177 (O_177,N_19149,N_19926);
xor UO_178 (O_178,N_19000,N_19726);
xnor UO_179 (O_179,N_18602,N_19861);
and UO_180 (O_180,N_18987,N_19035);
and UO_181 (O_181,N_19970,N_18210);
and UO_182 (O_182,N_18139,N_19245);
nand UO_183 (O_183,N_19961,N_18415);
or UO_184 (O_184,N_19021,N_18611);
nor UO_185 (O_185,N_18101,N_19472);
nand UO_186 (O_186,N_18283,N_19875);
nor UO_187 (O_187,N_19374,N_19564);
and UO_188 (O_188,N_18939,N_18563);
or UO_189 (O_189,N_19900,N_19431);
nor UO_190 (O_190,N_19138,N_19849);
nand UO_191 (O_191,N_18053,N_19546);
or UO_192 (O_192,N_19379,N_19091);
nor UO_193 (O_193,N_18966,N_18320);
xnor UO_194 (O_194,N_19223,N_18867);
nor UO_195 (O_195,N_19837,N_18827);
and UO_196 (O_196,N_18313,N_19582);
nand UO_197 (O_197,N_19998,N_18617);
xnor UO_198 (O_198,N_19637,N_19392);
and UO_199 (O_199,N_18676,N_18556);
xnor UO_200 (O_200,N_19159,N_19314);
nand UO_201 (O_201,N_19295,N_19642);
nor UO_202 (O_202,N_18636,N_18840);
nor UO_203 (O_203,N_19051,N_18363);
nor UO_204 (O_204,N_19309,N_19154);
nor UO_205 (O_205,N_19343,N_18273);
or UO_206 (O_206,N_18935,N_19852);
xor UO_207 (O_207,N_18331,N_18176);
nand UO_208 (O_208,N_19885,N_18562);
and UO_209 (O_209,N_18658,N_19506);
xor UO_210 (O_210,N_19460,N_18748);
or UO_211 (O_211,N_18068,N_19658);
nand UO_212 (O_212,N_19005,N_19025);
nand UO_213 (O_213,N_18622,N_18796);
and UO_214 (O_214,N_18765,N_18167);
and UO_215 (O_215,N_19358,N_18976);
or UO_216 (O_216,N_19356,N_18166);
nand UO_217 (O_217,N_18461,N_19703);
xor UO_218 (O_218,N_18306,N_18143);
xnor UO_219 (O_219,N_18512,N_18807);
nand UO_220 (O_220,N_18707,N_18403);
xor UO_221 (O_221,N_19718,N_19121);
and UO_222 (O_222,N_19886,N_19954);
nor UO_223 (O_223,N_19740,N_18309);
and UO_224 (O_224,N_18782,N_18673);
or UO_225 (O_225,N_19409,N_19252);
xor UO_226 (O_226,N_18576,N_19345);
and UO_227 (O_227,N_18930,N_18488);
or UO_228 (O_228,N_19968,N_19694);
and UO_229 (O_229,N_19473,N_19368);
nand UO_230 (O_230,N_18040,N_19161);
nand UO_231 (O_231,N_19535,N_18417);
or UO_232 (O_232,N_19213,N_19673);
nand UO_233 (O_233,N_18757,N_19884);
or UO_234 (O_234,N_19462,N_19329);
nor UO_235 (O_235,N_19423,N_19247);
and UO_236 (O_236,N_18380,N_19254);
xnor UO_237 (O_237,N_19128,N_18299);
and UO_238 (O_238,N_19384,N_19242);
and UO_239 (O_239,N_18937,N_19847);
and UO_240 (O_240,N_19895,N_19300);
xor UO_241 (O_241,N_19555,N_19933);
or UO_242 (O_242,N_18804,N_18260);
nor UO_243 (O_243,N_19032,N_19483);
or UO_244 (O_244,N_18195,N_19854);
xnor UO_245 (O_245,N_18206,N_19516);
nor UO_246 (O_246,N_19130,N_18785);
and UO_247 (O_247,N_18307,N_19169);
nor UO_248 (O_248,N_18995,N_19378);
nand UO_249 (O_249,N_18057,N_18039);
xnor UO_250 (O_250,N_19140,N_19283);
and UO_251 (O_251,N_19271,N_18669);
nor UO_252 (O_252,N_19267,N_18469);
nor UO_253 (O_253,N_18247,N_19668);
or UO_254 (O_254,N_19545,N_19214);
nor UO_255 (O_255,N_19839,N_18416);
xnor UO_256 (O_256,N_18910,N_19988);
xnor UO_257 (O_257,N_18508,N_18546);
xnor UO_258 (O_258,N_19304,N_18940);
nand UO_259 (O_259,N_19621,N_19602);
xor UO_260 (O_260,N_19299,N_18760);
xor UO_261 (O_261,N_19565,N_19235);
and UO_262 (O_262,N_18866,N_18504);
nand UO_263 (O_263,N_18409,N_19678);
xor UO_264 (O_264,N_18670,N_18718);
or UO_265 (O_265,N_19879,N_19313);
nor UO_266 (O_266,N_19874,N_19061);
and UO_267 (O_267,N_19205,N_19147);
and UO_268 (O_268,N_18975,N_19561);
or UO_269 (O_269,N_18879,N_18705);
xnor UO_270 (O_270,N_19671,N_18366);
nor UO_271 (O_271,N_18745,N_18296);
and UO_272 (O_272,N_18250,N_18810);
xnor UO_273 (O_273,N_18829,N_19292);
or UO_274 (O_274,N_18565,N_19665);
and UO_275 (O_275,N_18844,N_18475);
and UO_276 (O_276,N_19576,N_18405);
and UO_277 (O_277,N_18657,N_19232);
nor UO_278 (O_278,N_18689,N_19350);
nor UO_279 (O_279,N_18732,N_18759);
or UO_280 (O_280,N_19054,N_18316);
nand UO_281 (O_281,N_19201,N_18900);
and UO_282 (O_282,N_19008,N_18656);
nor UO_283 (O_283,N_18708,N_18446);
xnor UO_284 (O_284,N_18062,N_18245);
nand UO_285 (O_285,N_18973,N_18198);
xnor UO_286 (O_286,N_18384,N_18594);
nand UO_287 (O_287,N_18980,N_18996);
nand UO_288 (O_288,N_18823,N_19769);
or UO_289 (O_289,N_18152,N_18613);
nor UO_290 (O_290,N_19361,N_18158);
and UO_291 (O_291,N_19444,N_19189);
nor UO_292 (O_292,N_18984,N_18625);
xnor UO_293 (O_293,N_18780,N_19820);
xor UO_294 (O_294,N_19167,N_19604);
nor UO_295 (O_295,N_18826,N_19790);
nand UO_296 (O_296,N_19238,N_19112);
and UO_297 (O_297,N_18303,N_18375);
or UO_298 (O_298,N_19386,N_19873);
xnor UO_299 (O_299,N_18955,N_19479);
xnor UO_300 (O_300,N_18237,N_18680);
nand UO_301 (O_301,N_19596,N_18928);
or UO_302 (O_302,N_18411,N_18100);
or UO_303 (O_303,N_19901,N_19484);
or UO_304 (O_304,N_19544,N_18507);
nor UO_305 (O_305,N_18125,N_18408);
nor UO_306 (O_306,N_18942,N_19806);
or UO_307 (O_307,N_19690,N_19768);
or UO_308 (O_308,N_18184,N_19794);
or UO_309 (O_309,N_18836,N_19089);
nor UO_310 (O_310,N_19397,N_19367);
nand UO_311 (O_311,N_18242,N_18216);
and UO_312 (O_312,N_18775,N_19796);
or UO_313 (O_313,N_18333,N_18948);
nor UO_314 (O_314,N_18609,N_19759);
or UO_315 (O_315,N_19600,N_19615);
and UO_316 (O_316,N_19524,N_18186);
and UO_317 (O_317,N_18025,N_19904);
xor UO_318 (O_318,N_18542,N_19276);
xnor UO_319 (O_319,N_18227,N_19571);
xor UO_320 (O_320,N_19691,N_18898);
xor UO_321 (O_321,N_19783,N_19919);
and UO_322 (O_322,N_19653,N_18941);
or UO_323 (O_323,N_18281,N_18054);
or UO_324 (O_324,N_18683,N_19994);
and UO_325 (O_325,N_19542,N_18773);
xnor UO_326 (O_326,N_19370,N_19279);
nand UO_327 (O_327,N_18805,N_18425);
nand UO_328 (O_328,N_19991,N_18820);
or UO_329 (O_329,N_19083,N_19509);
xor UO_330 (O_330,N_19210,N_19754);
xor UO_331 (O_331,N_18906,N_18394);
or UO_332 (O_332,N_19017,N_18357);
and UO_333 (O_333,N_19046,N_19757);
and UO_334 (O_334,N_18870,N_18257);
nor UO_335 (O_335,N_19711,N_19940);
and UO_336 (O_336,N_19644,N_18515);
nor UO_337 (O_337,N_19027,N_19699);
xnor UO_338 (O_338,N_18259,N_18005);
xnor UO_339 (O_339,N_19340,N_19053);
or UO_340 (O_340,N_18477,N_18322);
nor UO_341 (O_341,N_19779,N_19323);
and UO_342 (O_342,N_19725,N_18058);
nor UO_343 (O_343,N_18630,N_18115);
nor UO_344 (O_344,N_19139,N_19448);
and UO_345 (O_345,N_18754,N_18350);
xnor UO_346 (O_346,N_19995,N_18261);
or UO_347 (O_347,N_19118,N_18571);
and UO_348 (O_348,N_19955,N_19770);
or UO_349 (O_349,N_19499,N_18457);
or UO_350 (O_350,N_18330,N_18233);
nand UO_351 (O_351,N_18361,N_19402);
and UO_352 (O_352,N_18126,N_19823);
and UO_353 (O_353,N_19262,N_19424);
nor UO_354 (O_354,N_18949,N_19212);
nand UO_355 (O_355,N_18076,N_18922);
xnor UO_356 (O_356,N_18885,N_19960);
and UO_357 (O_357,N_19168,N_19335);
xor UO_358 (O_358,N_18497,N_18816);
xor UO_359 (O_359,N_19490,N_18323);
and UO_360 (O_360,N_18926,N_19024);
nand UO_361 (O_361,N_19714,N_19579);
nor UO_362 (O_362,N_18493,N_18693);
and UO_363 (O_363,N_19048,N_18480);
or UO_364 (O_364,N_19391,N_18346);
nor UO_365 (O_365,N_18831,N_18451);
nand UO_366 (O_366,N_19916,N_18050);
or UO_367 (O_367,N_19897,N_19601);
nor UO_368 (O_368,N_18383,N_19778);
and UO_369 (O_369,N_19657,N_18977);
nor UO_370 (O_370,N_19716,N_18097);
nand UO_371 (O_371,N_19488,N_18726);
xnor UO_372 (O_372,N_18919,N_18519);
and UO_373 (O_373,N_18790,N_18716);
or UO_374 (O_374,N_18501,N_19105);
nand UO_375 (O_375,N_18231,N_18654);
and UO_376 (O_376,N_19734,N_18679);
nor UO_377 (O_377,N_18243,N_19286);
or UO_378 (O_378,N_18205,N_19037);
nor UO_379 (O_379,N_18249,N_18254);
nand UO_380 (O_380,N_19018,N_19889);
or UO_381 (O_381,N_19684,N_19928);
nand UO_382 (O_382,N_18318,N_18762);
xor UO_383 (O_383,N_18448,N_18217);
and UO_384 (O_384,N_18356,N_18138);
or UO_385 (O_385,N_18612,N_18899);
xnor UO_386 (O_386,N_18777,N_19505);
nand UO_387 (O_387,N_19194,N_19202);
or UO_388 (O_388,N_19294,N_19193);
and UO_389 (O_389,N_18616,N_18567);
nand UO_390 (O_390,N_18621,N_19459);
nand UO_391 (O_391,N_19447,N_18557);
or UO_392 (O_392,N_19296,N_18767);
and UO_393 (O_393,N_19641,N_18514);
and UO_394 (O_394,N_19563,N_19532);
or UO_395 (O_395,N_18694,N_19939);
and UO_396 (O_396,N_19016,N_18859);
xor UO_397 (O_397,N_18441,N_19815);
nor UO_398 (O_398,N_19844,N_18344);
nor UO_399 (O_399,N_18099,N_18107);
nor UO_400 (O_400,N_18098,N_19110);
nand UO_401 (O_401,N_19765,N_18015);
or UO_402 (O_402,N_19869,N_19631);
nor UO_403 (O_403,N_19133,N_19209);
or UO_404 (O_404,N_19945,N_19570);
nand UO_405 (O_405,N_18029,N_18338);
nor UO_406 (O_406,N_19775,N_19382);
xnor UO_407 (O_407,N_19708,N_18578);
xnor UO_408 (O_408,N_19148,N_19744);
nor UO_409 (O_409,N_18596,N_18456);
and UO_410 (O_410,N_18848,N_18925);
or UO_411 (O_411,N_19530,N_18304);
and UO_412 (O_412,N_18644,N_18687);
nor UO_413 (O_413,N_19619,N_18505);
nand UO_414 (O_414,N_19060,N_18791);
nor UO_415 (O_415,N_18155,N_19648);
or UO_416 (O_416,N_19371,N_19115);
and UO_417 (O_417,N_18806,N_19317);
nor UO_418 (O_418,N_19075,N_18963);
and UO_419 (O_419,N_18655,N_19249);
nand UO_420 (O_420,N_19297,N_18606);
and UO_421 (O_421,N_19104,N_18122);
and UO_422 (O_422,N_18641,N_19364);
nor UO_423 (O_423,N_18704,N_19143);
nor UO_424 (O_424,N_18174,N_19415);
nor UO_425 (O_425,N_19578,N_19191);
and UO_426 (O_426,N_18300,N_18714);
nand UO_427 (O_427,N_19050,N_18862);
and UO_428 (O_428,N_19446,N_18539);
nand UO_429 (O_429,N_19131,N_18903);
xor UO_430 (O_430,N_19261,N_18482);
and UO_431 (O_431,N_18141,N_19750);
xnor UO_432 (O_432,N_18197,N_19129);
xnor UO_433 (O_433,N_18834,N_18353);
and UO_434 (O_434,N_18802,N_18873);
and UO_435 (O_435,N_19015,N_18631);
and UO_436 (O_436,N_18302,N_19738);
or UO_437 (O_437,N_18581,N_18579);
nor UO_438 (O_438,N_19751,N_18439);
and UO_439 (O_439,N_18496,N_19905);
nor UO_440 (O_440,N_18467,N_18023);
and UO_441 (O_441,N_18758,N_18525);
nor UO_442 (O_442,N_19971,N_19562);
and UO_443 (O_443,N_19181,N_19301);
and UO_444 (O_444,N_19127,N_18494);
nand UO_445 (O_445,N_18920,N_19422);
and UO_446 (O_446,N_19306,N_19743);
and UO_447 (O_447,N_19650,N_19513);
xor UO_448 (O_448,N_18997,N_18583);
or UO_449 (O_449,N_18845,N_19515);
nor UO_450 (O_450,N_19825,N_18341);
nand UO_451 (O_451,N_19863,N_19855);
or UO_452 (O_452,N_19200,N_19256);
or UO_453 (O_453,N_18855,N_19589);
and UO_454 (O_454,N_19913,N_18552);
and UO_455 (O_455,N_18487,N_18466);
or UO_456 (O_456,N_19157,N_19872);
nand UO_457 (O_457,N_19399,N_19425);
xnor UO_458 (O_458,N_18559,N_18607);
xor UO_459 (O_459,N_18004,N_18096);
xor UO_460 (O_460,N_19470,N_19476);
nor UO_461 (O_461,N_19377,N_19938);
xnor UO_462 (O_462,N_18352,N_18854);
nand UO_463 (O_463,N_18886,N_19966);
or UO_464 (O_464,N_19272,N_19344);
xor UO_465 (O_465,N_19330,N_19116);
xor UO_466 (O_466,N_18114,N_18763);
xnor UO_467 (O_467,N_18248,N_19693);
or UO_468 (O_468,N_19067,N_18124);
nor UO_469 (O_469,N_18002,N_19163);
or UO_470 (O_470,N_19722,N_19248);
nand UO_471 (O_471,N_19643,N_19942);
nor UO_472 (O_472,N_18933,N_19792);
nand UO_473 (O_473,N_19174,N_18913);
nand UO_474 (O_474,N_19927,N_18016);
xnor UO_475 (O_475,N_19676,N_19848);
nor UO_476 (O_476,N_19526,N_19132);
nor UO_477 (O_477,N_19723,N_19092);
and UO_478 (O_478,N_19022,N_19903);
nand UO_479 (O_479,N_19443,N_18684);
nand UO_480 (O_480,N_19100,N_18236);
nand UO_481 (O_481,N_18189,N_18036);
nand UO_482 (O_482,N_18747,N_18998);
nor UO_483 (O_483,N_18358,N_18355);
or UO_484 (O_484,N_19353,N_18083);
or UO_485 (O_485,N_19059,N_18490);
or UO_486 (O_486,N_18882,N_19956);
nand UO_487 (O_487,N_19857,N_19537);
nor UO_488 (O_488,N_18725,N_18332);
and UO_489 (O_489,N_18799,N_18373);
or UO_490 (O_490,N_18218,N_18841);
nor UO_491 (O_491,N_19931,N_19211);
nor UO_492 (O_492,N_19574,N_19780);
and UO_493 (O_493,N_19357,N_18137);
or UO_494 (O_494,N_19992,N_19660);
xor UO_495 (O_495,N_19491,N_18713);
nor UO_496 (O_496,N_19772,N_19303);
nor UO_497 (O_497,N_18988,N_18442);
and UO_498 (O_498,N_19395,N_18968);
and UO_499 (O_499,N_18811,N_19834);
and UO_500 (O_500,N_19222,N_18824);
and UO_501 (O_501,N_19649,N_19289);
nor UO_502 (O_502,N_18190,N_19947);
nor UO_503 (O_503,N_19598,N_18298);
nor UO_504 (O_504,N_18749,N_19049);
or UO_505 (O_505,N_18674,N_19228);
and UO_506 (O_506,N_19039,N_18069);
xor UO_507 (O_507,N_19681,N_18117);
xor UO_508 (O_508,N_18499,N_19707);
nor UO_509 (O_509,N_19669,N_18251);
or UO_510 (O_510,N_19625,N_19103);
xor UO_511 (O_511,N_18709,N_19071);
nand UO_512 (O_512,N_18258,N_19466);
nor UO_513 (O_513,N_19702,N_18093);
xnor UO_514 (O_514,N_18364,N_19534);
xor UO_515 (O_515,N_18500,N_19097);
nand UO_516 (O_516,N_19811,N_18177);
or UO_517 (O_517,N_19456,N_18809);
or UO_518 (O_518,N_18957,N_19113);
nor UO_519 (O_519,N_18381,N_18554);
or UO_520 (O_520,N_19822,N_19805);
nor UO_521 (O_521,N_19924,N_19023);
xor UO_522 (O_522,N_18424,N_19220);
nand UO_523 (O_523,N_19120,N_19106);
nand UO_524 (O_524,N_19529,N_19063);
xor UO_525 (O_525,N_19412,N_18821);
nor UO_526 (O_526,N_18215,N_18904);
nor UO_527 (O_527,N_19003,N_19146);
xor UO_528 (O_528,N_18407,N_18502);
and UO_529 (O_529,N_19733,N_19042);
nand UO_530 (O_530,N_19705,N_19153);
nor UO_531 (O_531,N_19477,N_18603);
and UO_532 (O_532,N_19094,N_18929);
or UO_533 (O_533,N_18429,N_19922);
or UO_534 (O_534,N_18084,N_19251);
nor UO_535 (O_535,N_18413,N_18287);
and UO_536 (O_536,N_19566,N_18045);
or UO_537 (O_537,N_18812,N_18856);
or UO_538 (O_538,N_19514,N_19004);
xor UO_539 (O_539,N_19311,N_19799);
nor UO_540 (O_540,N_18706,N_18839);
xor UO_541 (O_541,N_18030,N_18464);
nor UO_542 (O_542,N_19917,N_19581);
and UO_543 (O_543,N_19162,N_19797);
nor UO_544 (O_544,N_18401,N_19700);
and UO_545 (O_545,N_18746,N_19760);
nor UO_546 (O_546,N_18468,N_19013);
or UO_547 (O_547,N_18648,N_19033);
nand UO_548 (O_548,N_19259,N_18647);
nand UO_549 (O_549,N_19936,N_19123);
nand UO_550 (O_550,N_18454,N_19429);
nand UO_551 (O_551,N_18604,N_18325);
nor UO_552 (O_552,N_19244,N_18883);
xor UO_553 (O_553,N_18006,N_18327);
and UO_554 (O_554,N_18819,N_18288);
nor UO_555 (O_555,N_19107,N_18048);
xor UO_556 (O_556,N_18314,N_19645);
or UO_557 (O_557,N_19859,N_19417);
and UO_558 (O_558,N_18328,N_19072);
nor UO_559 (O_559,N_19197,N_19972);
nand UO_560 (O_560,N_19045,N_18774);
nand UO_561 (O_561,N_19178,N_18723);
xor UO_562 (O_562,N_18428,N_18530);
and UO_563 (O_563,N_18538,N_19554);
or UO_564 (O_564,N_19287,N_18440);
and UO_565 (O_565,N_19930,N_19420);
or UO_566 (O_566,N_18147,N_19932);
and UO_567 (O_567,N_18872,N_18792);
or UO_568 (O_568,N_18289,N_18768);
xnor UO_569 (O_569,N_19275,N_19481);
xnor UO_570 (O_570,N_18209,N_19270);
nand UO_571 (O_571,N_19426,N_18169);
nand UO_572 (O_572,N_18239,N_18060);
and UO_573 (O_573,N_19260,N_18640);
nor UO_574 (O_574,N_18479,N_18212);
or UO_575 (O_575,N_19941,N_18574);
nand UO_576 (O_576,N_19503,N_18085);
nor UO_577 (O_577,N_19549,N_18183);
nor UO_578 (O_578,N_19073,N_19504);
xor UO_579 (O_579,N_18887,N_18985);
or UO_580 (O_580,N_19082,N_19605);
or UO_581 (O_581,N_18865,N_18367);
nor UO_582 (O_582,N_19332,N_18540);
xnor UO_583 (O_583,N_19558,N_19677);
and UO_584 (O_584,N_18950,N_19858);
or UO_585 (O_585,N_19099,N_18779);
or UO_586 (O_586,N_19666,N_18526);
nand UO_587 (O_587,N_18896,N_18761);
and UO_588 (O_588,N_19553,N_18894);
nand UO_589 (O_589,N_19366,N_19647);
and UO_590 (O_590,N_18907,N_19728);
or UO_591 (O_591,N_19285,N_19620);
or UO_592 (O_592,N_19298,N_18014);
and UO_593 (O_593,N_18776,N_19550);
or UO_594 (O_594,N_19243,N_19512);
nand UO_595 (O_595,N_18850,N_18619);
nand UO_596 (O_596,N_19080,N_18597);
nor UO_597 (O_597,N_18982,N_19019);
or UO_598 (O_598,N_19468,N_18498);
nor UO_599 (O_599,N_18295,N_19177);
or UO_600 (O_600,N_18228,N_18527);
nor UO_601 (O_601,N_18359,N_19326);
xor UO_602 (O_602,N_19438,N_18610);
nand UO_603 (O_603,N_18080,N_18222);
nand UO_604 (O_604,N_18091,N_19328);
and UO_605 (O_605,N_18422,N_19679);
and UO_606 (O_606,N_18244,N_19795);
nand UO_607 (O_607,N_19065,N_18520);
nor UO_608 (O_608,N_18362,N_18864);
or UO_609 (O_609,N_18614,N_18529);
xnor UO_610 (O_610,N_18635,N_19119);
or UO_611 (O_611,N_19675,N_18756);
or UO_612 (O_612,N_19437,N_19788);
or UO_613 (O_613,N_19727,N_18695);
nor UO_614 (O_614,N_19958,N_19890);
or UO_615 (O_615,N_18842,N_18801);
nor UO_616 (O_616,N_19845,N_18967);
and UO_617 (O_617,N_18503,N_19748);
nand UO_618 (O_618,N_19052,N_19831);
and UO_619 (O_619,N_19777,N_19749);
xor UO_620 (O_620,N_18652,N_19766);
or UO_621 (O_621,N_18161,N_18550);
xnor UO_622 (O_622,N_19755,N_18590);
xor UO_623 (O_623,N_19567,N_18431);
nand UO_624 (O_624,N_18875,N_19518);
xnor UO_625 (O_625,N_19030,N_18324);
nor UO_626 (O_626,N_19626,N_19548);
and UO_627 (O_627,N_19055,N_18561);
and UO_628 (O_628,N_18743,N_18962);
or UO_629 (O_629,N_18017,N_18524);
or UO_630 (O_630,N_19686,N_19179);
nor UO_631 (O_631,N_19293,N_19282);
or UO_632 (O_632,N_18193,N_18019);
xor UO_633 (O_633,N_18001,N_19523);
xor UO_634 (O_634,N_18102,N_19894);
xnor UO_635 (O_635,N_18666,N_18786);
and UO_636 (O_636,N_19983,N_19712);
nand UO_637 (O_637,N_18593,N_19102);
xor UO_638 (O_638,N_19624,N_19160);
or UO_639 (O_639,N_19934,N_19719);
and UO_640 (O_640,N_18665,N_18889);
nand UO_641 (O_641,N_18135,N_19569);
or UO_642 (O_642,N_19419,N_19451);
xor UO_643 (O_643,N_18551,N_18698);
nor UO_644 (O_644,N_19173,N_18981);
nor UO_645 (O_645,N_19188,N_18427);
and UO_646 (O_646,N_19882,N_19737);
nor UO_647 (O_647,N_18165,N_18418);
nor UO_648 (O_648,N_19830,N_18934);
xnor UO_649 (O_649,N_18382,N_18691);
or UO_650 (O_650,N_19950,N_19069);
and UO_651 (O_651,N_18110,N_19635);
xor UO_652 (O_652,N_19590,N_18031);
xnor UO_653 (O_653,N_18204,N_18119);
nand UO_654 (O_654,N_19661,N_18591);
xor UO_655 (O_655,N_19172,N_18878);
nor UO_656 (O_656,N_18742,N_19898);
xnor UO_657 (O_657,N_18010,N_18589);
xnor UO_658 (O_658,N_19697,N_18034);
or UO_659 (O_659,N_18489,N_19501);
nand UO_660 (O_660,N_18917,N_18191);
or UO_661 (O_661,N_18835,N_19454);
xnor UO_662 (O_662,N_18784,N_18664);
xor UO_663 (O_663,N_18340,N_18595);
nor UO_664 (O_664,N_19006,N_19521);
or UO_665 (O_665,N_18989,N_19720);
nand UO_666 (O_666,N_19891,N_19312);
xor UO_667 (O_667,N_19203,N_18131);
nand UO_668 (O_668,N_19592,N_19465);
xor UO_669 (O_669,N_19014,N_19012);
and UO_670 (O_670,N_18046,N_19843);
or UO_671 (O_671,N_18545,N_18815);
or UO_672 (O_672,N_18092,N_19856);
nand UO_673 (O_673,N_18719,N_19056);
xnor UO_674 (O_674,N_18912,N_19226);
nand UO_675 (O_675,N_18430,N_19064);
nand UO_676 (O_676,N_18476,N_19176);
and UO_677 (O_677,N_18132,N_18452);
or UO_678 (O_678,N_18443,N_18319);
nand UO_679 (O_679,N_19682,N_19835);
and UO_680 (O_680,N_18280,N_19784);
xor UO_681 (O_681,N_19321,N_19497);
and UO_682 (O_682,N_19170,N_18857);
xnor UO_683 (O_683,N_19892,N_19606);
or UO_684 (O_684,N_19414,N_18753);
nand UO_685 (O_685,N_18895,N_19840);
nand UO_686 (O_686,N_18293,N_18171);
nand UO_687 (O_687,N_18678,N_18662);
or UO_688 (O_688,N_18954,N_19616);
nor UO_689 (O_689,N_18404,N_19587);
xnor UO_690 (O_690,N_18628,N_18783);
and UO_691 (O_691,N_18992,N_19352);
nor UO_692 (O_692,N_19959,N_19519);
and UO_693 (O_693,N_18633,N_19763);
and UO_694 (O_694,N_19973,N_19029);
nand UO_695 (O_695,N_18156,N_18414);
xnor UO_696 (O_696,N_18435,N_18129);
xnor UO_697 (O_697,N_18639,N_19632);
or UO_698 (O_698,N_19654,N_19320);
xor UO_699 (O_699,N_18537,N_19908);
nand UO_700 (O_700,N_19469,N_18979);
nand UO_701 (O_701,N_19918,N_19250);
nor UO_702 (O_702,N_18470,N_19237);
nand UO_703 (O_703,N_18916,N_18696);
nand UO_704 (O_704,N_19911,N_18047);
nand UO_705 (O_705,N_19977,N_18710);
nor UO_706 (O_706,N_18423,N_18884);
nor UO_707 (O_707,N_19584,N_19230);
or UO_708 (O_708,N_19439,N_19851);
nand UO_709 (O_709,N_18112,N_18371);
xor UO_710 (O_710,N_19338,N_18553);
or UO_711 (O_711,N_18379,N_19921);
or UO_712 (O_712,N_19841,N_19236);
or UO_713 (O_713,N_18651,N_18724);
nand UO_714 (O_714,N_18400,N_18246);
nand UO_715 (O_715,N_18959,N_18142);
nor UO_716 (O_716,N_19111,N_19434);
xor UO_717 (O_717,N_18225,N_19079);
or UO_718 (O_718,N_19081,N_19990);
nor UO_719 (O_719,N_18262,N_19240);
nor UO_720 (O_720,N_19929,N_18170);
and UO_721 (O_721,N_18860,N_19633);
nand UO_722 (O_722,N_18741,N_18924);
nor UO_723 (O_723,N_19441,N_18052);
and UO_724 (O_724,N_18203,N_18065);
xor UO_725 (O_725,N_19817,N_18305);
xnor UO_726 (O_726,N_19322,N_18993);
xor UO_727 (O_727,N_19278,N_19195);
xnor UO_728 (O_728,N_19583,N_18555);
or UO_729 (O_729,N_18566,N_18219);
nor UO_730 (O_730,N_18858,N_18463);
or UO_731 (O_731,N_18410,N_18232);
or UO_732 (O_732,N_19651,N_19388);
nand UO_733 (O_733,N_19342,N_19427);
nand UO_734 (O_734,N_19151,N_19225);
nand UO_735 (O_735,N_18269,N_19180);
xor UO_736 (O_736,N_19077,N_18123);
nand UO_737 (O_737,N_19246,N_18412);
xor UO_738 (O_738,N_18116,N_18090);
or UO_739 (O_739,N_18702,N_19277);
xnor UO_740 (O_740,N_18157,N_18234);
nand UO_741 (O_741,N_18008,N_18509);
nand UO_742 (O_742,N_18626,N_18095);
nor UO_743 (O_743,N_18339,N_19442);
nor UO_744 (O_744,N_19372,N_19096);
xor UO_745 (O_745,N_18522,N_18560);
xor UO_746 (O_746,N_19088,N_18055);
or UO_747 (O_747,N_19066,N_19381);
nor UO_748 (O_748,N_19341,N_18241);
or UO_749 (O_749,N_18618,N_18587);
or UO_750 (O_750,N_19229,N_18436);
nor UO_751 (O_751,N_19164,N_19406);
nor UO_752 (O_752,N_19655,N_18391);
and UO_753 (O_753,N_18642,N_18632);
or UO_754 (O_754,N_18682,N_18214);
nor UO_755 (O_755,N_18830,N_19864);
and UO_756 (O_756,N_19560,N_18105);
or UO_757 (O_757,N_18661,N_18677);
or UO_758 (O_758,N_18033,N_18064);
nand UO_759 (O_759,N_18472,N_19597);
xnor UO_760 (O_760,N_19935,N_19944);
nor UO_761 (O_761,N_19528,N_18229);
nand UO_762 (O_762,N_18274,N_18252);
xor UO_763 (O_763,N_19302,N_18822);
and UO_764 (O_764,N_18089,N_19539);
xor UO_765 (O_765,N_19745,N_19349);
or UO_766 (O_766,N_19325,N_19867);
xor UO_767 (O_767,N_18453,N_19319);
nand UO_768 (O_768,N_19982,N_18159);
nor UO_769 (O_769,N_19281,N_18310);
xnor UO_770 (O_770,N_18086,N_19688);
xor UO_771 (O_771,N_19196,N_19802);
or UO_772 (O_772,N_18351,N_19333);
xnor UO_773 (O_773,N_18458,N_19706);
nand UO_774 (O_774,N_19593,N_19047);
or UO_775 (O_775,N_18931,N_19360);
or UO_776 (O_776,N_18825,N_19398);
xnor UO_777 (O_777,N_19031,N_19517);
and UO_778 (O_778,N_19906,N_18770);
or UO_779 (O_779,N_19362,N_19752);
and UO_780 (O_780,N_19618,N_19984);
xor UO_781 (O_781,N_19324,N_18511);
and UO_782 (O_782,N_18905,N_19450);
nor UO_783 (O_783,N_18485,N_18668);
xnor UO_784 (O_784,N_18733,N_19363);
or UO_785 (O_785,N_19827,N_19963);
nor UO_786 (O_786,N_19108,N_18070);
xnor UO_787 (O_787,N_18276,N_18853);
nor UO_788 (O_788,N_19401,N_18111);
nand UO_789 (O_789,N_18267,N_18455);
nor UO_790 (O_790,N_19776,N_19141);
or UO_791 (O_791,N_19756,N_18543);
and UO_792 (O_792,N_19206,N_19732);
or UO_793 (O_793,N_18377,N_19810);
nor UO_794 (O_794,N_18927,N_19533);
or UO_795 (O_795,N_19307,N_18334);
or UO_796 (O_796,N_19798,N_18437);
nor UO_797 (O_797,N_18253,N_19028);
and UO_798 (O_798,N_19573,N_19964);
and UO_799 (O_799,N_18374,N_18558);
xor UO_800 (O_800,N_18523,N_19920);
xnor UO_801 (O_801,N_18335,N_18659);
xor UO_802 (O_802,N_18717,N_18868);
nor UO_803 (O_803,N_18268,N_18044);
and UO_804 (O_804,N_19800,N_19407);
xor UO_805 (O_805,N_19865,N_18521);
nor UO_806 (O_806,N_18000,N_18385);
xnor UO_807 (O_807,N_18368,N_19492);
and UO_808 (O_808,N_18740,N_19449);
xnor UO_809 (O_809,N_18735,N_19753);
and UO_810 (O_810,N_19692,N_19062);
or UO_811 (O_811,N_18035,N_18162);
or UO_812 (O_812,N_18766,N_18202);
xor UO_813 (O_813,N_18369,N_19588);
xnor UO_814 (O_814,N_18301,N_19853);
xor UO_815 (O_815,N_18360,N_19552);
or UO_816 (O_816,N_18365,N_19761);
and UO_817 (O_817,N_19171,N_18297);
or UO_818 (O_818,N_18149,N_18275);
xor UO_819 (O_819,N_18386,N_18675);
xnor UO_820 (O_820,N_18729,N_18196);
and UO_821 (O_821,N_18650,N_19764);
xnor UO_822 (O_822,N_18946,N_19385);
or UO_823 (O_823,N_18434,N_19816);
xor UO_824 (O_824,N_19663,N_19832);
nand UO_825 (O_825,N_18600,N_18952);
nor UO_826 (O_826,N_19603,N_18270);
or UO_827 (O_827,N_19710,N_19627);
nand UO_828 (O_828,N_19198,N_19383);
nand UO_829 (O_829,N_19674,N_19359);
and UO_830 (O_830,N_19253,N_19416);
nor UO_831 (O_831,N_18317,N_19979);
xnor UO_832 (O_832,N_19522,N_19134);
xor UO_833 (O_833,N_18549,N_18943);
nand UO_834 (O_834,N_19152,N_19418);
or UO_835 (O_835,N_18106,N_19883);
nor UO_836 (O_836,N_18343,N_19002);
or UO_837 (O_837,N_18781,N_19870);
and UO_838 (O_838,N_19997,N_19951);
nor UO_839 (O_839,N_18956,N_19531);
nand UO_840 (O_840,N_19925,N_19782);
or UO_841 (O_841,N_19489,N_19337);
and UO_842 (O_842,N_19150,N_19387);
or UO_843 (O_843,N_18471,N_18315);
or UO_844 (O_844,N_19351,N_19793);
nor UO_845 (O_845,N_18182,N_18342);
nor UO_846 (O_846,N_18432,N_18711);
xnor UO_847 (O_847,N_18832,N_18851);
nand UO_848 (O_848,N_18983,N_18902);
or UO_849 (O_849,N_18345,N_18108);
xor UO_850 (O_850,N_18564,N_19527);
nor UO_851 (O_851,N_18752,N_18888);
or UO_852 (O_852,N_18971,N_19485);
nor UO_853 (O_853,N_19762,N_19680);
or UO_854 (O_854,N_18970,N_19500);
xnor UO_855 (O_855,N_19672,N_19440);
nor UO_856 (O_856,N_18290,N_18311);
xor UO_857 (O_857,N_18154,N_19403);
nor UO_858 (O_858,N_18978,N_18199);
nand UO_859 (O_859,N_18063,N_19536);
nor UO_860 (O_860,N_18846,N_19393);
and UO_861 (O_861,N_18038,N_18185);
xnor UO_862 (O_862,N_18751,N_19656);
nor UO_863 (O_863,N_19907,N_19551);
and UO_864 (O_864,N_19455,N_19136);
or UO_865 (O_865,N_19394,N_18043);
or UO_866 (O_866,N_18179,N_18392);
nand UO_867 (O_867,N_18547,N_19880);
or UO_868 (O_868,N_19068,N_18582);
xor UO_869 (O_869,N_18953,N_19638);
nor UO_870 (O_870,N_18175,N_18728);
or UO_871 (O_871,N_19999,N_19824);
or UO_872 (O_872,N_18798,N_18881);
xnor UO_873 (O_873,N_18120,N_18876);
xnor UO_874 (O_874,N_19771,N_19090);
nand UO_875 (O_875,N_18688,N_19785);
or UO_876 (O_876,N_19953,N_19609);
xor UO_877 (O_877,N_18601,N_19978);
or UO_878 (O_878,N_18336,N_18459);
and UO_879 (O_879,N_18387,N_19833);
or UO_880 (O_880,N_18308,N_18049);
nor UO_881 (O_881,N_19985,N_18282);
nor UO_882 (O_882,N_19125,N_18667);
nor UO_883 (O_883,N_18570,N_18445);
or UO_884 (O_884,N_19158,N_18769);
xnor UO_885 (O_885,N_19098,N_18945);
nor UO_886 (O_886,N_18398,N_19182);
or UO_887 (O_887,N_18513,N_18389);
or UO_888 (O_888,N_19348,N_18230);
or UO_889 (O_889,N_19084,N_19595);
or UO_890 (O_890,N_18235,N_19862);
and UO_891 (O_891,N_18692,N_19787);
nand UO_892 (O_892,N_19607,N_19709);
nand UO_893 (O_893,N_19636,N_18506);
or UO_894 (O_894,N_19233,N_18278);
and UO_895 (O_895,N_19813,N_19204);
nor UO_896 (O_896,N_18892,N_19801);
or UO_897 (O_897,N_19453,N_18492);
or UO_898 (O_898,N_19511,N_19486);
xnor UO_899 (O_899,N_19975,N_18637);
nor UO_900 (O_900,N_19556,N_18921);
and UO_901 (O_901,N_18965,N_19034);
nor UO_902 (O_902,N_18541,N_19346);
nand UO_903 (O_903,N_18370,N_18127);
or UO_904 (O_904,N_19142,N_18200);
or UO_905 (O_905,N_19117,N_18932);
xnor UO_906 (O_906,N_19433,N_19291);
xor UO_907 (O_907,N_19613,N_19234);
or UO_908 (O_908,N_18188,N_19789);
and UO_909 (O_909,N_18592,N_19836);
and UO_910 (O_910,N_18286,N_18376);
xor UO_911 (O_911,N_18211,N_18240);
or UO_912 (O_912,N_19639,N_18624);
nand UO_913 (O_913,N_19610,N_19058);
nor UO_914 (O_914,N_19538,N_18877);
nor UO_915 (O_915,N_18018,N_19070);
xor UO_916 (O_916,N_19475,N_19011);
nor UO_917 (O_917,N_18372,N_18042);
or UO_918 (O_918,N_19662,N_19114);
or UO_919 (O_919,N_18321,N_18312);
nand UO_920 (O_920,N_19614,N_18013);
nor UO_921 (O_921,N_19804,N_18737);
nand UO_922 (O_922,N_19866,N_18535);
nor UO_923 (O_923,N_18794,N_18588);
nor UO_924 (O_924,N_19731,N_19217);
nor UO_925 (O_925,N_18663,N_18911);
nor UO_926 (O_926,N_18736,N_18536);
xnor UO_927 (O_927,N_19255,N_18646);
or UO_928 (O_928,N_18026,N_18088);
xor UO_929 (O_929,N_19949,N_19767);
or UO_930 (O_930,N_19411,N_19464);
nor UO_931 (O_931,N_19730,N_18264);
and UO_932 (O_932,N_18081,N_19495);
nor UO_933 (O_933,N_18059,N_18643);
or UO_934 (O_934,N_19818,N_19001);
nand UO_935 (O_935,N_18738,N_19967);
or UO_936 (O_936,N_18104,N_19318);
nor UO_937 (O_937,N_18638,N_19715);
nor UO_938 (O_938,N_18140,N_18266);
and UO_939 (O_939,N_18337,N_18548);
xnor UO_940 (O_940,N_19273,N_18837);
xor UO_941 (O_941,N_18474,N_18121);
and UO_942 (O_942,N_19667,N_19078);
nor UO_943 (O_943,N_18395,N_19594);
nor UO_944 (O_944,N_19670,N_19445);
nand UO_945 (O_945,N_18145,N_19520);
nand UO_946 (O_946,N_19987,N_19809);
xor UO_947 (O_947,N_18294,N_18011);
and UO_948 (O_948,N_18071,N_18620);
xnor UO_949 (O_949,N_19746,N_19192);
or UO_950 (O_950,N_19910,N_18915);
nand UO_951 (O_951,N_18712,N_18438);
nor UO_952 (O_952,N_19241,N_19786);
xnor UO_953 (O_953,N_18730,N_19239);
and UO_954 (O_954,N_19375,N_19724);
nand UO_955 (O_955,N_19041,N_18685);
xnor UO_956 (O_956,N_18893,N_18974);
nand UO_957 (O_957,N_19496,N_19623);
xor UO_958 (O_958,N_19828,N_18991);
nor UO_959 (O_959,N_19902,N_19876);
nand UO_960 (O_960,N_19215,N_19404);
nand UO_961 (O_961,N_18201,N_19044);
and UO_962 (O_962,N_19868,N_19948);
nand UO_963 (O_963,N_19269,N_19467);
nand UO_964 (O_964,N_19400,N_18771);
nand UO_965 (O_965,N_18627,N_19316);
and UO_966 (O_966,N_18516,N_18532);
xnor UO_967 (O_967,N_19122,N_18094);
nor UO_968 (O_968,N_19373,N_18041);
xnor UO_969 (O_969,N_18402,N_19135);
or UO_970 (O_970,N_19696,N_18569);
nor UO_971 (O_971,N_18354,N_18575);
and UO_972 (O_972,N_19976,N_18510);
and UO_973 (O_973,N_18491,N_19199);
and UO_974 (O_974,N_18028,N_18192);
xor UO_975 (O_975,N_18388,N_18168);
xor UO_976 (O_976,N_19057,N_18852);
and UO_977 (O_977,N_19510,N_18223);
nand UO_978 (O_978,N_19878,N_19888);
nor UO_979 (O_979,N_19452,N_19376);
or UO_980 (O_980,N_18022,N_19396);
nand UO_981 (O_981,N_19208,N_18079);
nand UO_982 (O_982,N_19432,N_19586);
and UO_983 (O_983,N_19310,N_19218);
nor UO_984 (O_984,N_19557,N_18960);
nor UO_985 (O_985,N_18958,N_18279);
xnor UO_986 (O_986,N_19227,N_19899);
nor UO_987 (O_987,N_19701,N_18213);
nor UO_988 (O_988,N_18486,N_18849);
nand UO_989 (O_989,N_19580,N_19428);
xor UO_990 (O_990,N_18481,N_18936);
and UO_991 (O_991,N_19268,N_18686);
or UO_992 (O_992,N_18901,N_19887);
nor UO_993 (O_993,N_18599,N_19190);
or UO_994 (O_994,N_19390,N_18961);
xnor UO_995 (O_995,N_19721,N_18164);
xor UO_996 (O_996,N_18734,N_18833);
nand UO_997 (O_997,N_19405,N_19846);
nor UO_998 (O_998,N_19735,N_19421);
xnor UO_999 (O_999,N_18151,N_19183);
or UO_1000 (O_1000,N_19088,N_19273);
nor UO_1001 (O_1001,N_19774,N_19459);
or UO_1002 (O_1002,N_18826,N_18572);
nor UO_1003 (O_1003,N_18637,N_19905);
nor UO_1004 (O_1004,N_18922,N_18565);
xnor UO_1005 (O_1005,N_19679,N_18204);
nor UO_1006 (O_1006,N_19400,N_18121);
xor UO_1007 (O_1007,N_18721,N_19312);
nor UO_1008 (O_1008,N_19679,N_18607);
and UO_1009 (O_1009,N_19557,N_18703);
or UO_1010 (O_1010,N_19493,N_18425);
and UO_1011 (O_1011,N_19416,N_19242);
nor UO_1012 (O_1012,N_19916,N_19569);
xnor UO_1013 (O_1013,N_18187,N_19875);
nand UO_1014 (O_1014,N_18119,N_19811);
nor UO_1015 (O_1015,N_19575,N_19757);
nand UO_1016 (O_1016,N_19679,N_19399);
xnor UO_1017 (O_1017,N_19191,N_19629);
nand UO_1018 (O_1018,N_18090,N_19555);
or UO_1019 (O_1019,N_18202,N_19069);
and UO_1020 (O_1020,N_18436,N_18893);
and UO_1021 (O_1021,N_19101,N_19378);
nand UO_1022 (O_1022,N_19182,N_18562);
nand UO_1023 (O_1023,N_19471,N_19485);
xnor UO_1024 (O_1024,N_19488,N_19179);
and UO_1025 (O_1025,N_19222,N_19953);
nand UO_1026 (O_1026,N_19046,N_19485);
xnor UO_1027 (O_1027,N_18200,N_18025);
and UO_1028 (O_1028,N_18773,N_19234);
or UO_1029 (O_1029,N_19205,N_19622);
xnor UO_1030 (O_1030,N_18977,N_18557);
or UO_1031 (O_1031,N_18528,N_19497);
xnor UO_1032 (O_1032,N_18799,N_19417);
or UO_1033 (O_1033,N_18409,N_19394);
nor UO_1034 (O_1034,N_18756,N_19460);
and UO_1035 (O_1035,N_18927,N_18437);
or UO_1036 (O_1036,N_19141,N_18859);
nand UO_1037 (O_1037,N_18185,N_19854);
xor UO_1038 (O_1038,N_19077,N_19614);
and UO_1039 (O_1039,N_18403,N_18031);
or UO_1040 (O_1040,N_19406,N_19574);
and UO_1041 (O_1041,N_19889,N_18403);
or UO_1042 (O_1042,N_19312,N_19607);
and UO_1043 (O_1043,N_18296,N_19601);
nor UO_1044 (O_1044,N_18371,N_19617);
or UO_1045 (O_1045,N_19893,N_18527);
nor UO_1046 (O_1046,N_18336,N_18155);
nor UO_1047 (O_1047,N_19724,N_18044);
nor UO_1048 (O_1048,N_18826,N_19061);
nor UO_1049 (O_1049,N_18350,N_19794);
nand UO_1050 (O_1050,N_19210,N_19175);
xor UO_1051 (O_1051,N_18273,N_18092);
nand UO_1052 (O_1052,N_18463,N_19804);
or UO_1053 (O_1053,N_18360,N_18311);
nand UO_1054 (O_1054,N_19807,N_19672);
or UO_1055 (O_1055,N_18007,N_19645);
nand UO_1056 (O_1056,N_18486,N_19178);
nor UO_1057 (O_1057,N_19293,N_19700);
nor UO_1058 (O_1058,N_19471,N_19119);
xnor UO_1059 (O_1059,N_18307,N_18736);
and UO_1060 (O_1060,N_18182,N_19130);
nand UO_1061 (O_1061,N_19792,N_18688);
nand UO_1062 (O_1062,N_18032,N_19364);
nor UO_1063 (O_1063,N_18939,N_19072);
nor UO_1064 (O_1064,N_18567,N_19843);
nor UO_1065 (O_1065,N_19170,N_19129);
or UO_1066 (O_1066,N_19184,N_18166);
nand UO_1067 (O_1067,N_18551,N_19867);
nor UO_1068 (O_1068,N_19332,N_18381);
and UO_1069 (O_1069,N_19662,N_19478);
and UO_1070 (O_1070,N_18165,N_19206);
and UO_1071 (O_1071,N_18431,N_18527);
nand UO_1072 (O_1072,N_18541,N_18985);
xor UO_1073 (O_1073,N_19174,N_18631);
xnor UO_1074 (O_1074,N_18436,N_19327);
or UO_1075 (O_1075,N_19461,N_19222);
xor UO_1076 (O_1076,N_18825,N_18816);
and UO_1077 (O_1077,N_18203,N_18838);
and UO_1078 (O_1078,N_18924,N_18560);
nor UO_1079 (O_1079,N_19806,N_18465);
and UO_1080 (O_1080,N_19806,N_19963);
xor UO_1081 (O_1081,N_18590,N_19038);
and UO_1082 (O_1082,N_19400,N_18862);
nand UO_1083 (O_1083,N_19215,N_19750);
or UO_1084 (O_1084,N_18799,N_19122);
or UO_1085 (O_1085,N_19511,N_19458);
and UO_1086 (O_1086,N_19140,N_19249);
xor UO_1087 (O_1087,N_19712,N_19407);
nand UO_1088 (O_1088,N_18582,N_18921);
or UO_1089 (O_1089,N_18251,N_18761);
and UO_1090 (O_1090,N_19028,N_19180);
nor UO_1091 (O_1091,N_19015,N_18624);
xor UO_1092 (O_1092,N_18334,N_19806);
and UO_1093 (O_1093,N_18769,N_18701);
nor UO_1094 (O_1094,N_19536,N_18610);
and UO_1095 (O_1095,N_19281,N_19335);
and UO_1096 (O_1096,N_18779,N_18842);
and UO_1097 (O_1097,N_18524,N_19368);
or UO_1098 (O_1098,N_18950,N_18587);
or UO_1099 (O_1099,N_19253,N_19122);
and UO_1100 (O_1100,N_18642,N_18448);
nand UO_1101 (O_1101,N_19464,N_18214);
xor UO_1102 (O_1102,N_19767,N_18158);
nor UO_1103 (O_1103,N_18948,N_19970);
nor UO_1104 (O_1104,N_19723,N_19705);
nand UO_1105 (O_1105,N_18297,N_18091);
nand UO_1106 (O_1106,N_18907,N_18651);
nand UO_1107 (O_1107,N_19471,N_19758);
xor UO_1108 (O_1108,N_18324,N_18778);
and UO_1109 (O_1109,N_18551,N_19148);
xor UO_1110 (O_1110,N_18816,N_19705);
or UO_1111 (O_1111,N_18698,N_18348);
xnor UO_1112 (O_1112,N_18514,N_19020);
xor UO_1113 (O_1113,N_19856,N_18089);
xnor UO_1114 (O_1114,N_18826,N_19276);
or UO_1115 (O_1115,N_18720,N_18043);
nand UO_1116 (O_1116,N_19003,N_18113);
xor UO_1117 (O_1117,N_19189,N_18455);
nand UO_1118 (O_1118,N_19312,N_19122);
nand UO_1119 (O_1119,N_18454,N_18509);
and UO_1120 (O_1120,N_18161,N_19016);
or UO_1121 (O_1121,N_19450,N_19014);
nand UO_1122 (O_1122,N_19108,N_18089);
and UO_1123 (O_1123,N_18768,N_18781);
or UO_1124 (O_1124,N_19679,N_19478);
nand UO_1125 (O_1125,N_18127,N_18083);
or UO_1126 (O_1126,N_18577,N_19487);
nor UO_1127 (O_1127,N_18754,N_18453);
and UO_1128 (O_1128,N_18704,N_19537);
or UO_1129 (O_1129,N_18283,N_18343);
xnor UO_1130 (O_1130,N_18999,N_19612);
xor UO_1131 (O_1131,N_18525,N_19440);
and UO_1132 (O_1132,N_19723,N_19455);
nor UO_1133 (O_1133,N_18735,N_18517);
xor UO_1134 (O_1134,N_18361,N_19083);
nor UO_1135 (O_1135,N_19338,N_18417);
nand UO_1136 (O_1136,N_19009,N_19884);
nand UO_1137 (O_1137,N_19488,N_18542);
nor UO_1138 (O_1138,N_18853,N_18232);
xor UO_1139 (O_1139,N_19321,N_19873);
nor UO_1140 (O_1140,N_18524,N_18837);
and UO_1141 (O_1141,N_18277,N_19864);
or UO_1142 (O_1142,N_19494,N_19988);
xor UO_1143 (O_1143,N_19196,N_18666);
and UO_1144 (O_1144,N_19893,N_18323);
nor UO_1145 (O_1145,N_19929,N_18334);
nand UO_1146 (O_1146,N_19653,N_19205);
nor UO_1147 (O_1147,N_19693,N_18466);
xnor UO_1148 (O_1148,N_19975,N_19527);
nor UO_1149 (O_1149,N_19981,N_19210);
nor UO_1150 (O_1150,N_18458,N_18796);
and UO_1151 (O_1151,N_18705,N_18960);
nand UO_1152 (O_1152,N_18483,N_19996);
xor UO_1153 (O_1153,N_19845,N_19111);
nor UO_1154 (O_1154,N_18011,N_18663);
and UO_1155 (O_1155,N_18392,N_18102);
nand UO_1156 (O_1156,N_18754,N_19242);
xnor UO_1157 (O_1157,N_19150,N_18098);
and UO_1158 (O_1158,N_19385,N_19333);
and UO_1159 (O_1159,N_19693,N_19066);
xor UO_1160 (O_1160,N_19667,N_19957);
nor UO_1161 (O_1161,N_19066,N_18937);
xnor UO_1162 (O_1162,N_18590,N_19042);
nor UO_1163 (O_1163,N_19462,N_18544);
and UO_1164 (O_1164,N_19220,N_19813);
or UO_1165 (O_1165,N_19459,N_19717);
and UO_1166 (O_1166,N_19035,N_18177);
or UO_1167 (O_1167,N_18593,N_18684);
xor UO_1168 (O_1168,N_19182,N_18524);
nor UO_1169 (O_1169,N_18583,N_19759);
or UO_1170 (O_1170,N_18716,N_19515);
and UO_1171 (O_1171,N_18937,N_19437);
and UO_1172 (O_1172,N_18165,N_18510);
xnor UO_1173 (O_1173,N_19171,N_19449);
and UO_1174 (O_1174,N_18862,N_18375);
and UO_1175 (O_1175,N_18917,N_18338);
xnor UO_1176 (O_1176,N_19230,N_19814);
xor UO_1177 (O_1177,N_18291,N_19984);
and UO_1178 (O_1178,N_18166,N_18966);
and UO_1179 (O_1179,N_18550,N_18918);
and UO_1180 (O_1180,N_19160,N_19182);
or UO_1181 (O_1181,N_18958,N_18731);
nor UO_1182 (O_1182,N_19563,N_18424);
nor UO_1183 (O_1183,N_18550,N_18514);
xnor UO_1184 (O_1184,N_19262,N_19944);
or UO_1185 (O_1185,N_19275,N_19451);
xor UO_1186 (O_1186,N_18691,N_18881);
or UO_1187 (O_1187,N_19567,N_19125);
xnor UO_1188 (O_1188,N_18773,N_18553);
nor UO_1189 (O_1189,N_18443,N_19093);
or UO_1190 (O_1190,N_19723,N_18395);
nand UO_1191 (O_1191,N_19334,N_19741);
nand UO_1192 (O_1192,N_19010,N_19479);
nor UO_1193 (O_1193,N_18344,N_18782);
or UO_1194 (O_1194,N_18174,N_18451);
xnor UO_1195 (O_1195,N_18442,N_19956);
nor UO_1196 (O_1196,N_18691,N_19440);
xor UO_1197 (O_1197,N_18266,N_19515);
nor UO_1198 (O_1198,N_19461,N_18647);
or UO_1199 (O_1199,N_19086,N_19133);
and UO_1200 (O_1200,N_18180,N_18839);
nand UO_1201 (O_1201,N_19669,N_19504);
or UO_1202 (O_1202,N_19107,N_19386);
or UO_1203 (O_1203,N_19809,N_18944);
nor UO_1204 (O_1204,N_18911,N_18422);
or UO_1205 (O_1205,N_18922,N_18096);
nand UO_1206 (O_1206,N_18856,N_18366);
or UO_1207 (O_1207,N_18764,N_18230);
xnor UO_1208 (O_1208,N_19293,N_18111);
nor UO_1209 (O_1209,N_18410,N_19480);
nor UO_1210 (O_1210,N_18927,N_19078);
and UO_1211 (O_1211,N_18431,N_18068);
nand UO_1212 (O_1212,N_19225,N_19242);
and UO_1213 (O_1213,N_19219,N_18511);
nor UO_1214 (O_1214,N_18778,N_19956);
nand UO_1215 (O_1215,N_19898,N_19910);
xor UO_1216 (O_1216,N_19833,N_19636);
nor UO_1217 (O_1217,N_18431,N_18353);
and UO_1218 (O_1218,N_18535,N_19529);
nor UO_1219 (O_1219,N_18168,N_19321);
nor UO_1220 (O_1220,N_19430,N_19650);
nand UO_1221 (O_1221,N_18706,N_19564);
nor UO_1222 (O_1222,N_19677,N_18430);
nor UO_1223 (O_1223,N_19560,N_18964);
xnor UO_1224 (O_1224,N_18746,N_19389);
nor UO_1225 (O_1225,N_19843,N_19575);
nand UO_1226 (O_1226,N_19794,N_18984);
or UO_1227 (O_1227,N_19593,N_19286);
nor UO_1228 (O_1228,N_18971,N_18859);
nor UO_1229 (O_1229,N_18409,N_18683);
xnor UO_1230 (O_1230,N_19471,N_19554);
and UO_1231 (O_1231,N_18621,N_19875);
nor UO_1232 (O_1232,N_18895,N_19026);
nand UO_1233 (O_1233,N_18073,N_18067);
xnor UO_1234 (O_1234,N_18718,N_19444);
xor UO_1235 (O_1235,N_18894,N_18825);
nor UO_1236 (O_1236,N_19950,N_18030);
nor UO_1237 (O_1237,N_18357,N_18015);
and UO_1238 (O_1238,N_19535,N_18788);
nand UO_1239 (O_1239,N_18012,N_19597);
xnor UO_1240 (O_1240,N_19225,N_19132);
or UO_1241 (O_1241,N_19955,N_18712);
xor UO_1242 (O_1242,N_19095,N_19858);
or UO_1243 (O_1243,N_18516,N_19552);
nand UO_1244 (O_1244,N_18526,N_19880);
nor UO_1245 (O_1245,N_19267,N_19358);
nor UO_1246 (O_1246,N_19432,N_18151);
or UO_1247 (O_1247,N_18578,N_19438);
and UO_1248 (O_1248,N_18867,N_18203);
nor UO_1249 (O_1249,N_18333,N_19229);
nor UO_1250 (O_1250,N_19962,N_18481);
nor UO_1251 (O_1251,N_19858,N_19984);
or UO_1252 (O_1252,N_19229,N_19581);
and UO_1253 (O_1253,N_19415,N_18151);
and UO_1254 (O_1254,N_19971,N_19765);
xor UO_1255 (O_1255,N_18722,N_18739);
nand UO_1256 (O_1256,N_19301,N_18688);
or UO_1257 (O_1257,N_19988,N_19038);
or UO_1258 (O_1258,N_18195,N_19462);
xnor UO_1259 (O_1259,N_19220,N_18515);
and UO_1260 (O_1260,N_18702,N_19566);
nor UO_1261 (O_1261,N_19403,N_18693);
nor UO_1262 (O_1262,N_19561,N_19588);
or UO_1263 (O_1263,N_18550,N_18985);
or UO_1264 (O_1264,N_19588,N_18623);
nand UO_1265 (O_1265,N_19987,N_18479);
xor UO_1266 (O_1266,N_19534,N_19420);
and UO_1267 (O_1267,N_19909,N_19403);
and UO_1268 (O_1268,N_18468,N_18338);
nand UO_1269 (O_1269,N_19051,N_18603);
and UO_1270 (O_1270,N_19856,N_18543);
or UO_1271 (O_1271,N_18546,N_18659);
or UO_1272 (O_1272,N_19477,N_18727);
nand UO_1273 (O_1273,N_19779,N_18105);
and UO_1274 (O_1274,N_19644,N_19540);
xnor UO_1275 (O_1275,N_18174,N_18419);
nand UO_1276 (O_1276,N_19083,N_18437);
and UO_1277 (O_1277,N_18513,N_18198);
and UO_1278 (O_1278,N_18854,N_18790);
nor UO_1279 (O_1279,N_18953,N_19444);
or UO_1280 (O_1280,N_18594,N_18731);
xor UO_1281 (O_1281,N_18658,N_18722);
nor UO_1282 (O_1282,N_18546,N_18196);
xor UO_1283 (O_1283,N_18632,N_18343);
nor UO_1284 (O_1284,N_19855,N_18028);
nand UO_1285 (O_1285,N_18782,N_18062);
nand UO_1286 (O_1286,N_18814,N_19423);
and UO_1287 (O_1287,N_18882,N_18249);
xnor UO_1288 (O_1288,N_19078,N_18207);
nor UO_1289 (O_1289,N_18949,N_19060);
or UO_1290 (O_1290,N_18560,N_19512);
nor UO_1291 (O_1291,N_19685,N_18431);
xor UO_1292 (O_1292,N_19509,N_19646);
and UO_1293 (O_1293,N_18944,N_19344);
nor UO_1294 (O_1294,N_18808,N_18038);
and UO_1295 (O_1295,N_19718,N_18858);
nor UO_1296 (O_1296,N_19512,N_19664);
xor UO_1297 (O_1297,N_19365,N_19018);
xnor UO_1298 (O_1298,N_19004,N_18830);
nand UO_1299 (O_1299,N_18283,N_19556);
nand UO_1300 (O_1300,N_19084,N_18832);
or UO_1301 (O_1301,N_19754,N_19072);
nand UO_1302 (O_1302,N_18251,N_18294);
nor UO_1303 (O_1303,N_18589,N_19659);
nand UO_1304 (O_1304,N_18416,N_19764);
xnor UO_1305 (O_1305,N_19307,N_19538);
xnor UO_1306 (O_1306,N_18400,N_18336);
nand UO_1307 (O_1307,N_19113,N_19882);
nor UO_1308 (O_1308,N_18980,N_19612);
xor UO_1309 (O_1309,N_19668,N_19967);
or UO_1310 (O_1310,N_19741,N_18471);
or UO_1311 (O_1311,N_18566,N_19841);
or UO_1312 (O_1312,N_19171,N_19064);
nand UO_1313 (O_1313,N_18295,N_18612);
and UO_1314 (O_1314,N_19084,N_19826);
nand UO_1315 (O_1315,N_18230,N_19192);
and UO_1316 (O_1316,N_19753,N_18908);
nor UO_1317 (O_1317,N_19174,N_19119);
xnor UO_1318 (O_1318,N_18647,N_19889);
nand UO_1319 (O_1319,N_19198,N_19360);
or UO_1320 (O_1320,N_18809,N_19264);
and UO_1321 (O_1321,N_18408,N_19585);
nor UO_1322 (O_1322,N_19194,N_18525);
xor UO_1323 (O_1323,N_18166,N_19811);
or UO_1324 (O_1324,N_19384,N_19099);
xnor UO_1325 (O_1325,N_18109,N_18499);
xor UO_1326 (O_1326,N_19408,N_18706);
and UO_1327 (O_1327,N_18909,N_18356);
and UO_1328 (O_1328,N_18027,N_19963);
nor UO_1329 (O_1329,N_18948,N_19446);
and UO_1330 (O_1330,N_18683,N_19930);
nand UO_1331 (O_1331,N_18300,N_19695);
nor UO_1332 (O_1332,N_19966,N_19285);
or UO_1333 (O_1333,N_18709,N_18763);
or UO_1334 (O_1334,N_19094,N_19730);
nand UO_1335 (O_1335,N_18129,N_18146);
or UO_1336 (O_1336,N_18653,N_19157);
xnor UO_1337 (O_1337,N_19828,N_19363);
or UO_1338 (O_1338,N_18001,N_19469);
xor UO_1339 (O_1339,N_19060,N_19842);
or UO_1340 (O_1340,N_18940,N_18563);
nor UO_1341 (O_1341,N_18054,N_18248);
or UO_1342 (O_1342,N_19766,N_18820);
nand UO_1343 (O_1343,N_18936,N_18880);
or UO_1344 (O_1344,N_19211,N_19796);
nor UO_1345 (O_1345,N_18412,N_19051);
nand UO_1346 (O_1346,N_19935,N_19783);
and UO_1347 (O_1347,N_18833,N_19015);
xor UO_1348 (O_1348,N_18373,N_18778);
nor UO_1349 (O_1349,N_19114,N_19497);
xnor UO_1350 (O_1350,N_18940,N_18566);
nand UO_1351 (O_1351,N_19927,N_19309);
nor UO_1352 (O_1352,N_18951,N_18115);
nor UO_1353 (O_1353,N_18449,N_19391);
or UO_1354 (O_1354,N_18885,N_19961);
nand UO_1355 (O_1355,N_18477,N_19072);
and UO_1356 (O_1356,N_18715,N_18532);
nand UO_1357 (O_1357,N_18109,N_18072);
or UO_1358 (O_1358,N_18882,N_19203);
and UO_1359 (O_1359,N_18783,N_19736);
nand UO_1360 (O_1360,N_19176,N_19270);
and UO_1361 (O_1361,N_19205,N_19094);
or UO_1362 (O_1362,N_18318,N_19276);
xor UO_1363 (O_1363,N_18959,N_19001);
or UO_1364 (O_1364,N_19302,N_18645);
and UO_1365 (O_1365,N_18870,N_19093);
nand UO_1366 (O_1366,N_18308,N_18297);
or UO_1367 (O_1367,N_18149,N_18197);
xnor UO_1368 (O_1368,N_18212,N_18418);
and UO_1369 (O_1369,N_18930,N_19787);
or UO_1370 (O_1370,N_19157,N_18883);
and UO_1371 (O_1371,N_18203,N_19524);
nand UO_1372 (O_1372,N_18904,N_19657);
nand UO_1373 (O_1373,N_18572,N_19802);
nand UO_1374 (O_1374,N_19481,N_19658);
nor UO_1375 (O_1375,N_18928,N_19276);
nor UO_1376 (O_1376,N_19405,N_18805);
nand UO_1377 (O_1377,N_19489,N_18728);
nand UO_1378 (O_1378,N_18914,N_18390);
or UO_1379 (O_1379,N_19313,N_19340);
xor UO_1380 (O_1380,N_18909,N_19664);
xnor UO_1381 (O_1381,N_18670,N_18503);
xnor UO_1382 (O_1382,N_18819,N_19453);
and UO_1383 (O_1383,N_18561,N_18517);
and UO_1384 (O_1384,N_19310,N_19587);
and UO_1385 (O_1385,N_19188,N_19087);
xnor UO_1386 (O_1386,N_18252,N_19126);
nor UO_1387 (O_1387,N_19476,N_18092);
nand UO_1388 (O_1388,N_19495,N_18672);
xor UO_1389 (O_1389,N_18781,N_19679);
xnor UO_1390 (O_1390,N_19634,N_18227);
and UO_1391 (O_1391,N_19695,N_18531);
or UO_1392 (O_1392,N_19154,N_19337);
xor UO_1393 (O_1393,N_19839,N_18261);
xor UO_1394 (O_1394,N_18757,N_19625);
or UO_1395 (O_1395,N_18765,N_18060);
nand UO_1396 (O_1396,N_18766,N_18272);
and UO_1397 (O_1397,N_18372,N_18032);
nand UO_1398 (O_1398,N_18520,N_18391);
and UO_1399 (O_1399,N_18623,N_18555);
or UO_1400 (O_1400,N_18949,N_18256);
or UO_1401 (O_1401,N_19461,N_18532);
nand UO_1402 (O_1402,N_19085,N_18575);
xor UO_1403 (O_1403,N_19097,N_19246);
nand UO_1404 (O_1404,N_18020,N_18869);
or UO_1405 (O_1405,N_18363,N_18943);
nor UO_1406 (O_1406,N_19998,N_18709);
nand UO_1407 (O_1407,N_19584,N_19822);
nand UO_1408 (O_1408,N_19783,N_19726);
or UO_1409 (O_1409,N_19253,N_19455);
nor UO_1410 (O_1410,N_18280,N_18893);
and UO_1411 (O_1411,N_19244,N_19155);
nand UO_1412 (O_1412,N_19082,N_18443);
nor UO_1413 (O_1413,N_18338,N_18122);
nand UO_1414 (O_1414,N_19005,N_18370);
and UO_1415 (O_1415,N_19658,N_19283);
xor UO_1416 (O_1416,N_18807,N_19455);
xnor UO_1417 (O_1417,N_19254,N_18605);
or UO_1418 (O_1418,N_18204,N_18289);
nor UO_1419 (O_1419,N_18831,N_18016);
and UO_1420 (O_1420,N_19354,N_19805);
or UO_1421 (O_1421,N_18177,N_19690);
xor UO_1422 (O_1422,N_18338,N_18983);
and UO_1423 (O_1423,N_19916,N_19876);
and UO_1424 (O_1424,N_19002,N_19585);
or UO_1425 (O_1425,N_18747,N_19026);
nand UO_1426 (O_1426,N_19975,N_18154);
nor UO_1427 (O_1427,N_19896,N_18298);
or UO_1428 (O_1428,N_18732,N_19408);
nor UO_1429 (O_1429,N_18723,N_19152);
xor UO_1430 (O_1430,N_19308,N_18738);
or UO_1431 (O_1431,N_19667,N_19676);
nor UO_1432 (O_1432,N_19517,N_18496);
or UO_1433 (O_1433,N_18125,N_19603);
xor UO_1434 (O_1434,N_18825,N_18567);
and UO_1435 (O_1435,N_18352,N_19271);
or UO_1436 (O_1436,N_18891,N_19783);
or UO_1437 (O_1437,N_18367,N_19163);
xnor UO_1438 (O_1438,N_19245,N_19130);
nand UO_1439 (O_1439,N_18544,N_19351);
nor UO_1440 (O_1440,N_18764,N_18794);
nor UO_1441 (O_1441,N_19405,N_19184);
xor UO_1442 (O_1442,N_19625,N_18124);
xnor UO_1443 (O_1443,N_19962,N_19780);
nand UO_1444 (O_1444,N_18730,N_19693);
nand UO_1445 (O_1445,N_18408,N_18748);
nor UO_1446 (O_1446,N_19121,N_19057);
and UO_1447 (O_1447,N_18072,N_19088);
xnor UO_1448 (O_1448,N_19582,N_18114);
or UO_1449 (O_1449,N_19356,N_19629);
nor UO_1450 (O_1450,N_18639,N_18977);
nor UO_1451 (O_1451,N_18709,N_18654);
and UO_1452 (O_1452,N_19710,N_19771);
nand UO_1453 (O_1453,N_18363,N_18102);
nor UO_1454 (O_1454,N_18928,N_19344);
nand UO_1455 (O_1455,N_18177,N_19618);
or UO_1456 (O_1456,N_18762,N_19140);
nor UO_1457 (O_1457,N_19836,N_18504);
nand UO_1458 (O_1458,N_18134,N_18257);
nor UO_1459 (O_1459,N_19669,N_18092);
nor UO_1460 (O_1460,N_18460,N_18188);
xnor UO_1461 (O_1461,N_19654,N_18076);
or UO_1462 (O_1462,N_18537,N_18639);
or UO_1463 (O_1463,N_18970,N_18001);
xnor UO_1464 (O_1464,N_19592,N_18197);
xnor UO_1465 (O_1465,N_18560,N_18188);
nor UO_1466 (O_1466,N_19205,N_19658);
nor UO_1467 (O_1467,N_18829,N_19212);
and UO_1468 (O_1468,N_19009,N_18424);
nor UO_1469 (O_1469,N_18574,N_18789);
xnor UO_1470 (O_1470,N_19502,N_19255);
nor UO_1471 (O_1471,N_18530,N_18878);
or UO_1472 (O_1472,N_18479,N_19373);
and UO_1473 (O_1473,N_18247,N_19076);
xor UO_1474 (O_1474,N_18709,N_18575);
nand UO_1475 (O_1475,N_19778,N_19408);
and UO_1476 (O_1476,N_19621,N_19561);
nand UO_1477 (O_1477,N_19125,N_19032);
or UO_1478 (O_1478,N_18306,N_19419);
or UO_1479 (O_1479,N_18736,N_19367);
nand UO_1480 (O_1480,N_18004,N_18318);
nor UO_1481 (O_1481,N_19745,N_19585);
nand UO_1482 (O_1482,N_19578,N_18560);
xnor UO_1483 (O_1483,N_19399,N_18958);
xor UO_1484 (O_1484,N_18526,N_19814);
or UO_1485 (O_1485,N_18025,N_19935);
nor UO_1486 (O_1486,N_18072,N_19801);
or UO_1487 (O_1487,N_18543,N_19491);
nor UO_1488 (O_1488,N_19135,N_19677);
or UO_1489 (O_1489,N_19912,N_19282);
or UO_1490 (O_1490,N_18436,N_19663);
and UO_1491 (O_1491,N_19686,N_18496);
and UO_1492 (O_1492,N_18143,N_18081);
or UO_1493 (O_1493,N_18025,N_18627);
nor UO_1494 (O_1494,N_19313,N_19491);
nand UO_1495 (O_1495,N_19769,N_19079);
nand UO_1496 (O_1496,N_18315,N_18263);
nand UO_1497 (O_1497,N_18584,N_18413);
nand UO_1498 (O_1498,N_18780,N_18781);
nand UO_1499 (O_1499,N_18476,N_19171);
nor UO_1500 (O_1500,N_18966,N_18825);
xnor UO_1501 (O_1501,N_19478,N_18707);
or UO_1502 (O_1502,N_18278,N_19708);
or UO_1503 (O_1503,N_19808,N_18241);
nor UO_1504 (O_1504,N_18255,N_18093);
and UO_1505 (O_1505,N_18993,N_18388);
or UO_1506 (O_1506,N_18494,N_19450);
and UO_1507 (O_1507,N_18244,N_19992);
xnor UO_1508 (O_1508,N_18145,N_19191);
or UO_1509 (O_1509,N_19786,N_19873);
nand UO_1510 (O_1510,N_18560,N_18218);
and UO_1511 (O_1511,N_18571,N_18779);
or UO_1512 (O_1512,N_19603,N_18470);
xnor UO_1513 (O_1513,N_19594,N_19145);
and UO_1514 (O_1514,N_18510,N_19624);
xor UO_1515 (O_1515,N_18177,N_19084);
nor UO_1516 (O_1516,N_18816,N_19944);
nand UO_1517 (O_1517,N_18066,N_18749);
or UO_1518 (O_1518,N_18144,N_18579);
xor UO_1519 (O_1519,N_18416,N_19750);
or UO_1520 (O_1520,N_18812,N_19511);
nor UO_1521 (O_1521,N_18692,N_18482);
or UO_1522 (O_1522,N_18392,N_18036);
and UO_1523 (O_1523,N_18066,N_19156);
or UO_1524 (O_1524,N_19402,N_19617);
and UO_1525 (O_1525,N_18147,N_19553);
nor UO_1526 (O_1526,N_18116,N_19686);
and UO_1527 (O_1527,N_18859,N_18447);
or UO_1528 (O_1528,N_18326,N_18707);
xor UO_1529 (O_1529,N_19723,N_19606);
xnor UO_1530 (O_1530,N_18580,N_19973);
nor UO_1531 (O_1531,N_18050,N_18899);
and UO_1532 (O_1532,N_18765,N_19800);
or UO_1533 (O_1533,N_19651,N_19051);
and UO_1534 (O_1534,N_18648,N_19580);
nor UO_1535 (O_1535,N_19415,N_19792);
nand UO_1536 (O_1536,N_18020,N_19030);
xnor UO_1537 (O_1537,N_18610,N_19306);
nor UO_1538 (O_1538,N_18820,N_19140);
nor UO_1539 (O_1539,N_19537,N_19988);
nand UO_1540 (O_1540,N_18888,N_19653);
nor UO_1541 (O_1541,N_19072,N_18586);
and UO_1542 (O_1542,N_19236,N_18976);
xnor UO_1543 (O_1543,N_18447,N_19239);
nand UO_1544 (O_1544,N_19647,N_19604);
or UO_1545 (O_1545,N_19056,N_19876);
nand UO_1546 (O_1546,N_19157,N_18432);
xor UO_1547 (O_1547,N_18061,N_19215);
nor UO_1548 (O_1548,N_19184,N_18281);
xnor UO_1549 (O_1549,N_18451,N_18749);
nor UO_1550 (O_1550,N_18594,N_19780);
and UO_1551 (O_1551,N_19499,N_18778);
or UO_1552 (O_1552,N_18032,N_18253);
and UO_1553 (O_1553,N_19656,N_18975);
xor UO_1554 (O_1554,N_19519,N_19438);
or UO_1555 (O_1555,N_19480,N_19492);
xor UO_1556 (O_1556,N_19720,N_18533);
xnor UO_1557 (O_1557,N_19546,N_19357);
nor UO_1558 (O_1558,N_18003,N_18984);
nor UO_1559 (O_1559,N_19121,N_19427);
xnor UO_1560 (O_1560,N_19502,N_19005);
or UO_1561 (O_1561,N_19659,N_19299);
xnor UO_1562 (O_1562,N_19300,N_19031);
xnor UO_1563 (O_1563,N_19283,N_19700);
xor UO_1564 (O_1564,N_18621,N_19870);
or UO_1565 (O_1565,N_19423,N_19806);
nand UO_1566 (O_1566,N_18398,N_19194);
or UO_1567 (O_1567,N_19515,N_18914);
xor UO_1568 (O_1568,N_18329,N_18635);
and UO_1569 (O_1569,N_18051,N_18420);
xor UO_1570 (O_1570,N_18432,N_19145);
and UO_1571 (O_1571,N_18046,N_18555);
nor UO_1572 (O_1572,N_19147,N_18597);
xnor UO_1573 (O_1573,N_18905,N_19195);
and UO_1574 (O_1574,N_18247,N_18285);
and UO_1575 (O_1575,N_18871,N_19874);
and UO_1576 (O_1576,N_19309,N_19051);
xor UO_1577 (O_1577,N_19686,N_19242);
nand UO_1578 (O_1578,N_19083,N_18000);
nand UO_1579 (O_1579,N_19748,N_18219);
nand UO_1580 (O_1580,N_18333,N_18358);
or UO_1581 (O_1581,N_19003,N_18093);
or UO_1582 (O_1582,N_19862,N_19063);
xor UO_1583 (O_1583,N_19632,N_19007);
nand UO_1584 (O_1584,N_18115,N_18494);
nor UO_1585 (O_1585,N_18303,N_19409);
or UO_1586 (O_1586,N_18225,N_19101);
nand UO_1587 (O_1587,N_18099,N_19239);
or UO_1588 (O_1588,N_18954,N_18641);
and UO_1589 (O_1589,N_19644,N_19412);
xor UO_1590 (O_1590,N_19234,N_19811);
nor UO_1591 (O_1591,N_18031,N_19855);
and UO_1592 (O_1592,N_19666,N_18258);
nand UO_1593 (O_1593,N_18603,N_18490);
or UO_1594 (O_1594,N_19218,N_19015);
xor UO_1595 (O_1595,N_18324,N_19142);
xor UO_1596 (O_1596,N_18891,N_18070);
and UO_1597 (O_1597,N_19880,N_19882);
or UO_1598 (O_1598,N_19401,N_19797);
and UO_1599 (O_1599,N_18025,N_18976);
nor UO_1600 (O_1600,N_19997,N_19646);
and UO_1601 (O_1601,N_19974,N_19211);
nand UO_1602 (O_1602,N_19051,N_18135);
or UO_1603 (O_1603,N_19658,N_18111);
nand UO_1604 (O_1604,N_19854,N_18044);
nor UO_1605 (O_1605,N_19856,N_18663);
xnor UO_1606 (O_1606,N_19806,N_18140);
or UO_1607 (O_1607,N_18411,N_19023);
nor UO_1608 (O_1608,N_19629,N_19908);
xnor UO_1609 (O_1609,N_19791,N_18098);
xnor UO_1610 (O_1610,N_19492,N_19369);
nand UO_1611 (O_1611,N_18520,N_18445);
and UO_1612 (O_1612,N_19318,N_19512);
nor UO_1613 (O_1613,N_19197,N_19819);
and UO_1614 (O_1614,N_18169,N_19889);
nor UO_1615 (O_1615,N_19853,N_18207);
and UO_1616 (O_1616,N_18933,N_19012);
xnor UO_1617 (O_1617,N_19698,N_19033);
and UO_1618 (O_1618,N_19042,N_19129);
nand UO_1619 (O_1619,N_19560,N_19200);
nor UO_1620 (O_1620,N_19848,N_18513);
or UO_1621 (O_1621,N_18176,N_18957);
xnor UO_1622 (O_1622,N_18077,N_19266);
xor UO_1623 (O_1623,N_18910,N_18121);
xor UO_1624 (O_1624,N_18353,N_19278);
or UO_1625 (O_1625,N_18628,N_18285);
nor UO_1626 (O_1626,N_18972,N_18672);
and UO_1627 (O_1627,N_19972,N_19048);
nor UO_1628 (O_1628,N_19240,N_18048);
nand UO_1629 (O_1629,N_19425,N_19314);
nand UO_1630 (O_1630,N_19473,N_18753);
nand UO_1631 (O_1631,N_19557,N_18655);
and UO_1632 (O_1632,N_18759,N_18884);
and UO_1633 (O_1633,N_19910,N_18014);
nor UO_1634 (O_1634,N_19349,N_19630);
nor UO_1635 (O_1635,N_18377,N_19154);
nor UO_1636 (O_1636,N_18700,N_18678);
nor UO_1637 (O_1637,N_19623,N_18435);
and UO_1638 (O_1638,N_18299,N_19228);
and UO_1639 (O_1639,N_19262,N_18207);
nor UO_1640 (O_1640,N_19285,N_19023);
nor UO_1641 (O_1641,N_19273,N_19897);
nor UO_1642 (O_1642,N_19925,N_19755);
xnor UO_1643 (O_1643,N_18506,N_18359);
and UO_1644 (O_1644,N_19802,N_18505);
or UO_1645 (O_1645,N_18109,N_18913);
xor UO_1646 (O_1646,N_18845,N_18216);
and UO_1647 (O_1647,N_19115,N_18807);
or UO_1648 (O_1648,N_18807,N_19957);
or UO_1649 (O_1649,N_19713,N_18334);
and UO_1650 (O_1650,N_18159,N_18560);
and UO_1651 (O_1651,N_19464,N_19366);
nand UO_1652 (O_1652,N_19716,N_19918);
or UO_1653 (O_1653,N_18018,N_18276);
or UO_1654 (O_1654,N_19273,N_19994);
nand UO_1655 (O_1655,N_19458,N_18604);
xnor UO_1656 (O_1656,N_18303,N_19312);
or UO_1657 (O_1657,N_19465,N_18971);
nand UO_1658 (O_1658,N_18129,N_19278);
or UO_1659 (O_1659,N_19083,N_18582);
xnor UO_1660 (O_1660,N_18819,N_18641);
or UO_1661 (O_1661,N_19588,N_18838);
nor UO_1662 (O_1662,N_19276,N_19223);
and UO_1663 (O_1663,N_19161,N_18484);
and UO_1664 (O_1664,N_18343,N_18752);
xor UO_1665 (O_1665,N_19080,N_18181);
nor UO_1666 (O_1666,N_18695,N_19632);
nor UO_1667 (O_1667,N_18881,N_18526);
and UO_1668 (O_1668,N_19366,N_18120);
or UO_1669 (O_1669,N_18408,N_18219);
nor UO_1670 (O_1670,N_19293,N_18548);
or UO_1671 (O_1671,N_18619,N_19858);
and UO_1672 (O_1672,N_18147,N_18947);
xor UO_1673 (O_1673,N_18929,N_19031);
and UO_1674 (O_1674,N_19083,N_18907);
and UO_1675 (O_1675,N_18168,N_19846);
nand UO_1676 (O_1676,N_18684,N_19569);
nand UO_1677 (O_1677,N_19203,N_19937);
nand UO_1678 (O_1678,N_18417,N_18877);
or UO_1679 (O_1679,N_19736,N_18621);
and UO_1680 (O_1680,N_18517,N_19519);
or UO_1681 (O_1681,N_18443,N_19477);
or UO_1682 (O_1682,N_18862,N_19814);
nand UO_1683 (O_1683,N_19005,N_18973);
and UO_1684 (O_1684,N_18676,N_18871);
or UO_1685 (O_1685,N_18163,N_18557);
or UO_1686 (O_1686,N_19128,N_18795);
or UO_1687 (O_1687,N_18135,N_19303);
nand UO_1688 (O_1688,N_18864,N_18193);
or UO_1689 (O_1689,N_19130,N_18469);
or UO_1690 (O_1690,N_18874,N_18389);
nand UO_1691 (O_1691,N_18397,N_19687);
nor UO_1692 (O_1692,N_18166,N_18824);
nand UO_1693 (O_1693,N_18436,N_18128);
or UO_1694 (O_1694,N_18118,N_18721);
nor UO_1695 (O_1695,N_18958,N_19404);
nand UO_1696 (O_1696,N_19232,N_18733);
nor UO_1697 (O_1697,N_19348,N_19943);
and UO_1698 (O_1698,N_18069,N_19449);
nand UO_1699 (O_1699,N_19834,N_18738);
or UO_1700 (O_1700,N_19135,N_18959);
xor UO_1701 (O_1701,N_18551,N_18512);
and UO_1702 (O_1702,N_18914,N_18088);
or UO_1703 (O_1703,N_19362,N_19053);
and UO_1704 (O_1704,N_19980,N_19973);
xor UO_1705 (O_1705,N_19369,N_18814);
nor UO_1706 (O_1706,N_18926,N_18831);
nor UO_1707 (O_1707,N_19377,N_18956);
nor UO_1708 (O_1708,N_19307,N_18022);
nor UO_1709 (O_1709,N_18720,N_19040);
xnor UO_1710 (O_1710,N_18008,N_18936);
nand UO_1711 (O_1711,N_19408,N_18850);
xor UO_1712 (O_1712,N_18042,N_19557);
nor UO_1713 (O_1713,N_18364,N_19891);
and UO_1714 (O_1714,N_18784,N_18193);
nand UO_1715 (O_1715,N_19607,N_19040);
nand UO_1716 (O_1716,N_19585,N_18860);
and UO_1717 (O_1717,N_19763,N_19659);
xnor UO_1718 (O_1718,N_19122,N_19509);
and UO_1719 (O_1719,N_19580,N_18974);
xnor UO_1720 (O_1720,N_19145,N_18349);
nand UO_1721 (O_1721,N_18101,N_18772);
and UO_1722 (O_1722,N_19910,N_19726);
and UO_1723 (O_1723,N_19193,N_18424);
xnor UO_1724 (O_1724,N_18859,N_19430);
and UO_1725 (O_1725,N_19379,N_19899);
nand UO_1726 (O_1726,N_18055,N_18528);
nor UO_1727 (O_1727,N_19833,N_18054);
or UO_1728 (O_1728,N_19126,N_18955);
nor UO_1729 (O_1729,N_18590,N_18667);
and UO_1730 (O_1730,N_19799,N_19616);
or UO_1731 (O_1731,N_18406,N_18232);
or UO_1732 (O_1732,N_18380,N_18709);
and UO_1733 (O_1733,N_19982,N_19173);
xnor UO_1734 (O_1734,N_18921,N_18327);
or UO_1735 (O_1735,N_18567,N_18454);
or UO_1736 (O_1736,N_18849,N_19658);
nand UO_1737 (O_1737,N_18196,N_19703);
or UO_1738 (O_1738,N_18809,N_19428);
or UO_1739 (O_1739,N_18899,N_18535);
nor UO_1740 (O_1740,N_18447,N_18208);
nand UO_1741 (O_1741,N_19686,N_19434);
or UO_1742 (O_1742,N_18219,N_19279);
or UO_1743 (O_1743,N_18536,N_18236);
or UO_1744 (O_1744,N_18110,N_18221);
nand UO_1745 (O_1745,N_18467,N_18730);
and UO_1746 (O_1746,N_18177,N_18986);
and UO_1747 (O_1747,N_18174,N_18195);
nor UO_1748 (O_1748,N_18177,N_19945);
nand UO_1749 (O_1749,N_19897,N_19807);
or UO_1750 (O_1750,N_18167,N_19449);
xnor UO_1751 (O_1751,N_18324,N_19615);
xnor UO_1752 (O_1752,N_19043,N_18506);
nor UO_1753 (O_1753,N_19234,N_19164);
xnor UO_1754 (O_1754,N_18397,N_19927);
nor UO_1755 (O_1755,N_19121,N_19443);
and UO_1756 (O_1756,N_18509,N_19733);
and UO_1757 (O_1757,N_19703,N_19261);
and UO_1758 (O_1758,N_19390,N_18005);
nor UO_1759 (O_1759,N_18894,N_18537);
xor UO_1760 (O_1760,N_19448,N_19641);
nor UO_1761 (O_1761,N_19186,N_19709);
xnor UO_1762 (O_1762,N_18334,N_19028);
nand UO_1763 (O_1763,N_19880,N_18062);
nor UO_1764 (O_1764,N_18180,N_19514);
and UO_1765 (O_1765,N_18519,N_19247);
nand UO_1766 (O_1766,N_18197,N_18846);
or UO_1767 (O_1767,N_19189,N_19669);
or UO_1768 (O_1768,N_18666,N_18300);
nor UO_1769 (O_1769,N_19868,N_19414);
xor UO_1770 (O_1770,N_19669,N_18385);
nand UO_1771 (O_1771,N_19845,N_18496);
and UO_1772 (O_1772,N_18422,N_18418);
nand UO_1773 (O_1773,N_18377,N_18371);
nor UO_1774 (O_1774,N_19209,N_19899);
or UO_1775 (O_1775,N_18174,N_19332);
xor UO_1776 (O_1776,N_18119,N_18599);
nand UO_1777 (O_1777,N_19343,N_18618);
nor UO_1778 (O_1778,N_19058,N_19632);
nand UO_1779 (O_1779,N_18925,N_19095);
xor UO_1780 (O_1780,N_19283,N_18788);
nand UO_1781 (O_1781,N_18596,N_19546);
xnor UO_1782 (O_1782,N_19426,N_18029);
xor UO_1783 (O_1783,N_19482,N_18670);
or UO_1784 (O_1784,N_18851,N_18987);
xor UO_1785 (O_1785,N_18822,N_18512);
xor UO_1786 (O_1786,N_19159,N_18514);
nand UO_1787 (O_1787,N_19467,N_18504);
nand UO_1788 (O_1788,N_19821,N_18181);
and UO_1789 (O_1789,N_18012,N_18653);
xnor UO_1790 (O_1790,N_19867,N_19349);
nand UO_1791 (O_1791,N_18055,N_18977);
xor UO_1792 (O_1792,N_19627,N_19123);
and UO_1793 (O_1793,N_19979,N_19530);
nand UO_1794 (O_1794,N_18045,N_19879);
nor UO_1795 (O_1795,N_19077,N_19309);
and UO_1796 (O_1796,N_19143,N_19927);
nand UO_1797 (O_1797,N_19556,N_19199);
or UO_1798 (O_1798,N_18198,N_19456);
nand UO_1799 (O_1799,N_18723,N_19201);
or UO_1800 (O_1800,N_18156,N_19246);
and UO_1801 (O_1801,N_19458,N_18655);
nand UO_1802 (O_1802,N_18510,N_19507);
nor UO_1803 (O_1803,N_19210,N_18073);
nand UO_1804 (O_1804,N_18024,N_19290);
and UO_1805 (O_1805,N_18204,N_18391);
nand UO_1806 (O_1806,N_18944,N_19394);
or UO_1807 (O_1807,N_18977,N_19764);
or UO_1808 (O_1808,N_19359,N_18875);
or UO_1809 (O_1809,N_18726,N_19044);
nor UO_1810 (O_1810,N_18732,N_18438);
and UO_1811 (O_1811,N_19966,N_18245);
nor UO_1812 (O_1812,N_18472,N_19211);
nor UO_1813 (O_1813,N_18410,N_19706);
nand UO_1814 (O_1814,N_18320,N_19426);
nand UO_1815 (O_1815,N_18926,N_19418);
xnor UO_1816 (O_1816,N_18159,N_18249);
and UO_1817 (O_1817,N_18581,N_18634);
xnor UO_1818 (O_1818,N_19663,N_19873);
xnor UO_1819 (O_1819,N_19086,N_18609);
nand UO_1820 (O_1820,N_18407,N_18083);
nand UO_1821 (O_1821,N_19912,N_19286);
nor UO_1822 (O_1822,N_19144,N_18487);
and UO_1823 (O_1823,N_18442,N_18452);
nand UO_1824 (O_1824,N_18169,N_19739);
nor UO_1825 (O_1825,N_19966,N_19424);
xnor UO_1826 (O_1826,N_18549,N_19605);
nand UO_1827 (O_1827,N_19372,N_19227);
and UO_1828 (O_1828,N_18243,N_19064);
nor UO_1829 (O_1829,N_18361,N_18404);
or UO_1830 (O_1830,N_18138,N_18160);
nand UO_1831 (O_1831,N_19299,N_18465);
and UO_1832 (O_1832,N_18284,N_19530);
nor UO_1833 (O_1833,N_18497,N_19038);
or UO_1834 (O_1834,N_18617,N_18318);
and UO_1835 (O_1835,N_19772,N_18980);
xor UO_1836 (O_1836,N_18809,N_19137);
xor UO_1837 (O_1837,N_19306,N_18684);
nand UO_1838 (O_1838,N_19454,N_19359);
or UO_1839 (O_1839,N_18723,N_19184);
nor UO_1840 (O_1840,N_19472,N_18863);
nand UO_1841 (O_1841,N_19825,N_18635);
or UO_1842 (O_1842,N_18081,N_19681);
nor UO_1843 (O_1843,N_19337,N_19929);
and UO_1844 (O_1844,N_19664,N_18987);
xnor UO_1845 (O_1845,N_18816,N_18723);
nor UO_1846 (O_1846,N_19032,N_19149);
and UO_1847 (O_1847,N_19900,N_19517);
or UO_1848 (O_1848,N_18174,N_19759);
nor UO_1849 (O_1849,N_19201,N_18350);
or UO_1850 (O_1850,N_18917,N_19244);
nand UO_1851 (O_1851,N_18923,N_19309);
xor UO_1852 (O_1852,N_19571,N_18295);
xnor UO_1853 (O_1853,N_19942,N_18672);
nand UO_1854 (O_1854,N_18915,N_19809);
and UO_1855 (O_1855,N_18254,N_18025);
and UO_1856 (O_1856,N_19237,N_19435);
xnor UO_1857 (O_1857,N_19974,N_19262);
xor UO_1858 (O_1858,N_18000,N_19470);
xnor UO_1859 (O_1859,N_19420,N_18338);
or UO_1860 (O_1860,N_19334,N_18547);
nand UO_1861 (O_1861,N_19909,N_19658);
and UO_1862 (O_1862,N_19655,N_18825);
xnor UO_1863 (O_1863,N_19797,N_19026);
and UO_1864 (O_1864,N_19920,N_19863);
and UO_1865 (O_1865,N_19542,N_19551);
and UO_1866 (O_1866,N_19325,N_19419);
xor UO_1867 (O_1867,N_19186,N_18881);
nand UO_1868 (O_1868,N_18388,N_19984);
xnor UO_1869 (O_1869,N_19925,N_18683);
nor UO_1870 (O_1870,N_18976,N_19544);
or UO_1871 (O_1871,N_19062,N_18413);
and UO_1872 (O_1872,N_18557,N_18695);
nor UO_1873 (O_1873,N_19532,N_18484);
or UO_1874 (O_1874,N_19222,N_19296);
or UO_1875 (O_1875,N_18708,N_18245);
xnor UO_1876 (O_1876,N_19944,N_18290);
or UO_1877 (O_1877,N_19001,N_18049);
nor UO_1878 (O_1878,N_18838,N_19867);
nand UO_1879 (O_1879,N_19527,N_18810);
nor UO_1880 (O_1880,N_18284,N_19445);
and UO_1881 (O_1881,N_19514,N_19942);
xnor UO_1882 (O_1882,N_18501,N_19522);
nor UO_1883 (O_1883,N_18493,N_18300);
nor UO_1884 (O_1884,N_19853,N_18962);
nand UO_1885 (O_1885,N_18977,N_19363);
nor UO_1886 (O_1886,N_18993,N_19194);
xnor UO_1887 (O_1887,N_18074,N_18067);
nand UO_1888 (O_1888,N_18326,N_18680);
xor UO_1889 (O_1889,N_19218,N_18571);
and UO_1890 (O_1890,N_19650,N_18321);
xnor UO_1891 (O_1891,N_19949,N_18727);
xor UO_1892 (O_1892,N_19414,N_18111);
nor UO_1893 (O_1893,N_19041,N_19005);
or UO_1894 (O_1894,N_18330,N_19669);
nand UO_1895 (O_1895,N_18015,N_19328);
xnor UO_1896 (O_1896,N_18493,N_19526);
nand UO_1897 (O_1897,N_19833,N_18660);
or UO_1898 (O_1898,N_18960,N_18911);
or UO_1899 (O_1899,N_19746,N_18598);
and UO_1900 (O_1900,N_19799,N_19195);
and UO_1901 (O_1901,N_18877,N_18443);
and UO_1902 (O_1902,N_19679,N_19672);
or UO_1903 (O_1903,N_19049,N_19007);
xnor UO_1904 (O_1904,N_19557,N_19774);
and UO_1905 (O_1905,N_19778,N_18098);
nand UO_1906 (O_1906,N_19545,N_18450);
xnor UO_1907 (O_1907,N_19239,N_19005);
xor UO_1908 (O_1908,N_19642,N_19051);
or UO_1909 (O_1909,N_19873,N_18010);
and UO_1910 (O_1910,N_18830,N_18811);
and UO_1911 (O_1911,N_18162,N_18183);
nand UO_1912 (O_1912,N_19064,N_18270);
or UO_1913 (O_1913,N_19218,N_19079);
nand UO_1914 (O_1914,N_18473,N_18500);
nand UO_1915 (O_1915,N_18808,N_19552);
and UO_1916 (O_1916,N_19463,N_18971);
nor UO_1917 (O_1917,N_19071,N_18103);
and UO_1918 (O_1918,N_18234,N_19488);
and UO_1919 (O_1919,N_18604,N_18380);
or UO_1920 (O_1920,N_18117,N_18981);
and UO_1921 (O_1921,N_19419,N_19438);
nand UO_1922 (O_1922,N_19972,N_19543);
and UO_1923 (O_1923,N_19491,N_18761);
or UO_1924 (O_1924,N_19680,N_18831);
nand UO_1925 (O_1925,N_19870,N_18646);
nor UO_1926 (O_1926,N_19826,N_18479);
xor UO_1927 (O_1927,N_19291,N_18759);
nand UO_1928 (O_1928,N_19303,N_19705);
nor UO_1929 (O_1929,N_18098,N_19991);
xor UO_1930 (O_1930,N_18014,N_18343);
xor UO_1931 (O_1931,N_18938,N_18352);
and UO_1932 (O_1932,N_18140,N_18261);
nor UO_1933 (O_1933,N_19850,N_18152);
and UO_1934 (O_1934,N_19613,N_19840);
nor UO_1935 (O_1935,N_19079,N_19893);
nor UO_1936 (O_1936,N_19581,N_19777);
xor UO_1937 (O_1937,N_18481,N_19578);
nor UO_1938 (O_1938,N_18250,N_19076);
nand UO_1939 (O_1939,N_19962,N_19335);
or UO_1940 (O_1940,N_19020,N_18285);
nand UO_1941 (O_1941,N_19510,N_18514);
and UO_1942 (O_1942,N_19717,N_18800);
and UO_1943 (O_1943,N_19546,N_19290);
nand UO_1944 (O_1944,N_18951,N_19979);
nor UO_1945 (O_1945,N_18359,N_19903);
nor UO_1946 (O_1946,N_19482,N_19856);
nor UO_1947 (O_1947,N_18932,N_18492);
or UO_1948 (O_1948,N_19489,N_19809);
nor UO_1949 (O_1949,N_19010,N_18111);
or UO_1950 (O_1950,N_18390,N_18071);
or UO_1951 (O_1951,N_18522,N_19369);
or UO_1952 (O_1952,N_19967,N_19341);
nor UO_1953 (O_1953,N_18853,N_19628);
or UO_1954 (O_1954,N_18303,N_18231);
or UO_1955 (O_1955,N_18070,N_18811);
and UO_1956 (O_1956,N_19752,N_18739);
nand UO_1957 (O_1957,N_19962,N_18895);
nand UO_1958 (O_1958,N_19096,N_19789);
nand UO_1959 (O_1959,N_18991,N_18604);
xnor UO_1960 (O_1960,N_18698,N_19946);
nor UO_1961 (O_1961,N_19120,N_18137);
nand UO_1962 (O_1962,N_18950,N_18455);
xor UO_1963 (O_1963,N_19478,N_19284);
and UO_1964 (O_1964,N_18390,N_18392);
nand UO_1965 (O_1965,N_18959,N_18498);
or UO_1966 (O_1966,N_18044,N_18679);
xnor UO_1967 (O_1967,N_18395,N_19958);
nor UO_1968 (O_1968,N_18903,N_18574);
or UO_1969 (O_1969,N_18295,N_19982);
and UO_1970 (O_1970,N_18015,N_18294);
nand UO_1971 (O_1971,N_18286,N_18562);
and UO_1972 (O_1972,N_19348,N_19842);
nand UO_1973 (O_1973,N_19963,N_18026);
nor UO_1974 (O_1974,N_18465,N_18010);
nor UO_1975 (O_1975,N_18921,N_18093);
and UO_1976 (O_1976,N_18314,N_18229);
nor UO_1977 (O_1977,N_18521,N_18549);
xor UO_1978 (O_1978,N_19463,N_18719);
nand UO_1979 (O_1979,N_18552,N_19089);
xor UO_1980 (O_1980,N_18770,N_19228);
xor UO_1981 (O_1981,N_18921,N_18594);
nor UO_1982 (O_1982,N_19327,N_18169);
nand UO_1983 (O_1983,N_18381,N_19551);
or UO_1984 (O_1984,N_18741,N_19954);
xnor UO_1985 (O_1985,N_18798,N_18678);
nand UO_1986 (O_1986,N_19051,N_18904);
xor UO_1987 (O_1987,N_19906,N_19801);
xnor UO_1988 (O_1988,N_19863,N_19410);
nand UO_1989 (O_1989,N_19582,N_19383);
xnor UO_1990 (O_1990,N_19041,N_19815);
or UO_1991 (O_1991,N_18773,N_18132);
nor UO_1992 (O_1992,N_19382,N_19803);
or UO_1993 (O_1993,N_19440,N_18241);
nor UO_1994 (O_1994,N_19524,N_18379);
nor UO_1995 (O_1995,N_19337,N_18119);
nand UO_1996 (O_1996,N_19504,N_19632);
or UO_1997 (O_1997,N_18370,N_19968);
nand UO_1998 (O_1998,N_18747,N_19299);
xor UO_1999 (O_1999,N_19018,N_18435);
nor UO_2000 (O_2000,N_19140,N_18083);
and UO_2001 (O_2001,N_19349,N_18496);
or UO_2002 (O_2002,N_19452,N_19445);
nor UO_2003 (O_2003,N_18150,N_18903);
and UO_2004 (O_2004,N_18541,N_18399);
and UO_2005 (O_2005,N_18140,N_19260);
or UO_2006 (O_2006,N_19377,N_18233);
nor UO_2007 (O_2007,N_19279,N_19572);
and UO_2008 (O_2008,N_19795,N_18045);
or UO_2009 (O_2009,N_19826,N_19960);
xor UO_2010 (O_2010,N_19406,N_19700);
nand UO_2011 (O_2011,N_19410,N_19198);
and UO_2012 (O_2012,N_18549,N_18204);
nor UO_2013 (O_2013,N_18195,N_19412);
nand UO_2014 (O_2014,N_18699,N_18460);
xor UO_2015 (O_2015,N_19661,N_18940);
nor UO_2016 (O_2016,N_19878,N_19155);
and UO_2017 (O_2017,N_19526,N_19992);
nand UO_2018 (O_2018,N_18809,N_18299);
xnor UO_2019 (O_2019,N_18093,N_19094);
or UO_2020 (O_2020,N_19970,N_19827);
nor UO_2021 (O_2021,N_19054,N_18077);
and UO_2022 (O_2022,N_18447,N_19160);
and UO_2023 (O_2023,N_18250,N_19481);
or UO_2024 (O_2024,N_19778,N_19935);
nor UO_2025 (O_2025,N_19207,N_19028);
or UO_2026 (O_2026,N_19302,N_19007);
or UO_2027 (O_2027,N_18765,N_19125);
nor UO_2028 (O_2028,N_19756,N_18095);
nand UO_2029 (O_2029,N_18120,N_18093);
nor UO_2030 (O_2030,N_19797,N_18570);
xor UO_2031 (O_2031,N_18952,N_18885);
and UO_2032 (O_2032,N_18964,N_19806);
xor UO_2033 (O_2033,N_19694,N_19317);
xnor UO_2034 (O_2034,N_18490,N_19138);
nor UO_2035 (O_2035,N_18351,N_18865);
xor UO_2036 (O_2036,N_19577,N_18715);
nor UO_2037 (O_2037,N_18032,N_19393);
or UO_2038 (O_2038,N_19045,N_19945);
xor UO_2039 (O_2039,N_19984,N_19959);
nand UO_2040 (O_2040,N_19448,N_18654);
and UO_2041 (O_2041,N_18808,N_19382);
nor UO_2042 (O_2042,N_18269,N_19557);
and UO_2043 (O_2043,N_18505,N_18581);
nand UO_2044 (O_2044,N_19641,N_18218);
nand UO_2045 (O_2045,N_19024,N_19844);
nand UO_2046 (O_2046,N_19127,N_19685);
and UO_2047 (O_2047,N_19751,N_19322);
or UO_2048 (O_2048,N_19676,N_19561);
xnor UO_2049 (O_2049,N_19910,N_18551);
nor UO_2050 (O_2050,N_18788,N_18772);
nor UO_2051 (O_2051,N_18338,N_18330);
or UO_2052 (O_2052,N_19610,N_19237);
nor UO_2053 (O_2053,N_18046,N_19770);
nand UO_2054 (O_2054,N_18574,N_18174);
xor UO_2055 (O_2055,N_18643,N_18604);
nand UO_2056 (O_2056,N_19649,N_19671);
xnor UO_2057 (O_2057,N_18974,N_19911);
or UO_2058 (O_2058,N_19349,N_18422);
xor UO_2059 (O_2059,N_19324,N_18786);
xnor UO_2060 (O_2060,N_18406,N_19146);
nand UO_2061 (O_2061,N_18986,N_18157);
or UO_2062 (O_2062,N_19914,N_19470);
or UO_2063 (O_2063,N_18446,N_18971);
xnor UO_2064 (O_2064,N_19791,N_19216);
xor UO_2065 (O_2065,N_18656,N_18070);
xnor UO_2066 (O_2066,N_18238,N_18754);
xor UO_2067 (O_2067,N_19177,N_19676);
and UO_2068 (O_2068,N_19885,N_18712);
nor UO_2069 (O_2069,N_18844,N_18065);
and UO_2070 (O_2070,N_19110,N_19380);
nor UO_2071 (O_2071,N_18193,N_19315);
xor UO_2072 (O_2072,N_19447,N_18756);
and UO_2073 (O_2073,N_19617,N_19395);
nand UO_2074 (O_2074,N_19647,N_18496);
nand UO_2075 (O_2075,N_19867,N_19933);
xnor UO_2076 (O_2076,N_19131,N_18137);
nand UO_2077 (O_2077,N_19591,N_19710);
nand UO_2078 (O_2078,N_19312,N_18604);
xor UO_2079 (O_2079,N_18829,N_19322);
nor UO_2080 (O_2080,N_18377,N_19677);
xnor UO_2081 (O_2081,N_18344,N_18893);
nand UO_2082 (O_2082,N_19759,N_19932);
nor UO_2083 (O_2083,N_19237,N_18811);
nand UO_2084 (O_2084,N_18837,N_19730);
and UO_2085 (O_2085,N_19244,N_18463);
nand UO_2086 (O_2086,N_19702,N_18172);
xor UO_2087 (O_2087,N_19274,N_19661);
nand UO_2088 (O_2088,N_18797,N_19388);
nor UO_2089 (O_2089,N_19509,N_19988);
or UO_2090 (O_2090,N_18809,N_18633);
nand UO_2091 (O_2091,N_18146,N_19111);
nand UO_2092 (O_2092,N_19667,N_18121);
xnor UO_2093 (O_2093,N_18868,N_18124);
and UO_2094 (O_2094,N_18765,N_19335);
xnor UO_2095 (O_2095,N_18247,N_19987);
nor UO_2096 (O_2096,N_19920,N_18461);
nand UO_2097 (O_2097,N_19017,N_18266);
nor UO_2098 (O_2098,N_18763,N_19746);
and UO_2099 (O_2099,N_19124,N_18677);
and UO_2100 (O_2100,N_18831,N_19490);
and UO_2101 (O_2101,N_18449,N_19406);
xnor UO_2102 (O_2102,N_18862,N_18624);
xnor UO_2103 (O_2103,N_19112,N_18807);
and UO_2104 (O_2104,N_18179,N_18909);
nor UO_2105 (O_2105,N_19967,N_19816);
nand UO_2106 (O_2106,N_18990,N_18936);
and UO_2107 (O_2107,N_19023,N_19038);
or UO_2108 (O_2108,N_19017,N_19185);
or UO_2109 (O_2109,N_19765,N_18579);
nor UO_2110 (O_2110,N_18047,N_19751);
or UO_2111 (O_2111,N_18622,N_19683);
and UO_2112 (O_2112,N_18125,N_18486);
or UO_2113 (O_2113,N_18065,N_19468);
or UO_2114 (O_2114,N_18529,N_19922);
nand UO_2115 (O_2115,N_18966,N_19304);
and UO_2116 (O_2116,N_18176,N_18204);
or UO_2117 (O_2117,N_18213,N_18798);
or UO_2118 (O_2118,N_18545,N_19895);
nand UO_2119 (O_2119,N_18192,N_18515);
or UO_2120 (O_2120,N_19209,N_18687);
xnor UO_2121 (O_2121,N_18669,N_19983);
nor UO_2122 (O_2122,N_18763,N_19292);
and UO_2123 (O_2123,N_18385,N_19463);
nor UO_2124 (O_2124,N_18099,N_19021);
xor UO_2125 (O_2125,N_19075,N_18781);
nor UO_2126 (O_2126,N_19327,N_18552);
nor UO_2127 (O_2127,N_18019,N_18410);
xor UO_2128 (O_2128,N_19081,N_19603);
xor UO_2129 (O_2129,N_19168,N_18590);
xnor UO_2130 (O_2130,N_19525,N_18908);
xnor UO_2131 (O_2131,N_18545,N_19130);
and UO_2132 (O_2132,N_18348,N_18954);
or UO_2133 (O_2133,N_19939,N_19270);
xor UO_2134 (O_2134,N_19619,N_18041);
and UO_2135 (O_2135,N_19964,N_19540);
nand UO_2136 (O_2136,N_18526,N_18506);
or UO_2137 (O_2137,N_18806,N_19681);
xor UO_2138 (O_2138,N_19189,N_18148);
nand UO_2139 (O_2139,N_19676,N_19453);
or UO_2140 (O_2140,N_18253,N_18207);
or UO_2141 (O_2141,N_19026,N_19214);
xnor UO_2142 (O_2142,N_19845,N_18887);
xor UO_2143 (O_2143,N_19567,N_18537);
or UO_2144 (O_2144,N_19959,N_18712);
or UO_2145 (O_2145,N_19593,N_18700);
and UO_2146 (O_2146,N_19613,N_19102);
xnor UO_2147 (O_2147,N_19161,N_18703);
nor UO_2148 (O_2148,N_18353,N_18003);
and UO_2149 (O_2149,N_18665,N_19353);
xnor UO_2150 (O_2150,N_19136,N_19359);
or UO_2151 (O_2151,N_18868,N_18506);
nor UO_2152 (O_2152,N_19312,N_19625);
nor UO_2153 (O_2153,N_18309,N_19147);
nor UO_2154 (O_2154,N_18108,N_18586);
xnor UO_2155 (O_2155,N_19969,N_19975);
nand UO_2156 (O_2156,N_18013,N_19932);
or UO_2157 (O_2157,N_19528,N_19347);
nand UO_2158 (O_2158,N_18478,N_19559);
and UO_2159 (O_2159,N_18330,N_18258);
or UO_2160 (O_2160,N_18686,N_18092);
and UO_2161 (O_2161,N_18889,N_18763);
and UO_2162 (O_2162,N_18544,N_19205);
and UO_2163 (O_2163,N_19684,N_19230);
nand UO_2164 (O_2164,N_19011,N_19442);
nor UO_2165 (O_2165,N_18285,N_18827);
or UO_2166 (O_2166,N_18199,N_18128);
xor UO_2167 (O_2167,N_19776,N_18214);
xor UO_2168 (O_2168,N_19907,N_19890);
xnor UO_2169 (O_2169,N_19992,N_18178);
nand UO_2170 (O_2170,N_19062,N_18549);
or UO_2171 (O_2171,N_19481,N_19429);
xnor UO_2172 (O_2172,N_18412,N_19454);
xnor UO_2173 (O_2173,N_18507,N_18017);
xor UO_2174 (O_2174,N_19487,N_19763);
and UO_2175 (O_2175,N_18174,N_19682);
or UO_2176 (O_2176,N_19744,N_18042);
xor UO_2177 (O_2177,N_19437,N_19440);
nor UO_2178 (O_2178,N_19838,N_18928);
xor UO_2179 (O_2179,N_19280,N_19294);
and UO_2180 (O_2180,N_18817,N_19809);
nor UO_2181 (O_2181,N_18894,N_18987);
nand UO_2182 (O_2182,N_18716,N_18656);
and UO_2183 (O_2183,N_19844,N_19730);
nor UO_2184 (O_2184,N_18799,N_18224);
xor UO_2185 (O_2185,N_19903,N_18054);
xnor UO_2186 (O_2186,N_19216,N_18577);
xor UO_2187 (O_2187,N_18738,N_19351);
and UO_2188 (O_2188,N_18556,N_19063);
xor UO_2189 (O_2189,N_18175,N_18299);
or UO_2190 (O_2190,N_19233,N_18507);
xor UO_2191 (O_2191,N_18951,N_19522);
xnor UO_2192 (O_2192,N_19146,N_18792);
nand UO_2193 (O_2193,N_18804,N_18315);
or UO_2194 (O_2194,N_19698,N_19512);
xnor UO_2195 (O_2195,N_19619,N_19108);
xnor UO_2196 (O_2196,N_18261,N_18547);
xnor UO_2197 (O_2197,N_18997,N_18745);
or UO_2198 (O_2198,N_19700,N_19048);
xnor UO_2199 (O_2199,N_18361,N_18812);
nor UO_2200 (O_2200,N_19075,N_18686);
nor UO_2201 (O_2201,N_19947,N_18218);
nor UO_2202 (O_2202,N_19734,N_19633);
xor UO_2203 (O_2203,N_18152,N_19747);
nor UO_2204 (O_2204,N_18176,N_18615);
xor UO_2205 (O_2205,N_18353,N_19041);
and UO_2206 (O_2206,N_18224,N_18400);
xor UO_2207 (O_2207,N_19426,N_19336);
nand UO_2208 (O_2208,N_18526,N_19040);
xnor UO_2209 (O_2209,N_18219,N_19484);
nand UO_2210 (O_2210,N_19211,N_18755);
and UO_2211 (O_2211,N_19663,N_18856);
nand UO_2212 (O_2212,N_19059,N_18189);
xnor UO_2213 (O_2213,N_18887,N_19872);
nor UO_2214 (O_2214,N_18814,N_18897);
nor UO_2215 (O_2215,N_18215,N_18135);
nor UO_2216 (O_2216,N_19159,N_18618);
nand UO_2217 (O_2217,N_18533,N_19089);
or UO_2218 (O_2218,N_18365,N_19640);
or UO_2219 (O_2219,N_18376,N_19692);
and UO_2220 (O_2220,N_18020,N_19028);
and UO_2221 (O_2221,N_19343,N_18029);
xor UO_2222 (O_2222,N_18693,N_19572);
and UO_2223 (O_2223,N_19496,N_19083);
or UO_2224 (O_2224,N_19055,N_19946);
nand UO_2225 (O_2225,N_19824,N_18159);
nand UO_2226 (O_2226,N_18773,N_18681);
or UO_2227 (O_2227,N_19086,N_19251);
nor UO_2228 (O_2228,N_19647,N_19365);
nand UO_2229 (O_2229,N_19350,N_18310);
and UO_2230 (O_2230,N_18887,N_18441);
nand UO_2231 (O_2231,N_19323,N_19107);
or UO_2232 (O_2232,N_19088,N_19157);
nand UO_2233 (O_2233,N_18020,N_19299);
or UO_2234 (O_2234,N_19814,N_18568);
nand UO_2235 (O_2235,N_19054,N_18585);
nor UO_2236 (O_2236,N_19687,N_19187);
nor UO_2237 (O_2237,N_19280,N_18753);
or UO_2238 (O_2238,N_18148,N_19692);
or UO_2239 (O_2239,N_19624,N_19765);
nand UO_2240 (O_2240,N_18881,N_18263);
nor UO_2241 (O_2241,N_19212,N_19868);
nand UO_2242 (O_2242,N_19267,N_19247);
xor UO_2243 (O_2243,N_19959,N_18540);
xor UO_2244 (O_2244,N_19508,N_18719);
xnor UO_2245 (O_2245,N_18438,N_19944);
nand UO_2246 (O_2246,N_18418,N_18289);
nand UO_2247 (O_2247,N_19520,N_19974);
nor UO_2248 (O_2248,N_19636,N_19134);
nor UO_2249 (O_2249,N_18559,N_18502);
and UO_2250 (O_2250,N_19052,N_18716);
xor UO_2251 (O_2251,N_18931,N_19157);
or UO_2252 (O_2252,N_18557,N_19295);
or UO_2253 (O_2253,N_19483,N_18831);
xor UO_2254 (O_2254,N_18392,N_19323);
nor UO_2255 (O_2255,N_19652,N_19038);
and UO_2256 (O_2256,N_18103,N_18346);
nand UO_2257 (O_2257,N_19966,N_18297);
nor UO_2258 (O_2258,N_18247,N_19794);
nand UO_2259 (O_2259,N_18778,N_19319);
nand UO_2260 (O_2260,N_19400,N_19177);
or UO_2261 (O_2261,N_18088,N_18851);
xor UO_2262 (O_2262,N_19790,N_18491);
xnor UO_2263 (O_2263,N_19806,N_18180);
nand UO_2264 (O_2264,N_18015,N_19837);
and UO_2265 (O_2265,N_18655,N_18142);
xor UO_2266 (O_2266,N_18689,N_19542);
or UO_2267 (O_2267,N_19271,N_18650);
nand UO_2268 (O_2268,N_18279,N_18948);
and UO_2269 (O_2269,N_19390,N_19900);
and UO_2270 (O_2270,N_18877,N_19353);
and UO_2271 (O_2271,N_18318,N_19082);
or UO_2272 (O_2272,N_18417,N_19299);
nor UO_2273 (O_2273,N_18292,N_19624);
nor UO_2274 (O_2274,N_18464,N_18641);
or UO_2275 (O_2275,N_18430,N_19218);
and UO_2276 (O_2276,N_19443,N_19036);
or UO_2277 (O_2277,N_19235,N_18330);
or UO_2278 (O_2278,N_19181,N_18163);
xnor UO_2279 (O_2279,N_19326,N_18409);
and UO_2280 (O_2280,N_19845,N_19161);
nand UO_2281 (O_2281,N_18077,N_19194);
and UO_2282 (O_2282,N_19027,N_18650);
and UO_2283 (O_2283,N_18310,N_18225);
or UO_2284 (O_2284,N_18386,N_18123);
and UO_2285 (O_2285,N_19528,N_18391);
nand UO_2286 (O_2286,N_18219,N_19466);
nor UO_2287 (O_2287,N_18700,N_18953);
or UO_2288 (O_2288,N_18030,N_19566);
and UO_2289 (O_2289,N_19409,N_18608);
nand UO_2290 (O_2290,N_19767,N_19094);
xnor UO_2291 (O_2291,N_19211,N_19680);
nand UO_2292 (O_2292,N_19573,N_18202);
nand UO_2293 (O_2293,N_19988,N_18123);
nor UO_2294 (O_2294,N_18687,N_19680);
xor UO_2295 (O_2295,N_19743,N_19553);
and UO_2296 (O_2296,N_19506,N_19249);
nand UO_2297 (O_2297,N_18800,N_19285);
nor UO_2298 (O_2298,N_19208,N_18615);
nor UO_2299 (O_2299,N_18867,N_19838);
and UO_2300 (O_2300,N_18441,N_19772);
nand UO_2301 (O_2301,N_19932,N_19163);
or UO_2302 (O_2302,N_19323,N_18892);
xnor UO_2303 (O_2303,N_19904,N_19592);
nand UO_2304 (O_2304,N_19336,N_18993);
nand UO_2305 (O_2305,N_18562,N_19991);
nor UO_2306 (O_2306,N_19471,N_19081);
and UO_2307 (O_2307,N_19653,N_19204);
nand UO_2308 (O_2308,N_18207,N_18155);
or UO_2309 (O_2309,N_18474,N_18447);
or UO_2310 (O_2310,N_19402,N_18904);
or UO_2311 (O_2311,N_19427,N_18893);
or UO_2312 (O_2312,N_19225,N_19062);
nor UO_2313 (O_2313,N_19922,N_18656);
nand UO_2314 (O_2314,N_19611,N_18222);
nor UO_2315 (O_2315,N_19807,N_19037);
xor UO_2316 (O_2316,N_18770,N_18323);
nand UO_2317 (O_2317,N_18907,N_19429);
xnor UO_2318 (O_2318,N_19581,N_19912);
nand UO_2319 (O_2319,N_19860,N_19300);
and UO_2320 (O_2320,N_19555,N_18286);
nand UO_2321 (O_2321,N_18145,N_19700);
and UO_2322 (O_2322,N_19395,N_18540);
and UO_2323 (O_2323,N_18856,N_18917);
nand UO_2324 (O_2324,N_18891,N_18931);
nor UO_2325 (O_2325,N_19221,N_18324);
and UO_2326 (O_2326,N_19262,N_19796);
or UO_2327 (O_2327,N_18103,N_18658);
nand UO_2328 (O_2328,N_19614,N_19012);
or UO_2329 (O_2329,N_19055,N_18387);
xor UO_2330 (O_2330,N_18021,N_18077);
or UO_2331 (O_2331,N_19978,N_18208);
nand UO_2332 (O_2332,N_18744,N_18624);
xnor UO_2333 (O_2333,N_19873,N_19229);
nand UO_2334 (O_2334,N_18017,N_19770);
or UO_2335 (O_2335,N_18118,N_19063);
and UO_2336 (O_2336,N_18030,N_18924);
xnor UO_2337 (O_2337,N_18995,N_18010);
nand UO_2338 (O_2338,N_19008,N_18064);
nor UO_2339 (O_2339,N_19837,N_18637);
or UO_2340 (O_2340,N_18332,N_19013);
or UO_2341 (O_2341,N_18531,N_18738);
nor UO_2342 (O_2342,N_19137,N_18457);
and UO_2343 (O_2343,N_18783,N_18617);
nand UO_2344 (O_2344,N_19731,N_19319);
xnor UO_2345 (O_2345,N_19982,N_18186);
xnor UO_2346 (O_2346,N_18840,N_18484);
or UO_2347 (O_2347,N_19777,N_19892);
nor UO_2348 (O_2348,N_19650,N_19041);
xnor UO_2349 (O_2349,N_18638,N_18840);
nor UO_2350 (O_2350,N_19686,N_19500);
nor UO_2351 (O_2351,N_19811,N_19951);
xnor UO_2352 (O_2352,N_19140,N_18526);
nand UO_2353 (O_2353,N_18126,N_18383);
or UO_2354 (O_2354,N_18550,N_19493);
nor UO_2355 (O_2355,N_18477,N_19742);
and UO_2356 (O_2356,N_18660,N_19259);
and UO_2357 (O_2357,N_19916,N_18235);
nor UO_2358 (O_2358,N_19595,N_19016);
nand UO_2359 (O_2359,N_18930,N_19414);
nand UO_2360 (O_2360,N_18061,N_19858);
nor UO_2361 (O_2361,N_19901,N_18836);
or UO_2362 (O_2362,N_19315,N_18880);
nand UO_2363 (O_2363,N_19672,N_19191);
and UO_2364 (O_2364,N_18016,N_18403);
nand UO_2365 (O_2365,N_18128,N_19324);
and UO_2366 (O_2366,N_18982,N_18417);
nor UO_2367 (O_2367,N_18906,N_19944);
nor UO_2368 (O_2368,N_19661,N_19734);
and UO_2369 (O_2369,N_19472,N_19971);
nor UO_2370 (O_2370,N_19390,N_19120);
nor UO_2371 (O_2371,N_18934,N_19019);
or UO_2372 (O_2372,N_18179,N_18566);
or UO_2373 (O_2373,N_18675,N_19857);
nor UO_2374 (O_2374,N_19894,N_19013);
and UO_2375 (O_2375,N_19540,N_19180);
nand UO_2376 (O_2376,N_19827,N_19647);
xnor UO_2377 (O_2377,N_19278,N_19044);
nor UO_2378 (O_2378,N_18627,N_19318);
nor UO_2379 (O_2379,N_19539,N_18032);
or UO_2380 (O_2380,N_18112,N_19381);
and UO_2381 (O_2381,N_19611,N_19521);
and UO_2382 (O_2382,N_18574,N_18205);
nand UO_2383 (O_2383,N_19872,N_19628);
and UO_2384 (O_2384,N_19757,N_18208);
nand UO_2385 (O_2385,N_19134,N_19608);
and UO_2386 (O_2386,N_18494,N_19331);
nand UO_2387 (O_2387,N_19371,N_19885);
or UO_2388 (O_2388,N_18276,N_18015);
xor UO_2389 (O_2389,N_18803,N_18327);
nand UO_2390 (O_2390,N_18681,N_18740);
nand UO_2391 (O_2391,N_19166,N_18894);
nor UO_2392 (O_2392,N_18292,N_18616);
nor UO_2393 (O_2393,N_18329,N_19579);
and UO_2394 (O_2394,N_19720,N_18888);
xor UO_2395 (O_2395,N_18741,N_19337);
and UO_2396 (O_2396,N_18414,N_19654);
or UO_2397 (O_2397,N_18490,N_19722);
and UO_2398 (O_2398,N_19468,N_19242);
xnor UO_2399 (O_2399,N_18616,N_19673);
or UO_2400 (O_2400,N_19564,N_18904);
nand UO_2401 (O_2401,N_18938,N_19118);
nand UO_2402 (O_2402,N_18183,N_19810);
xor UO_2403 (O_2403,N_19033,N_18367);
nand UO_2404 (O_2404,N_19516,N_18258);
or UO_2405 (O_2405,N_19192,N_19106);
nor UO_2406 (O_2406,N_18800,N_19168);
nor UO_2407 (O_2407,N_19268,N_19375);
and UO_2408 (O_2408,N_18509,N_18188);
or UO_2409 (O_2409,N_18816,N_19067);
or UO_2410 (O_2410,N_18154,N_19781);
nand UO_2411 (O_2411,N_19165,N_18259);
xor UO_2412 (O_2412,N_18380,N_18643);
nor UO_2413 (O_2413,N_18211,N_18361);
and UO_2414 (O_2414,N_19138,N_18306);
nor UO_2415 (O_2415,N_19627,N_18117);
xor UO_2416 (O_2416,N_19142,N_18216);
nand UO_2417 (O_2417,N_18887,N_19530);
or UO_2418 (O_2418,N_19168,N_18905);
and UO_2419 (O_2419,N_19676,N_18072);
xor UO_2420 (O_2420,N_18231,N_19179);
xor UO_2421 (O_2421,N_19335,N_19218);
nand UO_2422 (O_2422,N_19310,N_19215);
nor UO_2423 (O_2423,N_18068,N_18923);
nor UO_2424 (O_2424,N_18819,N_19887);
nor UO_2425 (O_2425,N_19989,N_19847);
and UO_2426 (O_2426,N_18434,N_18281);
xnor UO_2427 (O_2427,N_19596,N_19237);
nor UO_2428 (O_2428,N_19137,N_19438);
nor UO_2429 (O_2429,N_19969,N_18162);
nor UO_2430 (O_2430,N_18923,N_19526);
xor UO_2431 (O_2431,N_18027,N_19750);
nor UO_2432 (O_2432,N_18391,N_18557);
and UO_2433 (O_2433,N_18719,N_19512);
nor UO_2434 (O_2434,N_18048,N_18404);
xnor UO_2435 (O_2435,N_18161,N_18215);
nand UO_2436 (O_2436,N_18698,N_19468);
and UO_2437 (O_2437,N_19674,N_19848);
or UO_2438 (O_2438,N_19014,N_19333);
nand UO_2439 (O_2439,N_18465,N_18117);
and UO_2440 (O_2440,N_18584,N_18230);
nor UO_2441 (O_2441,N_18966,N_19563);
nor UO_2442 (O_2442,N_19510,N_18538);
nand UO_2443 (O_2443,N_19334,N_18558);
or UO_2444 (O_2444,N_19449,N_19946);
nor UO_2445 (O_2445,N_19909,N_18341);
and UO_2446 (O_2446,N_19672,N_18799);
and UO_2447 (O_2447,N_18821,N_18473);
xor UO_2448 (O_2448,N_19123,N_19812);
and UO_2449 (O_2449,N_18998,N_19374);
or UO_2450 (O_2450,N_18481,N_19149);
or UO_2451 (O_2451,N_18395,N_19770);
or UO_2452 (O_2452,N_19522,N_19500);
and UO_2453 (O_2453,N_18051,N_18907);
xnor UO_2454 (O_2454,N_18924,N_19807);
or UO_2455 (O_2455,N_19304,N_18015);
and UO_2456 (O_2456,N_18022,N_18408);
nand UO_2457 (O_2457,N_19823,N_18595);
nor UO_2458 (O_2458,N_19027,N_19806);
xor UO_2459 (O_2459,N_19381,N_18453);
nand UO_2460 (O_2460,N_18685,N_18002);
nor UO_2461 (O_2461,N_19331,N_18667);
or UO_2462 (O_2462,N_19466,N_19851);
xnor UO_2463 (O_2463,N_19675,N_18053);
and UO_2464 (O_2464,N_19127,N_18834);
nor UO_2465 (O_2465,N_19736,N_19616);
or UO_2466 (O_2466,N_19245,N_19098);
nor UO_2467 (O_2467,N_19769,N_19131);
and UO_2468 (O_2468,N_18148,N_18334);
xor UO_2469 (O_2469,N_18891,N_18537);
nand UO_2470 (O_2470,N_19714,N_18008);
xnor UO_2471 (O_2471,N_18981,N_19684);
xnor UO_2472 (O_2472,N_19384,N_19130);
xor UO_2473 (O_2473,N_19389,N_18807);
or UO_2474 (O_2474,N_18369,N_19849);
nor UO_2475 (O_2475,N_18198,N_18358);
or UO_2476 (O_2476,N_18258,N_19373);
and UO_2477 (O_2477,N_18902,N_19631);
nand UO_2478 (O_2478,N_18254,N_18727);
or UO_2479 (O_2479,N_18365,N_19063);
or UO_2480 (O_2480,N_19679,N_18149);
nor UO_2481 (O_2481,N_18398,N_19882);
nor UO_2482 (O_2482,N_19435,N_18373);
or UO_2483 (O_2483,N_18322,N_18756);
or UO_2484 (O_2484,N_19709,N_19471);
nor UO_2485 (O_2485,N_18115,N_19809);
nor UO_2486 (O_2486,N_19551,N_18362);
xor UO_2487 (O_2487,N_18094,N_18393);
xor UO_2488 (O_2488,N_19485,N_19657);
xor UO_2489 (O_2489,N_19355,N_19865);
or UO_2490 (O_2490,N_19048,N_18160);
nand UO_2491 (O_2491,N_19958,N_18729);
nand UO_2492 (O_2492,N_19509,N_19804);
or UO_2493 (O_2493,N_19672,N_18333);
nand UO_2494 (O_2494,N_18931,N_18804);
nand UO_2495 (O_2495,N_18616,N_19880);
or UO_2496 (O_2496,N_18187,N_19345);
and UO_2497 (O_2497,N_18858,N_19582);
or UO_2498 (O_2498,N_19014,N_19168);
xnor UO_2499 (O_2499,N_19015,N_18911);
endmodule